module min_hash(
  input wire [319:0] set1,
  input wire [319:0] set2,
  output wire [655:0] out
);
  // lint_off MULTIPLY
  function automatic [21:0] umul22b_16b_x_6b (input reg [15:0] lhs, input reg [5:0] rhs);
    begin
      umul22b_16b_x_6b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  // lint_off MULTIPLY
  function automatic [22:0] umul23b_16b_x_7b (input reg [15:0] lhs, input reg [6:0] rhs);
    begin
      umul23b_16b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [15:0] set1_unflattened[20];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  wire [15:0] set2_unflattened[20];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  wire [15:0] array_index_35223;
  wire [15:0] array_index_35225;
  wire [21:0] umul_35227;
  wire [21:0] umul_35228;
  wire [21:0] umul_35237;
  wire [21:0] umul_35238;
  wire [15:0] array_index_35239;
  wire [15:0] array_index_35243;
  wire [21:0] umul_35251;
  wire [15:0] add_35253;
  wire [21:0] umul_35255;
  wire [15:0] add_35257;
  wire [21:0] umul_35277;
  wire [21:0] umul_35278;
  wire [21:0] umul_35279;
  wire [21:0] add_35281;
  wire [21:0] umul_35283;
  wire [21:0] add_35285;
  wire [15:0] array_index_35287;
  wire [31:0] smod_35291;
  wire [15:0] array_index_35292;
  wire [31:0] smod_35296;
  wire [21:0] umul_35309;
  wire [15:0] add_35311;
  wire [21:0] umul_35315;
  wire [15:0] add_35317;
  wire [31:0] smod_35332;
  wire [31:0] smod_35336;
  wire [22:0] umul_35351;
  wire [22:0] umul_35352;
  wire [21:0] umul_35353;
  wire [20:0] add_35355;
  wire [21:0] umul_35357;
  wire [20:0] add_35359;
  wire [21:0] umul_35361;
  wire [21:0] add_35363;
  wire [21:0] umul_35367;
  wire [21:0] add_35369;
  wire [15:0] array_index_35373;
  wire [31:0] smod_35377;
  wire [15:0] array_index_35380;
  wire [31:0] smod_35384;
  wire [21:0] umul_35411;
  wire [15:0] add_35413;
  wire [15:0] sel_35418;
  wire [21:0] umul_35419;
  wire [15:0] add_35421;
  wire [15:0] sel_35426;
  wire [31:0] smod_35438;
  wire [31:0] smod_35442;
  wire [31:0] smod_35446;
  wire [31:0] smod_35452;
  wire [22:0] umul_35469;
  wire [22:0] umul_35470;
  wire [22:0] umul_35471;
  wire [22:0] add_35473;
  wire [22:0] umul_35475;
  wire [22:0] add_35477;
  wire [21:0] umul_35479;
  wire [20:0] add_35481;
  wire [21:0] umul_35485;
  wire [20:0] add_35487;
  wire [21:0] umul_35491;
  wire [21:0] add_35493;
  wire [15:0] sel_35498;
  wire [21:0] umul_35499;
  wire [21:0] add_35501;
  wire [15:0] sel_35506;
  wire [15:0] array_index_35507;
  wire [31:0] smod_35511;
  wire [15:0] array_index_35513;
  wire [31:0] smod_35517;
  wire [21:0] umul_35555;
  wire [15:0] add_35557;
  wire [15:0] sel_35562;
  wire [21:0] umul_35563;
  wire [15:0] add_35565;
  wire [15:0] sel_35570;
  wire [31:0] smod_35580;
  wire [31:0] smod_35584;
  wire [31:0] smod_35588;
  wire [31:0] smod_35594;
  wire [31:0] smod_35600;
  wire [31:0] smod_35605;
  wire [22:0] umul_35621;
  wire [20:0] add_35623;
  wire [22:0] umul_35625;
  wire [20:0] add_35627;
  wire [22:0] umul_35629;
  wire [22:0] add_35631;
  wire [22:0] umul_35635;
  wire [22:0] add_35637;
  wire [21:0] umul_35641;
  wire [20:0] add_35643;
  wire [15:0] sel_35648;
  wire [21:0] umul_35649;
  wire [20:0] add_35651;
  wire [15:0] sel_35656;
  wire [21:0] umul_35657;
  wire [21:0] add_35659;
  wire [15:0] sel_35664;
  wire [21:0] umul_35665;
  wire [21:0] add_35667;
  wire [15:0] sel_35672;
  wire [15:0] array_index_35673;
  wire [31:0] smod_35677;
  wire [15:0] array_index_35679;
  wire [31:0] smod_35683;
  wire [21:0] umul_35729;
  wire [15:0] add_35731;
  wire [15:0] sel_35736;
  wire [21:0] umul_35737;
  wire [15:0] add_35739;
  wire [15:0] sel_35744;
  wire [31:0] smod_35748;
  wire [31:0] smod_35752;
  wire [31:0] smod_35756;
  wire [31:0] smod_35762;
  wire [31:0] smod_35768;
  wire [31:0] smod_35773;
  wire [31:0] smod_35778;
  wire [31:0] smod_35783;
  wire [22:0] umul_35799;
  wire [20:0] add_35801;
  wire [22:0] umul_35805;
  wire [20:0] add_35807;
  wire [22:0] umul_35811;
  wire [22:0] add_35813;
  wire [15:0] sel_35818;
  wire [22:0] umul_35819;
  wire [22:0] add_35821;
  wire [15:0] sel_35826;
  wire [21:0] umul_35827;
  wire [20:0] add_35829;
  wire [15:0] sel_35834;
  wire [21:0] umul_35835;
  wire [20:0] add_35837;
  wire [15:0] sel_35842;
  wire [21:0] umul_35843;
  wire [21:0] add_35845;
  wire [15:0] sel_35850;
  wire [21:0] umul_35851;
  wire [21:0] add_35853;
  wire [15:0] sel_35858;
  wire [15:0] array_index_35859;
  wire [31:0] smod_35863;
  wire [15:0] array_index_35865;
  wire [31:0] smod_35869;
  wire [21:0] umul_35919;
  wire [15:0] add_35921;
  wire [15:0] sel_35926;
  wire [21:0] umul_35927;
  wire [15:0] add_35929;
  wire [15:0] sel_35934;
  wire [31:0] smod_35938;
  wire [31:0] smod_35944;
  wire [31:0] smod_35950;
  wire [31:0] smod_35955;
  wire [31:0] smod_35960;
  wire [31:0] smod_35965;
  wire [31:0] smod_35970;
  wire [31:0] smod_35975;
  wire [22:0] umul_35991;
  wire [20:0] add_35993;
  wire [15:0] sel_35998;
  wire [22:0] umul_35999;
  wire [20:0] add_36001;
  wire [15:0] sel_36006;
  wire [22:0] umul_36007;
  wire [22:0] add_36009;
  wire [15:0] sel_36014;
  wire [22:0] umul_36015;
  wire [22:0] add_36017;
  wire [15:0] sel_36022;
  wire [21:0] umul_36023;
  wire [20:0] add_36025;
  wire [15:0] sel_36030;
  wire [21:0] umul_36031;
  wire [20:0] add_36033;
  wire [15:0] sel_36038;
  wire [21:0] umul_36039;
  wire [21:0] add_36041;
  wire [15:0] sel_36046;
  wire [21:0] umul_36047;
  wire [21:0] add_36049;
  wire [15:0] sel_36054;
  wire [15:0] array_index_36055;
  wire [31:0] smod_36059;
  wire [15:0] array_index_36061;
  wire [31:0] smod_36065;
  wire [21:0] umul_36115;
  wire [15:0] add_36117;
  wire [15:0] sel_36122;
  wire [21:0] umul_36123;
  wire [15:0] add_36125;
  wire [15:0] sel_36130;
  wire [31:0] smod_36134;
  wire [31:0] smod_36139;
  wire [31:0] smod_36144;
  wire [31:0] smod_36149;
  wire [31:0] smod_36154;
  wire [31:0] smod_36159;
  wire [31:0] smod_36164;
  wire [31:0] smod_36169;
  wire [22:0] umul_36185;
  wire [20:0] add_36187;
  wire [15:0] sel_36192;
  wire [22:0] umul_36193;
  wire [20:0] add_36195;
  wire [15:0] sel_36200;
  wire [22:0] umul_36201;
  wire [22:0] add_36203;
  wire [15:0] sel_36208;
  wire [22:0] umul_36209;
  wire [22:0] add_36211;
  wire [15:0] sel_36216;
  wire [21:0] umul_36217;
  wire [20:0] add_36219;
  wire [15:0] sel_36224;
  wire [21:0] umul_36225;
  wire [20:0] add_36227;
  wire [15:0] sel_36232;
  wire [21:0] umul_36233;
  wire [21:0] add_36235;
  wire [15:0] sel_36240;
  wire [21:0] umul_36241;
  wire [21:0] add_36243;
  wire [15:0] sel_36248;
  wire [15:0] array_index_36249;
  wire [31:0] smod_36253;
  wire [15:0] array_index_36255;
  wire [31:0] smod_36259;
  wire [21:0] umul_36309;
  wire [15:0] add_36311;
  wire [15:0] sel_36316;
  wire [21:0] umul_36317;
  wire [15:0] add_36319;
  wire [15:0] sel_36324;
  wire [31:0] smod_36328;
  wire [31:0] smod_36333;
  wire [31:0] smod_36338;
  wire [31:0] smod_36343;
  wire [31:0] smod_36348;
  wire [31:0] smod_36353;
  wire [31:0] smod_36358;
  wire [31:0] smod_36363;
  wire [22:0] umul_36379;
  wire [20:0] add_36381;
  wire [15:0] sel_36386;
  wire [22:0] umul_36387;
  wire [20:0] add_36389;
  wire [15:0] sel_36394;
  wire [22:0] umul_36395;
  wire [22:0] add_36397;
  wire [15:0] sel_36402;
  wire [22:0] umul_36403;
  wire [22:0] add_36405;
  wire [15:0] sel_36410;
  wire [21:0] umul_36411;
  wire [20:0] add_36413;
  wire [15:0] sel_36418;
  wire [21:0] umul_36419;
  wire [20:0] add_36421;
  wire [15:0] sel_36426;
  wire [21:0] umul_36427;
  wire [21:0] add_36429;
  wire [15:0] sel_36434;
  wire [21:0] umul_36435;
  wire [21:0] add_36437;
  wire [15:0] sel_36442;
  wire [15:0] array_index_36443;
  wire [31:0] smod_36447;
  wire [15:0] array_index_36449;
  wire [31:0] smod_36453;
  wire [21:0] umul_36503;
  wire [15:0] add_36505;
  wire [15:0] sel_36510;
  wire [21:0] umul_36511;
  wire [15:0] add_36513;
  wire [15:0] sel_36518;
  wire [31:0] smod_36522;
  wire [31:0] smod_36527;
  wire [31:0] smod_36532;
  wire [31:0] smod_36537;
  wire [31:0] smod_36542;
  wire [31:0] smod_36547;
  wire [31:0] smod_36552;
  wire [31:0] smod_36557;
  wire [22:0] umul_36573;
  wire [20:0] add_36575;
  wire [15:0] sel_36580;
  wire [22:0] umul_36581;
  wire [20:0] add_36583;
  wire [15:0] sel_36588;
  wire [22:0] umul_36589;
  wire [22:0] add_36591;
  wire [15:0] sel_36596;
  wire [22:0] umul_36597;
  wire [22:0] add_36599;
  wire [15:0] sel_36604;
  wire [21:0] umul_36605;
  wire [20:0] add_36607;
  wire [15:0] sel_36612;
  wire [21:0] umul_36613;
  wire [20:0] add_36615;
  wire [15:0] sel_36620;
  wire [21:0] umul_36621;
  wire [21:0] add_36623;
  wire [15:0] sel_36628;
  wire [21:0] umul_36629;
  wire [21:0] add_36631;
  wire [15:0] sel_36636;
  wire [15:0] array_index_36637;
  wire [31:0] smod_36641;
  wire [15:0] array_index_36643;
  wire [31:0] smod_36647;
  wire [21:0] umul_36697;
  wire [15:0] add_36699;
  wire [15:0] sel_36704;
  wire [21:0] umul_36705;
  wire [15:0] add_36707;
  wire [15:0] sel_36712;
  wire [31:0] smod_36716;
  wire [31:0] smod_36721;
  wire [31:0] smod_36726;
  wire [31:0] smod_36731;
  wire [31:0] smod_36736;
  wire [31:0] smod_36741;
  wire [31:0] smod_36746;
  wire [31:0] smod_36751;
  wire [22:0] umul_36767;
  wire [20:0] add_36769;
  wire [15:0] sel_36774;
  wire [22:0] umul_36775;
  wire [20:0] add_36777;
  wire [15:0] sel_36782;
  wire [22:0] umul_36783;
  wire [22:0] add_36785;
  wire [15:0] sel_36790;
  wire [22:0] umul_36791;
  wire [22:0] add_36793;
  wire [15:0] sel_36798;
  wire [21:0] umul_36799;
  wire [20:0] add_36801;
  wire [15:0] sel_36806;
  wire [21:0] umul_36807;
  wire [20:0] add_36809;
  wire [15:0] sel_36814;
  wire [21:0] umul_36815;
  wire [21:0] add_36817;
  wire [15:0] sel_36822;
  wire [21:0] umul_36823;
  wire [21:0] add_36825;
  wire [15:0] sel_36830;
  wire [15:0] array_index_36831;
  wire [31:0] smod_36835;
  wire [15:0] array_index_36837;
  wire [31:0] smod_36841;
  wire [21:0] umul_36891;
  wire [15:0] add_36893;
  wire [15:0] sel_36898;
  wire [21:0] umul_36899;
  wire [15:0] add_36901;
  wire [15:0] sel_36906;
  wire [31:0] smod_36910;
  wire [31:0] smod_36915;
  wire [31:0] smod_36920;
  wire [31:0] smod_36925;
  wire [31:0] smod_36930;
  wire [31:0] smod_36935;
  wire [31:0] smod_36940;
  wire [31:0] smod_36945;
  wire [22:0] umul_36961;
  wire [20:0] add_36963;
  wire [15:0] sel_36968;
  wire [22:0] umul_36969;
  wire [20:0] add_36971;
  wire [15:0] sel_36976;
  wire [22:0] umul_36977;
  wire [22:0] add_36979;
  wire [15:0] sel_36984;
  wire [22:0] umul_36985;
  wire [22:0] add_36987;
  wire [15:0] sel_36992;
  wire [21:0] umul_36993;
  wire [20:0] add_36995;
  wire [15:0] sel_37000;
  wire [21:0] umul_37001;
  wire [20:0] add_37003;
  wire [15:0] sel_37008;
  wire [21:0] umul_37009;
  wire [21:0] add_37011;
  wire [15:0] sel_37016;
  wire [21:0] umul_37017;
  wire [21:0] add_37019;
  wire [15:0] sel_37024;
  wire [15:0] array_index_37025;
  wire [31:0] smod_37029;
  wire [15:0] array_index_37031;
  wire [31:0] smod_37035;
  wire [21:0] umul_37085;
  wire [15:0] add_37087;
  wire [15:0] sel_37092;
  wire [21:0] umul_37093;
  wire [15:0] add_37095;
  wire [15:0] sel_37100;
  wire [31:0] smod_37104;
  wire [31:0] smod_37109;
  wire [31:0] smod_37114;
  wire [31:0] smod_37119;
  wire [31:0] smod_37124;
  wire [31:0] smod_37129;
  wire [31:0] smod_37134;
  wire [31:0] smod_37139;
  wire [22:0] umul_37155;
  wire [20:0] add_37157;
  wire [15:0] sel_37162;
  wire [22:0] umul_37163;
  wire [20:0] add_37165;
  wire [15:0] sel_37170;
  wire [22:0] umul_37171;
  wire [22:0] add_37173;
  wire [15:0] sel_37178;
  wire [22:0] umul_37179;
  wire [22:0] add_37181;
  wire [15:0] sel_37186;
  wire [21:0] umul_37187;
  wire [20:0] add_37189;
  wire [15:0] sel_37194;
  wire [21:0] umul_37195;
  wire [20:0] add_37197;
  wire [15:0] sel_37202;
  wire [21:0] umul_37203;
  wire [21:0] add_37205;
  wire [15:0] sel_37210;
  wire [21:0] umul_37211;
  wire [21:0] add_37213;
  wire [15:0] sel_37218;
  wire [15:0] array_index_37219;
  wire [31:0] smod_37223;
  wire [15:0] array_index_37225;
  wire [31:0] smod_37229;
  wire [21:0] umul_37279;
  wire [15:0] add_37281;
  wire [15:0] sel_37286;
  wire [21:0] umul_37287;
  wire [15:0] add_37289;
  wire [15:0] sel_37294;
  wire [31:0] smod_37298;
  wire [31:0] smod_37303;
  wire [31:0] smod_37308;
  wire [31:0] smod_37313;
  wire [31:0] smod_37318;
  wire [31:0] smod_37323;
  wire [31:0] smod_37328;
  wire [31:0] smod_37333;
  wire [22:0] umul_37349;
  wire [20:0] add_37351;
  wire [15:0] sel_37356;
  wire [22:0] umul_37357;
  wire [20:0] add_37359;
  wire [15:0] sel_37364;
  wire [22:0] umul_37365;
  wire [22:0] add_37367;
  wire [15:0] sel_37372;
  wire [22:0] umul_37373;
  wire [22:0] add_37375;
  wire [15:0] sel_37380;
  wire [21:0] umul_37381;
  wire [20:0] add_37383;
  wire [15:0] sel_37388;
  wire [21:0] umul_37389;
  wire [20:0] add_37391;
  wire [15:0] sel_37396;
  wire [21:0] umul_37397;
  wire [21:0] add_37399;
  wire [15:0] sel_37404;
  wire [21:0] umul_37405;
  wire [21:0] add_37407;
  wire [15:0] sel_37412;
  wire [15:0] array_index_37413;
  wire [31:0] smod_37417;
  wire [15:0] array_index_37419;
  wire [31:0] smod_37423;
  wire [21:0] umul_37473;
  wire [15:0] add_37475;
  wire [15:0] sel_37480;
  wire [21:0] umul_37481;
  wire [15:0] add_37483;
  wire [15:0] sel_37488;
  wire [31:0] smod_37492;
  wire [31:0] smod_37497;
  wire [31:0] smod_37502;
  wire [31:0] smod_37507;
  wire [31:0] smod_37512;
  wire [31:0] smod_37517;
  wire [31:0] smod_37522;
  wire [31:0] smod_37527;
  wire [22:0] umul_37543;
  wire [20:0] add_37545;
  wire [15:0] sel_37550;
  wire [22:0] umul_37551;
  wire [20:0] add_37553;
  wire [15:0] sel_37558;
  wire [22:0] umul_37559;
  wire [22:0] add_37561;
  wire [15:0] sel_37566;
  wire [22:0] umul_37567;
  wire [22:0] add_37569;
  wire [15:0] sel_37574;
  wire [21:0] umul_37575;
  wire [20:0] add_37577;
  wire [15:0] sel_37582;
  wire [21:0] umul_37583;
  wire [20:0] add_37585;
  wire [15:0] sel_37590;
  wire [21:0] umul_37591;
  wire [21:0] add_37593;
  wire [15:0] sel_37598;
  wire [21:0] umul_37599;
  wire [21:0] add_37601;
  wire [15:0] sel_37606;
  wire [15:0] array_index_37607;
  wire [31:0] smod_37611;
  wire [15:0] array_index_37613;
  wire [31:0] smod_37617;
  wire [21:0] umul_37667;
  wire [15:0] add_37669;
  wire [15:0] sel_37674;
  wire [21:0] umul_37675;
  wire [15:0] add_37677;
  wire [15:0] sel_37682;
  wire [31:0] smod_37686;
  wire [31:0] smod_37691;
  wire [31:0] smod_37696;
  wire [31:0] smod_37701;
  wire [31:0] smod_37706;
  wire [31:0] smod_37711;
  wire [31:0] smod_37716;
  wire [31:0] smod_37721;
  wire [22:0] umul_37737;
  wire [20:0] add_37739;
  wire [15:0] sel_37744;
  wire [22:0] umul_37745;
  wire [20:0] add_37747;
  wire [15:0] sel_37752;
  wire [22:0] umul_37753;
  wire [22:0] add_37755;
  wire [15:0] sel_37760;
  wire [22:0] umul_37761;
  wire [22:0] add_37763;
  wire [15:0] sel_37768;
  wire [21:0] umul_37769;
  wire [20:0] add_37771;
  wire [15:0] sel_37776;
  wire [21:0] umul_37777;
  wire [20:0] add_37779;
  wire [15:0] sel_37784;
  wire [21:0] umul_37785;
  wire [21:0] add_37787;
  wire [15:0] sel_37792;
  wire [21:0] umul_37793;
  wire [21:0] add_37795;
  wire [15:0] sel_37800;
  wire [15:0] array_index_37801;
  wire [31:0] smod_37805;
  wire [15:0] array_index_37807;
  wire [31:0] smod_37811;
  wire [21:0] umul_37861;
  wire [15:0] add_37863;
  wire [15:0] sel_37868;
  wire [21:0] umul_37869;
  wire [15:0] add_37871;
  wire [15:0] sel_37876;
  wire [31:0] smod_37880;
  wire [31:0] smod_37885;
  wire [31:0] smod_37890;
  wire [31:0] smod_37895;
  wire [31:0] smod_37900;
  wire [31:0] smod_37905;
  wire [31:0] smod_37910;
  wire [31:0] smod_37915;
  wire [22:0] umul_37931;
  wire [20:0] add_37933;
  wire [15:0] sel_37938;
  wire [22:0] umul_37939;
  wire [20:0] add_37941;
  wire [15:0] sel_37946;
  wire [22:0] umul_37947;
  wire [22:0] add_37949;
  wire [15:0] sel_37954;
  wire [22:0] umul_37955;
  wire [22:0] add_37957;
  wire [15:0] sel_37962;
  wire [21:0] umul_37963;
  wire [20:0] add_37965;
  wire [15:0] sel_37970;
  wire [21:0] umul_37971;
  wire [20:0] add_37973;
  wire [15:0] sel_37978;
  wire [21:0] umul_37979;
  wire [21:0] add_37981;
  wire [15:0] sel_37986;
  wire [21:0] umul_37987;
  wire [21:0] add_37989;
  wire [15:0] sel_37994;
  wire [15:0] array_index_37995;
  wire [31:0] smod_37999;
  wire [15:0] array_index_38001;
  wire [31:0] smod_38005;
  wire [21:0] umul_38055;
  wire [15:0] add_38057;
  wire [15:0] sel_38062;
  wire [21:0] umul_38063;
  wire [15:0] add_38065;
  wire [15:0] sel_38070;
  wire [31:0] smod_38074;
  wire [31:0] smod_38079;
  wire [31:0] smod_38084;
  wire [31:0] smod_38089;
  wire [31:0] smod_38094;
  wire [31:0] smod_38099;
  wire [31:0] smod_38104;
  wire [31:0] smod_38109;
  wire [22:0] umul_38125;
  wire [20:0] add_38127;
  wire [15:0] sel_38132;
  wire [22:0] umul_38133;
  wire [20:0] add_38135;
  wire [15:0] sel_38140;
  wire [22:0] umul_38141;
  wire [22:0] add_38143;
  wire [15:0] sel_38148;
  wire [22:0] umul_38149;
  wire [22:0] add_38151;
  wire [15:0] sel_38156;
  wire [21:0] umul_38157;
  wire [20:0] add_38159;
  wire [15:0] sel_38164;
  wire [21:0] umul_38165;
  wire [20:0] add_38167;
  wire [15:0] sel_38172;
  wire [21:0] umul_38173;
  wire [21:0] add_38175;
  wire [15:0] sel_38180;
  wire [21:0] umul_38181;
  wire [21:0] add_38183;
  wire [15:0] sel_38188;
  wire [15:0] array_index_38189;
  wire [31:0] smod_38193;
  wire [15:0] array_index_38195;
  wire [31:0] smod_38199;
  wire [21:0] umul_38249;
  wire [15:0] add_38251;
  wire [15:0] sel_38256;
  wire [21:0] umul_38257;
  wire [15:0] add_38259;
  wire [15:0] sel_38264;
  wire [31:0] smod_38268;
  wire [31:0] smod_38273;
  wire [31:0] smod_38278;
  wire [31:0] smod_38283;
  wire [31:0] smod_38288;
  wire [31:0] smod_38293;
  wire [31:0] smod_38298;
  wire [31:0] smod_38303;
  wire [22:0] umul_38319;
  wire [20:0] add_38321;
  wire [15:0] sel_38326;
  wire [22:0] umul_38327;
  wire [20:0] add_38329;
  wire [15:0] sel_38334;
  wire [22:0] umul_38335;
  wire [22:0] add_38337;
  wire [15:0] sel_38342;
  wire [22:0] umul_38343;
  wire [22:0] add_38345;
  wire [15:0] sel_38350;
  wire [21:0] umul_38351;
  wire [20:0] add_38353;
  wire [15:0] sel_38358;
  wire [21:0] umul_38359;
  wire [20:0] add_38361;
  wire [15:0] sel_38366;
  wire [21:0] umul_38367;
  wire [21:0] add_38369;
  wire [15:0] sel_38374;
  wire [21:0] umul_38375;
  wire [21:0] add_38377;
  wire [15:0] sel_38382;
  wire [15:0] array_index_38383;
  wire [31:0] smod_38387;
  wire [15:0] array_index_38389;
  wire [31:0] smod_38393;
  wire [21:0] umul_38443;
  wire [15:0] add_38445;
  wire [15:0] sel_38450;
  wire [21:0] umul_38451;
  wire [15:0] add_38453;
  wire [15:0] sel_38458;
  wire [31:0] smod_38462;
  wire [31:0] smod_38467;
  wire [31:0] smod_38472;
  wire [31:0] smod_38477;
  wire [31:0] smod_38482;
  wire [31:0] smod_38487;
  wire [31:0] smod_38492;
  wire [31:0] smod_38497;
  wire [22:0] umul_38511;
  wire [20:0] add_38513;
  wire [15:0] sel_38518;
  wire [22:0] umul_38519;
  wire [20:0] add_38521;
  wire [15:0] sel_38526;
  wire [22:0] umul_38527;
  wire [22:0] add_38529;
  wire [15:0] sel_38534;
  wire [22:0] umul_38535;
  wire [22:0] add_38537;
  wire [15:0] sel_38542;
  wire [21:0] umul_38543;
  wire [20:0] add_38545;
  wire [15:0] sel_38550;
  wire [21:0] umul_38551;
  wire [20:0] add_38553;
  wire [15:0] sel_38558;
  wire [21:0] umul_38559;
  wire [21:0] add_38561;
  wire [15:0] sel_38566;
  wire [21:0] umul_38567;
  wire [21:0] add_38569;
  wire [15:0] sel_38574;
  wire [31:0] smod_38577;
  wire [31:0] smod_38581;
  wire [15:0] add_38632;
  wire [15:0] sel_38637;
  wire [15:0] add_38639;
  wire [15:0] sel_38644;
  wire [31:0] smod_38648;
  wire [31:0] smod_38653;
  wire [31:0] smod_38658;
  wire [31:0] smod_38663;
  wire [31:0] smod_38668;
  wire [31:0] smod_38673;
  wire [31:0] smod_38677;
  wire [31:0] smod_38681;
  wire [22:0] umul_38691;
  wire [20:0] add_38693;
  wire [15:0] sel_38698;
  wire [22:0] umul_38699;
  wire [20:0] add_38701;
  wire [15:0] sel_38706;
  wire [22:0] umul_38707;
  wire [22:0] add_38709;
  wire [15:0] sel_38714;
  wire [22:0] umul_38715;
  wire [22:0] add_38717;
  wire [15:0] sel_38722;
  wire [21:0] umul_38723;
  wire [20:0] add_38725;
  wire [15:0] sel_38730;
  wire [21:0] umul_38731;
  wire [20:0] add_38733;
  wire [15:0] sel_38738;
  wire [21:0] add_38740;
  wire [15:0] sel_38745;
  wire [21:0] add_38747;
  wire [15:0] sel_38752;
  wire [31:0] smod_38753;
  wire [31:0] smod_38755;
  wire [15:0] sel_38804;
  wire [15:0] sel_38808;
  wire [31:0] smod_38812;
  wire [31:0] smod_38817;
  wire [31:0] smod_38822;
  wire [31:0] smod_38827;
  wire [31:0] smod_38831;
  wire [31:0] smod_38835;
  wire [31:0] smod_38837;
  wire [31:0] smod_38839;
  wire [22:0] umul_38845;
  wire [20:0] add_38847;
  wire [15:0] sel_38852;
  wire [22:0] umul_38853;
  wire [20:0] add_38855;
  wire [15:0] sel_38860;
  wire [22:0] umul_38861;
  wire [22:0] add_38863;
  wire [15:0] sel_38868;
  wire [22:0] umul_38869;
  wire [22:0] add_38871;
  wire [15:0] sel_38876;
  wire [20:0] add_38878;
  wire [15:0] sel_38883;
  wire [20:0] add_38885;
  wire [15:0] sel_38890;
  wire [15:0] sel_38894;
  wire [15:0] sel_38898;
  wire [31:0] smod_38942;
  wire [31:0] smod_38947;
  wire [31:0] smod_38951;
  wire [31:0] smod_38955;
  wire [31:0] smod_38957;
  wire [31:0] smod_38959;
  wire [22:0] umul_38965;
  wire [20:0] add_38967;
  wire [15:0] sel_38972;
  wire [22:0] umul_38973;
  wire [20:0] add_38975;
  wire [15:0] sel_38980;
  wire [22:0] add_38982;
  wire [15:0] sel_38987;
  wire [22:0] add_38989;
  wire [15:0] sel_38994;
  wire [15:0] sel_38998;
  wire [15:0] sel_39002;
  wire [1:0] concat_39005;
  wire [1:0] add_39032;
  wire [31:0] smod_39035;
  wire [31:0] smod_39039;
  wire [31:0] smod_39041;
  wire [31:0] smod_39043;
  wire [20:0] add_39050;
  wire [15:0] sel_39055;
  wire [20:0] add_39057;
  wire [15:0] sel_39062;
  wire [15:0] sel_39066;
  wire [15:0] sel_39070;
  wire [2:0] concat_39073;
  wire [2:0] add_39088;
  wire [31:0] smod_39089;
  wire [31:0] smod_39091;
  wire [15:0] sel_39100;
  wire [15:0] sel_39104;
  wire [3:0] concat_39107;
  wire [3:0] add_39114;
  wire [4:0] concat_39121;
  wire [4:0] add_39124;
  assign array_index_35223 = set1_unflattened[5'h00];
  assign array_index_35225 = set2_unflattened[5'h00];
  assign umul_35227 = umul22b_16b_x_6b(array_index_35223, 6'h35);
  assign umul_35228 = umul22b_16b_x_6b(array_index_35225, 6'h35);
  assign umul_35237 = umul22b_16b_x_6b(array_index_35223, 6'h3b);
  assign umul_35238 = umul22b_16b_x_6b(array_index_35225, 6'h3b);
  assign array_index_35239 = set1_unflattened[5'h01];
  assign array_index_35243 = set2_unflattened[5'h01];
  assign umul_35251 = umul22b_16b_x_6b(array_index_35239, 6'h35);
  assign add_35253 = {1'h0, umul_35227[21:7]} + 16'h007d;
  assign umul_35255 = umul22b_16b_x_6b(array_index_35243, 6'h35);
  assign add_35257 = {1'h0, umul_35228[21:7]} + 16'h007d;
  assign umul_35277 = umul22b_16b_x_6b(array_index_35223, 6'h3d);
  assign umul_35278 = umul22b_16b_x_6b(array_index_35225, 6'h3d);
  assign umul_35279 = umul22b_16b_x_6b(array_index_35239, 6'h3b);
  assign add_35281 = {1'h0, umul_35237[21:1]} + 22'h00_1f59;
  assign umul_35283 = umul22b_16b_x_6b(array_index_35243, 6'h3b);
  assign add_35285 = {1'h0, umul_35238[21:1]} + 22'h00_1f59;
  assign array_index_35287 = set1_unflattened[5'h02];
  assign smod_35291 = $unsigned($signed({9'h000, add_35253, umul_35227[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_35292 = set2_unflattened[5'h02];
  assign smod_35296 = $unsigned($signed({9'h000, add_35257, umul_35228[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_35309 = umul22b_16b_x_6b(array_index_35287, 6'h35);
  assign add_35311 = {1'h0, umul_35251[21:7]} + 16'h007d;
  assign umul_35315 = umul22b_16b_x_6b(array_index_35292, 6'h35);
  assign add_35317 = {1'h0, umul_35255[21:7]} + 16'h007d;
  assign smod_35332 = $unsigned($signed({9'h000, add_35281, umul_35237[0]}) % $signed(32'h0000_3ffd));
  assign smod_35336 = $unsigned($signed({9'h000, add_35285, umul_35238[0]}) % $signed(32'h0000_3ffd));
  assign umul_35351 = umul23b_16b_x_7b(array_index_35223, 7'h47);
  assign umul_35352 = umul23b_16b_x_7b(array_index_35225, 7'h47);
  assign umul_35353 = umul22b_16b_x_6b(array_index_35239, 6'h3d);
  assign add_35355 = {1'h0, umul_35277[21:2]} + 21'h00_0fb9;
  assign umul_35357 = umul22b_16b_x_6b(array_index_35243, 6'h3d);
  assign add_35359 = {1'h0, umul_35278[21:2]} + 21'h00_0fb9;
  assign umul_35361 = umul22b_16b_x_6b(array_index_35287, 6'h3b);
  assign add_35363 = {1'h0, umul_35279[21:1]} + 22'h00_1f59;
  assign umul_35367 = umul22b_16b_x_6b(array_index_35292, 6'h3b);
  assign add_35369 = {1'h0, umul_35283[21:1]} + 22'h00_1f59;
  assign array_index_35373 = set1_unflattened[5'h03];
  assign smod_35377 = $unsigned($signed({9'h000, add_35311, umul_35251[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_35380 = set2_unflattened[5'h03];
  assign smod_35384 = $unsigned($signed({9'h000, add_35317, umul_35255[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_35411 = umul22b_16b_x_6b(array_index_35373, 6'h35);
  assign add_35413 = {1'h0, umul_35309[21:7]} + 16'h007d;
  assign sel_35418 = $signed({1'h0, smod_35291[15:0]}) < $signed(17'h0_3ffd) ? smod_35291[15:0] : 16'h3ffd;
  assign umul_35419 = umul22b_16b_x_6b(array_index_35380, 6'h35);
  assign add_35421 = {1'h0, umul_35315[21:7]} + 16'h007d;
  assign sel_35426 = $signed({1'h0, smod_35296[15:0]}) < $signed(17'h0_3ffd) ? smod_35296[15:0] : 16'h3ffd;
  assign smod_35438 = $unsigned($signed({9'h000, add_35355, umul_35277[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_35442 = $unsigned($signed({9'h000, add_35359, umul_35278[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_35446 = $unsigned($signed({9'h000, add_35363, umul_35279[0]}) % $signed(32'h0000_3ffd));
  assign smod_35452 = $unsigned($signed({9'h000, add_35369, umul_35283[0]}) % $signed(32'h0000_3ffd));
  assign umul_35469 = umul23b_16b_x_7b(array_index_35223, 7'h49);
  assign umul_35470 = umul23b_16b_x_7b(array_index_35225, 7'h49);
  assign umul_35471 = umul23b_16b_x_7b(array_index_35239, 7'h47);
  assign add_35473 = {1'h0, umul_35351[22:1]} + 23'h00_1f8b;
  assign umul_35475 = umul23b_16b_x_7b(array_index_35243, 7'h47);
  assign add_35477 = {1'h0, umul_35352[22:1]} + 23'h00_1f8b;
  assign umul_35479 = umul22b_16b_x_6b(array_index_35287, 6'h3d);
  assign add_35481 = {1'h0, umul_35353[21:2]} + 21'h00_0fb9;
  assign umul_35485 = umul22b_16b_x_6b(array_index_35292, 6'h3d);
  assign add_35487 = {1'h0, umul_35357[21:2]} + 21'h00_0fb9;
  assign umul_35491 = umul22b_16b_x_6b(array_index_35373, 6'h3b);
  assign add_35493 = {1'h0, umul_35361[21:1]} + 22'h00_1f59;
  assign sel_35498 = $signed({1'h0, smod_35332[15:0]}) < $signed(17'h0_3ffd) ? smod_35332[15:0] : 16'h3ffd;
  assign umul_35499 = umul22b_16b_x_6b(array_index_35380, 6'h3b);
  assign add_35501 = {1'h0, umul_35367[21:1]} + 22'h00_1f59;
  assign sel_35506 = $signed({1'h0, smod_35336[15:0]}) < $signed(17'h0_3ffd) ? smod_35336[15:0] : 16'h3ffd;
  assign array_index_35507 = set1_unflattened[5'h04];
  assign smod_35511 = $unsigned($signed({9'h000, add_35413, umul_35309[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_35513 = set2_unflattened[5'h04];
  assign smod_35517 = $unsigned($signed({9'h000, add_35421, umul_35315[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_35555 = umul22b_16b_x_6b(array_index_35507, 6'h35);
  assign add_35557 = {1'h0, umul_35411[21:7]} + 16'h007d;
  assign sel_35562 = $signed({1'h0, smod_35377[15:0]}) < $signed({1'h0, sel_35418}) ? smod_35377[15:0] : sel_35418;
  assign umul_35563 = umul22b_16b_x_6b(array_index_35513, 6'h35);
  assign add_35565 = {1'h0, umul_35419[21:7]} + 16'h007d;
  assign sel_35570 = $signed({1'h0, smod_35384[15:0]}) < $signed({1'h0, sel_35426}) ? smod_35384[15:0] : sel_35426;
  assign smod_35580 = $unsigned($signed({8'h00, add_35473, umul_35351[0]}) % $signed(32'h0000_3ffd));
  assign smod_35584 = $unsigned($signed({8'h00, add_35477, umul_35352[0]}) % $signed(32'h0000_3ffd));
  assign smod_35588 = $unsigned($signed({9'h000, add_35481, umul_35353[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_35594 = $unsigned($signed({9'h000, add_35487, umul_35357[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_35600 = $unsigned($signed({9'h000, add_35493, umul_35361[0]}) % $signed(32'h0000_3ffd));
  assign smod_35605 = $unsigned($signed({9'h000, add_35501, umul_35367[0]}) % $signed(32'h0000_3ffd));
  assign umul_35621 = umul23b_16b_x_7b(array_index_35239, 7'h49);
  assign add_35623 = {1'h0, umul_35469[22:3]} + 21'h00_07e9;
  assign umul_35625 = umul23b_16b_x_7b(array_index_35243, 7'h49);
  assign add_35627 = {1'h0, umul_35470[22:3]} + 21'h00_07e9;
  assign umul_35629 = umul23b_16b_x_7b(array_index_35287, 7'h47);
  assign add_35631 = {1'h0, umul_35471[22:1]} + 23'h00_1f8b;
  assign umul_35635 = umul23b_16b_x_7b(array_index_35292, 7'h47);
  assign add_35637 = {1'h0, umul_35475[22:1]} + 23'h00_1f8b;
  assign umul_35641 = umul22b_16b_x_6b(array_index_35373, 6'h3d);
  assign add_35643 = {1'h0, umul_35479[21:2]} + 21'h00_0fb9;
  assign sel_35648 = $signed({1'h0, smod_35438[15:0]}) < $signed(17'h0_3ffd) ? smod_35438[15:0] : 16'h3ffd;
  assign umul_35649 = umul22b_16b_x_6b(array_index_35380, 6'h3d);
  assign add_35651 = {1'h0, umul_35485[21:2]} + 21'h00_0fb9;
  assign sel_35656 = $signed({1'h0, smod_35442[15:0]}) < $signed(17'h0_3ffd) ? smod_35442[15:0] : 16'h3ffd;
  assign umul_35657 = umul22b_16b_x_6b(array_index_35507, 6'h3b);
  assign add_35659 = {1'h0, umul_35491[21:1]} + 22'h00_1f59;
  assign sel_35664 = $signed({1'h0, smod_35446[15:0]}) < $signed({1'h0, sel_35498}) ? smod_35446[15:0] : sel_35498;
  assign umul_35665 = umul22b_16b_x_6b(array_index_35513, 6'h3b);
  assign add_35667 = {1'h0, umul_35499[21:1]} + 22'h00_1f59;
  assign sel_35672 = $signed({1'h0, smod_35452[15:0]}) < $signed({1'h0, sel_35506}) ? smod_35452[15:0] : sel_35506;
  assign array_index_35673 = set1_unflattened[5'h05];
  assign smod_35677 = $unsigned($signed({9'h000, add_35557, umul_35411[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_35679 = set2_unflattened[5'h05];
  assign smod_35683 = $unsigned($signed({9'h000, add_35565, umul_35419[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_35729 = umul22b_16b_x_6b(array_index_35673, 6'h35);
  assign add_35731 = {1'h0, umul_35555[21:7]} + 16'h007d;
  assign sel_35736 = $signed({1'h0, smod_35511[15:0]}) < $signed({1'h0, sel_35562}) ? smod_35511[15:0] : sel_35562;
  assign umul_35737 = umul22b_16b_x_6b(array_index_35679, 6'h35);
  assign add_35739 = {1'h0, umul_35563[21:7]} + 16'h007d;
  assign sel_35744 = $signed({1'h0, smod_35517[15:0]}) < $signed({1'h0, sel_35570}) ? smod_35517[15:0] : sel_35570;
  assign smod_35748 = $unsigned($signed({8'h00, add_35623, umul_35469[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_35752 = $unsigned($signed({8'h00, add_35627, umul_35470[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_35756 = $unsigned($signed({8'h00, add_35631, umul_35471[0]}) % $signed(32'h0000_3ffd));
  assign smod_35762 = $unsigned($signed({8'h00, add_35637, umul_35475[0]}) % $signed(32'h0000_3ffd));
  assign smod_35768 = $unsigned($signed({9'h000, add_35643, umul_35479[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_35773 = $unsigned($signed({9'h000, add_35651, umul_35485[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_35778 = $unsigned($signed({9'h000, add_35659, umul_35491[0]}) % $signed(32'h0000_3ffd));
  assign smod_35783 = $unsigned($signed({9'h000, add_35667, umul_35499[0]}) % $signed(32'h0000_3ffd));
  assign umul_35799 = umul23b_16b_x_7b(array_index_35287, 7'h49);
  assign add_35801 = {1'h0, umul_35621[22:3]} + 21'h00_07e9;
  assign umul_35805 = umul23b_16b_x_7b(array_index_35292, 7'h49);
  assign add_35807 = {1'h0, umul_35625[22:3]} + 21'h00_07e9;
  assign umul_35811 = umul23b_16b_x_7b(array_index_35373, 7'h47);
  assign add_35813 = {1'h0, umul_35629[22:1]} + 23'h00_1f8b;
  assign sel_35818 = $signed({1'h0, smod_35580[15:0]}) < $signed(17'h0_3ffd) ? smod_35580[15:0] : 16'h3ffd;
  assign umul_35819 = umul23b_16b_x_7b(array_index_35380, 7'h47);
  assign add_35821 = {1'h0, umul_35635[22:1]} + 23'h00_1f8b;
  assign sel_35826 = $signed({1'h0, smod_35584[15:0]}) < $signed(17'h0_3ffd) ? smod_35584[15:0] : 16'h3ffd;
  assign umul_35827 = umul22b_16b_x_6b(array_index_35507, 6'h3d);
  assign add_35829 = {1'h0, umul_35641[21:2]} + 21'h00_0fb9;
  assign sel_35834 = $signed({1'h0, smod_35588[15:0]}) < $signed({1'h0, sel_35648}) ? smod_35588[15:0] : sel_35648;
  assign umul_35835 = umul22b_16b_x_6b(array_index_35513, 6'h3d);
  assign add_35837 = {1'h0, umul_35649[21:2]} + 21'h00_0fb9;
  assign sel_35842 = $signed({1'h0, smod_35594[15:0]}) < $signed({1'h0, sel_35656}) ? smod_35594[15:0] : sel_35656;
  assign umul_35843 = umul22b_16b_x_6b(array_index_35673, 6'h3b);
  assign add_35845 = {1'h0, umul_35657[21:1]} + 22'h00_1f59;
  assign sel_35850 = $signed({1'h0, smod_35600[15:0]}) < $signed({1'h0, sel_35664}) ? smod_35600[15:0] : sel_35664;
  assign umul_35851 = umul22b_16b_x_6b(array_index_35679, 6'h3b);
  assign add_35853 = {1'h0, umul_35665[21:1]} + 22'h00_1f59;
  assign sel_35858 = $signed({1'h0, smod_35605[15:0]}) < $signed({1'h0, sel_35672}) ? smod_35605[15:0] : sel_35672;
  assign array_index_35859 = set1_unflattened[5'h06];
  assign smod_35863 = $unsigned($signed({9'h000, add_35731, umul_35555[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_35865 = set2_unflattened[5'h06];
  assign smod_35869 = $unsigned($signed({9'h000, add_35739, umul_35563[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_35919 = umul22b_16b_x_6b(array_index_35859, 6'h35);
  assign add_35921 = {1'h0, umul_35729[21:7]} + 16'h007d;
  assign sel_35926 = $signed({1'h0, smod_35677[15:0]}) < $signed({1'h0, sel_35736}) ? smod_35677[15:0] : sel_35736;
  assign umul_35927 = umul22b_16b_x_6b(array_index_35865, 6'h35);
  assign add_35929 = {1'h0, umul_35737[21:7]} + 16'h007d;
  assign sel_35934 = $signed({1'h0, smod_35683[15:0]}) < $signed({1'h0, sel_35744}) ? smod_35683[15:0] : sel_35744;
  assign smod_35938 = $unsigned($signed({8'h00, add_35801, umul_35621[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_35944 = $unsigned($signed({8'h00, add_35807, umul_35625[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_35950 = $unsigned($signed({8'h00, add_35813, umul_35629[0]}) % $signed(32'h0000_3ffd));
  assign smod_35955 = $unsigned($signed({8'h00, add_35821, umul_35635[0]}) % $signed(32'h0000_3ffd));
  assign smod_35960 = $unsigned($signed({9'h000, add_35829, umul_35641[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_35965 = $unsigned($signed({9'h000, add_35837, umul_35649[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_35970 = $unsigned($signed({9'h000, add_35845, umul_35657[0]}) % $signed(32'h0000_3ffd));
  assign smod_35975 = $unsigned($signed({9'h000, add_35853, umul_35665[0]}) % $signed(32'h0000_3ffd));
  assign umul_35991 = umul23b_16b_x_7b(array_index_35373, 7'h49);
  assign add_35993 = {1'h0, umul_35799[22:3]} + 21'h00_07e9;
  assign sel_35998 = $signed({1'h0, smod_35748[15:0]}) < $signed(17'h0_3ffd) ? smod_35748[15:0] : 16'h3ffd;
  assign umul_35999 = umul23b_16b_x_7b(array_index_35380, 7'h49);
  assign add_36001 = {1'h0, umul_35805[22:3]} + 21'h00_07e9;
  assign sel_36006 = $signed({1'h0, smod_35752[15:0]}) < $signed(17'h0_3ffd) ? smod_35752[15:0] : 16'h3ffd;
  assign umul_36007 = umul23b_16b_x_7b(array_index_35507, 7'h47);
  assign add_36009 = {1'h0, umul_35811[22:1]} + 23'h00_1f8b;
  assign sel_36014 = $signed({1'h0, smod_35756[15:0]}) < $signed({1'h0, sel_35818}) ? smod_35756[15:0] : sel_35818;
  assign umul_36015 = umul23b_16b_x_7b(array_index_35513, 7'h47);
  assign add_36017 = {1'h0, umul_35819[22:1]} + 23'h00_1f8b;
  assign sel_36022 = $signed({1'h0, smod_35762[15:0]}) < $signed({1'h0, sel_35826}) ? smod_35762[15:0] : sel_35826;
  assign umul_36023 = umul22b_16b_x_6b(array_index_35673, 6'h3d);
  assign add_36025 = {1'h0, umul_35827[21:2]} + 21'h00_0fb9;
  assign sel_36030 = $signed({1'h0, smod_35768[15:0]}) < $signed({1'h0, sel_35834}) ? smod_35768[15:0] : sel_35834;
  assign umul_36031 = umul22b_16b_x_6b(array_index_35679, 6'h3d);
  assign add_36033 = {1'h0, umul_35835[21:2]} + 21'h00_0fb9;
  assign sel_36038 = $signed({1'h0, smod_35773[15:0]}) < $signed({1'h0, sel_35842}) ? smod_35773[15:0] : sel_35842;
  assign umul_36039 = umul22b_16b_x_6b(array_index_35859, 6'h3b);
  assign add_36041 = {1'h0, umul_35843[21:1]} + 22'h00_1f59;
  assign sel_36046 = $signed({1'h0, smod_35778[15:0]}) < $signed({1'h0, sel_35850}) ? smod_35778[15:0] : sel_35850;
  assign umul_36047 = umul22b_16b_x_6b(array_index_35865, 6'h3b);
  assign add_36049 = {1'h0, umul_35851[21:1]} + 22'h00_1f59;
  assign sel_36054 = $signed({1'h0, smod_35783[15:0]}) < $signed({1'h0, sel_35858}) ? smod_35783[15:0] : sel_35858;
  assign array_index_36055 = set1_unflattened[5'h07];
  assign smod_36059 = $unsigned($signed({9'h000, add_35921, umul_35729[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_36061 = set2_unflattened[5'h07];
  assign smod_36065 = $unsigned($signed({9'h000, add_35929, umul_35737[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_36115 = umul22b_16b_x_6b(array_index_36055, 6'h35);
  assign add_36117 = {1'h0, umul_35919[21:7]} + 16'h007d;
  assign sel_36122 = $signed({1'h0, smod_35863[15:0]}) < $signed({1'h0, sel_35926}) ? smod_35863[15:0] : sel_35926;
  assign umul_36123 = umul22b_16b_x_6b(array_index_36061, 6'h35);
  assign add_36125 = {1'h0, umul_35927[21:7]} + 16'h007d;
  assign sel_36130 = $signed({1'h0, smod_35869[15:0]}) < $signed({1'h0, sel_35934}) ? smod_35869[15:0] : sel_35934;
  assign smod_36134 = $unsigned($signed({8'h00, add_35993, umul_35799[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_36139 = $unsigned($signed({8'h00, add_36001, umul_35805[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_36144 = $unsigned($signed({8'h00, add_36009, umul_35811[0]}) % $signed(32'h0000_3ffd));
  assign smod_36149 = $unsigned($signed({8'h00, add_36017, umul_35819[0]}) % $signed(32'h0000_3ffd));
  assign smod_36154 = $unsigned($signed({9'h000, add_36025, umul_35827[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_36159 = $unsigned($signed({9'h000, add_36033, umul_35835[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_36164 = $unsigned($signed({9'h000, add_36041, umul_35843[0]}) % $signed(32'h0000_3ffd));
  assign smod_36169 = $unsigned($signed({9'h000, add_36049, umul_35851[0]}) % $signed(32'h0000_3ffd));
  assign umul_36185 = umul23b_16b_x_7b(array_index_35507, 7'h49);
  assign add_36187 = {1'h0, umul_35991[22:3]} + 21'h00_07e9;
  assign sel_36192 = $signed({1'h0, smod_35938[15:0]}) < $signed({1'h0, sel_35998}) ? smod_35938[15:0] : sel_35998;
  assign umul_36193 = umul23b_16b_x_7b(array_index_35513, 7'h49);
  assign add_36195 = {1'h0, umul_35999[22:3]} + 21'h00_07e9;
  assign sel_36200 = $signed({1'h0, smod_35944[15:0]}) < $signed({1'h0, sel_36006}) ? smod_35944[15:0] : sel_36006;
  assign umul_36201 = umul23b_16b_x_7b(array_index_35673, 7'h47);
  assign add_36203 = {1'h0, umul_36007[22:1]} + 23'h00_1f8b;
  assign sel_36208 = $signed({1'h0, smod_35950[15:0]}) < $signed({1'h0, sel_36014}) ? smod_35950[15:0] : sel_36014;
  assign umul_36209 = umul23b_16b_x_7b(array_index_35679, 7'h47);
  assign add_36211 = {1'h0, umul_36015[22:1]} + 23'h00_1f8b;
  assign sel_36216 = $signed({1'h0, smod_35955[15:0]}) < $signed({1'h0, sel_36022}) ? smod_35955[15:0] : sel_36022;
  assign umul_36217 = umul22b_16b_x_6b(array_index_35859, 6'h3d);
  assign add_36219 = {1'h0, umul_36023[21:2]} + 21'h00_0fb9;
  assign sel_36224 = $signed({1'h0, smod_35960[15:0]}) < $signed({1'h0, sel_36030}) ? smod_35960[15:0] : sel_36030;
  assign umul_36225 = umul22b_16b_x_6b(array_index_35865, 6'h3d);
  assign add_36227 = {1'h0, umul_36031[21:2]} + 21'h00_0fb9;
  assign sel_36232 = $signed({1'h0, smod_35965[15:0]}) < $signed({1'h0, sel_36038}) ? smod_35965[15:0] : sel_36038;
  assign umul_36233 = umul22b_16b_x_6b(array_index_36055, 6'h3b);
  assign add_36235 = {1'h0, umul_36039[21:1]} + 22'h00_1f59;
  assign sel_36240 = $signed({1'h0, smod_35970[15:0]}) < $signed({1'h0, sel_36046}) ? smod_35970[15:0] : sel_36046;
  assign umul_36241 = umul22b_16b_x_6b(array_index_36061, 6'h3b);
  assign add_36243 = {1'h0, umul_36047[21:1]} + 22'h00_1f59;
  assign sel_36248 = $signed({1'h0, smod_35975[15:0]}) < $signed({1'h0, sel_36054}) ? smod_35975[15:0] : sel_36054;
  assign array_index_36249 = set1_unflattened[5'h08];
  assign smod_36253 = $unsigned($signed({9'h000, add_36117, umul_35919[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_36255 = set2_unflattened[5'h08];
  assign smod_36259 = $unsigned($signed({9'h000, add_36125, umul_35927[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_36309 = umul22b_16b_x_6b(array_index_36249, 6'h35);
  assign add_36311 = {1'h0, umul_36115[21:7]} + 16'h007d;
  assign sel_36316 = $signed({1'h0, smod_36059[15:0]}) < $signed({1'h0, sel_36122}) ? smod_36059[15:0] : sel_36122;
  assign umul_36317 = umul22b_16b_x_6b(array_index_36255, 6'h35);
  assign add_36319 = {1'h0, umul_36123[21:7]} + 16'h007d;
  assign sel_36324 = $signed({1'h0, smod_36065[15:0]}) < $signed({1'h0, sel_36130}) ? smod_36065[15:0] : sel_36130;
  assign smod_36328 = $unsigned($signed({8'h00, add_36187, umul_35991[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_36333 = $unsigned($signed({8'h00, add_36195, umul_35999[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_36338 = $unsigned($signed({8'h00, add_36203, umul_36007[0]}) % $signed(32'h0000_3ffd));
  assign smod_36343 = $unsigned($signed({8'h00, add_36211, umul_36015[0]}) % $signed(32'h0000_3ffd));
  assign smod_36348 = $unsigned($signed({9'h000, add_36219, umul_36023[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_36353 = $unsigned($signed({9'h000, add_36227, umul_36031[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_36358 = $unsigned($signed({9'h000, add_36235, umul_36039[0]}) % $signed(32'h0000_3ffd));
  assign smod_36363 = $unsigned($signed({9'h000, add_36243, umul_36047[0]}) % $signed(32'h0000_3ffd));
  assign umul_36379 = umul23b_16b_x_7b(array_index_35673, 7'h49);
  assign add_36381 = {1'h0, umul_36185[22:3]} + 21'h00_07e9;
  assign sel_36386 = $signed({1'h0, smod_36134[15:0]}) < $signed({1'h0, sel_36192}) ? smod_36134[15:0] : sel_36192;
  assign umul_36387 = umul23b_16b_x_7b(array_index_35679, 7'h49);
  assign add_36389 = {1'h0, umul_36193[22:3]} + 21'h00_07e9;
  assign sel_36394 = $signed({1'h0, smod_36139[15:0]}) < $signed({1'h0, sel_36200}) ? smod_36139[15:0] : sel_36200;
  assign umul_36395 = umul23b_16b_x_7b(array_index_35859, 7'h47);
  assign add_36397 = {1'h0, umul_36201[22:1]} + 23'h00_1f8b;
  assign sel_36402 = $signed({1'h0, smod_36144[15:0]}) < $signed({1'h0, sel_36208}) ? smod_36144[15:0] : sel_36208;
  assign umul_36403 = umul23b_16b_x_7b(array_index_35865, 7'h47);
  assign add_36405 = {1'h0, umul_36209[22:1]} + 23'h00_1f8b;
  assign sel_36410 = $signed({1'h0, smod_36149[15:0]}) < $signed({1'h0, sel_36216}) ? smod_36149[15:0] : sel_36216;
  assign umul_36411 = umul22b_16b_x_6b(array_index_36055, 6'h3d);
  assign add_36413 = {1'h0, umul_36217[21:2]} + 21'h00_0fb9;
  assign sel_36418 = $signed({1'h0, smod_36154[15:0]}) < $signed({1'h0, sel_36224}) ? smod_36154[15:0] : sel_36224;
  assign umul_36419 = umul22b_16b_x_6b(array_index_36061, 6'h3d);
  assign add_36421 = {1'h0, umul_36225[21:2]} + 21'h00_0fb9;
  assign sel_36426 = $signed({1'h0, smod_36159[15:0]}) < $signed({1'h0, sel_36232}) ? smod_36159[15:0] : sel_36232;
  assign umul_36427 = umul22b_16b_x_6b(array_index_36249, 6'h3b);
  assign add_36429 = {1'h0, umul_36233[21:1]} + 22'h00_1f59;
  assign sel_36434 = $signed({1'h0, smod_36164[15:0]}) < $signed({1'h0, sel_36240}) ? smod_36164[15:0] : sel_36240;
  assign umul_36435 = umul22b_16b_x_6b(array_index_36255, 6'h3b);
  assign add_36437 = {1'h0, umul_36241[21:1]} + 22'h00_1f59;
  assign sel_36442 = $signed({1'h0, smod_36169[15:0]}) < $signed({1'h0, sel_36248}) ? smod_36169[15:0] : sel_36248;
  assign array_index_36443 = set1_unflattened[5'h09];
  assign smod_36447 = $unsigned($signed({9'h000, add_36311, umul_36115[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_36449 = set2_unflattened[5'h09];
  assign smod_36453 = $unsigned($signed({9'h000, add_36319, umul_36123[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_36503 = umul22b_16b_x_6b(array_index_36443, 6'h35);
  assign add_36505 = {1'h0, umul_36309[21:7]} + 16'h007d;
  assign sel_36510 = $signed({1'h0, smod_36253[15:0]}) < $signed({1'h0, sel_36316}) ? smod_36253[15:0] : sel_36316;
  assign umul_36511 = umul22b_16b_x_6b(array_index_36449, 6'h35);
  assign add_36513 = {1'h0, umul_36317[21:7]} + 16'h007d;
  assign sel_36518 = $signed({1'h0, smod_36259[15:0]}) < $signed({1'h0, sel_36324}) ? smod_36259[15:0] : sel_36324;
  assign smod_36522 = $unsigned($signed({8'h00, add_36381, umul_36185[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_36527 = $unsigned($signed({8'h00, add_36389, umul_36193[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_36532 = $unsigned($signed({8'h00, add_36397, umul_36201[0]}) % $signed(32'h0000_3ffd));
  assign smod_36537 = $unsigned($signed({8'h00, add_36405, umul_36209[0]}) % $signed(32'h0000_3ffd));
  assign smod_36542 = $unsigned($signed({9'h000, add_36413, umul_36217[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_36547 = $unsigned($signed({9'h000, add_36421, umul_36225[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_36552 = $unsigned($signed({9'h000, add_36429, umul_36233[0]}) % $signed(32'h0000_3ffd));
  assign smod_36557 = $unsigned($signed({9'h000, add_36437, umul_36241[0]}) % $signed(32'h0000_3ffd));
  assign umul_36573 = umul23b_16b_x_7b(array_index_35859, 7'h49);
  assign add_36575 = {1'h0, umul_36379[22:3]} + 21'h00_07e9;
  assign sel_36580 = $signed({1'h0, smod_36328[15:0]}) < $signed({1'h0, sel_36386}) ? smod_36328[15:0] : sel_36386;
  assign umul_36581 = umul23b_16b_x_7b(array_index_35865, 7'h49);
  assign add_36583 = {1'h0, umul_36387[22:3]} + 21'h00_07e9;
  assign sel_36588 = $signed({1'h0, smod_36333[15:0]}) < $signed({1'h0, sel_36394}) ? smod_36333[15:0] : sel_36394;
  assign umul_36589 = umul23b_16b_x_7b(array_index_36055, 7'h47);
  assign add_36591 = {1'h0, umul_36395[22:1]} + 23'h00_1f8b;
  assign sel_36596 = $signed({1'h0, smod_36338[15:0]}) < $signed({1'h0, sel_36402}) ? smod_36338[15:0] : sel_36402;
  assign umul_36597 = umul23b_16b_x_7b(array_index_36061, 7'h47);
  assign add_36599 = {1'h0, umul_36403[22:1]} + 23'h00_1f8b;
  assign sel_36604 = $signed({1'h0, smod_36343[15:0]}) < $signed({1'h0, sel_36410}) ? smod_36343[15:0] : sel_36410;
  assign umul_36605 = umul22b_16b_x_6b(array_index_36249, 6'h3d);
  assign add_36607 = {1'h0, umul_36411[21:2]} + 21'h00_0fb9;
  assign sel_36612 = $signed({1'h0, smod_36348[15:0]}) < $signed({1'h0, sel_36418}) ? smod_36348[15:0] : sel_36418;
  assign umul_36613 = umul22b_16b_x_6b(array_index_36255, 6'h3d);
  assign add_36615 = {1'h0, umul_36419[21:2]} + 21'h00_0fb9;
  assign sel_36620 = $signed({1'h0, smod_36353[15:0]}) < $signed({1'h0, sel_36426}) ? smod_36353[15:0] : sel_36426;
  assign umul_36621 = umul22b_16b_x_6b(array_index_36443, 6'h3b);
  assign add_36623 = {1'h0, umul_36427[21:1]} + 22'h00_1f59;
  assign sel_36628 = $signed({1'h0, smod_36358[15:0]}) < $signed({1'h0, sel_36434}) ? smod_36358[15:0] : sel_36434;
  assign umul_36629 = umul22b_16b_x_6b(array_index_36449, 6'h3b);
  assign add_36631 = {1'h0, umul_36435[21:1]} + 22'h00_1f59;
  assign sel_36636 = $signed({1'h0, smod_36363[15:0]}) < $signed({1'h0, sel_36442}) ? smod_36363[15:0] : sel_36442;
  assign array_index_36637 = set1_unflattened[5'h0a];
  assign smod_36641 = $unsigned($signed({9'h000, add_36505, umul_36309[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_36643 = set2_unflattened[5'h0a];
  assign smod_36647 = $unsigned($signed({9'h000, add_36513, umul_36317[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_36697 = umul22b_16b_x_6b(array_index_36637, 6'h35);
  assign add_36699 = {1'h0, umul_36503[21:7]} + 16'h007d;
  assign sel_36704 = $signed({1'h0, smod_36447[15:0]}) < $signed({1'h0, sel_36510}) ? smod_36447[15:0] : sel_36510;
  assign umul_36705 = umul22b_16b_x_6b(array_index_36643, 6'h35);
  assign add_36707 = {1'h0, umul_36511[21:7]} + 16'h007d;
  assign sel_36712 = $signed({1'h0, smod_36453[15:0]}) < $signed({1'h0, sel_36518}) ? smod_36453[15:0] : sel_36518;
  assign smod_36716 = $unsigned($signed({8'h00, add_36575, umul_36379[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_36721 = $unsigned($signed({8'h00, add_36583, umul_36387[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_36726 = $unsigned($signed({8'h00, add_36591, umul_36395[0]}) % $signed(32'h0000_3ffd));
  assign smod_36731 = $unsigned($signed({8'h00, add_36599, umul_36403[0]}) % $signed(32'h0000_3ffd));
  assign smod_36736 = $unsigned($signed({9'h000, add_36607, umul_36411[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_36741 = $unsigned($signed({9'h000, add_36615, umul_36419[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_36746 = $unsigned($signed({9'h000, add_36623, umul_36427[0]}) % $signed(32'h0000_3ffd));
  assign smod_36751 = $unsigned($signed({9'h000, add_36631, umul_36435[0]}) % $signed(32'h0000_3ffd));
  assign umul_36767 = umul23b_16b_x_7b(array_index_36055, 7'h49);
  assign add_36769 = {1'h0, umul_36573[22:3]} + 21'h00_07e9;
  assign sel_36774 = $signed({1'h0, smod_36522[15:0]}) < $signed({1'h0, sel_36580}) ? smod_36522[15:0] : sel_36580;
  assign umul_36775 = umul23b_16b_x_7b(array_index_36061, 7'h49);
  assign add_36777 = {1'h0, umul_36581[22:3]} + 21'h00_07e9;
  assign sel_36782 = $signed({1'h0, smod_36527[15:0]}) < $signed({1'h0, sel_36588}) ? smod_36527[15:0] : sel_36588;
  assign umul_36783 = umul23b_16b_x_7b(array_index_36249, 7'h47);
  assign add_36785 = {1'h0, umul_36589[22:1]} + 23'h00_1f8b;
  assign sel_36790 = $signed({1'h0, smod_36532[15:0]}) < $signed({1'h0, sel_36596}) ? smod_36532[15:0] : sel_36596;
  assign umul_36791 = umul23b_16b_x_7b(array_index_36255, 7'h47);
  assign add_36793 = {1'h0, umul_36597[22:1]} + 23'h00_1f8b;
  assign sel_36798 = $signed({1'h0, smod_36537[15:0]}) < $signed({1'h0, sel_36604}) ? smod_36537[15:0] : sel_36604;
  assign umul_36799 = umul22b_16b_x_6b(array_index_36443, 6'h3d);
  assign add_36801 = {1'h0, umul_36605[21:2]} + 21'h00_0fb9;
  assign sel_36806 = $signed({1'h0, smod_36542[15:0]}) < $signed({1'h0, sel_36612}) ? smod_36542[15:0] : sel_36612;
  assign umul_36807 = umul22b_16b_x_6b(array_index_36449, 6'h3d);
  assign add_36809 = {1'h0, umul_36613[21:2]} + 21'h00_0fb9;
  assign sel_36814 = $signed({1'h0, smod_36547[15:0]}) < $signed({1'h0, sel_36620}) ? smod_36547[15:0] : sel_36620;
  assign umul_36815 = umul22b_16b_x_6b(array_index_36637, 6'h3b);
  assign add_36817 = {1'h0, umul_36621[21:1]} + 22'h00_1f59;
  assign sel_36822 = $signed({1'h0, smod_36552[15:0]}) < $signed({1'h0, sel_36628}) ? smod_36552[15:0] : sel_36628;
  assign umul_36823 = umul22b_16b_x_6b(array_index_36643, 6'h3b);
  assign add_36825 = {1'h0, umul_36629[21:1]} + 22'h00_1f59;
  assign sel_36830 = $signed({1'h0, smod_36557[15:0]}) < $signed({1'h0, sel_36636}) ? smod_36557[15:0] : sel_36636;
  assign array_index_36831 = set1_unflattened[5'h0b];
  assign smod_36835 = $unsigned($signed({9'h000, add_36699, umul_36503[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_36837 = set2_unflattened[5'h0b];
  assign smod_36841 = $unsigned($signed({9'h000, add_36707, umul_36511[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_36891 = umul22b_16b_x_6b(array_index_36831, 6'h35);
  assign add_36893 = {1'h0, umul_36697[21:7]} + 16'h007d;
  assign sel_36898 = $signed({1'h0, smod_36641[15:0]}) < $signed({1'h0, sel_36704}) ? smod_36641[15:0] : sel_36704;
  assign umul_36899 = umul22b_16b_x_6b(array_index_36837, 6'h35);
  assign add_36901 = {1'h0, umul_36705[21:7]} + 16'h007d;
  assign sel_36906 = $signed({1'h0, smod_36647[15:0]}) < $signed({1'h0, sel_36712}) ? smod_36647[15:0] : sel_36712;
  assign smod_36910 = $unsigned($signed({8'h00, add_36769, umul_36573[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_36915 = $unsigned($signed({8'h00, add_36777, umul_36581[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_36920 = $unsigned($signed({8'h00, add_36785, umul_36589[0]}) % $signed(32'h0000_3ffd));
  assign smod_36925 = $unsigned($signed({8'h00, add_36793, umul_36597[0]}) % $signed(32'h0000_3ffd));
  assign smod_36930 = $unsigned($signed({9'h000, add_36801, umul_36605[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_36935 = $unsigned($signed({9'h000, add_36809, umul_36613[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_36940 = $unsigned($signed({9'h000, add_36817, umul_36621[0]}) % $signed(32'h0000_3ffd));
  assign smod_36945 = $unsigned($signed({9'h000, add_36825, umul_36629[0]}) % $signed(32'h0000_3ffd));
  assign umul_36961 = umul23b_16b_x_7b(array_index_36249, 7'h49);
  assign add_36963 = {1'h0, umul_36767[22:3]} + 21'h00_07e9;
  assign sel_36968 = $signed({1'h0, smod_36716[15:0]}) < $signed({1'h0, sel_36774}) ? smod_36716[15:0] : sel_36774;
  assign umul_36969 = umul23b_16b_x_7b(array_index_36255, 7'h49);
  assign add_36971 = {1'h0, umul_36775[22:3]} + 21'h00_07e9;
  assign sel_36976 = $signed({1'h0, smod_36721[15:0]}) < $signed({1'h0, sel_36782}) ? smod_36721[15:0] : sel_36782;
  assign umul_36977 = umul23b_16b_x_7b(array_index_36443, 7'h47);
  assign add_36979 = {1'h0, umul_36783[22:1]} + 23'h00_1f8b;
  assign sel_36984 = $signed({1'h0, smod_36726[15:0]}) < $signed({1'h0, sel_36790}) ? smod_36726[15:0] : sel_36790;
  assign umul_36985 = umul23b_16b_x_7b(array_index_36449, 7'h47);
  assign add_36987 = {1'h0, umul_36791[22:1]} + 23'h00_1f8b;
  assign sel_36992 = $signed({1'h0, smod_36731[15:0]}) < $signed({1'h0, sel_36798}) ? smod_36731[15:0] : sel_36798;
  assign umul_36993 = umul22b_16b_x_6b(array_index_36637, 6'h3d);
  assign add_36995 = {1'h0, umul_36799[21:2]} + 21'h00_0fb9;
  assign sel_37000 = $signed({1'h0, smod_36736[15:0]}) < $signed({1'h0, sel_36806}) ? smod_36736[15:0] : sel_36806;
  assign umul_37001 = umul22b_16b_x_6b(array_index_36643, 6'h3d);
  assign add_37003 = {1'h0, umul_36807[21:2]} + 21'h00_0fb9;
  assign sel_37008 = $signed({1'h0, smod_36741[15:0]}) < $signed({1'h0, sel_36814}) ? smod_36741[15:0] : sel_36814;
  assign umul_37009 = umul22b_16b_x_6b(array_index_36831, 6'h3b);
  assign add_37011 = {1'h0, umul_36815[21:1]} + 22'h00_1f59;
  assign sel_37016 = $signed({1'h0, smod_36746[15:0]}) < $signed({1'h0, sel_36822}) ? smod_36746[15:0] : sel_36822;
  assign umul_37017 = umul22b_16b_x_6b(array_index_36837, 6'h3b);
  assign add_37019 = {1'h0, umul_36823[21:1]} + 22'h00_1f59;
  assign sel_37024 = $signed({1'h0, smod_36751[15:0]}) < $signed({1'h0, sel_36830}) ? smod_36751[15:0] : sel_36830;
  assign array_index_37025 = set1_unflattened[5'h0c];
  assign smod_37029 = $unsigned($signed({9'h000, add_36893, umul_36697[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_37031 = set2_unflattened[5'h0c];
  assign smod_37035 = $unsigned($signed({9'h000, add_36901, umul_36705[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_37085 = umul22b_16b_x_6b(array_index_37025, 6'h35);
  assign add_37087 = {1'h0, umul_36891[21:7]} + 16'h007d;
  assign sel_37092 = $signed({1'h0, smod_36835[15:0]}) < $signed({1'h0, sel_36898}) ? smod_36835[15:0] : sel_36898;
  assign umul_37093 = umul22b_16b_x_6b(array_index_37031, 6'h35);
  assign add_37095 = {1'h0, umul_36899[21:7]} + 16'h007d;
  assign sel_37100 = $signed({1'h0, smod_36841[15:0]}) < $signed({1'h0, sel_36906}) ? smod_36841[15:0] : sel_36906;
  assign smod_37104 = $unsigned($signed({8'h00, add_36963, umul_36767[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_37109 = $unsigned($signed({8'h00, add_36971, umul_36775[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_37114 = $unsigned($signed({8'h00, add_36979, umul_36783[0]}) % $signed(32'h0000_3ffd));
  assign smod_37119 = $unsigned($signed({8'h00, add_36987, umul_36791[0]}) % $signed(32'h0000_3ffd));
  assign smod_37124 = $unsigned($signed({9'h000, add_36995, umul_36799[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_37129 = $unsigned($signed({9'h000, add_37003, umul_36807[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_37134 = $unsigned($signed({9'h000, add_37011, umul_36815[0]}) % $signed(32'h0000_3ffd));
  assign smod_37139 = $unsigned($signed({9'h000, add_37019, umul_36823[0]}) % $signed(32'h0000_3ffd));
  assign umul_37155 = umul23b_16b_x_7b(array_index_36443, 7'h49);
  assign add_37157 = {1'h0, umul_36961[22:3]} + 21'h00_07e9;
  assign sel_37162 = $signed({1'h0, smod_36910[15:0]}) < $signed({1'h0, sel_36968}) ? smod_36910[15:0] : sel_36968;
  assign umul_37163 = umul23b_16b_x_7b(array_index_36449, 7'h49);
  assign add_37165 = {1'h0, umul_36969[22:3]} + 21'h00_07e9;
  assign sel_37170 = $signed({1'h0, smod_36915[15:0]}) < $signed({1'h0, sel_36976}) ? smod_36915[15:0] : sel_36976;
  assign umul_37171 = umul23b_16b_x_7b(array_index_36637, 7'h47);
  assign add_37173 = {1'h0, umul_36977[22:1]} + 23'h00_1f8b;
  assign sel_37178 = $signed({1'h0, smod_36920[15:0]}) < $signed({1'h0, sel_36984}) ? smod_36920[15:0] : sel_36984;
  assign umul_37179 = umul23b_16b_x_7b(array_index_36643, 7'h47);
  assign add_37181 = {1'h0, umul_36985[22:1]} + 23'h00_1f8b;
  assign sel_37186 = $signed({1'h0, smod_36925[15:0]}) < $signed({1'h0, sel_36992}) ? smod_36925[15:0] : sel_36992;
  assign umul_37187 = umul22b_16b_x_6b(array_index_36831, 6'h3d);
  assign add_37189 = {1'h0, umul_36993[21:2]} + 21'h00_0fb9;
  assign sel_37194 = $signed({1'h0, smod_36930[15:0]}) < $signed({1'h0, sel_37000}) ? smod_36930[15:0] : sel_37000;
  assign umul_37195 = umul22b_16b_x_6b(array_index_36837, 6'h3d);
  assign add_37197 = {1'h0, umul_37001[21:2]} + 21'h00_0fb9;
  assign sel_37202 = $signed({1'h0, smod_36935[15:0]}) < $signed({1'h0, sel_37008}) ? smod_36935[15:0] : sel_37008;
  assign umul_37203 = umul22b_16b_x_6b(array_index_37025, 6'h3b);
  assign add_37205 = {1'h0, umul_37009[21:1]} + 22'h00_1f59;
  assign sel_37210 = $signed({1'h0, smod_36940[15:0]}) < $signed({1'h0, sel_37016}) ? smod_36940[15:0] : sel_37016;
  assign umul_37211 = umul22b_16b_x_6b(array_index_37031, 6'h3b);
  assign add_37213 = {1'h0, umul_37017[21:1]} + 22'h00_1f59;
  assign sel_37218 = $signed({1'h0, smod_36945[15:0]}) < $signed({1'h0, sel_37024}) ? smod_36945[15:0] : sel_37024;
  assign array_index_37219 = set1_unflattened[5'h0d];
  assign smod_37223 = $unsigned($signed({9'h000, add_37087, umul_36891[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_37225 = set2_unflattened[5'h0d];
  assign smod_37229 = $unsigned($signed({9'h000, add_37095, umul_36899[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_37279 = umul22b_16b_x_6b(array_index_37219, 6'h35);
  assign add_37281 = {1'h0, umul_37085[21:7]} + 16'h007d;
  assign sel_37286 = $signed({1'h0, smod_37029[15:0]}) < $signed({1'h0, sel_37092}) ? smod_37029[15:0] : sel_37092;
  assign umul_37287 = umul22b_16b_x_6b(array_index_37225, 6'h35);
  assign add_37289 = {1'h0, umul_37093[21:7]} + 16'h007d;
  assign sel_37294 = $signed({1'h0, smod_37035[15:0]}) < $signed({1'h0, sel_37100}) ? smod_37035[15:0] : sel_37100;
  assign smod_37298 = $unsigned($signed({8'h00, add_37157, umul_36961[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_37303 = $unsigned($signed({8'h00, add_37165, umul_36969[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_37308 = $unsigned($signed({8'h00, add_37173, umul_36977[0]}) % $signed(32'h0000_3ffd));
  assign smod_37313 = $unsigned($signed({8'h00, add_37181, umul_36985[0]}) % $signed(32'h0000_3ffd));
  assign smod_37318 = $unsigned($signed({9'h000, add_37189, umul_36993[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_37323 = $unsigned($signed({9'h000, add_37197, umul_37001[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_37328 = $unsigned($signed({9'h000, add_37205, umul_37009[0]}) % $signed(32'h0000_3ffd));
  assign smod_37333 = $unsigned($signed({9'h000, add_37213, umul_37017[0]}) % $signed(32'h0000_3ffd));
  assign umul_37349 = umul23b_16b_x_7b(array_index_36637, 7'h49);
  assign add_37351 = {1'h0, umul_37155[22:3]} + 21'h00_07e9;
  assign sel_37356 = $signed({1'h0, smod_37104[15:0]}) < $signed({1'h0, sel_37162}) ? smod_37104[15:0] : sel_37162;
  assign umul_37357 = umul23b_16b_x_7b(array_index_36643, 7'h49);
  assign add_37359 = {1'h0, umul_37163[22:3]} + 21'h00_07e9;
  assign sel_37364 = $signed({1'h0, smod_37109[15:0]}) < $signed({1'h0, sel_37170}) ? smod_37109[15:0] : sel_37170;
  assign umul_37365 = umul23b_16b_x_7b(array_index_36831, 7'h47);
  assign add_37367 = {1'h0, umul_37171[22:1]} + 23'h00_1f8b;
  assign sel_37372 = $signed({1'h0, smod_37114[15:0]}) < $signed({1'h0, sel_37178}) ? smod_37114[15:0] : sel_37178;
  assign umul_37373 = umul23b_16b_x_7b(array_index_36837, 7'h47);
  assign add_37375 = {1'h0, umul_37179[22:1]} + 23'h00_1f8b;
  assign sel_37380 = $signed({1'h0, smod_37119[15:0]}) < $signed({1'h0, sel_37186}) ? smod_37119[15:0] : sel_37186;
  assign umul_37381 = umul22b_16b_x_6b(array_index_37025, 6'h3d);
  assign add_37383 = {1'h0, umul_37187[21:2]} + 21'h00_0fb9;
  assign sel_37388 = $signed({1'h0, smod_37124[15:0]}) < $signed({1'h0, sel_37194}) ? smod_37124[15:0] : sel_37194;
  assign umul_37389 = umul22b_16b_x_6b(array_index_37031, 6'h3d);
  assign add_37391 = {1'h0, umul_37195[21:2]} + 21'h00_0fb9;
  assign sel_37396 = $signed({1'h0, smod_37129[15:0]}) < $signed({1'h0, sel_37202}) ? smod_37129[15:0] : sel_37202;
  assign umul_37397 = umul22b_16b_x_6b(array_index_37219, 6'h3b);
  assign add_37399 = {1'h0, umul_37203[21:1]} + 22'h00_1f59;
  assign sel_37404 = $signed({1'h0, smod_37134[15:0]}) < $signed({1'h0, sel_37210}) ? smod_37134[15:0] : sel_37210;
  assign umul_37405 = umul22b_16b_x_6b(array_index_37225, 6'h3b);
  assign add_37407 = {1'h0, umul_37211[21:1]} + 22'h00_1f59;
  assign sel_37412 = $signed({1'h0, smod_37139[15:0]}) < $signed({1'h0, sel_37218}) ? smod_37139[15:0] : sel_37218;
  assign array_index_37413 = set1_unflattened[5'h0e];
  assign smod_37417 = $unsigned($signed({9'h000, add_37281, umul_37085[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_37419 = set2_unflattened[5'h0e];
  assign smod_37423 = $unsigned($signed({9'h000, add_37289, umul_37093[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_37473 = umul22b_16b_x_6b(array_index_37413, 6'h35);
  assign add_37475 = {1'h0, umul_37279[21:7]} + 16'h007d;
  assign sel_37480 = $signed({1'h0, smod_37223[15:0]}) < $signed({1'h0, sel_37286}) ? smod_37223[15:0] : sel_37286;
  assign umul_37481 = umul22b_16b_x_6b(array_index_37419, 6'h35);
  assign add_37483 = {1'h0, umul_37287[21:7]} + 16'h007d;
  assign sel_37488 = $signed({1'h0, smod_37229[15:0]}) < $signed({1'h0, sel_37294}) ? smod_37229[15:0] : sel_37294;
  assign smod_37492 = $unsigned($signed({8'h00, add_37351, umul_37155[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_37497 = $unsigned($signed({8'h00, add_37359, umul_37163[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_37502 = $unsigned($signed({8'h00, add_37367, umul_37171[0]}) % $signed(32'h0000_3ffd));
  assign smod_37507 = $unsigned($signed({8'h00, add_37375, umul_37179[0]}) % $signed(32'h0000_3ffd));
  assign smod_37512 = $unsigned($signed({9'h000, add_37383, umul_37187[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_37517 = $unsigned($signed({9'h000, add_37391, umul_37195[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_37522 = $unsigned($signed({9'h000, add_37399, umul_37203[0]}) % $signed(32'h0000_3ffd));
  assign smod_37527 = $unsigned($signed({9'h000, add_37407, umul_37211[0]}) % $signed(32'h0000_3ffd));
  assign umul_37543 = umul23b_16b_x_7b(array_index_36831, 7'h49);
  assign add_37545 = {1'h0, umul_37349[22:3]} + 21'h00_07e9;
  assign sel_37550 = $signed({1'h0, smod_37298[15:0]}) < $signed({1'h0, sel_37356}) ? smod_37298[15:0] : sel_37356;
  assign umul_37551 = umul23b_16b_x_7b(array_index_36837, 7'h49);
  assign add_37553 = {1'h0, umul_37357[22:3]} + 21'h00_07e9;
  assign sel_37558 = $signed({1'h0, smod_37303[15:0]}) < $signed({1'h0, sel_37364}) ? smod_37303[15:0] : sel_37364;
  assign umul_37559 = umul23b_16b_x_7b(array_index_37025, 7'h47);
  assign add_37561 = {1'h0, umul_37365[22:1]} + 23'h00_1f8b;
  assign sel_37566 = $signed({1'h0, smod_37308[15:0]}) < $signed({1'h0, sel_37372}) ? smod_37308[15:0] : sel_37372;
  assign umul_37567 = umul23b_16b_x_7b(array_index_37031, 7'h47);
  assign add_37569 = {1'h0, umul_37373[22:1]} + 23'h00_1f8b;
  assign sel_37574 = $signed({1'h0, smod_37313[15:0]}) < $signed({1'h0, sel_37380}) ? smod_37313[15:0] : sel_37380;
  assign umul_37575 = umul22b_16b_x_6b(array_index_37219, 6'h3d);
  assign add_37577 = {1'h0, umul_37381[21:2]} + 21'h00_0fb9;
  assign sel_37582 = $signed({1'h0, smod_37318[15:0]}) < $signed({1'h0, sel_37388}) ? smod_37318[15:0] : sel_37388;
  assign umul_37583 = umul22b_16b_x_6b(array_index_37225, 6'h3d);
  assign add_37585 = {1'h0, umul_37389[21:2]} + 21'h00_0fb9;
  assign sel_37590 = $signed({1'h0, smod_37323[15:0]}) < $signed({1'h0, sel_37396}) ? smod_37323[15:0] : sel_37396;
  assign umul_37591 = umul22b_16b_x_6b(array_index_37413, 6'h3b);
  assign add_37593 = {1'h0, umul_37397[21:1]} + 22'h00_1f59;
  assign sel_37598 = $signed({1'h0, smod_37328[15:0]}) < $signed({1'h0, sel_37404}) ? smod_37328[15:0] : sel_37404;
  assign umul_37599 = umul22b_16b_x_6b(array_index_37419, 6'h3b);
  assign add_37601 = {1'h0, umul_37405[21:1]} + 22'h00_1f59;
  assign sel_37606 = $signed({1'h0, smod_37333[15:0]}) < $signed({1'h0, sel_37412}) ? smod_37333[15:0] : sel_37412;
  assign array_index_37607 = set1_unflattened[5'h0f];
  assign smod_37611 = $unsigned($signed({9'h000, add_37475, umul_37279[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_37613 = set2_unflattened[5'h0f];
  assign smod_37617 = $unsigned($signed({9'h000, add_37483, umul_37287[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_37667 = umul22b_16b_x_6b(array_index_37607, 6'h35);
  assign add_37669 = {1'h0, umul_37473[21:7]} + 16'h007d;
  assign sel_37674 = $signed({1'h0, smod_37417[15:0]}) < $signed({1'h0, sel_37480}) ? smod_37417[15:0] : sel_37480;
  assign umul_37675 = umul22b_16b_x_6b(array_index_37613, 6'h35);
  assign add_37677 = {1'h0, umul_37481[21:7]} + 16'h007d;
  assign sel_37682 = $signed({1'h0, smod_37423[15:0]}) < $signed({1'h0, sel_37488}) ? smod_37423[15:0] : sel_37488;
  assign smod_37686 = $unsigned($signed({8'h00, add_37545, umul_37349[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_37691 = $unsigned($signed({8'h00, add_37553, umul_37357[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_37696 = $unsigned($signed({8'h00, add_37561, umul_37365[0]}) % $signed(32'h0000_3ffd));
  assign smod_37701 = $unsigned($signed({8'h00, add_37569, umul_37373[0]}) % $signed(32'h0000_3ffd));
  assign smod_37706 = $unsigned($signed({9'h000, add_37577, umul_37381[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_37711 = $unsigned($signed({9'h000, add_37585, umul_37389[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_37716 = $unsigned($signed({9'h000, add_37593, umul_37397[0]}) % $signed(32'h0000_3ffd));
  assign smod_37721 = $unsigned($signed({9'h000, add_37601, umul_37405[0]}) % $signed(32'h0000_3ffd));
  assign umul_37737 = umul23b_16b_x_7b(array_index_37025, 7'h49);
  assign add_37739 = {1'h0, umul_37543[22:3]} + 21'h00_07e9;
  assign sel_37744 = $signed({1'h0, smod_37492[15:0]}) < $signed({1'h0, sel_37550}) ? smod_37492[15:0] : sel_37550;
  assign umul_37745 = umul23b_16b_x_7b(array_index_37031, 7'h49);
  assign add_37747 = {1'h0, umul_37551[22:3]} + 21'h00_07e9;
  assign sel_37752 = $signed({1'h0, smod_37497[15:0]}) < $signed({1'h0, sel_37558}) ? smod_37497[15:0] : sel_37558;
  assign umul_37753 = umul23b_16b_x_7b(array_index_37219, 7'h47);
  assign add_37755 = {1'h0, umul_37559[22:1]} + 23'h00_1f8b;
  assign sel_37760 = $signed({1'h0, smod_37502[15:0]}) < $signed({1'h0, sel_37566}) ? smod_37502[15:0] : sel_37566;
  assign umul_37761 = umul23b_16b_x_7b(array_index_37225, 7'h47);
  assign add_37763 = {1'h0, umul_37567[22:1]} + 23'h00_1f8b;
  assign sel_37768 = $signed({1'h0, smod_37507[15:0]}) < $signed({1'h0, sel_37574}) ? smod_37507[15:0] : sel_37574;
  assign umul_37769 = umul22b_16b_x_6b(array_index_37413, 6'h3d);
  assign add_37771 = {1'h0, umul_37575[21:2]} + 21'h00_0fb9;
  assign sel_37776 = $signed({1'h0, smod_37512[15:0]}) < $signed({1'h0, sel_37582}) ? smod_37512[15:0] : sel_37582;
  assign umul_37777 = umul22b_16b_x_6b(array_index_37419, 6'h3d);
  assign add_37779 = {1'h0, umul_37583[21:2]} + 21'h00_0fb9;
  assign sel_37784 = $signed({1'h0, smod_37517[15:0]}) < $signed({1'h0, sel_37590}) ? smod_37517[15:0] : sel_37590;
  assign umul_37785 = umul22b_16b_x_6b(array_index_37607, 6'h3b);
  assign add_37787 = {1'h0, umul_37591[21:1]} + 22'h00_1f59;
  assign sel_37792 = $signed({1'h0, smod_37522[15:0]}) < $signed({1'h0, sel_37598}) ? smod_37522[15:0] : sel_37598;
  assign umul_37793 = umul22b_16b_x_6b(array_index_37613, 6'h3b);
  assign add_37795 = {1'h0, umul_37599[21:1]} + 22'h00_1f59;
  assign sel_37800 = $signed({1'h0, smod_37527[15:0]}) < $signed({1'h0, sel_37606}) ? smod_37527[15:0] : sel_37606;
  assign array_index_37801 = set1_unflattened[5'h10];
  assign smod_37805 = $unsigned($signed({9'h000, add_37669, umul_37473[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_37807 = set2_unflattened[5'h10];
  assign smod_37811 = $unsigned($signed({9'h000, add_37677, umul_37481[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_37861 = umul22b_16b_x_6b(array_index_37801, 6'h35);
  assign add_37863 = {1'h0, umul_37667[21:7]} + 16'h007d;
  assign sel_37868 = $signed({1'h0, smod_37611[15:0]}) < $signed({1'h0, sel_37674}) ? smod_37611[15:0] : sel_37674;
  assign umul_37869 = umul22b_16b_x_6b(array_index_37807, 6'h35);
  assign add_37871 = {1'h0, umul_37675[21:7]} + 16'h007d;
  assign sel_37876 = $signed({1'h0, smod_37617[15:0]}) < $signed({1'h0, sel_37682}) ? smod_37617[15:0] : sel_37682;
  assign smod_37880 = $unsigned($signed({8'h00, add_37739, umul_37543[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_37885 = $unsigned($signed({8'h00, add_37747, umul_37551[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_37890 = $unsigned($signed({8'h00, add_37755, umul_37559[0]}) % $signed(32'h0000_3ffd));
  assign smod_37895 = $unsigned($signed({8'h00, add_37763, umul_37567[0]}) % $signed(32'h0000_3ffd));
  assign smod_37900 = $unsigned($signed({9'h000, add_37771, umul_37575[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_37905 = $unsigned($signed({9'h000, add_37779, umul_37583[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_37910 = $unsigned($signed({9'h000, add_37787, umul_37591[0]}) % $signed(32'h0000_3ffd));
  assign smod_37915 = $unsigned($signed({9'h000, add_37795, umul_37599[0]}) % $signed(32'h0000_3ffd));
  assign umul_37931 = umul23b_16b_x_7b(array_index_37219, 7'h49);
  assign add_37933 = {1'h0, umul_37737[22:3]} + 21'h00_07e9;
  assign sel_37938 = $signed({1'h0, smod_37686[15:0]}) < $signed({1'h0, sel_37744}) ? smod_37686[15:0] : sel_37744;
  assign umul_37939 = umul23b_16b_x_7b(array_index_37225, 7'h49);
  assign add_37941 = {1'h0, umul_37745[22:3]} + 21'h00_07e9;
  assign sel_37946 = $signed({1'h0, smod_37691[15:0]}) < $signed({1'h0, sel_37752}) ? smod_37691[15:0] : sel_37752;
  assign umul_37947 = umul23b_16b_x_7b(array_index_37413, 7'h47);
  assign add_37949 = {1'h0, umul_37753[22:1]} + 23'h00_1f8b;
  assign sel_37954 = $signed({1'h0, smod_37696[15:0]}) < $signed({1'h0, sel_37760}) ? smod_37696[15:0] : sel_37760;
  assign umul_37955 = umul23b_16b_x_7b(array_index_37419, 7'h47);
  assign add_37957 = {1'h0, umul_37761[22:1]} + 23'h00_1f8b;
  assign sel_37962 = $signed({1'h0, smod_37701[15:0]}) < $signed({1'h0, sel_37768}) ? smod_37701[15:0] : sel_37768;
  assign umul_37963 = umul22b_16b_x_6b(array_index_37607, 6'h3d);
  assign add_37965 = {1'h0, umul_37769[21:2]} + 21'h00_0fb9;
  assign sel_37970 = $signed({1'h0, smod_37706[15:0]}) < $signed({1'h0, sel_37776}) ? smod_37706[15:0] : sel_37776;
  assign umul_37971 = umul22b_16b_x_6b(array_index_37613, 6'h3d);
  assign add_37973 = {1'h0, umul_37777[21:2]} + 21'h00_0fb9;
  assign sel_37978 = $signed({1'h0, smod_37711[15:0]}) < $signed({1'h0, sel_37784}) ? smod_37711[15:0] : sel_37784;
  assign umul_37979 = umul22b_16b_x_6b(array_index_37801, 6'h3b);
  assign add_37981 = {1'h0, umul_37785[21:1]} + 22'h00_1f59;
  assign sel_37986 = $signed({1'h0, smod_37716[15:0]}) < $signed({1'h0, sel_37792}) ? smod_37716[15:0] : sel_37792;
  assign umul_37987 = umul22b_16b_x_6b(array_index_37807, 6'h3b);
  assign add_37989 = {1'h0, umul_37793[21:1]} + 22'h00_1f59;
  assign sel_37994 = $signed({1'h0, smod_37721[15:0]}) < $signed({1'h0, sel_37800}) ? smod_37721[15:0] : sel_37800;
  assign array_index_37995 = set1_unflattened[5'h11];
  assign smod_37999 = $unsigned($signed({9'h000, add_37863, umul_37667[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_38001 = set2_unflattened[5'h11];
  assign smod_38005 = $unsigned($signed({9'h000, add_37871, umul_37675[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_38055 = umul22b_16b_x_6b(array_index_37995, 6'h35);
  assign add_38057 = {1'h0, umul_37861[21:7]} + 16'h007d;
  assign sel_38062 = $signed({1'h0, smod_37805[15:0]}) < $signed({1'h0, sel_37868}) ? smod_37805[15:0] : sel_37868;
  assign umul_38063 = umul22b_16b_x_6b(array_index_38001, 6'h35);
  assign add_38065 = {1'h0, umul_37869[21:7]} + 16'h007d;
  assign sel_38070 = $signed({1'h0, smod_37811[15:0]}) < $signed({1'h0, sel_37876}) ? smod_37811[15:0] : sel_37876;
  assign smod_38074 = $unsigned($signed({8'h00, add_37933, umul_37737[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38079 = $unsigned($signed({8'h00, add_37941, umul_37745[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38084 = $unsigned($signed({8'h00, add_37949, umul_37753[0]}) % $signed(32'h0000_3ffd));
  assign smod_38089 = $unsigned($signed({8'h00, add_37957, umul_37761[0]}) % $signed(32'h0000_3ffd));
  assign smod_38094 = $unsigned($signed({9'h000, add_37965, umul_37769[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_38099 = $unsigned($signed({9'h000, add_37973, umul_37777[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_38104 = $unsigned($signed({9'h000, add_37981, umul_37785[0]}) % $signed(32'h0000_3ffd));
  assign smod_38109 = $unsigned($signed({9'h000, add_37989, umul_37793[0]}) % $signed(32'h0000_3ffd));
  assign umul_38125 = umul23b_16b_x_7b(array_index_37413, 7'h49);
  assign add_38127 = {1'h0, umul_37931[22:3]} + 21'h00_07e9;
  assign sel_38132 = $signed({1'h0, smod_37880[15:0]}) < $signed({1'h0, sel_37938}) ? smod_37880[15:0] : sel_37938;
  assign umul_38133 = umul23b_16b_x_7b(array_index_37419, 7'h49);
  assign add_38135 = {1'h0, umul_37939[22:3]} + 21'h00_07e9;
  assign sel_38140 = $signed({1'h0, smod_37885[15:0]}) < $signed({1'h0, sel_37946}) ? smod_37885[15:0] : sel_37946;
  assign umul_38141 = umul23b_16b_x_7b(array_index_37607, 7'h47);
  assign add_38143 = {1'h0, umul_37947[22:1]} + 23'h00_1f8b;
  assign sel_38148 = $signed({1'h0, smod_37890[15:0]}) < $signed({1'h0, sel_37954}) ? smod_37890[15:0] : sel_37954;
  assign umul_38149 = umul23b_16b_x_7b(array_index_37613, 7'h47);
  assign add_38151 = {1'h0, umul_37955[22:1]} + 23'h00_1f8b;
  assign sel_38156 = $signed({1'h0, smod_37895[15:0]}) < $signed({1'h0, sel_37962}) ? smod_37895[15:0] : sel_37962;
  assign umul_38157 = umul22b_16b_x_6b(array_index_37801, 6'h3d);
  assign add_38159 = {1'h0, umul_37963[21:2]} + 21'h00_0fb9;
  assign sel_38164 = $signed({1'h0, smod_37900[15:0]}) < $signed({1'h0, sel_37970}) ? smod_37900[15:0] : sel_37970;
  assign umul_38165 = umul22b_16b_x_6b(array_index_37807, 6'h3d);
  assign add_38167 = {1'h0, umul_37971[21:2]} + 21'h00_0fb9;
  assign sel_38172 = $signed({1'h0, smod_37905[15:0]}) < $signed({1'h0, sel_37978}) ? smod_37905[15:0] : sel_37978;
  assign umul_38173 = umul22b_16b_x_6b(array_index_37995, 6'h3b);
  assign add_38175 = {1'h0, umul_37979[21:1]} + 22'h00_1f59;
  assign sel_38180 = $signed({1'h0, smod_37910[15:0]}) < $signed({1'h0, sel_37986}) ? smod_37910[15:0] : sel_37986;
  assign umul_38181 = umul22b_16b_x_6b(array_index_38001, 6'h3b);
  assign add_38183 = {1'h0, umul_37987[21:1]} + 22'h00_1f59;
  assign sel_38188 = $signed({1'h0, smod_37915[15:0]}) < $signed({1'h0, sel_37994}) ? smod_37915[15:0] : sel_37994;
  assign array_index_38189 = set1_unflattened[5'h12];
  assign smod_38193 = $unsigned($signed({9'h000, add_38057, umul_37861[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_38195 = set2_unflattened[5'h12];
  assign smod_38199 = $unsigned($signed({9'h000, add_38065, umul_37869[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_38249 = umul22b_16b_x_6b(array_index_38189, 6'h35);
  assign add_38251 = {1'h0, umul_38055[21:7]} + 16'h007d;
  assign sel_38256 = $signed({1'h0, smod_37999[15:0]}) < $signed({1'h0, sel_38062}) ? smod_37999[15:0] : sel_38062;
  assign umul_38257 = umul22b_16b_x_6b(array_index_38195, 6'h35);
  assign add_38259 = {1'h0, umul_38063[21:7]} + 16'h007d;
  assign sel_38264 = $signed({1'h0, smod_38005[15:0]}) < $signed({1'h0, sel_38070}) ? smod_38005[15:0] : sel_38070;
  assign smod_38268 = $unsigned($signed({8'h00, add_38127, umul_37931[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38273 = $unsigned($signed({8'h00, add_38135, umul_37939[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38278 = $unsigned($signed({8'h00, add_38143, umul_37947[0]}) % $signed(32'h0000_3ffd));
  assign smod_38283 = $unsigned($signed({8'h00, add_38151, umul_37955[0]}) % $signed(32'h0000_3ffd));
  assign smod_38288 = $unsigned($signed({9'h000, add_38159, umul_37963[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_38293 = $unsigned($signed({9'h000, add_38167, umul_37971[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_38298 = $unsigned($signed({9'h000, add_38175, umul_37979[0]}) % $signed(32'h0000_3ffd));
  assign smod_38303 = $unsigned($signed({9'h000, add_38183, umul_37987[0]}) % $signed(32'h0000_3ffd));
  assign umul_38319 = umul23b_16b_x_7b(array_index_37607, 7'h49);
  assign add_38321 = {1'h0, umul_38125[22:3]} + 21'h00_07e9;
  assign sel_38326 = $signed({1'h0, smod_38074[15:0]}) < $signed({1'h0, sel_38132}) ? smod_38074[15:0] : sel_38132;
  assign umul_38327 = umul23b_16b_x_7b(array_index_37613, 7'h49);
  assign add_38329 = {1'h0, umul_38133[22:3]} + 21'h00_07e9;
  assign sel_38334 = $signed({1'h0, smod_38079[15:0]}) < $signed({1'h0, sel_38140}) ? smod_38079[15:0] : sel_38140;
  assign umul_38335 = umul23b_16b_x_7b(array_index_37801, 7'h47);
  assign add_38337 = {1'h0, umul_38141[22:1]} + 23'h00_1f8b;
  assign sel_38342 = $signed({1'h0, smod_38084[15:0]}) < $signed({1'h0, sel_38148}) ? smod_38084[15:0] : sel_38148;
  assign umul_38343 = umul23b_16b_x_7b(array_index_37807, 7'h47);
  assign add_38345 = {1'h0, umul_38149[22:1]} + 23'h00_1f8b;
  assign sel_38350 = $signed({1'h0, smod_38089[15:0]}) < $signed({1'h0, sel_38156}) ? smod_38089[15:0] : sel_38156;
  assign umul_38351 = umul22b_16b_x_6b(array_index_37995, 6'h3d);
  assign add_38353 = {1'h0, umul_38157[21:2]} + 21'h00_0fb9;
  assign sel_38358 = $signed({1'h0, smod_38094[15:0]}) < $signed({1'h0, sel_38164}) ? smod_38094[15:0] : sel_38164;
  assign umul_38359 = umul22b_16b_x_6b(array_index_38001, 6'h3d);
  assign add_38361 = {1'h0, umul_38165[21:2]} + 21'h00_0fb9;
  assign sel_38366 = $signed({1'h0, smod_38099[15:0]}) < $signed({1'h0, sel_38172}) ? smod_38099[15:0] : sel_38172;
  assign umul_38367 = umul22b_16b_x_6b(array_index_38189, 6'h3b);
  assign add_38369 = {1'h0, umul_38173[21:1]} + 22'h00_1f59;
  assign sel_38374 = $signed({1'h0, smod_38104[15:0]}) < $signed({1'h0, sel_38180}) ? smod_38104[15:0] : sel_38180;
  assign umul_38375 = umul22b_16b_x_6b(array_index_38195, 6'h3b);
  assign add_38377 = {1'h0, umul_38181[21:1]} + 22'h00_1f59;
  assign sel_38382 = $signed({1'h0, smod_38109[15:0]}) < $signed({1'h0, sel_38188}) ? smod_38109[15:0] : sel_38188;
  assign array_index_38383 = set1_unflattened[5'h13];
  assign smod_38387 = $unsigned($signed({9'h000, add_38251, umul_38055[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_38389 = set2_unflattened[5'h13];
  assign smod_38393 = $unsigned($signed({9'h000, add_38259, umul_38063[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_38443 = umul22b_16b_x_6b(array_index_38383, 6'h35);
  assign add_38445 = {1'h0, umul_38249[21:7]} + 16'h007d;
  assign sel_38450 = $signed({1'h0, smod_38193[15:0]}) < $signed({1'h0, sel_38256}) ? smod_38193[15:0] : sel_38256;
  assign umul_38451 = umul22b_16b_x_6b(array_index_38389, 6'h35);
  assign add_38453 = {1'h0, umul_38257[21:7]} + 16'h007d;
  assign sel_38458 = $signed({1'h0, smod_38199[15:0]}) < $signed({1'h0, sel_38264}) ? smod_38199[15:0] : sel_38264;
  assign smod_38462 = $unsigned($signed({8'h00, add_38321, umul_38125[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38467 = $unsigned($signed({8'h00, add_38329, umul_38133[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38472 = $unsigned($signed({8'h00, add_38337, umul_38141[0]}) % $signed(32'h0000_3ffd));
  assign smod_38477 = $unsigned($signed({8'h00, add_38345, umul_38149[0]}) % $signed(32'h0000_3ffd));
  assign smod_38482 = $unsigned($signed({9'h000, add_38353, umul_38157[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_38487 = $unsigned($signed({9'h000, add_38361, umul_38165[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_38492 = $unsigned($signed({9'h000, add_38369, umul_38173[0]}) % $signed(32'h0000_3ffd));
  assign smod_38497 = $unsigned($signed({9'h000, add_38377, umul_38181[0]}) % $signed(32'h0000_3ffd));
  assign umul_38511 = umul23b_16b_x_7b(array_index_37801, 7'h49);
  assign add_38513 = {1'h0, umul_38319[22:3]} + 21'h00_07e9;
  assign sel_38518 = $signed({1'h0, smod_38268[15:0]}) < $signed({1'h0, sel_38326}) ? smod_38268[15:0] : sel_38326;
  assign umul_38519 = umul23b_16b_x_7b(array_index_37807, 7'h49);
  assign add_38521 = {1'h0, umul_38327[22:3]} + 21'h00_07e9;
  assign sel_38526 = $signed({1'h0, smod_38273[15:0]}) < $signed({1'h0, sel_38334}) ? smod_38273[15:0] : sel_38334;
  assign umul_38527 = umul23b_16b_x_7b(array_index_37995, 7'h47);
  assign add_38529 = {1'h0, umul_38335[22:1]} + 23'h00_1f8b;
  assign sel_38534 = $signed({1'h0, smod_38278[15:0]}) < $signed({1'h0, sel_38342}) ? smod_38278[15:0] : sel_38342;
  assign umul_38535 = umul23b_16b_x_7b(array_index_38001, 7'h47);
  assign add_38537 = {1'h0, umul_38343[22:1]} + 23'h00_1f8b;
  assign sel_38542 = $signed({1'h0, smod_38283[15:0]}) < $signed({1'h0, sel_38350}) ? smod_38283[15:0] : sel_38350;
  assign umul_38543 = umul22b_16b_x_6b(array_index_38189, 6'h3d);
  assign add_38545 = {1'h0, umul_38351[21:2]} + 21'h00_0fb9;
  assign sel_38550 = $signed({1'h0, smod_38288[15:0]}) < $signed({1'h0, sel_38358}) ? smod_38288[15:0] : sel_38358;
  assign umul_38551 = umul22b_16b_x_6b(array_index_38195, 6'h3d);
  assign add_38553 = {1'h0, umul_38359[21:2]} + 21'h00_0fb9;
  assign sel_38558 = $signed({1'h0, smod_38293[15:0]}) < $signed({1'h0, sel_38366}) ? smod_38293[15:0] : sel_38366;
  assign umul_38559 = umul22b_16b_x_6b(array_index_38383, 6'h3b);
  assign add_38561 = {1'h0, umul_38367[21:1]} + 22'h00_1f59;
  assign sel_38566 = $signed({1'h0, smod_38298[15:0]}) < $signed({1'h0, sel_38374}) ? smod_38298[15:0] : sel_38374;
  assign umul_38567 = umul22b_16b_x_6b(array_index_38389, 6'h3b);
  assign add_38569 = {1'h0, umul_38375[21:1]} + 22'h00_1f59;
  assign sel_38574 = $signed({1'h0, smod_38303[15:0]}) < $signed({1'h0, sel_38382}) ? smod_38303[15:0] : sel_38382;
  assign smod_38577 = $unsigned($signed({9'h000, add_38445, umul_38249[6:0]}) % $signed(32'h0000_3ffd));
  assign smod_38581 = $unsigned($signed({9'h000, add_38453, umul_38257[6:0]}) % $signed(32'h0000_3ffd));
  assign add_38632 = {1'h0, umul_38443[21:7]} + 16'h007d;
  assign sel_38637 = $signed({1'h0, smod_38387[15:0]}) < $signed({1'h0, sel_38450}) ? smod_38387[15:0] : sel_38450;
  assign add_38639 = {1'h0, umul_38451[21:7]} + 16'h007d;
  assign sel_38644 = $signed({1'h0, smod_38393[15:0]}) < $signed({1'h0, sel_38458}) ? smod_38393[15:0] : sel_38458;
  assign smod_38648 = $unsigned($signed({8'h00, add_38513, umul_38319[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38653 = $unsigned($signed({8'h00, add_38521, umul_38327[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38658 = $unsigned($signed({8'h00, add_38529, umul_38335[0]}) % $signed(32'h0000_3ffd));
  assign smod_38663 = $unsigned($signed({8'h00, add_38537, umul_38343[0]}) % $signed(32'h0000_3ffd));
  assign smod_38668 = $unsigned($signed({9'h000, add_38545, umul_38351[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_38673 = $unsigned($signed({9'h000, add_38553, umul_38359[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_38677 = $unsigned($signed({9'h000, add_38561, umul_38367[0]}) % $signed(32'h0000_3ffd));
  assign smod_38681 = $unsigned($signed({9'h000, add_38569, umul_38375[0]}) % $signed(32'h0000_3ffd));
  assign umul_38691 = umul23b_16b_x_7b(array_index_37995, 7'h49);
  assign add_38693 = {1'h0, umul_38511[22:3]} + 21'h00_07e9;
  assign sel_38698 = $signed({1'h0, smod_38462[15:0]}) < $signed({1'h0, sel_38518}) ? smod_38462[15:0] : sel_38518;
  assign umul_38699 = umul23b_16b_x_7b(array_index_38001, 7'h49);
  assign add_38701 = {1'h0, umul_38519[22:3]} + 21'h00_07e9;
  assign sel_38706 = $signed({1'h0, smod_38467[15:0]}) < $signed({1'h0, sel_38526}) ? smod_38467[15:0] : sel_38526;
  assign umul_38707 = umul23b_16b_x_7b(array_index_38189, 7'h47);
  assign add_38709 = {1'h0, umul_38527[22:1]} + 23'h00_1f8b;
  assign sel_38714 = $signed({1'h0, smod_38472[15:0]}) < $signed({1'h0, sel_38534}) ? smod_38472[15:0] : sel_38534;
  assign umul_38715 = umul23b_16b_x_7b(array_index_38195, 7'h47);
  assign add_38717 = {1'h0, umul_38535[22:1]} + 23'h00_1f8b;
  assign sel_38722 = $signed({1'h0, smod_38477[15:0]}) < $signed({1'h0, sel_38542}) ? smod_38477[15:0] : sel_38542;
  assign umul_38723 = umul22b_16b_x_6b(array_index_38383, 6'h3d);
  assign add_38725 = {1'h0, umul_38543[21:2]} + 21'h00_0fb9;
  assign sel_38730 = $signed({1'h0, smod_38482[15:0]}) < $signed({1'h0, sel_38550}) ? smod_38482[15:0] : sel_38550;
  assign umul_38731 = umul22b_16b_x_6b(array_index_38389, 6'h3d);
  assign add_38733 = {1'h0, umul_38551[21:2]} + 21'h00_0fb9;
  assign sel_38738 = $signed({1'h0, smod_38487[15:0]}) < $signed({1'h0, sel_38558}) ? smod_38487[15:0] : sel_38558;
  assign add_38740 = {1'h0, umul_38559[21:1]} + 22'h00_1f59;
  assign sel_38745 = $signed({1'h0, smod_38492[15:0]}) < $signed({1'h0, sel_38566}) ? smod_38492[15:0] : sel_38566;
  assign add_38747 = {1'h0, umul_38567[21:1]} + 22'h00_1f59;
  assign sel_38752 = $signed({1'h0, smod_38497[15:0]}) < $signed({1'h0, sel_38574}) ? smod_38497[15:0] : sel_38574;
  assign smod_38753 = $unsigned($signed({9'h000, add_38632, umul_38443[6:0]}) % $signed(32'h0000_3ffd));
  assign smod_38755 = $unsigned($signed({9'h000, add_38639, umul_38451[6:0]}) % $signed(32'h0000_3ffd));
  assign sel_38804 = $signed({1'h0, smod_38577[15:0]}) < $signed({1'h0, sel_38637}) ? smod_38577[15:0] : sel_38637;
  assign sel_38808 = $signed({1'h0, smod_38581[15:0]}) < $signed({1'h0, sel_38644}) ? smod_38581[15:0] : sel_38644;
  assign smod_38812 = $unsigned($signed({8'h00, add_38693, umul_38511[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38817 = $unsigned($signed({8'h00, add_38701, umul_38519[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38822 = $unsigned($signed({8'h00, add_38709, umul_38527[0]}) % $signed(32'h0000_3ffd));
  assign smod_38827 = $unsigned($signed({8'h00, add_38717, umul_38535[0]}) % $signed(32'h0000_3ffd));
  assign smod_38831 = $unsigned($signed({9'h000, add_38725, umul_38543[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_38835 = $unsigned($signed({9'h000, add_38733, umul_38551[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_38837 = $unsigned($signed({9'h000, add_38740, umul_38559[0]}) % $signed(32'h0000_3ffd));
  assign smod_38839 = $unsigned($signed({9'h000, add_38747, umul_38567[0]}) % $signed(32'h0000_3ffd));
  assign umul_38845 = umul23b_16b_x_7b(array_index_38189, 7'h49);
  assign add_38847 = {1'h0, umul_38691[22:3]} + 21'h00_07e9;
  assign sel_38852 = $signed({1'h0, smod_38648[15:0]}) < $signed({1'h0, sel_38698}) ? smod_38648[15:0] : sel_38698;
  assign umul_38853 = umul23b_16b_x_7b(array_index_38195, 7'h49);
  assign add_38855 = {1'h0, umul_38699[22:3]} + 21'h00_07e9;
  assign sel_38860 = $signed({1'h0, smod_38653[15:0]}) < $signed({1'h0, sel_38706}) ? smod_38653[15:0] : sel_38706;
  assign umul_38861 = umul23b_16b_x_7b(array_index_38383, 7'h47);
  assign add_38863 = {1'h0, umul_38707[22:1]} + 23'h00_1f8b;
  assign sel_38868 = $signed({1'h0, smod_38658[15:0]}) < $signed({1'h0, sel_38714}) ? smod_38658[15:0] : sel_38714;
  assign umul_38869 = umul23b_16b_x_7b(array_index_38389, 7'h47);
  assign add_38871 = {1'h0, umul_38715[22:1]} + 23'h00_1f8b;
  assign sel_38876 = $signed({1'h0, smod_38663[15:0]}) < $signed({1'h0, sel_38722}) ? smod_38663[15:0] : sel_38722;
  assign add_38878 = {1'h0, umul_38723[21:2]} + 21'h00_0fb9;
  assign sel_38883 = $signed({1'h0, smod_38668[15:0]}) < $signed({1'h0, sel_38730}) ? smod_38668[15:0] : sel_38730;
  assign add_38885 = {1'h0, umul_38731[21:2]} + 21'h00_0fb9;
  assign sel_38890 = $signed({1'h0, smod_38673[15:0]}) < $signed({1'h0, sel_38738}) ? smod_38673[15:0] : sel_38738;
  assign sel_38894 = $signed({1'h0, smod_38677[15:0]}) < $signed({1'h0, sel_38745}) ? smod_38677[15:0] : sel_38745;
  assign sel_38898 = $signed({1'h0, smod_38681[15:0]}) < $signed({1'h0, sel_38752}) ? smod_38681[15:0] : sel_38752;
  assign smod_38942 = $unsigned($signed({8'h00, add_38847, umul_38691[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38947 = $unsigned($signed({8'h00, add_38855, umul_38699[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_38951 = $unsigned($signed({8'h00, add_38863, umul_38707[0]}) % $signed(32'h0000_3ffd));
  assign smod_38955 = $unsigned($signed({8'h00, add_38871, umul_38715[0]}) % $signed(32'h0000_3ffd));
  assign smod_38957 = $unsigned($signed({9'h000, add_38878, umul_38723[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_38959 = $unsigned($signed({9'h000, add_38885, umul_38731[1:0]}) % $signed(32'h0000_3ffd));
  assign umul_38965 = umul23b_16b_x_7b(array_index_38383, 7'h49);
  assign add_38967 = {1'h0, umul_38845[22:3]} + 21'h00_07e9;
  assign sel_38972 = $signed({1'h0, smod_38812[15:0]}) < $signed({1'h0, sel_38852}) ? smod_38812[15:0] : sel_38852;
  assign umul_38973 = umul23b_16b_x_7b(array_index_38389, 7'h49);
  assign add_38975 = {1'h0, umul_38853[22:3]} + 21'h00_07e9;
  assign sel_38980 = $signed({1'h0, smod_38817[15:0]}) < $signed({1'h0, sel_38860}) ? smod_38817[15:0] : sel_38860;
  assign add_38982 = {1'h0, umul_38861[22:1]} + 23'h00_1f8b;
  assign sel_38987 = $signed({1'h0, smod_38822[15:0]}) < $signed({1'h0, sel_38868}) ? smod_38822[15:0] : sel_38868;
  assign add_38989 = {1'h0, umul_38869[22:1]} + 23'h00_1f8b;
  assign sel_38994 = $signed({1'h0, smod_38827[15:0]}) < $signed({1'h0, sel_38876}) ? smod_38827[15:0] : sel_38876;
  assign sel_38998 = $signed({1'h0, smod_38831[15:0]}) < $signed({1'h0, sel_38883}) ? smod_38831[15:0] : sel_38883;
  assign sel_39002 = $signed({1'h0, smod_38835[15:0]}) < $signed({1'h0, sel_38890}) ? smod_38835[15:0] : sel_38890;
  assign concat_39005 = {1'h0, ($signed({1'h0, smod_38753[15:0]}) < $signed({1'h0, sel_38804}) ? smod_38753[15:0] : sel_38804) == ($signed({1'h0, smod_38755[15:0]}) < $signed({1'h0, sel_38808}) ? smod_38755[15:0] : sel_38808)};
  assign add_39032 = concat_39005 + 2'h1;
  assign smod_39035 = $unsigned($signed({8'h00, add_38967, umul_38845[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_39039 = $unsigned($signed({8'h00, add_38975, umul_38853[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_39041 = $unsigned($signed({8'h00, add_38982, umul_38861[0]}) % $signed(32'h0000_3ffd));
  assign smod_39043 = $unsigned($signed({8'h00, add_38989, umul_38869[0]}) % $signed(32'h0000_3ffd));
  assign add_39050 = {1'h0, umul_38965[22:3]} + 21'h00_07e9;
  assign sel_39055 = $signed({1'h0, smod_38942[15:0]}) < $signed({1'h0, sel_38972}) ? smod_38942[15:0] : sel_38972;
  assign add_39057 = {1'h0, umul_38973[22:3]} + 21'h00_07e9;
  assign sel_39062 = $signed({1'h0, smod_38947[15:0]}) < $signed({1'h0, sel_38980}) ? smod_38947[15:0] : sel_38980;
  assign sel_39066 = $signed({1'h0, smod_38951[15:0]}) < $signed({1'h0, sel_38987}) ? smod_38951[15:0] : sel_38987;
  assign sel_39070 = $signed({1'h0, smod_38955[15:0]}) < $signed({1'h0, sel_38994}) ? smod_38955[15:0] : sel_38994;
  assign concat_39073 = {1'h0, ($signed({1'h0, smod_38837[15:0]}) < $signed({1'h0, sel_38894}) ? smod_38837[15:0] : sel_38894) == ($signed({1'h0, smod_38839[15:0]}) < $signed({1'h0, sel_38898}) ? smod_38839[15:0] : sel_38898) ? add_39032 : concat_39005};
  assign add_39088 = concat_39073 + 3'h1;
  assign smod_39089 = $unsigned($signed({8'h00, add_39050, umul_38965[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_39091 = $unsigned($signed({8'h00, add_39057, umul_38973[2:0]}) % $signed(32'h0000_3ffd));
  assign sel_39100 = $signed({1'h0, smod_39035[15:0]}) < $signed({1'h0, sel_39055}) ? smod_39035[15:0] : sel_39055;
  assign sel_39104 = $signed({1'h0, smod_39039[15:0]}) < $signed({1'h0, sel_39062}) ? smod_39039[15:0] : sel_39062;
  assign concat_39107 = {1'h0, ($signed({1'h0, smod_38957[15:0]}) < $signed({1'h0, sel_38998}) ? smod_38957[15:0] : sel_38998) == ($signed({1'h0, smod_38959[15:0]}) < $signed({1'h0, sel_39002}) ? smod_38959[15:0] : sel_39002) ? add_39088 : concat_39073};
  assign add_39114 = concat_39107 + 4'h1;
  assign concat_39121 = {1'h0, ($signed({1'h0, smod_39041[15:0]}) < $signed({1'h0, sel_39066}) ? smod_39041[15:0] : sel_39066) == ($signed({1'h0, smod_39043[15:0]}) < $signed({1'h0, sel_39070}) ? smod_39043[15:0] : sel_39070) ? add_39114 : concat_39107};
  assign add_39124 = concat_39121 + 5'h01;
  assign out = {{11'h000, ($signed({1'h0, smod_39089[15:0]}) < $signed({1'h0, sel_39100}) ? smod_39089[15:0] : sel_39100) == ($signed({1'h0, smod_39091[15:0]}) < $signed({1'h0, sel_39104}) ? smod_39091[15:0] : sel_39104) ? add_39124 : concat_39121}, {set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
