module min_hash(set1, set2, out);
  wire _00000_, _00001_, _00002_, _00003_, _00004_, _00005_, _00006_, _00007_, _00008_, _00009_, _00010_, _00011_, _00012_, _00013_, _00014_, _00015_, _00016_, _00017_, _00018_, _00019_, _00020_, _00021_, _00022_, _00023_, _00024_, _00025_, _00026_, _00027_, _00028_, _00029_, _00030_, _00031_, _00032_, _00033_, _00034_, _00035_, _00036_, _00037_, _00038_, _00039_, _00040_, _00041_, _00042_, _00043_, _00044_, _00045_, _00046_, _00047_, _00048_, _00049_, _00050_, _00051_, _00052_, _00053_, _00054_, _00055_, _00056_, _00057_, _00058_, _00059_, _00060_, _00061_, _00062_, _00063_, _00064_, _00065_, _00066_, _00067_, _00068_, _00069_, _00070_, _00071_, _00072_, _00073_, _00074_, _00075_, _00076_, _00077_, _00078_, _00079_, _00080_, _00081_, _00082_, _00083_, _00084_, _00085_, _00086_, _00087_, _00088_, _00089_, _00090_, _00091_, _00092_, _00093_, _00094_, _00095_, _00096_, _00097_, _00098_, _00099_, _00100_, _00101_, _00102_, _00103_, _00104_, _00105_, _00106_, _00107_, _00108_, _00109_, _00110_, _00111_, _00112_, _00113_, _00114_, _00115_, _00116_, _00117_, _00118_, _00119_, _00120_, _00121_, _00122_, _00123_, _00124_, _00125_, _00126_, _00127_, _00128_, _00129_, _00130_, _00131_, _00132_, _00133_, _00134_, _00135_, _00136_, _00137_, _00138_, _00139_, _00140_, _00141_, _00142_, _00143_, _00144_, _00145_, _00146_, _00147_, _00148_, _00149_, _00150_, _00151_, _00152_, _00153_, _00154_, _00155_, _00156_, _00157_, _00158_, _00159_, _00160_, _00161_, _00162_, _00163_, _00164_, _00165_, _00166_, _00167_, _00168_, _00169_, _00170_, _00171_, _00172_, _00173_, _00174_, _00175_, _00176_, _00177_, _00178_, _00179_, _00180_, _00181_, _00182_, _00183_, _00184_, _00185_, _00186_, _00187_, _00188_, _00189_, _00190_, _00191_, _00192_, _00193_, _00194_, _00195_, _00196_, _00197_, _00198_, _00199_, _00200_, _00201_, _00202_, _00203_, _00204_, _00205_, _00206_, _00207_, _00208_, _00209_, _00210_, _00211_, _00212_, _00213_, _00214_, _00215_, _00216_, _00217_, _00218_, _00219_, _00220_, _00221_, _00222_, _00223_, _00224_, _00225_, _00226_, _00227_, _00228_, _00229_, _00230_, _00231_, _00232_, _00233_, _00234_, _00235_, _00236_, _00237_, _00238_, _00239_, _00240_, _00241_, _00242_, _00243_, _00244_, _00245_, _00246_, _00247_, _00248_, _00249_, _00250_, _00251_, _00252_, _00253_, _00254_, _00255_, _00256_, _00257_, _00258_, _00259_, _00260_, _00261_, _00262_, _00263_, _00264_, _00265_, _00266_, _00267_, _00268_, _00269_, _00270_, _00271_, _00272_, _00273_, _00274_, _00275_, _00276_, _00277_, _00278_, _00279_, _00280_, _00281_, _00282_, _00283_, _00284_, _00285_, _00286_, _00287_, _00288_, _00289_, _00290_, _00291_, _00292_, _00293_, _00294_, _00295_, _00296_, _00297_, _00298_, _00299_, _00300_, _00301_, _00302_, _00303_, _00304_, _00305_, _00306_, _00307_, _00308_, _00309_, _00310_, _00311_, _00312_, _00313_, _00314_, _00315_, _00316_, _00317_, _00318_, _00319_, _00320_, _00321_, _00322_, _00323_, _00324_, _00325_, _00326_, _00327_, _00328_, _00329_, _00330_, _00331_, _00332_, _00333_, _00334_, _00335_, _00336_, _00337_, _00338_, _00339_, _00340_, _00341_, _00342_, _00343_, _00344_, _00345_, _00346_, _00347_, _00348_, _00349_, _00350_, _00351_, _00352_, _00353_, _00354_, _00355_, _00356_, _00357_, _00358_, _00359_, _00360_, _00361_, _00362_, _00363_, _00364_, _00365_, _00366_, _00367_, _00368_, _00369_, _00370_, _00371_, _00372_, _00373_, _00374_, _00375_, _00376_, _00377_, _00378_, _00379_, _00380_, _00381_, _00382_, _00383_, _00384_, _00385_, _00386_, _00387_, _00388_, _00389_, _00390_, _00391_, _00392_, _00393_, _00394_, _00395_, _00396_, _00397_, _00398_, _00399_, _00400_, _00401_, _00402_, _00403_, _00404_, _00405_, _00406_, _00407_, _00408_, _00409_, _00410_, _00411_, _00412_, _00413_, _00414_, _00415_, _00416_, _00417_, _00418_, _00419_, _00420_, _00421_, _00422_, _00423_, _00424_, _00425_, _00426_, _00427_, _00428_, _00429_, _00430_, _00431_, _00432_, _00433_, _00434_, _00435_, _00436_, _00437_, _00438_, _00439_, _00440_, _00441_, _00442_, _00443_, _00444_, _00445_, _00446_, _00447_, _00448_, _00449_, _00450_, _00451_, _00452_, _00453_, _00454_, _00455_, _00456_, _00457_, _00458_, _00459_, _00460_, _00461_, _00462_, _00463_, _00464_, _00465_, _00466_, _00467_, _00468_, _00469_, _00470_, _00471_, _00472_, _00473_, _00474_, _00475_, _00476_, _00477_, _00478_, _00479_, _00480_, _00481_, _00482_, _00483_, _00484_, _00485_, _00486_, _00487_, _00488_, _00489_, _00490_, _00491_, _00492_, _00493_, _00494_, _00495_, _00496_, _00497_, _00498_, _00499_, _00500_, _00501_, _00502_, _00503_, _00504_, _00505_, _00506_, _00507_, _00508_, _00509_, _00510_, _00511_, _00512_, _00513_, _00514_, _00515_, _00516_, _00517_, _00518_, _00519_, _00520_, _00521_, _00522_, _00523_, _00524_, _00525_, _00526_, _00527_, _00528_, _00529_, _00530_, _00531_, _00532_, _00533_, _00534_, _00535_, _00536_, _00537_, _00538_, _00539_, _00540_, _00541_, _00542_, _00543_, _00544_, _00545_, _00546_, _00547_, _00548_, _00549_, _00550_, _00551_, _00552_, _00553_, _00554_, _00555_, _00556_, _00557_, _00558_, _00559_, _00560_, _00561_, _00562_, _00563_, _00564_, _00565_, _00566_, _00567_, _00568_, _00569_, _00570_, _00571_, _00572_, _00573_, _00574_, _00575_, _00576_, _00577_, _00578_, _00579_, _00580_, _00581_, _00582_, _00583_, _00584_, _00585_, _00586_, _00587_, _00588_, _00589_, _00590_, _00591_, _00592_, _00593_, _00594_, _00595_, _00596_, _00597_, _00598_, _00599_, _00600_, _00601_, _00602_, _00603_, _00604_, _00605_, _00606_, _00607_, _00608_, _00609_, _00610_, _00611_, _00612_, _00613_, _00614_, _00615_, _00616_, _00617_, _00618_, _00619_, _00620_, _00621_, _00622_, _00623_, _00624_, _00625_, _00626_, _00627_, _00628_, _00629_, _00630_, _00631_, _00632_, _00633_, _00634_, _00635_, _00636_, _00637_, _00638_, _00639_, _00640_, _00641_, _00642_, _00643_, _00644_, _00645_, _00646_, _00647_, _00648_, _00649_, _00650_, _00651_, _00652_, _00653_, _00654_, _00655_, _00656_, _00657_, _00658_, _00659_, _00660_, _00661_, _00662_, _00663_, _00664_, _00665_, _00666_, _00667_, _00668_, _00669_, _00670_, _00671_, _00672_, _00673_, _00674_, _00675_, _00676_, _00677_, _00678_, _00679_, _00680_, _00681_, _00682_, _00683_, _00684_, _00685_, _00686_, _00687_, _00688_, _00689_, _00690_, _00691_, _00692_, _00693_, _00694_, _00695_, _00696_, _00697_, _00698_, _00699_, _00700_, _00701_, _00702_, _00703_, _00704_, _00705_, _00706_, _00707_, _00708_, _00709_, _00710_, _00711_, _00712_, _00713_, _00714_, _00715_, _00716_, _00717_, _00718_, _00719_, _00720_, _00721_, _00722_, _00723_, _00724_, _00725_, _00726_, _00727_, _00728_, _00729_, _00730_, _00731_, _00732_, _00733_, _00734_, _00735_, _00736_, _00737_, _00738_, _00739_, _00740_, _00741_, _00742_, _00743_, _00744_, _00745_, _00746_, _00747_, _00748_, _00749_, _00750_, _00751_, _00752_, _00753_, _00754_, _00755_, _00756_, _00757_, _00758_, _00759_, _00760_, _00761_, _00762_, _00763_, _00764_, _00765_, _00766_, _00767_, _00768_, _00769_, _00770_, _00771_, _00772_, _00773_, _00774_, _00775_, _00776_, _00777_, _00778_, _00779_, _00780_, _00781_, _00782_, _00783_, _00784_, _00785_, _00786_, _00787_, _00788_, _00789_, _00790_, _00791_, _00792_, _00793_, _00794_, _00795_, _00796_, _00797_, _00798_, _00799_, _00800_, _00801_, _00802_, _00803_, _00804_, _00805_, _00806_, _00807_, _00808_, _00809_, _00810_, _00811_, _00812_, _00813_, _00814_, _00815_, _00816_, _00817_, _00818_, _00819_, _00820_, _00821_, _00822_, _00823_, _00824_, _00825_, _00826_, _00827_, _00828_, _00829_, _00830_, _00831_, _00832_, _00833_, _00834_, _00835_, _00836_, _00837_, _00838_, _00839_, _00840_, _00841_, _00842_, _00843_, _00844_, _00845_, _00846_, _00847_, _00848_, _00849_, _00850_, _00851_, _00852_, _00853_, _00854_, _00855_, _00856_, _00857_, _00858_, _00859_, _00860_, _00861_, _00862_, _00863_, _00864_, _00865_, _00866_, _00867_, _00868_, _00869_, _00870_, _00871_, _00872_, _00873_, _00874_, _00875_, _00876_, _00877_, _00878_, _00879_, _00880_, _00881_, _00882_, _00883_, _00884_, _00885_, _00886_, _00887_, _00888_, _00889_, _00890_, _00891_, _00892_, _00893_, _00894_, _00895_, _00896_, _00897_, _00898_, _00899_, _00900_, _00901_, _00902_, _00903_, _00904_, _00905_, _00906_, _00907_, _00908_, _00909_, _00910_, _00911_, _00912_, _00913_, _00914_, _00915_, _00916_, _00917_, _00918_, _00919_, _00920_, _00921_, _00922_, _00923_, _00924_, _00925_, _00926_, _00927_, _00928_, _00929_, _00930_, _00931_, _00932_, _00933_, _00934_, _00935_, _00936_, _00937_, _00938_, _00939_, _00940_, _00941_, _00942_, _00943_, _00944_, _00945_, _00946_, _00947_, _00948_, _00949_, _00950_, _00951_, _00952_, _00953_, _00954_, _00955_, _00956_, _00957_, _00958_, _00959_, _00960_, _00961_, _00962_, _00963_, _00964_, _00965_, _00966_, _00967_, _00968_, _00969_, _00970_, _00971_, _00972_, _00973_, _00974_, _00975_, _00976_, _00977_, _00978_, _00979_, _00980_, _00981_, _00982_, _00983_, _00984_, _00985_, _00986_, _00987_, _00988_, _00989_, _00990_, _00991_, _00992_, _00993_, _00994_, _00995_, _00996_, _00997_, _00998_, _00999_, _01000_, _01001_, _01002_, _01003_, _01004_, _01005_, _01006_, _01007_, _01008_, _01009_, _01010_, _01011_, _01012_, _01013_, _01014_, _01015_, _01016_, _01017_, _01018_, _01019_, _01020_, _01021_, _01022_, _01023_, _01024_, _01025_, _01026_, _01027_, _01028_, _01029_, _01030_, _01031_, _01032_, _01033_, _01034_, _01035_, _01036_, _01037_, _01038_, _01039_, _01040_, _01041_, _01042_, _01043_, _01044_, _01045_, _01046_, _01047_, _01048_, _01049_, _01050_, _01051_, _01052_, _01053_, _01054_, _01055_, _01056_, _01057_, _01058_, _01059_, _01060_, _01061_, _01062_, _01063_, _01064_, _01065_, _01066_, _01067_, _01068_, _01069_, _01070_, _01071_, _01072_, _01073_, _01074_, _01075_, _01076_, _01077_, _01078_, _01079_, _01080_, _01081_, _01082_, _01083_, _01084_, _01085_, _01086_, _01087_, _01088_, _01089_, _01090_, _01091_, _01092_, _01093_, _01094_, _01095_, _01096_, _01097_, _01098_, _01099_, _01100_, _01101_, _01102_, _01103_, _01104_, _01105_, _01106_, _01107_, _01108_, _01109_, _01110_, _01111_, _01112_, _01113_, _01114_, _01115_, _01116_, _01117_, _01118_, _01119_, _01120_, _01121_, _01122_, _01123_, _01124_, _01125_, _01126_, _01127_, _01128_, _01129_, _01130_, _01131_, _01132_, _01133_, _01134_, _01135_, _01136_, _01137_, _01138_, _01139_, _01140_, _01141_, _01142_, _01143_, _01144_, _01145_, _01146_, _01147_, _01148_, _01149_, _01150_, _01151_, _01152_, _01153_, _01154_, _01155_, _01156_, _01157_, _01158_, _01159_, _01160_, _01161_, _01162_, _01163_, _01164_, _01165_, _01166_, _01167_, _01168_, _01169_, _01170_, _01171_, _01172_, _01173_, _01174_, _01175_, _01176_, _01177_, _01178_, _01179_, _01180_, _01181_, _01182_, _01183_, _01184_, _01185_, _01186_, _01187_, _01188_, _01189_, _01190_, _01191_, _01192_, _01193_, _01194_, _01195_, _01196_, _01197_, _01198_, _01199_, _01200_, _01201_, _01202_, _01203_, _01204_, _01205_, _01206_, _01207_, _01208_, _01209_, _01210_, _01211_, _01212_, _01213_, _01214_, _01215_, _01216_, _01217_, _01218_, _01219_, _01220_, _01221_, _01222_, _01223_, _01224_, _01225_, _01226_, _01227_, _01228_, _01229_, _01230_, _01231_, _01232_, _01233_, _01234_, _01235_, _01236_, _01237_, _01238_, _01239_, _01240_, _01241_, _01242_, _01243_, _01244_, _01245_, _01246_, _01247_, _01248_, _01249_, _01250_, _01251_, _01252_, _01253_, _01254_, _01255_, _01256_, _01257_, _01258_, _01259_, _01260_, _01261_, _01262_, _01263_, _01264_, _01265_, _01266_, _01267_, _01268_, _01269_, _01270_, _01271_, _01272_, _01273_, _01274_, _01275_, _01276_, _01277_, _01278_, _01279_, _01280_, _01281_, _01282_, _01283_, _01284_, _01285_, _01286_, _01287_, _01288_, _01289_, _01290_, _01291_, _01292_, _01293_, _01294_, _01295_, _01296_, _01297_, _01298_, _01299_, _01300_, _01301_, _01302_, _01303_, _01304_, _01305_, _01306_, _01307_, _01308_, _01309_, _01310_, _01311_, _01312_, _01313_, _01314_, _01315_, _01316_, _01317_, _01318_, _01319_, _01320_, _01321_, _01322_, _01323_, _01324_, _01325_, _01326_, _01327_, _01328_, _01329_, _01330_, _01331_, _01332_, _01333_, _01334_, _01335_, _01336_, _01337_, _01338_, _01339_, _01340_, _01341_, _01342_, _01343_, _01344_, _01345_, _01346_, _01347_, _01348_, _01349_, _01350_, _01351_, _01352_, _01353_, _01354_, _01355_, _01356_, _01357_, _01358_, _01359_, _01360_, _01361_, _01362_, _01363_, _01364_, _01365_, _01366_, _01367_, _01368_, _01369_, _01370_, _01371_, _01372_, _01373_, _01374_, _01375_, _01376_, _01377_, _01378_, _01379_, _01380_, _01381_, _01382_, _01383_, _01384_, _01385_, _01386_, _01387_, _01388_, _01389_, _01390_, _01391_, _01392_, _01393_, _01394_, _01395_, _01396_, _01397_, _01398_, _01399_, _01400_, _01401_, _01402_, _01403_, _01404_, _01405_, _01406_, _01407_, _01408_, _01409_, _01410_, _01411_, _01412_, _01413_, _01414_, _01415_, _01416_, _01417_, _01418_, _01419_, _01420_, _01421_, _01422_, _01423_, _01424_, _01425_, _01426_, _01427_, _01428_, _01429_, _01430_, _01431_, _01432_, _01433_, _01434_, _01435_, _01436_, _01437_, _01438_, _01439_, _01440_, _01441_, _01442_, _01443_, _01444_, _01445_, _01446_, _01447_, _01448_, _01449_, _01450_, _01451_, _01452_, _01453_, _01454_, _01455_, _01456_, _01457_, _01458_, _01459_, _01460_, _01461_, _01462_, _01463_, _01464_, _01465_, _01466_, _01467_, _01468_, _01469_, _01470_, _01471_, _01472_, _01473_, _01474_, _01475_, _01476_, _01477_, _01478_, _01479_, _01480_, _01481_, _01482_, _01483_, _01484_, _01485_, _01486_, _01487_, _01488_, _01489_, _01490_, _01491_, _01492_, _01493_, _01494_, _01495_, _01496_, _01497_, _01498_, _01499_, _01500_, _01501_, _01502_, _01503_, _01504_, _01505_, _01506_, _01507_, _01508_, _01509_, _01510_, _01511_, _01512_, _01513_, _01514_, _01515_, _01516_, _01517_, _01518_, _01519_, _01520_, _01521_, _01522_, _01523_, _01524_, _01525_, _01526_, _01527_, _01528_, _01529_, _01530_, _01531_, _01532_, _01533_, _01534_, _01535_, _01536_, _01537_, _01538_, _01539_, _01540_, _01541_, _01542_, _01543_, _01544_, _01545_, _01546_, _01547_, _01548_, _01549_, _01550_, _01551_, _01552_, _01553_, _01554_, _01555_, _01556_, _01557_, _01558_, _01559_, _01560_, _01561_, _01562_, _01563_, _01564_, _01565_, _01566_, _01567_, _01568_, _01569_, _01570_, _01571_, _01572_, _01573_, _01574_, _01575_, _01576_, _01577_, _01578_, _01579_, _01580_, _01581_, _01582_, _01583_, _01584_, _01585_, _01586_, _01587_, _01588_, _01589_, _01590_, _01591_, _01592_, _01593_, _01594_, _01595_, _01596_, _01597_, _01598_, _01599_, _01600_, _01601_, _01602_, _01603_, _01604_, _01605_, _01606_, _01607_, _01608_, _01609_, _01610_, _01611_, _01612_, _01613_, _01614_, _01615_, _01616_, _01617_, _01618_, _01619_, _01620_, _01621_, _01622_, _01623_, _01624_, _01625_, _01626_, _01627_, _01628_, _01629_, _01630_, _01631_, _01632_, _01633_, _01634_, _01635_, _01636_, _01637_, _01638_, _01639_, _01640_, _01641_, _01642_, _01643_, _01644_, _01645_, _01646_, _01647_, _01648_, _01649_, _01650_, _01651_, _01652_, _01653_, _01654_, _01655_, _01656_, _01657_, _01658_, _01659_, _01660_, _01661_, _01662_, _01663_, _01664_, _01665_, _01666_, _01667_, _01668_, _01669_, _01670_, _01671_, _01672_, _01673_, _01674_, _01675_, _01676_, _01677_, _01678_, _01679_, _01680_, _01681_, _01682_, _01683_, _01684_, _01685_, _01686_, _01687_, _01688_, _01689_, _01690_, _01691_, _01692_, _01693_, _01694_, _01695_, _01696_, _01697_, _01698_, _01699_, _01700_, _01701_, _01702_, _01703_, _01704_, _01705_, _01706_, _01707_, _01708_, _01709_, _01710_, _01711_, _01712_, _01713_, _01714_, _01715_, _01716_, _01717_, _01718_, _01719_, _01720_, _01721_, _01722_, _01723_, _01724_, _01725_, _01726_, _01727_, _01728_, _01729_, _01730_, _01731_, _01732_, _01733_, _01734_, _01735_, _01736_, _01737_, _01738_, _01739_, _01740_, _01741_, _01742_, _01743_, _01744_, _01745_, _01746_, _01747_, _01748_, _01749_, _01750_, _01751_, _01752_, _01753_, _01754_, _01755_, _01756_, _01757_, _01758_, _01759_, _01760_, _01761_, _01762_, _01763_, _01764_, _01765_, _01766_, _01767_, _01768_, _01769_, _01770_, _01771_, _01772_, _01773_, _01774_, _01775_, _01776_, _01777_, _01778_, _01779_, _01780_, _01781_, _01782_, _01783_, _01784_, _01785_, _01786_, _01787_, _01788_, _01789_, _01790_, _01791_, _01792_, _01793_, _01794_, _01795_, _01796_, _01797_, _01798_, _01799_, _01800_, _01801_, _01802_, _01803_, _01804_, _01805_, _01806_, _01807_, _01808_, _01809_, _01810_, _01811_, _01812_, _01813_, _01814_, _01815_, _01816_, _01817_, _01818_, _01819_, _01820_, _01821_, _01822_, _01823_, _01824_, _01825_, _01826_, _01827_, _01828_, _01829_, _01830_, _01831_, _01832_, _01833_, _01834_, _01835_, _01836_, _01837_, _01838_, _01839_, _01840_, _01841_, _01842_, _01843_, _01844_, _01845_, _01846_, _01847_, _01848_, _01849_, _01850_, _01851_, _01852_, _01853_, _01854_, _01855_, _01856_, _01857_, _01858_, _01859_, _01860_, _01861_, _01862_, _01863_, _01864_, _01865_, _01866_, _01867_, _01868_, _01869_, _01870_, _01871_, _01872_, _01873_, _01874_, _01875_, _01876_, _01877_, _01878_, _01879_, _01880_, _01881_, _01882_, _01883_, _01884_, _01885_, _01886_, _01887_, _01888_, _01889_, _01890_, _01891_, _01892_, _01893_, _01894_, _01895_, _01896_, _01897_, _01898_, _01899_, _01900_, _01901_, _01902_, _01903_, _01904_, _01905_, _01906_, _01907_, _01908_, _01909_, _01910_, _01911_, _01912_, _01913_, _01914_, _01915_, _01916_, _01917_, _01918_, _01919_, _01920_, _01921_, _01922_, _01923_, _01924_, _01925_, _01926_, _01927_, _01928_, _01929_, _01930_, _01931_, _01932_, _01933_, _01934_, _01935_, _01936_, _01937_, _01938_, _01939_, _01940_, _01941_, _01942_, _01943_, _01944_, _01945_, _01946_, _01947_, _01948_, _01949_, _01950_, _01951_, _01952_, _01953_, _01954_, _01955_, _01956_, _01957_, _01958_, _01959_, _01960_, _01961_, _01962_, _01963_, _01964_, _01965_, _01966_, _01967_, _01968_, _01969_, _01970_, _01971_, _01972_, _01973_, _01974_, _01975_, _01976_, _01977_, _01978_, _01979_, _01980_, _01981_, _01982_, _01983_, _01984_, _01985_, _01986_, _01987_, _01988_, _01989_, _01990_, _01991_, _01992_, _01993_, _01994_, _01995_, _01996_, _01997_, _01998_, _01999_, _02000_, _02001_, _02002_, _02003_, _02004_, _02005_, _02006_, _02007_, _02008_, _02009_, _02010_, _02011_, _02012_, _02013_, _02014_, _02015_, _02016_, _02017_, _02018_, _02019_, _02020_, _02021_, _02022_, _02023_, _02024_, _02025_, _02026_, _02027_, _02028_, _02029_, _02030_, _02031_, _02032_, _02033_, _02034_, _02035_, _02036_, _02037_, _02038_, _02039_, _02040_, _02041_, _02042_, _02043_, _02044_, _02045_, _02046_, _02047_, _02048_, _02049_, _02050_, _02051_, _02052_, _02053_, _02054_, _02055_, _02056_, _02057_, _02058_, _02059_, _02060_, _02061_, _02062_, _02063_, _02064_, _02065_, _02066_, _02067_, _02068_, _02069_, _02070_, _02071_, _02072_, _02073_, _02074_, _02075_, _02076_, _02077_, _02078_, _02079_, _02080_, _02081_, _02082_, _02083_, _02084_, _02085_, _02086_, _02087_, _02088_, _02089_, _02090_, _02091_, _02092_, _02093_, _02094_, _02095_, _02096_, _02097_, _02098_, _02099_, _02100_, _02101_, _02102_, _02103_, _02104_, _02105_, _02106_, _02107_, _02108_, _02109_, _02110_, _02111_, _02112_, _02113_, _02114_, _02115_, _02116_, _02117_, _02118_, _02119_, _02120_, _02121_, _02122_, _02123_, _02124_, _02125_, _02126_, _02127_, _02128_, _02129_, _02130_, _02131_, _02132_, _02133_, _02134_, _02135_, _02136_, _02137_, _02138_, _02139_, _02140_, _02141_, _02142_, _02143_, _02144_, _02145_, _02146_, _02147_, _02148_, _02149_, _02150_, _02151_, _02152_, _02153_, _02154_, _02155_, _02156_, _02157_, _02158_, _02159_, _02160_, _02161_, _02162_, _02163_, _02164_, _02165_, _02166_, _02167_, _02168_, _02169_, _02170_, _02171_, _02172_, _02173_, _02174_, _02175_, _02176_, _02177_, _02178_, _02179_, _02180_, _02181_, _02182_, _02183_, _02184_, _02185_, _02186_, _02187_, _02188_, _02189_, _02190_, _02191_, _02192_, _02193_, _02194_, _02195_, _02196_, _02197_, _02198_, _02199_, _02200_, _02201_, _02202_, _02203_, _02204_, _02205_, _02206_, _02207_, _02208_, _02209_, _02210_, _02211_, _02212_, _02213_, _02214_, _02215_, _02216_, _02217_, _02218_, _02219_, _02220_, _02221_, _02222_, _02223_, _02224_, _02225_, _02226_, _02227_, _02228_, _02229_, _02230_, _02231_, _02232_, _02233_, _02234_, _02235_, _02236_, _02237_, _02238_, _02239_, _02240_, _02241_, _02242_, _02243_, _02244_, _02245_, _02246_, _02247_, _02248_, _02249_, _02250_, _02251_, _02252_, _02253_, _02254_, _02255_, _02256_, _02257_, _02258_, _02259_, _02260_, _02261_, _02262_, _02263_, _02264_, _02265_, _02266_, _02267_, _02268_, _02269_, _02270_, _02271_, _02272_, _02273_, _02274_, _02275_, _02276_, _02277_, _02278_, _02279_, _02280_, _02281_, _02282_, _02283_, _02284_, _02285_, _02286_, _02287_, _02288_, _02289_, _02290_, _02291_, _02292_, _02293_, _02294_, _02295_, _02296_, _02297_, _02298_, _02299_, _02300_, _02301_, _02302_, _02303_, _02304_, _02305_, _02306_, _02307_, _02308_, _02309_, _02310_, _02311_, _02312_, _02313_, _02314_, _02315_, _02316_, _02317_, _02318_, _02319_, _02320_, _02321_, _02322_, _02323_, _02324_, _02325_, _02326_, _02327_, _02328_, _02329_, _02330_, _02331_, _02332_, _02333_, _02334_, _02335_, _02336_, _02337_, _02338_, _02339_, _02340_, _02341_, _02342_, _02343_, _02344_, _02345_, _02346_, _02347_, _02348_, _02349_, _02350_, _02351_, _02352_, _02353_, _02354_, _02355_, _02356_, _02357_, _02358_, _02359_, _02360_, _02361_, _02362_, _02363_, _02364_, _02365_, _02366_, _02367_, _02368_, _02369_, _02370_, _02371_, _02372_, _02373_, _02374_, _02375_, _02376_, _02377_, _02378_, _02379_, _02380_, _02381_, _02382_, _02383_, _02384_, _02385_, _02386_, _02387_, _02388_, _02389_, _02390_, _02391_, _02392_, _02393_, _02394_, _02395_, _02396_, _02397_, _02398_, _02399_, _02400_, _02401_, _02402_, _02403_, _02404_, _02405_, _02406_, _02407_, _02408_, _02409_, _02410_, _02411_, _02412_, _02413_, _02414_, _02415_, _02416_, _02417_, _02418_, _02419_, _02420_, _02421_, _02422_, _02423_, _02424_, _02425_, _02426_, _02427_, _02428_, _02429_, _02430_, _02431_, _02432_, _02433_, _02434_, _02435_, _02436_, _02437_, _02438_, _02439_, _02440_, _02441_, _02442_, _02443_, _02444_, _02445_, _02446_, _02447_, _02448_, _02449_, _02450_, _02451_, _02452_, _02453_, _02454_, _02455_, _02456_, _02457_, _02458_, _02459_, _02460_, _02461_, _02462_, _02463_, _02464_, _02465_, _02466_, _02467_, _02468_, _02469_, _02470_, _02471_, _02472_, _02473_, _02474_, _02475_, _02476_, _02477_, _02478_, _02479_, _02480_, _02481_, _02482_, _02483_, _02484_, _02485_, _02486_, _02487_, _02488_, _02489_, _02490_, _02491_, _02492_, _02493_, _02494_, _02495_, _02496_, _02497_, _02498_, _02499_, _02500_, _02501_, _02502_, _02503_, _02504_, _02505_, _02506_, _02507_, _02508_, _02509_, _02510_, _02511_, _02512_, _02513_, _02514_, _02515_, _02516_, _02517_, _02518_, _02519_, _02520_, _02521_, _02522_, _02523_, _02524_, _02525_, _02526_, _02527_, _02528_, _02529_, _02530_, _02531_, _02532_, _02533_, _02534_, _02535_, _02536_, _02537_, _02538_, _02539_, _02540_, _02541_, _02542_, _02543_, _02544_, _02545_, _02546_, _02547_, _02548_, _02549_, _02550_, _02551_, _02552_, _02553_, _02554_, _02555_, _02556_, _02557_, _02558_, _02559_, _02560_, _02561_, _02562_, _02563_, _02564_, _02565_, _02566_, _02567_, _02568_, _02569_, _02570_, _02571_, _02572_, _02573_, _02574_, _02575_, _02576_, _02577_, _02578_, _02579_, _02580_, _02581_, _02582_, _02583_, _02584_, _02585_, _02586_, _02587_, _02588_, _02589_, _02590_, _02591_, _02592_, _02593_, _02594_, _02595_, _02596_, _02597_, _02598_, _02599_, _02600_, _02601_, _02602_, _02603_, _02604_, _02605_, _02606_, _02607_, _02608_, _02609_, _02610_, _02611_, _02612_, _02613_, _02614_, _02615_, _02616_, _02617_, _02618_, _02619_, _02620_, _02621_, _02622_, _02623_, _02624_, _02625_, _02626_, _02627_, _02628_, _02629_, _02630_, _02631_, _02632_, _02633_, _02634_, _02635_, _02636_, _02637_, _02638_, _02639_, _02640_, _02641_, _02642_, _02643_, _02644_, _02645_, _02646_, _02647_, _02648_, _02649_, _02650_, _02651_, _02652_, _02653_, _02654_, _02655_, _02656_, _02657_, _02658_, _02659_, _02660_, _02661_, _02662_, _02663_, _02664_, _02665_, _02666_, _02667_, _02668_, _02669_, _02670_, _02671_, _02672_, _02673_, _02674_, _02675_, _02676_, _02677_, _02678_, _02679_, _02680_, _02681_, _02682_, _02683_, _02684_, _02685_, _02686_, _02687_, _02688_, _02689_, _02690_, _02691_, _02692_, _02693_, _02694_, _02695_, _02696_, _02697_, _02698_, _02699_, _02700_, _02701_, _02702_, _02703_, _02704_, _02705_, _02706_, _02707_, _02708_, _02709_, _02710_, _02711_, _02712_, _02713_, _02714_, _02715_, _02716_, _02717_, _02718_, _02719_, _02720_, _02721_, _02722_, _02723_, _02724_, _02725_, _02726_, _02727_, _02728_, _02729_, _02730_, _02731_, _02732_, _02733_, _02734_, _02735_, _02736_, _02737_, _02738_, _02739_, _02740_, _02741_, _02742_, _02743_, _02744_, _02745_, _02746_, _02747_, _02748_, _02749_, _02750_, _02751_, _02752_, _02753_, _02754_, _02755_, _02756_, _02757_, _02758_, _02759_, _02760_, _02761_, _02762_, _02763_, _02764_, _02765_, _02766_, _02767_, _02768_, _02769_, _02770_, _02771_, _02772_, _02773_, _02774_, _02775_, _02776_, _02777_, _02778_, _02779_, _02780_, _02781_, _02782_, _02783_, _02784_, _02785_, _02786_, _02787_, _02788_, _02789_, _02790_, _02791_, _02792_, _02793_, _02794_, _02795_, _02796_, _02797_, _02798_, _02799_, _02800_, _02801_, _02802_, _02803_, _02804_, _02805_, _02806_, _02807_, _02808_, _02809_, _02810_, _02811_, _02812_, _02813_, _02814_, _02815_, _02816_, _02817_, _02818_, _02819_, _02820_, _02821_, _02822_, _02823_, _02824_, _02825_, _02826_, _02827_, _02828_, _02829_, _02830_, _02831_, _02832_, _02833_, _02834_, _02835_, _02836_, _02837_, _02838_, _02839_, _02840_, _02841_, _02842_, _02843_, _02844_, _02845_, _02846_, _02847_, _02848_, _02849_, _02850_, _02851_, _02852_, _02853_, _02854_, _02855_, _02856_, _02857_, _02858_, _02859_, _02860_, _02861_, _02862_, _02863_, _02864_, _02865_, _02866_, _02867_, _02868_, _02869_, _02870_, _02871_, _02872_, _02873_, _02874_, _02875_, _02876_, _02877_, _02878_, _02879_, _02880_, _02881_, _02882_, _02883_, _02884_, _02885_, _02886_, _02887_, _02888_, _02889_, _02890_, _02891_, _02892_, _02893_, _02894_, _02895_, _02896_, _02897_, _02898_, _02899_, _02900_, _02901_, _02902_, _02903_, _02904_, _02905_, _02906_, _02907_, _02908_, _02909_, _02910_, _02911_, _02912_, _02913_, _02914_, _02915_, _02916_, _02917_, _02918_, _02919_, _02920_, _02921_, _02922_, _02923_, _02924_, _02925_, _02926_, _02927_, _02928_, _02929_, _02930_, _02931_, _02932_, _02933_, _02934_, _02935_, _02936_, _02937_, _02938_, _02939_, _02940_, _02941_, _02942_, _02943_, _02944_, _02945_, _02946_, _02947_, _02948_, _02949_, _02950_, _02951_, _02952_, _02953_, _02954_, _02955_, _02956_, _02957_, _02958_, _02959_, _02960_, _02961_, _02962_, _02963_, _02964_, _02965_, _02966_, _02967_, _02968_, _02969_, _02970_, _02971_, _02972_, _02973_, _02974_, _02975_, _02976_, _02977_, _02978_, _02979_, _02980_, _02981_, _02982_, _02983_, _02984_, _02985_, _02986_, _02987_, _02988_, _02989_, _02990_, _02991_, _02992_, _02993_, _02994_, _02995_, _02996_, _02997_, _02998_, _02999_, _03000_, _03001_, _03002_, _03003_, _03004_, _03005_, _03006_, _03007_, _03008_, _03009_, _03010_, _03011_, _03012_, _03013_, _03014_, _03015_, _03016_, _03017_, _03018_, _03019_, _03020_, _03021_, _03022_, _03023_, _03024_, _03025_, _03026_, _03027_, _03028_, _03029_, _03030_, _03031_, _03032_, _03033_, _03034_, _03035_, _03036_, _03037_, _03038_, _03039_, _03040_, _03041_, _03042_, _03043_, _03044_, _03045_, _03046_, _03047_, _03048_, _03049_, _03050_, _03051_, _03052_, _03053_, _03054_, _03055_, _03056_, _03057_, _03058_, _03059_, _03060_, _03061_, _03062_, _03063_, _03064_, _03065_, _03066_, _03067_, _03068_, _03069_, _03070_, _03071_, _03072_, _03073_, _03074_, _03075_, _03076_, _03077_, _03078_, _03079_, _03080_, _03081_, _03082_, _03083_, _03084_, _03085_, _03086_, _03087_, _03088_, _03089_, _03090_, _03091_, _03092_, _03093_, _03094_, _03095_, _03096_, _03097_, _03098_, _03099_, _03100_, _03101_, _03102_, _03103_, _03104_, _03105_, _03106_, _03107_, _03108_, _03109_, _03110_, _03111_, _03112_, _03113_, _03114_, _03115_, _03116_, _03117_, _03118_, _03119_, _03120_, _03121_, _03122_, _03123_, _03124_, _03125_, _03126_, _03127_, _03128_, _03129_, _03130_, _03131_, _03132_, _03133_, _03134_, _03135_, _03136_, _03137_, _03138_, _03139_, _03140_, _03141_, _03142_, _03143_, _03144_, _03145_, _03146_, _03147_, _03148_, _03149_, _03150_, _03151_, _03152_, _03153_, _03154_, _03155_, _03156_, _03157_, _03158_, _03159_, _03160_, _03161_, _03162_, _03163_, _03164_, _03165_, _03166_, _03167_, _03168_, _03169_, _03170_, _03171_, _03172_, _03173_, _03174_, _03175_, _03176_, _03177_, _03178_, _03179_, _03180_, _03181_, _03182_, _03183_, _03184_, _03185_, _03186_, _03187_, _03188_, _03189_, _03190_, _03191_, _03192_, _03193_, _03194_, _03195_, _03196_, _03197_, _03198_, _03199_, _03200_, _03201_, _03202_, _03203_, _03204_, _03205_, _03206_, _03207_, _03208_, _03209_, _03210_, _03211_, _03212_, _03213_, _03214_, _03215_, _03216_, _03217_, _03218_, _03219_, _03220_, _03221_, _03222_, _03223_, _03224_, _03225_, _03226_, _03227_, _03228_, _03229_, _03230_, _03231_, _03232_, _03233_, _03234_, _03235_, _03236_, _03237_, _03238_, _03239_, _03240_, _03241_, _03242_, _03243_, _03244_, _03245_, _03246_, _03247_, _03248_, _03249_, _03250_, _03251_, _03252_, _03253_, _03254_, _03255_, _03256_, _03257_, _03258_, _03259_, _03260_, _03261_, _03262_, _03263_, _03264_, _03265_, _03266_, _03267_, _03268_, _03269_, _03270_, _03271_, _03272_, _03273_, _03274_, _03275_, _03276_, _03277_, _03278_, _03279_, _03280_, _03281_, _03282_, _03283_, _03284_, _03285_, _03286_, _03287_, _03288_, _03289_, _03290_, _03291_, _03292_, _03293_, _03294_, _03295_, _03296_, _03297_, _03298_, _03299_, _03300_, _03301_, _03302_, _03303_, _03304_, _03305_, _03306_, _03307_, _03308_, _03309_, _03310_, _03311_, _03312_, _03313_, _03314_, _03315_, _03316_, _03317_, _03318_, _03319_, _03320_, _03321_, _03322_, _03323_, _03324_, _03325_, _03326_, _03327_, _03328_, _03329_, _03330_, _03331_, _03332_, _03333_, _03334_, _03335_, _03336_, _03337_, _03338_, _03339_, _03340_, _03341_, _03342_, _03343_, _03344_, _03345_, _03346_, _03347_, _03348_, _03349_, _03350_, _03351_, _03352_, _03353_, _03354_, _03355_, _03356_, _03357_, _03358_, _03359_, _03360_, _03361_, _03362_, _03363_, _03364_, _03365_, _03366_, _03367_, _03368_, _03369_, _03370_, _03371_, _03372_, _03373_, _03374_, _03375_, _03376_, _03377_, _03378_, _03379_, _03380_, _03381_, _03382_, _03383_, _03384_, _03385_, _03386_, _03387_, _03388_, _03389_, _03390_, _03391_, _03392_, _03393_, _03394_, _03395_, _03396_, _03397_, _03398_, _03399_, _03400_, _03401_, _03402_, _03403_, _03404_, _03405_, _03406_, _03407_, _03408_, _03409_, _03410_, _03411_, _03412_, _03413_, _03414_, _03415_, _03416_, _03417_, _03418_, _03419_, _03420_, _03421_, _03422_, _03423_, _03424_, _03425_, _03426_, _03427_, _03428_, _03429_, _03430_, _03431_, _03432_, _03433_, _03434_, _03435_, _03436_, _03437_, _03438_, _03439_, _03440_, _03441_, _03442_, _03443_, _03444_, _03445_, _03446_, _03447_, _03448_, _03449_, _03450_, _03451_, _03452_, _03453_, _03454_, _03455_, _03456_, _03457_, _03458_, _03459_, _03460_, _03461_, _03462_, _03463_, _03464_, _03465_, _03466_, _03467_, _03468_, _03469_, _03470_, _03471_, _03472_, _03473_, _03474_, _03475_, _03476_, _03477_, _03478_, _03479_, _03480_, _03481_, _03482_, _03483_, _03484_, _03485_, _03486_, _03487_, _03488_, _03489_, _03490_, _03491_, _03492_, _03493_, _03494_, _03495_, _03496_, _03497_, _03498_, _03499_, _03500_, _03501_, _03502_, _03503_, _03504_, _03505_, _03506_, _03507_, _03508_, _03509_, _03510_, _03511_, _03512_, _03513_, _03514_, _03515_, _03516_, _03517_, _03518_, _03519_, _03520_, _03521_, _03522_, _03523_, _03524_, _03525_, _03526_, _03527_, _03528_, _03529_, _03530_, _03531_, _03532_, _03533_, _03534_, _03535_, _03536_, _03537_, _03538_, _03539_, _03540_, _03541_, _03542_, _03543_, _03544_, _03545_, _03546_, _03547_, _03548_, _03549_, _03550_, _03551_, _03552_, _03553_, _03554_, _03555_, _03556_, _03557_, _03558_, _03559_, _03560_, _03561_, _03562_, _03563_, _03564_, _03565_, _03566_, _03567_, _03568_, _03569_, _03570_, _03571_, _03572_, _03573_, _03574_, _03575_, _03576_, _03577_, _03578_, _03579_, _03580_, _03581_, _03582_, _03583_, _03584_, _03585_, _03586_, _03587_, _03588_, _03589_, _03590_, _03591_, _03592_, _03593_, _03594_, _03595_, _03596_, _03597_, _03598_, _03599_, _03600_, _03601_, _03602_, _03603_, _03604_, _03605_, _03606_, _03607_, _03608_, _03609_, _03610_, _03611_, _03612_, _03613_, _03614_, _03615_, _03616_, _03617_, _03618_, _03619_, _03620_, _03621_, _03622_, _03623_, _03624_, _03625_, _03626_, _03627_, _03628_, _03629_, _03630_, _03631_, _03632_, _03633_, _03634_, _03635_, _03636_, _03637_, _03638_, _03639_, _03640_, _03641_, _03642_, _03643_, _03644_, _03645_, _03646_, _03647_, _03648_, _03649_, _03650_, _03651_, _03652_, _03653_, _03654_, _03655_, _03656_, _03657_, _03658_, _03659_, _03660_, _03661_, _03662_, _03663_, _03664_, _03665_, _03666_, _03667_, _03668_, _03669_, _03670_, _03671_, _03672_, _03673_, _03674_, _03675_, _03676_, _03677_, _03678_, _03679_, _03680_, _03681_, _03682_, _03683_, _03684_, _03685_, _03686_, _03687_, _03688_, _03689_, _03690_, _03691_, _03692_, _03693_, _03694_, _03695_, _03696_, _03697_, _03698_, _03699_, _03700_, _03701_, _03702_, _03703_, _03704_, _03705_, _03706_, _03707_, _03708_, _03709_, _03710_, _03711_, _03712_, _03713_, _03714_, _03715_, _03716_, _03717_, _03718_, _03719_, _03720_, _03721_, _03722_, _03723_, _03724_, _03725_, _03726_, _03727_, _03728_, _03729_, _03730_, _03731_, _03732_, _03733_, _03734_, _03735_, _03736_, _03737_, _03738_, _03739_, _03740_, _03741_, _03742_, _03743_, _03744_, _03745_, _03746_, _03747_, _03748_, _03749_, _03750_, _03751_, _03752_, _03753_, _03754_, _03755_, _03756_, _03757_, _03758_, _03759_, _03760_, _03761_, _03762_, _03763_, _03764_, _03765_, _03766_, _03767_, _03768_, _03769_, _03770_, _03771_, _03772_, _03773_, _03774_, _03775_, _03776_, _03777_, _03778_, _03779_, _03780_, _03781_, _03782_, _03783_, _03784_, _03785_, _03786_, _03787_, _03788_, _03789_, _03790_, _03791_, _03792_, _03793_, _03794_, _03795_, _03796_, _03797_, _03798_, _03799_, _03800_, _03801_, _03802_, _03803_, _03804_, _03805_, _03806_, _03807_, _03808_, _03809_, _03810_, _03811_, _03812_, _03813_, _03814_, _03815_, _03816_, _03817_, _03818_, _03819_, _03820_, _03821_, _03822_, _03823_, _03824_, _03825_, _03826_, _03827_, _03828_, _03829_, _03830_, _03831_, _03832_, _03833_, _03834_, _03835_, _03836_, _03837_, _03838_, _03839_, _03840_, _03841_, _03842_, _03843_, _03844_, _03845_, _03846_, _03847_, _03848_, _03849_, _03850_, _03851_, _03852_, _03853_, _03854_, _03855_, _03856_, _03857_, _03858_, _03859_, _03860_, _03861_, _03862_, _03863_, _03864_, _03865_, _03866_, _03867_, _03868_, _03869_, _03870_, _03871_, _03872_, _03873_, _03874_, _03875_, _03876_, _03877_, _03878_, _03879_, _03880_, _03881_, _03882_, _03883_, _03884_, _03885_, _03886_, _03887_, _03888_, _03889_, _03890_, _03891_, _03892_, _03893_, _03894_, _03895_, _03896_, _03897_, _03898_, _03899_, _03900_, _03901_, _03902_, _03903_, _03904_, _03905_, _03906_, _03907_, _03908_, _03909_, _03910_, _03911_, _03912_, _03913_, _03914_, _03915_, _03916_, _03917_, _03918_, _03919_, _03920_, _03921_, _03922_, _03923_, _03924_, _03925_, _03926_, _03927_, _03928_, _03929_, _03930_, _03931_, _03932_, _03933_, _03934_, _03935_, _03936_, _03937_, _03938_, _03939_, _03940_, _03941_, _03942_, _03943_, _03944_, _03945_, _03946_, _03947_, _03948_, _03949_, _03950_, _03951_, _03952_, _03953_, _03954_, _03955_, _03956_, _03957_, _03958_, _03959_, _03960_, _03961_, _03962_, _03963_, _03964_, _03965_, _03966_, _03967_, _03968_, _03969_, _03970_, _03971_, _03972_, _03973_, _03974_, _03975_, _03976_, _03977_, _03978_, _03979_, _03980_, _03981_, _03982_, _03983_, _03984_, _03985_, _03986_, _03987_, _03988_, _03989_, _03990_, _03991_, _03992_, _03993_, _03994_, _03995_, _03996_, _03997_, _03998_, _03999_, _04000_, _04001_, _04002_, _04003_, _04004_, _04005_, _04006_, _04007_, _04008_, _04009_, _04010_, _04011_, _04012_, _04013_, _04014_, _04015_, _04016_, _04017_, _04018_, _04019_, _04020_, _04021_, _04022_, _04023_, _04024_, _04025_, _04026_, _04027_, _04028_, _04029_, _04030_, _04031_, _04032_, _04033_, _04034_, _04035_, _04036_, _04037_, _04038_, _04039_, _04040_, _04041_, _04042_, _04043_, _04044_, _04045_, _04046_, _04047_, _04048_, _04049_, _04050_, _04051_, _04052_, _04053_, _04054_, _04055_, _04056_, _04057_, _04058_, _04059_, _04060_, _04061_, _04062_, _04063_, _04064_, _04065_, _04066_, _04067_, _04068_, _04069_, _04070_, _04071_, _04072_, _04073_, _04074_, _04075_, _04076_, _04077_, _04078_, _04079_, _04080_, _04081_, _04082_, _04083_, _04084_, _04085_, _04086_, _04087_, _04088_, _04089_, _04090_, _04091_, _04092_, _04093_, _04094_, _04095_, _04096_, _04097_, _04098_, _04099_, _04100_, _04101_, _04102_, _04103_, _04104_, _04105_, _04106_, _04107_, _04108_, _04109_, _04110_, _04111_, _04112_, _04113_, _04114_, _04115_, _04116_, _04117_, _04118_, _04119_, _04120_, _04121_, _04122_, _04123_, _04124_, _04125_, _04126_, _04127_, _04128_, _04129_, _04130_, _04131_, _04132_, _04133_, _04134_, _04135_, _04136_, _04137_, _04138_, _04139_, _04140_, _04141_, _04142_, _04143_, _04144_, _04145_, _04146_, _04147_, _04148_, _04149_, _04150_, _04151_, _04152_, _04153_, _04154_, _04155_, _04156_, _04157_, _04158_, _04159_, _04160_, _04161_, _04162_, _04163_, _04164_, _04165_, _04166_, _04167_, _04168_, _04169_, _04170_, _04171_, _04172_, _04173_, _04174_, _04175_, _04176_, _04177_, _04178_, _04179_, _04180_, _04181_, _04182_, _04183_, _04184_, _04185_, _04186_, _04187_, _04188_, _04189_, _04190_, _04191_, _04192_, _04193_, _04194_, _04195_, _04196_, _04197_, _04198_, _04199_, _04200_, _04201_, _04202_, _04203_, _04204_, _04205_, _04206_, _04207_, _04208_, _04209_, _04210_, _04211_, _04212_, _04213_, _04214_, _04215_, _04216_, _04217_, _04218_, _04219_, _04220_, _04221_, _04222_, _04223_, _04224_, _04225_, _04226_, _04227_, _04228_, _04229_, _04230_, _04231_, _04232_, _04233_, _04234_, _04235_, _04236_, _04237_, _04238_, _04239_, _04240_, _04241_, _04242_, _04243_, _04244_, _04245_, _04246_, _04247_, _04248_, _04249_, _04250_, _04251_, _04252_, _04253_, _04254_, _04255_, _04256_, _04257_, _04258_, _04259_, _04260_, _04261_, _04262_, _04263_, _04264_, _04265_, _04266_, _04267_, _04268_, _04269_, _04270_, _04271_, _04272_, _04273_, _04274_, _04275_, _04276_, _04277_, _04278_, _04279_, _04280_, _04281_, _04282_, _04283_, _04284_, _04285_, _04286_, _04287_, _04288_, _04289_, _04290_, _04291_, _04292_, _04293_, _04294_, _04295_, _04296_, _04297_, _04298_, _04299_, _04300_, _04301_, _04302_, _04303_, _04304_, _04305_, _04306_, _04307_, _04308_, _04309_, _04310_, _04311_, _04312_, _04313_, _04314_, _04315_, _04316_, _04317_, _04318_, _04319_, _04320_, _04321_, _04322_, _04323_, _04324_, _04325_, _04326_, _04327_, _04328_, _04329_, _04330_, _04331_, _04332_, _04333_, _04334_, _04335_, _04336_, _04337_, _04338_, _04339_, _04340_, _04341_, _04342_, _04343_, _04344_, _04345_, _04346_, _04347_, _04348_, _04349_, _04350_, _04351_, _04352_, _04353_, _04354_, _04355_, _04356_, _04357_, _04358_, _04359_, _04360_, _04361_, _04362_, _04363_, _04364_, _04365_, _04366_, _04367_, _04368_, _04369_, _04370_, _04371_, _04372_, _04373_, _04374_, _04375_, _04376_, _04377_, _04378_, _04379_, _04380_, _04381_, _04382_, _04383_, _04384_, _04385_, _04386_, _04387_, _04388_, _04389_, _04390_, _04391_, _04392_, _04393_, _04394_, _04395_, _04396_, _04397_, _04398_, _04399_, _04400_, _04401_, _04402_, _04403_, _04404_, _04405_, _04406_, _04407_, _04408_, _04409_, _04410_, _04411_, _04412_, _04413_, _04414_, _04415_, _04416_, _04417_, _04418_, _04419_, _04420_, _04421_, _04422_, _04423_, _04424_, _04425_, _04426_, _04427_, _04428_, _04429_, _04430_, _04431_, _04432_, _04433_, _04434_, _04435_, _04436_, _04437_, _04438_, _04439_, _04440_, _04441_, _04442_, _04443_, _04444_, _04445_, _04446_, _04447_, _04448_, _04449_, _04450_, _04451_, _04452_, _04453_, _04454_, _04455_, _04456_, _04457_, _04458_, _04459_, _04460_, _04461_, _04462_, _04463_, _04464_, _04465_, _04466_, _04467_, _04468_, _04469_, _04470_, _04471_, _04472_, _04473_, _04474_, _04475_, _04476_, _04477_, _04478_, _04479_, _04480_, _04481_, _04482_, _04483_, _04484_, _04485_, _04486_, _04487_, _04488_, _04489_, _04490_, _04491_, _04492_, _04493_, _04494_, _04495_, _04496_, _04497_, _04498_, _04499_, _04500_, _04501_, _04502_, _04503_, _04504_, _04505_, _04506_, _04507_, _04508_, _04509_, _04510_, _04511_, _04512_, _04513_, _04514_, _04515_, _04516_, _04517_, _04518_, _04519_, _04520_, _04521_, _04522_, _04523_, _04524_, _04525_, _04526_, _04527_, _04528_, _04529_, _04530_, _04531_, _04532_, _04533_, _04534_, _04535_, _04536_, _04537_, _04538_, _04539_, _04540_, _04541_, _04542_, _04543_, _04544_, _04545_, _04546_, _04547_, _04548_, _04549_, _04550_, _04551_, _04552_, _04553_, _04554_, _04555_, _04556_, _04557_, _04558_, _04559_, _04560_, _04561_, _04562_, _04563_, _04564_, _04565_, _04566_, _04567_, _04568_, _04569_, _04570_, _04571_, _04572_, _04573_, _04574_, _04575_, _04576_, _04577_, _04578_, _04579_, _04580_, _04581_, _04582_, _04583_, _04584_, _04585_, _04586_, _04587_, _04588_, _04589_, _04590_, _04591_, _04592_, _04593_, _04594_, _04595_, _04596_, _04597_, _04598_, _04599_, _04600_, _04601_, _04602_, _04603_, _04604_, _04605_, _04606_, _04607_, _04608_, _04609_, _04610_, _04611_, _04612_, _04613_, _04614_, _04615_, _04616_, _04617_, _04618_, _04619_, _04620_, _04621_, _04622_, _04623_, _04624_, _04625_, _04626_, _04627_, _04628_, _04629_, _04630_, _04631_, _04632_, _04633_, _04634_, _04635_, _04636_, _04637_, _04638_, _04639_, _04640_, _04641_, _04642_, _04643_, _04644_, _04645_, _04646_, _04647_, _04648_, _04649_, _04650_, _04651_, _04652_, _04653_, _04654_, _04655_, _04656_, _04657_, _04658_, _04659_, _04660_, _04661_, _04662_, _04663_, _04664_, _04665_, _04666_, _04667_, _04668_, _04669_, _04670_, _04671_, _04672_, _04673_, _04674_, _04675_, _04676_, _04677_, _04678_, _04679_, _04680_, _04681_, _04682_, _04683_, _04684_, _04685_, _04686_, _04687_, _04688_, _04689_, _04690_, _04691_, _04692_, _04693_, _04694_, _04695_, _04696_, _04697_, _04698_, _04699_, _04700_, _04701_, _04702_, _04703_, _04704_, _04705_, _04706_, _04707_, _04708_, _04709_, _04710_, _04711_, _04712_, _04713_, _04714_, _04715_, _04716_, _04717_, _04718_, _04719_, _04720_, _04721_, _04722_, _04723_, _04724_, _04725_, _04726_, _04727_, _04728_, _04729_, _04730_, _04731_, _04732_, _04733_, _04734_, _04735_, _04736_, _04737_, _04738_, _04739_, _04740_, _04741_, _04742_, _04743_, _04744_, _04745_, _04746_, _04747_, _04748_, _04749_, _04750_, _04751_, _04752_, _04753_, _04754_, _04755_, _04756_, _04757_, _04758_, _04759_, _04760_, _04761_, _04762_, _04763_, _04764_, _04765_, _04766_, _04767_, _04768_, _04769_, _04770_, _04771_, _04772_, _04773_, _04774_, _04775_, _04776_, _04777_, _04778_, _04779_, _04780_, _04781_, _04782_, _04783_, _04784_, _04785_, _04786_, _04787_, _04788_, _04789_, _04790_, _04791_, _04792_, _04793_, _04794_, _04795_, _04796_, _04797_, _04798_, _04799_, _04800_, _04801_, _04802_, _04803_, _04804_, _04805_, _04806_, _04807_, _04808_, _04809_, _04810_, _04811_, _04812_, _04813_, _04814_, _04815_, _04816_, _04817_, _04818_, _04819_, _04820_, _04821_, _04822_, _04823_, _04824_, _04825_, _04826_, _04827_, _04828_, _04829_, _04830_, _04831_, _04832_, _04833_, _04834_, _04835_, _04836_, _04837_, _04838_, _04839_, _04840_, _04841_, _04842_, _04843_, _04844_, _04845_, _04846_, _04847_, _04848_, _04849_, _04850_, _04851_, _04852_, _04853_, _04854_, _04855_, _04856_, _04857_, _04858_, _04859_, _04860_, _04861_, _04862_, _04863_, _04864_, _04865_, _04866_, _04867_, _04868_, _04869_, _04870_, _04871_, _04872_, _04873_, _04874_, _04875_, _04876_, _04877_, _04878_, _04879_, _04880_, _04881_, _04882_, _04883_, _04884_, _04885_, _04886_, _04887_, _04888_, _04889_, _04890_, _04891_, _04892_, _04893_, _04894_, _04895_, _04896_, _04897_, _04898_, _04899_, _04900_, _04901_, _04902_, _04903_, _04904_, _04905_, _04906_, _04907_, _04908_, _04909_, _04910_, _04911_, _04912_, _04913_, _04914_, _04915_, _04916_, _04917_, _04918_, _04919_, _04920_, _04921_, _04922_, _04923_, _04924_, _04925_, _04926_, _04927_, _04928_, _04929_, _04930_, _04931_, _04932_, _04933_, _04934_, _04935_, _04936_, _04937_, _04938_, _04939_, _04940_, _04941_, _04942_, _04943_, _04944_, _04945_, _04946_, _04947_, _04948_, _04949_, _04950_, _04951_, _04952_, _04953_, _04954_, _04955_, _04956_, _04957_, _04958_, _04959_, _04960_, _04961_, _04962_, _04963_, _04964_, _04965_, _04966_, _04967_, _04968_, _04969_, _04970_, _04971_, _04972_, _04973_, _04974_, _04975_, _04976_, _04977_, _04978_, _04979_, _04980_, _04981_, _04982_, _04983_, _04984_, _04985_, _04986_, _04987_, _04988_, _04989_, _04990_, _04991_, _04992_, _04993_, _04994_, _04995_, _04996_, _04997_, _04998_, _04999_, _05000_, _05001_, _05002_, _05003_, _05004_, _05005_, _05006_, _05007_, _05008_, _05009_, _05010_, _05011_, _05012_, _05013_, _05014_, _05015_, _05016_, _05017_, _05018_, _05019_, _05020_, _05021_, _05022_, _05023_, _05024_, _05025_, _05026_, _05027_, _05028_, _05029_, _05030_, _05031_, _05032_, _05033_, _05034_, _05035_, _05036_, _05037_, _05038_, _05039_, _05040_, _05041_, _05042_, _05043_, _05044_, _05045_, _05046_, _05047_, _05048_, _05049_, _05050_, _05051_, _05052_, _05053_, _05054_, _05055_, _05056_, _05057_, _05058_, _05059_, _05060_, _05061_, _05062_, _05063_, _05064_, _05065_, _05066_, _05067_, _05068_, _05069_, _05070_, _05071_, _05072_, _05073_, _05074_, _05075_, _05076_, _05077_, _05078_, _05079_, _05080_, _05081_, _05082_, _05083_, _05084_, _05085_, _05086_, _05087_, _05088_, _05089_, _05090_, _05091_, _05092_, _05093_, _05094_, _05095_, _05096_, _05097_, _05098_, _05099_, _05100_, _05101_, _05102_, _05103_, _05104_, _05105_, _05106_, _05107_, _05108_, _05109_, _05110_, _05111_, _05112_, _05113_, _05114_, _05115_, _05116_, _05117_, _05118_, _05119_, _05120_, _05121_, _05122_, _05123_, _05124_, _05125_, _05126_, _05127_, _05128_, _05129_, _05130_, _05131_, _05132_, _05133_, _05134_, _05135_, _05136_, _05137_, _05138_, _05139_, _05140_, _05141_, _05142_, _05143_, _05144_, _05145_, _05146_, _05147_, _05148_, _05149_, _05150_, _05151_, _05152_, _05153_, _05154_, _05155_, _05156_, _05157_, _05158_, _05159_, _05160_, _05161_, _05162_, _05163_, _05164_, _05165_, _05166_, _05167_, _05168_, _05169_, _05170_, _05171_, _05172_, _05173_, _05174_, _05175_, _05176_, _05177_, _05178_, _05179_, _05180_, _05181_, _05182_, _05183_, _05184_, _05185_, _05186_, _05187_, _05188_, _05189_, _05190_, _05191_, _05192_, _05193_, _05194_, _05195_, _05196_, _05197_, _05198_, _05199_, _05200_, _05201_, _05202_, _05203_, _05204_, _05205_, _05206_, _05207_, _05208_, _05209_, _05210_, _05211_, _05212_, _05213_, _05214_, _05215_, _05216_, _05217_, _05218_, _05219_, _05220_, _05221_, _05222_, _05223_, _05224_, _05225_, _05226_, _05227_, _05228_, _05229_, _05230_, _05231_, _05232_, _05233_, _05234_, _05235_, _05236_, _05237_, _05238_, _05239_, _05240_, _05241_, _05242_, _05243_, _05244_, _05245_, _05246_, _05247_, _05248_, _05249_, _05250_, _05251_, _05252_, _05253_, _05254_, _05255_, _05256_, _05257_, _05258_, _05259_, _05260_, _05261_, _05262_, _05263_, _05264_, _05265_, _05266_, _05267_, _05268_, _05269_, _05270_, _05271_, _05272_, _05273_, _05274_, _05275_, _05276_, _05277_, _05278_, _05279_, _05280_, _05281_, _05282_, _05283_, _05284_, _05285_, _05286_, _05287_, _05288_, _05289_, _05290_, _05291_, _05292_, _05293_, _05294_, _05295_, _05296_, _05297_, _05298_, _05299_, _05300_, _05301_, _05302_, _05303_, _05304_, _05305_, _05306_, _05307_, _05308_, _05309_, _05310_, _05311_, _05312_, _05313_, _05314_, _05315_, _05316_, _05317_, _05318_, _05319_, _05320_, _05321_, _05322_, _05323_, _05324_, _05325_, _05326_, _05327_, _05328_, _05329_, _05330_, _05331_, _05332_, _05333_, _05334_, _05335_, _05336_, _05337_, _05338_, _05339_, _05340_, _05341_, _05342_, _05343_, _05344_, _05345_, _05346_, _05347_, _05348_, _05349_, _05350_, _05351_, _05352_, _05353_, _05354_, _05355_, _05356_, _05357_, _05358_, _05359_, _05360_, _05361_, _05362_, _05363_, _05364_, _05365_, _05366_, _05367_, _05368_, _05369_, _05370_, _05371_, _05372_, _05373_, _05374_, _05375_, _05376_, _05377_, _05378_, _05379_, _05380_, _05381_, _05382_, _05383_, _05384_, _05385_, _05386_, _05387_, _05388_, _05389_, _05390_, _05391_, _05392_, _05393_, _05394_, _05395_, _05396_, _05397_, _05398_, _05399_, _05400_, _05401_, _05402_, _05403_, _05404_, _05405_, _05406_, _05407_, _05408_, _05409_, _05410_, _05411_, _05412_, _05413_, _05414_, _05415_, _05416_, _05417_, _05418_, _05419_, _05420_, _05421_, _05422_, _05423_, _05424_, _05425_, _05426_, _05427_, _05428_, _05429_, _05430_, _05431_, _05432_, _05433_, _05434_, _05435_, _05436_, _05437_, _05438_, _05439_, _05440_, _05441_, _05442_, _05443_, _05444_, _05445_, _05446_, _05447_, _05448_, _05449_, _05450_, _05451_, _05452_, _05453_, _05454_, _05455_, _05456_, _05457_, _05458_, _05459_, _05460_, _05461_, _05462_, _05463_, _05464_, _05465_, _05466_, _05467_, _05468_, _05469_, _05470_, _05471_, _05472_, _05473_, _05474_, _05475_, _05476_, _05477_, _05478_, _05479_, _05480_, _05481_, _05482_, _05483_, _05484_, _05485_, _05486_, _05487_, _05488_, _05489_, _05490_, _05491_, _05492_, _05493_, _05494_, _05495_, _05496_, _05497_, _05498_, _05499_, _05500_, _05501_, _05502_, _05503_, _05504_, _05505_, _05506_, _05507_, _05508_, _05509_, _05510_, _05511_, _05512_, _05513_, _05514_, _05515_, _05516_, _05517_, _05518_, _05519_, _05520_, _05521_, _05522_, _05523_, _05524_, _05525_, _05526_, _05527_, _05528_, _05529_, _05530_, _05531_, _05532_, _05533_, _05534_, _05535_, _05536_, _05537_, _05538_, _05539_, _05540_, _05541_, _05542_, _05543_, _05544_, _05545_, _05546_, _05547_, _05548_, _05549_, _05550_, _05551_, _05552_, _05553_, _05554_, _05555_, _05556_, _05557_, _05558_, _05559_, _05560_, _05561_, _05562_, _05563_, _05564_, _05565_, _05566_, _05567_, _05568_, _05569_, _05570_, _05571_, _05572_, _05573_, _05574_, _05575_, _05576_, _05577_, _05578_, _05579_, _05580_, _05581_, _05582_, _05583_, _05584_, _05585_, _05586_, _05587_, _05588_, _05589_, _05590_, _05591_, _05592_, _05593_, _05594_, _05595_, _05596_, _05597_, _05598_, _05599_, _05600_, _05601_, _05602_, _05603_, _05604_, _05605_, _05606_, _05607_, _05608_, _05609_, _05610_, _05611_, _05612_, _05613_, _05614_, _05615_, _05616_, _05617_, _05618_, _05619_, _05620_, _05621_, _05622_, _05623_, _05624_, _05625_, _05626_, _05627_, _05628_, _05629_, _05630_, _05631_, _05632_, _05633_, _05634_, _05635_, _05636_, _05637_, _05638_, _05639_, _05640_, _05641_, _05642_, _05643_, _05644_, _05645_, _05646_, _05647_, _05648_, _05649_, _05650_, _05651_, _05652_, _05653_, _05654_, _05655_, _05656_, _05657_, _05658_, _05659_, _05660_, _05661_, _05662_, _05663_, _05664_, _05665_, _05666_, _05667_, _05668_, _05669_, _05670_, _05671_, _05672_, _05673_, _05674_, _05675_, _05676_, _05677_, _05678_, _05679_, _05680_, _05681_, _05682_, _05683_, _05684_, _05685_, _05686_, _05687_, _05688_, _05689_, _05690_, _05691_, _05692_, _05693_, _05694_, _05695_, _05696_, _05697_, _05698_, _05699_, _05700_, _05701_, _05702_, _05703_, _05704_, _05705_, _05706_, _05707_, _05708_, _05709_, _05710_, _05711_, _05712_, _05713_, _05714_, _05715_, _05716_, _05717_, _05718_, _05719_, _05720_, _05721_, _05722_, _05723_, _05724_, _05725_, _05726_, _05727_, _05728_, _05729_, _05730_, _05731_, _05732_, _05733_, _05734_, _05735_, _05736_, _05737_, _05738_, _05739_, _05740_, _05741_, _05742_, _05743_, _05744_, _05745_, _05746_, _05747_, _05748_, _05749_, _05750_, _05751_, _05752_, _05753_, _05754_, _05755_, _05756_, _05757_, _05758_, _05759_, _05760_, _05761_, _05762_, _05763_, _05764_, _05765_, _05766_, _05767_, _05768_, _05769_, _05770_, _05771_, _05772_, _05773_, _05774_, _05775_, _05776_, _05777_, _05778_, _05779_, _05780_, _05781_, _05782_, _05783_, _05784_, _05785_, _05786_, _05787_, _05788_, _05789_, _05790_, _05791_, _05792_, _05793_, _05794_, _05795_, _05796_, _05797_, _05798_, _05799_, _05800_, _05801_, _05802_, _05803_, _05804_, _05805_, _05806_, _05807_, _05808_, _05809_, _05810_, _05811_, _05812_, _05813_, _05814_, _05815_, _05816_, _05817_, _05818_, _05819_, _05820_, _05821_, _05822_, _05823_, _05824_, _05825_, _05826_, _05827_, _05828_, _05829_, _05830_, _05831_, _05832_, _05833_, _05834_, _05835_, _05836_, _05837_, _05838_, _05839_, _05840_, _05841_, _05842_, _05843_, _05844_, _05845_, _05846_, _05847_, _05848_, _05849_, _05850_, _05851_, _05852_, _05853_, _05854_, _05855_, _05856_, _05857_, _05858_, _05859_, _05860_, _05861_, _05862_, _05863_, _05864_, _05865_, _05866_, _05867_, _05868_, _05869_, _05870_, _05871_, _05872_, _05873_, _05874_, _05875_, _05876_, _05877_, _05878_, _05879_, _05880_, _05881_, _05882_, _05883_, _05884_, _05885_, _05886_, _05887_, _05888_, _05889_, _05890_, _05891_, _05892_, _05893_, _05894_, _05895_, _05896_, _05897_, _05898_, _05899_, _05900_, _05901_, _05902_, _05903_, _05904_, _05905_, _05906_, _05907_, _05908_, _05909_, _05910_, _05911_, _05912_, _05913_, _05914_, _05915_, _05916_, _05917_, _05918_, _05919_, _05920_, _05921_, _05922_, _05923_, _05924_, _05925_, _05926_, _05927_, _05928_, _05929_, _05930_, _05931_, _05932_, _05933_, _05934_, _05935_, _05936_, _05937_, _05938_, _05939_, _05940_, _05941_, _05942_, _05943_, _05944_, _05945_, _05946_, _05947_, _05948_, _05949_, _05950_, _05951_, _05952_, _05953_, _05954_, _05955_, _05956_, _05957_, _05958_, _05959_, _05960_, _05961_, _05962_, _05963_, _05964_, _05965_, _05966_, _05967_, _05968_, _05969_, _05970_, _05971_, _05972_, _05973_, _05974_, _05975_, _05976_, _05977_, _05978_, _05979_, _05980_, _05981_, _05982_, _05983_, _05984_, _05985_, _05986_, _05987_, _05988_, _05989_, _05990_, _05991_, _05992_, _05993_, _05994_, _05995_, _05996_, _05997_, _05998_, _05999_, _06000_, _06001_, _06002_, _06003_, _06004_, _06005_, _06006_, _06007_, _06008_, _06009_, _06010_, _06011_, _06012_, _06013_, _06014_, _06015_, _06016_, _06017_, _06018_, _06019_, _06020_, _06021_, _06022_, _06023_, _06024_, _06025_, _06026_, _06027_, _06028_, _06029_, _06030_, _06031_, _06032_, _06033_, _06034_, _06035_, _06036_, _06037_, _06038_, _06039_, _06040_, _06041_, _06042_, _06043_, _06044_, _06045_, _06046_, _06047_, _06048_, _06049_, _06050_, _06051_, _06052_, _06053_, _06054_, _06055_, _06056_, _06057_, _06058_, _06059_, _06060_, _06061_, _06062_, _06063_, _06064_, _06065_, _06066_, _06067_, _06068_, _06069_, _06070_, _06071_, _06072_, _06073_, _06074_, _06075_, _06076_, _06077_, _06078_, _06079_, _06080_, _06081_, _06082_, _06083_, _06084_, _06085_, _06086_, _06087_, _06088_, _06089_, _06090_, _06091_, _06092_, _06093_, _06094_, _06095_, _06096_, _06097_, _06098_, _06099_, _06100_, _06101_, _06102_, _06103_, _06104_, _06105_, _06106_, _06107_, _06108_, _06109_, _06110_, _06111_, _06112_, _06113_, _06114_, _06115_, _06116_, _06117_, _06118_, _06119_, _06120_, _06121_, _06122_, _06123_, _06124_, _06125_, _06126_, _06127_, _06128_, _06129_, _06130_, _06131_, _06132_, _06133_, _06134_, _06135_, _06136_, _06137_, _06138_, _06139_, _06140_, _06141_, _06142_, _06143_, _06144_, _06145_, _06146_, _06147_, _06148_, _06149_, _06150_, _06151_, _06152_, _06153_, _06154_, _06155_, _06156_, _06157_, _06158_, _06159_, _06160_, _06161_, _06162_, _06163_, _06164_, _06165_, _06166_, _06167_, _06168_, _06169_, _06170_, _06171_, _06172_, _06173_, _06174_, _06175_, _06176_, _06177_, _06178_, _06179_, _06180_, _06181_, _06182_, _06183_, _06184_, _06185_, _06186_, _06187_, _06188_, _06189_, _06190_, _06191_, _06192_, _06193_, _06194_, _06195_, _06196_, _06197_, _06198_, _06199_, _06200_, _06201_, _06202_, _06203_, _06204_, _06205_, _06206_, _06207_, _06208_, _06209_, _06210_, _06211_, _06212_, _06213_, _06214_, _06215_, _06216_, _06217_, _06218_, _06219_, _06220_, _06221_, _06222_, _06223_, _06224_, _06225_, _06226_, _06227_, _06228_, _06229_, _06230_, _06231_, _06232_, _06233_, _06234_, _06235_, _06236_, _06237_, _06238_, _06239_, _06240_, _06241_, _06242_, _06243_, _06244_, _06245_, _06246_, _06247_, _06248_, _06249_, _06250_, _06251_, _06252_, _06253_, _06254_, _06255_, _06256_, _06257_, _06258_, _06259_, _06260_, _06261_, _06262_, _06263_, _06264_, _06265_, _06266_, _06267_, _06268_, _06269_, _06270_, _06271_, _06272_, _06273_, _06274_, _06275_, _06276_, _06277_, _06278_, _06279_, _06280_, _06281_, _06282_, _06283_, _06284_, _06285_, _06286_, _06287_, _06288_, _06289_, _06290_, _06291_, _06292_, _06293_, _06294_, _06295_, _06296_, _06297_, _06298_, _06299_, _06300_, _06301_, _06302_, _06303_, _06304_, _06305_, _06306_, _06307_, _06308_, _06309_, _06310_, _06311_, _06312_, _06313_, _06314_, _06315_, _06316_, _06317_, _06318_, _06319_, _06320_, _06321_, _06322_, _06323_, _06324_, _06325_, _06326_, _06327_, _06328_, _06329_, _06330_, _06331_, _06332_, _06333_, _06334_, _06335_, _06336_, _06337_, _06338_, _06339_, _06340_, _06341_, _06342_, _06343_, _06344_, _06345_, _06346_, _06347_, _06348_, _06349_, _06350_, _06351_, _06352_, _06353_, _06354_, _06355_, _06356_, _06357_, _06358_, _06359_, _06360_, _06361_, _06362_, _06363_, _06364_, _06365_, _06366_, _06367_, _06368_, _06369_, _06370_, _06371_, _06372_, _06373_, _06374_, _06375_, _06376_, _06377_, _06378_, _06379_, _06380_, _06381_, _06382_, _06383_, _06384_, _06385_, _06386_, _06387_, _06388_, _06389_, _06390_, _06391_, _06392_, _06393_, _06394_, _06395_, _06396_, _06397_, _06398_, _06399_, _06400_, _06401_, _06402_, _06403_, _06404_, _06405_, _06406_, _06407_, _06408_, _06409_, _06410_, _06411_, _06412_, _06413_, _06414_, _06415_, _06416_, _06417_, _06418_, _06419_, _06420_, _06421_, _06422_, _06423_, _06424_, _06425_, _06426_, _06427_, _06428_, _06429_, _06430_, _06431_, _06432_, _06433_, _06434_, _06435_, _06436_, _06437_, _06438_, _06439_, _06440_, _06441_, _06442_, _06443_, _06444_, _06445_, _06446_, _06447_, _06448_, _06449_, _06450_, _06451_, _06452_, _06453_, _06454_, _06455_, _06456_, _06457_, _06458_, _06459_, _06460_, _06461_, _06462_, _06463_, _06464_, _06465_, _06466_, _06467_, _06468_, _06469_, _06470_, _06471_, _06472_, _06473_, _06474_, _06475_, _06476_, _06477_, _06478_, _06479_, _06480_, _06481_, _06482_, _06483_, _06484_, _06485_, _06486_, _06487_, _06488_, _06489_, _06490_, _06491_, _06492_, _06493_, _06494_, _06495_, _06496_, _06497_, _06498_, _06499_, _06500_, _06501_, _06502_, _06503_, _06504_, _06505_, _06506_, _06507_, _06508_, _06509_, _06510_, _06511_, _06512_, _06513_, _06514_, _06515_, _06516_, _06517_, _06518_, _06519_, _06520_, _06521_, _06522_, _06523_, _06524_, _06525_, _06526_, _06527_, _06528_, _06529_, _06530_, _06531_, _06532_, _06533_, _06534_, _06535_, _06536_, _06537_, _06538_, _06539_, _06540_, _06541_, _06542_, _06543_, _06544_, _06545_, _06546_, _06547_, _06548_, _06549_, _06550_, _06551_, _06552_, _06553_, _06554_, _06555_, _06556_, _06557_, _06558_, _06559_, _06560_, _06561_, _06562_, _06563_, _06564_, _06565_, _06566_, _06567_, _06568_, _06569_, _06570_, _06571_, _06572_, _06573_, _06574_, _06575_, _06576_, _06577_, _06578_, _06579_, _06580_, _06581_, _06582_, _06583_, _06584_, _06585_, _06586_, _06587_, _06588_, _06589_, _06590_, _06591_, _06592_, _06593_, _06594_, _06595_, _06596_, _06597_, _06598_, _06599_, _06600_, _06601_, _06602_, _06603_, _06604_, _06605_, _06606_, _06607_, _06608_, _06609_, _06610_, _06611_, _06612_, _06613_, _06614_, _06615_, _06616_, _06617_, _06618_, _06619_, _06620_, _06621_, _06622_, _06623_, _06624_, _06625_, _06626_, _06627_, _06628_, _06629_, _06630_, _06631_, _06632_, _06633_, _06634_, _06635_, _06636_, _06637_, _06638_, _06639_, _06640_, _06641_, _06642_, _06643_, _06644_, _06645_, _06646_, _06647_, _06648_, _06649_, _06650_, _06651_, _06652_, _06653_, _06654_, _06655_, _06656_, _06657_, _06658_, _06659_, _06660_, _06661_, _06662_, _06663_, _06664_, _06665_, _06666_, _06667_, _06668_, _06669_, _06670_, _06671_, _06672_, _06673_, _06674_, _06675_, _06676_, _06677_, _06678_, _06679_, _06680_, _06681_, _06682_, _06683_, _06684_, _06685_, _06686_, _06687_, _06688_, _06689_, _06690_, _06691_, _06692_, _06693_, _06694_, _06695_, _06696_, _06697_, _06698_, _06699_, _06700_, _06701_, _06702_, _06703_, _06704_, _06705_, _06706_, _06707_, _06708_, _06709_, _06710_, _06711_, _06712_, _06713_, _06714_, _06715_, _06716_, _06717_, _06718_, _06719_, _06720_, _06721_, _06722_, _06723_, _06724_, _06725_, _06726_, _06727_, _06728_, _06729_, _06730_, _06731_, _06732_, _06733_, _06734_, _06735_, _06736_, _06737_, _06738_, _06739_, _06740_, _06741_, _06742_, _06743_, _06744_, _06745_, _06746_, _06747_, _06748_, _06749_, _06750_, _06751_, _06752_, _06753_, _06754_, _06755_, _06756_, _06757_, _06758_, _06759_, _06760_, _06761_, _06762_, _06763_, _06764_, _06765_, _06766_, _06767_, _06768_, _06769_, _06770_, _06771_, _06772_, _06773_, _06774_, _06775_, _06776_, _06777_, _06778_, _06779_, _06780_, _06781_, _06782_, _06783_, _06784_, _06785_, _06786_, _06787_, _06788_, _06789_, _06790_, _06791_, _06792_, _06793_, _06794_, _06795_, _06796_, _06797_, _06798_, _06799_, _06800_, _06801_, _06802_, _06803_, _06804_, _06805_, _06806_, _06807_, _06808_, _06809_, _06810_, _06811_, _06812_, _06813_, _06814_, _06815_, _06816_, _06817_, _06818_, _06819_, _06820_, _06821_, _06822_, _06823_, _06824_, _06825_, _06826_, _06827_, _06828_, _06829_, _06830_, _06831_, _06832_, _06833_, _06834_, _06835_, _06836_, _06837_, _06838_, _06839_, _06840_, _06841_, _06842_, _06843_, _06844_, _06845_, _06846_, _06847_, _06848_, _06849_, _06850_, _06851_, _06852_, _06853_, _06854_, _06855_, _06856_, _06857_, _06858_, _06859_, _06860_, _06861_, _06862_, _06863_, _06864_, _06865_, _06866_, _06867_, _06868_, _06869_, _06870_, _06871_, _06872_, _06873_, _06874_, _06875_, _06876_, _06877_, _06878_, _06879_, _06880_, _06881_, _06882_, _06883_, _06884_, _06885_, _06886_, _06887_, _06888_, _06889_, _06890_, _06891_, _06892_, _06893_, _06894_, _06895_, _06896_, _06897_, _06898_, _06899_, _06900_, _06901_, _06902_, _06903_, _06904_, _06905_, _06906_, _06907_, _06908_, _06909_, _06910_, _06911_, _06912_, _06913_, _06914_, _06915_, _06916_, _06917_, _06918_, _06919_, _06920_, _06921_, _06922_, _06923_, _06924_, _06925_, _06926_, _06927_, _06928_, _06929_, _06930_, _06931_, _06932_, _06933_, _06934_, _06935_, _06936_, _06937_, _06938_, _06939_, _06940_, _06941_, _06942_, _06943_, _06944_, _06945_, _06946_, _06947_, _06948_, _06949_, _06950_, _06951_, _06952_, _06953_, _06954_, _06955_, _06956_, _06957_, _06958_, _06959_, _06960_, _06961_, _06962_, _06963_, _06964_, _06965_, _06966_, _06967_, _06968_, _06969_, _06970_, _06971_, _06972_, _06973_, _06974_, _06975_, _06976_, _06977_, _06978_, _06979_, _06980_, _06981_, _06982_, _06983_, _06984_, _06985_, _06986_, _06987_, _06988_, _06989_, _06990_, _06991_, _06992_, _06993_, _06994_, _06995_, _06996_, _06997_, _06998_, _06999_, _07000_, _07001_, _07002_, _07003_, _07004_, _07005_, _07006_, _07007_, _07008_, _07009_, _07010_, _07011_, _07012_, _07013_, _07014_, _07015_, _07016_, _07017_, _07018_, _07019_, _07020_, _07021_, _07022_, _07023_, _07024_, _07025_, _07026_, _07027_, _07028_, _07029_, _07030_, _07031_, _07032_, _07033_, _07034_, _07035_, _07036_, _07037_, _07038_, _07039_, _07040_, _07041_, _07042_, _07043_, _07044_, _07045_, _07046_, _07047_, _07048_, _07049_, _07050_, _07051_, _07052_, _07053_, _07054_, _07055_, _07056_, _07057_, _07058_, _07059_, _07060_, _07061_, _07062_, _07063_, _07064_, _07065_, _07066_, _07067_, _07068_, _07069_, _07070_, _07071_, _07072_, _07073_, _07074_, _07075_, _07076_, _07077_, _07078_, _07079_, _07080_, _07081_, _07082_, _07083_, _07084_, _07085_, _07086_, _07087_, _07088_, _07089_, _07090_, _07091_, _07092_, _07093_, _07094_, _07095_, _07096_, _07097_, _07098_, _07099_, _07100_, _07101_, _07102_, _07103_, _07104_, _07105_, _07106_, _07107_, _07108_, _07109_, _07110_, _07111_, _07112_, _07113_, _07114_, _07115_, _07116_, _07117_, _07118_, _07119_, _07120_, _07121_, _07122_, _07123_, _07124_, _07125_, _07126_, _07127_, _07128_, _07129_, _07130_, _07131_, _07132_, _07133_, _07134_, _07135_, _07136_, _07137_, _07138_, _07139_, _07140_, _07141_, _07142_, _07143_, _07144_, _07145_, _07146_, _07147_, _07148_, _07149_, _07150_, _07151_, _07152_, _07153_, _07154_, _07155_, _07156_, _07157_, _07158_, _07159_, _07160_, _07161_, _07162_, _07163_, _07164_, _07165_, _07166_, _07167_, _07168_, _07169_, _07170_, _07171_, _07172_, _07173_, _07174_, _07175_, _07176_, _07177_, _07178_, _07179_, _07180_, _07181_, _07182_, _07183_, _07184_, _07185_, _07186_, _07187_, _07188_, _07189_, _07190_, _07191_, _07192_, _07193_, _07194_, _07195_, _07196_, _07197_, _07198_, _07199_, _07200_, _07201_, _07202_, _07203_, _07204_, _07205_, _07206_, _07207_, _07208_, _07209_, _07210_, _07211_, _07212_, _07213_, _07214_, _07215_, _07216_, _07217_, _07218_, _07219_, _07220_, _07221_, _07222_, _07223_, _07224_, _07225_, _07226_, _07227_, _07228_, _07229_, _07230_, _07231_, _07232_, _07233_, _07234_, _07235_, _07236_, _07237_, _07238_, _07239_, _07240_, _07241_, _07242_, _07243_, _07244_, _07245_, _07246_, _07247_, _07248_, _07249_, _07250_, _07251_, _07252_, _07253_, _07254_, _07255_, _07256_, _07257_, _07258_, _07259_, _07260_, _07261_, _07262_, _07263_, _07264_, _07265_, _07266_, _07267_, _07268_, _07269_, _07270_, _07271_, _07272_, _07273_, _07274_, _07275_, _07276_, _07277_, _07278_, _07279_, _07280_, _07281_, _07282_, _07283_, _07284_, _07285_, _07286_, _07287_, _07288_, _07289_, _07290_, _07291_, _07292_, _07293_, _07294_, _07295_, _07296_, _07297_, _07298_, _07299_, _07300_, _07301_, _07302_, _07303_, _07304_, _07305_, _07306_, _07307_, _07308_, _07309_, _07310_, _07311_, _07312_, _07313_, _07314_, _07315_, _07316_, _07317_, _07318_, _07319_, _07320_, _07321_, _07322_, _07323_, _07324_, _07325_, _07326_, _07327_, _07328_, _07329_, _07330_, _07331_, _07332_, _07333_, _07334_, _07335_, _07336_, _07337_, _07338_, _07339_, _07340_, _07341_, _07342_, _07343_, _07344_, _07345_, _07346_, _07347_, _07348_, _07349_, _07350_, _07351_, _07352_, _07353_, _07354_, _07355_, _07356_, _07357_, _07358_, _07359_, _07360_, _07361_, _07362_, _07363_, _07364_, _07365_, _07366_, _07367_, _07368_, _07369_, _07370_, _07371_, _07372_, _07373_, _07374_, _07375_, _07376_, _07377_, _07378_, _07379_, _07380_, _07381_, _07382_, _07383_, _07384_, _07385_, _07386_, _07387_, _07388_, _07389_, _07390_, _07391_, _07392_, _07393_, _07394_, _07395_, _07396_, _07397_, _07398_, _07399_, _07400_, _07401_, _07402_, _07403_, _07404_, _07405_, _07406_, _07407_, _07408_, _07409_, _07410_, _07411_, _07412_, _07413_, _07414_, _07415_, _07416_, _07417_, _07418_, _07419_, _07420_, _07421_, _07422_, _07423_, _07424_, _07425_, _07426_, _07427_, _07428_, _07429_, _07430_, _07431_, _07432_, _07433_, _07434_, _07435_, _07436_, _07437_, _07438_, _07439_, _07440_, _07441_, _07442_, _07443_, _07444_, _07445_, _07446_, _07447_, _07448_, _07449_, _07450_, _07451_, _07452_, _07453_, _07454_, _07455_, _07456_, _07457_, _07458_, _07459_, _07460_, _07461_, _07462_, _07463_, _07464_, _07465_, _07466_, _07467_, _07468_, _07469_, _07470_, _07471_, _07472_, _07473_, _07474_, _07475_, _07476_, _07477_, _07478_, _07479_, _07480_, _07481_, _07482_, _07483_, _07484_, _07485_, _07486_, _07487_, _07488_, _07489_, _07490_, _07491_, _07492_, _07493_, _07494_, _07495_, _07496_, _07497_, _07498_, _07499_, _07500_, _07501_, _07502_, _07503_, _07504_, _07505_, _07506_, _07507_, _07508_, _07509_, _07510_, _07511_, _07512_, _07513_, _07514_, _07515_, _07516_, _07517_, _07518_, _07519_, _07520_, _07521_, _07522_, _07523_, _07524_, _07525_, _07526_, _07527_, _07528_, _07529_, _07530_, _07531_, _07532_, _07533_, _07534_, _07535_, _07536_, _07537_, _07538_, _07539_, _07540_, _07541_, _07542_, _07543_, _07544_, _07545_, _07546_, _07547_, _07548_, _07549_, _07550_, _07551_, _07552_, _07553_, _07554_, _07555_, _07556_, _07557_, _07558_, _07559_, _07560_, _07561_, _07562_, _07563_, _07564_, _07565_, _07566_, _07567_, _07568_, _07569_, _07570_, _07571_, _07572_, _07573_, _07574_, _07575_, _07576_, _07577_, _07578_, _07579_, _07580_, _07581_, _07582_, _07583_, _07584_, _07585_, _07586_, _07587_, _07588_, _07589_, _07590_, _07591_, _07592_, _07593_, _07594_, _07595_, _07596_, _07597_, _07598_, _07599_, _07600_, _07601_, _07602_, _07603_, _07604_, _07605_, _07606_, _07607_, _07608_, _07609_, _07610_, _07611_, _07612_, _07613_, _07614_, _07615_, _07616_, _07617_, _07618_, _07619_, _07620_, _07621_, _07622_, _07623_, _07624_, _07625_, _07626_, _07627_, _07628_, _07629_, _07630_, _07631_, _07632_, _07633_, _07634_, _07635_, _07636_, _07637_, _07638_, _07639_, _07640_, _07641_, _07642_, _07643_, _07644_, _07645_, _07646_, _07647_, _07648_, _07649_, _07650_, _07651_, _07652_, _07653_, _07654_, _07655_, _07656_, _07657_, _07658_, _07659_, _07660_, _07661_, _07662_, _07663_, _07664_, _07665_, _07666_, _07667_, _07668_, _07669_, _07670_, _07671_, _07672_, _07673_, _07674_, _07675_, _07676_, _07677_, _07678_, _07679_, _07680_, _07681_, _07682_, _07683_, _07684_, _07685_, _07686_, _07687_, _07688_, _07689_, _07690_, _07691_, _07692_, _07693_, _07694_, _07695_, _07696_, _07697_, _07698_, _07699_, _07700_, _07701_, _07702_, _07703_, _07704_, _07705_, _07706_, _07707_, _07708_, _07709_, _07710_, _07711_, _07712_, _07713_, _07714_, _07715_, _07716_, _07717_, _07718_, _07719_, _07720_, _07721_, _07722_, _07723_, _07724_, _07725_, _07726_, _07727_, _07728_, _07729_, _07730_, _07731_, _07732_, _07733_, _07734_, _07735_, _07736_, _07737_, _07738_, _07739_, _07740_, _07741_, _07742_, _07743_, _07744_, _07745_, _07746_, _07747_, _07748_, _07749_, _07750_, _07751_, _07752_, _07753_, _07754_, _07755_, _07756_, _07757_, _07758_, _07759_, _07760_, _07761_, _07762_, _07763_, _07764_, _07765_, _07766_, _07767_, _07768_, _07769_, _07770_, _07771_, _07772_, _07773_, _07774_, _07775_, _07776_, _07777_, _07778_, _07779_, _07780_, _07781_, _07782_, _07783_, _07784_, _07785_, _07786_, _07787_, _07788_, _07789_, _07790_, _07791_, _07792_, _07793_, _07794_, _07795_, _07796_, _07797_, _07798_, _07799_, _07800_, _07801_, _07802_, _07803_, _07804_, _07805_, _07806_, _07807_, _07808_, _07809_, _07810_, _07811_, _07812_, _07813_, _07814_, _07815_, _07816_, _07817_, _07818_, _07819_, _07820_, _07821_, _07822_, _07823_, _07824_, _07825_, _07826_, _07827_, _07828_, _07829_, _07830_, _07831_, _07832_, _07833_, _07834_, _07835_, _07836_, _07837_, _07838_, _07839_, _07840_, _07841_, _07842_, _07843_, _07844_, _07845_, _07846_, _07847_, _07848_, _07849_, _07850_, _07851_, _07852_, _07853_, _07854_, _07855_, _07856_, _07857_, _07858_, _07859_, _07860_, _07861_, _07862_, _07863_, _07864_, _07865_, _07866_, _07867_, _07868_, _07869_, _07870_, _07871_, _07872_, _07873_, _07874_, _07875_, _07876_, _07877_, _07878_, _07879_, _07880_, _07881_, _07882_, _07883_, _07884_, _07885_, _07886_, _07887_, _07888_, _07889_, _07890_, _07891_, _07892_, _07893_, _07894_, _07895_, _07896_, _07897_, _07898_, _07899_, _07900_, _07901_, _07902_, _07903_, _07904_, _07905_, _07906_, _07907_, _07908_, _07909_, _07910_, _07911_, _07912_, _07913_, _07914_, _07915_, _07916_, _07917_, _07918_, _07919_, _07920_, _07921_, _07922_, _07923_, _07924_, _07925_, _07926_, _07927_, _07928_, _07929_, _07930_, _07931_, _07932_, _07933_, _07934_, _07935_, _07936_, _07937_, _07938_, _07939_, _07940_, _07941_, _07942_, _07943_, _07944_, _07945_, _07946_, _07947_, _07948_, _07949_, _07950_, _07951_, _07952_, _07953_, _07954_, _07955_, _07956_, _07957_, _07958_, _07959_, _07960_, _07961_, _07962_, _07963_, _07964_, _07965_, _07966_, _07967_, _07968_, _07969_, _07970_, _07971_, _07972_, _07973_, _07974_, _07975_, _07976_, _07977_, _07978_, _07979_, _07980_, _07981_, _07982_, _07983_, _07984_, _07985_, _07986_, _07987_, _07988_, _07989_, _07990_, _07991_, _07992_, _07993_, _07994_, _07995_, _07996_, _07997_, _07998_, _07999_, _08000_, _08001_, _08002_, _08003_, _08004_, _08005_, _08006_, _08007_, _08008_, _08009_, _08010_, _08011_, _08012_, _08013_, _08014_, _08015_, _08016_, _08017_, _08018_, _08019_, _08020_, _08021_, _08022_, _08023_, _08024_, _08025_, _08026_, _08027_, _08028_, _08029_, _08030_, _08031_, _08032_, _08033_, _08034_, _08035_, _08036_, _08037_, _08038_, _08039_, _08040_, _08041_, _08042_, _08043_, _08044_, _08045_, _08046_, _08047_, _08048_, _08049_, _08050_, _08051_, _08052_, _08053_, _08054_, _08055_, _08056_, _08057_, _08058_, _08059_, _08060_, _08061_, _08062_, _08063_, _08064_, _08065_, _08066_, _08067_, _08068_, _08069_, _08070_, _08071_, _08072_, _08073_, _08074_, _08075_, _08076_, _08077_, _08078_, _08079_, _08080_, _08081_, _08082_, _08083_, _08084_, _08085_, _08086_, _08087_, _08088_, _08089_, _08090_, _08091_, _08092_, _08093_, _08094_, _08095_, _08096_, _08097_, _08098_, _08099_, _08100_, _08101_, _08102_, _08103_, _08104_, _08105_, _08106_, _08107_, _08108_, _08109_, _08110_, _08111_, _08112_, _08113_, _08114_, _08115_, _08116_, _08117_, _08118_, _08119_, _08120_, _08121_, _08122_, _08123_, _08124_, _08125_, _08126_, _08127_, _08128_, _08129_, _08130_, _08131_, _08132_, _08133_, _08134_, _08135_, _08136_, _08137_, _08138_, _08139_, _08140_, _08141_, _08142_, _08143_, _08144_, _08145_, _08146_, _08147_, _08148_, _08149_, _08150_, _08151_, _08152_, _08153_, _08154_, _08155_, _08156_, _08157_, _08158_, _08159_, _08160_, _08161_, _08162_, _08163_, _08164_, _08165_, _08166_, _08167_, _08168_, _08169_, _08170_, _08171_, _08172_, _08173_, _08174_, _08175_, _08176_, _08177_, _08178_, _08179_, _08180_, _08181_, _08182_, _08183_, _08184_, _08185_, _08186_, _08187_, _08188_, _08189_, _08190_, _08191_, _08192_, _08193_, _08194_, _08195_, _08196_, _08197_, _08198_, _08199_, _08200_, _08201_, _08202_, _08203_, _08204_, _08205_, _08206_, _08207_, _08208_, _08209_, _08210_, _08211_, _08212_, _08213_, _08214_, _08215_, _08216_, _08217_, _08218_, _08219_, _08220_, _08221_, _08222_, _08223_, _08224_, _08225_, _08226_, _08227_, _08228_, _08229_, _08230_, _08231_, _08232_, _08233_, _08234_, _08235_, _08236_, _08237_, _08238_, _08239_, _08240_, _08241_, _08242_, _08243_, _08244_, _08245_, _08246_, _08247_, _08248_, _08249_, _08250_, _08251_, _08252_, _08253_, _08254_, _08255_, _08256_, _08257_, _08258_, _08259_, _08260_, _08261_, _08262_, _08263_, _08264_, _08265_, _08266_, _08267_, _08268_, _08269_, _08270_, _08271_, _08272_, _08273_, _08274_, _08275_, _08276_, _08277_, _08278_, _08279_, _08280_, _08281_, _08282_, _08283_, _08284_, _08285_, _08286_, _08287_, _08288_, _08289_, _08290_, _08291_, _08292_, _08293_, _08294_, _08295_, _08296_, _08297_, _08298_, _08299_, _08300_, _08301_, _08302_, _08303_, _08304_, _08305_, _08306_, _08307_, _08308_, _08309_, _08310_, _08311_, _08312_, _08313_, _08314_, _08315_, _08316_, _08317_, _08318_, _08319_, _08320_, _08321_, _08322_, _08323_, _08324_, _08325_, _08326_, _08327_, _08328_, _08329_, _08330_, _08331_, _08332_, _08333_, _08334_, _08335_, _08336_, _08337_, _08338_, _08339_, _08340_, _08341_, _08342_, _08343_, _08344_, _08345_, _08346_, _08347_, _08348_, _08349_, _08350_, _08351_, _08352_, _08353_, _08354_, _08355_, _08356_, _08357_, _08358_, _08359_, _08360_, _08361_, _08362_, _08363_, _08364_, _08365_, _08366_, _08367_, _08368_, _08369_, _08370_, _08371_, _08372_, _08373_, _08374_, _08375_, _08376_, _08377_, _08378_, _08379_, _08380_, _08381_, _08382_, _08383_, _08384_, _08385_, _08386_, _08387_, _08388_, _08389_, _08390_, _08391_, _08392_, _08393_, _08394_, _08395_, _08396_, _08397_, _08398_, _08399_, _08400_, _08401_, _08402_, _08403_, _08404_, _08405_, _08406_, _08407_, _08408_, _08409_, _08410_, _08411_, _08412_, _08413_, _08414_, _08415_, _08416_, _08417_, _08418_, _08419_, _08420_, _08421_, _08422_, _08423_, _08424_, _08425_, _08426_, _08427_, _08428_, _08429_, _08430_, _08431_, _08432_, _08433_, _08434_, _08435_, _08436_, _08437_, _08438_, _08439_, _08440_, _08441_, _08442_, _08443_, _08444_, _08445_, _08446_, _08447_, _08448_, _08449_, _08450_, _08451_, _08452_, _08453_, _08454_, _08455_, _08456_, _08457_, _08458_, _08459_, _08460_, _08461_, _08462_, _08463_, _08464_, _08465_, _08466_, _08467_, _08468_, _08469_, _08470_, _08471_, _08472_, _08473_, _08474_, _08475_, _08476_, _08477_, _08478_, _08479_, _08480_, _08481_, _08482_, _08483_, _08484_, _08485_, _08486_, _08487_, _08488_, _08489_, _08490_, _08491_, _08492_, _08493_, _08494_, _08495_, _08496_, _08497_, _08498_, _08499_, _08500_, _08501_, _08502_, _08503_, _08504_, _08505_, _08506_, _08507_, _08508_, _08509_, _08510_, _08511_, _08512_, _08513_, _08514_, _08515_, _08516_, _08517_, _08518_, _08519_, _08520_, _08521_, _08522_, _08523_, _08524_, _08525_, _08526_, _08527_, _08528_, _08529_, _08530_, _08531_, _08532_, _08533_, _08534_, _08535_, _08536_, _08537_, _08538_, _08539_, _08540_, _08541_, _08542_, _08543_, _08544_, _08545_, _08546_, _08547_, _08548_, _08549_, _08550_, _08551_, _08552_, _08553_, _08554_, _08555_, _08556_, _08557_, _08558_, _08559_, _08560_, _08561_, _08562_, _08563_, _08564_, _08565_, _08566_, _08567_, _08568_, _08569_, _08570_, _08571_, _08572_, _08573_, _08574_, _08575_, _08576_, _08577_, _08578_, _08579_, _08580_, _08581_, _08582_, _08583_, _08584_, _08585_, _08586_, _08587_, _08588_, _08589_, _08590_, _08591_, _08592_, _08593_, _08594_, _08595_, _08596_, _08597_, _08598_, _08599_, _08600_, _08601_, _08602_, _08603_, _08604_, _08605_, _08606_, _08607_, _08608_, _08609_, _08610_, _08611_, _08612_, _08613_, _08614_, _08615_, _08616_, _08617_, _08618_, _08619_, _08620_, _08621_, _08622_, _08623_, _08624_, _08625_, _08626_, _08627_, _08628_, _08629_, _08630_, _08631_, _08632_, _08633_, _08634_, _08635_, _08636_, _08637_, _08638_, _08639_, _08640_, _08641_, _08642_, _08643_, _08644_, _08645_, _08646_, _08647_, _08648_, _08649_, _08650_, _08651_, _08652_, _08653_, _08654_, _08655_, _08656_, _08657_, _08658_, _08659_, _08660_, _08661_, _08662_, _08663_, _08664_, _08665_, _08666_, _08667_, _08668_, _08669_, _08670_, _08671_, _08672_, _08673_, _08674_, _08675_, _08676_, _08677_, _08678_, _08679_, _08680_, _08681_, _08682_, _08683_, _08684_, _08685_, _08686_, _08687_, _08688_, _08689_, _08690_, _08691_, _08692_, _08693_, _08694_, _08695_, _08696_, _08697_, _08698_, _08699_, _08700_, _08701_, _08702_, _08703_, _08704_, _08705_, _08706_, _08707_, _08708_, _08709_, _08710_, _08711_, _08712_, _08713_, _08714_, _08715_, _08716_, _08717_, _08718_, _08719_, _08720_, _08721_, _08722_, _08723_, _08724_, _08725_, _08726_, _08727_, _08728_, _08729_, _08730_, _08731_, _08732_, _08733_, _08734_, _08735_, _08736_, _08737_, _08738_, _08739_, _08740_, _08741_, _08742_, _08743_, _08744_, _08745_, _08746_, _08747_, _08748_, _08749_, _08750_, _08751_, _08752_, _08753_, _08754_, _08755_, _08756_, _08757_, _08758_, _08759_, _08760_, _08761_, _08762_, _08763_, _08764_, _08765_, _08766_, _08767_, _08768_, _08769_, _08770_, _08771_, _08772_, _08773_, _08774_, _08775_, _08776_, _08777_, _08778_, _08779_, _08780_, _08781_, _08782_, _08783_, _08784_, _08785_, _08786_, _08787_, _08788_, _08789_, _08790_, _08791_, _08792_, _08793_, _08794_, _08795_, _08796_, _08797_, _08798_, _08799_, _08800_, _08801_, _08802_, _08803_, _08804_, _08805_, _08806_, _08807_, _08808_, _08809_, _08810_, _08811_, _08812_, _08813_, _08814_, _08815_, _08816_, _08817_, _08818_, _08819_, _08820_, _08821_, _08822_, _08823_, _08824_, _08825_, _08826_, _08827_, _08828_, _08829_, _08830_, _08831_, _08832_, _08833_, _08834_, _08835_, _08836_, _08837_, _08838_, _08839_, _08840_, _08841_, _08842_, _08843_, _08844_, _08845_, _08846_, _08847_, _08848_, _08849_, _08850_, _08851_, _08852_, _08853_, _08854_, _08855_, _08856_, _08857_, _08858_, _08859_, _08860_, _08861_, _08862_, _08863_, _08864_, _08865_, _08866_, _08867_, _08868_, _08869_, _08870_, _08871_, _08872_, _08873_, _08874_, _08875_, _08876_, _08877_, _08878_, _08879_, _08880_, _08881_, _08882_, _08883_, _08884_, _08885_, _08886_, _08887_, _08888_, _08889_, _08890_, _08891_, _08892_, _08893_, _08894_, _08895_, _08896_, _08897_, _08898_, _08899_, _08900_, _08901_, _08902_, _08903_, _08904_, _08905_, _08906_, _08907_, _08908_, _08909_, _08910_, _08911_, _08912_, _08913_, _08914_, _08915_, _08916_, _08917_, _08918_, _08919_, _08920_, _08921_, _08922_, _08923_, _08924_, _08925_, _08926_, _08927_, _08928_, _08929_, _08930_, _08931_, _08932_, _08933_, _08934_, _08935_, _08936_, _08937_, _08938_, _08939_, _08940_, _08941_, _08942_, _08943_, _08944_, _08945_, _08946_, _08947_, _08948_, _08949_, _08950_, _08951_, _08952_, _08953_, _08954_, _08955_, _08956_, _08957_, _08958_, _08959_, _08960_, _08961_, _08962_, _08963_, _08964_, _08965_, _08966_, _08967_, _08968_, _08969_, _08970_, _08971_, _08972_, _08973_, _08974_, _08975_, _08976_, _08977_, _08978_, _08979_, _08980_, _08981_, _08982_, _08983_, _08984_, _08985_, _08986_, _08987_, _08988_, _08989_, _08990_, _08991_, _08992_, _08993_, _08994_, _08995_, _08996_, _08997_, _08998_, _08999_, _09000_, _09001_, _09002_, _09003_, _09004_, _09005_, _09006_, _09007_, _09008_, _09009_, _09010_, _09011_, _09012_, _09013_, _09014_, _09015_, _09016_, _09017_, _09018_, _09019_, _09020_, _09021_, _09022_, _09023_, _09024_, _09025_, _09026_, _09027_, _09028_, _09029_, _09030_, _09031_, _09032_, _09033_, _09034_, _09035_, _09036_, _09037_, _09038_, _09039_, _09040_, _09041_, _09042_, _09043_, _09044_, _09045_, _09046_, _09047_, _09048_, _09049_, _09050_, _09051_, _09052_, _09053_, _09054_, _09055_, _09056_, _09057_, _09058_, _09059_, _09060_, _09061_, _09062_, _09063_, _09064_, _09065_, _09066_, _09067_, _09068_, _09069_, _09070_, _09071_, _09072_, _09073_, _09074_, _09075_, _09076_, _09077_, _09078_, _09079_, _09080_, _09081_, _09082_, _09083_, _09084_, _09085_, _09086_, _09087_, _09088_, _09089_, _09090_, _09091_, _09092_, _09093_, _09094_, _09095_, _09096_, _09097_, _09098_, _09099_, _09100_, _09101_, _09102_, _09103_, _09104_, _09105_, _09106_, _09107_, _09108_, _09109_, _09110_, _09111_, _09112_, _09113_, _09114_, _09115_, _09116_, _09117_, _09118_, _09119_, _09120_, _09121_, _09122_, _09123_, _09124_, _09125_, _09126_, _09127_, _09128_, _09129_, _09130_, _09131_, _09132_, _09133_, _09134_, _09135_, _09136_, _09137_, _09138_, _09139_, _09140_, _09141_, _09142_, _09143_, _09144_, _09145_, _09146_, _09147_, _09148_, _09149_, _09150_, _09151_, _09152_, _09153_, _09154_, _09155_, _09156_, _09157_, _09158_, _09159_, _09160_, _09161_, _09162_, _09163_, _09164_, _09165_, _09166_, _09167_, _09168_, _09169_, _09170_, _09171_, _09172_, _09173_, _09174_, _09175_, _09176_, _09177_, _09178_, _09179_, _09180_, _09181_, _09182_, _09183_, _09184_, _09185_, _09186_, _09187_, _09188_, _09189_, _09190_, _09191_, _09192_, _09193_, _09194_, _09195_, _09196_, _09197_, _09198_, _09199_, _09200_, _09201_, _09202_, _09203_, _09204_, _09205_, _09206_, _09207_, _09208_, _09209_, _09210_, _09211_, _09212_, _09213_, _09214_, _09215_, _09216_, _09217_, _09218_, _09219_, _09220_, _09221_, _09222_, _09223_, _09224_, _09225_, _09226_, _09227_, _09228_, _09229_, _09230_, _09231_, _09232_, _09233_, _09234_, _09235_, _09236_, _09237_, _09238_, _09239_, _09240_, _09241_, _09242_, _09243_, _09244_, _09245_, _09246_, _09247_, _09248_, _09249_, _09250_, _09251_, _09252_, _09253_, _09254_, _09255_, _09256_, _09257_, _09258_, _09259_, _09260_, _09261_, _09262_, _09263_, _09264_, _09265_, _09266_, _09267_, _09268_, _09269_, _09270_, _09271_, _09272_, _09273_, _09274_, _09275_, _09276_, _09277_, _09278_, _09279_, _09280_, _09281_, _09282_, _09283_, _09284_, _09285_, _09286_, _09287_, _09288_, _09289_, _09290_, _09291_, _09292_, _09293_, _09294_, _09295_, _09296_, _09297_, _09298_, _09299_, _09300_, _09301_, _09302_, _09303_, _09304_, _09305_, _09306_, _09307_, _09308_, _09309_, _09310_, _09311_, _09312_, _09313_, _09314_, _09315_, _09316_, _09317_, _09318_, _09319_, _09320_, _09321_, _09322_, _09323_, _09324_, _09325_, _09326_, _09327_, _09328_, _09329_, _09330_, _09331_, _09332_, _09333_, _09334_, _09335_, _09336_, _09337_, _09338_, _09339_, _09340_, _09341_, _09342_, _09343_, _09344_, _09345_, _09346_, _09347_, _09348_, _09349_, _09350_, _09351_, _09352_, _09353_, _09354_, _09355_, _09356_, _09357_, _09358_, _09359_, _09360_, _09361_, _09362_, _09363_, _09364_, _09365_, _09366_, _09367_, _09368_, _09369_, _09370_, _09371_, _09372_, _09373_, _09374_, _09375_, _09376_, _09377_, _09378_, _09379_, _09380_, _09381_, _09382_, _09383_, _09384_, _09385_, _09386_, _09387_, _09388_, _09389_, _09390_, _09391_, _09392_, _09393_, _09394_, _09395_, _09396_, _09397_, _09398_, _09399_, _09400_, _09401_, _09402_, _09403_, _09404_, _09405_, _09406_, _09407_, _09408_, _09409_, _09410_, _09411_, _09412_, _09413_, _09414_, _09415_, _09416_, _09417_, _09418_, _09419_, _09420_, _09421_, _09422_, _09423_, _09424_, _09425_, _09426_, _09427_, _09428_, _09429_, _09430_, _09431_, _09432_, _09433_, _09434_, _09435_, _09436_, _09437_, _09438_, _09439_, _09440_, _09441_, _09442_, _09443_, _09444_, _09445_, _09446_, _09447_, _09448_, _09449_, _09450_, _09451_, _09452_, _09453_, _09454_, _09455_, _09456_, _09457_, _09458_, _09459_, _09460_, _09461_, _09462_, _09463_, _09464_, _09465_, _09466_, _09467_, _09468_, _09469_, _09470_, _09471_, _09472_, _09473_, _09474_, _09475_, _09476_, _09477_, _09478_, _09479_, _09480_, _09481_, _09482_, _09483_, _09484_, _09485_, _09486_, _09487_, _09488_, _09489_, _09490_, _09491_, _09492_, _09493_, _09494_, _09495_, _09496_, _09497_, _09498_, _09499_, _09500_, _09501_, _09502_, _09503_, _09504_, _09505_, _09506_, _09507_, _09508_, _09509_, _09510_, _09511_, _09512_, _09513_, _09514_, _09515_, _09516_, _09517_, _09518_, _09519_, _09520_, _09521_, _09522_, _09523_, _09524_, _09525_, _09526_, _09527_, _09528_, _09529_, _09530_, _09531_, _09532_, _09533_, _09534_, _09535_, _09536_, _09537_, _09538_, _09539_, _09540_, _09541_, _09542_, _09543_, _09544_, _09545_, _09546_, _09547_, _09548_, _09549_, _09550_, _09551_, _09552_, _09553_, _09554_, _09555_, _09556_, _09557_, _09558_, _09559_, _09560_, _09561_, _09562_, _09563_, _09564_, _09565_, _09566_, _09567_, _09568_, _09569_, _09570_, _09571_, _09572_, _09573_, _09574_, _09575_, _09576_, _09577_, _09578_, _09579_, _09580_, _09581_, _09582_, _09583_, _09584_, _09585_, _09586_, _09587_, _09588_, _09589_, _09590_, _09591_, _09592_, _09593_, _09594_, _09595_, _09596_, _09597_, _09598_, _09599_, _09600_, _09601_, _09602_, _09603_, _09604_, _09605_, _09606_, _09607_, _09608_, _09609_, _09610_, _09611_, _09612_, _09613_, _09614_, _09615_, _09616_, _09617_, _09618_, _09619_, _09620_, _09621_, _09622_, _09623_, _09624_, _09625_, _09626_, _09627_, _09628_, _09629_, _09630_, _09631_, _09632_, _09633_, _09634_, _09635_, _09636_, _09637_, _09638_, _09639_, _09640_, _09641_, _09642_, _09643_, _09644_, _09645_, _09646_, _09647_, _09648_, _09649_, _09650_, _09651_, _09652_, _09653_, _09654_, _09655_, _09656_, _09657_, _09658_, _09659_, _09660_, _09661_, _09662_, _09663_, _09664_, _09665_, _09666_, _09667_, _09668_, _09669_, _09670_, _09671_, _09672_, _09673_, _09674_, _09675_, _09676_, _09677_, _09678_, _09679_, _09680_, _09681_, _09682_, _09683_, _09684_, _09685_, _09686_, _09687_, _09688_, _09689_, _09690_, _09691_, _09692_, _09693_, _09694_, _09695_, _09696_, _09697_, _09698_, _09699_, _09700_, _09701_, _09702_, _09703_, _09704_, _09705_, _09706_, _09707_, _09708_, _09709_, _09710_, _09711_, _09712_, _09713_, _09714_, _09715_, _09716_, _09717_, _09718_, _09719_, _09720_, _09721_, _09722_, _09723_, _09724_, _09725_, _09726_, _09727_, _09728_, _09729_, _09730_, _09731_, _09732_, _09733_, _09734_, _09735_, _09736_, _09737_, _09738_, _09739_, _09740_, _09741_, _09742_, _09743_, _09744_, _09745_, _09746_, _09747_, _09748_, _09749_, _09750_, _09751_, _09752_, _09753_, _09754_, _09755_, _09756_, _09757_, _09758_, _09759_, _09760_, _09761_, _09762_, _09763_, _09764_, _09765_, _09766_, _09767_, _09768_, _09769_, _09770_, _09771_, _09772_, _09773_, _09774_, _09775_, _09776_, _09777_, _09778_, _09779_, _09780_, _09781_, _09782_, _09783_, _09784_, _09785_, _09786_, _09787_, _09788_, _09789_, _09790_, _09791_, _09792_, _09793_, _09794_, _09795_, _09796_, _09797_, _09798_, _09799_, _09800_, _09801_, _09802_, _09803_, _09804_, _09805_, _09806_, _09807_, _09808_, _09809_, _09810_, _09811_, _09812_, _09813_, _09814_, _09815_, _09816_, _09817_, _09818_, _09819_, _09820_, _09821_, _09822_, _09823_, _09824_, _09825_, _09826_, _09827_, _09828_, _09829_, _09830_, _09831_, _09832_, _09833_, _09834_, _09835_, _09836_, _09837_, _09838_, _09839_, _09840_, _09841_, _09842_, _09843_, _09844_, _09845_, _09846_, _09847_, _09848_, _09849_, _09850_, _09851_, _09852_, _09853_, _09854_, _09855_, _09856_, _09857_, _09858_, _09859_, _09860_, _09861_, _09862_, _09863_, _09864_, _09865_, _09866_, _09867_, _09868_, _09869_, _09870_, _09871_, _09872_, _09873_, _09874_, _09875_, _09876_, _09877_, _09878_, _09879_, _09880_, _09881_, _09882_, _09883_, _09884_, _09885_, _09886_, _09887_, _09888_, _09889_, _09890_, _09891_, _09892_, _09893_, _09894_, _09895_, _09896_, _09897_, _09898_, _09899_, _09900_, _09901_, _09902_, _09903_, _09904_, _09905_, _09906_, _09907_, _09908_, _09909_, _09910_, _09911_, _09912_, _09913_, _09914_, _09915_, _09916_, _09917_, _09918_, _09919_, _09920_, _09921_, _09922_, _09923_, _09924_, _09925_, _09926_, _09927_, _09928_, _09929_, _09930_, _09931_, _09932_, _09933_, _09934_, _09935_, _09936_, _09937_, _09938_, _09939_, _09940_, _09941_, _09942_, _09943_, _09944_, _09945_, _09946_, _09947_, _09948_, _09949_, _09950_, _09951_, _09952_, _09953_, _09954_, _09955_, _09956_, _09957_, _09958_, _09959_, _09960_, _09961_, _09962_, _09963_, _09964_, _09965_, _09966_, _09967_, _09968_, _09969_, _09970_, _09971_, _09972_, _09973_, _09974_, _09975_, _09976_, _09977_, _09978_, _09979_, _09980_, _09981_, _09982_, _09983_, _09984_, _09985_, _09986_, _09987_, _09988_, _09989_, _09990_, _09991_, _09992_, _09993_, _09994_, _09995_, _09996_, _09997_, _09998_, _09999_, _10000_, _10001_, _10002_, _10003_, _10004_, _10005_, _10006_, _10007_, _10008_, _10009_, _10010_, _10011_, _10012_, _10013_, _10014_, _10015_, _10016_, _10017_, _10018_, _10019_, _10020_, _10021_, _10022_, _10023_, _10024_, _10025_, _10026_, _10027_, _10028_, _10029_, _10030_, _10031_, _10032_, _10033_, _10034_, _10035_, _10036_, _10037_, _10038_, _10039_, _10040_, _10041_, _10042_, _10043_, _10044_, _10045_, _10046_, _10047_, _10048_, _10049_, _10050_, _10051_, _10052_, _10053_, _10054_, _10055_, _10056_, _10057_, _10058_, _10059_, _10060_, _10061_, _10062_, _10063_, _10064_, _10065_, _10066_, _10067_, _10068_, _10069_, _10070_, _10071_, _10072_, _10073_, _10074_, _10075_, _10076_, _10077_, _10078_, _10079_, _10080_, _10081_, _10082_, _10083_, _10084_, _10085_, _10086_, _10087_, _10088_, _10089_, _10090_, _10091_, _10092_, _10093_, _10094_, _10095_, _10096_, _10097_, _10098_, _10099_, _10100_, _10101_, _10102_, _10103_, _10104_, _10105_, _10106_, _10107_, _10108_, _10109_, _10110_, _10111_, _10112_, _10113_, _10114_, _10115_, _10116_, _10117_, _10118_, _10119_, _10120_, _10121_, _10122_, _10123_, _10124_, _10125_, _10126_, _10127_, _10128_, _10129_, _10130_, _10131_, _10132_, _10133_, _10134_, _10135_, _10136_, _10137_, _10138_, _10139_, _10140_, _10141_, _10142_, _10143_, _10144_, _10145_, _10146_, _10147_, _10148_, _10149_, _10150_, _10151_, _10152_, _10153_, _10154_, _10155_, _10156_, _10157_, _10158_, _10159_, _10160_, _10161_, _10162_, _10163_, _10164_, _10165_, _10166_, _10167_, _10168_, _10169_, _10170_, _10171_, _10172_, _10173_, _10174_, _10175_, _10176_, _10177_, _10178_, _10179_, _10180_, _10181_, _10182_, _10183_, _10184_, _10185_, _10186_, _10187_, _10188_, _10189_, _10190_, _10191_, _10192_, _10193_, _10194_, _10195_, _10196_, _10197_, _10198_, _10199_, _10200_, _10201_, _10202_, _10203_, _10204_, _10205_, _10206_, _10207_, _10208_, _10209_, _10210_, _10211_, _10212_, _10213_, _10214_, _10215_, _10216_, _10217_, _10218_, _10219_, _10220_, _10221_, _10222_, _10223_, _10224_, _10225_, _10226_, _10227_, _10228_, _10229_, _10230_, _10231_, _10232_, _10233_, _10234_, _10235_, _10236_, _10237_, _10238_, _10239_, _10240_, _10241_, _10242_, _10243_, _10244_, _10245_, _10246_, _10247_, _10248_, _10249_, _10250_, _10251_, _10252_, _10253_, _10254_, _10255_, _10256_, _10257_, _10258_, _10259_, _10260_, _10261_, _10262_, _10263_, _10264_, _10265_, _10266_, _10267_, _10268_, _10269_, _10270_, _10271_, _10272_, _10273_, _10274_, _10275_, _10276_, _10277_, _10278_, _10279_, _10280_, _10281_, _10282_, _10283_, _10284_, _10285_, _10286_, _10287_, _10288_, _10289_, _10290_, _10291_, _10292_, _10293_, _10294_, _10295_, _10296_, _10297_, _10298_, _10299_, _10300_, _10301_, _10302_, _10303_, _10304_, _10305_, _10306_, _10307_, _10308_, _10309_, _10310_, _10311_, _10312_, _10313_, _10314_, _10315_, _10316_, _10317_, _10318_, _10319_, _10320_, _10321_, _10322_, _10323_, _10324_, _10325_, _10326_, _10327_, _10328_, _10329_, _10330_, _10331_, _10332_, _10333_, _10334_, _10335_, _10336_, _10337_, _10338_, _10339_, _10340_, _10341_, _10342_, _10343_, _10344_, _10345_, _10346_, _10347_, _10348_, _10349_, _10350_, _10351_, _10352_, _10353_, _10354_, _10355_, _10356_, _10357_, _10358_, _10359_, _10360_, _10361_, _10362_, _10363_, _10364_, _10365_, _10366_, _10367_, _10368_, _10369_, _10370_, _10371_, _10372_, _10373_, _10374_, _10375_, _10376_, _10377_, _10378_, _10379_, _10380_, _10381_, _10382_, _10383_, _10384_, _10385_, _10386_, _10387_, _10388_, _10389_, _10390_, _10391_, _10392_, _10393_, _10394_, _10395_, _10396_, _10397_, _10398_, _10399_, _10400_, _10401_, _10402_, _10403_, _10404_, _10405_, _10406_, _10407_, _10408_, _10409_, _10410_, _10411_, _10412_, _10413_, _10414_, _10415_, _10416_, _10417_, _10418_, _10419_, _10420_, _10421_, _10422_, _10423_, _10424_, _10425_, _10426_, _10427_, _10428_, _10429_, _10430_, _10431_, _10432_, _10433_, _10434_, _10435_, _10436_, _10437_, _10438_, _10439_, _10440_, _10441_, _10442_, _10443_, _10444_, _10445_, _10446_, _10447_, _10448_, _10449_, _10450_, _10451_, _10452_, _10453_, _10454_, _10455_, _10456_, _10457_, _10458_, _10459_, _10460_, _10461_, _10462_, _10463_, _10464_, _10465_, _10466_, _10467_, _10468_, _10469_, _10470_, _10471_, _10472_, _10473_, _10474_, _10475_, _10476_, _10477_, _10478_, _10479_, _10480_, _10481_, _10482_, _10483_, _10484_, _10485_, _10486_, _10487_, _10488_, _10489_, _10490_, _10491_, _10492_, _10493_, _10494_, _10495_, _10496_, _10497_, _10498_, _10499_, _10500_, _10501_, _10502_, _10503_, _10504_, _10505_, _10506_, _10507_, _10508_, _10509_, _10510_, _10511_, _10512_, _10513_, _10514_, _10515_, _10516_, _10517_, _10518_, _10519_, _10520_, _10521_, _10522_, _10523_, _10524_, _10525_, _10526_, _10527_, _10528_, _10529_, _10530_, _10531_, _10532_, _10533_, _10534_, _10535_, _10536_, _10537_, _10538_, _10539_, _10540_, _10541_, _10542_, _10543_, _10544_, _10545_, _10546_, _10547_, _10548_, _10549_, _10550_, _10551_, _10552_, _10553_, _10554_, _10555_, _10556_, _10557_, _10558_, _10559_, _10560_, _10561_, _10562_, _10563_, _10564_, _10565_, _10566_, _10567_, _10568_, _10569_, _10570_, _10571_, _10572_, _10573_, _10574_, _10575_, _10576_, _10577_, _10578_, _10579_, _10580_, _10581_, _10582_, _10583_, _10584_, _10585_, _10586_, _10587_, _10588_, _10589_, _10590_, _10591_, _10592_, _10593_, _10594_, _10595_, _10596_, _10597_, _10598_, _10599_, _10600_, _10601_, _10602_, _10603_, _10604_, _10605_, _10606_, _10607_, _10608_, _10609_, _10610_, _10611_, _10612_, _10613_, _10614_, _10615_, _10616_, _10617_, _10618_, _10619_, _10620_, _10621_, _10622_, _10623_, _10624_, _10625_, _10626_, _10627_, _10628_, _10629_, _10630_, _10631_, _10632_, _10633_, _10634_, _10635_, _10636_, _10637_, _10638_, _10639_, _10640_, _10641_, _10642_, _10643_, _10644_, _10645_, _10646_, _10647_, _10648_, _10649_, _10650_, _10651_, _10652_, _10653_, _10654_, _10655_, _10656_, _10657_, _10658_, _10659_, _10660_, _10661_, _10662_, _10663_, _10664_, _10665_, _10666_, _10667_, _10668_, _10669_, _10670_, _10671_, _10672_, _10673_, _10674_, _10675_, _10676_, _10677_, _10678_, _10679_, _10680_, _10681_, _10682_, _10683_, _10684_, _10685_, _10686_, _10687_, _10688_, _10689_, _10690_, _10691_, _10692_, _10693_, _10694_, _10695_, _10696_, _10697_, _10698_, _10699_, _10700_, _10701_, _10702_, _10703_, _10704_, _10705_, _10706_, _10707_, _10708_, _10709_, _10710_, _10711_, _10712_, _10713_, _10714_, _10715_, _10716_, _10717_, _10718_, _10719_, _10720_, _10721_, _10722_, _10723_, _10724_, _10725_, _10726_, _10727_, _10728_, _10729_, _10730_, _10731_, _10732_, _10733_, _10734_, _10735_, _10736_, _10737_, _10738_, _10739_, _10740_, _10741_, _10742_, _10743_, _10744_, _10745_, _10746_, _10747_, _10748_, _10749_, _10750_, _10751_, _10752_, _10753_, _10754_, _10755_, _10756_, _10757_, _10758_, _10759_, _10760_, _10761_, _10762_, _10763_, _10764_, _10765_, _10766_, _10767_, _10768_, _10769_, _10770_, _10771_, _10772_, _10773_, _10774_, _10775_, _10776_, _10777_, _10778_, _10779_, _10780_, _10781_, _10782_, _10783_, _10784_, _10785_, _10786_, _10787_, _10788_, _10789_, _10790_, _10791_, _10792_, _10793_, _10794_, _10795_, _10796_, _10797_, _10798_, _10799_, _10800_, _10801_, _10802_, _10803_, _10804_, _10805_, _10806_, _10807_, _10808_, _10809_, _10810_, _10811_, _10812_, _10813_, _10814_, _10815_, _10816_, _10817_, _10818_, _10819_, _10820_, _10821_, _10822_, _10823_, _10824_, _10825_, _10826_, _10827_, _10828_, _10829_, _10830_, _10831_, _10832_, _10833_, _10834_, _10835_, _10836_, _10837_, _10838_, _10839_, _10840_, _10841_, _10842_, _10843_, _10844_, _10845_, _10846_, _10847_, _10848_, _10849_, _10850_, _10851_, _10852_, _10853_, _10854_, _10855_, _10856_, _10857_, _10858_, _10859_, _10860_, _10861_, _10862_, _10863_, _10864_, _10865_, _10866_, _10867_, _10868_, _10869_, _10870_, _10871_, _10872_, _10873_, _10874_, _10875_, _10876_, _10877_, _10878_, _10879_, _10880_, _10881_, _10882_, _10883_, _10884_, _10885_, _10886_, _10887_, _10888_, _10889_, _10890_, _10891_, _10892_, _10893_, _10894_, _10895_, _10896_, _10897_, _10898_, _10899_, _10900_, _10901_, _10902_, _10903_, _10904_, _10905_, _10906_, _10907_, _10908_, _10909_, _10910_, _10911_, _10912_, _10913_, _10914_, _10915_, _10916_, _10917_, _10918_, _10919_, _10920_, _10921_, _10922_, _10923_, _10924_, _10925_, _10926_, _10927_, _10928_, _10929_, _10930_, _10931_, _10932_, _10933_, _10934_, _10935_, _10936_, _10937_, _10938_, _10939_, _10940_, _10941_, _10942_, _10943_, _10944_, _10945_, _10946_, _10947_, _10948_, _10949_, _10950_, _10951_, _10952_, _10953_, _10954_, _10955_, _10956_, _10957_, _10958_, _10959_, _10960_, _10961_, _10962_, _10963_, _10964_, _10965_, _10966_, _10967_, _10968_, _10969_, _10970_, _10971_, _10972_, _10973_, _10974_, _10975_, _10976_, _10977_, _10978_, _10979_, _10980_, _10981_, _10982_, _10983_, _10984_, _10985_, _10986_, _10987_, _10988_, _10989_, _10990_, _10991_, _10992_, _10993_, _10994_, _10995_, _10996_, _10997_, _10998_, _10999_, _11000_, _11001_, _11002_, _11003_, _11004_, _11005_, _11006_, _11007_, _11008_, _11009_, _11010_, _11011_, _11012_, _11013_, _11014_, _11015_, _11016_, _11017_, _11018_, _11019_, _11020_, _11021_, _11022_, _11023_, _11024_, _11025_, _11026_, _11027_, _11028_, _11029_, _11030_, _11031_, _11032_, _11033_, _11034_, _11035_, _11036_, _11037_, _11038_, _11039_, _11040_, _11041_, _11042_, _11043_, _11044_, _11045_, _11046_, _11047_, _11048_, _11049_, _11050_, _11051_, _11052_, _11053_, _11054_, _11055_, _11056_, _11057_, _11058_, _11059_, _11060_, _11061_, _11062_, _11063_, _11064_, _11065_, _11066_, _11067_, _11068_, _11069_, _11070_, _11071_, _11072_, _11073_, _11074_, _11075_, _11076_, _11077_, _11078_, _11079_, _11080_, _11081_, _11082_, _11083_, _11084_, _11085_, _11086_, _11087_, _11088_, _11089_, _11090_, _11091_, _11092_, _11093_, _11094_, _11095_, _11096_, _11097_, _11098_, _11099_, _11100_, _11101_, _11102_, _11103_, _11104_, _11105_, _11106_, _11107_, _11108_, _11109_, _11110_, _11111_, _11112_, _11113_, _11114_, _11115_, _11116_, _11117_, _11118_, _11119_, _11120_, _11121_, _11122_, _11123_, _11124_, _11125_, _11126_, _11127_, _11128_, _11129_, _11130_, _11131_, _11132_, _11133_, _11134_, _11135_, _11136_, _11137_, _11138_, _11139_, _11140_, _11141_, _11142_, _11143_, _11144_, _11145_, _11146_, _11147_, _11148_, _11149_, _11150_, _11151_, _11152_, _11153_, _11154_, _11155_, _11156_, _11157_, _11158_, _11159_, _11160_, _11161_, _11162_, _11163_, _11164_, _11165_, _11166_, _11167_, _11168_, _11169_, _11170_, _11171_, _11172_, _11173_, _11174_, _11175_, _11176_, _11177_, _11178_, _11179_, _11180_, _11181_, _11182_, _11183_, _11184_, _11185_, _11186_, _11187_, _11188_, _11189_, _11190_, _11191_, _11192_, _11193_, _11194_, _11195_, _11196_, _11197_, _11198_, _11199_, _11200_, _11201_, _11202_, _11203_, _11204_, _11205_, _11206_, _11207_, _11208_, _11209_, _11210_, _11211_, _11212_, _11213_, _11214_, _11215_, _11216_, _11217_, _11218_, _11219_, _11220_, _11221_, _11222_, _11223_, _11224_, _11225_, _11226_, _11227_, _11228_, _11229_, _11230_, _11231_, _11232_, _11233_, _11234_, _11235_, _11236_, _11237_, _11238_, _11239_, _11240_, _11241_, _11242_, _11243_, _11244_, _11245_, _11246_, _11247_, _11248_, _11249_, _11250_, _11251_, _11252_, _11253_, _11254_, _11255_, _11256_, _11257_, _11258_, _11259_, _11260_, _11261_, _11262_, _11263_, _11264_, _11265_, _11266_, _11267_, _11268_, _11269_, _11270_, _11271_, _11272_, _11273_, _11274_, _11275_, _11276_, _11277_, _11278_, _11279_, _11280_, _11281_, _11282_, _11283_, _11284_, _11285_, _11286_, _11287_, _11288_, _11289_, _11290_, _11291_, _11292_, _11293_, _11294_, _11295_, _11296_, _11297_, _11298_, _11299_, _11300_, _11301_, _11302_, _11303_, _11304_, _11305_, _11306_, _11307_, _11308_, _11309_, _11310_, _11311_, _11312_, _11313_, _11314_, _11315_, _11316_, _11317_, _11318_, _11319_, _11320_, _11321_, _11322_, _11323_, _11324_, _11325_, _11326_, _11327_, _11328_, _11329_, _11330_, _11331_, _11332_, _11333_, _11334_, _11335_, _11336_, _11337_, _11338_, _11339_, _11340_, _11341_, _11342_, _11343_, _11344_, _11345_, _11346_, _11347_, _11348_, _11349_, _11350_, _11351_, _11352_, _11353_, _11354_, _11355_, _11356_, _11357_, _11358_, _11359_, _11360_, _11361_, _11362_, _11363_, _11364_, _11365_, _11366_, _11367_, _11368_, _11369_, _11370_, _11371_, _11372_, _11373_, _11374_, _11375_, _11376_, _11377_, _11378_, _11379_, _11380_, _11381_, _11382_, _11383_, _11384_, _11385_, _11386_, _11387_, _11388_, _11389_, _11390_, _11391_, _11392_, _11393_, _11394_, _11395_, _11396_, _11397_, _11398_, _11399_, _11400_, _11401_, _11402_, _11403_, _11404_, _11405_, _11406_, _11407_, _11408_, _11409_, _11410_, _11411_, _11412_, _11413_, _11414_, _11415_, _11416_, _11417_, _11418_, _11419_, _11420_, _11421_, _11422_, _11423_, _11424_, _11425_, _11426_, _11427_, _11428_, _11429_, _11430_, _11431_, _11432_, _11433_, _11434_, _11435_, _11436_, _11437_, _11438_, _11439_, _11440_, _11441_, _11442_, _11443_, _11444_, _11445_, _11446_, _11447_, _11448_, _11449_, _11450_, _11451_, _11452_, _11453_, _11454_, _11455_, _11456_, _11457_, _11458_, _11459_, _11460_, _11461_, _11462_, _11463_, _11464_, _11465_, _11466_, _11467_, _11468_, _11469_, _11470_, _11471_, _11472_, _11473_, _11474_, _11475_, _11476_, _11477_, _11478_, _11479_, _11480_, _11481_, _11482_, _11483_, _11484_, _11485_, _11486_, _11487_, _11488_, _11489_, _11490_, _11491_, _11492_, _11493_, _11494_, _11495_, _11496_, _11497_, _11498_, _11499_, _11500_, _11501_, _11502_, _11503_, _11504_, _11505_, _11506_, _11507_, _11508_, _11509_, _11510_, _11511_, _11512_, _11513_, _11514_, _11515_, _11516_, _11517_, _11518_, _11519_, _11520_, _11521_, _11522_, _11523_, _11524_, _11525_, _11526_, _11527_, _11528_, _11529_, _11530_, _11531_, _11532_, _11533_, _11534_, _11535_, _11536_, _11537_, _11538_, _11539_, _11540_, _11541_, _11542_, _11543_, _11544_, _11545_, _11546_, _11547_, _11548_, _11549_, _11550_, _11551_, _11552_, _11553_, _11554_, _11555_, _11556_, _11557_, _11558_, _11559_, _11560_, _11561_, _11562_, _11563_, _11564_, _11565_, _11566_, _11567_, _11568_, _11569_, _11570_, _11571_, _11572_, _11573_, _11574_, _11575_, _11576_, _11577_, _11578_, _11579_, _11580_, _11581_, _11582_, _11583_, _11584_, _11585_, _11586_, _11587_, _11588_, _11589_, _11590_, _11591_, _11592_, _11593_, _11594_, _11595_, _11596_, _11597_, _11598_, _11599_, _11600_, _11601_, _11602_, _11603_, _11604_, _11605_, _11606_, _11607_, _11608_, _11609_, _11610_, _11611_, _11612_, _11613_, _11614_, _11615_, _11616_, _11617_, _11618_, _11619_, _11620_, _11621_, _11622_, _11623_, _11624_, _11625_, _11626_, _11627_, _11628_, _11629_, _11630_, _11631_, _11632_, _11633_, _11634_, _11635_, _11636_, _11637_, _11638_, _11639_, _11640_, _11641_, _11642_, _11643_, _11644_, _11645_, _11646_, _11647_, _11648_, _11649_, _11650_, _11651_, _11652_, _11653_, _11654_, _11655_, _11656_, _11657_, _11658_, _11659_, _11660_, _11661_, _11662_, _11663_, _11664_, _11665_, _11666_, _11667_, _11668_, _11669_, _11670_, _11671_, _11672_, _11673_, _11674_, _11675_, _11676_, _11677_, _11678_, _11679_, _11680_, _11681_, _11682_, _11683_, _11684_, _11685_, _11686_, _11687_, _11688_, _11689_, _11690_, _11691_, _11692_, _11693_, _11694_, _11695_, _11696_, _11697_, _11698_, _11699_, _11700_, _11701_, _11702_, _11703_, _11704_, _11705_, _11706_, _11707_, _11708_, _11709_, _11710_, _11711_, _11712_, _11713_, _11714_, _11715_, _11716_, _11717_, _11718_, _11719_, _11720_, _11721_, _11722_, _11723_, _11724_, _11725_, _11726_, _11727_, _11728_, _11729_, _11730_, _11731_, _11732_, _11733_, _11734_, _11735_, _11736_, _11737_, _11738_, _11739_, _11740_, _11741_, _11742_, _11743_, _11744_, _11745_, _11746_, _11747_, _11748_, _11749_, _11750_, _11751_, _11752_, _11753_, _11754_, _11755_, _11756_, _11757_, _11758_, _11759_, _11760_, _11761_, _11762_, _11763_, _11764_, _11765_, _11766_, _11767_, _11768_, _11769_, _11770_, _11771_, _11772_, _11773_, _11774_, _11775_, _11776_, _11777_, _11778_, _11779_, _11780_, _11781_, _11782_, _11783_, _11784_, _11785_, _11786_, _11787_, _11788_, _11789_, _11790_, _11791_, _11792_, _11793_, _11794_, _11795_, _11796_, _11797_, _11798_, _11799_, _11800_, _11801_, _11802_, _11803_, _11804_, _11805_, _11806_, _11807_, _11808_, _11809_, _11810_, _11811_, _11812_, _11813_, _11814_, _11815_, _11816_, _11817_, _11818_, _11819_, _11820_, _11821_, _11822_, _11823_, _11824_, _11825_, _11826_, _11827_, _11828_, _11829_, _11830_, _11831_, _11832_, _11833_, _11834_, _11835_, _11836_, _11837_, _11838_, _11839_, _11840_, _11841_, _11842_, _11843_, _11844_, _11845_, _11846_, _11847_, _11848_, _11849_, _11850_, _11851_, _11852_, _11853_, _11854_, _11855_, _11856_, _11857_, _11858_, _11859_, _11860_, _11861_, _11862_, _11863_, _11864_, _11865_, _11866_, _11867_, _11868_, _11869_, _11870_, _11871_, _11872_, _11873_, _11874_, _11875_, _11876_, _11877_, _11878_, _11879_, _11880_, _11881_, _11882_, _11883_, _11884_, _11885_, _11886_, _11887_, _11888_, _11889_, _11890_, _11891_, _11892_, _11893_, _11894_, _11895_, _11896_, _11897_, _11898_, _11899_, _11900_, _11901_, _11902_, _11903_, _11904_, _11905_, _11906_, _11907_, _11908_, _11909_, _11910_, _11911_, _11912_, _11913_, _11914_, _11915_, _11916_, _11917_, _11918_, _11919_, _11920_, _11921_, _11922_, _11923_, _11924_, _11925_, _11926_, _11927_, _11928_, _11929_, _11930_, _11931_, _11932_, _11933_, _11934_, _11935_, _11936_, _11937_, _11938_, _11939_, _11940_, _11941_, _11942_, _11943_, _11944_, _11945_, _11946_, _11947_, _11948_, _11949_, _11950_, _11951_, _11952_, _11953_, _11954_, _11955_, _11956_, _11957_, _11958_, _11959_, _11960_, _11961_, _11962_, _11963_, _11964_, _11965_, _11966_, _11967_, _11968_, _11969_, _11970_, _11971_, _11972_, _11973_, _11974_, _11975_, _11976_, _11977_, _11978_, _11979_, _11980_, _11981_, _11982_, _11983_, _11984_, _11985_, _11986_, _11987_, _11988_, _11989_, _11990_, _11991_, _11992_, _11993_, _11994_, _11995_, _11996_, _11997_, _11998_, _11999_, _12000_, _12001_, _12002_, _12003_, _12004_, _12005_, _12006_, _12007_, _12008_, _12009_, _12010_, _12011_, _12012_, _12013_, _12014_, _12015_, _12016_, _12017_, _12018_, _12019_, _12020_, _12021_, _12022_, _12023_, _12024_, _12025_, _12026_, _12027_, _12028_, _12029_, _12030_, _12031_, _12032_, _12033_, _12034_, _12035_, _12036_, _12037_, _12038_, _12039_, _12040_, _12041_, _12042_, _12043_, _12044_, _12045_, _12046_, _12047_, _12048_, _12049_, _12050_, _12051_, _12052_, _12053_, _12054_, _12055_, _12056_, _12057_, _12058_, _12059_, _12060_, _12061_, _12062_, _12063_, _12064_, _12065_, _12066_, _12067_, _12068_, _12069_, _12070_, _12071_, _12072_, _12073_, _12074_, _12075_, _12076_, _12077_, _12078_, _12079_, _12080_, _12081_, _12082_, _12083_, _12084_, _12085_, _12086_, _12087_, _12088_, _12089_, _12090_, _12091_, _12092_, _12093_, _12094_, _12095_, _12096_, _12097_, _12098_, _12099_, _12100_, _12101_, _12102_, _12103_, _12104_, _12105_, _12106_, _12107_, _12108_, _12109_, _12110_, _12111_, _12112_, _12113_, _12114_, _12115_, _12116_, _12117_, _12118_, _12119_, _12120_, _12121_, _12122_, _12123_, _12124_, _12125_, _12126_, _12127_, _12128_, _12129_, _12130_, _12131_, _12132_, _12133_, _12134_, _12135_, _12136_, _12137_, _12138_, _12139_, _12140_, _12141_, _12142_, _12143_, _12144_, _12145_, _12146_, _12147_, _12148_, _12149_, _12150_, _12151_, _12152_, _12153_, _12154_, _12155_, _12156_, _12157_, _12158_, _12159_, _12160_, _12161_, _12162_, _12163_, _12164_, _12165_, _12166_, _12167_, _12168_, _12169_, _12170_, _12171_, _12172_, _12173_, _12174_, _12175_, _12176_, _12177_, _12178_, _12179_, _12180_, _12181_, _12182_, _12183_, _12184_, _12185_, _12186_, _12187_, _12188_, _12189_, _12190_, _12191_, _12192_, _12193_, _12194_, _12195_, _12196_, _12197_, _12198_, _12199_, _12200_, _12201_, _12202_, _12203_, _12204_, _12205_, _12206_, _12207_, _12208_, _12209_, _12210_, _12211_, _12212_, _12213_, _12214_, _12215_, _12216_, _12217_, _12218_, _12219_, _12220_, _12221_, _12222_, _12223_, _12224_, _12225_, _12226_, _12227_, _12228_, _12229_, _12230_, _12231_, _12232_, _12233_, _12234_, _12235_, _12236_, _12237_, _12238_, _12239_, _12240_, _12241_, _12242_, _12243_, _12244_, _12245_, _12246_, _12247_, _12248_, _12249_, _12250_, _12251_, _12252_, _12253_, _12254_, _12255_, _12256_, _12257_, _12258_, _12259_, _12260_, _12261_, _12262_, _12263_, _12264_, _12265_, _12266_, _12267_, _12268_, _12269_, _12270_, _12271_, _12272_, _12273_, _12274_, _12275_, _12276_, _12277_, _12278_, _12279_, _12280_, _12281_, _12282_, _12283_, _12284_, _12285_, _12286_, _12287_, _12288_, _12289_, _12290_, _12291_, _12292_, _12293_, _12294_, _12295_, _12296_, _12297_, _12298_, _12299_, _12300_, _12301_, _12302_, _12303_, _12304_, _12305_, _12306_, _12307_, _12308_, _12309_, _12310_, _12311_, _12312_, _12313_, _12314_, _12315_, _12316_, _12317_, _12318_, _12319_, _12320_, _12321_, _12322_, _12323_, _12324_, _12325_, _12326_, _12327_, _12328_, _12329_, _12330_, _12331_, _12332_, _12333_, _12334_, _12335_, _12336_, _12337_, _12338_, _12339_, _12340_, _12341_, _12342_, _12343_, _12344_, _12345_, _12346_, _12347_, _12348_, _12349_, _12350_, _12351_, _12352_, _12353_, _12354_, _12355_, _12356_, _12357_, _12358_, _12359_, _12360_, _12361_, _12362_, _12363_, _12364_, _12365_, _12366_, _12367_, _12368_, _12369_, _12370_, _12371_, _12372_, _12373_, _12374_, _12375_, _12376_, _12377_, _12378_, _12379_, _12380_, _12381_, _12382_, _12383_, _12384_, _12385_, _12386_, _12387_, _12388_, _12389_, _12390_, _12391_, _12392_, _12393_, _12394_, _12395_, _12396_, _12397_, _12398_, _12399_, _12400_, _12401_, _12402_, _12403_, _12404_, _12405_, _12406_, _12407_, _12408_, _12409_, _12410_, _12411_, _12412_, _12413_, _12414_, _12415_, _12416_, _12417_, _12418_, _12419_, _12420_, _12421_, _12422_, _12423_, _12424_, _12425_, _12426_, _12427_, _12428_, _12429_, _12430_, _12431_, _12432_, _12433_, _12434_, _12435_, _12436_, _12437_, _12438_, _12439_, _12440_, _12441_, _12442_, _12443_, _12444_, _12445_, _12446_, _12447_, _12448_, _12449_, _12450_, _12451_, _12452_, _12453_, _12454_, _12455_, _12456_, _12457_, _12458_, _12459_, _12460_, _12461_, _12462_, _12463_, _12464_, _12465_, _12466_, _12467_, _12468_, _12469_, _12470_, _12471_, _12472_, _12473_, _12474_, _12475_, _12476_, _12477_, _12478_, _12479_, _12480_, _12481_, _12482_, _12483_, _12484_, _12485_, _12486_, _12487_, _12488_, _12489_, _12490_, _12491_, _12492_, _12493_, _12494_, _12495_, _12496_, _12497_, _12498_, _12499_, _12500_, _12501_, _12502_, _12503_, _12504_, _12505_, _12506_, _12507_, _12508_, _12509_, _12510_, _12511_, _12512_, _12513_, _12514_, _12515_, _12516_, _12517_, _12518_, _12519_, _12520_, _12521_, _12522_, _12523_, _12524_, _12525_, _12526_, _12527_, _12528_, _12529_, _12530_, _12531_, _12532_, _12533_, _12534_, _12535_, _12536_, _12537_, _12538_, _12539_, _12540_, _12541_, _12542_, _12543_, _12544_, _12545_, _12546_, _12547_, _12548_, _12549_, _12550_, _12551_, _12552_, _12553_, _12554_, _12555_, _12556_, _12557_, _12558_, _12559_, _12560_, _12561_, _12562_, _12563_, _12564_, _12565_, _12566_, _12567_, _12568_, _12569_, _12570_, _12571_, _12572_, _12573_, _12574_, _12575_, _12576_, _12577_, _12578_, _12579_, _12580_, _12581_, _12582_, _12583_, _12584_, _12585_, _12586_, _12587_, _12588_, _12589_, _12590_, _12591_, _12592_, _12593_, _12594_, _12595_, _12596_, _12597_, _12598_, _12599_, _12600_, _12601_, _12602_, _12603_, _12604_, _12605_, _12606_, _12607_, _12608_, _12609_, _12610_, _12611_, _12612_, _12613_, _12614_, _12615_, _12616_, _12617_, _12618_, _12619_, _12620_, _12621_, _12622_, _12623_, _12624_, _12625_, _12626_, _12627_, _12628_, _12629_, _12630_, _12631_, _12632_, _12633_, _12634_, _12635_, _12636_, _12637_, _12638_, _12639_, _12640_, _12641_, _12642_, _12643_, _12644_, _12645_, _12646_, _12647_, _12648_, _12649_, _12650_, _12651_, _12652_, _12653_, _12654_, _12655_, _12656_, _12657_, _12658_, _12659_, _12660_, _12661_, _12662_, _12663_, _12664_, _12665_, _12666_, _12667_, _12668_, _12669_, _12670_, _12671_, _12672_, _12673_, _12674_, _12675_, _12676_, _12677_, _12678_, _12679_, _12680_, _12681_, _12682_, _12683_, _12684_, _12685_, _12686_, _12687_, _12688_, _12689_, _12690_, _12691_, _12692_, _12693_, _12694_, _12695_, _12696_, _12697_, _12698_, _12699_, _12700_, _12701_, _12702_, _12703_, _12704_, _12705_, _12706_, _12707_, _12708_, _12709_, _12710_, _12711_, _12712_, _12713_, _12714_, _12715_, _12716_, _12717_, _12718_, _12719_, _12720_, _12721_, _12722_, _12723_, _12724_, _12725_, _12726_, _12727_, _12728_, _12729_, _12730_, _12731_, _12732_, _12733_, _12734_, _12735_, _12736_, _12737_, _12738_, _12739_, _12740_, _12741_, _12742_, _12743_, _12744_, _12745_, _12746_, _12747_, _12748_, _12749_, _12750_, _12751_, _12752_, _12753_, _12754_, _12755_, _12756_, _12757_, _12758_, _12759_, _12760_, _12761_, _12762_, _12763_, _12764_, _12765_, _12766_, _12767_, _12768_, _12769_, _12770_, _12771_, _12772_, _12773_, _12774_, _12775_, _12776_, _12777_, _12778_, _12779_, _12780_, _12781_, _12782_, _12783_, _12784_, _12785_, _12786_, _12787_, _12788_, _12789_, _12790_, _12791_, _12792_, _12793_, _12794_, _12795_, _12796_, _12797_, _12798_, _12799_, _12800_, _12801_, _12802_, _12803_, _12804_, _12805_, _12806_, _12807_, _12808_, _12809_, _12810_, _12811_, _12812_, _12813_, _12814_, _12815_, _12816_, _12817_, _12818_, _12819_, _12820_, _12821_, _12822_, _12823_, _12824_, _12825_, _12826_, _12827_, _12828_, _12829_, _12830_, _12831_, _12832_, _12833_, _12834_, _12835_, _12836_, _12837_, _12838_, _12839_, _12840_, _12841_, _12842_, _12843_, _12844_, _12845_, _12846_, _12847_, _12848_, _12849_, _12850_, _12851_, _12852_, _12853_, _12854_, _12855_, _12856_, _12857_, _12858_, _12859_, _12860_, _12861_, _12862_, _12863_, _12864_, _12865_, _12866_, _12867_, _12868_, _12869_, _12870_, _12871_, _12872_, _12873_, _12874_, _12875_, _12876_, _12877_, _12878_, _12879_, _12880_, _12881_, _12882_, _12883_, _12884_, _12885_, _12886_, _12887_, _12888_, _12889_, _12890_, _12891_, _12892_, _12893_, _12894_, _12895_, _12896_, _12897_, _12898_, _12899_, _12900_, _12901_, _12902_, _12903_, _12904_, _12905_, _12906_, _12907_, _12908_, _12909_, _12910_, _12911_, _12912_, _12913_, _12914_, _12915_, _12916_, _12917_, _12918_, _12919_, _12920_, _12921_, _12922_, _12923_, _12924_, _12925_, _12926_, _12927_, _12928_, _12929_, _12930_, _12931_, _12932_, _12933_, _12934_, _12935_, _12936_, _12937_, _12938_, _12939_, _12940_, _12941_, _12942_, _12943_, _12944_, _12945_, _12946_, _12947_, _12948_, _12949_, _12950_, _12951_, _12952_, _12953_, _12954_, _12955_, _12956_, _12957_, _12958_, _12959_, _12960_, _12961_, _12962_, _12963_, _12964_, _12965_, _12966_, _12967_, _12968_, _12969_, _12970_, _12971_, _12972_, _12973_, _12974_, _12975_, _12976_, _12977_, _12978_, _12979_, _12980_, _12981_, _12982_, _12983_, _12984_, _12985_, _12986_, _12987_, _12988_, _12989_, _12990_, _12991_, _12992_, _12993_, _12994_, _12995_, _12996_, _12997_, _12998_, _12999_, _13000_, _13001_, _13002_, _13003_, _13004_, _13005_, _13006_, _13007_, _13008_, _13009_, _13010_, _13011_, _13012_, _13013_, _13014_, _13015_, _13016_, _13017_, _13018_, _13019_, _13020_, _13021_, _13022_, _13023_, _13024_, _13025_, _13026_, _13027_, _13028_, _13029_, _13030_, _13031_, _13032_, _13033_, _13034_, _13035_, _13036_, _13037_, _13038_, _13039_, _13040_, _13041_, _13042_, _13043_, _13044_, _13045_, _13046_, _13047_, _13048_, _13049_, _13050_, _13051_, _13052_, _13053_, _13054_, _13055_, _13056_, _13057_, _13058_, _13059_, _13060_, _13061_, _13062_, _13063_, _13064_, _13065_, _13066_, _13067_, _13068_, _13069_, _13070_, _13071_, _13072_, _13073_, _13074_, _13075_, _13076_, _13077_, _13078_, _13079_, _13080_, _13081_, _13082_, _13083_, _13084_, _13085_, _13086_, _13087_, _13088_, _13089_, _13090_, _13091_, _13092_, _13093_, _13094_, _13095_, _13096_, _13097_, _13098_, _13099_, _13100_, _13101_, _13102_, _13103_, _13104_, _13105_, _13106_, _13107_, _13108_, _13109_, _13110_, _13111_, _13112_, _13113_, _13114_, _13115_, _13116_, _13117_, _13118_, _13119_, _13120_, _13121_, _13122_, _13123_, _13124_, _13125_, _13126_, _13127_, _13128_, _13129_, _13130_, _13131_, _13132_, _13133_, _13134_, _13135_, _13136_, _13137_, _13138_, _13139_, _13140_, _13141_, _13142_, _13143_, _13144_, _13145_, _13146_, _13147_, _13148_, _13149_, _13150_, _13151_, _13152_, _13153_, _13154_, _13155_, _13156_, _13157_, _13158_, _13159_, _13160_, _13161_, _13162_, _13163_, _13164_, _13165_, _13166_, _13167_, _13168_, _13169_, _13170_, _13171_, _13172_, _13173_, _13174_, _13175_, _13176_, _13177_, _13178_, _13179_, _13180_, _13181_, _13182_, _13183_, _13184_, _13185_, _13186_, _13187_, _13188_, _13189_, _13190_, _13191_, _13192_, _13193_, _13194_, _13195_, _13196_, _13197_, _13198_, _13199_, _13200_, _13201_, _13202_, _13203_, _13204_, _13205_, _13206_, _13207_, _13208_, _13209_, _13210_, _13211_, _13212_, _13213_, _13214_, _13215_, _13216_, _13217_, _13218_, _13219_, _13220_, _13221_, _13222_, _13223_, _13224_, _13225_, _13226_, _13227_, _13228_, _13229_, _13230_, _13231_, _13232_, _13233_, _13234_, _13235_, _13236_, _13237_, _13238_, _13239_, _13240_, _13241_, _13242_, _13243_, _13244_, _13245_, _13246_, _13247_, _13248_, _13249_, _13250_, _13251_, _13252_, _13253_, _13254_, _13255_, _13256_, _13257_, _13258_, _13259_, _13260_, _13261_, _13262_, _13263_, _13264_, _13265_, _13266_, _13267_, _13268_, _13269_, _13270_, _13271_, _13272_, _13273_, _13274_, _13275_, _13276_, _13277_, _13278_, _13279_, _13280_, _13281_, _13282_, _13283_, _13284_, _13285_, _13286_, _13287_, _13288_, _13289_, _13290_, _13291_, _13292_, _13293_, _13294_, _13295_, _13296_, _13297_, _13298_, _13299_, _13300_, _13301_, _13302_, _13303_, _13304_, _13305_, _13306_, _13307_, _13308_, _13309_, _13310_, _13311_, _13312_, _13313_, _13314_, _13315_, _13316_, _13317_, _13318_, _13319_, _13320_, _13321_, _13322_, _13323_, _13324_, _13325_, _13326_, _13327_, _13328_, _13329_, _13330_, _13331_, _13332_, _13333_, _13334_, _13335_, _13336_, _13337_, _13338_, _13339_, _13340_, _13341_, _13342_, _13343_, _13344_, _13345_, _13346_, _13347_, _13348_, _13349_, _13350_, _13351_, _13352_, _13353_, _13354_, _13355_, _13356_, _13357_, _13358_, _13359_, _13360_, _13361_, _13362_, _13363_, _13364_, _13365_, _13366_, _13367_, _13368_, _13369_, _13370_, _13371_, _13372_, _13373_, _13374_, _13375_, _13376_, _13377_, _13378_, _13379_, _13380_, _13381_, _13382_, _13383_, _13384_, _13385_, _13386_, _13387_, _13388_, _13389_, _13390_, _13391_, _13392_, _13393_, _13394_, _13395_, _13396_, _13397_, _13398_, _13399_, _13400_, _13401_, _13402_, _13403_, _13404_, _13405_, _13406_, _13407_, _13408_, _13409_, _13410_, _13411_, _13412_, _13413_, _13414_, _13415_, _13416_, _13417_, _13418_, _13419_, _13420_, _13421_, _13422_, _13423_, _13424_, _13425_, _13426_, _13427_, _13428_, _13429_, _13430_, _13431_, _13432_, _13433_, _13434_, _13435_, _13436_, _13437_, _13438_, _13439_, _13440_, _13441_, _13442_, _13443_, _13444_, _13445_, _13446_, _13447_, _13448_, _13449_, _13450_, _13451_, _13452_, _13453_, _13454_, _13455_, _13456_, _13457_, _13458_, _13459_, _13460_, _13461_, _13462_, _13463_, _13464_, _13465_, _13466_, _13467_, _13468_, _13469_, _13470_, _13471_, _13472_, _13473_, _13474_, _13475_, _13476_, _13477_, _13478_, _13479_, _13480_, _13481_, _13482_, _13483_, _13484_, _13485_, _13486_, _13487_, _13488_, _13489_, _13490_, _13491_, _13492_, _13493_, _13494_, _13495_, _13496_, _13497_, _13498_, _13499_, _13500_, _13501_, _13502_, _13503_, _13504_, _13505_, _13506_, _13507_, _13508_, _13509_, _13510_, _13511_, _13512_, _13513_, _13514_, _13515_, _13516_, _13517_, _13518_, _13519_, _13520_, _13521_, _13522_, _13523_, _13524_, _13525_, _13526_, _13527_, _13528_, _13529_, _13530_, _13531_, _13532_, _13533_, _13534_, _13535_, _13536_, _13537_, _13538_, _13539_, _13540_, _13541_, _13542_, _13543_, _13544_, _13545_, _13546_, _13547_, _13548_, _13549_, _13550_, _13551_, _13552_, _13553_, _13554_, _13555_, _13556_, _13557_, _13558_, _13559_, _13560_, _13561_, _13562_, _13563_, _13564_, _13565_, _13566_, _13567_, _13568_, _13569_, _13570_, _13571_, _13572_, _13573_, _13574_, _13575_, _13576_, _13577_, _13578_, _13579_, _13580_, _13581_, _13582_, _13583_, _13584_, _13585_, _13586_, _13587_, _13588_, _13589_, _13590_, _13591_, _13592_, _13593_, _13594_, _13595_, _13596_, _13597_, _13598_, _13599_, _13600_, _13601_, _13602_, _13603_, _13604_, _13605_, _13606_, _13607_, _13608_, _13609_, _13610_, _13611_, _13612_, _13613_, _13614_, _13615_, _13616_, _13617_, _13618_, _13619_, _13620_, _13621_, _13622_, _13623_, _13624_, _13625_, _13626_, _13627_, _13628_, _13629_, _13630_, _13631_, _13632_, _13633_, _13634_, _13635_, _13636_, _13637_, _13638_, _13639_, _13640_, _13641_, _13642_, _13643_, _13644_, _13645_, _13646_, _13647_, _13648_, _13649_, _13650_, _13651_, _13652_, _13653_, _13654_, _13655_, _13656_, _13657_, _13658_, _13659_, _13660_, _13661_, _13662_, _13663_, _13664_, _13665_, _13666_, _13667_, _13668_, _13669_, _13670_, _13671_, _13672_, _13673_, _13674_, _13675_, _13676_, _13677_, _13678_, _13679_, _13680_, _13681_, _13682_, _13683_, _13684_, _13685_, _13686_, _13687_, _13688_, _13689_, _13690_, _13691_, _13692_, _13693_, _13694_, _13695_, _13696_, _13697_, _13698_, _13699_, _13700_, _13701_, _13702_, _13703_, _13704_, _13705_, _13706_, _13707_, _13708_, _13709_, _13710_, _13711_, _13712_, _13713_, _13714_, _13715_, _13716_, _13717_, _13718_, _13719_, _13720_, _13721_, _13722_, _13723_, _13724_, _13725_, _13726_, _13727_, _13728_, _13729_, _13730_, _13731_, _13732_, _13733_, _13734_, _13735_, _13736_, _13737_, _13738_, _13739_, _13740_, _13741_, _13742_, _13743_, _13744_, _13745_, _13746_, _13747_, _13748_, _13749_, _13750_, _13751_, _13752_, _13753_, _13754_, _13755_, _13756_, _13757_, _13758_, _13759_, _13760_, _13761_, _13762_, _13763_, _13764_, _13765_, _13766_, _13767_, _13768_, _13769_, _13770_, _13771_, _13772_, _13773_, _13774_, _13775_, _13776_, _13777_, _13778_, _13779_, _13780_, _13781_, _13782_, _13783_, _13784_, _13785_, _13786_, _13787_, _13788_, _13789_, _13790_, _13791_, _13792_, _13793_, _13794_, _13795_, _13796_, _13797_, _13798_, _13799_, _13800_, _13801_, _13802_, _13803_, _13804_, _13805_, _13806_, _13807_, _13808_, _13809_, _13810_, _13811_, _13812_, _13813_, _13814_, _13815_, _13816_, _13817_, _13818_, _13819_, _13820_, _13821_, _13822_, _13823_, _13824_, _13825_, _13826_, _13827_, _13828_, _13829_, _13830_, _13831_, _13832_, _13833_, _13834_, _13835_, _13836_, _13837_, _13838_, _13839_, _13840_, _13841_, _13842_, _13843_, _13844_, _13845_, _13846_, _13847_, _13848_, _13849_, _13850_, _13851_, _13852_, _13853_, _13854_, _13855_, _13856_, _13857_, _13858_, _13859_, _13860_, _13861_, _13862_, _13863_, _13864_, _13865_, _13866_, _13867_, _13868_, _13869_, _13870_, _13871_, _13872_, _13873_, _13874_, _13875_, _13876_, _13877_, _13878_, _13879_, _13880_, _13881_, _13882_, _13883_, _13884_, _13885_, _13886_, _13887_, _13888_, _13889_, _13890_, _13891_, _13892_, _13893_, _13894_, _13895_, _13896_, _13897_, _13898_, _13899_, _13900_, _13901_, _13902_, _13903_, _13904_, _13905_, _13906_, _13907_, _13908_, _13909_, _13910_, _13911_, _13912_, _13913_, _13914_, _13915_, _13916_, _13917_, _13918_, _13919_, _13920_, _13921_, _13922_, _13923_, _13924_, _13925_, _13926_, _13927_, _13928_, _13929_, _13930_, _13931_, _13932_, _13933_, _13934_, _13935_, _13936_, _13937_, _13938_, _13939_, _13940_, _13941_, _13942_, _13943_, _13944_, _13945_, _13946_, _13947_, _13948_, _13949_, _13950_, _13951_, _13952_, _13953_, _13954_, _13955_, _13956_, _13957_, _13958_, _13959_, _13960_, _13961_, _13962_, _13963_, _13964_, _13965_, _13966_, _13967_, _13968_, _13969_, _13970_, _13971_, _13972_, _13973_, _13974_, _13975_, _13976_, _13977_, _13978_, _13979_, _13980_, _13981_, _13982_, _13983_, _13984_, _13985_, _13986_, _13987_, _13988_, _13989_, _13990_, _13991_, _13992_, _13993_, _13994_, _13995_, _13996_, _13997_, _13998_, _13999_, _14000_, _14001_, _14002_, _14003_, _14004_, _14005_, _14006_, _14007_, _14008_, _14009_, _14010_, _14011_, _14012_, _14013_, _14014_, _14015_, _14016_, _14017_, _14018_, _14019_, _14020_, _14021_, _14022_, _14023_, _14024_, _14025_, _14026_, _14027_, _14028_, _14029_, _14030_, _14031_, _14032_, _14033_, _14034_, _14035_, _14036_, _14037_, _14038_, _14039_, _14040_, _14041_, _14042_, _14043_, _14044_, _14045_, _14046_, _14047_, _14048_, _14049_, _14050_, _14051_, _14052_, _14053_, _14054_, _14055_, _14056_, _14057_, _14058_, _14059_, _14060_, _14061_, _14062_, _14063_, _14064_, _14065_, _14066_, _14067_, _14068_, _14069_, _14070_, _14071_, _14072_, _14073_, _14074_, _14075_, _14076_, _14077_, _14078_, _14079_, _14080_, _14081_, _14082_, _14083_, _14084_, _14085_, _14086_, _14087_, _14088_, _14089_, _14090_, _14091_, _14092_, _14093_, _14094_, _14095_, _14096_, _14097_, _14098_, _14099_, _14100_, _14101_, _14102_, _14103_, _14104_, _14105_, _14106_, _14107_, _14108_, _14109_, _14110_, _14111_, _14112_, _14113_, _14114_, _14115_, _14116_, _14117_, _14118_, _14119_, _14120_, _14121_, _14122_, _14123_, _14124_, _14125_, _14126_, _14127_, _14128_, _14129_, _14130_, _14131_, _14132_, _14133_, _14134_, _14135_, _14136_, _14137_, _14138_, _14139_, _14140_, _14141_, _14142_, _14143_, _14144_, _14145_, _14146_, _14147_, _14148_, _14149_, _14150_, _14151_, _14152_, _14153_, _14154_, _14155_, _14156_, _14157_, _14158_, _14159_, _14160_, _14161_, _14162_, _14163_, _14164_, _14165_, _14166_, _14167_, _14168_, _14169_, _14170_, _14171_, _14172_, _14173_, _14174_, _14175_, _14176_, _14177_, _14178_, _14179_, _14180_, _14181_, _14182_, _14183_, _14184_, _14185_, _14186_, _14187_, _14188_, _14189_, _14190_, _14191_, _14192_, _14193_, _14194_, _14195_, _14196_, _14197_, _14198_, _14199_, _14200_, _14201_, _14202_, _14203_, _14204_, _14205_, _14206_, _14207_, _14208_, _14209_, _14210_, _14211_, _14212_, _14213_, _14214_, _14215_, _14216_, _14217_, _14218_, _14219_, _14220_, _14221_, _14222_, _14223_, _14224_, _14225_, _14226_, _14227_, _14228_, _14229_, _14230_, _14231_, _14232_, _14233_, _14234_, _14235_, _14236_, _14237_, _14238_, _14239_, _14240_, _14241_, _14242_, _14243_, _14244_, _14245_, _14246_, _14247_, _14248_, _14249_, _14250_, _14251_, _14252_, _14253_, _14254_, _14255_, _14256_, _14257_, _14258_, _14259_, _14260_, _14261_, _14262_, _14263_, _14264_, _14265_, _14266_, _14267_, _14268_, _14269_, _14270_, _14271_, _14272_, _14273_, _14274_, _14275_, _14276_, _14277_, _14278_, _14279_, _14280_, _14281_, _14282_, _14283_, _14284_, _14285_, _14286_, _14287_, _14288_, _14289_, _14290_, _14291_, _14292_, _14293_, _14294_, _14295_, _14296_, _14297_, _14298_, _14299_, _14300_, _14301_, _14302_, _14303_, _14304_, _14305_, _14306_, _14307_, _14308_, _14309_, _14310_, _14311_, _14312_, _14313_, _14314_, _14315_, _14316_, _14317_, _14318_, _14319_, _14320_, _14321_, _14322_, _14323_, _14324_, _14325_, _14326_, _14327_, _14328_, _14329_, _14330_, _14331_, _14332_, _14333_, _14334_, _14335_, _14336_, _14337_, _14338_, _14339_, _14340_, _14341_, _14342_, _14343_, _14344_, _14345_, _14346_, _14347_, _14348_, _14349_, _14350_, _14351_, _14352_, _14353_, _14354_, _14355_, _14356_, _14357_, _14358_, _14359_, _14360_, _14361_, _14362_, _14363_, _14364_, _14365_, _14366_, _14367_, _14368_, _14369_, _14370_, _14371_, _14372_, _14373_, _14374_, _14375_, _14376_, _14377_, _14378_, _14379_, _14380_, _14381_, _14382_, _14383_, _14384_, _14385_, _14386_, _14387_, _14388_, _14389_, _14390_, _14391_, _14392_, _14393_, _14394_, _14395_, _14396_, _14397_, _14398_, _14399_, _14400_, _14401_, _14402_, _14403_, _14404_, _14405_, _14406_, _14407_, _14408_, _14409_, _14410_, _14411_, _14412_, _14413_, _14414_, _14415_, _14416_, _14417_, _14418_, _14419_, _14420_, _14421_, _14422_, _14423_, _14424_, _14425_, _14426_, _14427_, _14428_, _14429_, _14430_, _14431_, _14432_, _14433_, _14434_, _14435_, _14436_, _14437_, _14438_, _14439_, _14440_, _14441_, _14442_, _14443_, _14444_, _14445_, _14446_, _14447_, _14448_, _14449_, _14450_, _14451_, _14452_, _14453_, _14454_, _14455_, _14456_, _14457_, _14458_, _14459_, _14460_, _14461_, _14462_, _14463_, _14464_, _14465_, _14466_, _14467_, _14468_, _14469_, _14470_, _14471_, _14472_, _14473_, _14474_, _14475_, _14476_, _14477_, _14478_, _14479_, _14480_, _14481_, _14482_, _14483_, _14484_, _14485_, _14486_, _14487_, _14488_, _14489_, _14490_, _14491_, _14492_, _14493_, _14494_, _14495_, _14496_, _14497_, _14498_, _14499_, _14500_, _14501_, _14502_, _14503_, _14504_, _14505_, _14506_, _14507_, _14508_, _14509_, _14510_, _14511_, _14512_, _14513_, _14514_, _14515_, _14516_, _14517_, _14518_, _14519_, _14520_, _14521_, _14522_, _14523_, _14524_, _14525_, _14526_, _14527_, _14528_, _14529_, _14530_, _14531_, _14532_, _14533_, _14534_, _14535_, _14536_, _14537_, _14538_, _14539_, _14540_, _14541_, _14542_, _14543_, _14544_, _14545_, _14546_, _14547_, _14548_, _14549_, _14550_, _14551_, _14552_, _14553_, _14554_, _14555_, _14556_, _14557_, _14558_, _14559_, _14560_, _14561_, _14562_, _14563_, _14564_, _14565_, _14566_, _14567_, _14568_, _14569_, _14570_, _14571_, _14572_, _14573_, _14574_, _14575_, _14576_, _14577_, _14578_, _14579_, _14580_, _14581_, _14582_, _14583_, _14584_, _14585_, _14586_, _14587_, _14588_, _14589_, _14590_, _14591_, _14592_, _14593_, _14594_, _14595_, _14596_, _14597_, _14598_, _14599_, _14600_, _14601_, _14602_, _14603_, _14604_, _14605_, _14606_, _14607_, _14608_, _14609_, _14610_, _14611_, _14612_, _14613_, _14614_, _14615_, _14616_, _14617_, _14618_, _14619_, _14620_, _14621_, _14622_, _14623_, _14624_, _14625_, _14626_, _14627_, _14628_, _14629_, _14630_, _14631_, _14632_, _14633_, _14634_, _14635_, _14636_, _14637_, _14638_, _14639_, _14640_, _14641_, _14642_, _14643_, _14644_, _14645_, _14646_, _14647_, _14648_, _14649_, _14650_, _14651_, _14652_, _14653_, _14654_, _14655_, _14656_, _14657_, _14658_, _14659_, _14660_, _14661_, _14662_, _14663_, _14664_, _14665_, _14666_, _14667_, _14668_, _14669_, _14670_, _14671_, _14672_, _14673_, _14674_, _14675_, _14676_, _14677_, _14678_, _14679_, _14680_, _14681_, _14682_, _14683_, _14684_, _14685_, _14686_, _14687_, _14688_, _14689_, _14690_, _14691_, _14692_, _14693_, _14694_, _14695_, _14696_, _14697_, _14698_, _14699_, _14700_, _14701_, _14702_, _14703_, _14704_, _14705_, _14706_, _14707_, _14708_, _14709_, _14710_, _14711_, _14712_, _14713_, _14714_, _14715_, _14716_, _14717_, _14718_, _14719_, _14720_, _14721_, _14722_, _14723_, _14724_, _14725_, _14726_, _14727_, _14728_, _14729_, _14730_, _14731_, _14732_, _14733_, _14734_, _14735_, _14736_, _14737_, _14738_, _14739_, _14740_, _14741_, _14742_, _14743_, _14744_, _14745_, _14746_, _14747_, _14748_, _14749_, _14750_, _14751_, _14752_, _14753_, _14754_, _14755_, _14756_, _14757_, _14758_, _14759_, _14760_, _14761_, _14762_, _14763_, _14764_, _14765_, _14766_, _14767_, _14768_, _14769_, _14770_, _14771_, _14772_, _14773_, _14774_, _14775_, _14776_, _14777_, _14778_, _14779_, _14780_, _14781_, _14782_, _14783_, _14784_, _14785_, _14786_, _14787_, _14788_, _14789_, _14790_, _14791_, _14792_, _14793_, _14794_, _14795_, _14796_, _14797_, _14798_, _14799_, _14800_, _14801_, _14802_, _14803_, _14804_, _14805_, _14806_, _14807_, _14808_, _14809_, _14810_, _14811_, _14812_, _14813_, _14814_, _14815_, _14816_, _14817_, _14818_, _14819_, _14820_, _14821_, _14822_, _14823_, _14824_, _14825_, _14826_, _14827_, _14828_, _14829_, _14830_, _14831_, _14832_, _14833_, _14834_, _14835_, _14836_, _14837_, _14838_, _14839_, _14840_, _14841_, _14842_, _14843_, _14844_, _14845_, _14846_, _14847_, _14848_, _14849_, _14850_, _14851_, _14852_, _14853_, _14854_, _14855_, _14856_, _14857_, _14858_, _14859_, _14860_, _14861_, _14862_, _14863_, _14864_, _14865_, _14866_, _14867_, _14868_, _14869_, _14870_, _14871_, _14872_, _14873_, _14874_, _14875_, _14876_, _14877_, _14878_, _14879_, _14880_, _14881_, _14882_, _14883_, _14884_, _14885_, _14886_, _14887_, _14888_, _14889_, _14890_, _14891_, _14892_, _14893_, _14894_, _14895_, _14896_, _14897_, _14898_, _14899_, _14900_, _14901_, _14902_, _14903_, _14904_, _14905_, _14906_, _14907_, _14908_, _14909_, _14910_, _14911_, _14912_, _14913_, _14914_, _14915_, _14916_, _14917_, _14918_, _14919_, _14920_, _14921_, _14922_, _14923_, _14924_, _14925_, _14926_, _14927_, _14928_, _14929_, _14930_, _14931_, _14932_, _14933_, _14934_, _14935_, _14936_, _14937_, _14938_, _14939_, _14940_, _14941_, _14942_, _14943_, _14944_, _14945_, _14946_, _14947_, _14948_, _14949_, _14950_, _14951_, _14952_, _14953_, _14954_, _14955_, _14956_, _14957_, _14958_, _14959_, _14960_, _14961_, _14962_, _14963_, _14964_, _14965_, _14966_, _14967_, _14968_, _14969_, _14970_, _14971_, _14972_, _14973_, _14974_, _14975_, _14976_, _14977_, _14978_, _14979_, _14980_, _14981_, _14982_, _14983_, _14984_, _14985_, _14986_, _14987_, _14988_, _14989_, _14990_, _14991_, _14992_, _14993_, _14994_, _14995_, _14996_, _14997_, _14998_, _14999_, _15000_, _15001_, _15002_, _15003_, _15004_, _15005_, _15006_, _15007_, _15008_, _15009_, _15010_, _15011_, _15012_, _15013_, _15014_, _15015_, _15016_, _15017_, _15018_, _15019_, _15020_, _15021_, _15022_, _15023_, _15024_, _15025_, _15026_, _15027_, _15028_, _15029_, _15030_, _15031_, _15032_, _15033_, _15034_, _15035_, _15036_, _15037_, _15038_, _15039_, _15040_, _15041_, _15042_, _15043_, _15044_, _15045_, _15046_, _15047_, _15048_, _15049_, _15050_, _15051_, _15052_, _15053_, _15054_, _15055_, _15056_, _15057_, _15058_, _15059_, _15060_, _15061_, _15062_, _15063_, _15064_, _15065_, _15066_, _15067_, _15068_, _15069_, _15070_, _15071_, _15072_, _15073_, _15074_, _15075_, _15076_, _15077_, _15078_, _15079_, _15080_, _15081_, _15082_, _15083_, _15084_, _15085_, _15086_, _15087_, _15088_, _15089_, _15090_, _15091_, _15092_, _15093_, _15094_, _15095_, _15096_, _15097_, _15098_, _15099_, _15100_, _15101_, _15102_, _15103_, _15104_, _15105_, _15106_, _15107_, _15108_, _15109_, _15110_, _15111_, _15112_, _15113_, _15114_, _15115_, _15116_, _15117_, _15118_, _15119_, _15120_, _15121_, _15122_, _15123_, _15124_, _15125_, _15126_, _15127_, _15128_, _15129_, _15130_, _15131_, _15132_, _15133_, _15134_, _15135_, _15136_, _15137_, _15138_, _15139_, _15140_, _15141_, _15142_, _15143_, _15144_, _15145_, _15146_, _15147_, _15148_, _15149_, _15150_, _15151_, _15152_, _15153_, _15154_, _15155_, _15156_, _15157_, _15158_, _15159_, _15160_, _15161_, _15162_, _15163_, _15164_, _15165_, _15166_, _15167_, _15168_, _15169_, _15170_, _15171_, _15172_, _15173_, _15174_, _15175_, _15176_, _15177_, _15178_, _15179_, _15180_, _15181_, _15182_, _15183_, _15184_, _15185_, _15186_, _15187_, _15188_, _15189_, _15190_, _15191_, _15192_, _15193_, _15194_, _15195_, _15196_, _15197_, _15198_, _15199_, _15200_, _15201_, _15202_, _15203_, _15204_, _15205_, _15206_, _15207_, _15208_, _15209_, _15210_, _15211_, _15212_, _15213_, _15214_, _15215_, _15216_, _15217_, _15218_, _15219_, _15220_, _15221_, _15222_, _15223_, _15224_, _15225_, _15226_, _15227_, _15228_, _15229_, _15230_, _15231_, _15232_, _15233_, _15234_, _15235_, _15236_, _15237_, _15238_, _15239_, _15240_, _15241_, _15242_, _15243_, _15244_, _15245_, _15246_, _15247_, _15248_, _15249_, _15250_, _15251_, _15252_, _15253_, _15254_, _15255_, _15256_, _15257_, _15258_, _15259_, _15260_, _15261_, _15262_, _15263_, _15264_, _15265_, _15266_, _15267_, _15268_, _15269_, _15270_, _15271_, _15272_, _15273_, _15274_, _15275_, _15276_, _15277_, _15278_, _15279_, _15280_, _15281_, _15282_, _15283_, _15284_, _15285_, _15286_, _15287_, _15288_, _15289_, _15290_, _15291_, _15292_, _15293_, _15294_, _15295_, _15296_, _15297_, _15298_, _15299_, _15300_, _15301_, _15302_, _15303_, _15304_, _15305_, _15306_, _15307_, _15308_, _15309_, _15310_, _15311_, _15312_, _15313_, _15314_, _15315_, _15316_, _15317_, _15318_, _15319_, _15320_, _15321_, _15322_, _15323_, _15324_, _15325_, _15326_, _15327_, _15328_, _15329_, _15330_, _15331_, _15332_, _15333_, _15334_, _15335_, _15336_, _15337_, _15338_, _15339_, _15340_, _15341_, _15342_, _15343_, _15344_, _15345_, _15346_, _15347_, _15348_, _15349_, _15350_, _15351_, _15352_, _15353_, _15354_, _15355_, _15356_, _15357_, _15358_, _15359_, _15360_, _15361_, _15362_, _15363_, _15364_, _15365_, _15366_, _15367_, _15368_, _15369_, _15370_, _15371_, _15372_, _15373_, _15374_, _15375_, _15376_, _15377_, _15378_, _15379_, _15380_, _15381_, _15382_, _15383_, _15384_, _15385_, _15386_, _15387_, _15388_, _15389_, _15390_, _15391_, _15392_, _15393_, _15394_, _15395_, _15396_, _15397_, _15398_, _15399_, _15400_, _15401_, _15402_, _15403_, _15404_, _15405_, _15406_, _15407_, _15408_, _15409_, _15410_, _15411_, _15412_, _15413_, _15414_, _15415_, _15416_, _15417_, _15418_, _15419_, _15420_, _15421_, _15422_, _15423_, _15424_, _15425_, _15426_, _15427_, _15428_, _15429_, _15430_, _15431_, _15432_, _15433_, _15434_, _15435_, _15436_, _15437_, _15438_, _15439_, _15440_, _15441_, _15442_, _15443_, _15444_, _15445_, _15446_, _15447_, _15448_, _15449_, _15450_, _15451_, _15452_, _15453_, _15454_, _15455_, _15456_, _15457_, _15458_, _15459_, _15460_, _15461_, _15462_, _15463_, _15464_, _15465_, _15466_, _15467_, _15468_, _15469_, _15470_, _15471_, _15472_, _15473_, _15474_, _15475_, _15476_, _15477_, _15478_, _15479_, _15480_, _15481_, _15482_, _15483_, _15484_, _15485_, _15486_, _15487_, _15488_, _15489_, _15490_, _15491_, _15492_, _15493_, _15494_, _15495_, _15496_, _15497_, _15498_, _15499_, _15500_, _15501_, _15502_, _15503_, _15504_, _15505_, _15506_, _15507_, _15508_, _15509_, _15510_, _15511_, _15512_, _15513_, _15514_, _15515_, _15516_, _15517_, _15518_, _15519_, _15520_, _15521_, _15522_, _15523_, _15524_, _15525_, _15526_, _15527_, _15528_, _15529_, _15530_, _15531_, _15532_, _15533_, _15534_, _15535_, _15536_, _15537_, _15538_, _15539_, _15540_, _15541_, _15542_, _15543_, _15544_, _15545_, _15546_, _15547_, _15548_, _15549_, _15550_, _15551_, _15552_, _15553_, _15554_, _15555_, _15556_, _15557_, _15558_, _15559_, _15560_, _15561_, _15562_, _15563_, _15564_, _15565_, _15566_, _15567_, _15568_, _15569_, _15570_, _15571_, _15572_, _15573_, _15574_, _15575_, _15576_, _15577_, _15578_, _15579_, _15580_, _15581_, _15582_, _15583_, _15584_, _15585_, _15586_, _15587_, _15588_, _15589_, _15590_, _15591_, _15592_, _15593_, _15594_, _15595_, _15596_, _15597_, _15598_, _15599_, _15600_, _15601_, _15602_, _15603_, _15604_, _15605_, _15606_, _15607_, _15608_, _15609_, _15610_, _15611_, _15612_, _15613_, _15614_, _15615_, _15616_, _15617_, _15618_, _15619_, _15620_, _15621_, _15622_, _15623_, _15624_, _15625_, _15626_, _15627_, _15628_, _15629_, _15630_, _15631_, _15632_, _15633_, _15634_, _15635_, _15636_, _15637_, _15638_, _15639_, _15640_, _15641_, _15642_, _15643_, _15644_, _15645_, _15646_, _15647_, _15648_, _15649_, _15650_, _15651_, _15652_, _15653_, _15654_, _15655_, _15656_, _15657_, _15658_, _15659_, _15660_, _15661_, _15662_, _15663_, _15664_, _15665_, _15666_, _15667_, _15668_, _15669_, _15670_, _15671_, _15672_, _15673_, _15674_, _15675_, _15676_, _15677_, _15678_, _15679_, _15680_, _15681_, _15682_, _15683_, _15684_, _15685_, _15686_, _15687_, _15688_, _15689_, _15690_, _15691_, _15692_, _15693_, _15694_, _15695_, _15696_, _15697_, _15698_, _15699_, _15700_, _15701_, _15702_, _15703_, _15704_, _15705_, _15706_, _15707_, _15708_, _15709_, _15710_, _15711_, _15712_, _15713_, _15714_, _15715_, _15716_, _15717_, _15718_, _15719_, _15720_, _15721_, _15722_, _15723_, _15724_, _15725_, _15726_, _15727_, _15728_, _15729_, _15730_, _15731_, _15732_, _15733_, _15734_, _15735_, _15736_, _15737_, _15738_, _15739_, _15740_, _15741_, _15742_, _15743_, _15744_, _15745_, _15746_, _15747_, _15748_, _15749_, _15750_, _15751_, _15752_, _15753_, _15754_, _15755_, _15756_, _15757_, _15758_, _15759_, _15760_, _15761_, _15762_, _15763_, _15764_, _15765_, _15766_, _15767_, _15768_, _15769_, _15770_, _15771_, _15772_, _15773_, _15774_, _15775_, _15776_, _15777_, _15778_, _15779_, _15780_, _15781_, _15782_, _15783_, _15784_, _15785_, _15786_, _15787_, _15788_, _15789_, _15790_, _15791_, _15792_, _15793_, _15794_, _15795_, _15796_, _15797_, _15798_, _15799_, _15800_, _15801_, _15802_, _15803_, _15804_, _15805_, _15806_, _15807_, _15808_, _15809_, _15810_, _15811_, _15812_, _15813_, _15814_, _15815_, _15816_, _15817_, _15818_, _15819_, _15820_, _15821_, _15822_, _15823_, _15824_, _15825_, _15826_, _15827_, _15828_, _15829_, _15830_, _15831_, _15832_, _15833_, _15834_, _15835_, _15836_, _15837_, _15838_, _15839_, _15840_, _15841_, _15842_, _15843_, _15844_, _15845_, _15846_, _15847_, _15848_, _15849_, _15850_, _15851_, _15852_, _15853_, _15854_, _15855_, _15856_, _15857_, _15858_, _15859_, _15860_, _15861_, _15862_, _15863_, _15864_, _15865_, _15866_, _15867_, _15868_, _15869_, _15870_, _15871_, _15872_, _15873_, _15874_, _15875_, _15876_, _15877_, _15878_, _15879_, _15880_, _15881_, _15882_, _15883_, _15884_, _15885_, _15886_, _15887_, _15888_, _15889_, _15890_, _15891_, _15892_, _15893_, _15894_, _15895_, _15896_, _15897_, _15898_, _15899_, _15900_, _15901_, _15902_, _15903_, _15904_, _15905_, _15906_, _15907_, _15908_, _15909_, _15910_, _15911_, _15912_, _15913_, _15914_, _15915_, _15916_, _15917_, _15918_, _15919_, _15920_, _15921_, _15922_, _15923_, _15924_, _15925_, _15926_, _15927_, _15928_, _15929_, _15930_, _15931_, _15932_, _15933_, _15934_, _15935_, _15936_, _15937_, _15938_, _15939_, _15940_, _15941_, _15942_, _15943_, _15944_, _15945_, _15946_, _15947_, _15948_, _15949_, _15950_, _15951_, _15952_, _15953_, _15954_, _15955_, _15956_, _15957_, _15958_, _15959_, _15960_, _15961_, _15962_, _15963_, _15964_, _15965_, _15966_, _15967_, _15968_, _15969_, _15970_, _15971_, _15972_, _15973_, _15974_, _15975_, _15976_, _15977_, _15978_, _15979_, _15980_, _15981_, _15982_, _15983_, _15984_, _15985_, _15986_, _15987_, _15988_, _15989_, _15990_, _15991_, _15992_, _15993_, _15994_, _15995_, _15996_, _15997_, _15998_, _15999_, _16000_, _16001_, _16002_, _16003_, _16004_, _16005_, _16006_, _16007_, _16008_, _16009_, _16010_, _16011_, _16012_, _16013_, _16014_, _16015_, _16016_, _16017_, _16018_, _16019_, _16020_, _16021_, _16022_, _16023_, _16024_, _16025_, _16026_, _16027_, _16028_, _16029_, _16030_, _16031_, _16032_, _16033_, _16034_, _16035_, _16036_, _16037_, _16038_, _16039_, _16040_, _16041_, _16042_, _16043_, _16044_, _16045_, _16046_, _16047_, _16048_, _16049_, _16050_, _16051_, _16052_, _16053_, _16054_, _16055_, _16056_, _16057_, _16058_, _16059_, _16060_, _16061_, _16062_, _16063_, _16064_, _16065_, _16066_, _16067_, _16068_, _16069_, _16070_, _16071_, _16072_, _16073_, _16074_, _16075_, _16076_, _16077_, _16078_, _16079_, _16080_, _16081_, _16082_, _16083_, _16084_, _16085_, _16086_, _16087_, _16088_, _16089_, _16090_, _16091_, _16092_, _16093_, _16094_, _16095_, _16096_, _16097_, _16098_, _16099_, _16100_, _16101_, _16102_, _16103_, _16104_, _16105_, _16106_, _16107_, _16108_, _16109_, _16110_, _16111_, _16112_, _16113_, _16114_, _16115_, _16116_, _16117_, _16118_, _16119_, _16120_, _16121_, _16122_, _16123_, _16124_, _16125_, _16126_, _16127_, _16128_, _16129_, _16130_, _16131_, _16132_, _16133_, _16134_, _16135_, _16136_, _16137_, _16138_, _16139_, _16140_, _16141_, _16142_, _16143_, _16144_, _16145_, _16146_, _16147_, _16148_, _16149_, _16150_, _16151_, _16152_, _16153_, _16154_, _16155_, _16156_, _16157_, _16158_, _16159_, _16160_, _16161_, _16162_, _16163_, _16164_, _16165_, _16166_, _16167_, _16168_, _16169_, _16170_, _16171_, _16172_, _16173_, _16174_, _16175_, _16176_, _16177_, _16178_, _16179_, _16180_, _16181_, _16182_, _16183_, _16184_, _16185_, _16186_, _16187_, _16188_, _16189_, _16190_, _16191_, _16192_, _16193_, _16194_, _16195_, _16196_, _16197_, _16198_, _16199_, _16200_, _16201_, _16202_, _16203_, _16204_, _16205_, _16206_, _16207_, _16208_, _16209_, _16210_, _16211_, _16212_, _16213_, _16214_, _16215_, _16216_, _16217_, _16218_, _16219_, _16220_, _16221_, _16222_, _16223_, _16224_, _16225_, _16226_, _16227_, _16228_, _16229_, _16230_, _16231_, _16232_, _16233_, _16234_, _16235_, _16236_, _16237_, _16238_, _16239_, _16240_, _16241_, _16242_, _16243_, _16244_, _16245_, _16246_, _16247_, _16248_, _16249_, _16250_, _16251_, _16252_, _16253_, _16254_, _16255_, _16256_, _16257_, _16258_, _16259_, _16260_, _16261_, _16262_, _16263_, _16264_, _16265_, _16266_, _16267_, _16268_, _16269_, _16270_, _16271_, _16272_, _16273_, _16274_, _16275_, _16276_, _16277_, _16278_, _16279_, _16280_, _16281_, _16282_, _16283_, _16284_, _16285_, _16286_, _16287_, _16288_, _16289_, _16290_, _16291_, _16292_, _16293_, _16294_, _16295_, _16296_, _16297_, _16298_, _16299_, _16300_, _16301_, _16302_, _16303_, _16304_, _16305_, _16306_, _16307_, _16308_, _16309_, _16310_, _16311_, _16312_, _16313_, _16314_, _16315_, _16316_, _16317_, _16318_, _16319_, _16320_, _16321_, _16322_, _16323_, _16324_, _16325_, _16326_, _16327_, _16328_, _16329_, _16330_, _16331_, _16332_, _16333_, _16334_, _16335_, _16336_, _16337_, _16338_, _16339_, _16340_, _16341_, _16342_, _16343_, _16344_, _16345_, _16346_, _16347_, _16348_, _16349_, _16350_, _16351_, _16352_, _16353_, _16354_, _16355_, _16356_, _16357_, _16358_, _16359_, _16360_, _16361_, _16362_, _16363_, _16364_, _16365_, _16366_, _16367_, _16368_, _16369_, _16370_, _16371_, _16372_, _16373_, _16374_, _16375_, _16376_, _16377_, _16378_, _16379_, _16380_, _16381_, _16382_, _16383_, _16384_, _16385_, _16386_, _16387_, _16388_, _16389_, _16390_, _16391_, _16392_, _16393_, _16394_, _16395_, _16396_, _16397_, _16398_, _16399_, _16400_, _16401_, _16402_, _16403_, _16404_, _16405_, _16406_, _16407_, _16408_, _16409_, _16410_, _16411_, _16412_, _16413_, _16414_, _16415_, _16416_, _16417_, _16418_, _16419_, _16420_, _16421_, _16422_, _16423_, _16424_, _16425_, _16426_, _16427_, _16428_, _16429_, _16430_, _16431_, _16432_, _16433_, _16434_, _16435_, _16436_, _16437_, _16438_, _16439_, _16440_, _16441_, _16442_, _16443_, _16444_, _16445_, _16446_, _16447_, _16448_, _16449_, _16450_, _16451_, _16452_, _16453_, _16454_, _16455_, _16456_, _16457_, _16458_, _16459_, _16460_, _16461_, _16462_, _16463_, _16464_, _16465_, _16466_, _16467_, _16468_, _16469_, _16470_, _16471_, _16472_, _16473_, _16474_, _16475_, _16476_, _16477_, _16478_, _16479_, _16480_, _16481_, _16482_, _16483_, _16484_, _16485_, _16486_, _16487_, _16488_, _16489_, _16490_, _16491_, _16492_, _16493_, _16494_, _16495_, _16496_, _16497_, _16498_, _16499_, _16500_, _16501_, _16502_, _16503_, _16504_, _16505_, _16506_, _16507_, _16508_, _16509_, _16510_, _16511_, _16512_, _16513_, _16514_, _16515_, _16516_, _16517_, _16518_, _16519_, _16520_, _16521_, _16522_, _16523_, _16524_, _16525_, _16526_, _16527_, _16528_, _16529_, _16530_, _16531_, _16532_, _16533_, _16534_, _16535_, _16536_, _16537_, _16538_, _16539_, _16540_, _16541_, _16542_, _16543_, _16544_, _16545_, _16546_, _16547_, _16548_, _16549_, _16550_, _16551_, _16552_, _16553_, _16554_, _16555_, _16556_, _16557_, _16558_, _16559_, _16560_, _16561_, _16562_, _16563_, _16564_, _16565_, _16566_, _16567_, _16568_, _16569_, _16570_, _16571_, _16572_, _16573_, _16574_, _16575_, _16576_, _16577_, _16578_, _16579_, _16580_, _16581_, _16582_, _16583_, _16584_, _16585_, _16586_, _16587_, _16588_, _16589_, _16590_, _16591_, _16592_, _16593_, _16594_, _16595_, _16596_, _16597_, _16598_, _16599_, _16600_, _16601_, _16602_, _16603_, _16604_, _16605_, _16606_, _16607_, _16608_, _16609_, _16610_, _16611_, _16612_, _16613_, _16614_, _16615_, _16616_, _16617_, _16618_, _16619_, _16620_, _16621_, _16622_, _16623_, _16624_, _16625_, _16626_, _16627_, _16628_, _16629_, _16630_, _16631_, _16632_, _16633_, _16634_, _16635_, _16636_, _16637_, _16638_, _16639_, _16640_, _16641_, _16642_, _16643_, _16644_, _16645_, _16646_, _16647_, _16648_, _16649_, _16650_, _16651_, _16652_, _16653_, _16654_, _16655_, _16656_, _16657_, _16658_, _16659_, _16660_, _16661_, _16662_, _16663_, _16664_, _16665_, _16666_, _16667_, _16668_, _16669_, _16670_, _16671_, _16672_, _16673_, _16674_, _16675_, _16676_, _16677_, _16678_, _16679_, _16680_, _16681_, _16682_, _16683_, _16684_, _16685_, _16686_, _16687_, _16688_, _16689_, _16690_, _16691_, _16692_, _16693_, _16694_, _16695_, _16696_, _16697_, _16698_, _16699_, _16700_, _16701_, _16702_, _16703_, _16704_, _16705_, _16706_, _16707_, _16708_, _16709_, _16710_, _16711_, _16712_, _16713_, _16714_, _16715_, _16716_, _16717_, _16718_, _16719_, _16720_, _16721_, _16722_, _16723_, _16724_, _16725_, _16726_, _16727_, _16728_, _16729_, _16730_, _16731_, _16732_, _16733_, _16734_, _16735_, _16736_, _16737_, _16738_, _16739_, _16740_, _16741_, _16742_, _16743_, _16744_, _16745_, _16746_, _16747_, _16748_, _16749_, _16750_, _16751_, _16752_, _16753_, _16754_, _16755_, _16756_, _16757_, _16758_, _16759_, _16760_, _16761_, _16762_, _16763_, _16764_, _16765_, _16766_, _16767_, _16768_, _16769_, _16770_, _16771_, _16772_, _16773_, _16774_, _16775_, _16776_, _16777_, _16778_, _16779_, _16780_, _16781_, _16782_, _16783_, _16784_, _16785_, _16786_, _16787_, _16788_, _16789_, _16790_, _16791_, _16792_, _16793_, _16794_, _16795_, _16796_, _16797_, _16798_, _16799_, _16800_, _16801_, _16802_, _16803_, _16804_, _16805_, _16806_, _16807_, _16808_, _16809_, _16810_, _16811_, _16812_, _16813_, _16814_, _16815_, _16816_, _16817_, _16818_, _16819_, _16820_, _16821_, _16822_, _16823_, _16824_, _16825_, _16826_, _16827_, _16828_, _16829_, _16830_, _16831_, _16832_, _16833_, _16834_, _16835_, _16836_, _16837_, _16838_, _16839_, _16840_, _16841_, _16842_, _16843_, _16844_, _16845_, _16846_, _16847_, _16848_, _16849_, _16850_, _16851_, _16852_, _16853_, _16854_, _16855_, _16856_, _16857_, _16858_, _16859_, _16860_, _16861_, _16862_, _16863_, _16864_, _16865_, _16866_, _16867_, _16868_, _16869_, _16870_, _16871_, _16872_, _16873_, _16874_, _16875_, _16876_, _16877_, _16878_, _16879_, _16880_, _16881_, _16882_, _16883_, _16884_, _16885_, _16886_, _16887_, _16888_, _16889_, _16890_, _16891_, _16892_, _16893_, _16894_, _16895_, _16896_, _16897_, _16898_, _16899_, _16900_, _16901_, _16902_, _16903_, _16904_, _16905_, _16906_, _16907_, _16908_, _16909_, _16910_, _16911_, _16912_, _16913_, _16914_, _16915_, _16916_, _16917_, _16918_, _16919_, _16920_, _16921_, _16922_, _16923_, _16924_, _16925_, _16926_, _16927_, _16928_, _16929_, _16930_, _16931_, _16932_, _16933_, _16934_, _16935_, _16936_, _16937_, _16938_, _16939_, _16940_, _16941_, _16942_, _16943_, _16944_, _16945_, _16946_, _16947_, _16948_, _16949_, _16950_, _16951_, _16952_, _16953_, _16954_, _16955_, _16956_, _16957_, _16958_, _16959_, _16960_, _16961_, _16962_, _16963_, _16964_, _16965_, _16966_, _16967_, _16968_, _16969_, _16970_, _16971_, _16972_, _16973_, _16974_, _16975_, _16976_, _16977_, _16978_, _16979_, _16980_, _16981_, _16982_, _16983_, _16984_, _16985_, _16986_, _16987_, _16988_, _16989_, _16990_, _16991_, _16992_, _16993_, _16994_, _16995_, _16996_, _16997_, _16998_, _16999_, _17000_, _17001_, _17002_, _17003_, _17004_, _17005_, _17006_, _17007_, _17008_, _17009_, _17010_, _17011_, _17012_, _17013_, _17014_, _17015_, _17016_, _17017_, _17018_, _17019_, _17020_, _17021_, _17022_, _17023_, _17024_, _17025_, _17026_, _17027_, _17028_, _17029_, _17030_, _17031_, _17032_, _17033_, _17034_, _17035_, _17036_, _17037_, _17038_, _17039_, _17040_, _17041_, _17042_, _17043_, _17044_, _17045_, _17046_, _17047_, _17048_, _17049_, _17050_, _17051_, _17052_, _17053_, _17054_, _17055_, _17056_, _17057_, _17058_, _17059_, _17060_, _17061_, _17062_, _17063_, _17064_, _17065_, _17066_, _17067_, _17068_, _17069_, _17070_, _17071_, _17072_, _17073_, _17074_, _17075_, _17076_, _17077_, _17078_, _17079_, _17080_, _17081_, _17082_, _17083_, _17084_, _17085_, _17086_, _17087_, _17088_, _17089_, _17090_, _17091_, _17092_, _17093_, _17094_, _17095_, _17096_, _17097_, _17098_, _17099_, _17100_, _17101_, _17102_, _17103_, _17104_, _17105_, _17106_, _17107_, _17108_, _17109_, _17110_, _17111_, _17112_, _17113_, _17114_, _17115_, _17116_, _17117_, _17118_, _17119_, _17120_, _17121_, _17122_, _17123_, _17124_, _17125_, _17126_, _17127_, _17128_, _17129_, _17130_, _17131_, _17132_, _17133_, _17134_, _17135_, _17136_, _17137_, _17138_, _17139_, _17140_, _17141_, _17142_, _17143_, _17144_, _17145_, _17146_, _17147_, _17148_, _17149_, _17150_, _17151_, _17152_, _17153_, _17154_, _17155_, _17156_, _17157_, _17158_, _17159_, _17160_, _17161_, _17162_, _17163_, _17164_, _17165_, _17166_, _17167_, _17168_, _17169_, _17170_, _17171_, _17172_, _17173_, _17174_, _17175_, _17176_, _17177_, _17178_, _17179_, _17180_, _17181_, _17182_, _17183_, _17184_, _17185_, _17186_, _17187_, _17188_, _17189_, _17190_, _17191_, _17192_, _17193_, _17194_, _17195_, _17196_, _17197_, _17198_, _17199_, _17200_, _17201_, _17202_, _17203_, _17204_, _17205_, _17206_, _17207_, _17208_, _17209_, _17210_, _17211_, _17212_, _17213_, _17214_, _17215_, _17216_, _17217_, _17218_, _17219_, _17220_, _17221_, _17222_, _17223_, _17224_, _17225_, _17226_, _17227_, _17228_, _17229_, _17230_, _17231_, _17232_, _17233_, _17234_, _17235_, _17236_, _17237_, _17238_, _17239_, _17240_, _17241_, _17242_, _17243_, _17244_, _17245_, _17246_, _17247_, _17248_, _17249_, _17250_, _17251_, _17252_, _17253_, _17254_, _17255_, _17256_, _17257_, _17258_, _17259_, _17260_, _17261_, _17262_, _17263_, _17264_, _17265_, _17266_, _17267_, _17268_, _17269_, _17270_, _17271_, _17272_, _17273_, _17274_, _17275_, _17276_, _17277_, _17278_, _17279_, _17280_, _17281_, _17282_, _17283_, _17284_, _17285_, _17286_, _17287_, _17288_, _17289_, _17290_, _17291_, _17292_, _17293_, _17294_, _17295_, _17296_, _17297_, _17298_, _17299_, _17300_, _17301_, _17302_, _17303_, _17304_, _17305_, _17306_, _17307_, _17308_, _17309_, _17310_, _17311_, _17312_, _17313_, _17314_, _17315_, _17316_, _17317_, _17318_, _17319_, _17320_, _17321_, _17322_, _17323_, _17324_, _17325_, _17326_, _17327_, _17328_, _17329_, _17330_, _17331_, _17332_, _17333_, _17334_, _17335_, _17336_, _17337_, _17338_, _17339_, _17340_, _17341_, _17342_, _17343_, _17344_, _17345_, _17346_, _17347_, _17348_, _17349_, _17350_, _17351_, _17352_, _17353_, _17354_, _17355_, _17356_, _17357_, _17358_, _17359_, _17360_, _17361_, _17362_, _17363_, _17364_, _17365_, _17366_, _17367_, _17368_, _17369_, _17370_, _17371_, _17372_, _17373_, _17374_, _17375_, _17376_, _17377_, _17378_, _17379_, _17380_, _17381_, _17382_, _17383_, _17384_, _17385_, _17386_, _17387_, _17388_, _17389_, _17390_, _17391_, _17392_, _17393_, _17394_, _17395_, _17396_, _17397_, _17398_, _17399_, _17400_, _17401_, _17402_, _17403_, _17404_, _17405_, _17406_, _17407_, _17408_, _17409_, _17410_, _17411_, _17412_, _17413_, _17414_, _17415_, _17416_, _17417_, _17418_, _17419_, _17420_, _17421_, _17422_, _17423_, _17424_, _17425_, _17426_, _17427_, _17428_, _17429_, _17430_, _17431_, _17432_, _17433_, _17434_, _17435_, _17436_, _17437_, _17438_, _17439_, _17440_, _17441_, _17442_, _17443_, _17444_, _17445_, _17446_, _17447_, _17448_, _17449_, _17450_, _17451_, _17452_, _17453_, _17454_, _17455_, _17456_, _17457_, _17458_, _17459_, _17460_, _17461_, _17462_, _17463_, _17464_, _17465_, _17466_, _17467_, _17468_, _17469_, _17470_, _17471_, _17472_, _17473_, _17474_, _17475_, _17476_, _17477_, _17478_, _17479_, _17480_, _17481_, _17482_, _17483_, _17484_, _17485_, _17486_, _17487_, _17488_, _17489_, _17490_, _17491_, _17492_, _17493_, _17494_, _17495_, _17496_, _17497_, _17498_, _17499_, _17500_, _17501_, _17502_, _17503_, _17504_, _17505_, _17506_, _17507_, _17508_, _17509_, _17510_, _17511_, _17512_, _17513_, _17514_, _17515_, _17516_, _17517_, _17518_, _17519_, _17520_, _17521_, _17522_, _17523_, _17524_, _17525_, _17526_, _17527_, _17528_, _17529_, _17530_, _17531_, _17532_, _17533_, _17534_, _17535_, _17536_, _17537_, _17538_, _17539_, _17540_, _17541_, _17542_, _17543_, _17544_, _17545_, _17546_, _17547_, _17548_, _17549_, _17550_, _17551_, _17552_, _17553_, _17554_, _17555_, _17556_, _17557_, _17558_, _17559_, _17560_, _17561_, _17562_, _17563_, _17564_, _17565_, _17566_, _17567_, _17568_, _17569_, _17570_, _17571_, _17572_, _17573_, _17574_, _17575_, _17576_, _17577_, _17578_, _17579_, _17580_, _17581_, _17582_, _17583_, _17584_, _17585_, _17586_, _17587_, _17588_, _17589_, _17590_, _17591_, _17592_, _17593_, _17594_, _17595_, _17596_, _17597_, _17598_, _17599_, _17600_, _17601_, _17602_, _17603_, _17604_, _17605_, _17606_, _17607_, _17608_, _17609_, _17610_, _17611_, _17612_, _17613_, _17614_, _17615_, _17616_, _17617_, _17618_, _17619_, _17620_, _17621_, _17622_, _17623_, _17624_, _17625_, _17626_, _17627_, _17628_, _17629_, _17630_, _17631_, _17632_, _17633_, _17634_, _17635_, _17636_, _17637_, _17638_, _17639_, _17640_, _17641_, _17642_, _17643_, _17644_, _17645_, _17646_, _17647_, _17648_, _17649_, _17650_, _17651_, _17652_, _17653_, _17654_, _17655_, _17656_, _17657_, _17658_, _17659_, _17660_, _17661_, _17662_, _17663_, _17664_, _17665_, _17666_, _17667_, _17668_, _17669_, _17670_, _17671_, _17672_, _17673_, _17674_, _17675_, _17676_, _17677_, _17678_, _17679_, _17680_, _17681_, _17682_, _17683_, _17684_, _17685_, _17686_, _17687_, _17688_, _17689_, _17690_, _17691_, _17692_, _17693_, _17694_, _17695_, _17696_, _17697_, _17698_, _17699_, _17700_, _17701_, _17702_, _17703_, _17704_, _17705_, _17706_, _17707_, _17708_, _17709_, _17710_, _17711_, _17712_, _17713_, _17714_, _17715_, _17716_, _17717_, _17718_, _17719_, _17720_, _17721_, _17722_, _17723_, _17724_, _17725_, _17726_, _17727_, _17728_, _17729_, _17730_, _17731_, _17732_, _17733_, _17734_, _17735_, _17736_, _17737_, _17738_, _17739_, _17740_, _17741_, _17742_, _17743_, _17744_, _17745_, _17746_, _17747_, _17748_, _17749_, _17750_, _17751_, _17752_, _17753_, _17754_, _17755_, _17756_, _17757_, _17758_, _17759_, _17760_, _17761_, _17762_, _17763_, _17764_, _17765_, _17766_, _17767_, _17768_, _17769_, _17770_, _17771_, _17772_, _17773_, _17774_, _17775_, _17776_, _17777_, _17778_, _17779_, _17780_, _17781_, _17782_, _17783_, _17784_, _17785_, _17786_, _17787_, _17788_, _17789_, _17790_, _17791_, _17792_, _17793_, _17794_, _17795_, _17796_, _17797_, _17798_, _17799_, _17800_, _17801_, _17802_, _17803_, _17804_, _17805_, _17806_, _17807_, _17808_, _17809_, _17810_, _17811_, _17812_, _17813_, _17814_, _17815_, _17816_, _17817_, _17818_, _17819_, _17820_, _17821_, _17822_, _17823_, _17824_, _17825_, _17826_, _17827_, _17828_, _17829_, _17830_, _17831_, _17832_, _17833_, _17834_, _17835_, _17836_, _17837_, _17838_, _17839_, _17840_, _17841_, _17842_, _17843_, _17844_, _17845_, _17846_, _17847_, _17848_, _17849_, _17850_, _17851_, _17852_, _17853_, _17854_, _17855_, _17856_, _17857_, _17858_, _17859_, _17860_, _17861_, _17862_, _17863_, _17864_, _17865_, _17866_, _17867_, _17868_, _17869_, _17870_, _17871_, _17872_, _17873_, _17874_, _17875_, _17876_, _17877_, _17878_, _17879_, _17880_, _17881_, _17882_, _17883_, _17884_, _17885_, _17886_, _17887_, _17888_, _17889_, _17890_, _17891_, _17892_, _17893_, _17894_, _17895_, _17896_, _17897_, _17898_, _17899_, _17900_, _17901_, _17902_, _17903_, _17904_, _17905_, _17906_, _17907_, _17908_, _17909_, _17910_, _17911_, _17912_, _17913_, _17914_, _17915_, _17916_, _17917_, _17918_, _17919_, _17920_, _17921_, _17922_, _17923_, _17924_, _17925_, _17926_, _17927_, _17928_, _17929_, _17930_, _17931_, _17932_, _17933_, _17934_, _17935_, _17936_, _17937_, _17938_, _17939_, _17940_, _17941_, _17942_, _17943_, _17944_, _17945_, _17946_, _17947_, _17948_, _17949_, _17950_, _17951_, _17952_, _17953_, _17954_, _17955_, _17956_, _17957_, _17958_, _17959_, _17960_, _17961_, _17962_, _17963_, _17964_, _17965_, _17966_, _17967_, _17968_, _17969_, _17970_, _17971_, _17972_, _17973_, _17974_, _17975_, _17976_, _17977_, _17978_, _17979_, _17980_, _17981_, _17982_, _17983_, _17984_, _17985_, _17986_, _17987_, _17988_, _17989_, _17990_, _17991_, _17992_, _17993_, _17994_, _17995_, _17996_, _17997_, _17998_, _17999_, _18000_, _18001_, _18002_, _18003_, _18004_, _18005_, _18006_, _18007_, _18008_, _18009_, _18010_, _18011_, _18012_, _18013_, _18014_, _18015_, _18016_, _18017_, _18018_, _18019_, _18020_, _18021_, _18022_, _18023_, _18024_, _18025_, _18026_, _18027_, _18028_, _18029_, _18030_, _18031_, _18032_, _18033_, _18034_, _18035_, _18036_, _18037_, _18038_, _18039_, _18040_, _18041_, _18042_, _18043_, _18044_, _18045_, _18046_, _18047_, _18048_, _18049_, _18050_, _18051_, _18052_, _18053_, _18054_, _18055_, _18056_, _18057_, _18058_, _18059_, _18060_, _18061_, _18062_, _18063_, _18064_, _18065_, _18066_, _18067_, _18068_, _18069_, _18070_, _18071_, _18072_, _18073_, _18074_, _18075_, _18076_, _18077_, _18078_, _18079_, _18080_, _18081_, _18082_, _18083_, _18084_, _18085_, _18086_, _18087_, _18088_, _18089_, _18090_, _18091_, _18092_, _18093_, _18094_, _18095_, _18096_, _18097_, _18098_, _18099_, _18100_, _18101_, _18102_, _18103_, _18104_, _18105_, _18106_, _18107_, _18108_, _18109_, _18110_, _18111_, _18112_, _18113_, _18114_, _18115_, _18116_, _18117_, _18118_, _18119_, _18120_, _18121_, _18122_, _18123_, _18124_, _18125_, _18126_, _18127_, _18128_, _18129_, _18130_, _18131_, _18132_, _18133_, _18134_, _18135_, _18136_, _18137_, _18138_, _18139_, _18140_, _18141_, _18142_, _18143_, _18144_, _18145_, _18146_, _18147_, _18148_, _18149_, _18150_, _18151_, _18152_, _18153_, _18154_, _18155_, _18156_, _18157_, _18158_, _18159_, _18160_, _18161_, _18162_, _18163_, _18164_, _18165_, _18166_, _18167_, _18168_, _18169_, _18170_, _18171_, _18172_, _18173_, _18174_, _18175_, _18176_, _18177_, _18178_, _18179_, _18180_, _18181_, _18182_, _18183_, _18184_, _18185_, _18186_, _18187_, _18188_, _18189_, _18190_, _18191_, _18192_, _18193_, _18194_, _18195_, _18196_, _18197_, _18198_, _18199_, _18200_, _18201_, _18202_, _18203_, _18204_, _18205_, _18206_, _18207_, _18208_, _18209_, _18210_, _18211_, _18212_, _18213_, _18214_, _18215_, _18216_, _18217_, _18218_, _18219_, _18220_, _18221_, _18222_, _18223_, _18224_, _18225_, _18226_, _18227_, _18228_, _18229_, _18230_, _18231_, _18232_, _18233_, _18234_, _18235_, _18236_, _18237_, _18238_, _18239_, _18240_, _18241_, _18242_, _18243_, _18244_, _18245_, _18246_, _18247_, _18248_, _18249_, _18250_, _18251_, _18252_, _18253_, _18254_, _18255_, _18256_, _18257_, _18258_, _18259_, _18260_, _18261_, _18262_, _18263_, _18264_, _18265_, _18266_, _18267_, _18268_, _18269_, _18270_, _18271_, _18272_, _18273_, _18274_, _18275_, _18276_, _18277_, _18278_, _18279_, _18280_, _18281_, _18282_, _18283_, _18284_, _18285_, _18286_, _18287_, _18288_, _18289_, _18290_, _18291_, _18292_, _18293_, _18294_, _18295_, _18296_, _18297_, _18298_, _18299_, _18300_, _18301_, _18302_, _18303_, _18304_, _18305_, _18306_, _18307_, _18308_, _18309_, _18310_, _18311_, _18312_, _18313_, _18314_, _18315_, _18316_, _18317_, _18318_, _18319_, _18320_, _18321_, _18322_, _18323_, _18324_, _18325_, _18326_, _18327_, _18328_, _18329_, _18330_, _18331_, _18332_, _18333_, _18334_, _18335_, _18336_, _18337_, _18338_, _18339_, _18340_, _18341_, _18342_, _18343_, _18344_, _18345_, _18346_, _18347_, _18348_, _18349_, _18350_, _18351_, _18352_, _18353_, _18354_, _18355_, _18356_, _18357_, _18358_, _18359_, _18360_, _18361_, _18362_, _18363_, _18364_, _18365_, _18366_, _18367_, _18368_, _18369_, _18370_, _18371_, _18372_, _18373_, _18374_, _18375_, _18376_, _18377_, _18378_, _18379_, _18380_, _18381_, _18382_, _18383_, _18384_, _18385_, _18386_, _18387_, _18388_, _18389_, _18390_, _18391_, _18392_, _18393_, _18394_, _18395_, _18396_, _18397_, _18398_, _18399_, _18400_, _18401_, _18402_, _18403_, _18404_, _18405_, _18406_, _18407_, _18408_, _18409_, _18410_, _18411_, _18412_, _18413_, _18414_, _18415_, _18416_, _18417_, _18418_, _18419_, _18420_, _18421_, _18422_, _18423_, _18424_, _18425_, _18426_, _18427_, _18428_, _18429_, _18430_, _18431_, _18432_, _18433_, _18434_, _18435_, _18436_, _18437_, _18438_, _18439_, _18440_, _18441_, _18442_, _18443_, _18444_, _18445_, _18446_, _18447_, _18448_, _18449_, _18450_, _18451_, _18452_, _18453_, _18454_, _18455_, _18456_, _18457_, _18458_, _18459_, _18460_, _18461_, _18462_, _18463_, _18464_, _18465_, _18466_, _18467_, _18468_, _18469_, _18470_, _18471_, _18472_, _18473_, _18474_, _18475_, _18476_, _18477_, _18478_, _18479_, _18480_, _18481_, _18482_, _18483_, _18484_, _18485_, _18486_, _18487_, _18488_, _18489_, _18490_, _18491_, _18492_, _18493_, _18494_, _18495_, _18496_, _18497_, _18498_, _18499_, _18500_, _18501_, _18502_, _18503_, _18504_, _18505_, _18506_, _18507_, _18508_, _18509_, _18510_, _18511_, _18512_, _18513_, _18514_, _18515_, _18516_, _18517_, _18518_, _18519_, _18520_, _18521_, _18522_, _18523_, _18524_, _18525_, _18526_, _18527_, _18528_, _18529_, _18530_, _18531_, _18532_, _18533_, _18534_, _18535_, _18536_, _18537_, _18538_, _18539_, _18540_, _18541_, _18542_, _18543_, _18544_, _18545_, _18546_, _18547_, _18548_, _18549_, _18550_, _18551_, _18552_, _18553_, _18554_, _18555_, _18556_, _18557_, _18558_, _18559_, _18560_, _18561_, _18562_, _18563_, _18564_, _18565_, _18566_, _18567_, _18568_, _18569_, _18570_, _18571_, _18572_, _18573_, _18574_, _18575_, _18576_, _18577_, _18578_, _18579_, _18580_, _18581_, _18582_, _18583_, _18584_, _18585_, _18586_, _18587_, _18588_, _18589_, _18590_, _18591_, _18592_, _18593_, _18594_, _18595_, _18596_, _18597_, _18598_, _18599_, _18600_, _18601_, _18602_, _18603_, _18604_, _18605_, _18606_, _18607_, _18608_, _18609_, _18610_, _18611_, _18612_, _18613_, _18614_, _18615_, _18616_, _18617_, _18618_, _18619_, _18620_, _18621_, _18622_, _18623_, _18624_, _18625_, _18626_, _18627_, _18628_, _18629_, _18630_, _18631_, _18632_, _18633_, _18634_, _18635_, _18636_, _18637_, _18638_, _18639_, _18640_, _18641_, _18642_, _18643_, _18644_, _18645_, _18646_, _18647_, _18648_, _18649_, _18650_, _18651_, _18652_, _18653_, _18654_, _18655_, _18656_, _18657_, _18658_, _18659_, _18660_, _18661_, _18662_, _18663_, _18664_, _18665_, _18666_, _18667_, _18668_, _18669_, _18670_, _18671_, _18672_, _18673_, _18674_, _18675_, _18676_, _18677_, _18678_, _18679_, _18680_, _18681_, _18682_, _18683_, _18684_, _18685_, _18686_, _18687_, _18688_, _18689_, _18690_, _18691_, _18692_, _18693_, _18694_, _18695_, _18696_, _18697_, _18698_, _18699_, _18700_, _18701_, _18702_, _18703_, _18704_, _18705_, _18706_, _18707_, _18708_, _18709_, _18710_, _18711_, _18712_, _18713_, _18714_, _18715_, _18716_, _18717_, _18718_, _18719_, _18720_, _18721_, _18722_, _18723_, _18724_, _18725_, _18726_, _18727_, _18728_, _18729_, _18730_, _18731_, _18732_, _18733_, _18734_, _18735_, _18736_, _18737_, _18738_, _18739_, _18740_, _18741_, _18742_, _18743_, _18744_, _18745_, _18746_, _18747_, _18748_, _18749_, _18750_, _18751_, _18752_, _18753_, _18754_, _18755_, _18756_, _18757_, _18758_, _18759_, _18760_, _18761_, _18762_, _18763_, _18764_, _18765_, _18766_, _18767_, _18768_, _18769_, _18770_, _18771_, _18772_, _18773_, _18774_, _18775_, _18776_, _18777_, _18778_, _18779_, _18780_, _18781_, _18782_, _18783_, _18784_, _18785_, _18786_, _18787_, _18788_, _18789_, _18790_, _18791_, _18792_, _18793_, _18794_, _18795_, _18796_, _18797_, _18798_, _18799_, _18800_, _18801_, _18802_, _18803_, _18804_, _18805_, _18806_, _18807_, _18808_, _18809_, _18810_, _18811_, _18812_, _18813_, _18814_, _18815_, _18816_, _18817_, _18818_, _18819_, _18820_, _18821_, _18822_, _18823_, _18824_, _18825_, _18826_, _18827_, _18828_, _18829_, _18830_, _18831_, _18832_, _18833_, _18834_, _18835_, _18836_, _18837_, _18838_, _18839_, _18840_, _18841_, _18842_, _18843_, _18844_, _18845_, _18846_, _18847_, _18848_, _18849_, _18850_, _18851_, _18852_, _18853_, _18854_, _18855_, _18856_, _18857_, _18858_, _18859_, _18860_, _18861_, _18862_, _18863_, _18864_, _18865_, _18866_, _18867_, _18868_, _18869_, _18870_, _18871_, _18872_, _18873_, _18874_, _18875_, _18876_, _18877_, _18878_, _18879_, _18880_, _18881_, _18882_, _18883_, _18884_, _18885_, _18886_, _18887_, _18888_, _18889_, _18890_, _18891_, _18892_, _18893_, _18894_, _18895_, _18896_, _18897_, _18898_, _18899_, _18900_, _18901_, _18902_, _18903_, _18904_, _18905_, _18906_, _18907_, _18908_, _18909_, _18910_, _18911_, _18912_, _18913_, _18914_, _18915_, _18916_, _18917_, _18918_, _18919_, _18920_, _18921_, _18922_, _18923_, _18924_, _18925_, _18926_, _18927_, _18928_, _18929_, _18930_, _18931_, _18932_, _18933_, _18934_, _18935_, _18936_, _18937_, _18938_, _18939_, _18940_, _18941_, _18942_, _18943_, _18944_, _18945_, _18946_, _18947_, _18948_, _18949_, _18950_, _18951_, _18952_, _18953_, _18954_, _18955_, _18956_, _18957_, _18958_, _18959_, _18960_, _18961_, _18962_, _18963_, _18964_, _18965_, _18966_, _18967_, _18968_, _18969_, _18970_, _18971_, _18972_, _18973_, _18974_, _18975_, _18976_, _18977_, _18978_, _18979_, _18980_, _18981_, _18982_, _18983_, _18984_, _18985_, _18986_, _18987_, _18988_, _18989_, _18990_, _18991_, _18992_, _18993_, _18994_, _18995_, _18996_, _18997_, _18998_, _18999_, _19000_, _19001_, _19002_, _19003_, _19004_, _19005_, _19006_, _19007_, _19008_, _19009_, _19010_, _19011_, _19012_, _19013_, _19014_, _19015_, _19016_, _19017_, _19018_, _19019_, _19020_, _19021_, _19022_, _19023_, _19024_, _19025_, _19026_, _19027_, _19028_, _19029_, _19030_, _19031_, _19032_, _19033_, _19034_, _19035_, _19036_, _19037_, _19038_, _19039_, _19040_, _19041_, _19042_, _19043_, _19044_, _19045_, _19046_, _19047_, _19048_, _19049_, _19050_, _19051_, _19052_, _19053_, _19054_, _19055_, _19056_, _19057_, _19058_, _19059_, _19060_, _19061_, _19062_, _19063_, _19064_, _19065_, _19066_, _19067_, _19068_, _19069_, _19070_, _19071_, _19072_, _19073_, _19074_, _19075_, _19076_, _19077_, _19078_, _19079_, _19080_, _19081_, _19082_, _19083_, _19084_, _19085_, _19086_, _19087_, _19088_, _19089_, _19090_, _19091_, _19092_, _19093_, _19094_, _19095_, _19096_, _19097_, _19098_, _19099_, _19100_, _19101_, _19102_, _19103_, _19104_, _19105_, _19106_, _19107_, _19108_, _19109_, _19110_, _19111_, _19112_, _19113_, _19114_, _19115_, _19116_, _19117_, _19118_, _19119_, _19120_, _19121_, _19122_, _19123_, _19124_, _19125_, _19126_, _19127_, _19128_, _19129_, _19130_, _19131_, _19132_, _19133_, _19134_, _19135_, _19136_, _19137_, _19138_, _19139_, _19140_, _19141_, _19142_, _19143_, _19144_, _19145_, _19146_, _19147_, _19148_, _19149_, _19150_, _19151_, _19152_, _19153_, _19154_, _19155_, _19156_, _19157_, _19158_, _19159_, _19160_, _19161_, _19162_, _19163_, _19164_, _19165_, _19166_, _19167_, _19168_, _19169_, _19170_, _19171_, _19172_, _19173_, _19174_, _19175_, _19176_, _19177_, _19178_, _19179_, _19180_, _19181_, _19182_, _19183_, _19184_, _19185_, _19186_, _19187_, _19188_, _19189_, _19190_, _19191_, _19192_, _19193_, _19194_, _19195_, _19196_, _19197_, _19198_, _19199_, _19200_, _19201_, _19202_, _19203_, _19204_, _19205_, _19206_, _19207_, _19208_, _19209_, _19210_, _19211_, _19212_, _19213_, _19214_, _19215_, _19216_, _19217_, _19218_, _19219_, _19220_, _19221_, _19222_, _19223_, _19224_, _19225_, _19226_, _19227_, _19228_, _19229_, _19230_, _19231_, _19232_, _19233_, _19234_, _19235_, _19236_, _19237_, _19238_, _19239_, _19240_, _19241_, _19242_, _19243_, _19244_, _19245_, _19246_, _19247_, _19248_, _19249_, _19250_, _19251_, _19252_, _19253_, _19254_, _19255_, _19256_, _19257_, _19258_, _19259_, _19260_, _19261_, _19262_, _19263_, _19264_, _19265_, _19266_, _19267_, _19268_, _19269_, _19270_, _19271_, _19272_, _19273_, _19274_, _19275_, _19276_, _19277_, _19278_, _19279_, _19280_, _19281_, _19282_, _19283_, _19284_, _19285_, _19286_, _19287_, _19288_, _19289_, _19290_, _19291_, _19292_, _19293_, _19294_, _19295_, _19296_, _19297_, _19298_, _19299_, _19300_, _19301_, _19302_, _19303_, _19304_, _19305_, _19306_, _19307_, _19308_, _19309_, _19310_, _19311_, _19312_, _19313_, _19314_, _19315_, _19316_, _19317_, _19318_, _19319_, _19320_, _19321_, _19322_, _19323_, _19324_, _19325_, _19326_, _19327_, _19328_, _19329_, _19330_, _19331_, _19332_, _19333_, _19334_, _19335_, _19336_, _19337_, _19338_, _19339_, _19340_, _19341_, _19342_, _19343_, _19344_, _19345_, _19346_, _19347_, _19348_, _19349_, _19350_, _19351_, _19352_, _19353_, _19354_, _19355_, _19356_, _19357_, _19358_, _19359_, _19360_, _19361_, _19362_, _19363_, _19364_, _19365_, _19366_, _19367_, _19368_, _19369_, _19370_, _19371_, _19372_, _19373_, _19374_, _19375_, _19376_, _19377_, _19378_, _19379_, _19380_, _19381_, _19382_, _19383_, _19384_, _19385_, _19386_, _19387_, _19388_, _19389_, _19390_, _19391_, _19392_, _19393_, _19394_, _19395_, _19396_, _19397_, _19398_, _19399_, _19400_, _19401_, _19402_, _19403_, _19404_, _19405_, _19406_, _19407_, _19408_, _19409_, _19410_, _19411_, _19412_, _19413_, _19414_, _19415_, _19416_, _19417_, _19418_, _19419_, _19420_, _19421_, _19422_, _19423_, _19424_, _19425_, _19426_, _19427_, _19428_, _19429_, _19430_, _19431_, _19432_, _19433_, _19434_, _19435_, _19436_, _19437_, _19438_, _19439_, _19440_, _19441_, _19442_, _19443_, _19444_, _19445_, _19446_, _19447_, _19448_, _19449_, _19450_, _19451_, _19452_, _19453_, _19454_, _19455_, _19456_, _19457_, _19458_, _19459_, _19460_, _19461_, _19462_, _19463_, _19464_, _19465_, _19466_, _19467_, _19468_, _19469_, _19470_, _19471_, _19472_, _19473_, _19474_, _19475_, _19476_, _19477_, _19478_, _19479_, _19480_, _19481_, _19482_, _19483_, _19484_, _19485_, _19486_, _19487_, _19488_, _19489_, _19490_, _19491_, _19492_, _19493_, _19494_, _19495_, _19496_, _19497_, _19498_, _19499_, _19500_, _19501_, _19502_, _19503_, _19504_, _19505_, _19506_, _19507_, _19508_, _19509_, _19510_, _19511_, _19512_, _19513_, _19514_, _19515_, _19516_, _19517_, _19518_, _19519_, _19520_, _19521_, _19522_, _19523_, _19524_, _19525_, _19526_, _19527_, _19528_, _19529_, _19530_, _19531_, _19532_, _19533_, _19534_, _19535_, _19536_, _19537_, _19538_, _19539_, _19540_, _19541_, _19542_, _19543_, _19544_, _19545_, _19546_, _19547_, _19548_, _19549_, _19550_, _19551_, _19552_, _19553_, _19554_, _19555_, _19556_, _19557_, _19558_, _19559_, _19560_, _19561_, _19562_, _19563_, _19564_, _19565_, _19566_, _19567_, _19568_, _19569_, _19570_, _19571_, _19572_, _19573_, _19574_, _19575_, _19576_, _19577_, _19578_, _19579_, _19580_, _19581_, _19582_, _19583_, _19584_, _19585_, _19586_, _19587_, _19588_, _19589_, _19590_, _19591_, _19592_, _19593_, _19594_, _19595_, _19596_, _19597_, _19598_, _19599_, _19600_, _19601_, _19602_, _19603_, _19604_, _19605_, _19606_, _19607_, _19608_, _19609_, _19610_, _19611_, _19612_, _19613_, _19614_, _19615_, _19616_, _19617_, _19618_, _19619_, _19620_, _19621_, _19622_, _19623_, _19624_, _19625_, _19626_, _19627_, _19628_, _19629_, _19630_, _19631_, _19632_, _19633_, _19634_, _19635_, _19636_, _19637_, _19638_, _19639_, _19640_, _19641_, _19642_, _19643_, _19644_, _19645_, _19646_, _19647_, _19648_, _19649_, _19650_, _19651_, _19652_, _19653_, _19654_, _19655_, _19656_, _19657_, _19658_, _19659_, _19660_, _19661_, _19662_, _19663_, _19664_, _19665_, _19666_, _19667_, _19668_, _19669_, _19670_, _19671_, _19672_, _19673_, _19674_, _19675_, _19676_, _19677_, _19678_, _19679_, _19680_, _19681_, _19682_, _19683_, _19684_, _19685_, _19686_, _19687_, _19688_, _19689_, _19690_, _19691_, _19692_, _19693_, _19694_, _19695_, _19696_, _19697_, _19698_, _19699_, _19700_, _19701_, _19702_, _19703_, _19704_, _19705_, _19706_, _19707_, _19708_, _19709_, _19710_, _19711_, _19712_, _19713_, _19714_, _19715_, _19716_, _19717_, _19718_, _19719_, _19720_, _19721_, _19722_, _19723_, _19724_, _19725_, _19726_, _19727_, _19728_, _19729_, _19730_, _19731_, _19732_, _19733_, _19734_, _19735_, _19736_, _19737_, _19738_, _19739_, _19740_, _19741_, _19742_, _19743_, _19744_, _19745_, _19746_, _19747_, _19748_, _19749_, _19750_, _19751_, _19752_, _19753_, _19754_, _19755_, _19756_, _19757_, _19758_, _19759_, _19760_, _19761_, _19762_, _19763_, _19764_, _19765_, _19766_, _19767_, _19768_, _19769_, _19770_, _19771_, _19772_, _19773_, _19774_, _19775_, _19776_, _19777_, _19778_, _19779_, _19780_, _19781_, _19782_, _19783_, _19784_, _19785_, _19786_, _19787_, _19788_, _19789_, _19790_, _19791_, _19792_, _19793_, _19794_, _19795_, _19796_, _19797_, _19798_, _19799_, _19800_, _19801_, _19802_, _19803_, _19804_, _19805_, _19806_, _19807_, _19808_, _19809_, _19810_, _19811_, _19812_, _19813_, _19814_, _19815_, _19816_, _19817_, _19818_, _19819_, _19820_, _19821_, _19822_, _19823_, _19824_, _19825_, _19826_, _19827_, _19828_, _19829_, _19830_, _19831_, _19832_, _19833_, _19834_, _19835_, _19836_, _19837_, _19838_, _19839_, _19840_, _19841_, _19842_, _19843_, _19844_, _19845_, _19846_, _19847_, _19848_, _19849_, _19850_, _19851_, _19852_, _19853_, _19854_, _19855_, _19856_, _19857_, _19858_, _19859_, _19860_, _19861_, _19862_, _19863_, _19864_, _19865_, _19866_, _19867_, _19868_, _19869_, _19870_, _19871_, _19872_, _19873_, _19874_, _19875_, _19876_, _19877_, _19878_, _19879_, _19880_, _19881_, _19882_, _19883_, _19884_, _19885_, _19886_, _19887_, _19888_, _19889_, _19890_, _19891_, _19892_, _19893_, _19894_, _19895_, _19896_, _19897_, _19898_, _19899_, _19900_, _19901_, _19902_, _19903_, _19904_, _19905_, _19906_, _19907_, _19908_, _19909_, _19910_, _19911_, _19912_, _19913_, _19914_, _19915_, _19916_, _19917_, _19918_, _19919_, _19920_, _19921_, _19922_, _19923_, _19924_, _19925_, _19926_, _19927_, _19928_, _19929_, _19930_, _19931_, _19932_, _19933_, _19934_, _19935_, _19936_, _19937_, _19938_, _19939_, _19940_, _19941_, _19942_, _19943_, _19944_, _19945_, _19946_, _19947_, _19948_, _19949_, _19950_, _19951_, _19952_, _19953_, _19954_, _19955_, _19956_, _19957_, _19958_, _19959_, _19960_, _19961_, _19962_, _19963_, _19964_, _19965_, _19966_, _19967_, _19968_, _19969_, _19970_, _19971_, _19972_, _19973_, _19974_, _19975_, _19976_, _19977_, _19978_, _19979_, _19980_, _19981_, _19982_, _19983_, _19984_, _19985_, _19986_, _19987_, _19988_, _19989_, _19990_, _19991_, _19992_, _19993_, _19994_, _19995_, _19996_, _19997_, _19998_, _19999_, _20000_, _20001_, _20002_, _20003_, _20004_, _20005_, _20006_, _20007_, _20008_, _20009_, _20010_, _20011_, _20012_, _20013_, _20014_, _20015_, _20016_, _20017_, _20018_, _20019_, _20020_, _20021_, _20022_, _20023_, _20024_, _20025_, _20026_, _20027_, _20028_, _20029_, _20030_, _20031_, _20032_, _20033_, _20034_, _20035_, _20036_, _20037_, _20038_, _20039_, _20040_, _20041_, _20042_, _20043_, _20044_, _20045_, _20046_, _20047_, _20048_, _20049_, _20050_, _20051_, _20052_, _20053_, _20054_, _20055_, _20056_, _20057_, _20058_, _20059_, _20060_, _20061_, _20062_, _20063_, _20064_, _20065_, _20066_, _20067_, _20068_, _20069_, _20070_, _20071_, _20072_, _20073_, _20074_, _20075_, _20076_, _20077_, _20078_, _20079_, _20080_, _20081_, _20082_, _20083_, _20084_, _20085_, _20086_, _20087_, _20088_, _20089_, _20090_, _20091_, _20092_, _20093_, _20094_, _20095_, _20096_, _20097_, _20098_, _20099_, _20100_, _20101_, _20102_, _20103_, _20104_, _20105_, _20106_, _20107_, _20108_, _20109_, _20110_, _20111_, _20112_, _20113_, _20114_, _20115_, _20116_, _20117_, _20118_, _20119_, _20120_, _20121_, _20122_, _20123_, _20124_, _20125_, _20126_, _20127_, _20128_, _20129_, _20130_, _20131_, _20132_, _20133_, _20134_, _20135_, _20136_, _20137_, _20138_, _20139_, _20140_, _20141_, _20142_, _20143_, _20144_, _20145_, _20146_, _20147_, _20148_, _20149_, _20150_, _20151_, _20152_, _20153_, _20154_, _20155_, _20156_, _20157_, _20158_, _20159_, _20160_, _20161_, _20162_, _20163_, _20164_, _20165_, _20166_, _20167_, _20168_, _20169_, _20170_, _20171_, _20172_, _20173_, _20174_, _20175_, _20176_, _20177_, _20178_, _20179_, _20180_, _20181_, _20182_, _20183_, _20184_, _20185_, _20186_, _20187_, _20188_, _20189_, _20190_, _20191_, _20192_, _20193_, _20194_, _20195_, _20196_, _20197_, _20198_, _20199_, _20200_, _20201_, _20202_, _20203_, _20204_, _20205_, _20206_, _20207_, _20208_, _20209_, _20210_, _20211_, _20212_, _20213_, _20214_, _20215_, _20216_, _20217_, _20218_, _20219_, _20220_, _20221_, _20222_, _20223_, _20224_, _20225_, _20226_, _20227_, _20228_, _20229_, _20230_, _20231_, _20232_, _20233_, _20234_, _20235_, _20236_, _20237_, _20238_, _20239_, _20240_, _20241_, _20242_, _20243_, _20244_, _20245_, _20246_, _20247_, _20248_, _20249_, _20250_, _20251_, _20252_, _20253_, _20254_, _20255_, _20256_, _20257_, _20258_, _20259_, _20260_, _20261_, _20262_, _20263_, _20264_, _20265_, _20266_, _20267_, _20268_, _20269_, _20270_, _20271_, _20272_, _20273_, _20274_, _20275_, _20276_, _20277_, _20278_, _20279_, _20280_, _20281_, _20282_, _20283_, _20284_, _20285_, _20286_, _20287_, _20288_, _20289_, _20290_, _20291_, _20292_, _20293_, _20294_, _20295_, _20296_, _20297_, _20298_, _20299_, _20300_, _20301_, _20302_, _20303_, _20304_, _20305_, _20306_, _20307_, _20308_, _20309_, _20310_, _20311_, _20312_, _20313_, _20314_, _20315_, _20316_, _20317_, _20318_, _20319_, _20320_, _20321_, _20322_, _20323_, _20324_, _20325_, _20326_, _20327_, _20328_, _20329_, _20330_, _20331_, _20332_, _20333_, _20334_, _20335_, _20336_, _20337_, _20338_, _20339_, _20340_, _20341_, _20342_, _20343_, _20344_, _20345_, _20346_, _20347_, _20348_, _20349_, _20350_, _20351_, _20352_, _20353_, _20354_, _20355_, _20356_, _20357_, _20358_, _20359_, _20360_, _20361_, _20362_, _20363_, _20364_, _20365_, _20366_, _20367_, _20368_, _20369_, _20370_, _20371_, _20372_, _20373_, _20374_, _20375_, _20376_, _20377_, _20378_, _20379_, _20380_, _20381_, _20382_, _20383_, _20384_, _20385_, _20386_, _20387_, _20388_, _20389_, _20390_, _20391_, _20392_, _20393_, _20394_, _20395_, _20396_, _20397_, _20398_, _20399_, _20400_, _20401_, _20402_, _20403_, _20404_, _20405_, _20406_, _20407_, _20408_, _20409_, _20410_, _20411_, _20412_, _20413_, _20414_, _20415_, _20416_, _20417_, _20418_, _20419_, _20420_, _20421_, _20422_, _20423_, _20424_, _20425_, _20426_, _20427_, _20428_, _20429_, _20430_, _20431_, _20432_, _20433_, _20434_, _20435_, _20436_, _20437_, _20438_, _20439_, _20440_, _20441_, _20442_, _20443_, _20444_, _20445_, _20446_, _20447_, _20448_, _20449_, _20450_, _20451_, _20452_, _20453_, _20454_, _20455_, _20456_, _20457_, _20458_, _20459_, _20460_, _20461_, _20462_, _20463_, _20464_, _20465_, _20466_, _20467_, _20468_, _20469_, _20470_, _20471_, _20472_, _20473_, _20474_, _20475_, _20476_, _20477_, _20478_, _20479_, _20480_, _20481_, _20482_, _20483_, _20484_, _20485_, _20486_, _20487_, _20488_, _20489_, _20490_, _20491_, _20492_, _20493_, _20494_, _20495_, _20496_, _20497_, _20498_, _20499_, _20500_, _20501_, _20502_, _20503_, _20504_, _20505_, _20506_, _20507_, _20508_, _20509_, _20510_, _20511_, _20512_, _20513_, _20514_, _20515_, _20516_, _20517_, _20518_, _20519_, _20520_, _20521_, _20522_, _20523_, _20524_, _20525_, _20526_, _20527_, _20528_, _20529_, _20530_, _20531_, _20532_, _20533_, _20534_, _20535_, _20536_, _20537_, _20538_, _20539_, _20540_, _20541_, _20542_, _20543_, _20544_, _20545_, _20546_, _20547_, _20548_, _20549_, _20550_, _20551_, _20552_, _20553_, _20554_, _20555_, _20556_, _20557_, _20558_, _20559_, _20560_, _20561_, _20562_, _20563_, _20564_, _20565_, _20566_, _20567_, _20568_, _20569_, _20570_, _20571_, _20572_, _20573_, _20574_, _20575_, _20576_, _20577_, _20578_, _20579_, _20580_, _20581_, _20582_, _20583_, _20584_, _20585_, _20586_, _20587_, _20588_, _20589_, _20590_, _20591_, _20592_, _20593_, _20594_, _20595_, _20596_, _20597_, _20598_, _20599_, _20600_, _20601_, _20602_, _20603_, _20604_, _20605_, _20606_, _20607_, _20608_, _20609_, _20610_, _20611_, _20612_, _20613_, _20614_, _20615_, _20616_, _20617_, _20618_, _20619_, _20620_, _20621_, _20622_, _20623_, _20624_, _20625_, _20626_, _20627_, _20628_, _20629_, _20630_, _20631_, _20632_, _20633_, _20634_, _20635_, _20636_, _20637_, _20638_, _20639_, _20640_, _20641_, _20642_, _20643_, _20644_, _20645_, _20646_, _20647_, _20648_, _20649_, _20650_, _20651_, _20652_, _20653_, _20654_, _20655_, _20656_, _20657_, _20658_, _20659_, _20660_, _20661_, _20662_, _20663_, _20664_, _20665_, _20666_, _20667_, _20668_, _20669_, _20670_, _20671_, _20672_, _20673_, _20674_, _20675_, _20676_, _20677_, _20678_, _20679_, _20680_, _20681_, _20682_, _20683_, _20684_, _20685_, _20686_, _20687_, _20688_, _20689_, _20690_, _20691_, _20692_, _20693_, _20694_, _20695_, _20696_, _20697_, _20698_, _20699_, _20700_, _20701_, _20702_, _20703_, _20704_, _20705_, _20706_, _20707_, _20708_, _20709_, _20710_, _20711_, _20712_, _20713_, _20714_, _20715_, _20716_, _20717_, _20718_, _20719_, _20720_, _20721_, _20722_, _20723_, _20724_, _20725_, _20726_, _20727_, _20728_, _20729_, _20730_, _20731_, _20732_, _20733_, _20734_, _20735_, _20736_, _20737_, _20738_, _20739_, _20740_, _20741_, _20742_, _20743_, _20744_, _20745_, _20746_, _20747_, _20748_, _20749_, _20750_, _20751_, _20752_, _20753_, _20754_, _20755_, _20756_, _20757_, _20758_, _20759_, _20760_, _20761_, _20762_, _20763_, _20764_, _20765_, _20766_, _20767_, _20768_, _20769_, _20770_, _20771_, _20772_, _20773_, _20774_, _20775_, _20776_, _20777_, _20778_, _20779_, _20780_, _20781_, _20782_, _20783_, _20784_, _20785_, _20786_, _20787_, _20788_, _20789_, _20790_, _20791_, _20792_, _20793_, _20794_, _20795_, _20796_, _20797_, _20798_, _20799_, _20800_, _20801_, _20802_, _20803_, _20804_, _20805_, _20806_, _20807_, _20808_, _20809_, _20810_, _20811_, _20812_, _20813_, _20814_, _20815_, _20816_, _20817_, _20818_, _20819_, _20820_, _20821_, _20822_, _20823_, _20824_, _20825_, _20826_, _20827_, _20828_, _20829_, _20830_, _20831_, _20832_, _20833_, _20834_, _20835_, _20836_, _20837_, _20838_, _20839_, _20840_, _20841_, _20842_, _20843_, _20844_, _20845_, _20846_, _20847_, _20848_, _20849_, _20850_, _20851_, _20852_, _20853_, _20854_, _20855_, _20856_, _20857_, _20858_, _20859_, _20860_, _20861_, _20862_, _20863_, _20864_, _20865_, _20866_, _20867_, _20868_, _20869_, _20870_, _20871_, _20872_, _20873_, _20874_, _20875_, _20876_, _20877_, _20878_, _20879_, _20880_, _20881_, _20882_, _20883_, _20884_, _20885_, _20886_, _20887_, _20888_, _20889_, _20890_, _20891_, _20892_, _20893_, _20894_, _20895_, _20896_, _20897_, _20898_, _20899_, _20900_, _20901_, _20902_, _20903_, _20904_, _20905_, _20906_, _20907_, _20908_, _20909_, _20910_, _20911_, _20912_, _20913_, _20914_, _20915_, _20916_, _20917_, _20918_, _20919_, _20920_, _20921_, _20922_, _20923_, _20924_, _20925_, _20926_, _20927_, _20928_, _20929_, _20930_, _20931_, _20932_, _20933_, _20934_, _20935_, _20936_, _20937_, _20938_, _20939_, _20940_, _20941_, _20942_, _20943_, _20944_, _20945_, _20946_, _20947_, _20948_, _20949_, _20950_, _20951_, _20952_, _20953_, _20954_, _20955_, _20956_, _20957_, _20958_, _20959_, _20960_, _20961_, _20962_, _20963_, _20964_, _20965_, _20966_, _20967_, _20968_, _20969_, _20970_, _20971_, _20972_, _20973_, _20974_, _20975_, _20976_, _20977_, _20978_, _20979_, _20980_, _20981_, _20982_, _20983_, _20984_, _20985_, _20986_, _20987_, _20988_, _20989_, _20990_, _20991_, _20992_, _20993_, _20994_, _20995_, _20996_, _20997_, _20998_, _20999_, _21000_, _21001_, _21002_, _21003_, _21004_, _21005_, _21006_, _21007_, _21008_, _21009_, _21010_, _21011_, _21012_, _21013_, _21014_, _21015_, _21016_, _21017_, _21018_, _21019_, _21020_, _21021_, _21022_, _21023_, _21024_, _21025_, _21026_, _21027_, _21028_, _21029_, _21030_, _21031_, _21032_, _21033_, _21034_, _21035_, _21036_, _21037_, _21038_, _21039_, _21040_, _21041_, _21042_, _21043_, _21044_, _21045_, _21046_, _21047_, _21048_, _21049_, _21050_, _21051_, _21052_, _21053_, _21054_, _21055_, _21056_, _21057_, _21058_, _21059_, _21060_, _21061_, _21062_, _21063_, _21064_, _21065_, _21066_, _21067_, _21068_, _21069_, _21070_, _21071_, _21072_, _21073_, _21074_, _21075_, _21076_, _21077_, _21078_, _21079_, _21080_, _21081_, _21082_, _21083_, _21084_, _21085_, _21086_, _21087_, _21088_, _21089_, _21090_, _21091_, _21092_, _21093_, _21094_, _21095_, _21096_, _21097_, _21098_, _21099_, _21100_, _21101_, _21102_, _21103_, _21104_, _21105_, _21106_, _21107_, _21108_, _21109_, _21110_, _21111_, _21112_, _21113_, _21114_, _21115_, _21116_, _21117_, _21118_, _21119_, _21120_, _21121_, _21122_, _21123_, _21124_, _21125_, _21126_, _21127_, _21128_, _21129_, _21130_, _21131_, _21132_, _21133_, _21134_, _21135_, _21136_, _21137_, _21138_, _21139_, _21140_, _21141_, _21142_, _21143_, _21144_, _21145_, _21146_, _21147_, _21148_, _21149_, _21150_, _21151_, _21152_, _21153_, _21154_, _21155_, _21156_, _21157_, _21158_, _21159_, _21160_, _21161_, _21162_, _21163_, _21164_, _21165_, _21166_, _21167_, _21168_, _21169_, _21170_, _21171_, _21172_, _21173_, _21174_, _21175_, _21176_, _21177_, _21178_, _21179_, _21180_, _21181_, _21182_, _21183_, _21184_, _21185_, _21186_, _21187_, _21188_, _21189_, _21190_, _21191_, _21192_, _21193_, _21194_, _21195_, _21196_, _21197_, _21198_, _21199_, _21200_, _21201_, _21202_, _21203_, _21204_, _21205_, _21206_, _21207_, _21208_, _21209_, _21210_, _21211_, _21212_, _21213_, _21214_, _21215_, _21216_, _21217_, _21218_, _21219_, _21220_, _21221_, _21222_, _21223_, _21224_, _21225_, _21226_, _21227_, _21228_, _21229_, _21230_, _21231_, _21232_, _21233_, _21234_, _21235_, _21236_, _21237_, _21238_, _21239_, _21240_, _21241_, _21242_, _21243_, _21244_, _21245_, _21246_, _21247_, _21248_, _21249_, _21250_, _21251_, _21252_, _21253_, _21254_, _21255_, _21256_, _21257_, _21258_, _21259_, _21260_, _21261_, _21262_, _21263_, _21264_, _21265_, _21266_, _21267_, _21268_, _21269_, _21270_, _21271_, _21272_, _21273_, _21274_, _21275_, _21276_, _21277_, _21278_, _21279_, _21280_, _21281_, _21282_, _21283_, _21284_, _21285_, _21286_, _21287_, _21288_, _21289_, _21290_, _21291_, _21292_, _21293_, _21294_, _21295_, _21296_, _21297_, _21298_, _21299_, _21300_, _21301_, _21302_, _21303_, _21304_, _21305_, _21306_, _21307_, _21308_, _21309_, _21310_, _21311_, _21312_, _21313_, _21314_, _21315_, _21316_, _21317_, _21318_, _21319_, _21320_, _21321_, _21322_, _21323_, _21324_, _21325_, _21326_, _21327_, _21328_, _21329_, _21330_, _21331_, _21332_, _21333_, _21334_, _21335_, _21336_, _21337_, _21338_, _21339_, _21340_, _21341_, _21342_, _21343_, _21344_, _21345_, _21346_, _21347_, _21348_, _21349_, _21350_, _21351_, _21352_, _21353_, _21354_, _21355_, _21356_, _21357_, _21358_, _21359_, _21360_, _21361_, _21362_, _21363_, _21364_, _21365_, _21366_, _21367_, _21368_, _21369_, _21370_, _21371_, _21372_, _21373_, _21374_, _21375_, _21376_, _21377_, _21378_, _21379_, _21380_, _21381_, _21382_, _21383_, _21384_, _21385_, _21386_, _21387_, _21388_, _21389_, _21390_, _21391_, _21392_, _21393_, _21394_, _21395_, _21396_, _21397_, _21398_, _21399_, _21400_, _21401_, _21402_, _21403_, _21404_, _21405_, _21406_, _21407_, _21408_, _21409_, _21410_, _21411_, _21412_, _21413_, _21414_, _21415_, _21416_, _21417_, _21418_, _21419_, _21420_, _21421_, _21422_, _21423_, _21424_, _21425_, _21426_, _21427_, _21428_, _21429_, _21430_, _21431_, _21432_, _21433_, _21434_, _21435_, _21436_, _21437_, _21438_, _21439_, _21440_, _21441_, _21442_, _21443_, _21444_, _21445_, _21446_, _21447_, _21448_, _21449_, _21450_, _21451_, _21452_, _21453_, _21454_, _21455_, _21456_, _21457_, _21458_, _21459_, _21460_, _21461_, _21462_, _21463_, _21464_, _21465_, _21466_, _21467_, _21468_, _21469_, _21470_, _21471_, _21472_, _21473_, _21474_, _21475_, _21476_, _21477_, _21478_, _21479_, _21480_, _21481_, _21482_, _21483_, _21484_, _21485_, _21486_, _21487_, _21488_, _21489_, _21490_, _21491_, _21492_, _21493_, _21494_, _21495_, _21496_, _21497_, _21498_, _21499_, _21500_, _21501_, _21502_, _21503_, _21504_, _21505_, _21506_, _21507_, _21508_, _21509_, _21510_, _21511_, _21512_, _21513_, _21514_, _21515_, _21516_, _21517_, _21518_, _21519_, _21520_, _21521_, _21522_, _21523_, _21524_, _21525_, _21526_, _21527_, _21528_, _21529_, _21530_, _21531_, _21532_, _21533_, _21534_, _21535_, _21536_, _21537_, _21538_, _21539_, _21540_, _21541_, _21542_, _21543_, _21544_, _21545_, _21546_, _21547_, _21548_, _21549_, _21550_, _21551_, _21552_, _21553_, _21554_, _21555_, _21556_, _21557_, _21558_, _21559_, _21560_, _21561_, _21562_, _21563_, _21564_, _21565_, _21566_, _21567_, _21568_, _21569_, _21570_, _21571_, _21572_, _21573_, _21574_, _21575_, _21576_, _21577_, _21578_, _21579_, _21580_, _21581_, _21582_, _21583_, _21584_, _21585_, _21586_, _21587_, _21588_, _21589_, _21590_, _21591_, _21592_, _21593_, _21594_, _21595_, _21596_, _21597_, _21598_, _21599_, _21600_, _21601_, _21602_, _21603_, _21604_, _21605_, _21606_, _21607_, _21608_, _21609_, _21610_, _21611_, _21612_, _21613_, _21614_, _21615_, _21616_, _21617_, _21618_, _21619_, _21620_, _21621_, _21622_, _21623_, _21624_, _21625_, _21626_, _21627_, _21628_, _21629_, _21630_, _21631_, _21632_, _21633_, _21634_, _21635_, _21636_, _21637_, _21638_, _21639_, _21640_, _21641_, _21642_, _21643_, _21644_, _21645_, _21646_, _21647_, _21648_, _21649_, _21650_, _21651_, _21652_, _21653_, _21654_, _21655_, _21656_, _21657_, _21658_, _21659_, _21660_, _21661_, _21662_, _21663_, _21664_, _21665_, _21666_, _21667_, _21668_, _21669_, _21670_, _21671_, _21672_, _21673_, _21674_, _21675_, _21676_, _21677_, _21678_, _21679_, _21680_, _21681_, _21682_, _21683_, _21684_, _21685_, _21686_, _21687_, _21688_, _21689_, _21690_, _21691_, _21692_, _21693_, _21694_, _21695_, _21696_, _21697_, _21698_, _21699_, _21700_, _21701_, _21702_, _21703_, _21704_, _21705_, _21706_, _21707_, _21708_, _21709_, _21710_, _21711_, _21712_, _21713_, _21714_, _21715_, _21716_, _21717_, _21718_, _21719_, _21720_, _21721_, _21722_, _21723_, _21724_, _21725_, _21726_, _21727_, _21728_, _21729_, _21730_, _21731_, _21732_, _21733_, _21734_, _21735_, _21736_, _21737_, _21738_, _21739_, _21740_, _21741_, _21742_, _21743_, _21744_, _21745_, _21746_, _21747_, _21748_, _21749_, _21750_, _21751_, _21752_, _21753_, _21754_, _21755_, _21756_, _21757_, _21758_, _21759_, _21760_, _21761_, _21762_, _21763_, _21764_, _21765_, _21766_, _21767_, _21768_, _21769_, _21770_, _21771_, _21772_, _21773_, _21774_, _21775_, _21776_, _21777_, _21778_, _21779_, _21780_, _21781_, _21782_, _21783_, _21784_, _21785_, _21786_, _21787_, _21788_, _21789_, _21790_, _21791_, _21792_, _21793_, _21794_, _21795_, _21796_, _21797_, _21798_, _21799_, _21800_, _21801_, _21802_, _21803_, _21804_, _21805_, _21806_, _21807_, _21808_, _21809_, _21810_, _21811_, _21812_, _21813_, _21814_, _21815_, _21816_, _21817_, _21818_, _21819_, _21820_, _21821_, _21822_, _21823_, _21824_, _21825_, _21826_, _21827_, _21828_, _21829_, _21830_, _21831_, _21832_, _21833_, _21834_, _21835_, _21836_, _21837_, _21838_, _21839_, _21840_, _21841_, _21842_, _21843_, _21844_, _21845_, _21846_, _21847_, _21848_, _21849_, _21850_, _21851_, _21852_, _21853_, _21854_, _21855_, _21856_, _21857_, _21858_, _21859_, _21860_, _21861_, _21862_, _21863_, _21864_, _21865_, _21866_, _21867_, _21868_, _21869_, _21870_, _21871_, _21872_, _21873_, _21874_, _21875_, _21876_, _21877_, _21878_, _21879_, _21880_, _21881_, _21882_, _21883_, _21884_, _21885_, _21886_, _21887_, _21888_, _21889_, _21890_, _21891_, _21892_, _21893_, _21894_, _21895_, _21896_, _21897_, _21898_, _21899_, _21900_, _21901_, _21902_, _21903_, _21904_, _21905_, _21906_, _21907_, _21908_, _21909_, _21910_, _21911_, _21912_, _21913_, _21914_, _21915_, _21916_, _21917_, _21918_, _21919_, _21920_, _21921_, _21922_, _21923_, _21924_, _21925_, _21926_, _21927_, _21928_, _21929_, _21930_, _21931_, _21932_, _21933_, _21934_, _21935_, _21936_, _21937_, _21938_, _21939_, _21940_, _21941_, _21942_, _21943_, _21944_, _21945_, _21946_, _21947_, _21948_, _21949_, _21950_, _21951_, _21952_, _21953_, _21954_, _21955_, _21956_, _21957_, _21958_, _21959_, _21960_, _21961_, _21962_, _21963_, _21964_, _21965_, _21966_, _21967_, _21968_, _21969_, _21970_, _21971_, _21972_, _21973_, _21974_, _21975_, _21976_, _21977_, _21978_, _21979_, _21980_, _21981_, _21982_, _21983_, _21984_, _21985_, _21986_, _21987_, _21988_, _21989_, _21990_, _21991_, _21992_, _21993_, _21994_, _21995_, _21996_, _21997_, _21998_, _21999_, _22000_, _22001_, _22002_, _22003_, _22004_, _22005_, _22006_, _22007_, _22008_, _22009_, _22010_, _22011_, _22012_, _22013_, _22014_, _22015_, _22016_, _22017_, _22018_, _22019_, _22020_, _22021_, _22022_, _22023_, _22024_, _22025_, _22026_, _22027_, _22028_, _22029_, _22030_, _22031_, _22032_, _22033_, _22034_, _22035_, _22036_, _22037_, _22038_, _22039_, _22040_, _22041_, _22042_, _22043_, _22044_, _22045_, _22046_, _22047_, _22048_, _22049_, _22050_, _22051_, _22052_, _22053_, _22054_, _22055_, _22056_, _22057_, _22058_, _22059_, _22060_, _22061_, _22062_, _22063_, _22064_, _22065_, _22066_, _22067_, _22068_, _22069_, _22070_, _22071_, _22072_, _22073_, _22074_, _22075_, _22076_, _22077_, _22078_, _22079_, _22080_, _22081_, _22082_, _22083_, _22084_, _22085_, _22086_, _22087_, _22088_, _22089_, _22090_, _22091_, _22092_, _22093_, _22094_, _22095_, _22096_, _22097_, _22098_, _22099_, _22100_, _22101_, _22102_, _22103_, _22104_, _22105_, _22106_, _22107_, _22108_, _22109_, _22110_, _22111_, _22112_, _22113_, _22114_, _22115_, _22116_, _22117_, _22118_, _22119_, _22120_, _22121_, _22122_, _22123_, _22124_, _22125_, _22126_, _22127_, _22128_, _22129_, _22130_, _22131_, _22132_, _22133_, _22134_, _22135_, _22136_, _22137_, _22138_, _22139_, _22140_, _22141_, _22142_, _22143_, _22144_, _22145_, _22146_, _22147_, _22148_, _22149_, _22150_, _22151_, _22152_, _22153_, _22154_, _22155_, _22156_, _22157_, _22158_, _22159_, _22160_, _22161_, _22162_, _22163_, _22164_, _22165_, _22166_, _22167_, _22168_, _22169_, _22170_, _22171_, _22172_, _22173_, _22174_, _22175_, _22176_, _22177_, _22178_, _22179_, _22180_, _22181_, _22182_, _22183_, _22184_, _22185_, _22186_, _22187_, _22188_, _22189_, _22190_, _22191_, _22192_, _22193_, _22194_, _22195_, _22196_, _22197_, _22198_, _22199_, _22200_, _22201_, _22202_, _22203_, _22204_, _22205_, _22206_, _22207_, _22208_, _22209_, _22210_, _22211_, _22212_, _22213_, _22214_, _22215_, _22216_, _22217_, _22218_, _22219_, _22220_, _22221_, _22222_, _22223_, _22224_, _22225_, _22226_, _22227_, _22228_, _22229_, _22230_, _22231_, _22232_, _22233_, _22234_, _22235_, _22236_, _22237_, _22238_, _22239_, _22240_, _22241_, _22242_, _22243_, _22244_, _22245_, _22246_, _22247_, _22248_, _22249_, _22250_, _22251_, _22252_, _22253_, _22254_, _22255_, _22256_, _22257_, _22258_, _22259_, _22260_, _22261_, _22262_, _22263_, _22264_, _22265_, _22266_, _22267_, _22268_, _22269_, _22270_, _22271_, _22272_, _22273_, _22274_, _22275_, _22276_, _22277_, _22278_, _22279_, _22280_, _22281_, _22282_, _22283_, _22284_, _22285_, _22286_, _22287_, _22288_, _22289_, _22290_, _22291_, _22292_, _22293_, _22294_, _22295_, _22296_, _22297_, _22298_, _22299_, _22300_, _22301_, _22302_, _22303_, _22304_, _22305_, _22306_, _22307_, _22308_, _22309_, _22310_, _22311_, _22312_, _22313_, _22314_, _22315_, _22316_, _22317_, _22318_, _22319_, _22320_, _22321_, _22322_, _22323_, _22324_, _22325_, _22326_, _22327_, _22328_, _22329_, _22330_, _22331_, _22332_, _22333_, _22334_, _22335_, _22336_, _22337_, _22338_, _22339_, _22340_, _22341_, _22342_, _22343_, _22344_, _22345_, _22346_, _22347_, _22348_, _22349_, _22350_, _22351_, _22352_, _22353_, _22354_, _22355_, _22356_, _22357_, _22358_, _22359_, _22360_, _22361_, _22362_, _22363_, _22364_, _22365_, _22366_, _22367_, _22368_, _22369_, _22370_, _22371_, _22372_, _22373_, _22374_, _22375_, _22376_, _22377_, _22378_, _22379_, _22380_, _22381_, _22382_, _22383_, _22384_, _22385_, _22386_, _22387_, _22388_, _22389_, _22390_, _22391_, _22392_, _22393_, _22394_, _22395_, _22396_, _22397_, _22398_, _22399_, _22400_, _22401_, _22402_, _22403_, _22404_, _22405_, _22406_, _22407_, _22408_, _22409_, _22410_, _22411_, _22412_, _22413_, _22414_, _22415_, _22416_, _22417_, _22418_, _22419_, _22420_, _22421_, _22422_, _22423_, _22424_, _22425_, _22426_, _22427_, _22428_, _22429_, _22430_, _22431_, _22432_, _22433_, _22434_, _22435_, _22436_, _22437_, _22438_, _22439_, _22440_, _22441_, _22442_, _22443_, _22444_, _22445_, _22446_, _22447_, _22448_, _22449_, _22450_, _22451_, _22452_, _22453_, _22454_, _22455_, _22456_, _22457_, _22458_, _22459_, _22460_, _22461_, _22462_, _22463_, _22464_, _22465_, _22466_, _22467_, _22468_, _22469_, _22470_, _22471_, _22472_, _22473_, _22474_, _22475_, _22476_, _22477_, _22478_, _22479_, _22480_, _22481_, _22482_, _22483_, _22484_, _22485_, _22486_, _22487_, _22488_, _22489_, _22490_, _22491_, _22492_, _22493_, _22494_, _22495_, _22496_, _22497_, _22498_, _22499_, _22500_, _22501_, _22502_, _22503_, _22504_, _22505_, _22506_, _22507_, _22508_, _22509_, _22510_, _22511_, _22512_, _22513_, _22514_, _22515_, _22516_, _22517_, _22518_, _22519_, _22520_, _22521_, _22522_, _22523_, _22524_, _22525_, _22526_, _22527_, _22528_, _22529_, _22530_, _22531_, _22532_, _22533_, _22534_, _22535_, _22536_, _22537_, _22538_, _22539_, _22540_, _22541_, _22542_, _22543_, _22544_, _22545_, _22546_, _22547_, _22548_, _22549_, _22550_, _22551_, _22552_, _22553_, _22554_, _22555_, _22556_, _22557_, _22558_, _22559_, _22560_, _22561_, _22562_, _22563_, _22564_, _22565_, _22566_, _22567_, _22568_, _22569_, _22570_, _22571_, _22572_, _22573_, _22574_, _22575_, _22576_, _22577_, _22578_, _22579_, _22580_, _22581_, _22582_, _22583_, _22584_, _22585_, _22586_, _22587_, _22588_, _22589_, _22590_, _22591_, _22592_, _22593_, _22594_, _22595_, _22596_, _22597_, _22598_, _22599_, _22600_, _22601_, _22602_, _22603_, _22604_, _22605_, _22606_, _22607_, _22608_, _22609_, _22610_, _22611_, _22612_, _22613_, _22614_, _22615_, _22616_, _22617_, _22618_, _22619_, _22620_, _22621_, _22622_, _22623_, _22624_, _22625_, _22626_, _22627_, _22628_, _22629_, _22630_, _22631_, _22632_, _22633_, _22634_, _22635_, _22636_, _22637_, _22638_, _22639_, _22640_, _22641_, _22642_, _22643_, _22644_, _22645_, _22646_, _22647_, _22648_, _22649_, _22650_, _22651_, _22652_, _22653_, _22654_, _22655_, _22656_, _22657_, _22658_, _22659_, _22660_, _22661_, _22662_, _22663_, _22664_, _22665_, _22666_, _22667_, _22668_, _22669_, _22670_, _22671_, _22672_, _22673_, _22674_, _22675_, _22676_, _22677_, _22678_, _22679_, _22680_, _22681_, _22682_, _22683_, _22684_, _22685_, _22686_, _22687_, _22688_, _22689_, _22690_, _22691_, _22692_, _22693_, _22694_, _22695_, _22696_, _22697_, _22698_, _22699_, _22700_, _22701_, _22702_, _22703_, _22704_, _22705_, _22706_, _22707_, _22708_, _22709_, _22710_, _22711_, _22712_, _22713_, _22714_, _22715_, _22716_, _22717_, _22718_, _22719_, _22720_, _22721_, _22722_, _22723_, _22724_, _22725_, _22726_, _22727_, _22728_, _22729_, _22730_, _22731_, _22732_, _22733_, _22734_, _22735_, _22736_, _22737_, _22738_, _22739_, _22740_, _22741_, _22742_, _22743_, _22744_, _22745_, _22746_, _22747_, _22748_, _22749_, _22750_, _22751_, _22752_, _22753_, _22754_, _22755_, _22756_, _22757_, _22758_, _22759_, _22760_, _22761_, _22762_, _22763_, _22764_, _22765_, _22766_, _22767_, _22768_, _22769_, _22770_, _22771_, _22772_, _22773_, _22774_, _22775_, _22776_, _22777_, _22778_, _22779_, _22780_, _22781_, _22782_, _22783_, _22784_, _22785_, _22786_, _22787_, _22788_, _22789_, _22790_, _22791_, _22792_, _22793_, _22794_, _22795_, _22796_, _22797_, _22798_, _22799_, _22800_, _22801_, _22802_, _22803_, _22804_, _22805_, _22806_, _22807_, _22808_, _22809_, _22810_, _22811_, _22812_, _22813_, _22814_, _22815_, _22816_, _22817_, _22818_, _22819_, _22820_, _22821_, _22822_, _22823_, _22824_, _22825_, _22826_, _22827_, _22828_, _22829_, _22830_, _22831_, _22832_, _22833_, _22834_, _22835_, _22836_, _22837_, _22838_, _22839_, _22840_, _22841_, _22842_, _22843_, _22844_, _22845_, _22846_, _22847_, _22848_, _22849_, _22850_, _22851_, _22852_, _22853_, _22854_, _22855_, _22856_, _22857_, _22858_, _22859_, _22860_, _22861_, _22862_, _22863_, _22864_, _22865_, _22866_, _22867_, _22868_, _22869_, _22870_, _22871_, _22872_, _22873_, _22874_, _22875_, _22876_, _22877_, _22878_, _22879_, _22880_, _22881_, _22882_, _22883_, _22884_, _22885_, _22886_, _22887_, _22888_, _22889_, _22890_, _22891_, _22892_, _22893_, _22894_, _22895_, _22896_, _22897_, _22898_, _22899_, _22900_, _22901_, _22902_, _22903_, _22904_, _22905_, _22906_, _22907_, _22908_, _22909_, _22910_, _22911_, _22912_, _22913_, _22914_, _22915_, _22916_, _22917_, _22918_, _22919_, _22920_, _22921_, _22922_, _22923_, _22924_, _22925_, _22926_, _22927_, _22928_, _22929_, _22930_, _22931_, _22932_, _22933_, _22934_, _22935_, _22936_, _22937_, _22938_, _22939_, _22940_, _22941_, _22942_, _22943_, _22944_, _22945_, _22946_, _22947_, _22948_, _22949_, _22950_, _22951_, _22952_, _22953_, _22954_, _22955_, _22956_, _22957_, _22958_, _22959_, _22960_, _22961_, _22962_, _22963_, _22964_, _22965_, _22966_, _22967_, _22968_, _22969_, _22970_, _22971_, _22972_, _22973_, _22974_, _22975_, _22976_, _22977_, _22978_, _22979_, _22980_, _22981_, _22982_, _22983_, _22984_, _22985_, _22986_, _22987_, _22988_, _22989_, _22990_, _22991_, _22992_, _22993_, _22994_, _22995_, _22996_, _22997_, _22998_, _22999_, _23000_, _23001_, _23002_, _23003_, _23004_, _23005_, _23006_, _23007_, _23008_, _23009_, _23010_, _23011_, _23012_, _23013_, _23014_, _23015_, _23016_, _23017_, _23018_, _23019_, _23020_, _23021_, _23022_, _23023_, _23024_, _23025_, _23026_, _23027_, _23028_, _23029_, _23030_, _23031_, _23032_, _23033_, _23034_, _23035_, _23036_, _23037_, _23038_, _23039_, _23040_, _23041_, _23042_, _23043_, _23044_, _23045_, _23046_, _23047_, _23048_, _23049_, _23050_, _23051_, _23052_, _23053_, _23054_, _23055_, _23056_, _23057_, _23058_, _23059_, _23060_, _23061_, _23062_, _23063_, _23064_, _23065_, _23066_, _23067_, _23068_, _23069_, _23070_, _23071_, _23072_, _23073_, _23074_, _23075_, _23076_, _23077_, _23078_, _23079_, _23080_, _23081_, _23082_, _23083_, _23084_, _23085_, _23086_, _23087_, _23088_, _23089_, _23090_, _23091_, _23092_, _23093_, _23094_, _23095_, _23096_, _23097_, _23098_, _23099_, _23100_, _23101_, _23102_, _23103_, _23104_, _23105_, _23106_, _23107_, _23108_, _23109_, _23110_, _23111_, _23112_, _23113_, _23114_, _23115_, _23116_, _23117_, _23118_, _23119_, _23120_, _23121_, _23122_, _23123_, _23124_, _23125_, _23126_, _23127_, _23128_, _23129_, _23130_, _23131_, _23132_, _23133_, _23134_, _23135_, _23136_, _23137_, _23138_, _23139_, _23140_, _23141_, _23142_, _23143_, _23144_, _23145_, _23146_, _23147_, _23148_, _23149_, _23150_, _23151_, _23152_, _23153_, _23154_, _23155_, _23156_, _23157_, _23158_, _23159_, _23160_, _23161_, _23162_, _23163_, _23164_, _23165_, _23166_, _23167_, _23168_, _23169_, _23170_, _23171_, _23172_, _23173_, _23174_, _23175_, _23176_, _23177_, _23178_, _23179_, _23180_, _23181_, _23182_, _23183_, _23184_, _23185_, _23186_, _23187_, _23188_, _23189_, _23190_, _23191_, _23192_, _23193_, _23194_, _23195_, _23196_, _23197_, _23198_, _23199_, _23200_, _23201_, _23202_, _23203_, _23204_, _23205_, _23206_, _23207_, _23208_, _23209_, _23210_, _23211_, _23212_, _23213_, _23214_, _23215_, _23216_, _23217_, _23218_, _23219_, _23220_, _23221_, _23222_, _23223_, _23224_, _23225_, _23226_, _23227_, _23228_, _23229_, _23230_, _23231_, _23232_, _23233_, _23234_, _23235_, _23236_, _23237_, _23238_, _23239_, _23240_, _23241_, _23242_, _23243_, _23244_, _23245_, _23246_, _23247_, _23248_, _23249_, _23250_, _23251_, _23252_, _23253_, _23254_, _23255_, _23256_, _23257_, _23258_, _23259_, _23260_, _23261_, _23262_, _23263_, _23264_, _23265_, _23266_, _23267_, _23268_, _23269_, _23270_, _23271_, _23272_, _23273_, _23274_, _23275_, _23276_, _23277_, _23278_, _23279_, _23280_, _23281_, _23282_, _23283_, _23284_, _23285_, _23286_, _23287_, _23288_, _23289_, _23290_, _23291_, _23292_, _23293_, _23294_, _23295_, _23296_, _23297_, _23298_, _23299_, _23300_, _23301_, _23302_, _23303_, _23304_, _23305_, _23306_, _23307_, _23308_, _23309_, _23310_, _23311_, _23312_, _23313_, _23314_, _23315_, _23316_, _23317_, _23318_, _23319_, _23320_, _23321_, _23322_, _23323_, _23324_, _23325_, _23326_, _23327_, _23328_, _23329_, _23330_, _23331_, _23332_, _23333_, _23334_, _23335_, _23336_, _23337_, _23338_, _23339_, _23340_, _23341_, _23342_, _23343_, _23344_, _23345_, _23346_, _23347_, _23348_, _23349_, _23350_, _23351_, _23352_, _23353_, _23354_, _23355_, _23356_, _23357_, _23358_, _23359_, _23360_, _23361_, _23362_, _23363_, _23364_, _23365_, _23366_, _23367_, _23368_, _23369_, _23370_, _23371_, _23372_, _23373_, _23374_, _23375_, _23376_, _23377_, _23378_, _23379_, _23380_, _23381_, _23382_, _23383_, _23384_, _23385_, _23386_, _23387_, _23388_, _23389_, _23390_, _23391_, _23392_, _23393_, _23394_, _23395_, _23396_, _23397_, _23398_, _23399_, _23400_, _23401_, _23402_, _23403_, _23404_, _23405_, _23406_, _23407_, _23408_, _23409_, _23410_, _23411_, _23412_, _23413_, _23414_, _23415_, _23416_, _23417_, _23418_, _23419_, _23420_, _23421_, _23422_, _23423_, _23424_, _23425_, _23426_, _23427_, _23428_, _23429_, _23430_, _23431_, _23432_, _23433_, _23434_, _23435_, _23436_, _23437_, _23438_, _23439_, _23440_, _23441_, _23442_, _23443_, _23444_, _23445_, _23446_, _23447_, _23448_, _23449_, _23450_, _23451_, _23452_, _23453_, _23454_, _23455_, _23456_, _23457_, _23458_, _23459_, _23460_, _23461_, _23462_, _23463_, _23464_, _23465_, _23466_, _23467_, _23468_, _23469_, _23470_, _23471_, _23472_, _23473_, _23474_, _23475_, _23476_, _23477_, _23478_, _23479_, _23480_, _23481_, _23482_, _23483_, _23484_, _23485_, _23486_, _23487_, _23488_, _23489_, _23490_, _23491_, _23492_, _23493_, _23494_, _23495_, _23496_, _23497_, _23498_, _23499_, _23500_, _23501_, _23502_, _23503_, _23504_, _23505_, _23506_, _23507_, _23508_, _23509_, _23510_, _23511_, _23512_, _23513_, _23514_, _23515_, _23516_, _23517_, _23518_, _23519_, _23520_, _23521_, _23522_, _23523_, _23524_, _23525_, _23526_, _23527_, _23528_, _23529_, _23530_, _23531_, _23532_, _23533_, _23534_, _23535_, _23536_, _23537_, _23538_, _23539_, _23540_, _23541_, _23542_, _23543_, _23544_, _23545_, _23546_, _23547_, _23548_, _23549_, _23550_, _23551_, _23552_, _23553_, _23554_, _23555_, _23556_, _23557_, _23558_, _23559_, _23560_, _23561_, _23562_, _23563_, _23564_, _23565_, _23566_, _23567_, _23568_, _23569_, _23570_, _23571_, _23572_, _23573_, _23574_, _23575_, _23576_, _23577_, _23578_, _23579_, _23580_, _23581_, _23582_, _23583_, _23584_, _23585_, _23586_, _23587_, _23588_, _23589_, _23590_, _23591_, _23592_, _23593_, _23594_, _23595_, _23596_, _23597_, _23598_, _23599_, _23600_, _23601_, _23602_, _23603_, _23604_, _23605_, _23606_, _23607_, _23608_, _23609_, _23610_, _23611_, _23612_, _23613_, _23614_, _23615_, _23616_, _23617_, _23618_, _23619_, _23620_, _23621_, _23622_, _23623_, _23624_, _23625_, _23626_, _23627_, _23628_, _23629_, _23630_, _23631_, _23632_, _23633_, _23634_, _23635_, _23636_, _23637_, _23638_, _23639_, _23640_, _23641_, _23642_, _23643_, _23644_, _23645_, _23646_, _23647_, _23648_, _23649_, _23650_, _23651_, _23652_, _23653_, _23654_, _23655_, _23656_, _23657_, _23658_, _23659_, _23660_, _23661_, _23662_, _23663_, _23664_, _23665_, _23666_, _23667_, _23668_, _23669_, _23670_, _23671_, _23672_, _23673_, _23674_, _23675_, _23676_, _23677_, _23678_, _23679_, _23680_, _23681_, _23682_, _23683_, _23684_, _23685_, _23686_, _23687_, _23688_, _23689_, _23690_, _23691_, _23692_, _23693_, _23694_, _23695_, _23696_, _23697_, _23698_, _23699_, _23700_, _23701_, _23702_, _23703_, _23704_, _23705_, _23706_, _23707_, _23708_, _23709_, _23710_, _23711_, _23712_, _23713_, _23714_, _23715_, _23716_, _23717_, _23718_, _23719_, _23720_, _23721_, _23722_, _23723_, _23724_, _23725_, _23726_, _23727_, _23728_, _23729_, _23730_, _23731_, _23732_, _23733_, _23734_, _23735_, _23736_, _23737_, _23738_, _23739_, _23740_, _23741_, _23742_, _23743_, _23744_, _23745_, _23746_, _23747_, _23748_, _23749_, _23750_, _23751_, _23752_, _23753_, _23754_, _23755_, _23756_, _23757_, _23758_, _23759_, _23760_, _23761_, _23762_, _23763_, _23764_, _23765_, _23766_, _23767_, _23768_, _23769_, _23770_, _23771_, _23772_, _23773_, _23774_, _23775_, _23776_, _23777_, _23778_, _23779_, _23780_, _23781_, _23782_, _23783_, _23784_, _23785_, _23786_, _23787_, _23788_, _23789_, _23790_, _23791_, _23792_, _23793_, _23794_, _23795_, _23796_, _23797_, _23798_, _23799_, _23800_, _23801_, _23802_, _23803_, _23804_, _23805_, _23806_, _23807_, _23808_, _23809_, _23810_, _23811_, _23812_, _23813_, _23814_, _23815_, _23816_, _23817_, _23818_, _23819_, _23820_, _23821_, _23822_, _23823_, _23824_, _23825_, _23826_, _23827_, _23828_, _23829_, _23830_, _23831_, _23832_, _23833_, _23834_, _23835_, _23836_, _23837_, _23838_, _23839_, _23840_, _23841_, _23842_, _23843_, _23844_, _23845_, _23846_, _23847_, _23848_, _23849_, _23850_, _23851_, _23852_, _23853_, _23854_, _23855_, _23856_, _23857_, _23858_, _23859_, _23860_, _23861_, _23862_, _23863_, _23864_, _23865_, _23866_, _23867_, _23868_, _23869_, _23870_, _23871_, _23872_, _23873_, _23874_, _23875_, _23876_, _23877_, _23878_, _23879_, _23880_, _23881_, _23882_, _23883_, _23884_, _23885_, _23886_, _23887_, _23888_, _23889_, _23890_, _23891_, _23892_, _23893_, _23894_, _23895_, _23896_, _23897_, _23898_, _23899_, _23900_, _23901_, _23902_, _23903_, _23904_, _23905_, _23906_, _23907_, _23908_, _23909_, _23910_, _23911_, _23912_, _23913_, _23914_, _23915_, _23916_, _23917_, _23918_, _23919_, _23920_, _23921_, _23922_, _23923_, _23924_, _23925_, _23926_, _23927_, _23928_, _23929_, _23930_, _23931_, _23932_, _23933_, _23934_, _23935_, _23936_, _23937_, _23938_, _23939_, _23940_, _23941_, _23942_, _23943_, _23944_, _23945_, _23946_, _23947_, _23948_, _23949_, _23950_, _23951_, _23952_, _23953_, _23954_, _23955_, _23956_, _23957_, _23958_, _23959_, _23960_, _23961_, _23962_, _23963_, _23964_, _23965_, _23966_, _23967_, _23968_, _23969_, _23970_, _23971_, _23972_, _23973_, _23974_, _23975_, _23976_, _23977_, _23978_, _23979_, _23980_, _23981_, _23982_, _23983_, _23984_, _23985_, _23986_, _23987_, _23988_, _23989_, _23990_, _23991_, _23992_, _23993_, _23994_, _23995_, _23996_, _23997_, _23998_, _23999_, _24000_, _24001_, _24002_, _24003_, _24004_, _24005_, _24006_, _24007_, _24008_, _24009_, _24010_, _24011_, _24012_, _24013_, _24014_, _24015_, _24016_, _24017_, _24018_, _24019_, _24020_, _24021_, _24022_, _24023_, _24024_, _24025_, _24026_, _24027_, _24028_, _24029_, _24030_, _24031_, _24032_, _24033_, _24034_, _24035_, _24036_, _24037_, _24038_, _24039_, _24040_, _24041_, _24042_, _24043_, _24044_, _24045_, _24046_, _24047_, _24048_, _24049_, _24050_, _24051_, _24052_, _24053_, _24054_, _24055_, _24056_, _24057_, _24058_, _24059_, _24060_, _24061_, _24062_, _24063_, _24064_, _24065_, _24066_, _24067_, _24068_, _24069_, _24070_, _24071_, _24072_, _24073_, _24074_, _24075_, _24076_, _24077_, _24078_, _24079_, _24080_, _24081_, _24082_, _24083_, _24084_, _24085_, _24086_, _24087_, _24088_, _24089_, _24090_, _24091_, _24092_, _24093_, _24094_, _24095_, _24096_, _24097_, _24098_, _24099_, _24100_, _24101_, _24102_, _24103_, _24104_, _24105_, _24106_, _24107_, _24108_, _24109_, _24110_, _24111_, _24112_, _24113_, _24114_, _24115_, _24116_, _24117_, _24118_, _24119_, _24120_, _24121_, _24122_, _24123_, _24124_, _24125_, _24126_, _24127_, _24128_, _24129_, _24130_, _24131_, _24132_, _24133_, _24134_, _24135_, _24136_, _24137_, _24138_, _24139_, _24140_, _24141_, _24142_, _24143_, _24144_, _24145_, _24146_, _24147_, _24148_, _24149_, _24150_, _24151_, _24152_, _24153_, _24154_, _24155_, _24156_, _24157_, _24158_, _24159_, _24160_, _24161_, _24162_, _24163_, _24164_, _24165_, _24166_, _24167_, _24168_, _24169_, _24170_, _24171_, _24172_, _24173_, _24174_, _24175_, _24176_, _24177_, _24178_, _24179_, _24180_, _24181_, _24182_, _24183_, _24184_, _24185_, _24186_, _24187_, _24188_, _24189_, _24190_, _24191_, _24192_, _24193_, _24194_, _24195_, _24196_, _24197_, _24198_, _24199_, _24200_, _24201_, _24202_, _24203_, _24204_, _24205_, _24206_, _24207_, _24208_, _24209_, _24210_, _24211_, _24212_, _24213_, _24214_, _24215_, _24216_, _24217_, _24218_, _24219_, _24220_, _24221_, _24222_, _24223_, _24224_, _24225_, _24226_, _24227_, _24228_, _24229_, _24230_, _24231_, _24232_, _24233_, _24234_, _24235_, _24236_, _24237_, _24238_, _24239_, _24240_, _24241_, _24242_, _24243_, _24244_, _24245_, _24246_, _24247_, _24248_, _24249_, _24250_, _24251_, _24252_, _24253_, _24254_, _24255_, _24256_, _24257_, _24258_, _24259_, _24260_, _24261_, _24262_, _24263_, _24264_, _24265_, _24266_, _24267_, _24268_, _24269_, _24270_, _24271_, _24272_, _24273_, _24274_, _24275_, _24276_, _24277_, _24278_, _24279_, _24280_, _24281_, _24282_, _24283_, _24284_, _24285_, _24286_, _24287_, _24288_, _24289_, _24290_, _24291_, _24292_, _24293_, _24294_, _24295_, _24296_, _24297_, _24298_, _24299_, _24300_, _24301_, _24302_, _24303_, _24304_, _24305_, _24306_, _24307_, _24308_, _24309_, _24310_, _24311_, _24312_, _24313_, _24314_, _24315_, _24316_, _24317_, _24318_, _24319_, _24320_, _24321_, _24322_, _24323_, _24324_, _24325_, _24326_, _24327_, _24328_, _24329_, _24330_, _24331_, _24332_, _24333_, _24334_, _24335_, _24336_, _24337_, _24338_, _24339_, _24340_, _24341_, _24342_, _24343_, _24344_, _24345_, _24346_, _24347_, _24348_, _24349_, _24350_, _24351_, _24352_, _24353_, _24354_, _24355_, _24356_, _24357_, _24358_, _24359_, _24360_, _24361_, _24362_, _24363_, _24364_, _24365_, _24366_, _24367_, _24368_, _24369_, _24370_, _24371_, _24372_, _24373_, _24374_, _24375_, _24376_, _24377_, _24378_, _24379_, _24380_, _24381_, _24382_, _24383_, _24384_, _24385_, _24386_, _24387_, _24388_, _24389_, _24390_, _24391_, _24392_, _24393_, _24394_, _24395_, _24396_, _24397_, _24398_, _24399_, _24400_, _24401_, _24402_, _24403_, _24404_, _24405_, _24406_, _24407_, _24408_, _24409_, _24410_, _24411_, _24412_, _24413_, _24414_, _24415_, _24416_, _24417_, _24418_, _24419_, _24420_, _24421_, _24422_, _24423_, _24424_, _24425_, _24426_, _24427_, _24428_, _24429_, _24430_, _24431_, _24432_, _24433_, _24434_, _24435_, _24436_, _24437_, _24438_, _24439_, _24440_, _24441_, _24442_, _24443_, _24444_, _24445_, _24446_, _24447_, _24448_, _24449_, _24450_, _24451_, _24452_, _24453_, _24454_, _24455_, _24456_, _24457_, _24458_, _24459_, _24460_, _24461_, _24462_, _24463_, _24464_, _24465_, _24466_, _24467_, _24468_, _24469_, _24470_, _24471_, _24472_, _24473_, _24474_, _24475_, _24476_, _24477_, _24478_, _24479_, _24480_, _24481_, _24482_, _24483_, _24484_, _24485_, _24486_, _24487_, _24488_, _24489_, _24490_, _24491_, _24492_, _24493_, _24494_, _24495_, _24496_, _24497_, _24498_, _24499_, _24500_, _24501_, _24502_, _24503_, _24504_, _24505_, _24506_, _24507_, _24508_, _24509_, _24510_, _24511_, _24512_, _24513_, _24514_, _24515_, _24516_, _24517_, _24518_, _24519_, _24520_, _24521_, _24522_, _24523_, _24524_, _24525_, _24526_, _24527_, _24528_, _24529_, _24530_, _24531_, _24532_, _24533_, _24534_, _24535_, _24536_, _24537_, _24538_, _24539_, _24540_, _24541_, _24542_, _24543_, _24544_, _24545_, _24546_, _24547_, _24548_, _24549_, _24550_, _24551_, _24552_, _24553_, _24554_, _24555_, _24556_, _24557_, _24558_, _24559_, _24560_, _24561_, _24562_, _24563_, _24564_, _24565_, _24566_, _24567_, _24568_, _24569_, _24570_, _24571_, _24572_, _24573_, _24574_, _24575_, _24576_, _24577_, _24578_, _24579_, _24580_, _24581_, _24582_, _24583_, _24584_, _24585_, _24586_, _24587_, _24588_, _24589_, _24590_, _24591_, _24592_, _24593_, _24594_, _24595_, _24596_, _24597_, _24598_, _24599_, _24600_, _24601_, _24602_, _24603_, _24604_, _24605_, _24606_, _24607_, _24608_, _24609_, _24610_, _24611_, _24612_, _24613_, _24614_, _24615_, _24616_, _24617_, _24618_, _24619_, _24620_, _24621_, _24622_, _24623_, _24624_, _24625_, _24626_, _24627_, _24628_, _24629_, _24630_, _24631_, _24632_, _24633_, _24634_, _24635_, _24636_, _24637_, _24638_, _24639_, _24640_, _24641_, _24642_, _24643_, _24644_, _24645_, _24646_, _24647_, _24648_, _24649_, _24650_, _24651_, _24652_, _24653_, _24654_, _24655_, _24656_, _24657_, _24658_, _24659_, _24660_, _24661_, _24662_, _24663_, _24664_, _24665_, _24666_, _24667_, _24668_, _24669_, _24670_, _24671_, _24672_, _24673_, _24674_, _24675_, _24676_, _24677_, _24678_, _24679_, _24680_, _24681_, _24682_, _24683_, _24684_, _24685_, _24686_, _24687_, _24688_, _24689_, _24690_, _24691_, _24692_, _24693_, _24694_, _24695_, _24696_, _24697_, _24698_, _24699_, _24700_, _24701_, _24702_, _24703_, _24704_, _24705_, _24706_, _24707_, _24708_, _24709_, _24710_, _24711_, _24712_, _24713_, _24714_, _24715_, _24716_, _24717_, _24718_, _24719_, _24720_, _24721_, _24722_, _24723_, _24724_, _24725_, _24726_, _24727_, _24728_, _24729_, _24730_, _24731_, _24732_, _24733_, _24734_, _24735_, _24736_, _24737_, _24738_, _24739_, _24740_, _24741_, _24742_, _24743_, _24744_, _24745_, _24746_, _24747_, _24748_, _24749_, _24750_, _24751_, _24752_, _24753_, _24754_, _24755_, _24756_, _24757_, _24758_, _24759_, _24760_, _24761_, _24762_, _24763_, _24764_, _24765_, _24766_, _24767_, _24768_, _24769_, _24770_, _24771_, _24772_, _24773_, _24774_, _24775_, _24776_, _24777_, _24778_, _24779_, _24780_, _24781_, _24782_, _24783_, _24784_, _24785_, _24786_, _24787_, _24788_, _24789_, _24790_, _24791_, _24792_, _24793_, _24794_, _24795_, _24796_, _24797_, _24798_, _24799_, _24800_, _24801_, _24802_, _24803_, _24804_, _24805_, _24806_, _24807_, _24808_, _24809_, _24810_, _24811_, _24812_, _24813_, _24814_, _24815_, _24816_, _24817_, _24818_, _24819_, _24820_, _24821_, _24822_, _24823_, _24824_, _24825_, _24826_, _24827_, _24828_, _24829_, _24830_, _24831_, _24832_, _24833_, _24834_, _24835_, _24836_, _24837_, _24838_, _24839_, _24840_, _24841_, _24842_, _24843_, _24844_, _24845_, _24846_, _24847_, _24848_, _24849_, _24850_, _24851_, _24852_, _24853_, _24854_, _24855_, _24856_, _24857_, _24858_, _24859_, _24860_, _24861_, _24862_, _24863_, _24864_, _24865_, _24866_, _24867_, _24868_, _24869_, _24870_, _24871_, _24872_, _24873_, _24874_, _24875_, _24876_, _24877_, _24878_, _24879_, _24880_, _24881_, _24882_, _24883_, _24884_, _24885_, _24886_, _24887_, _24888_, _24889_, _24890_, _24891_, _24892_, _24893_, _24894_, _24895_, _24896_, _24897_, _24898_, _24899_, _24900_, _24901_, _24902_, _24903_, _24904_, _24905_, _24906_, _24907_, _24908_, _24909_, _24910_, _24911_, _24912_, _24913_, _24914_, _24915_, _24916_, _24917_, _24918_, _24919_, _24920_, _24921_, _24922_, _24923_, _24924_, _24925_, _24926_, _24927_, _24928_, _24929_, _24930_, _24931_, _24932_, _24933_, _24934_, _24935_, _24936_, _24937_, _24938_, _24939_, _24940_, _24941_, _24942_, _24943_, _24944_, _24945_, _24946_, _24947_, _24948_, _24949_, _24950_, _24951_, _24952_, _24953_, _24954_, _24955_, _24956_, _24957_, _24958_, _24959_, _24960_, _24961_, _24962_, _24963_, _24964_, _24965_, _24966_, _24967_, _24968_, _24969_, _24970_, _24971_, _24972_, _24973_, _24974_, _24975_, _24976_, _24977_, _24978_, _24979_, _24980_, _24981_, _24982_, _24983_, _24984_, _24985_, _24986_, _24987_, _24988_, _24989_, _24990_, _24991_, _24992_, _24993_, _24994_, _24995_, _24996_, _24997_, _24998_, _24999_, _25000_, _25001_, _25002_, _25003_, _25004_, _25005_, _25006_, _25007_, _25008_, _25009_, _25010_, _25011_, _25012_, _25013_, _25014_, _25015_, _25016_, _25017_, _25018_, _25019_, _25020_, _25021_, _25022_, _25023_, _25024_, _25025_, _25026_, _25027_, _25028_, _25029_, _25030_, _25031_, _25032_, _25033_, _25034_, _25035_, _25036_, _25037_, _25038_, _25039_, _25040_, _25041_, _25042_, _25043_, _25044_, _25045_, _25046_, _25047_, _25048_, _25049_, _25050_, _25051_, _25052_, _25053_, _25054_, _25055_, _25056_, _25057_, _25058_, _25059_, _25060_, _25061_, _25062_, _25063_, _25064_, _25065_, _25066_, _25067_, _25068_, _25069_, _25070_, _25071_, _25072_, _25073_, _25074_, _25075_, _25076_, _25077_, _25078_, _25079_, _25080_, _25081_, _25082_, _25083_, _25084_, _25085_, _25086_, _25087_, _25088_, _25089_, _25090_, _25091_, _25092_, _25093_, _25094_, _25095_, _25096_, _25097_, _25098_, _25099_, _25100_, _25101_, _25102_, _25103_, _25104_, _25105_, _25106_, _25107_, _25108_, _25109_, _25110_, _25111_, _25112_, _25113_, _25114_, _25115_, _25116_, _25117_, _25118_, _25119_, _25120_, _25121_, _25122_, _25123_, _25124_, _25125_, _25126_, _25127_, _25128_, _25129_, _25130_, _25131_, _25132_, _25133_, _25134_, _25135_, _25136_, _25137_, _25138_, _25139_, _25140_, _25141_, _25142_, _25143_, _25144_, _25145_, _25146_, _25147_, _25148_, _25149_, _25150_, _25151_, _25152_, _25153_, _25154_, _25155_, _25156_, _25157_, _25158_, _25159_, _25160_, _25161_, _25162_, _25163_, _25164_, _25165_, _25166_, _25167_, _25168_, _25169_, _25170_, _25171_, _25172_, _25173_, _25174_, _25175_, _25176_, _25177_, _25178_, _25179_, _25180_, _25181_, _25182_, _25183_, _25184_, _25185_, _25186_, _25187_, _25188_, _25189_, _25190_, _25191_, _25192_, _25193_, _25194_, _25195_, _25196_, _25197_, _25198_, _25199_, _25200_, _25201_, _25202_, _25203_, _25204_, _25205_, _25206_, _25207_, _25208_, _25209_, _25210_, _25211_, _25212_, _25213_, _25214_, _25215_, _25216_, _25217_, _25218_, _25219_, _25220_, _25221_, _25222_, _25223_, _25224_, _25225_, _25226_, _25227_, _25228_, _25229_, _25230_, _25231_, _25232_, _25233_, _25234_, _25235_, _25236_, _25237_, _25238_, _25239_, _25240_, _25241_, _25242_, _25243_, _25244_, _25245_, _25246_, _25247_, _25248_, _25249_, _25250_, _25251_, _25252_, _25253_, _25254_, _25255_, _25256_, _25257_, _25258_, _25259_, _25260_, _25261_, _25262_, _25263_, _25264_, _25265_, _25266_, _25267_, _25268_, _25269_, _25270_, _25271_, _25272_, _25273_, _25274_, _25275_, _25276_, _25277_, _25278_, _25279_, _25280_, _25281_, _25282_, _25283_, _25284_, _25285_, _25286_, _25287_, _25288_, _25289_, _25290_, _25291_, _25292_, _25293_, _25294_, _25295_, _25296_, _25297_, _25298_, _25299_, _25300_, _25301_, _25302_, _25303_, _25304_, _25305_, _25306_, _25307_, _25308_, _25309_, _25310_, _25311_, _25312_, _25313_, _25314_, _25315_, _25316_, _25317_, _25318_, _25319_, _25320_, _25321_, _25322_, _25323_, _25324_, _25325_, _25326_, _25327_, _25328_, _25329_, _25330_, _25331_, _25332_, _25333_, _25334_, _25335_, _25336_, _25337_, _25338_, _25339_, _25340_, _25341_, _25342_, _25343_, _25344_, _25345_, _25346_, _25347_, _25348_, _25349_, _25350_, _25351_, _25352_, _25353_, _25354_, _25355_, _25356_, _25357_, _25358_, _25359_, _25360_, _25361_, _25362_, _25363_, _25364_, _25365_, _25366_, _25367_, _25368_, _25369_, _25370_, _25371_, _25372_, _25373_, _25374_, _25375_, _25376_, _25377_, _25378_, _25379_, _25380_, _25381_, _25382_, _25383_, _25384_, _25385_, _25386_, _25387_, _25388_, _25389_, _25390_, _25391_, _25392_, _25393_, _25394_, _25395_, _25396_, _25397_, _25398_, _25399_, _25400_, _25401_, _25402_, _25403_, _25404_, _25405_, _25406_, _25407_, _25408_, _25409_, _25410_, _25411_, _25412_, _25413_, _25414_, _25415_, _25416_, _25417_, _25418_, _25419_, _25420_, _25421_, _25422_, _25423_, _25424_, _25425_, _25426_, _25427_, _25428_, _25429_, _25430_, _25431_, _25432_, _25433_, _25434_, _25435_, _25436_, _25437_, _25438_, _25439_, _25440_, _25441_, _25442_, _25443_, _25444_, _25445_, _25446_, _25447_, _25448_, _25449_, _25450_, _25451_, _25452_, _25453_, _25454_, _25455_, _25456_, _25457_, _25458_, _25459_, _25460_, _25461_, _25462_, _25463_, _25464_, _25465_, _25466_, _25467_, _25468_, _25469_, _25470_, _25471_, _25472_, _25473_, _25474_, _25475_, _25476_, _25477_, _25478_, _25479_, _25480_, _25481_, _25482_, _25483_, _25484_, _25485_, _25486_, _25487_, _25488_, _25489_, _25490_, _25491_, _25492_, _25493_, _25494_, _25495_, _25496_, _25497_, _25498_, _25499_, _25500_, _25501_, _25502_, _25503_, _25504_, _25505_, _25506_, _25507_, _25508_, _25509_, _25510_, _25511_, _25512_, _25513_, _25514_, _25515_, _25516_, _25517_, _25518_, _25519_, _25520_, _25521_, _25522_, _25523_, _25524_, _25525_, _25526_, _25527_, _25528_, _25529_, _25530_, _25531_, _25532_, _25533_, _25534_, _25535_, _25536_, _25537_, _25538_, _25539_, _25540_, _25541_, _25542_, _25543_, _25544_, _25545_, _25546_, _25547_, _25548_, _25549_, _25550_, _25551_, _25552_, _25553_, _25554_, _25555_, _25556_, _25557_, _25558_, _25559_, _25560_, _25561_, _25562_, _25563_, _25564_, _25565_, _25566_, _25567_, _25568_, _25569_, _25570_, _25571_, _25572_, _25573_, _25574_, _25575_, _25576_, _25577_, _25578_, _25579_, _25580_, _25581_, _25582_, _25583_, _25584_, _25585_, _25586_, _25587_, _25588_, _25589_, _25590_, _25591_, _25592_, _25593_, _25594_, _25595_, _25596_, _25597_, _25598_, _25599_, _25600_, _25601_, _25602_, _25603_, _25604_, _25605_, _25606_, _25607_, _25608_, _25609_, _25610_, _25611_, _25612_, _25613_, _25614_, _25615_, _25616_, _25617_, _25618_, _25619_, _25620_, _25621_, _25622_, _25623_, _25624_, _25625_, _25626_, _25627_, _25628_, _25629_, _25630_, _25631_, _25632_, _25633_, _25634_, _25635_, _25636_, _25637_, _25638_, _25639_, _25640_, _25641_, _25642_, _25643_, _25644_, _25645_, _25646_, _25647_, _25648_, _25649_, _25650_, _25651_, _25652_, _25653_, _25654_, _25655_, _25656_, _25657_, _25658_, _25659_, _25660_, _25661_, _25662_, _25663_, _25664_, _25665_, _25666_, _25667_, _25668_, _25669_, _25670_, _25671_, _25672_, _25673_, _25674_, _25675_, _25676_, _25677_, _25678_, _25679_, _25680_, _25681_, _25682_, _25683_, _25684_, _25685_, _25686_, _25687_, _25688_, _25689_, _25690_, _25691_, _25692_, _25693_, _25694_, _25695_, _25696_, _25697_, _25698_, _25699_, _25700_, _25701_, _25702_, _25703_, _25704_, _25705_, _25706_, _25707_, _25708_, _25709_, _25710_, _25711_, _25712_, _25713_, _25714_, _25715_, _25716_, _25717_, _25718_, _25719_, _25720_, _25721_, _25722_, _25723_, _25724_, _25725_, _25726_, _25727_, _25728_, _25729_, _25730_, _25731_, _25732_, _25733_, _25734_, _25735_, _25736_, _25737_, _25738_, _25739_, _25740_, _25741_, _25742_, _25743_, _25744_, _25745_, _25746_, _25747_, _25748_, _25749_, _25750_, _25751_, _25752_, _25753_, _25754_, _25755_, _25756_, _25757_, _25758_, _25759_, _25760_, _25761_, _25762_, _25763_, _25764_, _25765_, _25766_, _25767_, _25768_, _25769_, _25770_, _25771_, _25772_, _25773_, _25774_, _25775_, _25776_, _25777_, _25778_, _25779_, _25780_, _25781_, _25782_, _25783_, _25784_, _25785_, _25786_, _25787_, _25788_, _25789_, _25790_, _25791_, _25792_, _25793_, _25794_, _25795_, _25796_, _25797_, _25798_, _25799_, _25800_, _25801_, _25802_, _25803_, _25804_, _25805_, _25806_, _25807_, _25808_, _25809_, _25810_, _25811_, _25812_, _25813_, _25814_, _25815_, _25816_, _25817_, _25818_, _25819_, _25820_, _25821_, _25822_, _25823_, _25824_, _25825_, _25826_, _25827_, _25828_, _25829_, _25830_, _25831_, _25832_, _25833_, _25834_, _25835_, _25836_, _25837_, _25838_, _25839_, _25840_, _25841_, _25842_, _25843_, _25844_, _25845_, _25846_, _25847_, _25848_, _25849_, _25850_, _25851_, _25852_, _25853_, _25854_, _25855_, _25856_, _25857_, _25858_, _25859_, _25860_, _25861_, _25862_, _25863_, _25864_, _25865_, _25866_, _25867_, _25868_, _25869_, _25870_, _25871_, _25872_, _25873_, _25874_, _25875_, _25876_, _25877_, _25878_, _25879_, _25880_, _25881_, _25882_, _25883_, _25884_, _25885_, _25886_, _25887_, _25888_, _25889_, _25890_, _25891_, _25892_, _25893_, _25894_, _25895_, _25896_, _25897_, _25898_, _25899_, _25900_, _25901_, _25902_, _25903_, _25904_, _25905_, _25906_, _25907_, _25908_, _25909_, _25910_, _25911_, _25912_, _25913_, _25914_, _25915_, _25916_, _25917_, _25918_, _25919_, _25920_, _25921_, _25922_, _25923_, _25924_, _25925_, _25926_, _25927_, _25928_, _25929_, _25930_, _25931_, _25932_, _25933_, _25934_, _25935_, _25936_, _25937_, _25938_, _25939_, _25940_, _25941_, _25942_, _25943_, _25944_, _25945_, _25946_, _25947_, _25948_, _25949_, _25950_, _25951_, _25952_, _25953_, _25954_, _25955_, _25956_, _25957_, _25958_, _25959_, _25960_, _25961_, _25962_, _25963_, _25964_, _25965_, _25966_, _25967_, _25968_, _25969_, _25970_, _25971_, _25972_, _25973_, _25974_, _25975_, _25976_, _25977_, _25978_, _25979_, _25980_, _25981_, _25982_, _25983_, _25984_, _25985_, _25986_, _25987_, _25988_, _25989_, _25990_, _25991_, _25992_, _25993_, _25994_, _25995_, _25996_, _25997_, _25998_, _25999_, _26000_, _26001_, _26002_, _26003_, _26004_, _26005_, _26006_, _26007_, _26008_, _26009_, _26010_, _26011_, _26012_, _26013_, _26014_, _26015_, _26016_, _26017_, _26018_, _26019_, _26020_, _26021_, _26022_, _26023_, _26024_, _26025_, _26026_, _26027_, _26028_, _26029_, _26030_, _26031_, _26032_, _26033_, _26034_, _26035_, _26036_, _26037_, _26038_, _26039_, _26040_, _26041_, _26042_, _26043_, _26044_, _26045_, _26046_, _26047_, _26048_, _26049_, _26050_, _26051_, _26052_, _26053_, _26054_, _26055_, _26056_, _26057_, _26058_, _26059_, _26060_, _26061_, _26062_, _26063_, _26064_, _26065_, _26066_, _26067_, _26068_, _26069_, _26070_, _26071_, _26072_, _26073_, _26074_, _26075_, _26076_, _26077_, _26078_, _26079_, _26080_, _26081_, _26082_, _26083_, _26084_, _26085_, _26086_, _26087_, _26088_, _26089_, _26090_, _26091_, _26092_, _26093_, _26094_, _26095_, _26096_, _26097_, _26098_, _26099_, _26100_, _26101_, _26102_, _26103_, _26104_, _26105_, _26106_, _26107_, _26108_, _26109_, _26110_, _26111_, _26112_, _26113_, _26114_, _26115_, _26116_, _26117_, _26118_, _26119_, _26120_, _26121_, _26122_, _26123_, _26124_, _26125_, _26126_, _26127_, _26128_, _26129_, _26130_, _26131_, _26132_, _26133_, _26134_, _26135_, _26136_, _26137_, _26138_, _26139_, _26140_, _26141_, _26142_, _26143_, _26144_, _26145_, _26146_, _26147_, _26148_, _26149_, _26150_, _26151_, _26152_, _26153_, _26154_, _26155_, _26156_, _26157_, _26158_, _26159_, _26160_, _26161_, _26162_, _26163_, _26164_, _26165_, _26166_, _26167_, _26168_, _26169_, _26170_, _26171_, _26172_, _26173_, _26174_, _26175_, _26176_, _26177_, _26178_, _26179_, _26180_, _26181_, _26182_, _26183_, _26184_, _26185_, _26186_, _26187_, _26188_, _26189_, _26190_, _26191_, _26192_, _26193_, _26194_, _26195_, _26196_, _26197_, _26198_, _26199_, _26200_, _26201_, _26202_, _26203_, _26204_, _26205_, _26206_, _26207_, _26208_, _26209_, _26210_, _26211_, _26212_, _26213_, _26214_, _26215_, _26216_, _26217_, _26218_, _26219_, _26220_, _26221_, _26222_, _26223_, _26224_, _26225_, _26226_, _26227_, _26228_, _26229_, _26230_, _26231_, _26232_, _26233_, _26234_, _26235_, _26236_, _26237_, _26238_, _26239_, _26240_, _26241_, _26242_, _26243_, _26244_, _26245_, _26246_, _26247_, _26248_, _26249_, _26250_, _26251_, _26252_, _26253_, _26254_, _26255_, _26256_, _26257_, _26258_, _26259_, _26260_, _26261_, _26262_, _26263_, _26264_, _26265_, _26266_, _26267_, _26268_, _26269_, _26270_, _26271_, _26272_, _26273_, _26274_, _26275_, _26276_, _26277_, _26278_, _26279_, _26280_, _26281_, _26282_, _26283_, _26284_, _26285_, _26286_, _26287_, _26288_, _26289_, _26290_, _26291_, _26292_, _26293_, _26294_, _26295_, _26296_, _26297_, _26298_, _26299_, _26300_, _26301_, _26302_, _26303_, _26304_, _26305_, _26306_, _26307_, _26308_, _26309_, _26310_, _26311_, _26312_, _26313_, _26314_, _26315_, _26316_, _26317_, _26318_, _26319_, _26320_, _26321_, _26322_, _26323_, _26324_, _26325_, _26326_, _26327_, _26328_, _26329_, _26330_, _26331_, _26332_, _26333_, _26334_, _26335_, _26336_, _26337_, _26338_, _26339_, _26340_, _26341_, _26342_, _26343_, _26344_, _26345_, _26346_, _26347_, _26348_, _26349_, _26350_, _26351_, _26352_, _26353_, _26354_, _26355_, _26356_, _26357_, _26358_, _26359_, _26360_, _26361_, _26362_, _26363_, _26364_, _26365_, _26366_, _26367_, _26368_, _26369_, _26370_, _26371_, _26372_, _26373_, _26374_, _26375_, _26376_, _26377_, _26378_, _26379_, _26380_, _26381_, _26382_, _26383_, _26384_, _26385_, _26386_, _26387_, _26388_, _26389_, _26390_, _26391_, _26392_, _26393_, _26394_, _26395_, _26396_, _26397_, _26398_, _26399_, _26400_, _26401_, _26402_, _26403_, _26404_, _26405_, _26406_, _26407_, _26408_, _26409_, _26410_, _26411_, _26412_, _26413_, _26414_, _26415_, _26416_, _26417_, _26418_, _26419_, _26420_, _26421_, _26422_, _26423_, _26424_, _26425_, _26426_, _26427_, _26428_, _26429_, _26430_, _26431_, _26432_, _26433_, _26434_, _26435_, _26436_, _26437_, _26438_, _26439_, _26440_, _26441_, _26442_, _26443_, _26444_, _26445_, _26446_, _26447_, _26448_, _26449_, _26450_, _26451_, _26452_, _26453_, _26454_, _26455_, _26456_, _26457_, _26458_, _26459_, _26460_, _26461_, _26462_, _26463_, _26464_, _26465_, _26466_, _26467_, _26468_, _26469_, _26470_, _26471_, _26472_, _26473_, _26474_, _26475_, _26476_, _26477_, _26478_, _26479_, _26480_, _26481_, _26482_, _26483_, _26484_, _26485_, _26486_, _26487_, _26488_, _26489_, _26490_, _26491_, _26492_, _26493_, _26494_, _26495_, _26496_, _26497_, _26498_, _26499_, _26500_, _26501_, _26502_, _26503_, _26504_, _26505_, _26506_, _26507_, _26508_, _26509_, _26510_, _26511_, _26512_, _26513_, _26514_, _26515_, _26516_, _26517_, _26518_, _26519_, _26520_, _26521_, _26522_, _26523_, _26524_, _26525_, _26526_, _26527_, _26528_, _26529_, _26530_, _26531_, _26532_, _26533_, _26534_, _26535_, _26536_, _26537_, _26538_, _26539_, _26540_, _26541_, _26542_, _26543_, _26544_, _26545_, _26546_, _26547_, _26548_, _26549_, _26550_, _26551_, _26552_, _26553_, _26554_, _26555_, _26556_, _26557_, _26558_, _26559_, _26560_, _26561_, _26562_, _26563_, _26564_, _26565_, _26566_, _26567_, _26568_, _26569_, _26570_, _26571_, _26572_, _26573_, _26574_, _26575_, _26576_, _26577_, _26578_, _26579_, _26580_, _26581_, _26582_, _26583_, _26584_, _26585_, _26586_, _26587_, _26588_, _26589_, _26590_, _26591_, _26592_, _26593_, _26594_, _26595_, _26596_, _26597_, _26598_, _26599_, _26600_, _26601_, _26602_, _26603_, _26604_, _26605_, _26606_, _26607_, _26608_, _26609_, _26610_, _26611_, _26612_, _26613_, _26614_, _26615_, _26616_, _26617_, _26618_, _26619_, _26620_, _26621_, _26622_, _26623_, _26624_, _26625_, _26626_, _26627_, _26628_, _26629_, _26630_, _26631_, _26632_, _26633_, _26634_, _26635_, _26636_, _26637_, _26638_, _26639_, _26640_, _26641_, _26642_, _26643_, _26644_, _26645_, _26646_, _26647_, _26648_, _26649_, _26650_, _26651_, _26652_, _26653_, _26654_, _26655_, _26656_, _26657_, _26658_, _26659_, _26660_, _26661_, _26662_, _26663_, _26664_, _26665_, _26666_, _26667_, _26668_, _26669_, _26670_, _26671_, _26672_, _26673_, _26674_, _26675_, _26676_, _26677_, _26678_, _26679_, _26680_, _26681_, _26682_, _26683_, _26684_, _26685_, _26686_, _26687_, _26688_, _26689_, _26690_, _26691_, _26692_, _26693_, _26694_, _26695_, _26696_, _26697_, _26698_, _26699_, _26700_, _26701_, _26702_, _26703_, _26704_, _26705_, _26706_, _26707_, _26708_, _26709_, _26710_, _26711_, _26712_, _26713_, _26714_, _26715_, _26716_, _26717_, _26718_, _26719_, _26720_, _26721_, _26722_, _26723_, _26724_, _26725_, _26726_, _26727_, _26728_, _26729_, _26730_, _26731_, _26732_, _26733_, _26734_, _26735_, _26736_, _26737_, _26738_, _26739_, _26740_, _26741_, _26742_, _26743_, _26744_, _26745_, _26746_, _26747_, _26748_, _26749_, _26750_, _26751_, _26752_, _26753_, _26754_, _26755_, _26756_, _26757_, _26758_, _26759_, _26760_, _26761_, _26762_, _26763_, _26764_, _26765_, _26766_, _26767_, _26768_, _26769_, _26770_, _26771_, _26772_, _26773_, _26774_, _26775_, _26776_, _26777_, _26778_, _26779_, _26780_, _26781_, _26782_, _26783_, _26784_, _26785_, _26786_, _26787_, _26788_, _26789_, _26790_, _26791_, _26792_, _26793_, _26794_, _26795_, _26796_, _26797_, _26798_, _26799_, _26800_, _26801_, _26802_, _26803_, _26804_, _26805_, _26806_, _26807_, _26808_, _26809_, _26810_, _26811_, _26812_, _26813_, _26814_, _26815_, _26816_, _26817_, _26818_, _26819_, _26820_, _26821_, _26822_, _26823_, _26824_, _26825_, _26826_, _26827_, _26828_, _26829_, _26830_, _26831_, _26832_, _26833_, _26834_, _26835_, _26836_, _26837_, _26838_, _26839_, _26840_, _26841_, _26842_, _26843_, _26844_, _26845_, _26846_, _26847_, _26848_, _26849_, _26850_, _26851_, _26852_, _26853_, _26854_, _26855_, _26856_, _26857_, _26858_, _26859_, _26860_, _26861_, _26862_, _26863_, _26864_, _26865_, _26866_, _26867_, _26868_, _26869_, _26870_, _26871_, _26872_, _26873_, _26874_, _26875_, _26876_, _26877_, _26878_, _26879_, _26880_, _26881_, _26882_, _26883_, _26884_, _26885_, _26886_, _26887_, _26888_, _26889_, _26890_, _26891_, _26892_, _26893_, _26894_, _26895_, _26896_, _26897_, _26898_, _26899_, _26900_, _26901_, _26902_, _26903_, _26904_, _26905_, _26906_, _26907_, _26908_, _26909_, _26910_, _26911_, _26912_, _26913_, _26914_, _26915_, _26916_, _26917_, _26918_, _26919_, _26920_, _26921_, _26922_, _26923_, _26924_, _26925_, _26926_, _26927_, _26928_, _26929_, _26930_, _26931_, _26932_, _26933_, _26934_, _26935_, _26936_, _26937_, _26938_, _26939_, _26940_, _26941_, _26942_, _26943_, _26944_, _26945_, _26946_, _26947_, _26948_, _26949_, _26950_, _26951_, _26952_, _26953_, _26954_, _26955_, _26956_, _26957_, _26958_, _26959_, _26960_, _26961_, _26962_, _26963_, _26964_, _26965_, _26966_, _26967_, _26968_, _26969_, _26970_, _26971_, _26972_, _26973_, _26974_, _26975_, _26976_, _26977_, _26978_, _26979_, _26980_, _26981_, _26982_, _26983_, _26984_, _26985_, _26986_, _26987_, _26988_, _26989_, _26990_, _26991_, _26992_, _26993_, _26994_, _26995_, _26996_, _26997_, _26998_, _26999_, _27000_, _27001_, _27002_, _27003_, _27004_, _27005_, _27006_, _27007_, _27008_, _27009_, _27010_, _27011_, _27012_, _27013_, _27014_, _27015_, _27016_, _27017_, _27018_, _27019_, _27020_, _27021_, _27022_, _27023_, _27024_, _27025_, _27026_, _27027_, _27028_, _27029_, _27030_, _27031_, _27032_, _27033_, _27034_, _27035_, _27036_, _27037_, _27038_, _27039_, _27040_, _27041_, _27042_, _27043_, _27044_, _27045_, _27046_, _27047_, _27048_, _27049_, _27050_, _27051_, _27052_, _27053_, _27054_, _27055_, _27056_, _27057_, _27058_, _27059_, _27060_, _27061_, _27062_, _27063_, _27064_, _27065_, _27066_, _27067_, _27068_, _27069_, _27070_, _27071_, _27072_, _27073_, _27074_, _27075_, _27076_, _27077_, _27078_, _27079_, _27080_, _27081_, _27082_, _27083_, _27084_, _27085_, _27086_, _27087_, _27088_, _27089_, _27090_, _27091_, _27092_, _27093_, _27094_, _27095_, _27096_, _27097_, _27098_, _27099_, _27100_, _27101_, _27102_, _27103_, _27104_, _27105_, _27106_, _27107_, _27108_, _27109_, _27110_, _27111_, _27112_, _27113_, _27114_, _27115_, _27116_, _27117_, _27118_, _27119_, _27120_, _27121_, _27122_, _27123_, _27124_, _27125_, _27126_, _27127_, _27128_, _27129_, _27130_, _27131_, _27132_, _27133_, _27134_, _27135_, _27136_, _27137_, _27138_, _27139_, _27140_, _27141_, _27142_, _27143_, _27144_, _27145_, _27146_, _27147_, _27148_, _27149_, _27150_, _27151_, _27152_, _27153_, _27154_, _27155_, _27156_, _27157_, _27158_, _27159_, _27160_, _27161_, _27162_, _27163_, _27164_, _27165_, _27166_, _27167_, _27168_, _27169_, _27170_, _27171_, _27172_, _27173_, _27174_, _27175_, _27176_, _27177_, _27178_, _27179_, _27180_, _27181_, _27182_, _27183_, _27184_, _27185_, _27186_, _27187_, _27188_, _27189_, _27190_, _27191_, _27192_, _27193_, _27194_, _27195_, _27196_, _27197_, _27198_, _27199_, _27200_, _27201_, _27202_, _27203_, _27204_, _27205_, _27206_, _27207_, _27208_, _27209_, _27210_, _27211_, _27212_, _27213_, _27214_, _27215_, _27216_, _27217_, _27218_, _27219_, _27220_, _27221_, _27222_, _27223_, _27224_, _27225_, _27226_, _27227_, _27228_, _27229_, _27230_, _27231_, _27232_, _27233_, _27234_, _27235_, _27236_, _27237_, _27238_, _27239_, _27240_, _27241_, _27242_, _27243_, _27244_, _27245_, _27246_, _27247_, _27248_, _27249_, _27250_, _27251_, _27252_, _27253_, _27254_, _27255_, _27256_, _27257_, _27258_, _27259_, _27260_, _27261_, _27262_, _27263_, _27264_, _27265_, _27266_, _27267_, _27268_, _27269_, _27270_, _27271_, _27272_, _27273_, _27274_, _27275_, _27276_, _27277_, _27278_, _27279_, _27280_, _27281_, _27282_, _27283_, _27284_, _27285_, _27286_, _27287_, _27288_, _27289_, _27290_, _27291_, _27292_, _27293_, _27294_, _27295_, _27296_, _27297_, _27298_, _27299_, _27300_, _27301_, _27302_, _27303_, _27304_, _27305_, _27306_, _27307_, _27308_, _27309_, _27310_, _27311_, _27312_, _27313_, _27314_, _27315_, _27316_, _27317_, _27318_, _27319_, _27320_, _27321_, _27322_, _27323_, _27324_, _27325_, _27326_, _27327_, _27328_, _27329_, _27330_, _27331_, _27332_, _27333_, _27334_, _27335_, _27336_, _27337_, _27338_, _27339_, _27340_, _27341_, _27342_, _27343_, _27344_, _27345_, _27346_, _27347_, _27348_, _27349_, _27350_, _27351_, _27352_, _27353_, _27354_, _27355_, _27356_, _27357_, _27358_, _27359_, _27360_, _27361_, _27362_, _27363_, _27364_, _27365_, _27366_, _27367_, _27368_, _27369_, _27370_, _27371_, _27372_, _27373_, _27374_, _27375_, _27376_, _27377_, _27378_, _27379_, _27380_, _27381_, _27382_, _27383_, _27384_, _27385_, _27386_, _27387_, _27388_, _27389_, _27390_, _27391_, _27392_, _27393_, _27394_, _27395_, _27396_, _27397_, _27398_, _27399_, _27400_, _27401_, _27402_, _27403_, _27404_, _27405_, _27406_, _27407_, _27408_, _27409_, _27410_, _27411_, _27412_, _27413_, _27414_, _27415_, _27416_, _27417_, _27418_, _27419_, _27420_, _27421_, _27422_, _27423_, _27424_, _27425_, _27426_, _27427_, _27428_, _27429_, _27430_, _27431_, _27432_, _27433_, _27434_, _27435_, _27436_, _27437_, _27438_, _27439_, _27440_, _27441_, _27442_, _27443_, _27444_, _27445_, _27446_, _27447_, _27448_, _27449_, _27450_, _27451_, _27452_, _27453_, _27454_, _27455_, _27456_, _27457_, _27458_, _27459_, _27460_, _27461_, _27462_, _27463_, _27464_, _27465_, _27466_, _27467_, _27468_, _27469_, _27470_, _27471_, _27472_, _27473_, _27474_, _27475_, _27476_, _27477_, _27478_, _27479_, _27480_, _27481_, _27482_, _27483_, _27484_, _27485_, _27486_, _27487_, _27488_, _27489_, _27490_, _27491_, _27492_, _27493_, _27494_, _27495_, _27496_, _27497_, _27498_, _27499_, _27500_, _27501_, _27502_, _27503_, _27504_, _27505_, _27506_, _27507_, _27508_, _27509_, _27510_, _27511_, _27512_, _27513_, _27514_, _27515_, _27516_, _27517_, _27518_, _27519_, _27520_, _27521_, _27522_, _27523_, _27524_, _27525_, _27526_, _27527_, _27528_, _27529_, _27530_, _27531_, _27532_, _27533_, _27534_, _27535_, _27536_, _27537_, _27538_, _27539_, _27540_, _27541_, _27542_, _27543_, _27544_, _27545_, _27546_, _27547_, _27548_, _27549_, _27550_, _27551_, _27552_, _27553_, _27554_, _27555_, _27556_, _27557_, _27558_, _27559_, _27560_, _27561_, _27562_, _27563_, _27564_, _27565_, _27566_, _27567_, _27568_, _27569_, _27570_, _27571_, _27572_, _27573_, _27574_, _27575_, _27576_, _27577_, _27578_, _27579_, _27580_, _27581_, _27582_, _27583_, _27584_, _27585_, _27586_, _27587_, _27588_, _27589_, _27590_, _27591_, _27592_, _27593_, _27594_, _27595_, _27596_, _27597_, _27598_, _27599_, _27600_, _27601_, _27602_, _27603_, _27604_, _27605_, _27606_, _27607_, _27608_, _27609_, _27610_, _27611_, _27612_, _27613_, _27614_, _27615_, _27616_, _27617_, _27618_, _27619_, _27620_, _27621_, _27622_, _27623_, _27624_, _27625_, _27626_, _27627_, _27628_, _27629_, _27630_, _27631_, _27632_, _27633_, _27634_, _27635_, _27636_, _27637_, _27638_, _27639_, _27640_, _27641_, _27642_, _27643_, _27644_, _27645_, _27646_, _27647_, _27648_, _27649_, _27650_, _27651_, _27652_, _27653_, _27654_, _27655_, _27656_, _27657_, _27658_, _27659_, _27660_, _27661_, _27662_, _27663_, _27664_, _27665_, _27666_, _27667_, _27668_, _27669_, _27670_, _27671_, _27672_, _27673_, _27674_, _27675_, _27676_, _27677_, _27678_, _27679_, _27680_, _27681_, _27682_, _27683_, _27684_, _27685_, _27686_, _27687_, _27688_, _27689_, _27690_, _27691_, _27692_, _27693_, _27694_, _27695_, _27696_, _27697_, _27698_, _27699_, _27700_, _27701_, _27702_, _27703_, _27704_, _27705_, _27706_, _27707_, _27708_, _27709_, _27710_, _27711_, _27712_, _27713_, _27714_, _27715_, _27716_, _27717_, _27718_, _27719_, _27720_, _27721_, _27722_, _27723_, _27724_, _27725_, _27726_, _27727_, _27728_, _27729_, _27730_, _27731_, _27732_, _27733_, _27734_, _27735_, _27736_, _27737_, _27738_, _27739_, _27740_, _27741_, _27742_, _27743_, _27744_, _27745_, _27746_, _27747_, _27748_, _27749_, _27750_, _27751_, _27752_, _27753_, _27754_, _27755_, _27756_, _27757_, _27758_, _27759_, _27760_, _27761_, _27762_, _27763_, _27764_, _27765_, _27766_, _27767_, _27768_, _27769_, _27770_, _27771_, _27772_, _27773_, _27774_, _27775_, _27776_, _27777_, _27778_, _27779_, _27780_, _27781_, _27782_, _27783_, _27784_, _27785_, _27786_, _27787_, _27788_, _27789_, _27790_, _27791_, _27792_, _27793_, _27794_, _27795_, _27796_, _27797_, _27798_, _27799_, _27800_, _27801_, _27802_, _27803_, _27804_, _27805_, _27806_, _27807_, _27808_, _27809_, _27810_, _27811_, _27812_, _27813_, _27814_, _27815_, _27816_, _27817_, _27818_, _27819_, _27820_, _27821_, _27822_, _27823_, _27824_, _27825_, _27826_, _27827_, _27828_, _27829_, _27830_, _27831_, _27832_, _27833_, _27834_, _27835_, _27836_, _27837_, _27838_, _27839_, _27840_, _27841_, _27842_, _27843_, _27844_, _27845_, _27846_, _27847_, _27848_, _27849_, _27850_, _27851_, _27852_, _27853_, _27854_, _27855_, _27856_, _27857_, _27858_, _27859_, _27860_, _27861_, _27862_, _27863_, _27864_, _27865_, _27866_, _27867_, _27868_, _27869_, _27870_, _27871_, _27872_, _27873_, _27874_, _27875_, _27876_, _27877_, _27878_, _27879_, _27880_, _27881_, _27882_, _27883_, _27884_, _27885_, _27886_, _27887_, _27888_, _27889_, _27890_, _27891_, _27892_, _27893_, _27894_, _27895_, _27896_, _27897_, _27898_, _27899_, _27900_, _27901_, _27902_, _27903_, _27904_, _27905_, _27906_, _27907_, _27908_, _27909_, _27910_, _27911_, _27912_, _27913_, _27914_, _27915_, _27916_, _27917_, _27918_, _27919_, _27920_, _27921_, _27922_, _27923_, _27924_, _27925_, _27926_, _27927_, _27928_, _27929_, _27930_, _27931_, _27932_, _27933_, _27934_, _27935_, _27936_, _27937_, _27938_, _27939_, _27940_, _27941_, _27942_, _27943_, _27944_, _27945_, _27946_, _27947_, _27948_, _27949_, _27950_, _27951_, _27952_, _27953_, _27954_, _27955_, _27956_, _27957_, _27958_, _27959_, _27960_, _27961_, _27962_, _27963_, _27964_, _27965_, _27966_, _27967_, _27968_, _27969_, _27970_, _27971_, _27972_, _27973_, _27974_, _27975_, _27976_, _27977_, _27978_, _27979_, _27980_, _27981_, _27982_, _27983_, _27984_, _27985_, _27986_, _27987_, _27988_, _27989_, _27990_, _27991_, _27992_, _27993_, _27994_, _27995_, _27996_, _27997_, _27998_, _27999_, _28000_, _28001_, _28002_, _28003_, _28004_, _28005_, _28006_, _28007_, _28008_, _28009_, _28010_, _28011_, _28012_, _28013_, _28014_, _28015_, _28016_, _28017_, _28018_, _28019_, _28020_, _28021_, _28022_, _28023_, _28024_, _28025_, _28026_, _28027_, _28028_, _28029_, _28030_, _28031_, _28032_, _28033_, _28034_, _28035_, _28036_, _28037_, _28038_, _28039_, _28040_, _28041_, _28042_, _28043_, _28044_, _28045_, _28046_, _28047_, _28048_, _28049_, _28050_, _28051_, _28052_, _28053_, _28054_, _28055_, _28056_, _28057_, _28058_, _28059_, _28060_, _28061_, _28062_, _28063_, _28064_, _28065_, _28066_, _28067_, _28068_, _28069_, _28070_, _28071_, _28072_, _28073_, _28074_, _28075_, _28076_, _28077_, _28078_, _28079_, _28080_, _28081_, _28082_, _28083_, _28084_, _28085_, _28086_, _28087_, _28088_, _28089_, _28090_, _28091_, _28092_, _28093_, _28094_, _28095_, _28096_, _28097_, _28098_, _28099_, _28100_, _28101_, _28102_, _28103_, _28104_, _28105_, _28106_, _28107_, _28108_, _28109_, _28110_, _28111_, _28112_, _28113_, _28114_, _28115_, _28116_, _28117_, _28118_, _28119_, _28120_, _28121_, _28122_, _28123_, _28124_, _28125_, _28126_, _28127_, _28128_, _28129_, _28130_, _28131_, _28132_, _28133_, _28134_, _28135_, _28136_, _28137_, _28138_, _28139_, _28140_, _28141_, _28142_, _28143_, _28144_, _28145_, _28146_, _28147_, _28148_, _28149_, _28150_, _28151_, _28152_, _28153_, _28154_, _28155_, _28156_, _28157_, _28158_, _28159_, _28160_, _28161_, _28162_, _28163_, _28164_, _28165_, _28166_, _28167_, _28168_, _28169_, _28170_, _28171_, _28172_, _28173_, _28174_, _28175_, _28176_, _28177_, _28178_, _28179_, _28180_, _28181_, _28182_, _28183_, _28184_, _28185_, _28186_, _28187_, _28188_, _28189_, _28190_, _28191_, _28192_, _28193_, _28194_, _28195_, _28196_, _28197_, _28198_, _28199_, _28200_, _28201_, _28202_, _28203_, _28204_, _28205_, _28206_, _28207_, _28208_, _28209_, _28210_, _28211_, _28212_, _28213_, _28214_, _28215_, _28216_, _28217_, _28218_, _28219_, _28220_, _28221_, _28222_, _28223_, _28224_, _28225_, _28226_, _28227_, _28228_, _28229_, _28230_, _28231_, _28232_, _28233_, _28234_, _28235_, _28236_, _28237_, _28238_, _28239_, _28240_, _28241_, _28242_, _28243_, _28244_, _28245_, _28246_, _28247_, _28248_, _28249_, _28250_, _28251_, _28252_, _28253_, _28254_, _28255_, _28256_, _28257_, _28258_, _28259_, _28260_, _28261_, _28262_, _28263_, _28264_, _28265_, _28266_, _28267_, _28268_, _28269_, _28270_, _28271_, _28272_, _28273_, _28274_, _28275_, _28276_, _28277_, _28278_, _28279_, _28280_, _28281_, _28282_, _28283_, _28284_, _28285_, _28286_, _28287_, _28288_, _28289_, _28290_, _28291_, _28292_, _28293_, _28294_, _28295_, _28296_, _28297_, _28298_, _28299_, _28300_, _28301_, _28302_, _28303_, _28304_, _28305_, _28306_, _28307_, _28308_, _28309_, _28310_, _28311_, _28312_, _28313_, _28314_, _28315_, _28316_, _28317_, _28318_, _28319_, _28320_, _28321_, _28322_, _28323_, _28324_, _28325_, _28326_, _28327_, _28328_, _28329_, _28330_, _28331_, _28332_, _28333_, _28334_, _28335_, _28336_, _28337_, _28338_, _28339_, _28340_, _28341_, _28342_, _28343_, _28344_, _28345_, _28346_, _28347_, _28348_, _28349_, _28350_, _28351_, _28352_, _28353_, _28354_, _28355_, _28356_, _28357_, _28358_, _28359_, _28360_, _28361_, _28362_, _28363_, _28364_, _28365_, _28366_, _28367_, _28368_, _28369_, _28370_, _28371_, _28372_, _28373_, _28374_, _28375_, _28376_, _28377_, _28378_, _28379_, _28380_, _28381_, _28382_, _28383_, _28384_, _28385_, _28386_, _28387_, _28388_, _28389_, _28390_, _28391_, _28392_, _28393_, _28394_, _28395_, _28396_, _28397_, _28398_, _28399_, _28400_, _28401_, _28402_, _28403_, _28404_, _28405_, _28406_, _28407_, _28408_, _28409_, _28410_, _28411_, _28412_, _28413_, _28414_, _28415_, _28416_, _28417_, _28418_, _28419_, _28420_, _28421_, _28422_, _28423_, _28424_, _28425_, _28426_, _28427_, _28428_, _28429_, _28430_, _28431_, _28432_, _28433_, _28434_, _28435_, _28436_, _28437_, _28438_, _28439_, _28440_, _28441_, _28442_, _28443_, _28444_, _28445_, _28446_, _28447_, _28448_, _28449_, _28450_, _28451_, _28452_, _28453_, _28454_, _28455_, _28456_, _28457_, _28458_, _28459_, _28460_, _28461_, _28462_, _28463_, _28464_, _28465_, _28466_, _28467_, _28468_, _28469_, _28470_, _28471_, _28472_, _28473_, _28474_, _28475_, _28476_, _28477_, _28478_, _28479_, _28480_, _28481_, _28482_, _28483_, _28484_, _28485_, _28486_, _28487_, _28488_, _28489_, _28490_, _28491_, _28492_, _28493_, _28494_, _28495_, _28496_, _28497_, _28498_, _28499_, _28500_, _28501_, _28502_, _28503_, _28504_, _28505_, _28506_, _28507_, _28508_, _28509_, _28510_, _28511_, _28512_, _28513_, _28514_, _28515_, _28516_, _28517_, _28518_, _28519_, _28520_, _28521_, _28522_, _28523_, _28524_, _28525_, _28526_, _28527_, _28528_, _28529_, _28530_, _28531_, _28532_, _28533_, _28534_, _28535_, _28536_, _28537_, _28538_, _28539_, _28540_, _28541_, _28542_, _28543_, _28544_, _28545_, _28546_, _28547_, _28548_, _28549_, _28550_, _28551_, _28552_, _28553_, _28554_, _28555_, _28556_, _28557_, _28558_, _28559_, _28560_, _28561_, _28562_, _28563_, _28564_, _28565_, _28566_, _28567_, _28568_, _28569_, _28570_, _28571_, _28572_, _28573_, _28574_, _28575_, _28576_, _28577_, _28578_, _28579_, _28580_, _28581_, _28582_, _28583_, _28584_, _28585_, _28586_, _28587_, _28588_, _28589_, _28590_, _28591_, _28592_, _28593_, _28594_, _28595_, _28596_, _28597_, _28598_, _28599_, _28600_, _28601_, _28602_, _28603_, _28604_, _28605_, _28606_, _28607_, _28608_, _28609_, _28610_, _28611_, _28612_, _28613_, _28614_, _28615_, _28616_, _28617_, _28618_, _28619_, _28620_, _28621_, _28622_, _28623_, _28624_, _28625_, _28626_, _28627_, _28628_, _28629_, _28630_, _28631_, _28632_, _28633_, _28634_, _28635_, _28636_, _28637_, _28638_, _28639_, _28640_, _28641_, _28642_, _28643_, _28644_, _28645_, _28646_, _28647_, _28648_, _28649_, _28650_, _28651_, _28652_, _28653_, _28654_, _28655_, _28656_, _28657_, _28658_, _28659_, _28660_, _28661_, _28662_, _28663_, _28664_, _28665_, _28666_, _28667_, _28668_, _28669_, _28670_, _28671_, _28672_, _28673_, _28674_, _28675_, _28676_, _28677_, _28678_, _28679_, _28680_, _28681_, _28682_, _28683_, _28684_, _28685_, _28686_, _28687_, _28688_, _28689_, _28690_, _28691_, _28692_, _28693_, _28694_, _28695_, _28696_, _28697_, _28698_, _28699_, _28700_, _28701_, _28702_, _28703_, _28704_, _28705_, _28706_, _28707_, _28708_, _28709_, _28710_, _28711_, _28712_, _28713_, _28714_, _28715_, _28716_, _28717_, _28718_, _28719_, _28720_, _28721_, _28722_, _28723_, _28724_, _28725_, _28726_, _28727_, _28728_, _28729_, _28730_, _28731_, _28732_, _28733_, _28734_, _28735_, _28736_, _28737_, _28738_, _28739_, _28740_, _28741_, _28742_, _28743_, _28744_, _28745_, _28746_, _28747_, _28748_, _28749_, _28750_, _28751_, _28752_, _28753_, _28754_, _28755_, _28756_, _28757_, _28758_, _28759_, _28760_, _28761_, _28762_, _28763_, _28764_, _28765_, _28766_, _28767_, _28768_, _28769_, _28770_, _28771_, _28772_, _28773_, _28774_, _28775_, _28776_, _28777_, _28778_, _28779_, _28780_, _28781_, _28782_, _28783_, _28784_, _28785_, _28786_, _28787_, _28788_, _28789_, _28790_, _28791_, _28792_, _28793_, _28794_, _28795_, _28796_, _28797_, _28798_, _28799_, _28800_, _28801_, _28802_, _28803_, _28804_, _28805_, _28806_, _28807_, _28808_, _28809_, _28810_, _28811_, _28812_, _28813_, _28814_, _28815_, _28816_, _28817_, _28818_, _28819_, _28820_, _28821_, _28822_, _28823_, _28824_, _28825_, _28826_, _28827_, _28828_, _28829_, _28830_, _28831_, _28832_, _28833_, _28834_, _28835_, _28836_, _28837_, _28838_, _28839_, _28840_, _28841_, _28842_, _28843_, _28844_, _28845_, _28846_, _28847_, _28848_, _28849_, _28850_, _28851_, _28852_, _28853_, _28854_, _28855_, _28856_, _28857_, _28858_, _28859_, _28860_, _28861_, _28862_, _28863_, _28864_, _28865_, _28866_, _28867_, _28868_, _28869_, _28870_, _28871_, _28872_, _28873_, _28874_, _28875_, _28876_, _28877_, _28878_, _28879_, _28880_, _28881_, _28882_, _28883_, _28884_, _28885_, _28886_, _28887_, _28888_, _28889_, _28890_, _28891_, _28892_, _28893_, _28894_, _28895_, _28896_, _28897_, _28898_, _28899_, _28900_, _28901_, _28902_, _28903_, _28904_, _28905_, _28906_, _28907_, _28908_, _28909_, _28910_, _28911_, _28912_, _28913_, _28914_, _28915_, _28916_, _28917_, _28918_, _28919_, _28920_, _28921_, _28922_, _28923_, _28924_, _28925_, _28926_, _28927_, _28928_, _28929_, _28930_, _28931_, _28932_, _28933_, _28934_, _28935_, _28936_, _28937_, _28938_, _28939_, _28940_, _28941_, _28942_, _28943_, _28944_, _28945_, _28946_, _28947_, _28948_, _28949_, _28950_, _28951_, _28952_, _28953_, _28954_, _28955_, _28956_, _28957_, _28958_, _28959_, _28960_, _28961_, _28962_, _28963_, _28964_, _28965_, _28966_, _28967_, _28968_, _28969_, _28970_, _28971_, _28972_, _28973_, _28974_, _28975_, _28976_, _28977_, _28978_, _28979_, _28980_, _28981_, _28982_, _28983_, _28984_, _28985_, _28986_, _28987_, _28988_, _28989_, _28990_, _28991_, _28992_, _28993_, _28994_, _28995_, _28996_, _28997_, _28998_, _28999_, _29000_, _29001_, _29002_, _29003_, _29004_, _29005_, _29006_, _29007_, _29008_, _29009_, _29010_, _29011_, _29012_, _29013_, _29014_, _29015_, _29016_, _29017_, _29018_, _29019_, _29020_, _29021_, _29022_, _29023_, _29024_, _29025_, _29026_, _29027_, _29028_, _29029_, _29030_, _29031_, _29032_, _29033_, _29034_, _29035_, _29036_, _29037_, _29038_, _29039_, _29040_, _29041_, _29042_, _29043_, _29044_, _29045_, _29046_, _29047_, _29048_, _29049_, _29050_, _29051_, _29052_, _29053_, _29054_, _29055_, _29056_, _29057_, _29058_, _29059_, _29060_, _29061_, _29062_, _29063_, _29064_, _29065_, _29066_, _29067_, _29068_, _29069_, _29070_, _29071_, _29072_, _29073_, _29074_, _29075_, _29076_, _29077_, _29078_, _29079_, _29080_, _29081_, _29082_, _29083_, _29084_, _29085_, _29086_, _29087_, _29088_, _29089_, _29090_, _29091_, _29092_, _29093_, _29094_, _29095_, _29096_, _29097_, _29098_, _29099_, _29100_, _29101_, _29102_, _29103_, _29104_, _29105_, _29106_, _29107_, _29108_, _29109_, _29110_, _29111_, _29112_, _29113_, _29114_, _29115_, _29116_, _29117_, _29118_, _29119_, _29120_, _29121_, _29122_, _29123_, _29124_, _29125_, _29126_, _29127_, _29128_, _29129_, _29130_, _29131_, _29132_, _29133_, _29134_, _29135_, _29136_, _29137_, _29138_, _29139_, _29140_, _29141_, _29142_, _29143_, _29144_, _29145_, _29146_, _29147_, _29148_, _29149_, _29150_, _29151_, _29152_, _29153_, _29154_, _29155_, _29156_, _29157_, _29158_, _29159_, _29160_, _29161_, _29162_, _29163_, _29164_, _29165_, _29166_, _29167_, _29168_, _29169_, _29170_, _29171_, _29172_, _29173_, _29174_, _29175_, _29176_, _29177_, _29178_, _29179_, _29180_, _29181_, _29182_, _29183_, _29184_, _29185_, _29186_, _29187_, _29188_, _29189_, _29190_, _29191_, _29192_, _29193_, _29194_, _29195_, _29196_, _29197_, _29198_, _29199_, _29200_, _29201_, _29202_, _29203_, _29204_, _29205_, _29206_, _29207_, _29208_, _29209_, _29210_, _29211_, _29212_, _29213_, _29214_, _29215_, _29216_, _29217_, _29218_, _29219_, _29220_, _29221_, _29222_, _29223_, _29224_, _29225_, _29226_, _29227_, _29228_, _29229_, _29230_, _29231_, _29232_, _29233_, _29234_, _29235_, _29236_, _29237_, _29238_, _29239_, _29240_, _29241_, _29242_, _29243_, _29244_, _29245_, _29246_, _29247_, _29248_, _29249_, _29250_, _29251_, _29252_, _29253_, _29254_, _29255_, _29256_, _29257_, _29258_, _29259_, _29260_, _29261_, _29262_, _29263_, _29264_, _29265_, _29266_, _29267_, _29268_, _29269_, _29270_, _29271_, _29272_, _29273_, _29274_, _29275_, _29276_, _29277_, _29278_, _29279_, _29280_, _29281_, _29282_, _29283_, _29284_, _29285_, _29286_, _29287_, _29288_, _29289_, _29290_, _29291_, _29292_, _29293_, _29294_, _29295_, _29296_, _29297_, _29298_, _29299_, _29300_, _29301_, _29302_, _29303_, _29304_, _29305_, _29306_, _29307_, _29308_, _29309_, _29310_, _29311_, _29312_, _29313_, _29314_, _29315_, _29316_, _29317_, _29318_, _29319_, _29320_, _29321_, _29322_, _29323_, _29324_, _29325_, _29326_, _29327_, _29328_, _29329_, _29330_, _29331_, _29332_, _29333_, _29334_, _29335_, _29336_, _29337_, _29338_, _29339_, _29340_, _29341_, _29342_, _29343_, _29344_, _29345_, _29346_, _29347_, _29348_, _29349_, _29350_, _29351_, _29352_, _29353_, _29354_, _29355_, _29356_, _29357_, _29358_, _29359_, _29360_, _29361_, _29362_, _29363_, _29364_, _29365_, _29366_, _29367_, _29368_, _29369_, _29370_, _29371_, _29372_, _29373_, _29374_, _29375_, _29376_, _29377_, _29378_, _29379_, _29380_, _29381_, _29382_, _29383_, _29384_, _29385_, _29386_, _29387_, _29388_, _29389_, _29390_, _29391_, _29392_, _29393_, _29394_, _29395_, _29396_, _29397_, _29398_, _29399_, _29400_, _29401_, _29402_, _29403_, _29404_, _29405_, _29406_, _29407_, _29408_, _29409_, _29410_, _29411_, _29412_, _29413_, _29414_, _29415_, _29416_, _29417_, _29418_, _29419_, _29420_, _29421_, _29422_, _29423_, _29424_, _29425_, _29426_, _29427_, _29428_, _29429_, _29430_, _29431_, _29432_, _29433_, _29434_, _29435_, _29436_, _29437_, _29438_, _29439_, _29440_, _29441_, _29442_, _29443_, _29444_, _29445_, _29446_, _29447_, _29448_, _29449_, _29450_, _29451_, _29452_, _29453_, _29454_, _29455_, _29456_, _29457_, _29458_, _29459_, _29460_, _29461_, _29462_, _29463_, _29464_, _29465_, _29466_, _29467_, _29468_, _29469_, _29470_, _29471_, _29472_, _29473_, _29474_, _29475_, _29476_, _29477_, _29478_, _29479_, _29480_, _29481_, _29482_, _29483_, _29484_, _29485_, _29486_, _29487_, _29488_, _29489_, _29490_, _29491_, _29492_, _29493_, _29494_, _29495_, _29496_, _29497_, _29498_, _29499_, _29500_, _29501_, _29502_, _29503_, _29504_, _29505_, _29506_, _29507_, _29508_, _29509_, _29510_, _29511_, _29512_, _29513_, _29514_, _29515_, _29516_, _29517_, _29518_, _29519_, _29520_, _29521_, _29522_, _29523_, _29524_, _29525_, _29526_, _29527_, _29528_, _29529_, _29530_, _29531_, _29532_, _29533_, _29534_, _29535_, _29536_, _29537_, _29538_, _29539_, _29540_, _29541_, _29542_, _29543_, _29544_, _29545_, _29546_, _29547_, _29548_, _29549_, _29550_, _29551_, _29552_, _29553_, _29554_, _29555_, _29556_, _29557_, _29558_, _29559_, _29560_, _29561_, _29562_, _29563_, _29564_, _29565_, _29566_, _29567_, _29568_, _29569_, _29570_, _29571_, _29572_, _29573_, _29574_, _29575_, _29576_, _29577_, _29578_, _29579_, _29580_, _29581_, _29582_, _29583_, _29584_, _29585_, _29586_, _29587_, _29588_, _29589_, _29590_, _29591_, _29592_, _29593_, _29594_, _29595_, _29596_, _29597_, _29598_, _29599_, _29600_, _29601_, _29602_, _29603_, _29604_, _29605_, _29606_, _29607_, _29608_, _29609_, _29610_, _29611_, _29612_, _29613_, _29614_, _29615_, _29616_, _29617_, _29618_, _29619_, _29620_, _29621_, _29622_, _29623_, _29624_, _29625_, _29626_, _29627_, _29628_, _29629_, _29630_, _29631_, _29632_, _29633_, _29634_, _29635_, _29636_, _29637_, _29638_, _29639_, _29640_, _29641_, _29642_, _29643_, _29644_, _29645_, _29646_, _29647_, _29648_, _29649_, _29650_, _29651_, _29652_, _29653_, _29654_, _29655_, _29656_, _29657_, _29658_, _29659_, _29660_, _29661_, _29662_, _29663_, _29664_, _29665_, _29666_, _29667_, _29668_, _29669_, _29670_, _29671_, _29672_, _29673_, _29674_, _29675_, _29676_, _29677_, _29678_, _29679_, _29680_, _29681_, _29682_, _29683_, _29684_, _29685_, _29686_, _29687_, _29688_, _29689_, _29690_, _29691_, _29692_, _29693_, _29694_, _29695_, _29696_, _29697_, _29698_, _29699_, _29700_, _29701_, _29702_, _29703_, _29704_, _29705_, _29706_, _29707_, _29708_, _29709_, _29710_, _29711_, _29712_, _29713_, _29714_, _29715_, _29716_, _29717_, _29718_, _29719_, _29720_, _29721_, _29722_, _29723_, _29724_, _29725_, _29726_, _29727_, _29728_, _29729_, _29730_, _29731_, _29732_, _29733_, _29734_, _29735_, _29736_, _29737_, _29738_, _29739_, _29740_, _29741_, _29742_, _29743_, _29744_, _29745_, _29746_, _29747_, _29748_, _29749_, _29750_, _29751_, _29752_, _29753_, _29754_, _29755_, _29756_, _29757_, _29758_, _29759_, _29760_, _29761_, _29762_, _29763_, _29764_, _29765_, _29766_, _29767_, _29768_, _29769_, _29770_, _29771_, _29772_, _29773_, _29774_, _29775_, _29776_, _29777_, _29778_, _29779_, _29780_, _29781_, _29782_, _29783_, _29784_, _29785_, _29786_, _29787_, _29788_, _29789_, _29790_, _29791_, _29792_, _29793_, _29794_, _29795_, _29796_, _29797_, _29798_, _29799_, _29800_, _29801_, _29802_, _29803_, _29804_, _29805_, _29806_, _29807_, _29808_, _29809_, _29810_, _29811_, _29812_, _29813_, _29814_, _29815_, _29816_, _29817_, _29818_, _29819_, _29820_, _29821_, _29822_, _29823_, _29824_, _29825_, _29826_, _29827_, _29828_, _29829_, _29830_, _29831_, _29832_, _29833_, _29834_, _29835_, _29836_, _29837_, _29838_, _29839_, _29840_, _29841_, _29842_, _29843_, _29844_, _29845_, _29846_, _29847_, _29848_, _29849_, _29850_, _29851_, _29852_, _29853_, _29854_, _29855_, _29856_, _29857_, _29858_, _29859_, _29860_, _29861_, _29862_, _29863_, _29864_, _29865_, _29866_, _29867_, _29868_, _29869_, _29870_, _29871_, _29872_, _29873_, _29874_, _29875_, _29876_, _29877_, _29878_, _29879_, _29880_, _29881_, _29882_, _29883_, _29884_, _29885_, _29886_, _29887_, _29888_, _29889_, _29890_, _29891_, _29892_, _29893_, _29894_, _29895_, _29896_, _29897_, _29898_, _29899_, _29900_, _29901_, _29902_, _29903_, _29904_, _29905_, _29906_, _29907_, _29908_, _29909_, _29910_, _29911_, _29912_, _29913_, _29914_, _29915_, _29916_, _29917_, _29918_, _29919_, _29920_, _29921_, _29922_, _29923_, _29924_, _29925_, _29926_, _29927_, _29928_, _29929_, _29930_, _29931_, _29932_, _29933_, _29934_, _29935_, _29936_, _29937_, _29938_, _29939_, _29940_, _29941_, _29942_, _29943_, _29944_, _29945_, _29946_, _29947_, _29948_, _29949_, _29950_, _29951_, _29952_, _29953_, _29954_, _29955_, _29956_, _29957_, _29958_, _29959_, _29960_, _29961_, _29962_, _29963_, _29964_, _29965_, _29966_, _29967_, _29968_, _29969_, _29970_, _29971_, _29972_, _29973_, _29974_, _29975_, _29976_, _29977_, _29978_, _29979_, _29980_, _29981_, _29982_, _29983_, _29984_, _29985_, _29986_, _29987_, _29988_, _29989_, _29990_, _29991_, _29992_, _29993_, _29994_, _29995_, _29996_, _29997_, _29998_, _29999_, _30000_, _30001_, _30002_, _30003_, _30004_, _30005_, _30006_, _30007_, _30008_, _30009_, _30010_, _30011_, _30012_, _30013_, _30014_, _30015_, _30016_, _30017_, _30018_, _30019_, _30020_, _30021_, _30022_, _30023_, _30024_, _30025_, _30026_, _30027_, _30028_, _30029_, _30030_, _30031_, _30032_, _30033_, _30034_, _30035_, _30036_, _30037_, _30038_, _30039_, _30040_, _30041_, _30042_, _30043_, _30044_, _30045_, _30046_, _30047_, _30048_, _30049_, _30050_, _30051_, _30052_, _30053_, _30054_, _30055_, _30056_, _30057_, _30058_, _30059_, _30060_, _30061_, _30062_, _30063_, _30064_, _30065_, _30066_, _30067_, _30068_, _30069_, _30070_, _30071_, _30072_, _30073_, _30074_, _30075_, _30076_, _30077_, _30078_, _30079_, _30080_, _30081_, _30082_, _30083_, _30084_, _30085_, _30086_, _30087_, _30088_, _30089_, _30090_, _30091_, _30092_, _30093_, _30094_, _30095_, _30096_, _30097_, _30098_, _30099_, _30100_, _30101_, _30102_, _30103_, _30104_, _30105_, _30106_, _30107_, _30108_, _30109_, _30110_, _30111_, _30112_, _30113_, _30114_, _30115_, _30116_, _30117_, _30118_, _30119_, _30120_, _30121_, _30122_, _30123_, _30124_, _30125_, _30126_, _30127_, _30128_, _30129_, _30130_, _30131_, _30132_, _30133_, _30134_, _30135_, _30136_, _30137_, _30138_, _30139_, _30140_, _30141_, _30142_, _30143_, _30144_, _30145_, _30146_, _30147_, _30148_, _30149_, _30150_, _30151_, _30152_, _30153_, _30154_, _30155_, _30156_, _30157_, _30158_, _30159_, _30160_, _30161_, _30162_, _30163_, _30164_, _30165_, _30166_, _30167_, _30168_, _30169_, _30170_, _30171_, _30172_, _30173_, _30174_, _30175_, _30176_, _30177_, _30178_, _30179_, _30180_, _30181_, _30182_, _30183_, _30184_, _30185_, _30186_, _30187_, _30188_, _30189_, _30190_, _30191_, _30192_, _30193_, _30194_, _30195_, _30196_, _30197_, _30198_, _30199_, _30200_, _30201_, _30202_, _30203_, _30204_, _30205_, _30206_, _30207_, _30208_, _30209_, _30210_, _30211_, _30212_, _30213_, _30214_, _30215_, _30216_, _30217_, _30218_, _30219_, _30220_, _30221_, _30222_, _30223_, _30224_, _30225_, _30226_, _30227_, _30228_, _30229_, _30230_, _30231_, _30232_, _30233_, _30234_, _30235_, _30236_, _30237_, _30238_, _30239_, _30240_, _30241_, _30242_, _30243_, _30244_, _30245_, _30246_, _30247_, _30248_, _30249_, _30250_, _30251_, _30252_, _30253_, _30254_, _30255_, _30256_, _30257_, _30258_, _30259_, _30260_, _30261_, _30262_, _30263_, _30264_, _30265_, _30266_, _30267_, _30268_, _30269_, _30270_, _30271_, _30272_, _30273_, _30274_, _30275_, _30276_, _30277_, _30278_, _30279_, _30280_, _30281_, _30282_, _30283_, _30284_, _30285_, _30286_, _30287_, _30288_, _30289_, _30290_, _30291_, _30292_, _30293_, _30294_, _30295_, _30296_, _30297_, _30298_, _30299_, _30300_, _30301_, _30302_, _30303_, _30304_, _30305_, _30306_, _30307_, _30308_, _30309_, _30310_, _30311_, _30312_, _30313_, _30314_, _30315_, _30316_, _30317_, _30318_, _30319_, _30320_, _30321_, _30322_, _30323_, _30324_, _30325_, _30326_, _30327_, _30328_, _30329_, _30330_, _30331_, _30332_, _30333_, _30334_, _30335_, _30336_, _30337_, _30338_, _30339_, _30340_, _30341_, _30342_, _30343_, _30344_, _30345_, _30346_, _30347_, _30348_, _30349_, _30350_, _30351_, _30352_, _30353_, _30354_, _30355_, _30356_, _30357_, _30358_, _30359_, _30360_, _30361_, _30362_, _30363_, _30364_, _30365_, _30366_, _30367_, _30368_, _30369_, _30370_, _30371_, _30372_, _30373_, _30374_, _30375_, _30376_, _30377_, _30378_, _30379_, _30380_, _30381_, _30382_, _30383_, _30384_, _30385_, _30386_, _30387_, _30388_, _30389_, _30390_, _30391_, _30392_, _30393_, _30394_, _30395_, _30396_, _30397_, _30398_, _30399_, _30400_, _30401_, _30402_, _30403_, _30404_, _30405_, _30406_, _30407_, _30408_, _30409_, _30410_, _30411_, _30412_, _30413_, _30414_, _30415_, _30416_, _30417_, _30418_, _30419_, _30420_, _30421_, _30422_, _30423_, _30424_, _30425_, _30426_, _30427_, _30428_, _30429_, _30430_, _30431_, _30432_, _30433_, _30434_, _30435_, _30436_, _30437_, _30438_, _30439_, _30440_, _30441_, _30442_, _30443_, _30444_, _30445_, _30446_, _30447_, _30448_, _30449_, _30450_, _30451_, _30452_, _30453_, _30454_, _30455_, _30456_, _30457_, _30458_, _30459_, _30460_, _30461_, _30462_, _30463_, _30464_, _30465_, _30466_, _30467_, _30468_, _30469_, _30470_, _30471_, _30472_, _30473_, _30474_, _30475_, _30476_, _30477_, _30478_, _30479_, _30480_, _30481_, _30482_, _30483_, _30484_, _30485_, _30486_, _30487_, _30488_, _30489_, _30490_, _30491_, _30492_, _30493_, _30494_, _30495_, _30496_, _30497_, _30498_, _30499_, _30500_, _30501_, _30502_, _30503_, _30504_, _30505_, _30506_, _30507_, _30508_, _30509_, _30510_, _30511_, _30512_, _30513_, _30514_, _30515_, _30516_, _30517_, _30518_, _30519_, _30520_, _30521_, _30522_, _30523_, _30524_, _30525_, _30526_, _30527_, _30528_, _30529_, _30530_, _30531_, _30532_, _30533_, _30534_, _30535_, _30536_, _30537_, _30538_, _30539_, _30540_, _30541_, _30542_, _30543_, _30544_, _30545_, _30546_, _30547_, _30548_, _30549_, _30550_, _30551_, _30552_, _30553_, _30554_, _30555_, _30556_, _30557_, _30558_, _30559_, _30560_, _30561_, _30562_, _30563_, _30564_, _30565_, _30566_, _30567_, _30568_, _30569_, _30570_, _30571_, _30572_, _30573_, _30574_, _30575_, _30576_, _30577_, _30578_, _30579_, _30580_, _30581_, _30582_, _30583_, _30584_, _30585_, _30586_, _30587_, _30588_, _30589_, _30590_, _30591_, _30592_, _30593_, _30594_, _30595_, _30596_, _30597_, _30598_, _30599_, _30600_, _30601_, _30602_, _30603_, _30604_, _30605_, _30606_, _30607_, _30608_, _30609_, _30610_, _30611_, _30612_, _30613_, _30614_, _30615_, _30616_, _30617_, _30618_, _30619_, _30620_, _30621_, _30622_, _30623_, _30624_, _30625_, _30626_, _30627_, _30628_, _30629_, _30630_, _30631_, _30632_, _30633_, _30634_, _30635_, _30636_, _30637_, _30638_, _30639_, _30640_, _30641_, _30642_, _30643_, _30644_, _30645_, _30646_, _30647_, _30648_, _30649_, _30650_, _30651_, _30652_, _30653_, _30654_, _30655_, _30656_, _30657_, _30658_, _30659_, _30660_, _30661_, _30662_, _30663_, _30664_, _30665_, _30666_, _30667_, _30668_, _30669_, _30670_, _30671_, _30672_, _30673_, _30674_, _30675_, _30676_, _30677_, _30678_, _30679_, _30680_, _30681_, _30682_, _30683_, _30684_, _30685_, _30686_, _30687_, _30688_, _30689_, _30690_, _30691_, _30692_, _30693_, _30694_, _30695_, _30696_, _30697_, _30698_, _30699_, _30700_, _30701_, _30702_, _30703_, _30704_, _30705_, _30706_, _30707_, _30708_, _30709_, _30710_, _30711_, _30712_, _30713_, _30714_, _30715_, _30716_, _30717_, _30718_, _30719_, _30720_, _30721_, _30722_, _30723_, _30724_, _30725_, _30726_, _30727_, _30728_, _30729_, _30730_, _30731_, _30732_, _30733_, _30734_, _30735_, _30736_, _30737_, _30738_, _30739_, _30740_, _30741_, _30742_, _30743_, _30744_, _30745_, _30746_, _30747_, _30748_, _30749_, _30750_, _30751_, _30752_, _30753_, _30754_, _30755_, _30756_, _30757_, _30758_, _30759_, _30760_, _30761_, _30762_, _30763_, _30764_, _30765_, _30766_, _30767_, _30768_, _30769_, _30770_, _30771_, _30772_, _30773_, _30774_, _30775_, _30776_, _30777_, _30778_, _30779_, _30780_, _30781_, _30782_, _30783_, _30784_, _30785_, _30786_, _30787_, _30788_, _30789_, _30790_, _30791_, _30792_, _30793_, _30794_, _30795_, _30796_, _30797_, _30798_, _30799_, _30800_, _30801_, _30802_, _30803_, _30804_, _30805_, _30806_, _30807_, _30808_, _30809_, _30810_, _30811_, _30812_, _30813_, _30814_, _30815_, _30816_, _30817_, _30818_, _30819_, _30820_, _30821_, _30822_, _30823_, _30824_, _30825_, _30826_, _30827_, _30828_, _30829_, _30830_, _30831_, _30832_, _30833_, _30834_, _30835_, _30836_, _30837_, _30838_, _30839_, _30840_, _30841_, _30842_, _30843_, _30844_, _30845_, _30846_, _30847_, _30848_, _30849_, _30850_, _30851_, _30852_, _30853_, _30854_, _30855_, _30856_, _30857_, _30858_, _30859_, _30860_, _30861_, _30862_, _30863_, _30864_, _30865_, _30866_, _30867_, _30868_, _30869_, _30870_, _30871_, _30872_, _30873_, _30874_, _30875_, _30876_, _30877_, _30878_, _30879_, _30880_, _30881_, _30882_, _30883_, _30884_, _30885_, _30886_, _30887_, _30888_, _30889_, _30890_, _30891_, _30892_, _30893_, _30894_, _30895_, _30896_, _30897_, _30898_, _30899_, _30900_, _30901_, _30902_, _30903_, _30904_, _30905_, _30906_, _30907_, _30908_, _30909_, _30910_, _30911_, _30912_, _30913_, _30914_, _30915_, _30916_, _30917_, _30918_, _30919_, _30920_, _30921_, _30922_, _30923_, _30924_, _30925_, _30926_, _30927_, _30928_, _30929_, _30930_, _30931_, _30932_, _30933_, _30934_, _30935_, _30936_, _30937_, _30938_, _30939_, _30940_, _30941_, _30942_, _30943_, _30944_, _30945_, _30946_, _30947_, _30948_, _30949_, _30950_, _30951_, _30952_, _30953_, _30954_, _30955_, _30956_, _30957_, _30958_, _30959_, _30960_, _30961_, _30962_, _30963_, _30964_, _30965_, _30966_, _30967_, _30968_, _30969_, _30970_, _30971_, _30972_, _30973_, _30974_, _30975_, _30976_, _30977_, _30978_, _30979_, _30980_, _30981_, _30982_, _30983_, _30984_, _30985_, _30986_, _30987_, _30988_, _30989_, _30990_, _30991_, _30992_, _30993_, _30994_, _30995_, _30996_, _30997_, _30998_, _30999_, _31000_, _31001_, _31002_, _31003_, _31004_, _31005_, _31006_, _31007_, _31008_, _31009_, _31010_, _31011_, _31012_, _31013_, _31014_, _31015_, _31016_, _31017_, _31018_, _31019_, _31020_, _31021_, _31022_, _31023_, _31024_, _31025_, _31026_, _31027_, _31028_, _31029_, _31030_, _31031_, _31032_, _31033_, _31034_, _31035_, _31036_, _31037_, _31038_, _31039_, _31040_, _31041_, _31042_, _31043_, _31044_, _31045_, _31046_, _31047_, _31048_, _31049_, _31050_, _31051_, _31052_, _31053_, _31054_, _31055_, _31056_, _31057_, _31058_, _31059_, _31060_, _31061_, _31062_, _31063_, _31064_, _31065_, _31066_, _31067_, _31068_, _31069_, _31070_, _31071_, _31072_, _31073_, _31074_, _31075_, _31076_, _31077_, _31078_, _31079_, _31080_, _31081_, _31082_, _31083_, _31084_, _31085_, _31086_, _31087_, _31088_, _31089_, _31090_, _31091_, _31092_, _31093_, _31094_, _31095_, _31096_, _31097_, _31098_, _31099_, _31100_, _31101_, _31102_, _31103_, _31104_, _31105_, _31106_, _31107_, _31108_, _31109_, _31110_, _31111_, _31112_, _31113_, _31114_, _31115_, _31116_, _31117_, _31118_, _31119_, _31120_, _31121_, _31122_, _31123_, _31124_, _31125_, _31126_, _31127_, _31128_, _31129_, _31130_, _31131_, _31132_, _31133_, _31134_, _31135_, _31136_, _31137_, _31138_, _31139_, _31140_, _31141_, _31142_, _31143_, _31144_, _31145_, _31146_, _31147_, _31148_, _31149_, _31150_, _31151_, _31152_, _31153_, _31154_, _31155_, _31156_, _31157_, _31158_, _31159_, _31160_, _31161_, _31162_, _31163_, _31164_, _31165_, _31166_, _31167_, _31168_, _31169_, _31170_, _31171_, _31172_, _31173_, _31174_, _31175_, _31176_, _31177_, _31178_, _31179_, _31180_, _31181_, _31182_, _31183_, _31184_, _31185_, _31186_, _31187_, _31188_, _31189_, _31190_, _31191_, _31192_, _31193_, _31194_, _31195_, _31196_, _31197_, _31198_, _31199_, _31200_, _31201_, _31202_, _31203_, _31204_, _31205_, _31206_, _31207_, _31208_, _31209_, _31210_, _31211_, _31212_, _31213_, _31214_, _31215_, _31216_, _31217_, _31218_, _31219_, _31220_, _31221_, _31222_, _31223_, _31224_, _31225_, _31226_, _31227_, _31228_, _31229_, _31230_, _31231_, _31232_, _31233_, _31234_, _31235_, _31236_, _31237_, _31238_, _31239_, _31240_, _31241_, _31242_, _31243_, _31244_, _31245_, _31246_, _31247_, _31248_, _31249_, _31250_, _31251_, _31252_, _31253_, _31254_, _31255_, _31256_, _31257_, _31258_, _31259_, _31260_, _31261_, _31262_, _31263_, _31264_, _31265_, _31266_, _31267_, _31268_, _31269_, _31270_, _31271_, _31272_, _31273_, _31274_, _31275_, _31276_, _31277_, _31278_, _31279_, _31280_, _31281_, _31282_, _31283_, _31284_, _31285_, _31286_, _31287_, _31288_, _31289_, _31290_, _31291_, _31292_, _31293_, _31294_, _31295_, _31296_, _31297_, _31298_, _31299_, _31300_, _31301_, _31302_, _31303_, _31304_, _31305_, _31306_, _31307_, _31308_, _31309_, _31310_, _31311_, _31312_, _31313_, _31314_, _31315_, _31316_, _31317_, _31318_, _31319_, _31320_, _31321_, _31322_, _31323_, _31324_, _31325_, _31326_, _31327_, _31328_, _31329_, _31330_, _31331_, _31332_, _31333_, _31334_, _31335_, _31336_, _31337_, _31338_, _31339_, _31340_, _31341_, _31342_, _31343_, _31344_, _31345_, _31346_, _31347_, _31348_, _31349_, _31350_, _31351_, _31352_, _31353_, _31354_, _31355_, _31356_, _31357_, _31358_, _31359_, _31360_, _31361_, _31362_, _31363_, _31364_, _31365_, _31366_, _31367_, _31368_, _31369_, _31370_, _31371_, _31372_, _31373_, _31374_, _31375_, _31376_, _31377_, _31378_, _31379_, _31380_, _31381_, _31382_, _31383_, _31384_, _31385_, _31386_, _31387_, _31388_, _31389_, _31390_, _31391_, _31392_, _31393_, _31394_, _31395_, _31396_, _31397_, _31398_, _31399_, _31400_, _31401_, _31402_, _31403_, _31404_, _31405_, _31406_, _31407_, _31408_, _31409_, _31410_, _31411_, _31412_, _31413_, _31414_, _31415_, _31416_, _31417_, _31418_, _31419_, _31420_, _31421_, _31422_, _31423_, _31424_, _31425_, _31426_, _31427_, _31428_, _31429_, _31430_, _31431_, _31432_, _31433_, _31434_, _31435_, _31436_, _31437_, _31438_, _31439_, _31440_, _31441_, _31442_, _31443_, _31444_, _31445_, _31446_, _31447_, _31448_, _31449_, _31450_, _31451_, _31452_, _31453_, _31454_, _31455_, _31456_, _31457_, _31458_, _31459_, _31460_, _31461_, _31462_, _31463_, _31464_, _31465_, _31466_, _31467_, _31468_, _31469_, _31470_, _31471_, _31472_, _31473_, _31474_, _31475_, _31476_, _31477_, _31478_, _31479_, _31480_, _31481_, _31482_, _31483_, _31484_, _31485_, _31486_, _31487_, _31488_, _31489_, _31490_, _31491_, _31492_, _31493_, _31494_, _31495_, _31496_, _31497_, _31498_, _31499_, _31500_, _31501_, _31502_, _31503_, _31504_, _31505_, _31506_, _31507_, _31508_, _31509_, _31510_, _31511_, _31512_, _31513_, _31514_, _31515_, _31516_, _31517_, _31518_, _31519_, _31520_, _31521_, _31522_, _31523_, _31524_, _31525_, _31526_, _31527_, _31528_, _31529_, _31530_, _31531_, _31532_, _31533_, _31534_, _31535_, _31536_, _31537_, _31538_, _31539_, _31540_, _31541_, _31542_, _31543_, _31544_, _31545_, _31546_, _31547_, _31548_, _31549_, _31550_, _31551_, _31552_, _31553_, _31554_, _31555_, _31556_, _31557_, _31558_, _31559_, _31560_, _31561_, _31562_, _31563_, _31564_, _31565_, _31566_, _31567_, _31568_, _31569_, _31570_, _31571_, _31572_, _31573_, _31574_, _31575_, _31576_, _31577_, _31578_, _31579_, _31580_, _31581_, _31582_, _31583_, _31584_, _31585_, _31586_, _31587_, _31588_, _31589_, _31590_, _31591_, _31592_, _31593_, _31594_, _31595_, _31596_, _31597_, _31598_, _31599_, _31600_, _31601_, _31602_, _31603_, _31604_, _31605_, _31606_, _31607_, _31608_, _31609_, _31610_, _31611_, _31612_, _31613_, _31614_, _31615_, _31616_, _31617_, _31618_, _31619_, _31620_, _31621_, _31622_, _31623_, _31624_, _31625_, _31626_, _31627_, _31628_, _31629_, _31630_, _31631_, _31632_, _31633_, _31634_, _31635_, _31636_, _31637_, _31638_, _31639_, _31640_, _31641_, _31642_, _31643_, _31644_, _31645_, _31646_, _31647_, _31648_, _31649_, _31650_, _31651_, _31652_, _31653_, _31654_, _31655_, _31656_, _31657_, _31658_, _31659_, _31660_, _31661_, _31662_, _31663_, _31664_, _31665_, _31666_, _31667_, _31668_, _31669_, _31670_, _31671_, _31672_, _31673_, _31674_, _31675_, _31676_, _31677_, _31678_, _31679_, _31680_, _31681_, _31682_, _31683_, _31684_, _31685_, _31686_, _31687_, _31688_, _31689_, _31690_, _31691_, _31692_, _31693_, _31694_, _31695_, _31696_, _31697_, _31698_, _31699_, _31700_, _31701_, _31702_, _31703_, _31704_, _31705_, _31706_, _31707_, _31708_, _31709_, _31710_, _31711_, _31712_, _31713_, _31714_, _31715_, _31716_, _31717_, _31718_, _31719_, _31720_, _31721_, _31722_, _31723_, _31724_, _31725_, _31726_, _31727_, _31728_, _31729_, _31730_, _31731_, _31732_, _31733_, _31734_, _31735_, _31736_, _31737_, _31738_, _31739_, _31740_, _31741_, _31742_, _31743_, _31744_, _31745_, _31746_, _31747_, _31748_, _31749_, _31750_, _31751_, _31752_, _31753_, _31754_, _31755_, _31756_, _31757_, _31758_, _31759_, _31760_, _31761_, _31762_, _31763_, _31764_, _31765_, _31766_, _31767_, _31768_, _31769_, _31770_, _31771_, _31772_, _31773_, _31774_, _31775_, _31776_, _31777_, _31778_, _31779_, _31780_, _31781_, _31782_, _31783_, _31784_, _31785_, _31786_, _31787_, _31788_, _31789_, _31790_, _31791_, _31792_, _31793_, _31794_, _31795_, _31796_, _31797_, _31798_, _31799_, _31800_, _31801_, _31802_, _31803_, _31804_, _31805_, _31806_, _31807_, _31808_, _31809_, _31810_, _31811_, _31812_, _31813_, _31814_, _31815_, _31816_, _31817_, _31818_, _31819_, _31820_, _31821_, _31822_, _31823_, _31824_, _31825_, _31826_, _31827_, _31828_, _31829_, _31830_, _31831_, _31832_, _31833_, _31834_, _31835_, _31836_, _31837_, _31838_, _31839_, _31840_, _31841_, _31842_, _31843_, _31844_, _31845_, _31846_, _31847_, _31848_, _31849_, _31850_, _31851_, _31852_, _31853_, _31854_, _31855_, _31856_, _31857_, _31858_, _31859_, _31860_, _31861_, _31862_, _31863_, _31864_, _31865_, _31866_, _31867_, _31868_, _31869_, _31870_, _31871_, _31872_, _31873_, _31874_, _31875_, _31876_, _31877_, _31878_, _31879_, _31880_, _31881_, _31882_, _31883_, _31884_, _31885_, _31886_, _31887_, _31888_, _31889_, _31890_, _31891_, _31892_, _31893_, _31894_, _31895_, _31896_, _31897_, _31898_, _31899_, _31900_, _31901_, _31902_, _31903_, _31904_, _31905_, _31906_, _31907_, _31908_, _31909_, _31910_, _31911_, _31912_, _31913_, _31914_, _31915_, _31916_, _31917_, _31918_, _31919_, _31920_, _31921_, _31922_, _31923_, _31924_, _31925_, _31926_, _31927_, _31928_, _31929_, _31930_, _31931_, _31932_, _31933_, _31934_, _31935_, _31936_, _31937_, _31938_, _31939_, _31940_, _31941_, _31942_, _31943_, _31944_, _31945_, _31946_, _31947_, _31948_, _31949_, _31950_, _31951_, _31952_, _31953_, _31954_, _31955_, _31956_, _31957_, _31958_, _31959_, _31960_, _31961_, _31962_, _31963_, _31964_, _31965_, _31966_, _31967_, _31968_, _31969_, _31970_, _31971_, _31972_, _31973_, _31974_, _31975_, _31976_, _31977_, _31978_, _31979_, _31980_, _31981_, _31982_, _31983_, _31984_, _31985_, _31986_, _31987_, _31988_, _31989_, _31990_, _31991_, _31992_, _31993_, _31994_, _31995_, _31996_, _31997_, _31998_, _31999_, _32000_, _32001_, _32002_, _32003_, _32004_, _32005_, _32006_, _32007_, _32008_, _32009_, _32010_, _32011_, _32012_, _32013_, _32014_, _32015_, _32016_, _32017_, _32018_, _32019_, _32020_, _32021_, _32022_, _32023_, _32024_, _32025_, _32026_, _32027_, _32028_, _32029_, _32030_, _32031_, _32032_, _32033_, _32034_, _32035_, _32036_, _32037_, _32038_, _32039_, _32040_, _32041_, _32042_, _32043_, _32044_, _32045_, _32046_, _32047_, _32048_, _32049_, _32050_, _32051_, _32052_, _32053_, _32054_, _32055_, _32056_, _32057_, _32058_, _32059_, _32060_, _32061_, _32062_, _32063_, _32064_, _32065_, _32066_, _32067_, _32068_, _32069_, _32070_, _32071_, _32072_, _32073_, _32074_, _32075_, _32076_, _32077_, _32078_, _32079_, _32080_, _32081_, _32082_, _32083_, _32084_, _32085_, _32086_, _32087_, _32088_, _32089_, _32090_, _32091_, _32092_, _32093_, _32094_, _32095_, _32096_, _32097_, _32098_, _32099_, _32100_, _32101_, _32102_, _32103_, _32104_, _32105_, _32106_, _32107_, _32108_, _32109_, _32110_, _32111_, _32112_, _32113_, _32114_, _32115_, _32116_, _32117_, _32118_, _32119_, _32120_, _32121_, _32122_, _32123_, _32124_, _32125_, _32126_, _32127_, _32128_, _32129_, _32130_, _32131_, _32132_, _32133_, _32134_, _32135_, _32136_, _32137_, _32138_, _32139_, _32140_, _32141_, _32142_, _32143_, _32144_, _32145_, _32146_, _32147_, _32148_, _32149_, _32150_, _32151_, _32152_, _32153_, _32154_, _32155_, _32156_, _32157_, _32158_, _32159_, _32160_, _32161_, _32162_, _32163_, _32164_, _32165_, _32166_, _32167_, _32168_, _32169_, _32170_, _32171_, _32172_, _32173_, _32174_, _32175_, _32176_, _32177_, _32178_, _32179_, _32180_, _32181_, _32182_, _32183_, _32184_, _32185_, _32186_, _32187_, _32188_, _32189_, _32190_, _32191_, _32192_, _32193_, _32194_, _32195_, _32196_, _32197_, _32198_, _32199_, _32200_, _32201_, _32202_, _32203_, _32204_, _32205_, _32206_, _32207_, _32208_, _32209_, _32210_, _32211_, _32212_, _32213_, _32214_, _32215_, _32216_, _32217_, _32218_, _32219_, _32220_, _32221_, _32222_, _32223_, _32224_, _32225_, _32226_, _32227_, _32228_, _32229_, _32230_, _32231_, _32232_, _32233_, _32234_, _32235_, _32236_, _32237_, _32238_, _32239_, _32240_, _32241_, _32242_, _32243_, _32244_, _32245_, _32246_, _32247_, _32248_, _32249_, _32250_, _32251_, _32252_, _32253_, _32254_, _32255_, _32256_, _32257_, _32258_, _32259_, _32260_, _32261_, _32262_, _32263_, _32264_, _32265_, _32266_, _32267_, _32268_, _32269_, _32270_, _32271_, _32272_, _32273_, _32274_, _32275_, _32276_, _32277_, _32278_, _32279_, _32280_, _32281_, _32282_, _32283_, _32284_, _32285_, _32286_, _32287_, _32288_, _32289_, _32290_, _32291_, _32292_, _32293_, _32294_, _32295_, _32296_, _32297_, _32298_, _32299_, _32300_, _32301_, _32302_, _32303_, _32304_, _32305_, _32306_, _32307_, _32308_, _32309_, _32310_, _32311_, _32312_, _32313_, _32314_, _32315_, _32316_, _32317_, _32318_, _32319_, _32320_, _32321_, _32322_, _32323_, _32324_, _32325_, _32326_, _32327_, _32328_, _32329_, _32330_, _32331_, _32332_, _32333_, _32334_, _32335_, _32336_, _32337_, _32338_, _32339_, _32340_, _32341_, _32342_, _32343_, _32344_, _32345_, _32346_, _32347_, _32348_, _32349_, _32350_, _32351_, _32352_, _32353_, _32354_, _32355_, _32356_, _32357_, _32358_, _32359_, _32360_, _32361_, _32362_, _32363_, _32364_, _32365_, _32366_, _32367_, _32368_, _32369_, _32370_, _32371_, _32372_, _32373_, _32374_, _32375_, _32376_, _32377_, _32378_, _32379_, _32380_, _32381_, _32382_, _32383_, _32384_, _32385_, _32386_, _32387_, _32388_, _32389_, _32390_, _32391_, _32392_, _32393_, _32394_, _32395_, _32396_, _32397_, _32398_, _32399_, _32400_, _32401_, _32402_, _32403_, _32404_, _32405_, _32406_, _32407_, _32408_, _32409_, _32410_, _32411_, _32412_, _32413_, _32414_, _32415_, _32416_, _32417_, _32418_, _32419_, _32420_, _32421_, _32422_, _32423_, _32424_, _32425_, _32426_, _32427_, _32428_, _32429_, _32430_, _32431_, _32432_, _32433_, _32434_, _32435_, _32436_, _32437_, _32438_, _32439_, _32440_, _32441_, _32442_, _32443_, _32444_, _32445_, _32446_, _32447_, _32448_, _32449_, _32450_, _32451_, _32452_, _32453_, _32454_, _32455_, _32456_, _32457_, _32458_, _32459_, _32460_, _32461_, _32462_, _32463_, _32464_, _32465_, _32466_, _32467_, _32468_, _32469_, _32470_, _32471_, _32472_, _32473_, _32474_, _32475_, _32476_, _32477_, _32478_, _32479_, _32480_, _32481_, _32482_, _32483_, _32484_, _32485_, _32486_, _32487_, _32488_, _32489_, _32490_, _32491_, _32492_, _32493_, _32494_, _32495_, _32496_, _32497_, _32498_, _32499_, _32500_, _32501_, _32502_, _32503_, _32504_, _32505_, _32506_, _32507_, _32508_, _32509_, _32510_, _32511_, _32512_, _32513_, _32514_, _32515_, _32516_, _32517_, _32518_, _32519_, _32520_, _32521_, _32522_, _32523_, _32524_, _32525_, _32526_, _32527_, _32528_, _32529_, _32530_, _32531_, _32532_, _32533_, _32534_, _32535_, _32536_, _32537_, _32538_, _32539_, _32540_, _32541_, _32542_, _32543_, _32544_, _32545_, _32546_, _32547_, _32548_, _32549_, _32550_, _32551_, _32552_, _32553_, _32554_, _32555_, _32556_, _32557_, _32558_, _32559_, _32560_, _32561_, _32562_, _32563_, _32564_, _32565_, _32566_, _32567_, _32568_, _32569_, _32570_, _32571_, _32572_, _32573_, _32574_, _32575_, _32576_, _32577_, _32578_, _32579_, _32580_, _32581_, _32582_, _32583_, _32584_, _32585_, _32586_, _32587_, _32588_, _32589_, _32590_, _32591_, _32592_, _32593_, _32594_, _32595_, _32596_, _32597_, _32598_, _32599_, _32600_, _32601_, _32602_, _32603_, _32604_, _32605_, _32606_, _32607_, _32608_, _32609_, _32610_, _32611_, _32612_, _32613_, _32614_, _32615_, _32616_, _32617_, _32618_, _32619_, _32620_, _32621_, _32622_, _32623_, _32624_, _32625_, _32626_, _32627_, _32628_, _32629_, _32630_, _32631_, _32632_, _32633_, _32634_, _32635_, _32636_, _32637_, _32638_, _32639_, _32640_, _32641_, _32642_, _32643_, _32644_, _32645_, _32646_, _32647_, _32648_, _32649_, _32650_, _32651_, _32652_, _32653_, _32654_, _32655_, _32656_, _32657_, _32658_, _32659_, _32660_, _32661_, _32662_, _32663_, _32664_, _32665_, _32666_, _32667_, _32668_, _32669_, _32670_, _32671_, _32672_, _32673_, _32674_, _32675_, _32676_, _32677_, _32678_, _32679_, _32680_, _32681_, _32682_, _32683_, _32684_, _32685_, _32686_, _32687_, _32688_, _32689_, _32690_, _32691_, _32692_, _32693_, _32694_, _32695_, _32696_, _32697_, _32698_, _32699_, _32700_, _32701_, _32702_, _32703_, _32704_, _32705_, _32706_, _32707_, _32708_, _32709_, _32710_, _32711_, _32712_, _32713_, _32714_, _32715_, _32716_, _32717_, _32718_, _32719_, _32720_, _32721_, _32722_, _32723_, _32724_, _32725_, _32726_, _32727_, _32728_, _32729_, _32730_, _32731_, _32732_, _32733_, _32734_, _32735_, _32736_, _32737_, _32738_, _32739_, _32740_, _32741_, _32742_, _32743_, _32744_, _32745_, _32746_, _32747_, _32748_, _32749_, _32750_, _32751_, _32752_, _32753_, _32754_, _32755_, _32756_, _32757_, _32758_, _32759_, _32760_, _32761_, _32762_, _32763_, _32764_, _32765_, _32766_, _32767_, _32768_, _32769_, _32770_, _32771_, _32772_, _32773_, _32774_, _32775_, _32776_, _32777_, _32778_, _32779_, _32780_, _32781_, _32782_, _32783_, _32784_, _32785_, _32786_, _32787_, _32788_, _32789_, _32790_, _32791_, _32792_, _32793_, _32794_, _32795_, _32796_, _32797_, _32798_, _32799_, _32800_, _32801_, _32802_, _32803_, _32804_, _32805_, _32806_, _32807_, _32808_, _32809_, _32810_, _32811_, _32812_, _32813_, _32814_, _32815_, _32816_, _32817_, _32818_, _32819_, _32820_, _32821_, _32822_, _32823_, _32824_, _32825_, _32826_, _32827_, _32828_, _32829_, _32830_, _32831_, _32832_, _32833_, _32834_, _32835_, _32836_, _32837_, _32838_, _32839_, _32840_, _32841_, _32842_, _32843_, _32844_, _32845_, _32846_, _32847_, _32848_, _32849_, _32850_, _32851_, _32852_, _32853_, _32854_, _32855_, _32856_, _32857_, _32858_, _32859_, _32860_, _32861_, _32862_, _32863_, _32864_, _32865_, _32866_, _32867_, _32868_, _32869_, _32870_, _32871_, _32872_, _32873_, _32874_, _32875_, _32876_, _32877_, _32878_, _32879_, _32880_, _32881_, _32882_, _32883_, _32884_, _32885_, _32886_, _32887_, _32888_, _32889_, _32890_, _32891_, _32892_, _32893_, _32894_, _32895_, _32896_, _32897_, _32898_, _32899_, _32900_, _32901_, _32902_, _32903_, _32904_, _32905_, _32906_, _32907_, _32908_, _32909_, _32910_, _32911_, _32912_, _32913_, _32914_, _32915_, _32916_, _32917_, _32918_, _32919_, _32920_, _32921_, _32922_, _32923_, _32924_, _32925_, _32926_, _32927_, _32928_, _32929_, _32930_, _32931_, _32932_, _32933_, _32934_, _32935_, _32936_, _32937_, _32938_, _32939_, _32940_, _32941_, _32942_, _32943_, _32944_, _32945_, _32946_, _32947_, _32948_, _32949_, _32950_, _32951_, _32952_, _32953_, _32954_, _32955_, _32956_, _32957_, _32958_, _32959_, _32960_, _32961_, _32962_, _32963_, _32964_, _32965_, _32966_, _32967_, _32968_, _32969_, _32970_, _32971_, _32972_, _32973_, _32974_, _32975_, _32976_, _32977_, _32978_, _32979_, _32980_, _32981_, _32982_, _32983_, _32984_, _32985_, _32986_, _32987_, _32988_, _32989_, _32990_, _32991_, _32992_, _32993_, _32994_, _32995_, _32996_, _32997_, _32998_, _32999_, _33000_, _33001_, _33002_, _33003_, _33004_, _33005_, _33006_, _33007_, _33008_, _33009_, _33010_, _33011_, _33012_, _33013_, _33014_, _33015_, _33016_, _33017_, _33018_, _33019_, _33020_, _33021_, _33022_, _33023_, _33024_, _33025_, _33026_, _33027_, _33028_, _33029_, _33030_, _33031_, _33032_, _33033_, _33034_, _33035_, _33036_, _33037_, _33038_, _33039_, _33040_, _33041_, _33042_, _33043_, _33044_, _33045_, _33046_, _33047_, _33048_, _33049_, _33050_, _33051_, _33052_, _33053_, _33054_, _33055_, _33056_, _33057_, _33058_, _33059_, _33060_, _33061_, _33062_, _33063_, _33064_, _33065_, _33066_, _33067_, _33068_, _33069_, _33070_, _33071_, _33072_, _33073_, _33074_, _33075_, _33076_, _33077_, _33078_, _33079_, _33080_, _33081_, _33082_, _33083_, _33084_, _33085_, _33086_, _33087_, _33088_, _33089_, _33090_, _33091_, _33092_, _33093_, _33094_, _33095_, _33096_, _33097_, _33098_, _33099_, _33100_, _33101_, _33102_, _33103_, _33104_, _33105_, _33106_, _33107_, _33108_, _33109_, _33110_, _33111_, _33112_, _33113_, _33114_, _33115_, _33116_, _33117_, _33118_, _33119_, _33120_, _33121_, _33122_, _33123_, _33124_, _33125_, _33126_, _33127_, _33128_, _33129_, _33130_, _33131_, _33132_, _33133_, _33134_, _33135_, _33136_, _33137_, _33138_, _33139_, _33140_, _33141_, _33142_, _33143_, _33144_, _33145_, _33146_, _33147_, _33148_, _33149_, _33150_, _33151_, _33152_, _33153_, _33154_, _33155_, _33156_, _33157_, _33158_, _33159_, _33160_, _33161_, _33162_, _33163_, _33164_, _33165_, _33166_, _33167_, _33168_, _33169_, _33170_, _33171_, _33172_, _33173_, _33174_, _33175_, _33176_, _33177_, _33178_, _33179_, _33180_, _33181_, _33182_, _33183_, _33184_, _33185_, _33186_, _33187_, _33188_, _33189_, _33190_, _33191_, _33192_, _33193_, _33194_, _33195_, _33196_, _33197_, _33198_, _33199_, _33200_, _33201_, _33202_, _33203_, _33204_, _33205_, _33206_, _33207_, _33208_, _33209_, _33210_, _33211_, _33212_, _33213_, _33214_, _33215_, _33216_, _33217_, _33218_, _33219_, _33220_, _33221_, _33222_, _33223_, _33224_, _33225_, _33226_, _33227_, _33228_, _33229_, _33230_, _33231_, _33232_, _33233_, _33234_, _33235_, _33236_, _33237_, _33238_, _33239_, _33240_, _33241_, _33242_, _33243_, _33244_, _33245_, _33246_, _33247_, _33248_, _33249_, _33250_, _33251_, _33252_, _33253_, _33254_, _33255_, _33256_, _33257_, _33258_, _33259_, _33260_, _33261_, _33262_, _33263_, _33264_, _33265_, _33266_, _33267_, _33268_, _33269_, _33270_, _33271_, _33272_, _33273_, _33274_, _33275_, _33276_, _33277_, _33278_, _33279_, _33280_, _33281_, _33282_, _33283_, _33284_, _33285_, _33286_, _33287_, _33288_, _33289_, _33290_, _33291_, _33292_, _33293_, _33294_, _33295_, _33296_, _33297_, _33298_, _33299_, _33300_, _33301_, _33302_, _33303_, _33304_, _33305_, _33306_, _33307_, _33308_, _33309_, _33310_, _33311_, _33312_, _33313_, _33314_, _33315_, _33316_, _33317_, _33318_, _33319_, _33320_, _33321_, _33322_, _33323_, _33324_, _33325_, _33326_, _33327_, _33328_, _33329_, _33330_, _33331_, _33332_, _33333_, _33334_, _33335_, _33336_, _33337_, _33338_, _33339_, _33340_, _33341_, _33342_, _33343_, _33344_, _33345_, _33346_, _33347_, _33348_, _33349_, _33350_, _33351_, _33352_, _33353_, _33354_, _33355_, _33356_, _33357_, _33358_, _33359_, _33360_, _33361_, _33362_, _33363_, _33364_, _33365_, _33366_, _33367_, _33368_, _33369_, _33370_, _33371_, _33372_, _33373_, _33374_, _33375_, _33376_, _33377_, _33378_, _33379_, _33380_, _33381_, _33382_, _33383_, _33384_, _33385_, _33386_, _33387_, _33388_, _33389_, _33390_, _33391_, _33392_, _33393_, _33394_, _33395_, _33396_, _33397_, _33398_, _33399_, _33400_, _33401_, _33402_, _33403_, _33404_, _33405_, _33406_, _33407_, _33408_, _33409_, _33410_, _33411_, _33412_, _33413_, _33414_, _33415_, _33416_, _33417_, _33418_, _33419_, _33420_, _33421_, _33422_, _33423_, _33424_, _33425_, _33426_, _33427_, _33428_, _33429_, _33430_, _33431_, _33432_, _33433_, _33434_, _33435_, _33436_, _33437_, _33438_, _33439_, _33440_, _33441_, _33442_, _33443_, _33444_, _33445_, _33446_, _33447_, _33448_, _33449_, _33450_, _33451_, _33452_, _33453_, _33454_, _33455_, _33456_, _33457_, _33458_, _33459_, _33460_, _33461_, _33462_, _33463_, _33464_, _33465_, _33466_, _33467_, _33468_, _33469_, _33470_, _33471_, _33472_, _33473_, _33474_, _33475_, _33476_, _33477_, _33478_, _33479_, _33480_, _33481_, _33482_, _33483_, _33484_, _33485_, _33486_, _33487_, _33488_, _33489_, _33490_, _33491_, _33492_, _33493_, _33494_, _33495_, _33496_, _33497_, _33498_, _33499_, _33500_, _33501_, _33502_, _33503_, _33504_, _33505_, _33506_, _33507_, _33508_, _33509_, _33510_, _33511_, _33512_, _33513_, _33514_, _33515_, _33516_, _33517_, _33518_, _33519_, _33520_, _33521_, _33522_, _33523_, _33524_, _33525_, _33526_, _33527_, _33528_, _33529_, _33530_, _33531_, _33532_, _33533_, _33534_, _33535_, _33536_, _33537_, _33538_, _33539_, _33540_, _33541_, _33542_, _33543_, _33544_, _33545_, _33546_, _33547_, _33548_, _33549_, _33550_, _33551_, _33552_, _33553_, _33554_, _33555_, _33556_, _33557_, _33558_, _33559_, _33560_, _33561_, _33562_, _33563_, _33564_, _33565_, _33566_, _33567_, _33568_, _33569_, _33570_, _33571_, _33572_, _33573_, _33574_, _33575_, _33576_, _33577_, _33578_, _33579_, _33580_, _33581_, _33582_, _33583_, _33584_, _33585_, _33586_, _33587_, _33588_, _33589_, _33590_, _33591_, _33592_, _33593_, _33594_, _33595_, _33596_, _33597_, _33598_, _33599_, _33600_, _33601_, _33602_, _33603_, _33604_, _33605_, _33606_, _33607_, _33608_, _33609_, _33610_, _33611_, _33612_, _33613_, _33614_, _33615_, _33616_, _33617_, _33618_, _33619_, _33620_, _33621_, _33622_, _33623_, _33624_, _33625_, _33626_, _33627_, _33628_, _33629_, _33630_, _33631_, _33632_, _33633_, _33634_, _33635_, _33636_, _33637_, _33638_, _33639_, _33640_, _33641_, _33642_, _33643_, _33644_, _33645_, _33646_, _33647_, _33648_, _33649_, _33650_, _33651_, _33652_, _33653_, _33654_, _33655_, _33656_, _33657_, _33658_, _33659_, _33660_, _33661_, _33662_, _33663_, _33664_, _33665_, _33666_, _33667_, _33668_, _33669_, _33670_, _33671_, _33672_, _33673_, _33674_, _33675_, _33676_, _33677_, _33678_, _33679_, _33680_, _33681_, _33682_, _33683_, _33684_, _33685_, _33686_, _33687_, _33688_, _33689_, _33690_, _33691_, _33692_, _33693_, _33694_, _33695_, _33696_, _33697_, _33698_, _33699_, _33700_, _33701_, _33702_, _33703_, _33704_, _33705_, _33706_, _33707_, _33708_, _33709_, _33710_, _33711_, _33712_, _33713_, _33714_, _33715_, _33716_, _33717_, _33718_, _33719_, _33720_, _33721_, _33722_, _33723_, _33724_, _33725_, _33726_, _33727_, _33728_, _33729_, _33730_, _33731_, _33732_, _33733_, _33734_, _33735_, _33736_, _33737_, _33738_, _33739_, _33740_, _33741_, _33742_, _33743_, _33744_, _33745_, _33746_, _33747_, _33748_, _33749_, _33750_, _33751_, _33752_, _33753_, _33754_, _33755_, _33756_, _33757_, _33758_, _33759_, _33760_, _33761_, _33762_, _33763_, _33764_, _33765_, _33766_, _33767_, _33768_, _33769_, _33770_, _33771_, _33772_, _33773_, _33774_, _33775_, _33776_, _33777_, _33778_, _33779_, _33780_, _33781_, _33782_, _33783_, _33784_, _33785_, _33786_, _33787_, _33788_, _33789_, _33790_, _33791_, _33792_, _33793_, _33794_, _33795_, _33796_, _33797_, _33798_, _33799_, _33800_, _33801_, _33802_, _33803_, _33804_, _33805_, _33806_, _33807_, _33808_, _33809_, _33810_, _33811_, _33812_, _33813_, _33814_, _33815_, _33816_, _33817_, _33818_, _33819_, _33820_, _33821_, _33822_, _33823_, _33824_, _33825_, _33826_, _33827_, _33828_, _33829_, _33830_, _33831_, _33832_, _33833_, _33834_, _33835_, _33836_, _33837_, _33838_, _33839_, _33840_, _33841_, _33842_, _33843_, _33844_, _33845_, _33846_, _33847_, _33848_, _33849_, _33850_, _33851_, _33852_, _33853_, _33854_, _33855_, _33856_, _33857_, _33858_, _33859_, _33860_, _33861_, _33862_, _33863_, _33864_, _33865_, _33866_, _33867_, _33868_, _33869_, _33870_, _33871_, _33872_, _33873_, _33874_, _33875_, _33876_, _33877_, _33878_, _33879_, _33880_, _33881_, _33882_, _33883_, _33884_, _33885_, _33886_, _33887_, _33888_, _33889_, _33890_, _33891_, _33892_, _33893_, _33894_, _33895_, _33896_, _33897_, _33898_, _33899_, _33900_, _33901_, _33902_, _33903_, _33904_, _33905_, _33906_, _33907_, _33908_, _33909_, _33910_, _33911_, _33912_, _33913_, _33914_, _33915_, _33916_, _33917_, _33918_, _33919_, _33920_, _33921_, _33922_, _33923_, _33924_, _33925_, _33926_, _33927_, _33928_, _33929_, _33930_, _33931_, _33932_, _33933_, _33934_, _33935_, _33936_, _33937_, _33938_, _33939_, _33940_, _33941_, _33942_, _33943_, _33944_, _33945_, _33946_, _33947_, _33948_, _33949_, _33950_, _33951_, _33952_, _33953_, _33954_, _33955_, _33956_, _33957_, _33958_, _33959_, _33960_, _33961_, _33962_, _33963_, _33964_, _33965_, _33966_, _33967_, _33968_, _33969_, _33970_, _33971_, _33972_, _33973_, _33974_, _33975_, _33976_, _33977_, _33978_, _33979_, _33980_, _33981_, _33982_, _33983_, _33984_, _33985_, _33986_, _33987_, _33988_, _33989_, _33990_, _33991_, _33992_, _33993_, _33994_, _33995_, _33996_, _33997_, _33998_, _33999_, _34000_, _34001_, _34002_, _34003_, _34004_, _34005_, _34006_, _34007_, _34008_, _34009_, _34010_, _34011_, _34012_, _34013_, _34014_, _34015_, _34016_, _34017_, _34018_, _34019_, _34020_, _34021_, _34022_, _34023_, _34024_, _34025_, _34026_, _34027_, _34028_, _34029_, _34030_, _34031_, _34032_, _34033_, _34034_, _34035_, _34036_, _34037_, _34038_, _34039_, _34040_, _34041_, _34042_, _34043_, _34044_, _34045_, _34046_, _34047_, _34048_, _34049_, _34050_, _34051_, _34052_, _34053_, _34054_, _34055_, _34056_, _34057_, _34058_, _34059_, _34060_, _34061_, _34062_, _34063_, _34064_, _34065_, _34066_, _34067_, _34068_, _34069_, _34070_, _34071_, _34072_, _34073_, _34074_, _34075_, _34076_, _34077_, _34078_, _34079_, _34080_, _34081_, _34082_, _34083_, _34084_, _34085_, _34086_, _34087_, _34088_, _34089_, _34090_, _34091_, _34092_, _34093_, _34094_, _34095_, _34096_, _34097_, _34098_, _34099_, _34100_, _34101_, _34102_, _34103_, _34104_, _34105_, _34106_, _34107_, _34108_, _34109_, _34110_, _34111_, _34112_, _34113_, _34114_, _34115_, _34116_, _34117_, _34118_, _34119_, _34120_, _34121_, _34122_, _34123_, _34124_, _34125_, _34126_, _34127_, _34128_, _34129_, _34130_, _34131_, _34132_, _34133_, _34134_, _34135_, _34136_, _34137_, _34138_, _34139_, _34140_, _34141_, _34142_, _34143_, _34144_, _34145_, _34146_, _34147_, _34148_, _34149_, _34150_, _34151_, _34152_, _34153_, _34154_, _34155_, _34156_, _34157_, _34158_, _34159_, _34160_, _34161_, _34162_, _34163_, _34164_, _34165_, _34166_, _34167_, _34168_, _34169_, _34170_, _34171_, _34172_, _34173_, _34174_, _34175_, _34176_, _34177_, _34178_, _34179_, _34180_, _34181_, _34182_, _34183_, _34184_, _34185_, _34186_, _34187_, _34188_, _34189_, _34190_, _34191_, _34192_, _34193_, _34194_, _34195_, _34196_, _34197_, _34198_, _34199_, _34200_, _34201_, _34202_, _34203_, _34204_, _34205_, _34206_, _34207_, _34208_, _34209_, _34210_, _34211_, _34212_, _34213_, _34214_, _34215_, _34216_, _34217_, _34218_, _34219_, _34220_, _34221_, _34222_, _34223_, _34224_, _34225_, _34226_, _34227_, _34228_, _34229_, _34230_, _34231_, _34232_, _34233_, _34234_, _34235_, _34236_, _34237_, _34238_, _34239_, _34240_, _34241_, _34242_, _34243_, _34244_, _34245_, _34246_, _34247_, _34248_, _34249_, _34250_, _34251_, _34252_, _34253_, _34254_, _34255_, _34256_, _34257_, _34258_, _34259_, _34260_, _34261_, _34262_, _34263_, _34264_, _34265_, _34266_, _34267_, _34268_, _34269_, _34270_, _34271_, _34272_, _34273_, _34274_, _34275_, _34276_, _34277_, _34278_, _34279_, _34280_, _34281_, _34282_, _34283_, _34284_, _34285_, _34286_, _34287_, _34288_, _34289_, _34290_, _34291_, _34292_, _34293_, _34294_, _34295_, _34296_, _34297_, _34298_, _34299_, _34300_, _34301_, _34302_, _34303_, _34304_, _34305_, _34306_, _34307_, _34308_, _34309_, _34310_, _34311_, _34312_, _34313_, _34314_, _34315_, _34316_, _34317_, _34318_, _34319_, _34320_, _34321_, _34322_, _34323_, _34324_, _34325_, _34326_, _34327_, _34328_, _34329_, _34330_, _34331_, _34332_, _34333_, _34334_, _34335_, _34336_, _34337_, _34338_, _34339_, _34340_, _34341_, _34342_, _34343_, _34344_, _34345_, _34346_, _34347_, _34348_, _34349_, _34350_, _34351_, _34352_, _34353_, _34354_, _34355_, _34356_, _34357_, _34358_, _34359_, _34360_, _34361_, _34362_, _34363_, _34364_, _34365_, _34366_, _34367_, _34368_, _34369_, _34370_, _34371_, _34372_, _34373_, _34374_, _34375_, _34376_, _34377_, _34378_, _34379_, _34380_, _34381_, _34382_, _34383_, _34384_, _34385_, _34386_, _34387_, _34388_, _34389_, _34390_, _34391_, _34392_, _34393_, _34394_, _34395_, _34396_, _34397_, _34398_, _34399_, _34400_, _34401_, _34402_, _34403_, _34404_, _34405_, _34406_, _34407_, _34408_, _34409_, _34410_, _34411_, _34412_, _34413_, _34414_, _34415_, _34416_, _34417_, _34418_, _34419_, _34420_, _34421_, _34422_, _34423_, _34424_, _34425_, _34426_, _34427_, _34428_, _34429_, _34430_, _34431_, _34432_, _34433_, _34434_, _34435_, _34436_, _34437_, _34438_, _34439_, _34440_, _34441_, _34442_, _34443_, _34444_, _34445_, _34446_, _34447_, _34448_, _34449_, _34450_, _34451_, _34452_, _34453_, _34454_, _34455_, _34456_, _34457_, _34458_, _34459_, _34460_, _34461_, _34462_, _34463_, _34464_, _34465_, _34466_, _34467_, _34468_, _34469_, _34470_, _34471_, _34472_, _34473_, _34474_, _34475_, _34476_, _34477_, _34478_, _34479_, _34480_, _34481_, _34482_, _34483_, _34484_, _34485_, _34486_, _34487_, _34488_, _34489_, _34490_, _34491_, _34492_, _34493_, _34494_, _34495_, _34496_, _34497_, _34498_, _34499_, _34500_, _34501_, _34502_, _34503_, _34504_, _34505_, _34506_, _34507_, _34508_, _34509_, _34510_, _34511_, _34512_, _34513_, _34514_, _34515_, _34516_, _34517_, _34518_, _34519_, _34520_, _34521_, _34522_, _34523_, _34524_, _34525_, _34526_, _34527_, _34528_, _34529_, _34530_, _34531_, _34532_, _34533_, _34534_, _34535_, _34536_, _34537_, _34538_, _34539_, _34540_, _34541_, _34542_, _34543_, _34544_, _34545_, _34546_, _34547_, _34548_, _34549_, _34550_, _34551_, _34552_, _34553_, _34554_, _34555_, _34556_, _34557_, _34558_, _34559_, _34560_, _34561_, _34562_, _34563_, _34564_, _34565_, _34566_, _34567_, _34568_, _34569_, _34570_, _34571_, _34572_, _34573_, _34574_, _34575_, _34576_, _34577_, _34578_, _34579_, _34580_, _34581_, _34582_, _34583_, _34584_, _34585_, _34586_, _34587_, _34588_, _34589_, _34590_, _34591_, _34592_, _34593_, _34594_, _34595_, _34596_, _34597_, _34598_, _34599_, _34600_, _34601_, _34602_, _34603_, _34604_, _34605_, _34606_, _34607_, _34608_, _34609_, _34610_, _34611_, _34612_, _34613_, _34614_, _34615_, _34616_, _34617_, _34618_, _34619_, _34620_, _34621_, _34622_, _34623_, _34624_, _34625_, _34626_, _34627_, _34628_, _34629_, _34630_, _34631_, _34632_, _34633_, _34634_, _34635_, _34636_, _34637_, _34638_, _34639_, _34640_, _34641_, _34642_, _34643_, _34644_, _34645_, _34646_, _34647_, _34648_, _34649_, _34650_, _34651_, _34652_, _34653_, _34654_, _34655_, _34656_, _34657_, _34658_, _34659_, _34660_, _34661_, _34662_, _34663_, _34664_, _34665_, _34666_, _34667_, _34668_, _34669_, _34670_, _34671_, _34672_, _34673_, _34674_, _34675_, _34676_, _34677_, _34678_, _34679_, _34680_, _34681_, _34682_, _34683_, _34684_, _34685_, _34686_, _34687_, _34688_, _34689_, _34690_, _34691_, _34692_, _34693_, _34694_, _34695_, _34696_, _34697_, _34698_, _34699_, _34700_, _34701_, _34702_, _34703_, _34704_, _34705_, _34706_, _34707_, _34708_, _34709_, _34710_, _34711_, _34712_, _34713_, _34714_, _34715_, _34716_, _34717_, _34718_, _34719_, _34720_, _34721_, _34722_, _34723_, _34724_, _34725_, _34726_, _34727_, _34728_, _34729_, _34730_, _34731_, _34732_, _34733_, _34734_, _34735_, _34736_, _34737_, _34738_, _34739_, _34740_, _34741_, _34742_, _34743_, _34744_, _34745_, _34746_, _34747_, _34748_, _34749_, _34750_, _34751_, _34752_, _34753_, _34754_, _34755_, _34756_, _34757_, _34758_, _34759_, _34760_, _34761_, _34762_, _34763_, _34764_, _34765_, _34766_, _34767_, _34768_, _34769_, _34770_, _34771_, _34772_, _34773_, _34774_, _34775_, _34776_, _34777_, _34778_, _34779_, _34780_, _34781_, _34782_, _34783_, _34784_, _34785_, _34786_, _34787_, _34788_, _34789_, _34790_, _34791_, _34792_, _34793_, _34794_, _34795_, _34796_, _34797_, _34798_, _34799_, _34800_, _34801_, _34802_, _34803_, _34804_, _34805_, _34806_, _34807_, _34808_, _34809_, _34810_, _34811_, _34812_, _34813_, _34814_, _34815_, _34816_, _34817_, _34818_, _34819_, _34820_, _34821_, _34822_, _34823_, _34824_, _34825_, _34826_, _34827_, _34828_, _34829_, _34830_, _34831_, _34832_, _34833_, _34834_, _34835_, _34836_, _34837_, _34838_, _34839_, _34840_, _34841_, _34842_, _34843_, _34844_, _34845_, _34846_, _34847_, _34848_, _34849_, _34850_, _34851_, _34852_, _34853_, _34854_, _34855_, _34856_, _34857_, _34858_, _34859_, _34860_, _34861_, _34862_, _34863_, _34864_, _34865_, _34866_, _34867_, _34868_, _34869_, _34870_, _34871_, _34872_, _34873_, _34874_, _34875_, _34876_, _34877_, _34878_, _34879_, _34880_, _34881_, _34882_, _34883_, _34884_, _34885_, _34886_, _34887_, _34888_, _34889_, _34890_, _34891_, _34892_, _34893_, _34894_, _34895_, _34896_, _34897_, _34898_, _34899_, _34900_, _34901_, _34902_, _34903_, _34904_, _34905_, _34906_, _34907_, _34908_, _34909_, _34910_, _34911_, _34912_, _34913_, _34914_, _34915_, _34916_, _34917_, _34918_, _34919_, _34920_, _34921_, _34922_, _34923_, _34924_, _34925_, _34926_, _34927_, _34928_, _34929_, _34930_, _34931_, _34932_, _34933_, _34934_, _34935_, _34936_, _34937_, _34938_, _34939_, _34940_, _34941_, _34942_, _34943_, _34944_, _34945_, _34946_, _34947_, _34948_, _34949_, _34950_, _34951_, _34952_, _34953_, _34954_, _34955_, _34956_, _34957_, _34958_, _34959_, _34960_, _34961_, _34962_, _34963_, _34964_, _34965_, _34966_, _34967_, _34968_, _34969_, _34970_, _34971_, _34972_, _34973_, _34974_, _34975_, _34976_, _34977_, _34978_, _34979_, _34980_, _34981_, _34982_, _34983_, _34984_, _34985_, _34986_, _34987_, _34988_, _34989_, _34990_, _34991_, _34992_, _34993_, _34994_, _34995_, _34996_, _34997_, _34998_, _34999_, _35000_, _35001_, _35002_, _35003_, _35004_, _35005_, _35006_, _35007_, _35008_, _35009_, _35010_, _35011_, _35012_, _35013_, _35014_, _35015_, _35016_, _35017_, _35018_, _35019_, _35020_, _35021_, _35022_, _35023_, _35024_, _35025_, _35026_, _35027_, _35028_, _35029_, _35030_, _35031_, _35032_, _35033_, _35034_, _35035_, _35036_, _35037_, _35038_, _35039_, _35040_, _35041_, _35042_, _35043_, _35044_, _35045_, _35046_, _35047_, _35048_, _35049_, _35050_, _35051_, _35052_, _35053_, _35054_, _35055_, _35056_, _35057_, _35058_, _35059_, _35060_, _35061_, _35062_, _35063_, _35064_, _35065_, _35066_, _35067_, _35068_, _35069_, _35070_, _35071_, _35072_, _35073_, _35074_, _35075_, _35076_, _35077_, _35078_, _35079_, _35080_, _35081_, _35082_, _35083_, _35084_, _35085_, _35086_, _35087_, _35088_, _35089_, _35090_, _35091_, _35092_, _35093_, _35094_, _35095_, _35096_, _35097_, _35098_, _35099_, _35100_, _35101_, _35102_, _35103_, _35104_, _35105_, _35106_, _35107_, _35108_, _35109_, _35110_, _35111_, _35112_, _35113_, _35114_, _35115_, _35116_, _35117_, _35118_, _35119_, _35120_, _35121_, _35122_, _35123_, _35124_, _35125_, _35126_, _35127_, _35128_, _35129_, _35130_, _35131_, _35132_, _35133_, _35134_, _35135_, _35136_, _35137_, _35138_, _35139_, _35140_, _35141_, _35142_, _35143_, _35144_, _35145_, _35146_, _35147_, _35148_, _35149_, _35150_, _35151_, _35152_, _35153_, _35154_, _35155_, _35156_, _35157_, _35158_, _35159_, _35160_, _35161_, _35162_, _35163_, _35164_, _35165_, _35166_, _35167_, _35168_, _35169_, _35170_, _35171_, _35172_, _35173_, _35174_, _35175_, _35176_, _35177_, _35178_, _35179_, _35180_, _35181_, _35182_, _35183_, _35184_, _35185_, _35186_, _35187_, _35188_, _35189_, _35190_, _35191_, _35192_, _35193_, _35194_, _35195_, _35196_, _35197_, _35198_, _35199_, _35200_, _35201_, _35202_, _35203_, _35204_, _35205_, _35206_, _35207_, _35208_, _35209_, _35210_, _35211_, _35212_, _35213_, _35214_, _35215_, _35216_, _35217_, _35218_, _35219_, _35220_, _35221_, _35222_, _35223_, _35224_, _35225_, _35226_, _35227_, _35228_, _35229_, _35230_, _35231_, _35232_, _35233_, _35234_, _35235_, _35236_, _35237_, _35238_, _35239_, _35240_, _35241_, _35242_, _35243_, _35244_, _35245_, _35246_, _35247_, _35248_, _35249_, _35250_, _35251_, _35252_, _35253_, _35254_, _35255_, _35256_, _35257_, _35258_, _35259_, _35260_, _35261_, _35262_, _35263_, _35264_, _35265_, _35266_, _35267_, _35268_, _35269_, _35270_, _35271_, _35272_, _35273_, _35274_, _35275_, _35276_, _35277_, _35278_, _35279_, _35280_, _35281_, _35282_, _35283_, _35284_, _35285_, _35286_, _35287_, _35288_, _35289_, _35290_, _35291_, _35292_, _35293_, _35294_, _35295_, _35296_, _35297_, _35298_, _35299_, _35300_, _35301_, _35302_, _35303_, _35304_, _35305_, _35306_, _35307_, _35308_, _35309_, _35310_, _35311_, _35312_, _35313_, _35314_, _35315_, _35316_, _35317_, _35318_, _35319_, _35320_, _35321_, _35322_, _35323_, _35324_, _35325_, _35326_, _35327_, _35328_, _35329_, _35330_, _35331_, _35332_, _35333_, _35334_, _35335_, _35336_, _35337_, _35338_, _35339_, _35340_, _35341_, _35342_, _35343_, _35344_, _35345_, _35346_, _35347_, _35348_, _35349_, _35350_, _35351_, _35352_, _35353_, _35354_, _35355_, _35356_, _35357_, _35358_, _35359_, _35360_, _35361_, _35362_, _35363_, _35364_, _35365_, _35366_, _35367_, _35368_, _35369_, _35370_, _35371_, _35372_, _35373_, _35374_, _35375_, _35376_, _35377_, _35378_, _35379_, _35380_, _35381_, _35382_, _35383_, _35384_, _35385_, _35386_, _35387_, _35388_, _35389_, _35390_, _35391_, _35392_, _35393_, _35394_, _35395_, _35396_, _35397_, _35398_, _35399_, _35400_, _35401_, _35402_, _35403_, _35404_, _35405_, _35406_, _35407_, _35408_, _35409_, _35410_, _35411_, _35412_, _35413_, _35414_, _35415_, _35416_, _35417_, _35418_, _35419_, _35420_, _35421_, _35422_, _35423_, _35424_, _35425_, _35426_, _35427_, _35428_, _35429_, _35430_, _35431_, _35432_, _35433_, _35434_, _35435_, _35436_, _35437_, _35438_, _35439_, _35440_, _35441_, _35442_, _35443_, _35444_, _35445_, _35446_, _35447_, _35448_, _35449_, _35450_, _35451_, _35452_, _35453_, _35454_, _35455_, _35456_, _35457_, _35458_, _35459_, _35460_, _35461_, _35462_, _35463_, _35464_, _35465_, _35466_, _35467_, _35468_, _35469_, _35470_, _35471_, _35472_, _35473_, _35474_, _35475_, _35476_, _35477_, _35478_, _35479_, _35480_, _35481_, _35482_, _35483_, _35484_, _35485_, _35486_, _35487_, _35488_, _35489_, _35490_, _35491_, _35492_, _35493_, _35494_, _35495_, _35496_, _35497_, _35498_, _35499_, _35500_, _35501_, _35502_, _35503_, _35504_, _35505_, _35506_, _35507_, _35508_, _35509_, _35510_, _35511_, _35512_, _35513_, _35514_, _35515_, _35516_, _35517_, _35518_, _35519_, _35520_, _35521_, _35522_, _35523_, _35524_, _35525_, _35526_, _35527_, _35528_, _35529_, _35530_, _35531_, _35532_, _35533_, _35534_, _35535_, _35536_, _35537_, _35538_, _35539_, _35540_, _35541_, _35542_, _35543_, _35544_, _35545_, _35546_, _35547_, _35548_, _35549_, _35550_, _35551_, _35552_, _35553_, _35554_, _35555_, _35556_, _35557_, _35558_, _35559_, _35560_, _35561_, _35562_, _35563_, _35564_, _35565_, _35566_, _35567_, _35568_, _35569_, _35570_, _35571_, _35572_, _35573_, _35574_, _35575_, _35576_, _35577_, _35578_, _35579_, _35580_, _35581_, _35582_, _35583_, _35584_, _35585_, _35586_, _35587_, _35588_, _35589_, _35590_, _35591_, _35592_, _35593_, _35594_, _35595_, _35596_, _35597_, _35598_, _35599_, _35600_, _35601_, _35602_, _35603_, _35604_, _35605_, _35606_, _35607_, _35608_, _35609_, _35610_, _35611_, _35612_, _35613_, _35614_, _35615_, _35616_, _35617_, _35618_, _35619_, _35620_, _35621_, _35622_, _35623_, _35624_, _35625_, _35626_, _35627_, _35628_, _35629_, _35630_, _35631_, _35632_, _35633_, _35634_, _35635_, _35636_, _35637_, _35638_, _35639_, _35640_, _35641_, _35642_, _35643_, _35644_, _35645_, _35646_, _35647_, _35648_, _35649_, _35650_, _35651_, _35652_, _35653_, _35654_, _35655_, _35656_, _35657_, _35658_, _35659_, _35660_, _35661_, _35662_, _35663_, _35664_, _35665_, _35666_, _35667_, _35668_, _35669_, _35670_, _35671_, _35672_, _35673_, _35674_, _35675_, _35676_, _35677_, _35678_, _35679_, _35680_, _35681_, _35682_, _35683_, _35684_, _35685_, _35686_, _35687_, _35688_, _35689_, _35690_, _35691_, _35692_, _35693_, _35694_, _35695_, _35696_, _35697_, _35698_, _35699_, _35700_, _35701_, _35702_, _35703_, _35704_, _35705_, _35706_, _35707_, _35708_, _35709_, _35710_, _35711_, _35712_, _35713_, _35714_, _35715_, _35716_, _35717_, _35718_, _35719_, _35720_, _35721_, _35722_, _35723_, _35724_, _35725_, _35726_, _35727_, _35728_, _35729_, _35730_, _35731_, _35732_, _35733_, _35734_, _35735_, _35736_, _35737_, _35738_, _35739_, _35740_, _35741_, _35742_, _35743_, _35744_, _35745_, _35746_, _35747_, _35748_, _35749_, _35750_, _35751_, _35752_, _35753_, _35754_, _35755_, _35756_, _35757_, _35758_, _35759_, _35760_, _35761_, _35762_, _35763_, _35764_, _35765_, _35766_, _35767_, _35768_, _35769_, _35770_, _35771_, _35772_, _35773_, _35774_, _35775_, _35776_, _35777_, _35778_, _35779_, _35780_, _35781_, _35782_, _35783_, _35784_, _35785_, _35786_, _35787_, _35788_, _35789_, _35790_, _35791_, _35792_, _35793_, _35794_, _35795_, _35796_, _35797_, _35798_, _35799_, _35800_, _35801_, _35802_, _35803_, _35804_, _35805_, _35806_, _35807_, _35808_, _35809_, _35810_, _35811_, _35812_, _35813_, _35814_, _35815_, _35816_, _35817_, _35818_, _35819_, _35820_, _35821_, _35822_, _35823_, _35824_, _35825_, _35826_, _35827_, _35828_, _35829_, _35830_, _35831_, _35832_, _35833_, _35834_, _35835_, _35836_, _35837_, _35838_, _35839_, _35840_, _35841_, _35842_, _35843_, _35844_, _35845_, _35846_, _35847_, _35848_, _35849_, _35850_, _35851_, _35852_, _35853_, _35854_, _35855_, _35856_, _35857_, _35858_, _35859_, _35860_, _35861_, _35862_, _35863_, _35864_, _35865_, _35866_, _35867_, _35868_, _35869_, _35870_, _35871_, _35872_, _35873_, _35874_, _35875_, _35876_, _35877_, _35878_, _35879_, _35880_, _35881_, _35882_, _35883_, _35884_, _35885_, _35886_, _35887_, _35888_, _35889_, _35890_, _35891_, _35892_, _35893_, _35894_, _35895_, _35896_, _35897_, _35898_, _35899_, _35900_, _35901_, _35902_, _35903_, _35904_, _35905_, _35906_, _35907_, _35908_, _35909_, _35910_, _35911_, _35912_, _35913_, _35914_, _35915_, _35916_, _35917_, _35918_, _35919_, _35920_, _35921_, _35922_, _35923_, _35924_, _35925_, _35926_, _35927_, _35928_, _35929_, _35930_, _35931_, _35932_, _35933_, _35934_, _35935_, _35936_, _35937_, _35938_, _35939_, _35940_, _35941_, _35942_, _35943_, _35944_, _35945_, _35946_, _35947_, _35948_, _35949_, _35950_, _35951_, _35952_, _35953_, _35954_, _35955_, _35956_, _35957_, _35958_, _35959_, _35960_, _35961_, _35962_, _35963_, _35964_, _35965_, _35966_, _35967_, _35968_, _35969_, _35970_, _35971_, _35972_, _35973_, _35974_, _35975_, _35976_, _35977_, _35978_, _35979_, _35980_, _35981_, _35982_, _35983_, _35984_, _35985_, _35986_, _35987_, _35988_, _35989_, _35990_, _35991_, _35992_, _35993_, _35994_, _35995_, _35996_, _35997_, _35998_, _35999_, _36000_, _36001_, _36002_, _36003_, _36004_, _36005_, _36006_, _36007_, _36008_, _36009_, _36010_, _36011_, _36012_, _36013_, _36014_, _36015_, _36016_, _36017_, _36018_, _36019_, _36020_, _36021_, _36022_, _36023_, _36024_, _36025_, _36026_, _36027_, _36028_, _36029_, _36030_, _36031_, _36032_, _36033_, _36034_, _36035_, _36036_, _36037_, _36038_, _36039_, _36040_, _36041_, _36042_, _36043_, _36044_, _36045_, _36046_, _36047_, _36048_, _36049_, _36050_, _36051_, _36052_, _36053_, _36054_, _36055_, _36056_, _36057_, _36058_, _36059_, _36060_, _36061_, _36062_, _36063_, _36064_, _36065_, _36066_, _36067_, _36068_, _36069_, _36070_, _36071_, _36072_, _36073_, _36074_, _36075_, _36076_, _36077_, _36078_, _36079_, _36080_, _36081_, _36082_, _36083_, _36084_, _36085_, _36086_, _36087_, _36088_, _36089_, _36090_, _36091_, _36092_, _36093_, _36094_, _36095_, _36096_, _36097_, _36098_, _36099_, _36100_, _36101_, _36102_, _36103_, _36104_, _36105_, _36106_, _36107_, _36108_, _36109_, _36110_, _36111_, _36112_, _36113_, _36114_, _36115_, _36116_, _36117_, _36118_, _36119_, _36120_, _36121_, _36122_, _36123_, _36124_, _36125_, _36126_, _36127_, _36128_, _36129_, _36130_, _36131_, _36132_, _36133_, _36134_, _36135_, _36136_, _36137_, _36138_, _36139_, _36140_, _36141_, _36142_, _36143_, _36144_, _36145_, _36146_, _36147_, _36148_, _36149_, _36150_, _36151_, _36152_, _36153_, _36154_, _36155_, _36156_, _36157_, _36158_, _36159_, _36160_, _36161_, _36162_, _36163_, _36164_, _36165_, _36166_, _36167_, _36168_, _36169_, _36170_, _36171_, _36172_, _36173_, _36174_, _36175_, _36176_, _36177_, _36178_, _36179_, _36180_, _36181_, _36182_, _36183_, _36184_, _36185_, _36186_, _36187_, _36188_, _36189_, _36190_, _36191_, _36192_, _36193_, _36194_, _36195_, _36196_, _36197_, _36198_, _36199_, _36200_, _36201_, _36202_, _36203_, _36204_, _36205_, _36206_, _36207_, _36208_, _36209_, _36210_, _36211_, _36212_, _36213_, _36214_, _36215_, _36216_, _36217_, _36218_, _36219_, _36220_, _36221_, _36222_, _36223_, _36224_, _36225_, _36226_, _36227_, _36228_, _36229_, _36230_, _36231_, _36232_, _36233_, _36234_, _36235_, _36236_, _36237_, _36238_, _36239_, _36240_, _36241_, _36242_, _36243_, _36244_, _36245_, _36246_, _36247_, _36248_, _36249_, _36250_, _36251_, _36252_, _36253_, _36254_, _36255_, _36256_, _36257_, _36258_, _36259_, _36260_, _36261_, _36262_, _36263_, _36264_, _36265_, _36266_, _36267_, _36268_, _36269_, _36270_, _36271_, _36272_, _36273_, _36274_, _36275_, _36276_, _36277_, _36278_, _36279_, _36280_, _36281_, _36282_, _36283_, _36284_, _36285_, _36286_, _36287_, _36288_, _36289_, _36290_, _36291_, _36292_, _36293_, _36294_, _36295_, _36296_, _36297_, _36298_, _36299_, _36300_, _36301_, _36302_, _36303_, _36304_, _36305_, _36306_, _36307_, _36308_, _36309_, _36310_, _36311_, _36312_, _36313_, _36314_, _36315_, _36316_, _36317_, _36318_, _36319_, _36320_, _36321_, _36322_, _36323_, _36324_, _36325_, _36326_, _36327_, _36328_, _36329_, _36330_, _36331_, _36332_, _36333_, _36334_, _36335_, _36336_, _36337_, _36338_, _36339_, _36340_, _36341_, _36342_, _36343_, _36344_, _36345_, _36346_, _36347_, _36348_, _36349_, _36350_, _36351_, _36352_, _36353_, _36354_, _36355_, _36356_, _36357_, _36358_, _36359_, _36360_, _36361_, _36362_, _36363_, _36364_, _36365_, _36366_, _36367_, _36368_, _36369_, _36370_, _36371_, _36372_, _36373_, _36374_, _36375_, _36376_, _36377_, _36378_, _36379_, _36380_, _36381_, _36382_, _36383_, _36384_, _36385_, _36386_, _36387_, _36388_, _36389_, _36390_, _36391_, _36392_, _36393_, _36394_, _36395_, _36396_, _36397_, _36398_, _36399_, _36400_, _36401_, _36402_, _36403_, _36404_, _36405_, _36406_, _36407_, _36408_, _36409_, _36410_, _36411_, _36412_, _36413_, _36414_, _36415_, _36416_, _36417_, _36418_, _36419_, _36420_, _36421_, _36422_, _36423_, _36424_, _36425_, _36426_, _36427_, _36428_, _36429_, _36430_, _36431_, _36432_, _36433_, _36434_, _36435_, _36436_, _36437_, _36438_, _36439_, _36440_, _36441_, _36442_, _36443_, _36444_, _36445_, _36446_, _36447_, _36448_, _36449_, _36450_, _36451_, _36452_, _36453_, _36454_, _36455_, _36456_, _36457_, _36458_, _36459_, _36460_, _36461_, _36462_, _36463_, _36464_, _36465_, _36466_, _36467_, _36468_, _36469_, _36470_, _36471_, _36472_, _36473_, _36474_, _36475_, _36476_, _36477_, _36478_, _36479_, _36480_, _36481_, _36482_, _36483_, _36484_, _36485_, _36486_, _36487_, _36488_, _36489_, _36490_, _36491_, _36492_, _36493_, _36494_, _36495_, _36496_, _36497_, _36498_, _36499_, _36500_, _36501_, _36502_, _36503_, _36504_, _36505_, _36506_, _36507_, _36508_, _36509_, _36510_, _36511_, _36512_, _36513_, _36514_, _36515_, _36516_, _36517_, _36518_, _36519_, _36520_, _36521_, _36522_, _36523_, _36524_, _36525_, _36526_, _36527_, _36528_, _36529_, _36530_, _36531_, _36532_, _36533_, _36534_, _36535_, _36536_, _36537_, _36538_, _36539_, _36540_, _36541_, _36542_, _36543_, _36544_, _36545_, _36546_, _36547_, _36548_, _36549_, _36550_, _36551_, _36552_, _36553_, _36554_, _36555_, _36556_, _36557_, _36558_, _36559_, _36560_, _36561_, _36562_, _36563_, _36564_, _36565_, _36566_, _36567_, _36568_, _36569_, _36570_, _36571_, _36572_, _36573_, _36574_, _36575_, _36576_, _36577_, _36578_, _36579_, _36580_, _36581_, _36582_, _36583_, _36584_, _36585_, _36586_, _36587_, _36588_, _36589_, _36590_, _36591_, _36592_, _36593_, _36594_, _36595_, _36596_, _36597_, _36598_, _36599_, _36600_, _36601_, _36602_, _36603_, _36604_, _36605_, _36606_, _36607_, _36608_, _36609_, _36610_, _36611_, _36612_, _36613_, _36614_, _36615_, _36616_, _36617_, _36618_, _36619_, _36620_, _36621_, _36622_, _36623_, _36624_, _36625_, _36626_, _36627_, _36628_, _36629_, _36630_, _36631_, _36632_, _36633_, _36634_, _36635_, _36636_, _36637_, _36638_, _36639_, _36640_, _36641_, _36642_, _36643_, _36644_, _36645_, _36646_, _36647_, _36648_, _36649_, _36650_, _36651_, _36652_, _36653_, _36654_, _36655_, _36656_, _36657_, _36658_, _36659_, _36660_, _36661_, _36662_, _36663_, _36664_, _36665_, _36666_, _36667_, _36668_, _36669_, _36670_, _36671_, _36672_, _36673_, _36674_, _36675_, _36676_, _36677_, _36678_, _36679_, _36680_, _36681_, _36682_, _36683_, _36684_, _36685_, _36686_, _36687_, _36688_, _36689_, _36690_, _36691_, _36692_, _36693_, _36694_, _36695_, _36696_, _36697_, _36698_, _36699_, _36700_, _36701_, _36702_, _36703_, _36704_, _36705_, _36706_, _36707_, _36708_, _36709_, _36710_, _36711_, _36712_, _36713_, _36714_, _36715_, _36716_, _36717_, _36718_, _36719_, _36720_, _36721_, _36722_, _36723_, _36724_, _36725_, _36726_, _36727_, _36728_, _36729_, _36730_, _36731_, _36732_, _36733_, _36734_, _36735_, _36736_, _36737_, _36738_, _36739_, _36740_, _36741_, _36742_, _36743_, _36744_, _36745_, _36746_, _36747_, _36748_, _36749_, _36750_, _36751_, _36752_, _36753_, _36754_, _36755_, _36756_, _36757_, _36758_, _36759_, _36760_, _36761_, _36762_, _36763_, _36764_, _36765_, _36766_, _36767_, _36768_, _36769_, _36770_, _36771_, _36772_, _36773_, _36774_, _36775_, _36776_, _36777_, _36778_, _36779_, _36780_, _36781_, _36782_, _36783_, _36784_, _36785_, _36786_, _36787_, _36788_, _36789_, _36790_, _36791_, _36792_, _36793_, _36794_, _36795_, _36796_, _36797_, _36798_, _36799_, _36800_, _36801_, _36802_, _36803_, _36804_, _36805_, _36806_, _36807_, _36808_, _36809_, _36810_, _36811_, _36812_, _36813_, _36814_, _36815_, _36816_, _36817_, _36818_, _36819_, _36820_, _36821_, _36822_, _36823_, _36824_, _36825_, _36826_, _36827_, _36828_, _36829_, _36830_, _36831_, _36832_, _36833_, _36834_, _36835_, _36836_, _36837_, _36838_, _36839_, _36840_, _36841_, _36842_, _36843_, _36844_, _36845_, _36846_, _36847_, _36848_, _36849_, _36850_, _36851_, _36852_, _36853_, _36854_, _36855_, _36856_, _36857_, _36858_, _36859_, _36860_, _36861_, _36862_, _36863_, _36864_, _36865_, _36866_, _36867_, _36868_, _36869_, _36870_, _36871_, _36872_, _36873_, _36874_, _36875_, _36876_, _36877_, _36878_, _36879_, _36880_, _36881_, _36882_, _36883_, _36884_, _36885_, _36886_, _36887_, _36888_, _36889_, _36890_, _36891_, _36892_, _36893_, _36894_, _36895_, _36896_, _36897_, _36898_, _36899_, _36900_, _36901_, _36902_, _36903_, _36904_, _36905_, _36906_, _36907_, _36908_, _36909_, _36910_, _36911_, _36912_, _36913_, _36914_, _36915_, _36916_, _36917_, _36918_, _36919_, _36920_, _36921_, _36922_, _36923_, _36924_, _36925_, _36926_, _36927_, _36928_, _36929_, _36930_, _36931_, _36932_, _36933_, _36934_, _36935_, _36936_, _36937_, _36938_, _36939_, _36940_, _36941_, _36942_, _36943_, _36944_, _36945_, _36946_, _36947_, _36948_, _36949_, _36950_, _36951_, _36952_, _36953_, _36954_, _36955_, _36956_, _36957_, _36958_, _36959_, _36960_, _36961_, _36962_, _36963_, _36964_, _36965_, _36966_, _36967_, _36968_, _36969_, _36970_, _36971_, _36972_, _36973_, _36974_, _36975_, _36976_, _36977_, _36978_, _36979_, _36980_, _36981_, _36982_, _36983_, _36984_, _36985_, _36986_, _36987_, _36988_, _36989_, _36990_, _36991_, _36992_, _36993_, _36994_, _36995_, _36996_, _36997_, _36998_, _36999_, _37000_, _37001_, _37002_, _37003_, _37004_, _37005_, _37006_, _37007_, _37008_, _37009_, _37010_, _37011_, _37012_, _37013_, _37014_, _37015_, _37016_, _37017_, _37018_, _37019_, _37020_, _37021_, _37022_, _37023_, _37024_, _37025_, _37026_, _37027_, _37028_, _37029_, _37030_, _37031_, _37032_, _37033_, _37034_, _37035_, _37036_, _37037_, _37038_, _37039_, _37040_, _37041_, _37042_, _37043_, _37044_, _37045_, _37046_, _37047_, _37048_, _37049_, _37050_, _37051_, _37052_, _37053_, _37054_, _37055_, _37056_, _37057_, _37058_, _37059_, _37060_, _37061_, _37062_, _37063_, _37064_, _37065_, _37066_, _37067_, _37068_, _37069_, _37070_, _37071_, _37072_, _37073_, _37074_, _37075_, _37076_, _37077_, _37078_, _37079_, _37080_, _37081_, _37082_, _37083_, _37084_, _37085_, _37086_, _37087_, _37088_, _37089_, _37090_, _37091_, _37092_, _37093_, _37094_, _37095_, _37096_, _37097_, _37098_, _37099_, _37100_, _37101_, _37102_, _37103_, _37104_, _37105_, _37106_, _37107_, _37108_, _37109_, _37110_, _37111_, _37112_, _37113_, _37114_, _37115_, _37116_, _37117_, _37118_, _37119_, _37120_, _37121_, _37122_, _37123_, _37124_, _37125_, _37126_, _37127_, _37128_, _37129_, _37130_, _37131_, _37132_, _37133_, _37134_, _37135_, _37136_, _37137_, _37138_, _37139_, _37140_, _37141_, _37142_, _37143_, _37144_, _37145_, _37146_, _37147_, _37148_, _37149_, _37150_, _37151_, _37152_, _37153_, _37154_, _37155_, _37156_, _37157_, _37158_, _37159_, _37160_, _37161_, _37162_, _37163_, _37164_, _37165_, _37166_, _37167_, _37168_, _37169_, _37170_, _37171_, _37172_, _37173_, _37174_, _37175_, _37176_, _37177_, _37178_, _37179_, _37180_, _37181_, _37182_, _37183_, _37184_, _37185_, _37186_, _37187_, _37188_, _37189_, _37190_, _37191_, _37192_, _37193_, _37194_, _37195_, _37196_, _37197_, _37198_, _37199_, _37200_, _37201_, _37202_, _37203_, _37204_, _37205_, _37206_, _37207_, _37208_, _37209_, _37210_, _37211_, _37212_, _37213_, _37214_, _37215_, _37216_, _37217_, _37218_, _37219_, _37220_, _37221_, _37222_, _37223_, _37224_, _37225_, _37226_, _37227_, _37228_, _37229_, _37230_, _37231_, _37232_, _37233_, _37234_, _37235_, _37236_, _37237_, _37238_, _37239_, _37240_, _37241_, _37242_, _37243_, _37244_, _37245_, _37246_, _37247_, _37248_, _37249_, _37250_, _37251_, _37252_, _37253_, _37254_, _37255_, _37256_, _37257_, _37258_, _37259_, _37260_, _37261_, _37262_, _37263_, _37264_, _37265_, _37266_, _37267_, _37268_, _37269_, _37270_, _37271_, _37272_, _37273_, _37274_, _37275_, _37276_, _37277_, _37278_, _37279_, _37280_, _37281_, _37282_, _37283_, _37284_, _37285_, _37286_, _37287_, _37288_, _37289_, _37290_, _37291_, _37292_, _37293_, _37294_, _37295_, _37296_, _37297_, _37298_, _37299_, _37300_, _37301_, _37302_, _37303_, _37304_, _37305_, _37306_, _37307_, _37308_, _37309_, _37310_, _37311_, _37312_, _37313_, _37314_, _37315_, _37316_, _37317_, _37318_, _37319_, _37320_, _37321_, _37322_, _37323_, _37324_, _37325_, _37326_, _37327_, _37328_, _37329_, _37330_, _37331_, _37332_, _37333_, _37334_, _37335_, _37336_, _37337_, _37338_, _37339_, _37340_, _37341_, _37342_, _37343_, _37344_, _37345_, _37346_, _37347_, _37348_, _37349_, _37350_, _37351_, _37352_, _37353_, _37354_, _37355_, _37356_, _37357_, _37358_, _37359_, _37360_, _37361_, _37362_, _37363_, _37364_, _37365_, _37366_, _37367_, _37368_, _37369_, _37370_, _37371_, _37372_, _37373_, _37374_, _37375_, _37376_, _37377_, _37378_, _37379_, _37380_, _37381_, _37382_, _37383_, _37384_, _37385_, _37386_, _37387_, _37388_, _37389_, _37390_, _37391_, _37392_, _37393_, _37394_, _37395_, _37396_, _37397_, _37398_, _37399_, _37400_, _37401_, _37402_, _37403_, _37404_, _37405_, _37406_, _37407_, _37408_, _37409_, _37410_, _37411_, _37412_, _37413_, _37414_, _37415_, _37416_, _37417_, _37418_, _37419_, _37420_, _37421_, _37422_, _37423_, _37424_, _37425_, _37426_, _37427_, _37428_, _37429_, _37430_, _37431_, _37432_, _37433_, _37434_, _37435_, _37436_, _37437_, _37438_, _37439_, _37440_, _37441_, _37442_, _37443_, _37444_, _37445_, _37446_, _37447_, _37448_, _37449_, _37450_, _37451_, _37452_, _37453_, _37454_, _37455_, _37456_, _37457_, _37458_, _37459_, _37460_, _37461_, _37462_, _37463_, _37464_, _37465_, _37466_, _37467_, _37468_, _37469_, _37470_, _37471_, _37472_, _37473_, _37474_, _37475_, _37476_, _37477_, _37478_, _37479_, _37480_, _37481_, _37482_, _37483_, _37484_, _37485_, _37486_, _37487_, _37488_, _37489_, _37490_, _37491_, _37492_, _37493_, _37494_, _37495_, _37496_, _37497_, _37498_, _37499_, _37500_, _37501_, _37502_, _37503_, _37504_, _37505_, _37506_, _37507_, _37508_, _37509_, _37510_, _37511_, _37512_, _37513_, _37514_, _37515_, _37516_, _37517_, _37518_, _37519_, _37520_, _37521_, _37522_, _37523_, _37524_, _37525_, _37526_, _37527_, _37528_, _37529_, _37530_, _37531_, _37532_, _37533_, _37534_, _37535_, _37536_, _37537_, _37538_, _37539_, _37540_, _37541_, _37542_, _37543_, _37544_, _37545_, _37546_, _37547_, _37548_, _37549_, _37550_, _37551_, _37552_, _37553_, _37554_, _37555_, _37556_, _37557_, _37558_, _37559_, _37560_, _37561_, _37562_, _37563_, _37564_, _37565_, _37566_, _37567_, _37568_, _37569_, _37570_, _37571_, _37572_, _37573_, _37574_, _37575_, _37576_, _37577_, _37578_, _37579_, _37580_, _37581_, _37582_, _37583_, _37584_, _37585_, _37586_, _37587_, _37588_, _37589_, _37590_, _37591_, _37592_, _37593_, _37594_, _37595_, _37596_, _37597_, _37598_, _37599_, _37600_, _37601_, _37602_, _37603_, _37604_, _37605_, _37606_, _37607_, _37608_, _37609_, _37610_, _37611_, _37612_, _37613_, _37614_, _37615_, _37616_, _37617_, _37618_, _37619_, _37620_, _37621_, _37622_, _37623_, _37624_, _37625_, _37626_, _37627_, _37628_, _37629_, _37630_, _37631_, _37632_, _37633_, _37634_, _37635_, _37636_, _37637_, _37638_, _37639_, _37640_, _37641_, _37642_, _37643_, _37644_, _37645_, _37646_, _37647_, _37648_, _37649_, _37650_, _37651_, _37652_, _37653_, _37654_, _37655_, _37656_, _37657_, _37658_, _37659_, _37660_, _37661_, _37662_, _37663_, _37664_, _37665_, _37666_, _37667_, _37668_, _37669_, _37670_, _37671_, _37672_, _37673_, _37674_, _37675_, _37676_, _37677_, _37678_, _37679_, _37680_, _37681_, _37682_, _37683_, _37684_, _37685_, _37686_, _37687_, _37688_, _37689_, _37690_, _37691_, _37692_, _37693_, _37694_, _37695_, _37696_, _37697_, _37698_, _37699_, _37700_, _37701_, _37702_, _37703_, _37704_, _37705_, _37706_, _37707_, _37708_, _37709_, _37710_, _37711_, _37712_, _37713_, _37714_, _37715_, _37716_, _37717_, _37718_, _37719_, _37720_, _37721_, _37722_, _37723_, _37724_, _37725_, _37726_, _37727_, _37728_, _37729_, _37730_, _37731_, _37732_, _37733_, _37734_, _37735_, _37736_, _37737_, _37738_, _37739_, _37740_, _37741_, _37742_, _37743_, _37744_, _37745_, _37746_, _37747_, _37748_, _37749_, _37750_, _37751_, _37752_, _37753_, _37754_, _37755_, _37756_, _37757_, _37758_, _37759_, _37760_, _37761_, _37762_, _37763_, _37764_, _37765_, _37766_, _37767_, _37768_, _37769_, _37770_, _37771_, _37772_, _37773_, _37774_, _37775_, _37776_, _37777_, _37778_, _37779_, _37780_, _37781_, _37782_, _37783_, _37784_, _37785_, _37786_, _37787_, _37788_, _37789_, _37790_, _37791_, _37792_, _37793_, _37794_, _37795_, _37796_, _37797_, _37798_, _37799_, _37800_, _37801_, _37802_, _37803_, _37804_, _37805_, _37806_, _37807_, _37808_, _37809_, _37810_, _37811_, _37812_, _37813_, _37814_, _37815_, _37816_, _37817_, _37818_, _37819_, _37820_, _37821_, _37822_, _37823_, _37824_, _37825_, _37826_, _37827_, _37828_, _37829_, _37830_, _37831_, _37832_, _37833_, _37834_, _37835_, _37836_, _37837_, _37838_, _37839_, _37840_, _37841_, _37842_, _37843_, _37844_, _37845_, _37846_, _37847_, _37848_, _37849_, _37850_, _37851_, _37852_, _37853_, _37854_, _37855_, _37856_, _37857_, _37858_, _37859_, _37860_, _37861_, _37862_, _37863_, _37864_, _37865_, _37866_, _37867_, _37868_, _37869_, _37870_, _37871_, _37872_, _37873_, _37874_, _37875_, _37876_, _37877_, _37878_, _37879_, _37880_, _37881_, _37882_, _37883_, _37884_, _37885_, _37886_, _37887_, _37888_, _37889_, _37890_, _37891_, _37892_, _37893_, _37894_, _37895_, _37896_, _37897_, _37898_, _37899_, _37900_, _37901_, _37902_, _37903_, _37904_, _37905_, _37906_, _37907_, _37908_, _37909_, _37910_, _37911_, _37912_, _37913_, _37914_, _37915_, _37916_, _37917_, _37918_, _37919_, _37920_, _37921_, _37922_, _37923_, _37924_, _37925_, _37926_, _37927_, _37928_, _37929_, _37930_, _37931_, _37932_, _37933_, _37934_, _37935_, _37936_, _37937_, _37938_, _37939_, _37940_, _37941_, _37942_, _37943_, _37944_, _37945_, _37946_, _37947_, _37948_, _37949_, _37950_, _37951_, _37952_, _37953_, _37954_, _37955_, _37956_, _37957_, _37958_, _37959_, _37960_, _37961_, _37962_, _37963_, _37964_, _37965_, _37966_, _37967_, _37968_, _37969_, _37970_, _37971_, _37972_, _37973_, _37974_, _37975_, _37976_, _37977_, _37978_, _37979_, _37980_, _37981_, _37982_, _37983_, _37984_, _37985_, _37986_, _37987_, _37988_, _37989_, _37990_, _37991_, _37992_, _37993_, _37994_, _37995_, _37996_, _37997_, _37998_, _37999_, _38000_, _38001_, _38002_, _38003_, _38004_, _38005_, _38006_, _38007_, _38008_, _38009_, _38010_, _38011_, _38012_, _38013_, _38014_, _38015_, _38016_, _38017_, _38018_, _38019_, _38020_, _38021_, _38022_, _38023_, _38024_, _38025_, _38026_, _38027_, _38028_, _38029_, _38030_, _38031_, _38032_, _38033_, _38034_, _38035_, _38036_, _38037_, _38038_, _38039_, _38040_, _38041_, _38042_, _38043_, _38044_, _38045_, _38046_, _38047_, _38048_, _38049_, _38050_, _38051_, _38052_, _38053_, _38054_, _38055_, _38056_, _38057_, _38058_, _38059_, _38060_, _38061_, _38062_, _38063_, _38064_, _38065_, _38066_, _38067_, _38068_, _38069_, _38070_, _38071_, _38072_, _38073_, _38074_, _38075_, _38076_, _38077_, _38078_, _38079_, _38080_, _38081_, _38082_, _38083_, _38084_, _38085_, _38086_, _38087_, _38088_, _38089_, _38090_, _38091_, _38092_, _38093_, _38094_, _38095_, _38096_, _38097_, _38098_, _38099_, _38100_, _38101_, _38102_, _38103_, _38104_, _38105_, _38106_, _38107_, _38108_, _38109_, _38110_, _38111_, _38112_, _38113_, _38114_, _38115_, _38116_, _38117_, _38118_, _38119_, _38120_, _38121_, _38122_, _38123_, _38124_, _38125_, _38126_, _38127_, _38128_, _38129_, _38130_, _38131_, _38132_, _38133_, _38134_, _38135_, _38136_, _38137_, _38138_, _38139_, _38140_, _38141_, _38142_, _38143_, _38144_, _38145_, _38146_, _38147_, _38148_, _38149_, _38150_, _38151_, _38152_, _38153_, _38154_, _38155_, _38156_, _38157_, _38158_, _38159_, _38160_, _38161_, _38162_, _38163_, _38164_, _38165_, _38166_, _38167_, _38168_, _38169_, _38170_, _38171_, _38172_, _38173_, _38174_, _38175_, _38176_, _38177_, _38178_, _38179_, _38180_, _38181_, _38182_, _38183_, _38184_, _38185_, _38186_, _38187_, _38188_, _38189_, _38190_, _38191_, _38192_, _38193_, _38194_, _38195_, _38196_, _38197_, _38198_, _38199_, _38200_, _38201_, _38202_, _38203_, _38204_, _38205_, _38206_, _38207_, _38208_, _38209_, _38210_, _38211_, _38212_, _38213_, _38214_, _38215_, _38216_, _38217_, _38218_, _38219_, _38220_, _38221_, _38222_, _38223_, _38224_, _38225_, _38226_, _38227_, _38228_, _38229_, _38230_, _38231_, _38232_, _38233_, _38234_, _38235_, _38236_, _38237_, _38238_, _38239_, _38240_, _38241_, _38242_, _38243_, _38244_, _38245_, _38246_, _38247_, _38248_, _38249_, _38250_, _38251_, _38252_, _38253_, _38254_, _38255_, _38256_, _38257_, _38258_, _38259_, _38260_, _38261_, _38262_, _38263_, _38264_, _38265_, _38266_, _38267_, _38268_, _38269_, _38270_, _38271_, _38272_, _38273_, _38274_, _38275_, _38276_, _38277_, _38278_, _38279_, _38280_, _38281_, _38282_, _38283_, _38284_, _38285_, _38286_, _38287_, _38288_, _38289_, _38290_, _38291_, _38292_, _38293_, _38294_, _38295_, _38296_, _38297_, _38298_, _38299_, _38300_, _38301_, _38302_, _38303_, _38304_, _38305_, _38306_, _38307_, _38308_, _38309_, _38310_, _38311_, _38312_, _38313_, _38314_, _38315_, _38316_, _38317_, _38318_, _38319_, _38320_, _38321_, _38322_, _38323_, _38324_, _38325_, _38326_, _38327_, _38328_, _38329_, _38330_, _38331_, _38332_, _38333_, _38334_, _38335_, _38336_, _38337_, _38338_, _38339_, _38340_, _38341_, _38342_, _38343_, _38344_, _38345_, _38346_, _38347_, _38348_, _38349_, _38350_, _38351_, _38352_, _38353_, _38354_, _38355_, _38356_, _38357_, _38358_, _38359_, _38360_, _38361_, _38362_, _38363_, _38364_, _38365_, _38366_, _38367_, _38368_, _38369_, _38370_, _38371_, _38372_, _38373_, _38374_, _38375_, _38376_, _38377_, _38378_, _38379_, _38380_, _38381_, _38382_, _38383_, _38384_, _38385_, _38386_, _38387_, _38388_, _38389_, _38390_, _38391_, _38392_, _38393_, _38394_, _38395_, _38396_, _38397_, _38398_, _38399_, _38400_, _38401_, _38402_, _38403_, _38404_, _38405_, _38406_, _38407_, _38408_, _38409_, _38410_, _38411_, _38412_, _38413_, _38414_, _38415_, _38416_, _38417_, _38418_, _38419_, _38420_, _38421_, _38422_, _38423_, _38424_, _38425_, _38426_, _38427_, _38428_, _38429_, _38430_, _38431_, _38432_, _38433_, _38434_, _38435_, _38436_, _38437_, _38438_, _38439_, _38440_, _38441_, _38442_, _38443_, _38444_, _38445_, _38446_, _38447_, _38448_, _38449_, _38450_, _38451_, _38452_, _38453_, _38454_, _38455_, _38456_, _38457_, _38458_, _38459_, _38460_, _38461_, _38462_, _38463_, _38464_, _38465_, _38466_, _38467_, _38468_, _38469_, _38470_, _38471_, _38472_, _38473_, _38474_, _38475_, _38476_, _38477_, _38478_, _38479_, _38480_, _38481_, _38482_, _38483_, _38484_, _38485_, _38486_, _38487_, _38488_, _38489_, _38490_, _38491_, _38492_, _38493_, _38494_, _38495_, _38496_, _38497_, _38498_, _38499_, _38500_, _38501_, _38502_, _38503_, _38504_, _38505_, _38506_, _38507_, _38508_, _38509_, _38510_, _38511_, _38512_, _38513_, _38514_, _38515_, _38516_, _38517_, _38518_, _38519_, _38520_, _38521_, _38522_, _38523_, _38524_, _38525_, _38526_, _38527_, _38528_, _38529_, _38530_, _38531_, _38532_, _38533_, _38534_, _38535_, _38536_, _38537_, _38538_, _38539_, _38540_, _38541_, _38542_, _38543_, _38544_, _38545_, _38546_, _38547_, _38548_, _38549_, _38550_, _38551_, _38552_, _38553_, _38554_, _38555_, _38556_, _38557_, _38558_, _38559_, _38560_, _38561_, _38562_, _38563_, _38564_, _38565_, _38566_, _38567_, _38568_, _38569_, _38570_, _38571_, _38572_, _38573_, _38574_, _38575_, _38576_, _38577_, _38578_, _38579_, _38580_, _38581_, _38582_, _38583_, _38584_, _38585_, _38586_, _38587_, _38588_, _38589_, _38590_, _38591_, _38592_, _38593_, _38594_, _38595_, _38596_, _38597_, _38598_, _38599_, _38600_, _38601_, _38602_, _38603_, _38604_, _38605_, _38606_, _38607_, _38608_, _38609_, _38610_, _38611_, _38612_, _38613_, _38614_, _38615_, _38616_, _38617_, _38618_, _38619_, _38620_, _38621_, _38622_, _38623_, _38624_, _38625_, _38626_, _38627_, _38628_, _38629_, _38630_, _38631_, _38632_, _38633_, _38634_, _38635_, _38636_, _38637_, _38638_, _38639_, _38640_, _38641_, _38642_, _38643_, _38644_, _38645_, _38646_, _38647_, _38648_, _38649_, _38650_, _38651_, _38652_, _38653_, _38654_, _38655_, _38656_, _38657_, _38658_, _38659_, _38660_, _38661_, _38662_, _38663_, _38664_, _38665_, _38666_, _38667_, _38668_, _38669_, _38670_, _38671_, _38672_, _38673_, _38674_, _38675_, _38676_, _38677_, _38678_, _38679_, _38680_, _38681_, _38682_, _38683_, _38684_, _38685_, _38686_, _38687_, _38688_, _38689_, _38690_, _38691_, _38692_, _38693_, _38694_, _38695_, _38696_, _38697_, _38698_, _38699_, _38700_, _38701_, _38702_, _38703_, _38704_, _38705_, _38706_, _38707_, _38708_, _38709_, _38710_, _38711_, _38712_, _38713_, _38714_, _38715_, _38716_, _38717_, _38718_, _38719_, _38720_, _38721_, _38722_, _38723_, _38724_, _38725_, _38726_, _38727_, _38728_, _38729_, _38730_, _38731_, _38732_, _38733_, _38734_, _38735_, _38736_, _38737_, _38738_, _38739_, _38740_, _38741_, _38742_, _38743_, _38744_, _38745_, _38746_, _38747_, _38748_, _38749_, _38750_, _38751_, _38752_, _38753_, _38754_, _38755_, _38756_, _38757_, _38758_, _38759_, _38760_, _38761_, _38762_, _38763_, _38764_, _38765_, _38766_, _38767_, _38768_, _38769_, _38770_, _38771_, _38772_, _38773_, _38774_, _38775_, _38776_, _38777_, _38778_, _38779_, _38780_, _38781_, _38782_, _38783_, _38784_, _38785_, _38786_, _38787_, _38788_, _38789_, _38790_, _38791_, _38792_, _38793_, _38794_, _38795_, _38796_, _38797_, _38798_, _38799_, _38800_, _38801_, _38802_, _38803_, _38804_, _38805_, _38806_, _38807_, _38808_, _38809_, _38810_, _38811_, _38812_, _38813_, _38814_, _38815_, _38816_, _38817_, _38818_, _38819_, _38820_, _38821_, _38822_, _38823_, _38824_, _38825_, _38826_, _38827_, _38828_, _38829_, _38830_, _38831_, _38832_, _38833_, _38834_, _38835_, _38836_, _38837_, _38838_, _38839_, _38840_, _38841_, _38842_, _38843_, _38844_, _38845_, _38846_, _38847_, _38848_, _38849_, _38850_, _38851_, _38852_, _38853_, _38854_, _38855_, _38856_, _38857_, _38858_, _38859_, _38860_, _38861_, _38862_, _38863_, _38864_, _38865_, _38866_, _38867_, _38868_, _38869_, _38870_, _38871_, _38872_, _38873_, _38874_, _38875_, _38876_, _38877_, _38878_, _38879_, _38880_, _38881_, _38882_, _38883_, _38884_, _38885_, _38886_, _38887_, _38888_, _38889_, _38890_, _38891_, _38892_, _38893_, _38894_, _38895_, _38896_, _38897_, _38898_, _38899_, _38900_, _38901_, _38902_, _38903_, _38904_, _38905_, _38906_, _38907_, _38908_, _38909_, _38910_, _38911_, _38912_, _38913_, _38914_, _38915_, _38916_, _38917_, _38918_, _38919_, _38920_, _38921_, _38922_, _38923_, _38924_, _38925_, _38926_, _38927_, _38928_, _38929_, _38930_, _38931_, _38932_, _38933_, _38934_, _38935_, _38936_, _38937_, _38938_, _38939_, _38940_, _38941_, _38942_, _38943_, _38944_, _38945_, _38946_, _38947_, _38948_, _38949_, _38950_, _38951_, _38952_, _38953_, _38954_, _38955_, _38956_, _38957_, _38958_, _38959_, _38960_, _38961_, _38962_, _38963_, _38964_, _38965_, _38966_, _38967_, _38968_, _38969_, _38970_, _38971_, _38972_, _38973_, _38974_, _38975_, _38976_, _38977_, _38978_, _38979_, _38980_, _38981_, _38982_, _38983_, _38984_, _38985_, _38986_, _38987_, _38988_, _38989_, _38990_, _38991_, _38992_, _38993_, _38994_, _38995_, _38996_, _38997_, _38998_, _38999_, _39000_, _39001_, _39002_, _39003_, _39004_, _39005_, _39006_, _39007_, _39008_, _39009_, _39010_, _39011_, _39012_, _39013_, _39014_, _39015_, _39016_, _39017_, _39018_, _39019_, _39020_, _39021_, _39022_, _39023_, _39024_, _39025_, _39026_, _39027_, _39028_, _39029_, _39030_, _39031_, _39032_, _39033_, _39034_, _39035_, _39036_, _39037_, _39038_, _39039_, _39040_, _39041_, _39042_, _39043_, _39044_, _39045_, _39046_, _39047_, _39048_, _39049_, _39050_, _39051_, _39052_, _39053_, _39054_, _39055_, _39056_, _39057_, _39058_, _39059_, _39060_, _39061_, _39062_, _39063_, _39064_, _39065_, _39066_, _39067_, _39068_, _39069_, _39070_, _39071_, _39072_, _39073_, _39074_, _39075_, _39076_, _39077_, _39078_, _39079_, _39080_, _39081_, _39082_, _39083_, _39084_, _39085_, _39086_, _39087_, _39088_, _39089_, _39090_, _39091_, _39092_, _39093_, _39094_, _39095_, _39096_, _39097_, _39098_, _39099_, _39100_, _39101_, _39102_, _39103_, _39104_, _39105_, _39106_, _39107_, _39108_, _39109_, _39110_, _39111_, _39112_, _39113_, _39114_, _39115_, _39116_, _39117_, _39118_, _39119_, _39120_, _39121_, _39122_, _39123_, _39124_, _39125_, _39126_, _39127_, _39128_, _39129_, _39130_, _39131_, _39132_, _39133_, _39134_, _39135_, _39136_, _39137_, _39138_, _39139_, _39140_, _39141_, _39142_, _39143_, _39144_, _39145_, _39146_, _39147_, _39148_, _39149_, _39150_, _39151_, _39152_, _39153_, _39154_, _39155_, _39156_, _39157_, _39158_, _39159_, _39160_, _39161_, _39162_, _39163_, _39164_, _39165_, _39166_, _39167_, _39168_, _39169_, _39170_, _39171_, _39172_, _39173_, _39174_, _39175_, _39176_, _39177_, _39178_, _39179_, _39180_, _39181_, _39182_, _39183_, _39184_, _39185_, _39186_, _39187_, _39188_, _39189_, _39190_, _39191_, _39192_, _39193_, _39194_, _39195_, _39196_, _39197_, _39198_, _39199_, _39200_, _39201_, _39202_, _39203_, _39204_, _39205_, _39206_, _39207_, _39208_, _39209_, _39210_, _39211_, _39212_, _39213_, _39214_, _39215_, _39216_, _39217_, _39218_, _39219_, _39220_, _39221_, _39222_, _39223_, _39224_, _39225_, _39226_, _39227_, _39228_, _39229_, _39230_, _39231_, _39232_, _39233_, _39234_, _39235_, _39236_, _39237_, _39238_, _39239_, _39240_, _39241_, _39242_, _39243_, _39244_, _39245_, _39246_, _39247_, _39248_, _39249_, _39250_, _39251_, _39252_, _39253_, _39254_, _39255_, _39256_, _39257_, _39258_, _39259_, _39260_, _39261_, _39262_, _39263_, _39264_, _39265_, _39266_, _39267_, _39268_, _39269_, _39270_, _39271_, _39272_, _39273_, _39274_, _39275_, _39276_, _39277_, _39278_, _39279_, _39280_, _39281_, _39282_, _39283_, _39284_, _39285_, _39286_, _39287_, _39288_, _39289_, _39290_, _39291_, _39292_, _39293_, _39294_, _39295_, _39296_, _39297_, _39298_, _39299_, _39300_, _39301_, _39302_, _39303_, _39304_, _39305_, _39306_, _39307_, _39308_, _39309_, _39310_, _39311_, _39312_, _39313_, _39314_, _39315_, _39316_, _39317_, _39318_, _39319_, _39320_, _39321_, _39322_, _39323_, _39324_, _39325_, _39326_, _39327_, _39328_, _39329_, _39330_, _39331_, _39332_, _39333_, _39334_, _39335_, _39336_, _39337_, _39338_, _39339_, _39340_, _39341_, _39342_, _39343_, _39344_, _39345_, _39346_, _39347_, _39348_, _39349_, _39350_, _39351_, _39352_, _39353_, _39354_, _39355_, _39356_, _39357_, _39358_, _39359_, _39360_, _39361_, _39362_, _39363_, _39364_, _39365_, _39366_, _39367_, _39368_, _39369_, _39370_, _39371_, _39372_, _39373_, _39374_, _39375_, _39376_, _39377_, _39378_, _39379_, _39380_, _39381_, _39382_, _39383_, _39384_, _39385_, _39386_, _39387_, _39388_, _39389_, _39390_, _39391_, _39392_, _39393_, _39394_, _39395_, _39396_, _39397_, _39398_, _39399_, _39400_, _39401_, _39402_, _39403_, _39404_, _39405_, _39406_, _39407_, _39408_, _39409_, _39410_, _39411_, _39412_, _39413_, _39414_, _39415_, _39416_, _39417_, _39418_, _39419_, _39420_, _39421_, _39422_, _39423_, _39424_, _39425_, _39426_, _39427_, _39428_, _39429_, _39430_, _39431_, _39432_, _39433_, _39434_, _39435_, _39436_, _39437_, _39438_, _39439_, _39440_, _39441_, _39442_, _39443_, _39444_, _39445_, _39446_, _39447_, _39448_, _39449_, _39450_, _39451_, _39452_, _39453_, _39454_, _39455_, _39456_, _39457_, _39458_, _39459_, _39460_, _39461_, _39462_, _39463_, _39464_, _39465_, _39466_, _39467_, _39468_, _39469_, _39470_, _39471_, _39472_, _39473_, _39474_, _39475_, _39476_, _39477_, _39478_, _39479_, _39480_, _39481_, _39482_, _39483_, _39484_, _39485_, _39486_, _39487_, _39488_, _39489_, _39490_, _39491_, _39492_, _39493_, _39494_, _39495_, _39496_, _39497_, _39498_, _39499_, _39500_, _39501_, _39502_, _39503_, _39504_, _39505_, _39506_, _39507_, _39508_, _39509_, _39510_, _39511_, _39512_, _39513_, _39514_, _39515_, _39516_, _39517_, _39518_, _39519_, _39520_, _39521_, _39522_, _39523_, _39524_, _39525_, _39526_, _39527_, _39528_, _39529_, _39530_, _39531_, _39532_, _39533_, _39534_, _39535_, _39536_, _39537_, _39538_, _39539_, _39540_, _39541_, _39542_, _39543_, _39544_, _39545_, _39546_, _39547_, _39548_, _39549_, _39550_, _39551_, _39552_, _39553_, _39554_, _39555_, _39556_, _39557_, _39558_, _39559_, _39560_, _39561_, _39562_, _39563_, _39564_, _39565_, _39566_, _39567_, _39568_, _39569_, _39570_, _39571_, _39572_, _39573_, _39574_, _39575_, _39576_, _39577_, _39578_, _39579_, _39580_, _39581_, _39582_, _39583_, _39584_, _39585_, _39586_, _39587_, _39588_, _39589_, _39590_, _39591_, _39592_, _39593_, _39594_, _39595_, _39596_, _39597_, _39598_, _39599_, _39600_, _39601_, _39602_, _39603_, _39604_, _39605_, _39606_, _39607_, _39608_, _39609_, _39610_, _39611_, _39612_, _39613_, _39614_, _39615_, _39616_, _39617_, _39618_, _39619_, _39620_, _39621_, _39622_, _39623_, _39624_, _39625_, _39626_, _39627_, _39628_, _39629_, _39630_, _39631_, _39632_, _39633_, _39634_, _39635_, _39636_, _39637_, _39638_, _39639_, _39640_, _39641_, _39642_, _39643_, _39644_, _39645_, _39646_, _39647_, _39648_, _39649_, _39650_, _39651_, _39652_, _39653_, _39654_, _39655_, _39656_, _39657_, _39658_, _39659_, _39660_, _39661_, _39662_, _39663_, _39664_, _39665_, _39666_, _39667_, _39668_, _39669_, _39670_, _39671_, _39672_, _39673_, _39674_, _39675_, _39676_, _39677_, _39678_, _39679_, _39680_, _39681_, _39682_, _39683_, _39684_, _39685_, _39686_, _39687_, _39688_, _39689_, _39690_, _39691_, _39692_, _39693_, _39694_, _39695_, _39696_, _39697_, _39698_, _39699_, _39700_, _39701_, _39702_, _39703_, _39704_, _39705_, _39706_, _39707_, _39708_, _39709_, _39710_, _39711_, _39712_, _39713_, _39714_, _39715_, _39716_, _39717_, _39718_, _39719_, _39720_, _39721_, _39722_, _39723_, _39724_, _39725_, _39726_, _39727_, _39728_, _39729_, _39730_, _39731_, _39732_, _39733_, _39734_, _39735_, _39736_, _39737_, _39738_, _39739_, _39740_, _39741_, _39742_, _39743_, _39744_, _39745_, _39746_, _39747_, _39748_, _39749_, _39750_, _39751_, _39752_, _39753_, _39754_, _39755_, _39756_, _39757_, _39758_, _39759_, _39760_, _39761_, _39762_, _39763_, _39764_, _39765_, _39766_, _39767_, _39768_, _39769_, _39770_, _39771_, _39772_, _39773_, _39774_, _39775_, _39776_, _39777_, _39778_, _39779_, _39780_, _39781_, _39782_, _39783_, _39784_, _39785_, _39786_, _39787_, _39788_, _39789_, _39790_, _39791_, _39792_, _39793_, _39794_, _39795_, _39796_, _39797_, _39798_, _39799_, _39800_, _39801_, _39802_, _39803_, _39804_, _39805_, _39806_, _39807_, _39808_, _39809_, _39810_, _39811_, _39812_, _39813_, _39814_, _39815_, _39816_, _39817_, _39818_, _39819_, _39820_, _39821_, _39822_, _39823_, _39824_, _39825_, _39826_, _39827_, _39828_, _39829_, _39830_, _39831_, _39832_, _39833_, _39834_, _39835_, _39836_, _39837_, _39838_, _39839_, _39840_, _39841_, _39842_, _39843_, _39844_, _39845_, _39846_, _39847_, _39848_, _39849_, _39850_, _39851_, _39852_, _39853_, _39854_, _39855_, _39856_, _39857_, _39858_, _39859_, _39860_, _39861_, _39862_, _39863_, _39864_, _39865_, _39866_, _39867_, _39868_, _39869_, _39870_, _39871_, _39872_, _39873_, _39874_, _39875_, _39876_, _39877_, _39878_, _39879_, _39880_, _39881_, _39882_, _39883_, _39884_, _39885_, _39886_, _39887_, _39888_, _39889_, _39890_, _39891_, _39892_, _39893_, _39894_, _39895_, _39896_, _39897_, _39898_, _39899_, _39900_, _39901_, _39902_, _39903_, _39904_, _39905_, _39906_, _39907_, _39908_, _39909_, _39910_, _39911_, _39912_, _39913_, _39914_, _39915_, _39916_, _39917_, _39918_, _39919_, _39920_, _39921_, _39922_, _39923_, _39924_, _39925_, _39926_, _39927_, _39928_, _39929_, _39930_, _39931_, _39932_, _39933_, _39934_, _39935_, _39936_, _39937_, _39938_, _39939_, _39940_, _39941_, _39942_, _39943_, _39944_, _39945_, _39946_, _39947_, _39948_, _39949_, _39950_, _39951_, _39952_, _39953_, _39954_, _39955_, _39956_, _39957_, _39958_, _39959_, _39960_, _39961_, _39962_, _39963_, _39964_, _39965_, _39966_, _39967_, _39968_, _39969_, _39970_, _39971_, _39972_, _39973_, _39974_, _39975_, _39976_, _39977_, _39978_, _39979_, _39980_, _39981_, _39982_, _39983_, _39984_, _39985_, _39986_, _39987_, _39988_, _39989_, _39990_, _39991_, _39992_, _39993_, _39994_, _39995_, _39996_, _39997_, _39998_, _39999_, _40000_, _40001_, _40002_, _40003_, _40004_, _40005_, _40006_, _40007_, _40008_, _40009_, _40010_, _40011_, _40012_, _40013_, _40014_, _40015_, _40016_, _40017_, _40018_, _40019_, _40020_, _40021_, _40022_, _40023_, _40024_, _40025_, _40026_, _40027_, _40028_, _40029_, _40030_, _40031_, _40032_, _40033_, _40034_, _40035_, _40036_, _40037_, _40038_, _40039_, _40040_, _40041_, _40042_, _40043_, _40044_, _40045_, _40046_, _40047_, _40048_, _40049_, _40050_, _40051_, _40052_, _40053_, _40054_, _40055_, _40056_, _40057_, _40058_, _40059_, _40060_, _40061_, _40062_, _40063_, _40064_, _40065_, _40066_, _40067_, _40068_, _40069_, _40070_, _40071_, _40072_, _40073_, _40074_, _40075_, _40076_, _40077_, _40078_, _40079_, _40080_, _40081_, _40082_, _40083_, _40084_, _40085_, _40086_, _40087_, _40088_, _40089_, _40090_, _40091_, _40092_, _40093_, _40094_, _40095_, _40096_, _40097_, _40098_, _40099_, _40100_, _40101_, _40102_, _40103_, _40104_, _40105_, _40106_, _40107_, _40108_, _40109_, _40110_, _40111_, _40112_, _40113_, _40114_, _40115_, _40116_, _40117_, _40118_, _40119_, _40120_, _40121_, _40122_, _40123_, _40124_, _40125_, _40126_, _40127_, _40128_, _40129_, _40130_, _40131_, _40132_, _40133_, _40134_, _40135_, _40136_, _40137_, _40138_, _40139_, _40140_, _40141_, _40142_, _40143_, _40144_, _40145_, _40146_, _40147_, _40148_, _40149_, _40150_, _40151_, _40152_, _40153_, _40154_, _40155_, _40156_, _40157_, _40158_, _40159_, _40160_, _40161_, _40162_, _40163_, _40164_, _40165_, _40166_, _40167_, _40168_, _40169_, _40170_, _40171_, _40172_, _40173_, _40174_, _40175_, _40176_, _40177_, _40178_, _40179_, _40180_, _40181_, _40182_, _40183_, _40184_, _40185_, _40186_, _40187_, _40188_, _40189_, _40190_, _40191_, _40192_, _40193_, _40194_, _40195_, _40196_, _40197_, _40198_, _40199_, _40200_, _40201_, _40202_, _40203_, _40204_, _40205_, _40206_, _40207_, _40208_, _40209_, _40210_, _40211_, _40212_, _40213_, _40214_, _40215_, _40216_, _40217_, _40218_, _40219_, _40220_, _40221_, _40222_, _40223_, _40224_, _40225_, _40226_, _40227_, _40228_, _40229_, _40230_, _40231_, _40232_, _40233_, _40234_, _40235_, _40236_, _40237_, _40238_, _40239_, _40240_, _40241_, _40242_, _40243_, _40244_, _40245_, _40246_, _40247_, _40248_, _40249_, _40250_, _40251_, _40252_, _40253_, _40254_, _40255_, _40256_, _40257_, _40258_, _40259_, _40260_, _40261_, _40262_, _40263_, _40264_, _40265_, _40266_, _40267_, _40268_, _40269_, _40270_, _40271_, _40272_, _40273_, _40274_, _40275_, _40276_, _40277_, _40278_, _40279_, _40280_, _40281_, _40282_, _40283_, _40284_, _40285_, _40286_, _40287_, _40288_, _40289_, _40290_, _40291_, _40292_, _40293_, _40294_, _40295_, _40296_, _40297_, _40298_, _40299_, _40300_, _40301_, _40302_, _40303_, _40304_, _40305_, _40306_, _40307_, _40308_, _40309_, _40310_, _40311_, _40312_, _40313_, _40314_, _40315_, _40316_, _40317_, _40318_, _40319_, _40320_, _40321_, _40322_, _40323_, _40324_, _40325_, _40326_, _40327_, _40328_, _40329_, _40330_, _40331_, _40332_, _40333_, _40334_, _40335_, _40336_, _40337_, _40338_, _40339_, _40340_, _40341_, _40342_, _40343_, _40344_, _40345_, _40346_, _40347_, _40348_, _40349_, _40350_, _40351_, _40352_, _40353_, _40354_, _40355_, _40356_, _40357_, _40358_, _40359_, _40360_, _40361_, _40362_, _40363_, _40364_, _40365_, _40366_, _40367_, _40368_, _40369_, _40370_, _40371_, _40372_, _40373_, _40374_, _40375_, _40376_, _40377_, _40378_, _40379_, _40380_, _40381_, _40382_, _40383_, _40384_, _40385_, _40386_, _40387_, _40388_, _40389_, _40390_, _40391_, _40392_, _40393_, _40394_, _40395_, _40396_, _40397_, _40398_, _40399_, _40400_, _40401_, _40402_, _40403_, _40404_, _40405_, _40406_, _40407_, _40408_, _40409_, _40410_, _40411_, _40412_, _40413_, _40414_, _40415_, _40416_, _40417_, _40418_, _40419_, _40420_, _40421_, _40422_, _40423_, _40424_, _40425_, _40426_, _40427_, _40428_, _40429_, _40430_, _40431_, _40432_, _40433_, _40434_, _40435_, _40436_, _40437_, _40438_, _40439_, _40440_, _40441_, _40442_, _40443_, _40444_, _40445_, _40446_, _40447_, _40448_, _40449_, _40450_, _40451_, _40452_, _40453_, _40454_, _40455_, _40456_, _40457_, _40458_, _40459_, _40460_, _40461_, _40462_, _40463_, _40464_, _40465_, _40466_, _40467_, _40468_, _40469_, _40470_, _40471_, _40472_, _40473_, _40474_, _40475_, _40476_, _40477_, _40478_, _40479_, _40480_, _40481_, _40482_, _40483_, _40484_, _40485_, _40486_, _40487_, _40488_, _40489_, _40490_, _40491_, _40492_, _40493_, _40494_, _40495_, _40496_, _40497_, _40498_, _40499_, _40500_, _40501_, _40502_, _40503_, _40504_, _40505_, _40506_, _40507_, _40508_, _40509_, _40510_, _40511_, _40512_, _40513_, _40514_, _40515_, _40516_, _40517_, _40518_, _40519_, _40520_, _40521_, _40522_, _40523_, _40524_, _40525_, _40526_, _40527_, _40528_, _40529_, _40530_, _40531_, _40532_, _40533_, _40534_, _40535_, _40536_, _40537_, _40538_, _40539_, _40540_, _40541_, _40542_, _40543_, _40544_, _40545_, _40546_, _40547_, _40548_, _40549_, _40550_, _40551_, _40552_, _40553_, _40554_, _40555_, _40556_, _40557_, _40558_, _40559_, _40560_, _40561_, _40562_, _40563_, _40564_, _40565_, _40566_, _40567_, _40568_, _40569_, _40570_, _40571_, _40572_, _40573_, _40574_, _40575_, _40576_, _40577_, _40578_, _40579_, _40580_, _40581_, _40582_, _40583_, _40584_, _40585_, _40586_, _40587_, _40588_, _40589_, _40590_, _40591_, _40592_, _40593_, _40594_, _40595_, _40596_, _40597_, _40598_, _40599_, _40600_, _40601_, _40602_, _40603_, _40604_, _40605_, _40606_, _40607_, _40608_, _40609_, _40610_, _40611_, _40612_, _40613_, _40614_, _40615_, _40616_, _40617_, _40618_, _40619_, _40620_, _40621_, _40622_, _40623_, _40624_, _40625_, _40626_, _40627_, _40628_, _40629_, _40630_, _40631_, _40632_, _40633_, _40634_, _40635_, _40636_, _40637_, _40638_, _40639_, _40640_, _40641_, _40642_, _40643_, _40644_, _40645_, _40646_, _40647_, _40648_, _40649_, _40650_, _40651_, _40652_, _40653_, _40654_, _40655_, _40656_, _40657_, _40658_, _40659_, _40660_, _40661_, _40662_, _40663_, _40664_, _40665_, _40666_, _40667_, _40668_, _40669_, _40670_, _40671_, _40672_, _40673_, _40674_, _40675_, _40676_, _40677_, _40678_, _40679_, _40680_, _40681_, _40682_, _40683_, _40684_, _40685_, _40686_, _40687_, _40688_, _40689_, _40690_, _40691_, _40692_, _40693_, _40694_, _40695_, _40696_, _40697_, _40698_, _40699_, _40700_, _40701_, _40702_, _40703_, _40704_, _40705_, _40706_, _40707_, _40708_, _40709_, _40710_, _40711_, _40712_, _40713_, _40714_, _40715_, _40716_, _40717_, _40718_, _40719_, _40720_, _40721_, _40722_, _40723_, _40724_, _40725_, _40726_, _40727_, _40728_, _40729_, _40730_, _40731_, _40732_, _40733_, _40734_, _40735_, _40736_, _40737_, _40738_, _40739_, _40740_, _40741_, _40742_, _40743_, _40744_, _40745_, _40746_, _40747_, _40748_, _40749_, _40750_, _40751_, _40752_, _40753_, _40754_, _40755_, _40756_, _40757_, _40758_, _40759_, _40760_, _40761_, _40762_, _40763_, _40764_, _40765_, _40766_, _40767_, _40768_, _40769_, _40770_, _40771_, _40772_, _40773_, _40774_, _40775_, _40776_, _40777_, _40778_, _40779_, _40780_, _40781_, _40782_, _40783_, _40784_, _40785_, _40786_, _40787_, _40788_, _40789_, _40790_, _40791_, _40792_, _40793_, _40794_, _40795_, _40796_, _40797_, _40798_, _40799_, _40800_, _40801_, _40802_, _40803_, _40804_, _40805_, _40806_, _40807_, _40808_, _40809_, _40810_, _40811_, _40812_, _40813_, _40814_, _40815_, _40816_, _40817_, _40818_, _40819_, _40820_, _40821_, _40822_, _40823_, _40824_, _40825_, _40826_, _40827_, _40828_, _40829_, _40830_, _40831_, _40832_, _40833_, _40834_, _40835_, _40836_, _40837_, _40838_, _40839_, _40840_, _40841_, _40842_, _40843_, _40844_, _40845_, _40846_, _40847_, _40848_, _40849_, _40850_, _40851_, _40852_, _40853_, _40854_, _40855_, _40856_, _40857_, _40858_, _40859_, _40860_, _40861_, _40862_, _40863_, _40864_, _40865_, _40866_, _40867_, _40868_, _40869_, _40870_, _40871_, _40872_, _40873_, _40874_, _40875_, _40876_, _40877_, _40878_, _40879_, _40880_, _40881_, _40882_, _40883_, _40884_, _40885_, _40886_, _40887_, _40888_, _40889_, _40890_, _40891_, _40892_, _40893_, _40894_, _40895_, _40896_, _40897_, _40898_, _40899_, _40900_, _40901_, _40902_, _40903_, _40904_, _40905_, _40906_, _40907_, _40908_, _40909_, _40910_, _40911_, _40912_, _40913_, _40914_, _40915_, _40916_, _40917_, _40918_, _40919_, _40920_, _40921_, _40922_, _40923_, _40924_, _40925_, _40926_, _40927_, _40928_, _40929_, _40930_, _40931_, _40932_, _40933_, _40934_, _40935_, _40936_, _40937_, _40938_, _40939_, _40940_, _40941_, _40942_, _40943_, _40944_, _40945_, _40946_, _40947_, _40948_, _40949_, _40950_, _40951_, _40952_, _40953_, _40954_, _40955_, _40956_, _40957_, _40958_, _40959_, _40960_, _40961_, _40962_, _40963_, _40964_, _40965_, _40966_, _40967_, _40968_, _40969_, _40970_, _40971_, _40972_, _40973_, _40974_, _40975_, _40976_, _40977_, _40978_, _40979_, _40980_, _40981_, _40982_, _40983_, _40984_, _40985_, _40986_, _40987_, _40988_, _40989_, _40990_, _40991_, _40992_, _40993_, _40994_, _40995_, _40996_, _40997_, _40998_, _40999_, _41000_, _41001_, _41002_, _41003_, _41004_, _41005_, _41006_, _41007_, _41008_, _41009_, _41010_, _41011_, _41012_, _41013_, _41014_, _41015_, _41016_, _41017_, _41018_, _41019_, _41020_, _41021_, _41022_, _41023_, _41024_, _41025_, _41026_, _41027_, _41028_, _41029_, _41030_, _41031_, _41032_, _41033_, _41034_, _41035_, _41036_, _41037_, _41038_, _41039_, _41040_, _41041_, _41042_, _41043_, _41044_, _41045_, _41046_, _41047_, _41048_, _41049_, _41050_, _41051_, _41052_, _41053_, _41054_, _41055_, _41056_, _41057_, _41058_, _41059_, _41060_, _41061_, _41062_, _41063_, _41064_, _41065_, _41066_, _41067_, _41068_, _41069_, _41070_, _41071_, _41072_, _41073_, _41074_, _41075_, _41076_, _41077_, _41078_, _41079_, _41080_, _41081_, _41082_, _41083_, _41084_, _41085_, _41086_, _41087_, _41088_, _41089_, _41090_, _41091_, _41092_, _41093_, _41094_, _41095_, _41096_, _41097_, _41098_, _41099_, _41100_, _41101_, _41102_, _41103_, _41104_, _41105_, _41106_, _41107_, _41108_, _41109_, _41110_, _41111_, _41112_, _41113_, _41114_, _41115_, _41116_, _41117_, _41118_, _41119_, _41120_, _41121_, _41122_, _41123_, _41124_, _41125_, _41126_, _41127_, _41128_, _41129_, _41130_, _41131_, _41132_, _41133_, _41134_, _41135_, _41136_, _41137_, _41138_, _41139_, _41140_, _41141_, _41142_, _41143_, _41144_, _41145_, _41146_, _41147_, _41148_, _41149_, _41150_, _41151_, _41152_, _41153_, _41154_, _41155_, _41156_, _41157_, _41158_, _41159_, _41160_, _41161_, _41162_, _41163_, _41164_, _41165_, _41166_, _41167_, _41168_, _41169_, _41170_, _41171_, _41172_, _41173_, _41174_, _41175_, _41176_, _41177_, _41178_, _41179_, _41180_, _41181_, _41182_, _41183_, _41184_, _41185_, _41186_, _41187_, _41188_, _41189_, _41190_, _41191_, _41192_, _41193_, _41194_, _41195_, _41196_, _41197_, _41198_, _41199_, _41200_, _41201_, _41202_, _41203_, _41204_, _41205_, _41206_, _41207_, _41208_, _41209_, _41210_, _41211_, _41212_, _41213_, _41214_, _41215_, _41216_, _41217_, _41218_, _41219_, _41220_, _41221_, _41222_, _41223_, _41224_, _41225_, _41226_, _41227_, _41228_, _41229_, _41230_, _41231_, _41232_, _41233_, _41234_, _41235_, _41236_, _41237_, _41238_, _41239_, _41240_, _41241_, _41242_, _41243_, _41244_, _41245_, _41246_, _41247_, _41248_, _41249_, _41250_, _41251_, _41252_, _41253_, _41254_, _41255_, _41256_, _41257_, _41258_, _41259_, _41260_, _41261_, _41262_, _41263_, _41264_, _41265_, _41266_, _41267_, _41268_, _41269_, _41270_, _41271_, _41272_, _41273_, _41274_, _41275_, _41276_, _41277_, _41278_, _41279_, _41280_, _41281_, _41282_, _41283_, _41284_, _41285_, _41286_, _41287_, _41288_, _41289_, _41290_, _41291_, _41292_, _41293_, _41294_, _41295_, _41296_, _41297_, _41298_, _41299_, _41300_, _41301_, _41302_, _41303_, _41304_, _41305_, _41306_, _41307_, _41308_, _41309_, _41310_, _41311_, _41312_, _41313_, _41314_, _41315_, _41316_, _41317_, _41318_, _41319_, _41320_, _41321_, _41322_, _41323_, _41324_, _41325_, _41326_, _41327_, _41328_, _41329_, _41330_, _41331_, _41332_, _41333_, _41334_, _41335_, _41336_, _41337_, _41338_, _41339_, _41340_, _41341_, _41342_, _41343_, _41344_, _41345_, _41346_, _41347_, _41348_, _41349_, _41350_, _41351_, _41352_, _41353_, _41354_, _41355_, _41356_, _41357_, _41358_, _41359_, _41360_, _41361_, _41362_, _41363_, _41364_, _41365_, _41366_, _41367_, _41368_, _41369_, _41370_, _41371_, _41372_, _41373_, _41374_, _41375_, _41376_, _41377_, _41378_, _41379_, _41380_, _41381_, _41382_, _41383_, _41384_, _41385_, _41386_, _41387_, _41388_, _41389_, _41390_, _41391_, _41392_, _41393_, _41394_, _41395_, _41396_, _41397_, _41398_, _41399_, _41400_, _41401_, _41402_, _41403_, _41404_, _41405_, _41406_, _41407_, _41408_, _41409_, _41410_, _41411_, _41412_, _41413_, _41414_, _41415_, _41416_, _41417_, _41418_, _41419_, _41420_, _41421_, _41422_, _41423_, _41424_, _41425_, _41426_, _41427_, _41428_, _41429_, _41430_, _41431_, _41432_, _41433_, _41434_, _41435_, _41436_, _41437_, _41438_, _41439_, _41440_, _41441_, _41442_, _41443_, _41444_, _41445_, _41446_, _41447_, _41448_, _41449_, _41450_, _41451_, _41452_, _41453_, _41454_, _41455_, _41456_, _41457_, _41458_, _41459_, _41460_, _41461_, _41462_, _41463_, _41464_, _41465_, _41466_, _41467_, _41468_, _41469_, _41470_, _41471_, _41472_, _41473_, _41474_, _41475_, _41476_, _41477_, _41478_, _41479_, _41480_, _41481_, _41482_, _41483_, _41484_, _41485_, _41486_, _41487_, _41488_, _41489_, _41490_, _41491_, _41492_, _41493_, _41494_, _41495_, _41496_, _41497_, _41498_, _41499_, _41500_, _41501_, _41502_, _41503_, _41504_, _41505_, _41506_, _41507_, _41508_, _41509_, _41510_, _41511_, _41512_, _41513_, _41514_, _41515_, _41516_, _41517_, _41518_, _41519_, _41520_, _41521_, _41522_, _41523_, _41524_, _41525_, _41526_, _41527_, _41528_, _41529_, _41530_, _41531_, _41532_, _41533_, _41534_, _41535_, _41536_, _41537_, _41538_, _41539_, _41540_, _41541_, _41542_, _41543_, _41544_, _41545_, _41546_, _41547_, _41548_, _41549_, _41550_, _41551_, _41552_, _41553_, _41554_, _41555_, _41556_, _41557_, _41558_, _41559_, _41560_, _41561_, _41562_, _41563_, _41564_, _41565_, _41566_, _41567_, _41568_, _41569_, _41570_, _41571_, _41572_, _41573_, _41574_, _41575_, _41576_, _41577_, _41578_, _41579_, _41580_, _41581_, _41582_, _41583_, _41584_, _41585_, _41586_, _41587_, _41588_, _41589_, _41590_, _41591_, _41592_, _41593_, _41594_, _41595_, _41596_, _41597_, _41598_, _41599_, _41600_, _41601_, _41602_, _41603_, _41604_, _41605_, _41606_, _41607_, _41608_, _41609_, _41610_, _41611_, _41612_, _41613_, _41614_, _41615_, _41616_, _41617_, _41618_, _41619_, _41620_, _41621_, _41622_, _41623_, _41624_, _41625_, _41626_, _41627_, _41628_, _41629_, _41630_, _41631_, _41632_, _41633_, _41634_, _41635_, _41636_, _41637_, _41638_, _41639_, _41640_, _41641_, _41642_, _41643_, _41644_, _41645_, _41646_, _41647_, _41648_, _41649_, _41650_, _41651_, _41652_, _41653_, _41654_, _41655_, _41656_, _41657_, _41658_, _41659_, _41660_, _41661_, _41662_, _41663_, _41664_, _41665_, _41666_, _41667_, _41668_, _41669_, _41670_, _41671_, _41672_, _41673_, _41674_, _41675_, _41676_, _41677_, _41678_, _41679_, _41680_, _41681_, _41682_, _41683_, _41684_, _41685_, _41686_, _41687_, _41688_, _41689_, _41690_, _41691_, _41692_, _41693_, _41694_, _41695_, _41696_, _41697_, _41698_, _41699_, _41700_, _41701_, _41702_, _41703_, _41704_, _41705_, _41706_, _41707_, _41708_, _41709_, _41710_, _41711_, _41712_, _41713_, _41714_, _41715_, _41716_, _41717_, _41718_, _41719_, _41720_, _41721_, _41722_, _41723_, _41724_, _41725_, _41726_, _41727_, _41728_, _41729_, _41730_, _41731_, _41732_, _41733_, _41734_, _41735_, _41736_, _41737_, _41738_, _41739_, _41740_, _41741_, _41742_, _41743_, _41744_, _41745_, _41746_, _41747_, _41748_, _41749_, _41750_, _41751_, _41752_, _41753_, _41754_, _41755_, _41756_, _41757_, _41758_, _41759_, _41760_, _41761_, _41762_, _41763_, _41764_, _41765_, _41766_, _41767_, _41768_, _41769_, _41770_, _41771_, _41772_, _41773_, _41774_, _41775_, _41776_, _41777_, _41778_, _41779_, _41780_, _41781_, _41782_, _41783_, _41784_, _41785_, _41786_, _41787_, _41788_, _41789_, _41790_, _41791_, _41792_, _41793_, _41794_, _41795_, _41796_, _41797_, _41798_, _41799_, _41800_, _41801_, _41802_, _41803_, _41804_, _41805_, _41806_, _41807_, _41808_, _41809_, _41810_, _41811_, _41812_, _41813_, _41814_, _41815_, _41816_, _41817_, _41818_, _41819_, _41820_, _41821_, _41822_, _41823_, _41824_, _41825_, _41826_, _41827_, _41828_, _41829_, _41830_, _41831_, _41832_, _41833_, _41834_, _41835_, _41836_, _41837_, _41838_, _41839_, _41840_, _41841_, _41842_, _41843_, _41844_, _41845_, _41846_, _41847_, _41848_, _41849_, _41850_, _41851_, _41852_, _41853_, _41854_, _41855_, _41856_, _41857_, _41858_, _41859_, _41860_, _41861_, _41862_, _41863_, _41864_, _41865_, _41866_, _41867_, _41868_, _41869_, _41870_, _41871_, _41872_, _41873_, _41874_, _41875_, _41876_, _41877_, _41878_, _41879_, _41880_, _41881_, _41882_, _41883_, _41884_, _41885_, _41886_, _41887_, _41888_, _41889_, _41890_, _41891_, _41892_, _41893_, _41894_, _41895_, _41896_, _41897_, _41898_, _41899_, _41900_, _41901_, _41902_, _41903_, _41904_, _41905_, _41906_, _41907_, _41908_, _41909_, _41910_, _41911_, _41912_, _41913_, _41914_, _41915_, _41916_, _41917_, _41918_, _41919_, _41920_, _41921_, _41922_, _41923_, _41924_, _41925_, _41926_, _41927_, _41928_, _41929_, _41930_, _41931_, _41932_, _41933_, _41934_, _41935_, _41936_, _41937_, _41938_, _41939_, _41940_, _41941_, _41942_, _41943_, _41944_, _41945_, _41946_, _41947_, _41948_, _41949_, _41950_, _41951_, _41952_, _41953_, _41954_, _41955_, _41956_, _41957_, _41958_, _41959_, _41960_, _41961_, _41962_, _41963_, _41964_, _41965_, _41966_, _41967_, _41968_, _41969_, _41970_, _41971_, _41972_, _41973_, _41974_, _41975_, _41976_, _41977_, _41978_, _41979_, _41980_, _41981_, _41982_, _41983_, _41984_, _41985_, _41986_, _41987_, _41988_, _41989_, _41990_, _41991_, _41992_, _41993_, _41994_, _41995_, _41996_, _41997_, _41998_, _41999_, _42000_, _42001_, _42002_, _42003_, _42004_, _42005_, _42006_, _42007_, _42008_, _42009_, _42010_, _42011_, _42012_, _42013_, _42014_, _42015_, _42016_, _42017_, _42018_, _42019_, _42020_, _42021_, _42022_, _42023_, _42024_, _42025_, _42026_, _42027_, _42028_, _42029_, _42030_, _42031_, _42032_, _42033_, _42034_, _42035_, _42036_, _42037_, _42038_, _42039_, _42040_, _42041_, _42042_, _42043_, _42044_, _42045_, _42046_, _42047_, _42048_, _42049_, _42050_, _42051_, _42052_, _42053_, _42054_, _42055_, _42056_, _42057_, _42058_, _42059_, _42060_, _42061_, _42062_, _42063_, _42064_, _42065_, _42066_, _42067_, _42068_, _42069_, _42070_, _42071_, _42072_, _42073_, _42074_, _42075_, _42076_, _42077_, _42078_, _42079_, _42080_, _42081_, _42082_, _42083_, _42084_, _42085_, _42086_, _42087_, _42088_, _42089_, _42090_, _42091_, _42092_, _42093_, _42094_, _42095_, _42096_, _42097_, _42098_, _42099_, _42100_, _42101_, _42102_, _42103_, _42104_, _42105_, _42106_, _42107_, _42108_, _42109_, _42110_, _42111_, _42112_, _42113_, _42114_, _42115_, _42116_, _42117_, _42118_, _42119_, _42120_, _42121_, _42122_, _42123_, _42124_, _42125_, _42126_, _42127_, _42128_, _42129_, _42130_, _42131_, _42132_, _42133_, _42134_, _42135_, _42136_, _42137_, _42138_, _42139_, _42140_, _42141_, _42142_, _42143_, _42144_, _42145_, _42146_, _42147_, _42148_, _42149_, _42150_, _42151_, _42152_, _42153_, _42154_, _42155_, _42156_, _42157_, _42158_, _42159_, _42160_, _42161_, _42162_, _42163_, _42164_, _42165_, _42166_, _42167_, _42168_, _42169_, _42170_, _42171_, _42172_, _42173_, _42174_, _42175_, _42176_, _42177_, _42178_, _42179_, _42180_, _42181_, _42182_, _42183_, _42184_, _42185_, _42186_, _42187_, _42188_, _42189_, _42190_, _42191_, _42192_, _42193_, _42194_, _42195_, _42196_, _42197_, _42198_, _42199_, _42200_, _42201_, _42202_, _42203_, _42204_, _42205_, _42206_, _42207_, _42208_, _42209_, _42210_, _42211_, _42212_, _42213_, _42214_, _42215_, _42216_, _42217_, _42218_, _42219_, _42220_, _42221_, _42222_, _42223_, _42224_, _42225_, _42226_, _42227_, _42228_, _42229_, _42230_, _42231_, _42232_, _42233_, _42234_, _42235_, _42236_, _42237_, _42238_, _42239_, _42240_, _42241_, _42242_, _42243_, _42244_, _42245_, _42246_, _42247_, _42248_, _42249_, _42250_, _42251_, _42252_, _42253_, _42254_, _42255_, _42256_, _42257_, _42258_, _42259_, _42260_, _42261_, _42262_, _42263_, _42264_, _42265_, _42266_, _42267_, _42268_, _42269_, _42270_, _42271_, _42272_, _42273_, _42274_, _42275_, _42276_, _42277_, _42278_, _42279_, _42280_, _42281_, _42282_, _42283_, _42284_, _42285_, _42286_, _42287_, _42288_, _42289_, _42290_, _42291_, _42292_, _42293_, _42294_, _42295_, _42296_, _42297_, _42298_, _42299_, _42300_, _42301_, _42302_, _42303_, _42304_, _42305_, _42306_, _42307_, _42308_, _42309_, _42310_, _42311_, _42312_, _42313_, _42314_, _42315_, _42316_, _42317_, _42318_, _42319_, _42320_, _42321_, _42322_, _42323_, _42324_, _42325_, _42326_, _42327_, _42328_, _42329_, _42330_, _42331_, _42332_, _42333_, _42334_, _42335_, _42336_, _42337_, _42338_, _42339_, _42340_, _42341_, _42342_, _42343_, _42344_, _42345_, _42346_, _42347_, _42348_, _42349_, _42350_, _42351_, _42352_, _42353_, _42354_, _42355_, _42356_, _42357_, _42358_, _42359_, _42360_, _42361_, _42362_, _42363_, _42364_, _42365_, _42366_, _42367_, _42368_, _42369_, _42370_, _42371_, _42372_, _42373_, _42374_, _42375_, _42376_, _42377_, _42378_, _42379_, _42380_, _42381_, _42382_, _42383_, _42384_, _42385_, _42386_, _42387_, _42388_, _42389_, _42390_, _42391_, _42392_, _42393_, _42394_, _42395_, _42396_, _42397_, _42398_, _42399_, _42400_, _42401_, _42402_, _42403_, _42404_, _42405_, _42406_, _42407_, _42408_, _42409_, _42410_, _42411_, _42412_, _42413_, _42414_, _42415_, _42416_, _42417_, _42418_, _42419_, _42420_, _42421_, _42422_, _42423_, _42424_, _42425_, _42426_, _42427_, _42428_, _42429_, _42430_, _42431_, _42432_, _42433_, _42434_, _42435_, _42436_, _42437_, _42438_, _42439_, _42440_, _42441_, _42442_, _42443_, _42444_, _42445_, _42446_, _42447_, _42448_, _42449_, _42450_, _42451_, _42452_, _42453_, _42454_, _42455_, _42456_, _42457_, _42458_, _42459_, _42460_, _42461_, _42462_, _42463_, _42464_, _42465_, _42466_, _42467_, _42468_, _42469_, _42470_, _42471_, _42472_, _42473_, _42474_, _42475_, _42476_, _42477_, _42478_, _42479_, _42480_, _42481_, _42482_, _42483_, _42484_, _42485_, _42486_, _42487_, _42488_, _42489_, _42490_, _42491_, _42492_, _42493_, _42494_, _42495_, _42496_, _42497_, _42498_, _42499_, _42500_, _42501_, _42502_, _42503_, _42504_, _42505_, _42506_, _42507_, _42508_, _42509_, _42510_, _42511_, _42512_, _42513_, _42514_, _42515_, _42516_, _42517_, _42518_, _42519_, _42520_, _42521_, _42522_, _42523_, _42524_, _42525_, _42526_, _42527_, _42528_, _42529_, _42530_, _42531_, _42532_, _42533_, _42534_, _42535_, _42536_, _42537_, _42538_, _42539_, _42540_, _42541_, _42542_, _42543_, _42544_, _42545_, _42546_, _42547_, _42548_, _42549_, _42550_, _42551_, _42552_, _42553_, _42554_, _42555_, _42556_, _42557_, _42558_, _42559_, _42560_, _42561_, _42562_, _42563_, _42564_, _42565_, _42566_, _42567_, _42568_, _42569_, _42570_, _42571_, _42572_, _42573_, _42574_, _42575_, _42576_, _42577_, _42578_, _42579_, _42580_, _42581_, _42582_, _42583_, _42584_, _42585_, _42586_, _42587_, _42588_, _42589_, _42590_, _42591_, _42592_, _42593_, _42594_, _42595_, _42596_, _42597_, _42598_, _42599_, _42600_, _42601_, _42602_, _42603_, _42604_, _42605_, _42606_, _42607_, _42608_, _42609_, _42610_, _42611_, _42612_, _42613_, _42614_, _42615_, _42616_, _42617_, _42618_, _42619_, _42620_, _42621_, _42622_, _42623_, _42624_, _42625_, _42626_, _42627_, _42628_, _42629_, _42630_, _42631_, _42632_, _42633_, _42634_, _42635_, _42636_, _42637_, _42638_, _42639_, _42640_, _42641_, _42642_, _42643_, _42644_, _42645_, _42646_, _42647_, _42648_, _42649_, _42650_, _42651_, _42652_, _42653_, _42654_, _42655_, _42656_, _42657_, _42658_, _42659_, _42660_, _42661_, _42662_, _42663_, _42664_, _42665_, _42666_, _42667_, _42668_, _42669_, _42670_, _42671_, _42672_, _42673_, _42674_, _42675_, _42676_, _42677_, _42678_, _42679_, _42680_, _42681_, _42682_, _42683_, _42684_, _42685_, _42686_, _42687_, _42688_, _42689_, _42690_, _42691_, _42692_, _42693_, _42694_, _42695_, _42696_, _42697_, _42698_, _42699_, _42700_, _42701_, _42702_, _42703_, _42704_, _42705_, _42706_, _42707_, _42708_, _42709_, _42710_, _42711_, _42712_, _42713_, _42714_, _42715_, _42716_, _42717_, _42718_, _42719_, _42720_, _42721_, _42722_, _42723_, _42724_, _42725_, _42726_, _42727_, _42728_, _42729_, _42730_, _42731_, _42732_, _42733_, _42734_, _42735_, _42736_, _42737_, _42738_, _42739_, _42740_, _42741_, _42742_, _42743_, _42744_, _42745_, _42746_, _42747_, _42748_, _42749_, _42750_, _42751_, _42752_, _42753_, _42754_, _42755_, _42756_, _42757_, _42758_, _42759_, _42760_, _42761_, _42762_, _42763_, _42764_, _42765_, _42766_, _42767_, _42768_, _42769_, _42770_, _42771_, _42772_, _42773_, _42774_, _42775_, _42776_, _42777_, _42778_, _42779_, _42780_, _42781_, _42782_, _42783_, _42784_, _42785_, _42786_, _42787_, _42788_, _42789_, _42790_, _42791_, _42792_, _42793_, _42794_, _42795_, _42796_, _42797_, _42798_, _42799_, _42800_, _42801_, _42802_, _42803_, _42804_, _42805_, _42806_, _42807_, _42808_, _42809_, _42810_, _42811_, _42812_, _42813_, _42814_, _42815_, _42816_, _42817_, _42818_, _42819_, _42820_, _42821_, _42822_, _42823_, _42824_, _42825_, _42826_, _42827_, _42828_, _42829_, _42830_, _42831_, _42832_, _42833_, _42834_, _42835_, _42836_, _42837_, _42838_, _42839_, _42840_, _42841_, _42842_, _42843_, _42844_, _42845_, _42846_, _42847_, _42848_, _42849_, _42850_, _42851_, _42852_, _42853_, _42854_, _42855_, _42856_, _42857_, _42858_, _42859_, _42860_, _42861_, _42862_, _42863_, _42864_, _42865_, _42866_, _42867_, _42868_, _42869_, _42870_, _42871_, _42872_, _42873_, _42874_, _42875_, _42876_, _42877_, _42878_, _42879_, _42880_, _42881_, _42882_, _42883_, _42884_, _42885_, _42886_, _42887_, _42888_, _42889_, _42890_, _42891_, _42892_, _42893_, _42894_, _42895_, _42896_, _42897_, _42898_, _42899_, _42900_, _42901_, _42902_, _42903_, _42904_, _42905_, _42906_, _42907_, _42908_, _42909_, _42910_, _42911_, _42912_, _42913_, _42914_, _42915_, _42916_, _42917_, _42918_, _42919_, _42920_, _42921_, _42922_, _42923_, _42924_, _42925_, _42926_, _42927_, _42928_, _42929_, _42930_, _42931_, _42932_, _42933_, _42934_, _42935_, _42936_, _42937_, _42938_, _42939_, _42940_, _42941_, _42942_, _42943_, _42944_, _42945_, _42946_, _42947_, _42948_, _42949_, _42950_, _42951_, _42952_, _42953_, _42954_, _42955_, _42956_, _42957_, _42958_, _42959_, _42960_, _42961_, _42962_, _42963_, _42964_, _42965_, _42966_, _42967_, _42968_, _42969_, _42970_, _42971_, _42972_, _42973_, _42974_, _42975_, _42976_, _42977_, _42978_, _42979_, _42980_, _42981_, _42982_, _42983_, _42984_, _42985_, _42986_, _42987_, _42988_, _42989_, _42990_, _42991_, _42992_, _42993_, _42994_, _42995_, _42996_, _42997_, _42998_, _42999_, _43000_, _43001_, _43002_, _43003_, _43004_, _43005_, _43006_, _43007_, _43008_, _43009_, _43010_, _43011_, _43012_, _43013_, _43014_, _43015_, _43016_, _43017_, _43018_, _43019_, _43020_, _43021_, _43022_, _43023_, _43024_, _43025_, _43026_, _43027_, _43028_, _43029_, _43030_, _43031_, _43032_, _43033_, _43034_, _43035_, _43036_, _43037_, _43038_, _43039_, _43040_, _43041_, _43042_, _43043_, _43044_, _43045_, _43046_, _43047_, _43048_, _43049_, _43050_, _43051_, _43052_, _43053_, _43054_, _43055_, _43056_, _43057_, _43058_, _43059_, _43060_, _43061_, _43062_, _43063_, _43064_, _43065_, _43066_, _43067_, _43068_, _43069_, _43070_, _43071_, _43072_, _43073_, _43074_, _43075_, _43076_, _43077_, _43078_, _43079_, _43080_, _43081_, _43082_, _43083_, _43084_, _43085_, _43086_, _43087_, _43088_, _43089_, _43090_, _43091_, _43092_, _43093_, _43094_, _43095_, _43096_, _43097_, _43098_, _43099_, _43100_, _43101_, _43102_, _43103_, _43104_, _43105_, _43106_, _43107_, _43108_, _43109_, _43110_, _43111_, _43112_, _43113_, _43114_, _43115_, _43116_, _43117_, _43118_, _43119_, _43120_, _43121_, _43122_, _43123_, _43124_, _43125_, _43126_, _43127_, _43128_, _43129_, _43130_, _43131_, _43132_, _43133_, _43134_, _43135_, _43136_, _43137_, _43138_, _43139_, _43140_, _43141_, _43142_, _43143_, _43144_, _43145_, _43146_, _43147_, _43148_, _43149_, _43150_, _43151_, _43152_, _43153_, _43154_, _43155_, _43156_, _43157_, _43158_, _43159_, _43160_, _43161_, _43162_, _43163_, _43164_, _43165_, _43166_, _43167_, _43168_, _43169_, _43170_, _43171_, _43172_, _43173_, _43174_, _43175_, _43176_, _43177_, _43178_, _43179_, _43180_, _43181_, _43182_, _43183_, _43184_, _43185_, _43186_, _43187_, _43188_, _43189_, _43190_, _43191_, _43192_, _43193_, _43194_, _43195_, _43196_, _43197_, _43198_, _43199_, _43200_, _43201_, _43202_, _43203_, _43204_, _43205_, _43206_, _43207_, _43208_, _43209_, _43210_, _43211_, _43212_, _43213_, _43214_, _43215_, _43216_, _43217_, _43218_, _43219_, _43220_, _43221_, _43222_, _43223_, _43224_, _43225_, _43226_, _43227_, _43228_, _43229_, _43230_, _43231_, _43232_, _43233_, _43234_, _43235_, _43236_, _43237_, _43238_, _43239_, _43240_, _43241_, _43242_, _43243_, _43244_, _43245_, _43246_, _43247_, _43248_, _43249_, _43250_, _43251_, _43252_, _43253_, _43254_, _43255_, _43256_, _43257_, _43258_, _43259_, _43260_, _43261_, _43262_, _43263_, _43264_, _43265_, _43266_, _43267_, _43268_, _43269_, _43270_, _43271_, _43272_, _43273_, _43274_, _43275_, _43276_, _43277_, _43278_, _43279_, _43280_, _43281_, _43282_, _43283_, _43284_, _43285_, _43286_, _43287_, _43288_, _43289_, _43290_, _43291_, _43292_, _43293_, _43294_, _43295_, _43296_, _43297_, _43298_, _43299_, _43300_, _43301_, _43302_, _43303_, _43304_, _43305_, _43306_, _43307_, _43308_, _43309_, _43310_, _43311_, _43312_, _43313_, _43314_, _43315_, _43316_, _43317_, _43318_, _43319_, _43320_, _43321_, _43322_, _43323_, _43324_, _43325_, _43326_, _43327_, _43328_, _43329_, _43330_, _43331_, _43332_, _43333_, _43334_, _43335_, _43336_, _43337_, _43338_, _43339_, _43340_, _43341_, _43342_, _43343_, _43344_, _43345_, _43346_, _43347_, _43348_, _43349_, _43350_, _43351_, _43352_, _43353_, _43354_, _43355_, _43356_, _43357_, _43358_, _43359_, _43360_, _43361_, _43362_, _43363_, _43364_, _43365_, _43366_, _43367_, _43368_, _43369_, _43370_, _43371_, _43372_, _43373_, _43374_, _43375_, _43376_, _43377_, _43378_, _43379_, _43380_, _43381_, _43382_, _43383_, _43384_, _43385_, _43386_, _43387_, _43388_, _43389_, _43390_, _43391_, _43392_, _43393_, _43394_, _43395_, _43396_, _43397_, _43398_, _43399_, _43400_, _43401_, _43402_, _43403_, _43404_, _43405_, _43406_, _43407_, _43408_, _43409_, _43410_, _43411_, _43412_, _43413_, _43414_, _43415_, _43416_, _43417_, _43418_, _43419_, _43420_, _43421_, _43422_, _43423_, _43424_, _43425_, _43426_, _43427_, _43428_, _43429_, _43430_, _43431_, _43432_, _43433_, _43434_, _43435_, _43436_, _43437_, _43438_, _43439_, _43440_, _43441_, _43442_, _43443_, _43444_, _43445_, _43446_, _43447_, _43448_, _43449_, _43450_, _43451_, _43452_, _43453_, _43454_, _43455_, _43456_, _43457_, _43458_, _43459_, _43460_, _43461_, _43462_, _43463_, _43464_, _43465_, _43466_, _43467_, _43468_, _43469_, _43470_, _43471_, _43472_, _43473_, _43474_, _43475_, _43476_, _43477_, _43478_, _43479_, _43480_, _43481_, _43482_, _43483_, _43484_, _43485_, _43486_, _43487_, _43488_, _43489_, _43490_, _43491_, _43492_, _43493_, _43494_, _43495_, _43496_, _43497_, _43498_, _43499_, _43500_, _43501_, _43502_, _43503_, _43504_, _43505_, _43506_, _43507_, _43508_, _43509_, _43510_, _43511_, _43512_, _43513_, _43514_, _43515_, _43516_, _43517_, _43518_, _43519_, _43520_, _43521_, _43522_, _43523_, _43524_, _43525_, _43526_, _43527_, _43528_, _43529_, _43530_, _43531_, _43532_, _43533_, _43534_, _43535_, _43536_, _43537_, _43538_, _43539_, _43540_, _43541_, _43542_, _43543_, _43544_, _43545_, _43546_, _43547_, _43548_, _43549_, _43550_, _43551_, _43552_, _43553_, _43554_, _43555_, _43556_, _43557_, _43558_, _43559_, _43560_, _43561_, _43562_, _43563_, _43564_, _43565_, _43566_, _43567_, _43568_, _43569_, _43570_, _43571_, _43572_, _43573_, _43574_, _43575_, _43576_, _43577_, _43578_, _43579_, _43580_, _43581_, _43582_, _43583_, _43584_, _43585_, _43586_, _43587_, _43588_, _43589_, _43590_, _43591_, _43592_, _43593_, _43594_, _43595_, _43596_, _43597_, _43598_, _43599_, _43600_, _43601_, _43602_, _43603_, _43604_, _43605_, _43606_, _43607_, _43608_, _43609_, _43610_, _43611_, _43612_, _43613_, _43614_, _43615_, _43616_, _43617_, _43618_, _43619_, _43620_, _43621_, _43622_, _43623_, _43624_, _43625_, _43626_, _43627_, _43628_, _43629_, _43630_, _43631_, _43632_, _43633_, _43634_, _43635_, _43636_, _43637_, _43638_, _43639_, _43640_, _43641_, _43642_, _43643_, _43644_, _43645_, _43646_, _43647_, _43648_, _43649_, _43650_, _43651_, _43652_, _43653_, _43654_, _43655_, _43656_, _43657_, _43658_, _43659_, _43660_, _43661_, _43662_, _43663_, _43664_, _43665_, _43666_, _43667_, _43668_, _43669_, _43670_, _43671_, _43672_, _43673_, _43674_, _43675_, _43676_, _43677_, _43678_, _43679_, _43680_, _43681_, _43682_, _43683_, _43684_, _43685_, _43686_, _43687_, _43688_, _43689_, _43690_, _43691_, _43692_, _43693_, _43694_, _43695_, _43696_, _43697_, _43698_, _43699_, _43700_, _43701_, _43702_, _43703_, _43704_, _43705_, _43706_, _43707_, _43708_, _43709_, _43710_, _43711_, _43712_, _43713_, _43714_, _43715_, _43716_, _43717_, _43718_, _43719_, _43720_, _43721_, _43722_, _43723_, _43724_, _43725_, _43726_, _43727_, _43728_, _43729_, _43730_, _43731_, _43732_, _43733_, _43734_, _43735_, _43736_, _43737_, _43738_, _43739_, _43740_, _43741_, _43742_, _43743_, _43744_, _43745_, _43746_, _43747_, _43748_, _43749_, _43750_, _43751_, _43752_, _43753_, _43754_, _43755_, _43756_, _43757_, _43758_, _43759_, _43760_, _43761_, _43762_, _43763_, _43764_, _43765_, _43766_, _43767_, _43768_, _43769_, _43770_, _43771_, _43772_, _43773_, _43774_, _43775_, _43776_, _43777_, _43778_, _43779_, _43780_, _43781_, _43782_, _43783_, _43784_, _43785_, _43786_, _43787_, _43788_, _43789_, _43790_, _43791_, _43792_, _43793_, , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , ;
  input [319:0] set1;
  input [319:0] set2;
  input set1[0], set1[1], set1[2], set1[3], set1[4], set1[5], set1[6], set1[7], set1[8], set1[9], set1[10], set1[11], set1[12], set1[13], set1[14], set1[15], set1[16], set1[17], set1[18], set1[19], set1[20], set1[21], set1[22], set1[23], set1[24], set1[25], set1[26], set1[27], set1[28], set1[29], set1[30], set1[31], set1[32], set1[33], set1[34], set1[35], set1[36], set1[37], set1[38], set1[39], set1[40], set1[41], set1[42], set1[43], set1[44], set1[45], set1[46], set1[47], set1[48], set1[49], set1[50], set1[51], set1[52], set1[53], set1[54], set1[55], set1[56], set1[57], set1[58], set1[59], set1[60], set1[61], set1[62], set1[63], set1[64], set1[65], set1[66], set1[67], set1[68], set1[69], set1[70], set1[71], set1[72], set1[73], set1[74], set1[75], set1[76], set1[77], set1[78], set1[79], set1[80], set1[81], set1[82], set1[83], set1[84], set1[85], set1[86], set1[87], set1[88], set1[89], set1[90], set1[91], set1[92], set1[93], set1[94], set1[95], set1[96], set1[97], set1[98], set1[99], set1[100], set1[101], set1[102], set1[103], set1[104], set1[105], set1[106], set1[107], set1[108], set1[109], set1[110], set1[111], set1[112], set1[113], set1[114], set1[115], set1[116], set1[117], set1[118], set1[119], set1[120], set1[121], set1[122], set1[123], set1[124], set1[125], set1[126], set1[127], set1[128], set1[129], set1[130], set1[131], set1[132], set1[133], set1[134], set1[135], set1[136], set1[137], set1[138], set1[139], set1[140], set1[141], set1[142], set1[143], set1[144], set1[145], set1[146], set1[147], set1[148], set1[149], set1[150], set1[151], set1[152], set1[153], set1[154], set1[155], set1[156], set1[157], set1[158], set1[159], set1[160], set1[161], set1[162], set1[163], set1[164], set1[165], set1[166], set1[167], set1[168], set1[169], set1[170], set1[171], set1[172], set1[173], set1[174], set1[175], set1[176], set1[177], set1[178], set1[179], set1[180], set1[181], set1[182], set1[183], set1[184], set1[185], set1[186], set1[187], set1[188], set1[189], set1[190], set1[191], set1[192], set1[193], set1[194], set1[195], set1[196], set1[197], set1[198], set1[199], set1[200], set1[201], set1[202], set1[203], set1[204], set1[205], set1[206], set1[207], set1[208], set1[209], set1[210], set1[211], set1[212], set1[213], set1[214], set1[215], set1[216], set1[217], set1[218], set1[219], set1[220], set1[221], set1[222], set1[223], set1[224], set1[225], set1[226], set1[227], set1[228], set1[229], set1[230], set1[231], set1[232], set1[233], set1[234], set1[235], set1[236], set1[237], set1[238], set1[239], set1[240], set1[241], set1[242], set1[243], set1[244], set1[245], set1[246], set1[247], set1[248], set1[249], set1[250], set1[251], set1[252], set1[253], set1[254], set1[255], set1[256], set1[257], set1[258], set1[259], set1[260], set1[261], set1[262], set1[263], set1[264], set1[265], set1[266], set1[267], set1[268], set1[269], set1[270], set1[271], set1[272], set1[273], set1[274], set1[275], set1[276], set1[277], set1[278], set1[279], set1[280], set1[281], set1[282], set1[283], set1[284], set1[285], set1[286], set1[287], set1[288], set1[289], set1[290], set1[291], set1[292], set1[293], set1[294], set1[295], set1[296], set1[297], set1[298], set1[299], set1[300], set1[301], set1[302], set1[303], set1[304], set1[305], set1[306], set1[307], set1[308], set1[309], set1[310], set1[311], set1[312], set1[313], set1[314], set1[315], set1[316], set1[317], set1[318], set1[319], set2[0], set2[1], set2[2], set2[3], set2[4], set2[5], set2[6], set2[7], set2[8], set2[9], set2[10], set2[11], set2[12], set2[13], set2[14], set2[15], set2[16], set2[17], set2[18], set2[19], set2[20], set2[21], set2[22], set2[23], set2[24], set2[25], set2[26], set2[27], set2[28], set2[29], set2[30], set2[31], set2[32], set2[33], set2[34], set2[35], set2[36], set2[37], set2[38], set2[39], set2[40], set2[41], set2[42], set2[43], set2[44], set2[45], set2[46], set2[47], set2[48], set2[49], set2[50], set2[51], set2[52], set2[53], set2[54], set2[55], set2[56], set2[57], set2[58], set2[59], set2[60], set2[61], set2[62], set2[63], set2[64], set2[65], set2[66], set2[67], set2[68], set2[69], set2[70], set2[71], set2[72], set2[73], set2[74], set2[75], set2[76], set2[77], set2[78], set2[79], set2[80], set2[81], set2[82], set2[83], set2[84], set2[85], set2[86], set2[87], set2[88], set2[89], set2[90], set2[91], set2[92], set2[93], set2[94], set2[95], set2[96], set2[97], set2[98], set2[99], set2[100], set2[101], set2[102], set2[103], set2[104], set2[105], set2[106], set2[107], set2[108], set2[109], set2[110], set2[111], set2[112], set2[113], set2[114], set2[115], set2[116], set2[117], set2[118], set2[119], set2[120], set2[121], set2[122], set2[123], set2[124], set2[125], set2[126], set2[127], set2[128], set2[129], set2[130], set2[131], set2[132], set2[133], set2[134], set2[135], set2[136], set2[137], set2[138], set2[139], set2[140], set2[141], set2[142], set2[143], set2[144], set2[145], set2[146], set2[147], set2[148], set2[149], set2[150], set2[151], set2[152], set2[153], set2[154], set2[155], set2[156], set2[157], set2[158], set2[159], set2[160], set2[161], set2[162], set2[163], set2[164], set2[165], set2[166], set2[167], set2[168], set2[169], set2[170], set2[171], set2[172], set2[173], set2[174], set2[175], set2[176], set2[177], set2[178], set2[179], set2[180], set2[181], set2[182], set2[183], set2[184], set2[185], set2[186], set2[187], set2[188], set2[189], set2[190], set2[191], set2[192], set2[193], set2[194], set2[195], set2[196], set2[197], set2[198], set2[199], set2[200], set2[201], set2[202], set2[203], set2[204], set2[205], set2[206], set2[207], set2[208], set2[209], set2[210], set2[211], set2[212], set2[213], set2[214], set2[215], set2[216], set2[217], set2[218], set2[219], set2[220], set2[221], set2[222], set2[223], set2[224], set2[225], set2[226], set2[227], set2[228], set2[229], set2[230], set2[231], set2[232], set2[233], set2[234], set2[235], set2[236], set2[237], set2[238], set2[239], set2[240], set2[241], set2[242], set2[243], set2[244], set2[245], set2[246], set2[247], set2[248], set2[249], set2[250], set2[251], set2[252], set2[253], set2[254], set2[255], set2[256], set2[257], set2[258], set2[259], set2[260], set2[261], set2[262], set2[263], set2[264], set2[265], set2[266], set2[267], set2[268], set2[269], set2[270], set2[271], set2[272], set2[273], set2[274], set2[275], set2[276], set2[277], set2[278], set2[279], set2[280], set2[281], set2[282], set2[283], set2[284], set2[285], set2[286], set2[287], set2[288], set2[289], set2[290], set2[291], set2[292], set2[293], set2[294], set2[295], set2[296], set2[297], set2[298], set2[299], set2[300], set2[301], set2[302], set2[303], set2[304], set2[305], set2[306], set2[307], set2[308], set2[309], set2[310], set2[311], set2[312], set2[313], set2[314], set2[315], set2[316], set2[317], set2[318], set2[319];
  output out[0], out[1], out[2], out[3], out[4], out[5], out[6], out[7], out[8], out[9], out[10], out[11], out[12], out[13], out[14], out[15], out[16], out[17], out[18], out[19], out[20], out[21], out[22], out[23], out[24], out[25], out[26], out[27], out[28], out[29], out[30], out[31], out[32], out[33], out[34], out[35], out[36], out[37], out[38], out[39], out[40], out[41], out[42], out[43], out[44], out[45], out[46], out[47], out[48], out[49], out[50], out[51], out[52], out[53], out[54], out[55], out[56], out[57], out[58], out[59], out[60], out[61], out[62], out[63], out[64], out[65], out[66], out[67], out[68], out[69], out[70], out[71], out[72], out[73], out[74], out[75], out[76], out[77], out[78], out[79], out[80], out[81], out[82], out[83], out[84], out[85], out[86], out[87], out[88], out[89], out[90], out[91], out[92], out[93], out[94], out[95], out[96], out[97], out[98], out[99], out[100], out[101], out[102], out[103], out[104], out[105], out[106], out[107], out[108], out[109], out[110], out[111], out[112], out[113], out[114], out[115], out[116], out[117], out[118], out[119], out[120], out[121], out[122], out[123], out[124], out[125], out[126], out[127], out[128], out[129], out[130], out[131], out[132], out[133], out[134], out[135], out[136], out[137], out[138], out[139], out[140], out[141], out[142], out[143], out[144], out[145], out[146], out[147], out[148], out[149], out[150], out[151], out[152], out[153], out[154], out[155], out[156], out[157], out[158], out[159], out[160], out[161], out[162], out[163], out[164], out[165], out[166], out[167], out[168], out[169], out[170], out[171], out[172], out[173], out[174], out[175], out[176], out[177], out[178], out[179], out[180], out[181], out[182], out[183], out[184], out[185], out[186], out[187], out[188], out[189], out[190], out[191], out[192], out[193], out[194], out[195], out[196], out[197], out[198], out[199], out[200], out[201], out[202], out[203], out[204], out[205], out[206], out[207], out[208], out[209], out[210], out[211], out[212], out[213], out[214], out[215], out[216], out[217], out[218], out[219], out[220], out[221], out[222], out[223], out[224], out[225], out[226], out[227], out[228], out[229], out[230], out[231], out[232], out[233], out[234], out[235], out[236], out[237], out[238], out[239], out[240], out[241], out[242], out[243], out[244], out[245], out[246], out[247], out[248], out[249], out[250], out[251], out[252], out[253], out[254], out[255], out[256], out[257], out[258], out[259], out[260], out[261], out[262], out[263], out[264], out[265], out[266], out[267], out[268], out[269], out[270], out[271], out[272], out[273], out[274], out[275], out[276], out[277], out[278], out[279], out[280], out[281], out[282], out[283], out[284], out[285], out[286], out[287], out[288], out[289], out[290], out[291], out[292], out[293], out[294], out[295], out[296], out[297], out[298], out[299], out[300], out[301], out[302], out[303], out[304], out[305], out[306], out[307], out[308], out[309], out[310], out[311], out[312], out[313], out[314], out[315], out[316], out[317], out[318], out[319], out[320], out[321], out[322], out[323], out[324], out[325], out[326], out[327], out[328], out[329], out[330], out[331], out[332], out[333], out[334], out[335], out[336], out[337], out[338], out[339], out[340], out[341], out[342], out[343], out[344], out[345], out[346], out[347], out[348], out[349], out[350], out[351], out[352], out[353], out[354], out[355], out[356], out[357], out[358], out[359], out[360], out[361], out[362], out[363], out[364], out[365], out[366], out[367], out[368], out[369], out[370], out[371], out[372], out[373], out[374], out[375], out[376], out[377], out[378], out[379], out[380], out[381], out[382], out[383], out[384], out[385], out[386], out[387], out[388], out[389], out[390], out[391], out[392], out[393], out[394], out[395], out[396], out[397], out[398], out[399], out[400], out[401], out[402], out[403], out[404], out[405], out[406], out[407], out[408], out[409], out[410], out[411], out[412], out[413], out[414], out[415], out[416], out[417], out[418], out[419], out[420], out[421], out[422], out[423], out[424], out[425], out[426], out[427], out[428], out[429], out[430], out[431], out[432], out[433], out[434], out[435], out[436], out[437], out[438], out[439], out[440], out[441], out[442], out[443], out[444], out[445], out[446], out[447], out[448], out[449], out[450], out[451], out[452], out[453], out[454], out[455], out[456], out[457], out[458], out[459], out[460], out[461], out[462], out[463], out[464], out[465], out[466], out[467], out[468], out[469], out[470], out[471], out[472], out[473], out[474], out[475], out[476], out[477], out[478], out[479], out[480], out[481], out[482], out[483], out[484], out[485], out[486], out[487], out[488], out[489], out[490], out[491], out[492], out[493], out[494], out[495], out[496], out[497], out[498], out[499], out[500], out[501], out[502], out[503], out[504], out[505], out[506], out[507], out[508], out[509], out[510], out[511], out[512], out[513], out[514], out[515], out[516], out[517], out[518], out[519], out[520], out[521], out[522], out[523], out[524], out[525], out[526], out[527], out[528], out[529], out[530], out[531], out[532], out[533], out[534], out[535], out[536], out[537], out[538], out[539], out[540], out[541], out[542], out[543], out[544], out[545], out[546], out[547], out[548], out[549], out[550], out[551], out[552], out[553], out[554], out[555], out[556], out[557], out[558], out[559], out[560], out[561], out[562], out[563], out[564], out[565], out[566], out[567], out[568], out[569], out[570], out[571], out[572], out[573], out[574], out[575], out[576], out[577], out[578], out[579], out[580], out[581], out[582], out[583], out[584], out[585], out[586], out[587], out[588], out[589], out[590], out[591], out[592], out[593], out[594], out[595], out[596], out[597], out[598], out[599], out[600], out[601], out[602], out[603], out[604], out[605], out[606], out[607], out[608], out[609], out[610], out[611], out[612], out[613], out[614], out[615], out[616], out[617], out[618], out[619], out[620], out[621], out[622], out[623], out[624], out[625], out[626], out[627], out[628], out[629], out[630], out[631], out[632], out[633], out[634], out[635], out[636], out[637], out[638], out[639], out[640], out[641], out[642], out[643], out[644], out[645], out[646], out[647];
  not g_43794_(out[320], _39295_);
  not g_43795_(out[321], _39306_);
  not g_43796_(out[322], _39317_);
  not g_43797_(out[323], _39328_);
  not g_43798_(out[324], _39339_);
  not g_43799_(out[325], _39350_);
  not g_43800_(out[326], _39361_);
  not g_43801_(out[327], _39372_);
  not g_43802_(out[7], _39383_);
  not g_43803_(out[328], _39394_);
  not g_43804_(out[329], _39405_);
  not g_43805_(out[330], _39416_);
  not g_43806_(out[331], _39427_);
  not g_43807_(out[11], _39438_);
  not g_43808_(out[332], _39449_);
  not g_43809_(out[333], _39460_);
  not g_43810_(out[334], _39471_);
  not g_43811_(out[335], _39482_);
  not g_43812_(out[27], _39493_);
  not g_43813_(out[28], _39504_);
  not g_43814_(out[39], _39515_);
  not g_43815_(out[43], _39526_);
  not g_43816_(out[59], _39537_);
  not g_43817_(out[75], _39548_);
  not g_43818_(out[91], _39559_);
  not g_43819_(out[107], _39570_);
  not g_43820_(out[123], _39581_);
  not g_43821_(out[139], _39592_);
  not g_43822_(out[155], _39603_);
  not g_43823_(out[171], _39614_);
  not g_43824_(out[187], _39625_);
  not g_43825_(out[203], _39636_);
  not g_43826_(out[219], _39647_);
  not g_43827_(out[235], _39658_);
  not g_43828_(out[251], _39669_);
  not g_43829_(out[267], _39680_);
  not g_43830_(out[283], _39691_);
  not g_43831_(out[299], _39702_);
  not g_43832_(out[311], _39713_);
  not g_43833_(out[315], _39724_);
  not g_43834_(out[347], _39735_);
  not g_43835_(out[363], _39746_);
  not g_43836_(out[379], _39757_);
  not g_43837_(out[395], _39768_);
  not g_43838_(out[411], _39779_);
  not g_43839_(out[427], _39790_);
  not g_43840_(out[443], _39801_);
  not g_43841_(out[459], _39812_);
  not g_43842_(out[475], _39823_);
  not g_43843_(out[491], _39834_);
  not g_43844_(out[507], _39845_);
  not g_43845_(out[523], _39856_);
  not g_43846_(out[539], _39867_);
  not g_43847_(out[555], _39878_);
  not g_43848_(out[571], _39889_);
  not g_43849_(out[587], _39900_);
  not g_43850_(out[603], _39911_);
  not g_43851_(out[619], _39922_);
  not g_43852_(out[631], _39933_);
  not g_43853_(out[635], _39944_);
  and g_43854_(_39713_, out[631], _39955_);
  and g_43855_(out[311], _39933_, _39966_);
  xor g_43856_(out[304], out[624], _39977_);
  xor g_43857_(out[319], out[639], _39988_);
  xor g_43858_(out[315], out[635], _39999_);
  xor g_43859_(out[308], out[628], _40010_);
  xor g_43860_(out[309], out[629], _40021_);
  xor g_43861_(out[314], out[634], _40032_);
  xor g_43862_(out[312], out[632], _40043_);
  xor g_43863_(out[307], out[627], _40054_);
  xor g_43864_(out[305], out[625], _40065_);
  xor g_43865_(out[317], out[637], _40076_);
  xor g_43866_(out[318], out[638], _40087_);
  xor g_43867_(out[310], out[630], _40098_);
  xor g_43868_(out[316], out[636], _40109_);
  or g_43869_(_40010_, _40054_, _40120_);
  xor g_43870_(out[313], out[633], _40131_);
  or g_43871_(_40032_, _40098_, _40142_);
  or g_43872_(_40120_, _40142_, _40153_);
  or g_43873_(_39999_, _40021_, _40164_);
  or g_43874_(_40076_, _40164_, _40175_);
  or g_43875_(_40153_, _40175_, _40186_);
  or g_43876_(_39977_, _40109_, _40197_);
  or g_43877_(_40186_, _40197_, _40208_);
  xor g_43878_(out[306], out[626], _40219_);
  or g_43879_(_39955_, _40219_, _40230_);
  or g_43880_(_39988_, _40087_, _40241_);
  or g_43881_(_40230_, _40241_, _40252_);
  or g_43882_(_39966_, _40131_, _40263_);
  or g_43883_(_40065_, _40263_, _40274_);
  or g_43884_(_40252_, _40274_, _40285_);
  or g_43885_(_40043_, _40285_, _40296_);
  or g_43886_(_40208_, _40296_, _40307_);
  xor g_43887_(out[295], out[631], _40318_);
  and g_43888_(_39702_, out[635], _40329_);
  xor g_43889_(out[302], out[638], _40340_);
  xor g_43890_(out[296], out[632], _40351_);
  xor g_43891_(out[289], out[625], _40362_);
  xor g_43892_(out[301], out[637], _40373_);
  xor g_43893_(out[297], out[633], _40384_);
  xor g_43894_(out[292], out[628], _40395_);
  xor g_43895_(out[290], out[626], _40406_);
  and g_43896_(out[299], _39944_, _40417_);
  xor g_43897_(out[291], out[627], _40428_);
  xor g_43898_(out[294], out[630], _40439_);
  xor g_43899_(out[303], out[639], _40450_);
  xor g_43900_(out[298], out[634], _40461_);
  xor g_43901_(out[293], out[629], _40472_);
  xor g_43902_(out[288], out[624], _40483_);
  or g_43903_(_40340_, _40395_, _40494_);
  or g_43904_(_40351_, _40373_, _40505_);
  or g_43905_(_40406_, _40461_, _40516_);
  or g_43906_(_40505_, _40516_, _40527_);
  or g_43907_(_40384_, _40428_, _40538_);
  or g_43908_(_40472_, _40483_, _40549_);
  or g_43909_(_40538_, _40549_, _40560_);
  or g_43910_(_40527_, _40560_, _40571_);
  xor g_43911_(out[300], out[636], _40582_);
  or g_43912_(_40329_, _40582_, _40593_);
  or g_43913_(_40318_, _40439_, _40604_);
  or g_43914_(_40593_, _40604_, _40615_);
  or g_43915_(_40362_, _40417_, _40626_);
  or g_43916_(_40450_, _40626_, _40637_);
  or g_43917_(_40615_, _40637_, _40648_);
  or g_43918_(_40571_, _40648_, _40659_);
  or g_43919_(_40494_, _40659_, _40670_);
  xor g_43920_(out[273], out[625], _40681_);
  and g_43921_(out[283], _39944_, _40692_);
  xor g_43922_(out[286], out[638], _40703_);
  xor g_43923_(out[275], out[627], _40714_);
  xor g_43924_(out[276], out[628], _40725_);
  xor g_43925_(out[274], out[626], _40736_);
  xor g_43926_(out[281], out[633], _40747_);
  xor g_43927_(out[272], out[624], _40758_);
  and g_43928_(_39691_, out[635], _40769_);
  xor g_43929_(out[278], out[630], _40780_);
  xor g_43930_(out[282], out[634], _40791_);
  xor g_43931_(out[277], out[629], _40802_);
  xor g_43932_(out[287], out[639], _40813_);
  xor g_43933_(out[285], out[637], _40824_);
  xor g_43934_(out[280], out[632], _40835_);
  or g_43935_(_40703_, _40725_, _40846_);
  or g_43936_(_40824_, _40835_, _40857_);
  or g_43937_(_40736_, _40791_, _40868_);
  or g_43938_(_40857_, _40868_, _40879_);
  or g_43939_(_40714_, _40747_, _40890_);
  or g_43940_(_40758_, _40802_, _40901_);
  or g_43941_(_40890_, _40901_, _40912_);
  or g_43942_(_40879_, _40912_, _40923_);
  xor g_43943_(out[284], out[636], _40934_);
  or g_43944_(_40769_, _40934_, _40945_);
  xor g_43945_(out[279], out[631], _40956_);
  or g_43946_(_40780_, _40956_, _40967_);
  or g_43947_(_40945_, _40967_, _40978_);
  or g_43948_(_40681_, _40692_, _40989_);
  or g_43949_(_40813_, _40989_, _41000_);
  or g_43950_(_40978_, _41000_, _41011_);
  or g_43951_(_40923_, _41011_, _41022_);
  or g_43952_(_40846_, _41022_, _41033_);
  xor g_43953_(out[263], out[631], _41044_);
  and g_43954_(_39680_, out[635], _41055_);
  xor g_43955_(out[270], out[638], _41066_);
  xor g_43956_(out[264], out[632], _41077_);
  xor g_43957_(out[257], out[625], _41088_);
  xor g_43958_(out[269], out[637], _41099_);
  xor g_43959_(out[265], out[633], _41110_);
  xor g_43960_(out[260], out[628], _41121_);
  xor g_43961_(out[258], out[626], _41132_);
  and g_43962_(out[267], _39944_, _41143_);
  xor g_43963_(out[259], out[627], _41154_);
  xor g_43964_(out[262], out[630], _41165_);
  xor g_43965_(out[271], out[639], _41176_);
  xor g_43966_(out[266], out[634], _41187_);
  xor g_43967_(out[261], out[629], _41198_);
  xor g_43968_(out[256], out[624], _41209_);
  or g_43969_(_41066_, _41121_, _41220_);
  or g_43970_(_41077_, _41099_, _41231_);
  or g_43971_(_41132_, _41187_, _41242_);
  or g_43972_(_41231_, _41242_, _41253_);
  or g_43973_(_41110_, _41154_, _41264_);
  or g_43974_(_41198_, _41209_, _41275_);
  or g_43975_(_41264_, _41275_, _41286_);
  or g_43976_(_41253_, _41286_, _41297_);
  xor g_43977_(out[268], out[636], _41308_);
  or g_43978_(_41055_, _41308_, _41319_);
  or g_43979_(_41044_, _41165_, _41330_);
  or g_43980_(_41319_, _41330_, _41341_);
  or g_43981_(_41088_, _41143_, _41352_);
  or g_43982_(_41176_, _41352_, _41363_);
  or g_43983_(_41341_, _41363_, _41374_);
  or g_43984_(_41297_, _41374_, _41385_);
  or g_43985_(_41220_, _41385_, _41396_);
  xor g_43986_(out[241], out[625], _41407_);
  and g_43987_(out[251], _39944_, _41418_);
  xor g_43988_(out[249], out[633], _41429_);
  xor g_43989_(out[240], out[624], _41440_);
  xor g_43990_(out[254], out[638], _41451_);
  xor g_43991_(out[244], out[628], _41462_);
  or g_43992_(_41451_, _41462_, _41473_);
  xor g_43993_(out[253], out[637], _41484_);
  xor g_43994_(out[243], out[627], _41495_);
  and g_43995_(_39669_, out[635], _41506_);
  xor g_43996_(out[246], out[630], _41517_);
  xor g_43997_(out[250], out[634], _41528_);
  xor g_43998_(out[245], out[629], _41539_);
  xor g_43999_(out[255], out[639], _41550_);
  xor g_44000_(out[248], out[632], _41561_);
  or g_44001_(_41484_, _41561_, _41572_);
  xor g_44002_(out[242], out[626], _41583_);
  or g_44003_(_41528_, _41583_, _41594_);
  or g_44004_(_41572_, _41594_, _41605_);
  or g_44005_(_41429_, _41495_, _41616_);
  or g_44006_(_41539_, _41616_, _41627_);
  or g_44007_(_41605_, _41627_, _41638_);
  or g_44008_(_41473_, _41638_, _41649_);
  xor g_44009_(out[252], out[636], _41660_);
  or g_44010_(_41506_, _41660_, _41671_);
  xor g_44011_(out[247], out[631], _41682_);
  or g_44012_(_41517_, _41682_, _41693_);
  or g_44013_(_41671_, _41693_, _41704_);
  or g_44014_(_41407_, _41418_, _41715_);
  or g_44015_(_41550_, _41715_, _41726_);
  or g_44016_(_41704_, _41726_, _41737_);
  or g_44017_(_41440_, _41737_, _41748_);
  or g_44018_(_41649_, _41748_, _41759_);
  xor g_44019_(out[231], out[631], _41770_);
  and g_44020_(_39658_, out[635], _41781_);
  xor g_44021_(out[238], out[638], _41792_);
  xor g_44022_(out[232], out[632], _41803_);
  xor g_44023_(out[225], out[625], _41814_);
  xor g_44024_(out[237], out[637], _41825_);
  xor g_44025_(out[233], out[633], _41836_);
  xor g_44026_(out[228], out[628], _41847_);
  xor g_44027_(out[226], out[626], _41858_);
  and g_44028_(out[235], _39944_, _41869_);
  xor g_44029_(out[227], out[627], _41880_);
  xor g_44030_(out[230], out[630], _41891_);
  xor g_44031_(out[239], out[639], _41902_);
  xor g_44032_(out[234], out[634], _41913_);
  xor g_44033_(out[229], out[629], _41924_);
  xor g_44034_(out[224], out[624], _41935_);
  or g_44035_(_41792_, _41847_, _41946_);
  or g_44036_(_41803_, _41825_, _41957_);
  or g_44037_(_41858_, _41913_, _41968_);
  or g_44038_(_41957_, _41968_, _41979_);
  or g_44039_(_41836_, _41880_, _41990_);
  or g_44040_(_41924_, _41935_, _42001_);
  or g_44041_(_41990_, _42001_, _42012_);
  or g_44042_(_41979_, _42012_, _42023_);
  xor g_44043_(out[236], out[636], _42034_);
  or g_44044_(_41781_, _42034_, _42045_);
  or g_44045_(_41770_, _41891_, _42056_);
  or g_44046_(_42045_, _42056_, _42067_);
  or g_44047_(_41814_, _41869_, _42078_);
  or g_44048_(_41902_, _42078_, _42089_);
  or g_44049_(_42067_, _42089_, _42100_);
  or g_44050_(_42023_, _42100_, _42111_);
  or g_44051_(_41946_, _42111_, _42122_);
  xor g_44052_(out[209], out[625], _42133_);
  and g_44053_(out[219], _39944_, _42144_);
  xor g_44054_(out[217], out[633], _42155_);
  xor g_44055_(out[208], out[624], _42166_);
  xor g_44056_(out[222], out[638], _42177_);
  xor g_44057_(out[212], out[628], _42188_);
  or g_44058_(_42177_, _42188_, _42199_);
  xor g_44059_(out[221], out[637], _42210_);
  xor g_44060_(out[211], out[627], _42221_);
  and g_44061_(_39647_, out[635], _42232_);
  xor g_44062_(out[214], out[630], _42243_);
  xor g_44063_(out[218], out[634], _42254_);
  xor g_44064_(out[213], out[629], _42265_);
  xor g_44065_(out[223], out[639], _42276_);
  xor g_44066_(out[216], out[632], _42287_);
  or g_44067_(_42210_, _42287_, _42298_);
  xor g_44068_(out[210], out[626], _42309_);
  or g_44069_(_42254_, _42309_, _42320_);
  or g_44070_(_42298_, _42320_, _42331_);
  or g_44071_(_42155_, _42221_, _42342_);
  or g_44072_(_42265_, _42342_, _42353_);
  or g_44073_(_42331_, _42353_, _42364_);
  or g_44074_(_42199_, _42364_, _42375_);
  xor g_44075_(out[220], out[636], _42386_);
  or g_44076_(_42232_, _42386_, _42397_);
  xor g_44077_(out[215], out[631], _42408_);
  or g_44078_(_42243_, _42408_, _42419_);
  or g_44079_(_42397_, _42419_, _42430_);
  or g_44080_(_42133_, _42144_, _42441_);
  or g_44081_(_42276_, _42441_, _42452_);
  or g_44082_(_42430_, _42452_, _42463_);
  or g_44083_(_42166_, _42463_, _42474_);
  or g_44084_(_42375_, _42474_, _42485_);
  xor g_44085_(out[199], out[631], _42496_);
  and g_44086_(_39636_, out[635], _42507_);
  xor g_44087_(out[206], out[638], _42518_);
  xor g_44088_(out[200], out[632], _42529_);
  xor g_44089_(out[193], out[625], _42540_);
  xor g_44090_(out[205], out[637], _42551_);
  xor g_44091_(out[201], out[633], _42562_);
  xor g_44092_(out[196], out[628], _42573_);
  xor g_44093_(out[194], out[626], _42584_);
  and g_44094_(out[203], _39944_, _42595_);
  xor g_44095_(out[195], out[627], _42606_);
  xor g_44096_(out[198], out[630], _42617_);
  xor g_44097_(out[207], out[639], _42628_);
  xor g_44098_(out[202], out[634], _42639_);
  xor g_44099_(out[197], out[629], _42650_);
  xor g_44100_(out[192], out[624], _42661_);
  or g_44101_(_42518_, _42573_, _42672_);
  or g_44102_(_42529_, _42551_, _42683_);
  or g_44103_(_42584_, _42639_, _42694_);
  or g_44104_(_42683_, _42694_, _42705_);
  or g_44105_(_42562_, _42606_, _42716_);
  or g_44106_(_42650_, _42661_, _42727_);
  or g_44107_(_42716_, _42727_, _42738_);
  or g_44108_(_42705_, _42738_, _42749_);
  xor g_44109_(out[204], out[636], _42760_);
  or g_44110_(_42507_, _42760_, _42771_);
  or g_44111_(_42496_, _42617_, _42782_);
  or g_44112_(_42771_, _42782_, _42793_);
  or g_44113_(_42540_, _42595_, _42804_);
  or g_44114_(_42628_, _42804_, _42815_);
  or g_44115_(_42793_, _42815_, _42826_);
  or g_44116_(_42749_, _42826_, _42837_);
  or g_44117_(_42672_, _42837_, _42848_);
  xor g_44118_(out[189], out[637], _42859_);
  xor g_44119_(out[178], out[626], _42870_);
  xor g_44120_(out[181], out[629], _42881_);
  xor g_44121_(out[185], out[633], _42892_);
  xor g_44122_(out[180], out[628], _42903_);
  xor g_44123_(out[184], out[632], _42914_);
  xor g_44124_(out[190], out[638], _42925_);
  xor g_44125_(out[182], out[630], _42936_);
  xor g_44126_(out[191], out[639], _42947_);
  xor g_44127_(out[186], out[634], _42958_);
  xor g_44128_(out[176], out[624], _42969_);
  xor g_44129_(out[179], out[627], _42980_);
  and g_44130_(_39625_, out[635], _42991_);
  and g_44131_(out[187], _39944_, _43002_);
  xor g_44132_(out[177], out[625], _43013_);
  or g_44133_(_42903_, _42925_, _43024_);
  or g_44134_(_42859_, _42914_, _43035_);
  or g_44135_(_42870_, _42958_, _43046_);
  or g_44136_(_43035_, _43046_, _43057_);
  or g_44137_(_42892_, _42980_, _43068_);
  or g_44138_(_42881_, _42969_, _43079_);
  or g_44139_(_43068_, _43079_, _43090_);
  or g_44140_(_43057_, _43090_, _43101_);
  xor g_44141_(out[188], out[636], _43112_);
  or g_44142_(_42991_, _43112_, _43123_);
  xor g_44143_(out[183], out[631], _43134_);
  or g_44144_(_42936_, _43134_, _43145_);
  or g_44145_(_43123_, _43145_, _21900_);
  or g_44146_(_43002_, _43013_, _21911_);
  or g_44147_(_42947_, _21911_, _21922_);
  or g_44148_(_21900_, _21922_, _21933_);
  or g_44149_(_43101_, _21933_, _21944_);
  or g_44150_(_43024_, _21944_, _21955_);
  xor g_44151_(out[167], out[631], _21966_);
  and g_44152_(_39614_, out[635], _21977_);
  xor g_44153_(out[174], out[638], _21988_);
  xor g_44154_(out[168], out[632], _21999_);
  xor g_44155_(out[161], out[625], _22010_);
  xor g_44156_(out[173], out[637], _22021_);
  xor g_44157_(out[169], out[633], _22032_);
  xor g_44158_(out[164], out[628], _22043_);
  xor g_44159_(out[162], out[626], _22054_);
  and g_44160_(out[171], _39944_, _22065_);
  xor g_44161_(out[163], out[627], _22076_);
  xor g_44162_(out[166], out[630], _22087_);
  xor g_44163_(out[175], out[639], _22098_);
  xor g_44164_(out[170], out[634], _22109_);
  xor g_44165_(out[165], out[629], _22120_);
  xor g_44166_(out[160], out[624], _22131_);
  or g_44167_(_21988_, _22043_, _22142_);
  or g_44168_(_21999_, _22021_, _22153_);
  or g_44169_(_22054_, _22109_, _22164_);
  or g_44170_(_22153_, _22164_, _22175_);
  or g_44171_(_22032_, _22076_, _22186_);
  or g_44172_(_22120_, _22131_, _22197_);
  or g_44173_(_22186_, _22197_, _22208_);
  or g_44174_(_22175_, _22208_, _22219_);
  xor g_44175_(out[172], out[636], _22230_);
  or g_44176_(_21977_, _22230_, _22241_);
  or g_44177_(_21966_, _22087_, _22252_);
  or g_44178_(_22241_, _22252_, _22263_);
  or g_44179_(_22010_, _22065_, _22274_);
  or g_44180_(_22098_, _22274_, _22285_);
  or g_44181_(_22263_, _22285_, _22296_);
  or g_44182_(_22219_, _22296_, _22307_);
  or g_44183_(_22142_, _22307_, _22318_);
  xor g_44184_(out[156], out[636], _22329_);
  and g_44185_(_39603_, out[635], _22340_);
  xor g_44186_(out[152], out[632], _22351_);
  xor g_44187_(out[150], out[630], _22362_);
  xor g_44188_(out[157], out[637], _22373_);
  xor g_44189_(out[158], out[638], _22384_);
  xor g_44190_(out[146], out[626], _22395_);
  xor g_44191_(out[153], out[633], _22406_);
  xor g_44192_(out[149], out[629], _22417_);
  xor g_44193_(out[145], out[625], _22428_);
  and g_44194_(out[155], _39944_, _22439_);
  or g_44195_(_22351_, _22373_, _22450_);
  xor g_44196_(out[159], out[639], _22461_);
  xor g_44197_(out[154], out[634], _22472_);
  xor g_44198_(out[148], out[628], _22483_);
  xor g_44199_(out[147], out[627], _22494_);
  xor g_44200_(out[144], out[624], _22505_);
  or g_44201_(_22395_, _22472_, _22516_);
  or g_44202_(_22450_, _22516_, _22527_);
  or g_44203_(_22406_, _22494_, _22538_);
  or g_44204_(_22417_, _22538_, _22549_);
  or g_44205_(_22527_, _22549_, _22560_);
  or g_44206_(_22384_, _22483_, _22571_);
  or g_44207_(_22560_, _22571_, _22582_);
  or g_44208_(_22329_, _22340_, _22593_);
  xor g_44209_(out[151], out[631], _22604_);
  or g_44210_(_22362_, _22604_, _22615_);
  or g_44211_(_22593_, _22615_, _22626_);
  or g_44212_(_22428_, _22439_, _22637_);
  or g_44213_(_22461_, _22637_, _22648_);
  or g_44214_(_22626_, _22648_, _22659_);
  or g_44215_(_22505_, _22659_, _22670_);
  or g_44216_(_22582_, _22670_, _22681_);
  xor g_44217_(out[135], out[631], _22692_);
  and g_44218_(_39592_, out[635], _22703_);
  xor g_44219_(out[142], out[638], _22714_);
  xor g_44220_(out[136], out[632], _22725_);
  xor g_44221_(out[129], out[625], _22736_);
  xor g_44222_(out[141], out[637], _22747_);
  xor g_44223_(out[137], out[633], _22758_);
  xor g_44224_(out[132], out[628], _22769_);
  xor g_44225_(out[130], out[626], _22780_);
  and g_44226_(out[139], _39944_, _22791_);
  xor g_44227_(out[131], out[627], _22802_);
  xor g_44228_(out[134], out[630], _22813_);
  xor g_44229_(out[143], out[639], _22824_);
  xor g_44230_(out[138], out[634], _22835_);
  xor g_44231_(out[133], out[629], _22846_);
  xor g_44232_(out[128], out[624], _22857_);
  or g_44233_(_22714_, _22769_, _22868_);
  or g_44234_(_22725_, _22747_, _22879_);
  or g_44235_(_22780_, _22835_, _22890_);
  or g_44236_(_22879_, _22890_, _22901_);
  or g_44237_(_22758_, _22802_, _22912_);
  or g_44238_(_22846_, _22857_, _22923_);
  or g_44239_(_22912_, _22923_, _22934_);
  or g_44240_(_22901_, _22934_, _22945_);
  xor g_44241_(out[140], out[636], _22956_);
  or g_44242_(_22703_, _22956_, _22967_);
  or g_44243_(_22692_, _22813_, _22978_);
  or g_44244_(_22967_, _22978_, _22989_);
  or g_44245_(_22736_, _22791_, _23000_);
  or g_44246_(_22824_, _23000_, _23011_);
  or g_44247_(_22989_, _23011_, _23022_);
  or g_44248_(_22945_, _23022_, _23033_);
  or g_44249_(_22868_, _23033_, _23044_);
  xor g_44250_(out[115], out[627], _23055_);
  xor g_44251_(out[116], out[628], _23066_);
  xor g_44252_(out[126], out[638], _23077_);
  xor g_44253_(out[114], out[626], _23088_);
  xor g_44254_(out[117], out[629], _23099_);
  xor g_44255_(out[121], out[633], _23110_);
  xor g_44256_(out[120], out[632], _23121_);
  xor g_44257_(out[127], out[639], _23132_);
  xor g_44258_(out[122], out[634], _23143_);
  xor g_44259_(out[118], out[630], _23154_);
  xor g_44260_(out[112], out[624], _23165_);
  and g_44261_(_39581_, out[635], _23176_);
  and g_44262_(out[123], _39944_, _23187_);
  xor g_44263_(out[125], out[637], _23198_);
  or g_44264_(_23121_, _23198_, _23209_);
  xor g_44265_(out[113], out[625], _23220_);
  or g_44266_(_23088_, _23143_, _23231_);
  or g_44267_(_23209_, _23231_, _23242_);
  or g_44268_(_23055_, _23110_, _23253_);
  or g_44269_(_23099_, _23253_, _23264_);
  or g_44270_(_23242_, _23264_, _23275_);
  or g_44271_(_23066_, _23077_, _23286_);
  or g_44272_(_23275_, _23286_, _23297_);
  xor g_44273_(out[124], out[636], _23308_);
  or g_44274_(_23176_, _23308_, _23319_);
  xor g_44275_(out[119], out[631], _23330_);
  or g_44276_(_23154_, _23330_, _23341_);
  or g_44277_(_23319_, _23341_, _23352_);
  or g_44278_(_23187_, _23220_, _23363_);
  or g_44279_(_23132_, _23363_, _23374_);
  or g_44280_(_23352_, _23374_, _23385_);
  or g_44281_(_23165_, _23385_, _23396_);
  or g_44282_(_23297_, _23396_, _23407_);
  xor g_44283_(out[103], out[631], _23418_);
  and g_44284_(_39570_, out[635], _23429_);
  xor g_44285_(out[110], out[638], _23440_);
  xor g_44286_(out[104], out[632], _23451_);
  xor g_44287_(out[97], out[625], _23462_);
  xor g_44288_(out[109], out[637], _23473_);
  xor g_44289_(out[105], out[633], _23484_);
  xor g_44290_(out[100], out[628], _23495_);
  xor g_44291_(out[98], out[626], _23506_);
  and g_44292_(out[107], _39944_, _23517_);
  xor g_44293_(out[99], out[627], _23528_);
  xor g_44294_(out[102], out[630], _23539_);
  xor g_44295_(out[111], out[639], _23550_);
  xor g_44296_(out[106], out[634], _23561_);
  xor g_44297_(out[101], out[629], _23572_);
  xor g_44298_(out[96], out[624], _23583_);
  or g_44299_(_23440_, _23495_, _23594_);
  or g_44300_(_23451_, _23473_, _23605_);
  or g_44301_(_23506_, _23561_, _23616_);
  or g_44302_(_23605_, _23616_, _23627_);
  or g_44303_(_23484_, _23528_, _23638_);
  or g_44304_(_23572_, _23583_, _23649_);
  or g_44305_(_23638_, _23649_, _23660_);
  or g_44306_(_23627_, _23660_, _23671_);
  xor g_44307_(out[108], out[636], _23682_);
  or g_44308_(_23429_, _23682_, _23693_);
  or g_44309_(_23418_, _23539_, _23704_);
  or g_44310_(_23693_, _23704_, _23715_);
  or g_44311_(_23462_, _23517_, _23726_);
  or g_44312_(_23550_, _23726_, _23737_);
  or g_44313_(_23715_, _23737_, _23748_);
  or g_44314_(_23671_, _23748_, _23759_);
  or g_44315_(_23594_, _23759_, _23770_);
  xor g_44316_(out[92], out[636], _23781_);
  and g_44317_(_39559_, out[635], _23792_);
  xor g_44318_(out[93], out[637], _23803_);
  xor g_44319_(out[86], out[630], _23814_);
  xor g_44320_(out[88], out[632], _23825_);
  xor g_44321_(out[89], out[633], _23836_);
  xor g_44322_(out[94], out[638], _23847_);
  xor g_44323_(out[84], out[628], _23858_);
  or g_44324_(_23847_, _23858_, _23869_);
  xor g_44325_(out[85], out[629], _23880_);
  xor g_44326_(out[81], out[625], _23891_);
  and g_44327_(out[91], _39944_, _23902_);
  xor g_44328_(out[95], out[639], _23913_);
  xor g_44329_(out[90], out[634], _23924_);
  xor g_44330_(out[80], out[624], _23935_);
  xor g_44331_(out[82], out[626], _23946_);
  xor g_44332_(out[83], out[627], _23957_);
  or g_44333_(_23803_, _23825_, _23968_);
  or g_44334_(_23924_, _23946_, _23979_);
  or g_44335_(_23968_, _23979_, _23990_);
  or g_44336_(_23836_, _23957_, _24001_);
  or g_44337_(_23880_, _23935_, _24012_);
  or g_44338_(_24001_, _24012_, _24023_);
  or g_44339_(_23990_, _24023_, _24034_);
  or g_44340_(_23781_, _23792_, _24045_);
  xor g_44341_(out[87], out[631], _24056_);
  or g_44342_(_23814_, _24056_, _24067_);
  or g_44343_(_24045_, _24067_, _24078_);
  or g_44344_(_23891_, _23902_, _24089_);
  or g_44345_(_23913_, _24089_, _24100_);
  or g_44346_(_24078_, _24100_, _24111_);
  or g_44347_(_24034_, _24111_, _24122_);
  or g_44348_(_23869_, _24122_, _24133_);
  xor g_44349_(out[71], out[631], _24144_);
  and g_44350_(_39548_, out[635], _24155_);
  xor g_44351_(out[78], out[638], _24166_);
  xor g_44352_(out[72], out[632], _24177_);
  xor g_44353_(out[65], out[625], _24188_);
  xor g_44354_(out[77], out[637], _24199_);
  xor g_44355_(out[73], out[633], _24210_);
  xor g_44356_(out[68], out[628], _24221_);
  xor g_44357_(out[66], out[626], _24232_);
  and g_44358_(out[75], _39944_, _24243_);
  xor g_44359_(out[67], out[627], _24254_);
  xor g_44360_(out[70], out[630], _24265_);
  xor g_44361_(out[79], out[639], _24276_);
  xor g_44362_(out[74], out[634], _24287_);
  xor g_44363_(out[69], out[629], _24298_);
  xor g_44364_(out[64], out[624], _24309_);
  or g_44365_(_24166_, _24221_, _24320_);
  or g_44366_(_24177_, _24199_, _24331_);
  or g_44367_(_24232_, _24287_, _24342_);
  or g_44368_(_24331_, _24342_, _24353_);
  or g_44369_(_24210_, _24254_, _24364_);
  or g_44370_(_24298_, _24309_, _24375_);
  or g_44371_(_24364_, _24375_, _24386_);
  or g_44372_(_24353_, _24386_, _24397_);
  xor g_44373_(out[76], out[636], _24408_);
  or g_44374_(_24155_, _24408_, _24419_);
  or g_44375_(_24144_, _24265_, _24430_);
  or g_44376_(_24419_, _24430_, _24441_);
  or g_44377_(_24188_, _24243_, _24452_);
  or g_44378_(_24276_, _24452_, _24463_);
  or g_44379_(_24441_, _24463_, _24474_);
  or g_44380_(_24397_, _24474_, _24485_);
  or g_44381_(_24320_, _24485_, _24496_);
  xor g_44382_(out[49], out[625], _24507_);
  and g_44383_(out[59], _39944_, _24518_);
  xor g_44384_(out[57], out[633], _24529_);
  xor g_44385_(out[48], out[624], _24540_);
  xor g_44386_(out[62], out[638], _24551_);
  xor g_44387_(out[52], out[628], _24562_);
  or g_44388_(_24551_, _24562_, _24573_);
  xor g_44389_(out[61], out[637], _24584_);
  xor g_44390_(out[51], out[627], _24595_);
  and g_44391_(_39537_, out[635], _24606_);
  xor g_44392_(out[54], out[630], _24617_);
  xor g_44393_(out[58], out[634], _24628_);
  xor g_44394_(out[53], out[629], _24639_);
  xor g_44395_(out[63], out[639], _24650_);
  xor g_44396_(out[56], out[632], _24661_);
  or g_44397_(_24584_, _24661_, _24672_);
  xor g_44398_(out[50], out[626], _24683_);
  or g_44399_(_24628_, _24683_, _24694_);
  or g_44400_(_24672_, _24694_, _24705_);
  or g_44401_(_24529_, _24595_, _24716_);
  or g_44402_(_24639_, _24716_, _24727_);
  or g_44403_(_24705_, _24727_, _24738_);
  or g_44404_(_24573_, _24738_, _24749_);
  xor g_44405_(out[60], out[636], _24760_);
  or g_44406_(_24606_, _24760_, _24771_);
  xor g_44407_(out[55], out[631], _24782_);
  or g_44408_(_24617_, _24782_, _24793_);
  or g_44409_(_24771_, _24793_, _24804_);
  or g_44410_(_24507_, _24518_, _24815_);
  or g_44411_(_24650_, _24815_, _24826_);
  or g_44412_(_24804_, _24826_, _24837_);
  or g_44413_(_24540_, _24837_, _24848_);
  or g_44414_(_24749_, _24848_, _24859_);
  xor g_44415_(out[39], out[631], _24870_);
  and g_44416_(_39526_, out[635], _24881_);
  xor g_44417_(out[46], out[638], _24892_);
  xor g_44418_(out[40], out[632], _24903_);
  xor g_44419_(out[33], out[625], _24914_);
  xor g_44420_(out[45], out[637], _24925_);
  xor g_44421_(out[41], out[633], _24936_);
  xor g_44422_(out[36], out[628], _24947_);
  xor g_44423_(out[34], out[626], _24958_);
  and g_44424_(out[43], _39944_, _24969_);
  xor g_44425_(out[35], out[627], _24980_);
  xor g_44426_(out[38], out[630], _24991_);
  xor g_44427_(out[47], out[639], _25002_);
  xor g_44428_(out[42], out[634], _25013_);
  xor g_44429_(out[37], out[629], _25024_);
  xor g_44430_(out[32], out[624], _25035_);
  or g_44431_(_24892_, _24947_, _25046_);
  or g_44432_(_24903_, _24925_, _25057_);
  or g_44433_(_24958_, _25013_, _25068_);
  or g_44434_(_25057_, _25068_, _25079_);
  or g_44435_(_24936_, _24980_, _25090_);
  or g_44436_(_25024_, _25035_, _25101_);
  or g_44437_(_25090_, _25101_, _25112_);
  or g_44438_(_25079_, _25112_, _25123_);
  xor g_44439_(out[44], out[636], _25134_);
  or g_44440_(_24881_, _25134_, _25145_);
  or g_44441_(_24870_, _24991_, _25156_);
  or g_44442_(_25145_, _25156_, _25167_);
  or g_44443_(_24914_, _24969_, _25178_);
  or g_44444_(_25002_, _25178_, _25189_);
  or g_44445_(_25167_, _25189_, _25200_);
  or g_44446_(_25123_, _25200_, _25211_);
  or g_44447_(_25046_, _25211_, _25222_);
  xor g_44448_(out[29], out[637], _25233_);
  xor g_44449_(out[18], out[626], _25244_);
  xor g_44450_(out[21], out[629], _25255_);
  xor g_44451_(out[25], out[633], _25266_);
  xor g_44452_(out[20], out[628], _25277_);
  xor g_44453_(out[24], out[632], _25288_);
  xor g_44454_(out[30], out[638], _25299_);
  xor g_44455_(out[22], out[630], _25310_);
  xor g_44456_(out[31], out[639], _25321_);
  xor g_44457_(out[26], out[634], _25332_);
  xor g_44458_(out[16], out[624], _25343_);
  xor g_44459_(out[19], out[627], _25354_);
  and g_44460_(_39493_, out[635], _25365_);
  and g_44461_(out[27], _39944_, _25376_);
  xor g_44462_(out[17], out[625], _25387_);
  or g_44463_(_25277_, _25299_, _25398_);
  or g_44464_(_25233_, _25288_, _25409_);
  or g_44465_(_25244_, _25332_, _25420_);
  or g_44466_(_25409_, _25420_, _25431_);
  or g_44467_(_25266_, _25354_, _25442_);
  or g_44468_(_25255_, _25343_, _25453_);
  or g_44469_(_25442_, _25453_, _25464_);
  or g_44470_(_25431_, _25464_, _25475_);
  xor g_44471_(out[28], out[636], _25486_);
  or g_44472_(_25365_, _25486_, _25497_);
  xor g_44473_(out[23], out[631], _25508_);
  or g_44474_(_25310_, _25508_, _25519_);
  or g_44475_(_25497_, _25519_, _25530_);
  or g_44476_(_25376_, _25387_, _25541_);
  or g_44477_(_25321_, _25541_, _25552_);
  or g_44478_(_25530_, _25552_, _25563_);
  or g_44479_(_25475_, _25563_, _25574_);
  or g_44480_(_25398_, _25574_, _25585_);
  xor g_44481_(out[1], out[625], _25596_);
  and g_44482_(out[11], _39944_, _25607_);
  xor g_44483_(out[9], out[633], _25618_);
  xor g_44484_(out[0], out[624], _25629_);
  xor g_44485_(out[14], out[638], _25640_);
  xor g_44486_(out[4], out[628], _25651_);
  or g_44487_(_25640_, _25651_, _25662_);
  xor g_44488_(out[13], out[637], _25673_);
  xor g_44489_(out[3], out[627], _25684_);
  and g_44490_(_39438_, out[635], _25695_);
  xor g_44491_(out[6], out[630], _25706_);
  xor g_44492_(out[10], out[634], _25717_);
  xor g_44493_(out[5], out[629], _25728_);
  xor g_44494_(out[15], out[639], _25739_);
  xor g_44495_(out[8], out[632], _25750_);
  or g_44496_(_25673_, _25750_, _25761_);
  xor g_44497_(out[2], out[626], _25772_);
  or g_44498_(_25717_, _25772_, _25783_);
  or g_44499_(_25761_, _25783_, _25794_);
  or g_44500_(_25618_, _25684_, _25805_);
  or g_44501_(_25728_, _25805_, _25816_);
  or g_44502_(_25794_, _25816_, _25827_);
  or g_44503_(_25662_, _25827_, _25838_);
  xor g_44504_(out[12], out[636], _25849_);
  or g_44505_(_25695_, _25849_, _25860_);
  xor g_44506_(out[7], out[631], _25871_);
  or g_44507_(_25706_, _25871_, _25882_);
  or g_44508_(_25860_, _25882_, _25893_);
  or g_44509_(_25596_, _25607_, _25904_);
  or g_44510_(_25739_, _25904_, _25915_);
  or g_44511_(_25893_, _25915_, _25926_);
  or g_44512_(_25629_, _25926_, _25937_);
  or g_44513_(_25838_, _25937_, _25948_);
  xor g_44514_(out[311], out[615], _25959_);
  and g_44515_(_39724_, out[619], _25970_);
  xor g_44516_(out[318], out[622], _25981_);
  xor g_44517_(out[312], out[616], _25992_);
  xor g_44518_(out[305], out[609], _26003_);
  xor g_44519_(out[317], out[621], _26014_);
  xor g_44520_(out[313], out[617], _26025_);
  xor g_44521_(out[308], out[612], _26036_);
  xor g_44522_(out[306], out[610], _26047_);
  and g_44523_(out[315], _39922_, _26058_);
  xor g_44524_(out[307], out[611], _26069_);
  xor g_44525_(out[310], out[614], _26080_);
  xor g_44526_(out[319], out[623], _26091_);
  xor g_44527_(out[314], out[618], _26102_);
  xor g_44528_(out[309], out[613], _26113_);
  xor g_44529_(out[304], out[608], _26124_);
  or g_44530_(_25981_, _26036_, _26135_);
  or g_44531_(_25992_, _26014_, _26146_);
  or g_44532_(_26047_, _26102_, _26157_);
  or g_44533_(_26146_, _26157_, _26168_);
  or g_44534_(_26025_, _26069_, _26179_);
  or g_44535_(_26113_, _26124_, _26190_);
  or g_44536_(_26179_, _26190_, _26201_);
  or g_44537_(_26168_, _26201_, _26212_);
  xor g_44538_(out[316], out[620], _26223_);
  or g_44539_(_25970_, _26223_, _26234_);
  or g_44540_(_25959_, _26080_, _26245_);
  or g_44541_(_26234_, _26245_, _26256_);
  or g_44542_(_26003_, _26058_, _26267_);
  or g_44543_(_26091_, _26267_, _26278_);
  or g_44544_(_26256_, _26278_, _26289_);
  or g_44545_(_26212_, _26289_, _26300_);
  or g_44546_(_26135_, _26300_, _26311_);
  not g_44547_(_26311_, _26322_);
  xor g_44548_(out[289], out[609], _26333_);
  and g_44549_(out[299], _39922_, _26344_);
  xor g_44550_(out[297], out[617], _26355_);
  xor g_44551_(out[288], out[608], _26366_);
  xor g_44552_(out[302], out[622], _26377_);
  xor g_44553_(out[292], out[612], _26388_);
  or g_44554_(_26377_, _26388_, _26399_);
  xor g_44555_(out[301], out[621], _26410_);
  xor g_44556_(out[291], out[611], _26421_);
  and g_44557_(_39702_, out[619], _26432_);
  xor g_44558_(out[294], out[614], _26443_);
  xor g_44559_(out[298], out[618], _26454_);
  xor g_44560_(out[293], out[613], _26465_);
  xor g_44561_(out[303], out[623], _26476_);
  xor g_44562_(out[296], out[616], _26487_);
  or g_44563_(_26410_, _26487_, _26498_);
  xor g_44564_(out[290], out[610], _26509_);
  or g_44565_(_26454_, _26509_, _26520_);
  or g_44566_(_26498_, _26520_, _26531_);
  or g_44567_(_26355_, _26421_, _26542_);
  or g_44568_(_26465_, _26542_, _26553_);
  or g_44569_(_26531_, _26553_, _26564_);
  or g_44570_(_26399_, _26564_, _26575_);
  xor g_44571_(out[300], out[620], _26586_);
  or g_44572_(_26432_, _26586_, _26597_);
  xor g_44573_(out[295], out[615], _26608_);
  or g_44574_(_26443_, _26608_, _26619_);
  or g_44575_(_26597_, _26619_, _26630_);
  or g_44576_(_26333_, _26344_, _26641_);
  or g_44577_(_26476_, _26641_, _26652_);
  or g_44578_(_26630_, _26652_, _26663_);
  or g_44579_(_26366_, _26663_, _26674_);
  or g_44580_(_26575_, _26674_, _26685_);
  xor g_44581_(out[279], out[615], _26696_);
  and g_44582_(_39691_, out[619], _26707_);
  xor g_44583_(out[286], out[622], _26718_);
  xor g_44584_(out[280], out[616], _26729_);
  xor g_44585_(out[273], out[609], _26740_);
  xor g_44586_(out[285], out[621], _26751_);
  xor g_44587_(out[281], out[617], _26762_);
  xor g_44588_(out[276], out[612], _26773_);
  xor g_44589_(out[274], out[610], _26784_);
  and g_44590_(out[283], _39922_, _26795_);
  xor g_44591_(out[275], out[611], _26806_);
  xor g_44592_(out[278], out[614], _26817_);
  xor g_44593_(out[287], out[623], _26828_);
  xor g_44594_(out[282], out[618], _26839_);
  xor g_44595_(out[277], out[613], _26850_);
  xor g_44596_(out[272], out[608], _26861_);
  or g_44597_(_26718_, _26773_, _26872_);
  or g_44598_(_26729_, _26751_, _26883_);
  or g_44599_(_26784_, _26839_, _26894_);
  or g_44600_(_26883_, _26894_, _26905_);
  or g_44601_(_26762_, _26806_, _26916_);
  or g_44602_(_26850_, _26861_, _26927_);
  or g_44603_(_26916_, _26927_, _26938_);
  or g_44604_(_26905_, _26938_, _26949_);
  xor g_44605_(out[284], out[620], _26960_);
  or g_44606_(_26707_, _26960_, _26971_);
  or g_44607_(_26696_, _26817_, _26982_);
  or g_44608_(_26971_, _26982_, _26993_);
  or g_44609_(_26740_, _26795_, _27004_);
  or g_44610_(_26828_, _27004_, _27015_);
  or g_44611_(_26993_, _27015_, _27026_);
  or g_44612_(_26949_, _27026_, _27037_);
  or g_44613_(_26872_, _27037_, _27048_);
  and g_44614_(out[267], _39922_, _27059_);
  xor g_44615_(out[260], out[612], _27070_);
  xor g_44616_(out[270], out[622], _27081_);
  or g_44617_(_27070_, _27081_, _27092_);
  xor g_44618_(out[269], out[621], _27103_);
  xor g_44619_(out[259], out[611], _27114_);
  xor g_44620_(out[256], out[608], _27125_);
  and g_44621_(_39680_, out[619], _27136_);
  xor g_44622_(out[266], out[618], _27147_);
  xor g_44623_(out[271], out[623], _27158_);
  xor g_44624_(out[262], out[614], _27169_);
  xor g_44625_(out[261], out[613], _27180_);
  xor g_44626_(out[264], out[616], _27191_);
  or g_44627_(_27103_, _27191_, _27202_);
  xor g_44628_(out[258], out[610], _27213_);
  xor g_44629_(out[265], out[617], _27224_);
  xor g_44630_(out[257], out[609], _27235_);
  or g_44631_(_27147_, _27213_, _27246_);
  or g_44632_(_27202_, _27246_, _27257_);
  or g_44633_(_27114_, _27224_, _27268_);
  or g_44634_(_27180_, _27268_, _27279_);
  or g_44635_(_27257_, _27279_, _27290_);
  or g_44636_(_27092_, _27290_, _27301_);
  xor g_44637_(out[268], out[620], _27312_);
  or g_44638_(_27136_, _27312_, _27323_);
  xor g_44639_(out[263], out[615], _27334_);
  or g_44640_(_27169_, _27334_, _27345_);
  or g_44641_(_27323_, _27345_, _27356_);
  or g_44642_(_27059_, _27235_, _27367_);
  or g_44643_(_27158_, _27367_, _27378_);
  or g_44644_(_27356_, _27378_, _27389_);
  or g_44645_(_27125_, _27389_, _27400_);
  or g_44646_(_27301_, _27400_, _27411_);
  xor g_44647_(out[247], out[615], _27422_);
  and g_44648_(_39669_, out[619], _27433_);
  xor g_44649_(out[254], out[622], _27444_);
  xor g_44650_(out[248], out[616], _27455_);
  xor g_44651_(out[241], out[609], _27466_);
  xor g_44652_(out[253], out[621], _27477_);
  xor g_44653_(out[249], out[617], _27488_);
  xor g_44654_(out[244], out[612], _27499_);
  xor g_44655_(out[242], out[610], _27510_);
  and g_44656_(out[251], _39922_, _27521_);
  xor g_44657_(out[243], out[611], _27532_);
  xor g_44658_(out[246], out[614], _27543_);
  xor g_44659_(out[255], out[623], _27554_);
  xor g_44660_(out[250], out[618], _27564_);
  xor g_44661_(out[245], out[613], _27575_);
  xor g_44662_(out[240], out[608], _27586_);
  or g_44663_(_27444_, _27499_, _27597_);
  or g_44664_(_27455_, _27477_, _27608_);
  or g_44665_(_27510_, _27564_, _27619_);
  or g_44666_(_27608_, _27619_, _27630_);
  or g_44667_(_27488_, _27532_, _27641_);
  or g_44668_(_27575_, _27586_, _27652_);
  or g_44669_(_27641_, _27652_, _27663_);
  or g_44670_(_27630_, _27663_, _27674_);
  xor g_44671_(out[252], out[620], _27685_);
  or g_44672_(_27433_, _27685_, _27696_);
  or g_44673_(_27422_, _27543_, _27707_);
  or g_44674_(_27696_, _27707_, _27718_);
  or g_44675_(_27466_, _27521_, _27729_);
  or g_44676_(_27554_, _27729_, _27740_);
  or g_44677_(_27718_, _27740_, _27751_);
  or g_44678_(_27674_, _27751_, _27762_);
  or g_44679_(_27597_, _27762_, _27773_);
  xor g_44680_(out[225], out[609], _27784_);
  and g_44681_(out[235], _39922_, _27795_);
  xor g_44682_(out[233], out[617], _27806_);
  xor g_44683_(out[224], out[608], _27817_);
  xor g_44684_(out[238], out[622], _27828_);
  xor g_44685_(out[228], out[612], _27839_);
  or g_44686_(_27828_, _27839_, _27850_);
  xor g_44687_(out[237], out[621], _27861_);
  xor g_44688_(out[227], out[611], _27872_);
  and g_44689_(_39658_, out[619], _27883_);
  xor g_44690_(out[230], out[614], _27894_);
  xor g_44691_(out[234], out[618], _27905_);
  xor g_44692_(out[229], out[613], _27916_);
  xor g_44693_(out[239], out[623], _27927_);
  xor g_44694_(out[232], out[616], _27938_);
  or g_44695_(_27861_, _27938_, _27949_);
  xor g_44696_(out[226], out[610], _27960_);
  or g_44697_(_27905_, _27960_, _27971_);
  or g_44698_(_27949_, _27971_, _27982_);
  or g_44699_(_27806_, _27872_, _27993_);
  or g_44700_(_27916_, _27993_, _28004_);
  or g_44701_(_27982_, _28004_, _28015_);
  or g_44702_(_27850_, _28015_, _28026_);
  xor g_44703_(out[236], out[620], _28037_);
  or g_44704_(_27883_, _28037_, _28048_);
  xor g_44705_(out[231], out[615], _28059_);
  or g_44706_(_27894_, _28059_, _28070_);
  or g_44707_(_28048_, _28070_, _28081_);
  or g_44708_(_27784_, _27795_, _28092_);
  or g_44709_(_27927_, _28092_, _28103_);
  or g_44710_(_28081_, _28103_, _28114_);
  or g_44711_(_27817_, _28114_, _28125_);
  or g_44712_(_28026_, _28125_, _28136_);
  xor g_44713_(out[215], out[615], _28147_);
  and g_44714_(_39647_, out[619], _28158_);
  xor g_44715_(out[222], out[622], _28169_);
  xor g_44716_(out[216], out[616], _28180_);
  xor g_44717_(out[209], out[609], _28191_);
  xor g_44718_(out[221], out[621], _28202_);
  xor g_44719_(out[217], out[617], _28213_);
  xor g_44720_(out[212], out[612], _28224_);
  xor g_44721_(out[210], out[610], _28235_);
  and g_44722_(out[219], _39922_, _28246_);
  xor g_44723_(out[211], out[611], _28257_);
  xor g_44724_(out[214], out[614], _28268_);
  xor g_44725_(out[223], out[623], _28279_);
  xor g_44726_(out[218], out[618], _28290_);
  xor g_44727_(out[213], out[613], _28301_);
  xor g_44728_(out[208], out[608], _28312_);
  or g_44729_(_28169_, _28224_, _28323_);
  or g_44730_(_28180_, _28202_, _28334_);
  or g_44731_(_28235_, _28290_, _28345_);
  or g_44732_(_28334_, _28345_, _28356_);
  or g_44733_(_28213_, _28257_, _28367_);
  or g_44734_(_28301_, _28312_, _28378_);
  or g_44735_(_28367_, _28378_, _28389_);
  or g_44736_(_28356_, _28389_, _28400_);
  xor g_44737_(out[220], out[620], _28411_);
  or g_44738_(_28158_, _28411_, _28422_);
  or g_44739_(_28147_, _28268_, _28433_);
  or g_44740_(_28422_, _28433_, _28444_);
  or g_44741_(_28191_, _28246_, _28455_);
  or g_44742_(_28279_, _28455_, _28466_);
  or g_44743_(_28444_, _28466_, _28477_);
  or g_44744_(_28400_, _28477_, _28488_);
  or g_44745_(_28323_, _28488_, _28499_);
  xor g_44746_(out[193], out[609], _28510_);
  and g_44747_(_39636_, out[619], _28521_);
  and g_44748_(out[203], _39922_, _28532_);
  xor g_44749_(out[201], out[617], _28543_);
  xor g_44750_(out[192], out[608], _28554_);
  xor g_44751_(out[206], out[622], _28565_);
  xor g_44752_(out[196], out[612], _28576_);
  or g_44753_(_28565_, _28576_, _28587_);
  xor g_44754_(out[205], out[621], _28598_);
  xor g_44755_(out[195], out[611], _28609_);
  xor g_44756_(out[204], out[620], _28620_);
  xor g_44757_(out[198], out[614], _28631_);
  xor g_44758_(out[202], out[618], _28642_);
  xor g_44759_(out[197], out[613], _28653_);
  xor g_44760_(out[207], out[623], _28664_);
  xor g_44761_(out[200], out[616], _28675_);
  or g_44762_(_28598_, _28675_, _28686_);
  xor g_44763_(out[194], out[610], _28697_);
  or g_44764_(_28642_, _28697_, _28708_);
  or g_44765_(_28686_, _28708_, _28719_);
  or g_44766_(_28543_, _28609_, _28730_);
  or g_44767_(_28653_, _28730_, _28740_);
  or g_44768_(_28719_, _28740_, _28751_);
  or g_44769_(_28587_, _28751_, _28762_);
  or g_44770_(_28521_, _28620_, _28773_);
  xor g_44771_(out[199], out[615], _28784_);
  or g_44772_(_28631_, _28784_, _28795_);
  or g_44773_(_28773_, _28795_, _28806_);
  or g_44774_(_28510_, _28532_, _28817_);
  or g_44775_(_28664_, _28817_, _28828_);
  or g_44776_(_28806_, _28828_, _28839_);
  or g_44777_(_28554_, _28839_, _28850_);
  or g_44778_(_28762_, _28850_, _28861_);
  xor g_44779_(out[183], out[615], _28872_);
  and g_44780_(_39625_, out[619], _28883_);
  xor g_44781_(out[190], out[622], _28894_);
  xor g_44782_(out[184], out[616], _28905_);
  xor g_44783_(out[177], out[609], _28916_);
  xor g_44784_(out[189], out[621], _28927_);
  xor g_44785_(out[185], out[617], _28938_);
  xor g_44786_(out[180], out[612], _28949_);
  xor g_44787_(out[178], out[610], _28960_);
  and g_44788_(out[187], _39922_, _28971_);
  xor g_44789_(out[179], out[611], _28982_);
  xor g_44790_(out[182], out[614], _28993_);
  xor g_44791_(out[191], out[623], _29004_);
  xor g_44792_(out[186], out[618], _29015_);
  xor g_44793_(out[181], out[613], _29026_);
  xor g_44794_(out[176], out[608], _29037_);
  or g_44795_(_28894_, _28949_, _29048_);
  or g_44796_(_28905_, _28927_, _29059_);
  or g_44797_(_28960_, _29015_, _29070_);
  or g_44798_(_29059_, _29070_, _29081_);
  or g_44799_(_28938_, _28982_, _29092_);
  or g_44800_(_29026_, _29037_, _29103_);
  or g_44801_(_29092_, _29103_, _29114_);
  or g_44802_(_29081_, _29114_, _29125_);
  xor g_44803_(out[188], out[620], _29136_);
  or g_44804_(_28883_, _29136_, _29147_);
  or g_44805_(_28872_, _28993_, _29158_);
  or g_44806_(_29147_, _29158_, _29169_);
  or g_44807_(_28916_, _28971_, _29180_);
  or g_44808_(_29004_, _29180_, _29191_);
  or g_44809_(_29169_, _29191_, _29202_);
  or g_44810_(_29125_, _29202_, _29213_);
  or g_44811_(_29048_, _29213_, _29224_);
  xor g_44812_(out[161], out[609], _29235_);
  and g_44813_(out[171], _39922_, _29246_);
  xor g_44814_(out[169], out[617], _29257_);
  xor g_44815_(out[160], out[608], _29268_);
  xor g_44816_(out[174], out[622], _29279_);
  xor g_44817_(out[164], out[612], _29290_);
  or g_44818_(_29279_, _29290_, _29301_);
  xor g_44819_(out[173], out[621], _29312_);
  xor g_44820_(out[163], out[611], _29323_);
  and g_44821_(_39614_, out[619], _29334_);
  xor g_44822_(out[166], out[614], _29345_);
  xor g_44823_(out[170], out[618], _29356_);
  xor g_44824_(out[165], out[613], _29367_);
  xor g_44825_(out[175], out[623], _29378_);
  xor g_44826_(out[168], out[616], _29389_);
  or g_44827_(_29312_, _29389_, _29400_);
  xor g_44828_(out[162], out[610], _29411_);
  or g_44829_(_29356_, _29411_, _29422_);
  or g_44830_(_29400_, _29422_, _29433_);
  or g_44831_(_29257_, _29323_, _29444_);
  or g_44832_(_29367_, _29444_, _29455_);
  or g_44833_(_29433_, _29455_, _29466_);
  or g_44834_(_29301_, _29466_, _29477_);
  xor g_44835_(out[172], out[620], _29488_);
  or g_44836_(_29334_, _29488_, _29499_);
  xor g_44837_(out[167], out[615], _29510_);
  or g_44838_(_29345_, _29510_, _29521_);
  or g_44839_(_29499_, _29521_, _29532_);
  or g_44840_(_29235_, _29246_, _29543_);
  or g_44841_(_29378_, _29543_, _29554_);
  or g_44842_(_29532_, _29554_, _29565_);
  or g_44843_(_29268_, _29565_, _29576_);
  or g_44844_(_29477_, _29576_, _29587_);
  xor g_44845_(out[151], out[615], _29598_);
  and g_44846_(_39603_, out[619], _29609_);
  xor g_44847_(out[158], out[622], _29620_);
  xor g_44848_(out[152], out[616], _29631_);
  xor g_44849_(out[145], out[609], _29642_);
  xor g_44850_(out[157], out[621], _29653_);
  xor g_44851_(out[153], out[617], _29664_);
  xor g_44852_(out[148], out[612], _29675_);
  xor g_44853_(out[146], out[610], _29686_);
  and g_44854_(out[155], _39922_, _29697_);
  xor g_44855_(out[147], out[611], _29708_);
  xor g_44856_(out[150], out[614], _29719_);
  xor g_44857_(out[159], out[623], _29730_);
  xor g_44858_(out[154], out[618], _29741_);
  xor g_44859_(out[149], out[613], _29752_);
  xor g_44860_(out[144], out[608], _29763_);
  or g_44861_(_29620_, _29675_, _29774_);
  or g_44862_(_29631_, _29653_, _29785_);
  or g_44863_(_29686_, _29741_, _29796_);
  or g_44864_(_29785_, _29796_, _29807_);
  or g_44865_(_29664_, _29708_, _29818_);
  or g_44866_(_29752_, _29763_, _29829_);
  or g_44867_(_29818_, _29829_, _29840_);
  or g_44868_(_29807_, _29840_, _29851_);
  xor g_44869_(out[156], out[620], _29862_);
  or g_44870_(_29609_, _29862_, _29873_);
  or g_44871_(_29598_, _29719_, _29884_);
  or g_44872_(_29873_, _29884_, _29895_);
  or g_44873_(_29642_, _29697_, _29906_);
  or g_44874_(_29730_, _29906_, _29917_);
  or g_44875_(_29895_, _29917_, _29928_);
  or g_44876_(_29851_, _29928_, _29939_);
  or g_44877_(_29774_, _29939_, _29949_);
  xor g_44878_(out[129], out[609], _29960_);
  and g_44879_(out[139], _39922_, _29971_);
  xor g_44880_(out[137], out[617], _29982_);
  xor g_44881_(out[128], out[608], _29993_);
  xor g_44882_(out[142], out[622], _30004_);
  xor g_44883_(out[132], out[612], _30015_);
  or g_44884_(_30004_, _30015_, _30026_);
  xor g_44885_(out[141], out[621], _30037_);
  xor g_44886_(out[131], out[611], _30048_);
  and g_44887_(_39592_, out[619], _30059_);
  xor g_44888_(out[134], out[614], _30070_);
  xor g_44889_(out[138], out[618], _30081_);
  xor g_44890_(out[133], out[613], _30092_);
  xor g_44891_(out[143], out[623], _30103_);
  xor g_44892_(out[136], out[616], _30114_);
  or g_44893_(_30037_, _30114_, _30125_);
  xor g_44894_(out[130], out[610], _30136_);
  or g_44895_(_30081_, _30136_, _30147_);
  or g_44896_(_30125_, _30147_, _30158_);
  or g_44897_(_29982_, _30048_, _30169_);
  or g_44898_(_30092_, _30169_, _30180_);
  or g_44899_(_30158_, _30180_, _30191_);
  or g_44900_(_30026_, _30191_, _30202_);
  xor g_44901_(out[140], out[620], _30213_);
  or g_44902_(_30059_, _30213_, _30224_);
  xor g_44903_(out[135], out[615], _30235_);
  or g_44904_(_30070_, _30235_, _30246_);
  or g_44905_(_30224_, _30246_, _30257_);
  or g_44906_(_29960_, _29971_, _30268_);
  or g_44907_(_30103_, _30268_, _30279_);
  or g_44908_(_30257_, _30279_, _30290_);
  or g_44909_(_29993_, _30290_, _30301_);
  or g_44910_(_30202_, _30301_, _30312_);
  xor g_44911_(out[119], out[615], _30323_);
  and g_44912_(_39581_, out[619], _30334_);
  xor g_44913_(out[126], out[622], _30345_);
  xor g_44914_(out[120], out[616], _30356_);
  xor g_44915_(out[113], out[609], _30367_);
  xor g_44916_(out[125], out[621], _30378_);
  xor g_44917_(out[121], out[617], _30389_);
  xor g_44918_(out[116], out[612], _30400_);
  xor g_44919_(out[114], out[610], _30411_);
  and g_44920_(out[123], _39922_, _30422_);
  xor g_44921_(out[115], out[611], _30433_);
  xor g_44922_(out[118], out[614], _30444_);
  xor g_44923_(out[127], out[623], _30455_);
  xor g_44924_(out[122], out[618], _30466_);
  xor g_44925_(out[117], out[613], _30477_);
  xor g_44926_(out[112], out[608], _30488_);
  or g_44927_(_30345_, _30400_, _30499_);
  or g_44928_(_30356_, _30378_, _30510_);
  or g_44929_(_30411_, _30466_, _30521_);
  or g_44930_(_30510_, _30521_, _30532_);
  or g_44931_(_30389_, _30433_, _30543_);
  or g_44932_(_30477_, _30488_, _30554_);
  or g_44933_(_30543_, _30554_, _30565_);
  or g_44934_(_30532_, _30565_, _30576_);
  xor g_44935_(out[124], out[620], _30587_);
  or g_44936_(_30334_, _30587_, _30598_);
  or g_44937_(_30323_, _30444_, _30609_);
  or g_44938_(_30598_, _30609_, _30620_);
  or g_44939_(_30367_, _30422_, _30631_);
  or g_44940_(_30455_, _30631_, _30642_);
  or g_44941_(_30620_, _30642_, _30653_);
  or g_44942_(_30576_, _30653_, _30664_);
  or g_44943_(_30499_, _30664_, _30675_);
  xor g_44944_(out[97], out[609], _30686_);
  and g_44945_(out[107], _39922_, _30697_);
  xor g_44946_(out[105], out[617], _30708_);
  xor g_44947_(out[96], out[608], _30719_);
  xor g_44948_(out[110], out[622], _30730_);
  xor g_44949_(out[100], out[612], _30741_);
  or g_44950_(_30730_, _30741_, _30752_);
  xor g_44951_(out[109], out[621], _30763_);
  xor g_44952_(out[99], out[611], _30774_);
  and g_44953_(_39570_, out[619], _30785_);
  xor g_44954_(out[102], out[614], _30796_);
  xor g_44955_(out[106], out[618], _30807_);
  xor g_44956_(out[101], out[613], _30818_);
  xor g_44957_(out[111], out[623], _30829_);
  xor g_44958_(out[104], out[616], _30840_);
  or g_44959_(_30763_, _30840_, _30851_);
  xor g_44960_(out[98], out[610], _30862_);
  or g_44961_(_30807_, _30862_, _30873_);
  or g_44962_(_30851_, _30873_, _30884_);
  or g_44963_(_30708_, _30774_, _30895_);
  or g_44964_(_30818_, _30895_, _30906_);
  or g_44965_(_30884_, _30906_, _30917_);
  or g_44966_(_30752_, _30917_, _30928_);
  xor g_44967_(out[108], out[620], _30939_);
  or g_44968_(_30785_, _30939_, _30950_);
  xor g_44969_(out[103], out[615], _30961_);
  or g_44970_(_30796_, _30961_, _30972_);
  or g_44971_(_30950_, _30972_, _30983_);
  or g_44972_(_30686_, _30697_, _30994_);
  or g_44973_(_30829_, _30994_, _31005_);
  or g_44974_(_30983_, _31005_, _31016_);
  or g_44975_(_30719_, _31016_, _31027_);
  or g_44976_(_30928_, _31027_, _31038_);
  xor g_44977_(out[87], out[615], _31049_);
  and g_44978_(_39559_, out[619], _31060_);
  xor g_44979_(out[94], out[622], _31071_);
  xor g_44980_(out[88], out[616], _31082_);
  xor g_44981_(out[81], out[609], _31093_);
  xor g_44982_(out[93], out[621], _31104_);
  xor g_44983_(out[89], out[617], _31115_);
  xor g_44984_(out[84], out[612], _31126_);
  xor g_44985_(out[82], out[610], _31137_);
  and g_44986_(out[91], _39922_, _31148_);
  xor g_44987_(out[83], out[611], _31159_);
  xor g_44988_(out[86], out[614], _31170_);
  xor g_44989_(out[95], out[623], _31181_);
  xor g_44990_(out[90], out[618], _31192_);
  xor g_44991_(out[85], out[613], _31202_);
  xor g_44992_(out[80], out[608], _31213_);
  or g_44993_(_31071_, _31126_, _31224_);
  or g_44994_(_31082_, _31104_, _31235_);
  or g_44995_(_31137_, _31192_, _31246_);
  or g_44996_(_31235_, _31246_, _31257_);
  or g_44997_(_31115_, _31159_, _31268_);
  or g_44998_(_31202_, _31213_, _31279_);
  or g_44999_(_31268_, _31279_, _31290_);
  or g_45000_(_31257_, _31290_, _31301_);
  xor g_45001_(out[92], out[620], _31312_);
  or g_45002_(_31060_, _31312_, _31323_);
  or g_45003_(_31049_, _31170_, _31334_);
  or g_45004_(_31323_, _31334_, _31345_);
  or g_45005_(_31093_, _31148_, _31356_);
  or g_45006_(_31181_, _31356_, _31367_);
  or g_45007_(_31345_, _31367_, _31378_);
  or g_45008_(_31301_, _31378_, _31389_);
  or g_45009_(_31224_, _31389_, _31400_);
  xor g_45010_(out[65], out[609], _31411_);
  and g_45011_(out[75], _39922_, _31422_);
  xor g_45012_(out[73], out[617], _31433_);
  xor g_45013_(out[64], out[608], _31444_);
  xor g_45014_(out[78], out[622], _31455_);
  xor g_45015_(out[68], out[612], _31466_);
  or g_45016_(_31455_, _31466_, _31477_);
  xor g_45017_(out[77], out[621], _31488_);
  xor g_45018_(out[67], out[611], _31499_);
  and g_45019_(_39548_, out[619], _31510_);
  xor g_45020_(out[70], out[614], _31521_);
  xor g_45021_(out[74], out[618], _31532_);
  xor g_45022_(out[69], out[613], _31543_);
  xor g_45023_(out[79], out[623], _31554_);
  xor g_45024_(out[72], out[616], _31565_);
  or g_45025_(_31488_, _31565_, _31576_);
  xor g_45026_(out[66], out[610], _31587_);
  or g_45027_(_31532_, _31587_, _31598_);
  or g_45028_(_31576_, _31598_, _31609_);
  or g_45029_(_31433_, _31499_, _31620_);
  or g_45030_(_31543_, _31620_, _31631_);
  or g_45031_(_31609_, _31631_, _31642_);
  or g_45032_(_31477_, _31642_, _31653_);
  xor g_45033_(out[76], out[620], _31664_);
  or g_45034_(_31510_, _31664_, _31675_);
  xor g_45035_(out[71], out[615], _31686_);
  or g_45036_(_31521_, _31686_, _31697_);
  or g_45037_(_31675_, _31697_, _31708_);
  or g_45038_(_31411_, _31422_, _31719_);
  or g_45039_(_31554_, _31719_, _31730_);
  or g_45040_(_31708_, _31730_, _31741_);
  or g_45041_(_31444_, _31741_, _31752_);
  or g_45042_(_31653_, _31752_, _31763_);
  xor g_45043_(out[55], out[615], _31774_);
  and g_45044_(_39537_, out[619], _31785_);
  xor g_45045_(out[62], out[622], _31796_);
  xor g_45046_(out[56], out[616], _31807_);
  xor g_45047_(out[49], out[609], _31818_);
  xor g_45048_(out[61], out[621], _31829_);
  xor g_45049_(out[57], out[617], _31840_);
  xor g_45050_(out[52], out[612], _31851_);
  xor g_45051_(out[50], out[610], _31862_);
  and g_45052_(out[59], _39922_, _31873_);
  xor g_45053_(out[51], out[611], _31884_);
  xor g_45054_(out[54], out[614], _31895_);
  xor g_45055_(out[63], out[623], _31906_);
  xor g_45056_(out[58], out[618], _31917_);
  xor g_45057_(out[53], out[613], _31928_);
  xor g_45058_(out[48], out[608], _31939_);
  or g_45059_(_31796_, _31851_, _31950_);
  or g_45060_(_31807_, _31829_, _31961_);
  or g_45061_(_31862_, _31917_, _31972_);
  or g_45062_(_31961_, _31972_, _31983_);
  or g_45063_(_31840_, _31884_, _31994_);
  or g_45064_(_31928_, _31939_, _32005_);
  or g_45065_(_31994_, _32005_, _32016_);
  or g_45066_(_31983_, _32016_, _32027_);
  xor g_45067_(out[60], out[620], _32038_);
  or g_45068_(_31785_, _32038_, _32049_);
  or g_45069_(_31774_, _31895_, _32060_);
  or g_45070_(_32049_, _32060_, _32071_);
  or g_45071_(_31818_, _31873_, _32082_);
  or g_45072_(_31906_, _32082_, _32093_);
  or g_45073_(_32071_, _32093_, _32104_);
  or g_45074_(_32027_, _32104_, _32115_);
  or g_45075_(_31950_, _32115_, _32126_);
  xor g_45076_(out[33], out[609], _32137_);
  and g_45077_(out[43], _39922_, _32148_);
  xor g_45078_(out[41], out[617], _32159_);
  xor g_45079_(out[32], out[608], _32170_);
  xor g_45080_(out[46], out[622], _32181_);
  xor g_45081_(out[36], out[612], _32192_);
  or g_45082_(_32181_, _32192_, _32203_);
  xor g_45083_(out[45], out[621], _32214_);
  xor g_45084_(out[35], out[611], _32225_);
  and g_45085_(_39526_, out[619], _32236_);
  xor g_45086_(out[38], out[614], _32247_);
  xor g_45087_(out[42], out[618], _32258_);
  xor g_45088_(out[37], out[613], _32269_);
  xor g_45089_(out[47], out[623], _32280_);
  xor g_45090_(out[40], out[616], _32291_);
  or g_45091_(_32214_, _32291_, _32302_);
  xor g_45092_(out[34], out[610], _32313_);
  or g_45093_(_32258_, _32313_, _32324_);
  or g_45094_(_32302_, _32324_, _32335_);
  or g_45095_(_32159_, _32225_, _32346_);
  or g_45096_(_32269_, _32346_, _32357_);
  or g_45097_(_32335_, _32357_, _32368_);
  or g_45098_(_32203_, _32368_, _32379_);
  xor g_45099_(out[44], out[620], _32390_);
  or g_45100_(_32236_, _32390_, _32401_);
  xor g_45101_(out[39], out[615], _32412_);
  or g_45102_(_32247_, _32412_, _32423_);
  or g_45103_(_32401_, _32423_, _32434_);
  or g_45104_(_32137_, _32148_, _32445_);
  or g_45105_(_32280_, _32445_, _32456_);
  or g_45106_(_32434_, _32456_, _32467_);
  or g_45107_(_32170_, _32467_, _32478_);
  or g_45108_(_32379_, _32478_, _32488_);
  xor g_45109_(out[23], out[615], _32499_);
  and g_45110_(_39493_, out[619], _32510_);
  xor g_45111_(out[30], out[622], _32521_);
  xor g_45112_(out[24], out[616], _32532_);
  xor g_45113_(out[17], out[609], _32543_);
  xor g_45114_(out[29], out[621], _32554_);
  xor g_45115_(out[25], out[617], _32565_);
  xor g_45116_(out[20], out[612], _32576_);
  xor g_45117_(out[18], out[610], _32587_);
  and g_45118_(out[27], _39922_, _32598_);
  xor g_45119_(out[19], out[611], _32609_);
  xor g_45120_(out[22], out[614], _32620_);
  xor g_45121_(out[31], out[623], _32631_);
  xor g_45122_(out[26], out[618], _32642_);
  xor g_45123_(out[21], out[613], _32653_);
  xor g_45124_(out[16], out[608], _32664_);
  or g_45125_(_32521_, _32576_, _32675_);
  or g_45126_(_32532_, _32554_, _32686_);
  or g_45127_(_32587_, _32642_, _32697_);
  or g_45128_(_32686_, _32697_, _32708_);
  or g_45129_(_32565_, _32609_, _32719_);
  or g_45130_(_32653_, _32664_, _32730_);
  or g_45131_(_32719_, _32730_, _32741_);
  or g_45132_(_32708_, _32741_, _32752_);
  xor g_45133_(out[28], out[620], _32763_);
  or g_45134_(_32510_, _32763_, _32774_);
  or g_45135_(_32499_, _32620_, _32785_);
  or g_45136_(_32774_, _32785_, _32796_);
  or g_45137_(_32543_, _32598_, _32807_);
  or g_45138_(_32631_, _32807_, _32818_);
  or g_45139_(_32796_, _32818_, _32829_);
  or g_45140_(_32752_, _32829_, _32840_);
  or g_45141_(_32675_, _32840_, _32851_);
  and g_45142_(out[11], _39922_, _32862_);
  xor g_45143_(out[4], out[612], _32873_);
  xor g_45144_(out[14], out[622], _32884_);
  or g_45145_(_32873_, _32884_, _32895_);
  xor g_45146_(out[13], out[621], _32906_);
  xor g_45147_(out[3], out[611], _32917_);
  xor g_45148_(out[0], out[608], _32928_);
  and g_45149_(_39438_, out[619], _32939_);
  xor g_45150_(out[10], out[618], _32950_);
  xor g_45151_(out[15], out[623], _32961_);
  xor g_45152_(out[6], out[614], _32972_);
  xor g_45153_(out[5], out[613], _32983_);
  xor g_45154_(out[8], out[616], _32994_);
  or g_45155_(_32906_, _32994_, _33005_);
  xor g_45156_(out[2], out[610], _33016_);
  xor g_45157_(out[9], out[617], _33027_);
  xor g_45158_(out[1], out[609], _33038_);
  or g_45159_(_32950_, _33016_, _33049_);
  or g_45160_(_33005_, _33049_, _33060_);
  or g_45161_(_32917_, _33027_, _33071_);
  or g_45162_(_32983_, _33071_, _33082_);
  or g_45163_(_33060_, _33082_, _33093_);
  or g_45164_(_32895_, _33093_, _33104_);
  xor g_45165_(out[12], out[620], _33115_);
  or g_45166_(_32939_, _33115_, _33126_);
  xor g_45167_(out[7], out[615], _33137_);
  or g_45168_(_32972_, _33137_, _33148_);
  or g_45169_(_33126_, _33148_, _33159_);
  or g_45170_(_32862_, _33038_, _33170_);
  or g_45171_(_32961_, _33170_, _33181_);
  or g_45172_(_33159_, _33181_, _33192_);
  or g_45173_(_32928_, _33192_, _33203_);
  or g_45174_(_33104_, _33203_, _33214_);
  not g_45175_(_33214_, _33225_);
  xor g_45176_(out[305], out[593], _33236_);
  and g_45177_(out[315], _39911_, _33247_);
  xor g_45178_(out[318], out[606], _33258_);
  xor g_45179_(out[307], out[595], _33269_);
  xor g_45180_(out[308], out[596], _33280_);
  xor g_45181_(out[306], out[594], _33291_);
  xor g_45182_(out[313], out[601], _33302_);
  xor g_45183_(out[304], out[592], _33313_);
  and g_45184_(_39724_, out[603], _33324_);
  xor g_45185_(out[310], out[598], _33335_);
  xor g_45186_(out[314], out[602], _33346_);
  xor g_45187_(out[309], out[597], _33357_);
  xor g_45188_(out[319], out[607], _33368_);
  xor g_45189_(out[317], out[605], _33379_);
  xor g_45190_(out[312], out[600], _33390_);
  or g_45191_(_33258_, _33280_, _33401_);
  or g_45192_(_33379_, _33390_, _33412_);
  or g_45193_(_33291_, _33346_, _33423_);
  or g_45194_(_33412_, _33423_, _33434_);
  or g_45195_(_33269_, _33302_, _33445_);
  or g_45196_(_33313_, _33357_, _33456_);
  or g_45197_(_33445_, _33456_, _33467_);
  or g_45198_(_33434_, _33467_, _33478_);
  xor g_45199_(out[316], out[604], _33489_);
  or g_45200_(_33324_, _33489_, _33500_);
  xor g_45201_(out[311], out[599], _33511_);
  or g_45202_(_33335_, _33511_, _33522_);
  or g_45203_(_33500_, _33522_, _33533_);
  or g_45204_(_33236_, _33247_, _33544_);
  or g_45205_(_33368_, _33544_, _33555_);
  or g_45206_(_33533_, _33555_, _33566_);
  or g_45207_(_33478_, _33566_, _33577_);
  or g_45208_(_33401_, _33577_, _33588_);
  xor g_45209_(out[295], out[599], _33599_);
  and g_45210_(_39702_, out[603], _33610_);
  xor g_45211_(out[302], out[606], _33621_);
  xor g_45212_(out[296], out[600], _33632_);
  xor g_45213_(out[289], out[593], _33643_);
  xor g_45214_(out[301], out[605], _33654_);
  xor g_45215_(out[297], out[601], _33665_);
  xor g_45216_(out[292], out[596], _33676_);
  xor g_45217_(out[290], out[594], _33686_);
  and g_45218_(out[299], _39911_, _33697_);
  xor g_45219_(out[291], out[595], _33708_);
  xor g_45220_(out[294], out[598], _33719_);
  xor g_45221_(out[303], out[607], _33730_);
  xor g_45222_(out[298], out[602], _33741_);
  xor g_45223_(out[293], out[597], _33752_);
  xor g_45224_(out[288], out[592], _33763_);
  or g_45225_(_33621_, _33676_, _33774_);
  or g_45226_(_33632_, _33654_, _33785_);
  or g_45227_(_33686_, _33741_, _33796_);
  or g_45228_(_33785_, _33796_, _33807_);
  or g_45229_(_33665_, _33708_, _33818_);
  or g_45230_(_33752_, _33763_, _33829_);
  or g_45231_(_33818_, _33829_, _33840_);
  or g_45232_(_33807_, _33840_, _33851_);
  xor g_45233_(out[300], out[604], _33862_);
  or g_45234_(_33610_, _33862_, _33873_);
  or g_45235_(_33599_, _33719_, _33884_);
  or g_45236_(_33873_, _33884_, _33895_);
  or g_45237_(_33643_, _33697_, _33906_);
  or g_45238_(_33730_, _33906_, _33917_);
  or g_45239_(_33895_, _33917_, _33928_);
  or g_45240_(_33851_, _33928_, _33939_);
  or g_45241_(_33774_, _33939_, _33950_);
  and g_45242_(out[283], _39911_, _33961_);
  and g_45243_(_39691_, out[603], _33972_);
  xor g_45244_(out[273], out[593], _33983_);
  xor g_45245_(out[275], out[595], _33994_);
  xor g_45246_(out[279], out[599], _34005_);
  xor g_45247_(out[281], out[601], _34016_);
  xor g_45248_(out[287], out[607], _34027_);
  xor g_45249_(out[274], out[594], _34038_);
  xor g_45250_(out[286], out[606], _34049_);
  xor g_45251_(out[285], out[605], _34060_);
  xor g_45252_(out[280], out[600], _34071_);
  or g_45253_(_34060_, _34071_, _34082_);
  xor g_45254_(out[276], out[596], _34093_);
  xor g_45255_(out[278], out[598], _34104_);
  xor g_45256_(out[282], out[602], _34115_);
  xor g_45257_(out[277], out[597], _34126_);
  xor g_45258_(out[272], out[592], _34137_);
  or g_45259_(_34038_, _34115_, _34148_);
  or g_45260_(_34082_, _34148_, _34159_);
  or g_45261_(_33994_, _34016_, _34170_);
  or g_45262_(_34126_, _34170_, _34181_);
  or g_45263_(_34159_, _34181_, _34192_);
  or g_45264_(_34049_, _34093_, _34203_);
  or g_45265_(_34192_, _34203_, _34214_);
  xor g_45266_(out[284], out[604], _34225_);
  or g_45267_(_33972_, _34225_, _34236_);
  or g_45268_(_34005_, _34104_, _34247_);
  or g_45269_(_34236_, _34247_, _34258_);
  or g_45270_(_33961_, _33983_, _34269_);
  or g_45271_(_34027_, _34269_, _34280_);
  or g_45272_(_34258_, _34280_, _34291_);
  or g_45273_(_34137_, _34291_, _34302_);
  or g_45274_(_34214_, _34302_, _34313_);
  not g_45275_(_34313_, _34324_);
  xor g_45276_(out[263], out[599], _34335_);
  and g_45277_(_39680_, out[603], _34346_);
  xor g_45278_(out[270], out[606], _34357_);
  xor g_45279_(out[264], out[600], _34368_);
  xor g_45280_(out[257], out[593], _34379_);
  xor g_45281_(out[269], out[605], _34390_);
  xor g_45282_(out[265], out[601], _34401_);
  xor g_45283_(out[260], out[596], _34412_);
  xor g_45284_(out[258], out[594], _34423_);
  and g_45285_(out[267], _39911_, _34434_);
  xor g_45286_(out[259], out[595], _34445_);
  xor g_45287_(out[262], out[598], _34456_);
  xor g_45288_(out[271], out[607], _34467_);
  xor g_45289_(out[266], out[602], _34478_);
  xor g_45290_(out[261], out[597], _34489_);
  xor g_45291_(out[256], out[592], _34500_);
  or g_45292_(_34357_, _34412_, _34511_);
  or g_45293_(_34368_, _34390_, _34522_);
  or g_45294_(_34423_, _34478_, _34533_);
  or g_45295_(_34522_, _34533_, _34544_);
  or g_45296_(_34401_, _34445_, _34555_);
  or g_45297_(_34489_, _34500_, _34566_);
  or g_45298_(_34555_, _34566_, _34577_);
  or g_45299_(_34544_, _34577_, _34588_);
  xor g_45300_(out[268], out[604], _34599_);
  or g_45301_(_34346_, _34599_, _34610_);
  or g_45302_(_34335_, _34456_, _34621_);
  or g_45303_(_34610_, _34621_, _34632_);
  or g_45304_(_34379_, _34434_, _34642_);
  or g_45305_(_34467_, _34642_, _34653_);
  or g_45306_(_34632_, _34653_, _34664_);
  or g_45307_(_34588_, _34664_, _34675_);
  or g_45308_(_34511_, _34675_, _34686_);
  xor g_45309_(out[250], out[602], _34697_);
  xor g_45310_(out[242], out[594], _34708_);
  xor g_45311_(out[241], out[593], _34719_);
  and g_45312_(_39669_, out[603], _34730_);
  and g_45313_(out[251], _39911_, _34741_);
  xor g_45314_(out[253], out[605], _34752_);
  xor g_45315_(out[243], out[595], _34763_);
  xor g_45316_(out[254], out[606], _34774_);
  xor g_45317_(out[252], out[604], _34785_);
  xor g_45318_(out[248], out[600], _34796_);
  xor g_45319_(out[255], out[607], _34807_);
  xor g_45320_(out[245], out[597], _34818_);
  xor g_45321_(out[246], out[598], _34829_);
  xor g_45322_(out[240], out[592], _34840_);
  xor g_45323_(out[244], out[596], _34851_);
  or g_45324_(_34752_, _34796_, _34862_);
  xor g_45325_(out[249], out[601], _34873_);
  or g_45326_(_34697_, _34708_, _34884_);
  or g_45327_(_34862_, _34884_, _34895_);
  or g_45328_(_34763_, _34873_, _34906_);
  or g_45329_(_34818_, _34906_, _34917_);
  or g_45330_(_34895_, _34917_, _34928_);
  or g_45331_(_34774_, _34851_, _34939_);
  or g_45332_(_34928_, _34939_, _34950_);
  or g_45333_(_34730_, _34785_, _34961_);
  xor g_45334_(out[247], out[599], _34972_);
  or g_45335_(_34829_, _34972_, _34983_);
  or g_45336_(_34961_, _34983_, _34986_);
  or g_45337_(_34719_, _34741_, _34987_);
  or g_45338_(_34807_, _34987_, _34988_);
  or g_45339_(_34986_, _34988_, _34989_);
  or g_45340_(_34840_, _34989_, _34990_);
  or g_45341_(_34950_, _34990_, _34991_);
  xor g_45342_(out[231], out[599], _34992_);
  and g_45343_(_39658_, out[603], _34993_);
  xor g_45344_(out[238], out[606], _34994_);
  xor g_45345_(out[232], out[600], _34995_);
  xor g_45346_(out[225], out[593], _34996_);
  xor g_45347_(out[237], out[605], _34997_);
  xor g_45348_(out[233], out[601], _34998_);
  xor g_45349_(out[228], out[596], _34999_);
  xor g_45350_(out[226], out[594], _35000_);
  and g_45351_(out[235], _39911_, _35001_);
  xor g_45352_(out[227], out[595], _35002_);
  xor g_45353_(out[230], out[598], _35003_);
  xor g_45354_(out[239], out[607], _35004_);
  xor g_45355_(out[234], out[602], _35005_);
  xor g_45356_(out[229], out[597], _35006_);
  xor g_45357_(out[224], out[592], _35007_);
  or g_45358_(_34994_, _34999_, _35008_);
  or g_45359_(_34995_, _34997_, _35009_);
  or g_45360_(_35000_, _35005_, _35010_);
  or g_45361_(_35009_, _35010_, _35011_);
  or g_45362_(_34998_, _35002_, _35012_);
  or g_45363_(_35006_, _35007_, _35013_);
  or g_45364_(_35012_, _35013_, _35014_);
  or g_45365_(_35011_, _35014_, _35015_);
  xor g_45366_(out[236], out[604], _35016_);
  or g_45367_(_34993_, _35016_, _35017_);
  or g_45368_(_34992_, _35003_, _35018_);
  or g_45369_(_35017_, _35018_, _35019_);
  or g_45370_(_34996_, _35001_, _35020_);
  or g_45371_(_35004_, _35020_, _35021_);
  or g_45372_(_35019_, _35021_, _35022_);
  or g_45373_(_35015_, _35022_, _35023_);
  or g_45374_(_35008_, _35023_, _35024_);
  xor g_45375_(out[216], out[600], _35025_);
  xor g_45376_(out[213], out[597], _35026_);
  xor g_45377_(out[211], out[595], _35027_);
  xor g_45378_(out[222], out[606], _35028_);
  xor g_45379_(out[221], out[605], _35029_);
  xor g_45380_(out[210], out[594], _35030_);
  xor g_45381_(out[217], out[601], _35031_);
  xor g_45382_(out[214], out[598], _35032_);
  xor g_45383_(out[223], out[607], _35033_);
  xor g_45384_(out[218], out[602], _35034_);
  xor g_45385_(out[212], out[596], _35035_);
  xor g_45386_(out[208], out[592], _35036_);
  and g_45387_(_39647_, out[603], _35037_);
  and g_45388_(out[219], _39911_, _35038_);
  or g_45389_(_35025_, _35029_, _35039_);
  xor g_45390_(out[209], out[593], _35040_);
  or g_45391_(_35030_, _35034_, _35041_);
  or g_45392_(_35039_, _35041_, _35042_);
  or g_45393_(_35027_, _35031_, _35043_);
  or g_45394_(_35026_, _35043_, _35044_);
  or g_45395_(_35042_, _35044_, _35045_);
  or g_45396_(_35028_, _35035_, _35046_);
  or g_45397_(_35045_, _35046_, _35047_);
  xor g_45398_(out[220], out[604], _35048_);
  or g_45399_(_35037_, _35048_, _35049_);
  xor g_45400_(out[215], out[599], _35050_);
  or g_45401_(_35032_, _35050_, _35051_);
  or g_45402_(_35049_, _35051_, _35052_);
  or g_45403_(_35038_, _35040_, _35053_);
  or g_45404_(_35033_, _35053_, _35054_);
  or g_45405_(_35052_, _35054_, _35055_);
  or g_45406_(_35036_, _35055_, _35056_);
  or g_45407_(_35047_, _35056_, _35057_);
  xor g_45408_(out[199], out[599], _35058_);
  and g_45409_(_39636_, out[603], _35059_);
  xor g_45410_(out[206], out[606], _35060_);
  xor g_45411_(out[200], out[600], _35061_);
  xor g_45412_(out[193], out[593], _35062_);
  xor g_45413_(out[205], out[605], _35063_);
  xor g_45414_(out[201], out[601], _35064_);
  xor g_45415_(out[196], out[596], _35065_);
  xor g_45416_(out[194], out[594], _35066_);
  and g_45417_(out[203], _39911_, _35067_);
  xor g_45418_(out[195], out[595], _35068_);
  xor g_45419_(out[198], out[598], _35069_);
  xor g_45420_(out[207], out[607], _35070_);
  xor g_45421_(out[202], out[602], _35071_);
  xor g_45422_(out[197], out[597], _35072_);
  xor g_45423_(out[192], out[592], _35073_);
  or g_45424_(_35060_, _35065_, _35074_);
  not g_45425_(_35074_, _35075_);
  or g_45426_(_35061_, _35063_, _35076_);
  or g_45427_(_35066_, _35071_, _35077_);
  or g_45428_(_35076_, _35077_, _35078_);
  or g_45429_(_35064_, _35068_, _35079_);
  or g_45430_(_35072_, _35073_, _35080_);
  or g_45431_(_35079_, _35080_, _35081_);
  or g_45432_(_35078_, _35081_, _35082_);
  xor g_45433_(out[204], out[604], _35083_);
  or g_45434_(_35059_, _35083_, _35084_);
  or g_45435_(_35058_, _35069_, _35085_);
  or g_45436_(_35084_, _35085_, _35086_);
  or g_45437_(_35062_, _35067_, _35087_);
  or g_45438_(_35070_, _35087_, _35088_);
  or g_45439_(_35086_, _35088_, _35089_);
  or g_45440_(_35082_, _35089_, _35090_);
  not g_45441_(_35090_, _35091_);
  and g_45442_(_35075_, _35091_, _35092_);
  not g_45443_(_35092_, _35093_);
  xor g_45444_(out[177], out[593], _35094_);
  and g_45445_(out[187], _39911_, _35095_);
  xor g_45446_(out[185], out[601], _35096_);
  xor g_45447_(out[176], out[592], _35097_);
  xor g_45448_(out[190], out[606], _35098_);
  xor g_45449_(out[180], out[596], _35099_);
  or g_45450_(_35098_, _35099_, _35100_);
  xor g_45451_(out[189], out[605], _35101_);
  xor g_45452_(out[179], out[595], _35102_);
  and g_45453_(_39625_, out[603], _35103_);
  xor g_45454_(out[182], out[598], _35104_);
  xor g_45455_(out[186], out[602], _35105_);
  xor g_45456_(out[181], out[597], _35106_);
  xor g_45457_(out[191], out[607], _35107_);
  xor g_45458_(out[184], out[600], _35108_);
  or g_45459_(_35101_, _35108_, _35109_);
  xor g_45460_(out[178], out[594], _35110_);
  or g_45461_(_35105_, _35110_, _35111_);
  or g_45462_(_35109_, _35111_, _35112_);
  or g_45463_(_35096_, _35102_, _35113_);
  or g_45464_(_35106_, _35113_, _35114_);
  or g_45465_(_35112_, _35114_, _35115_);
  or g_45466_(_35100_, _35115_, _35116_);
  xor g_45467_(out[188], out[604], _35117_);
  or g_45468_(_35103_, _35117_, _35118_);
  xor g_45469_(out[183], out[599], _35119_);
  or g_45470_(_35104_, _35119_, _35120_);
  or g_45471_(_35118_, _35120_, _35121_);
  or g_45472_(_35094_, _35095_, _35122_);
  or g_45473_(_35107_, _35122_, _35123_);
  or g_45474_(_35121_, _35123_, _35124_);
  or g_45475_(_35097_, _35124_, _35125_);
  or g_45476_(_35116_, _35125_, _35126_);
  xor g_45477_(out[167], out[599], _35127_);
  and g_45478_(_39614_, out[603], _35128_);
  xor g_45479_(out[174], out[606], _35129_);
  xor g_45480_(out[168], out[600], _35130_);
  xor g_45481_(out[161], out[593], _35131_);
  xor g_45482_(out[173], out[605], _35132_);
  xor g_45483_(out[169], out[601], _35133_);
  xor g_45484_(out[164], out[596], _35134_);
  xor g_45485_(out[162], out[594], _35135_);
  and g_45486_(out[171], _39911_, _35136_);
  xor g_45487_(out[163], out[595], _35137_);
  xor g_45488_(out[166], out[598], _35138_);
  xor g_45489_(out[175], out[607], _35139_);
  xor g_45490_(out[170], out[602], _35140_);
  xor g_45491_(out[165], out[597], _35141_);
  xor g_45492_(out[160], out[592], _35142_);
  or g_45493_(_35129_, _35134_, _35143_);
  or g_45494_(_35130_, _35132_, _35144_);
  or g_45495_(_35135_, _35140_, _35145_);
  or g_45496_(_35144_, _35145_, _35146_);
  or g_45497_(_35133_, _35137_, _35147_);
  or g_45498_(_35141_, _35142_, _35148_);
  or g_45499_(_35147_, _35148_, _35149_);
  or g_45500_(_35146_, _35149_, _35150_);
  xor g_45501_(out[172], out[604], _35151_);
  or g_45502_(_35128_, _35151_, _35152_);
  or g_45503_(_35127_, _35138_, _35153_);
  or g_45504_(_35152_, _35153_, _35154_);
  or g_45505_(_35131_, _35136_, _35155_);
  or g_45506_(_35139_, _35155_, _35156_);
  or g_45507_(_35154_, _35156_, _35157_);
  or g_45508_(_35150_, _35157_, _35158_);
  or g_45509_(_35143_, _35158_, _35159_);
  and g_45510_(out[155], _39911_, _35160_);
  and g_45511_(_39603_, out[603], _35161_);
  xor g_45512_(out[157], out[605], _35162_);
  xor g_45513_(out[159], out[607], _35163_);
  xor g_45514_(out[145], out[593], _35164_);
  xor g_45515_(out[148], out[596], _35165_);
  xor g_45516_(out[158], out[606], _35166_);
  or g_45517_(_35165_, _35166_, _35167_);
  xor g_45518_(out[152], out[600], _35168_);
  xor g_45519_(out[144], out[592], _35169_);
  xor g_45520_(out[146], out[594], _35170_);
  xor g_45521_(out[153], out[601], _35171_);
  xor g_45522_(out[149], out[597], _35172_);
  xor g_45523_(out[147], out[595], _35173_);
  xor g_45524_(out[154], out[602], _35174_);
  xor g_45525_(out[150], out[598], _35175_);
  or g_45526_(_35162_, _35168_, _35176_);
  or g_45527_(_35170_, _35174_, _35177_);
  or g_45528_(_35176_, _35177_, _35178_);
  or g_45529_(_35171_, _35173_, _35179_);
  or g_45530_(_35169_, _35172_, _35180_);
  or g_45531_(_35179_, _35180_, _35181_);
  or g_45532_(_35178_, _35181_, _35182_);
  xor g_45533_(out[156], out[604], _35183_);
  or g_45534_(_35161_, _35183_, _35184_);
  xor g_45535_(out[151], out[599], _35185_);
  or g_45536_(_35175_, _35185_, _35186_);
  or g_45537_(_35184_, _35186_, _35187_);
  or g_45538_(_35160_, _35164_, _35188_);
  or g_45539_(_35163_, _35188_, _35189_);
  or g_45540_(_35187_, _35189_, _35190_);
  or g_45541_(_35182_, _35190_, _35191_);
  or g_45542_(_35167_, _35191_, _35192_);
  not g_45543_(_35192_, _35193_);
  xor g_45544_(out[135], out[599], _35194_);
  and g_45545_(_39592_, out[603], _35195_);
  xor g_45546_(out[142], out[606], _35196_);
  xor g_45547_(out[136], out[600], _35197_);
  xor g_45548_(out[129], out[593], _35198_);
  xor g_45549_(out[141], out[605], _35199_);
  xor g_45550_(out[137], out[601], _35200_);
  xor g_45551_(out[132], out[596], _35201_);
  xor g_45552_(out[130], out[594], _35202_);
  and g_45553_(out[139], _39911_, _35203_);
  xor g_45554_(out[131], out[595], _35204_);
  xor g_45555_(out[134], out[598], _35205_);
  xor g_45556_(out[143], out[607], _35206_);
  xor g_45557_(out[138], out[602], _35207_);
  xor g_45558_(out[133], out[597], _35208_);
  xor g_45559_(out[128], out[592], _35209_);
  or g_45560_(_35196_, _35201_, _35210_);
  or g_45561_(_35197_, _35199_, _35211_);
  or g_45562_(_35202_, _35207_, _35212_);
  or g_45563_(_35211_, _35212_, _35213_);
  or g_45564_(_35200_, _35204_, _35214_);
  or g_45565_(_35208_, _35209_, _35215_);
  or g_45566_(_35214_, _35215_, _35216_);
  or g_45567_(_35213_, _35216_, _35217_);
  xor g_45568_(out[140], out[604], _35218_);
  or g_45569_(_35195_, _35218_, _35219_);
  or g_45570_(_35194_, _35205_, _35220_);
  or g_45571_(_35219_, _35220_, _35221_);
  or g_45572_(_35198_, _35203_, _35222_);
  or g_45573_(_35206_, _35222_, _35223_);
  or g_45574_(_35221_, _35223_, _35224_);
  or g_45575_(_35217_, _35224_, _35225_);
  or g_45576_(_35210_, _35225_, _35226_);
  and g_45577_(out[123], _39911_, _35227_);
  and g_45578_(_39581_, out[603], _35228_);
  xor g_45579_(out[125], out[605], _35229_);
  xor g_45580_(out[122], out[602], _35230_);
  xor g_45581_(out[117], out[597], _35231_);
  xor g_45582_(out[124], out[604], _35232_);
  xor g_45583_(out[112], out[592], _35233_);
  xor g_45584_(out[114], out[594], _35234_);
  xor g_45585_(out[115], out[595], _35235_);
  xor g_45586_(out[121], out[601], _35236_);
  xor g_45587_(out[126], out[606], _35237_);
  xor g_45588_(out[127], out[607], _35238_);
  xor g_45589_(out[113], out[593], _35239_);
  xor g_45590_(out[118], out[598], _35240_);
  xor g_45591_(out[116], out[596], _35241_);
  xor g_45592_(out[120], out[600], _35242_);
  or g_45593_(_35229_, _35242_, _35243_);
  or g_45594_(_35230_, _35234_, _35244_);
  or g_45595_(_35243_, _35244_, _35245_);
  or g_45596_(_35235_, _35236_, _35246_);
  or g_45597_(_35231_, _35246_, _35247_);
  or g_45598_(_35245_, _35247_, _35248_);
  or g_45599_(_35237_, _35241_, _35249_);
  or g_45600_(_35248_, _35249_, _35250_);
  or g_45601_(_35228_, _35232_, _35251_);
  xor g_45602_(out[119], out[599], _35252_);
  or g_45603_(_35240_, _35252_, _35253_);
  or g_45604_(_35251_, _35253_, _35254_);
  or g_45605_(_35227_, _35239_, _35255_);
  or g_45606_(_35238_, _35255_, _35256_);
  or g_45607_(_35254_, _35256_, _35257_);
  or g_45608_(_35233_, _35257_, _35258_);
  or g_45609_(_35250_, _35258_, _35259_);
  xor g_45610_(out[103], out[599], _35260_);
  and g_45611_(_39570_, out[603], _35261_);
  xor g_45612_(out[110], out[606], _35262_);
  xor g_45613_(out[104], out[600], _35263_);
  xor g_45614_(out[97], out[593], _35264_);
  xor g_45615_(out[109], out[605], _35265_);
  xor g_45616_(out[105], out[601], _35266_);
  xor g_45617_(out[100], out[596], _35267_);
  xor g_45618_(out[98], out[594], _35268_);
  and g_45619_(out[107], _39911_, _35269_);
  xor g_45620_(out[99], out[595], _35270_);
  xor g_45621_(out[102], out[598], _35271_);
  xor g_45622_(out[111], out[607], _35272_);
  xor g_45623_(out[106], out[602], _35273_);
  xor g_45624_(out[101], out[597], _35274_);
  xor g_45625_(out[96], out[592], _35275_);
  or g_45626_(_35262_, _35267_, _35276_);
  or g_45627_(_35263_, _35265_, _35277_);
  or g_45628_(_35268_, _35273_, _35278_);
  or g_45629_(_35277_, _35278_, _35279_);
  or g_45630_(_35266_, _35270_, _35280_);
  or g_45631_(_35274_, _35275_, _35281_);
  or g_45632_(_35280_, _35281_, _35282_);
  or g_45633_(_35279_, _35282_, _35283_);
  xor g_45634_(out[108], out[604], _35284_);
  or g_45635_(_35261_, _35284_, _35285_);
  or g_45636_(_35260_, _35271_, _35286_);
  or g_45637_(_35285_, _35286_, _35287_);
  or g_45638_(_35264_, _35269_, _35288_);
  or g_45639_(_35272_, _35288_, _35289_);
  or g_45640_(_35287_, _35289_, _35290_);
  or g_45641_(_35283_, _35290_, _35291_);
  or g_45642_(_35276_, _35291_, _35292_);
  xor g_45643_(out[81], out[593], _35293_);
  and g_45644_(out[91], _39911_, _35294_);
  xor g_45645_(out[89], out[601], _35295_);
  xor g_45646_(out[80], out[592], _35296_);
  xor g_45647_(out[94], out[606], _35297_);
  xor g_45648_(out[84], out[596], _35298_);
  or g_45649_(_35297_, _35298_, _35299_);
  xor g_45650_(out[93], out[605], _35300_);
  xor g_45651_(out[83], out[595], _35301_);
  and g_45652_(_39559_, out[603], _35302_);
  xor g_45653_(out[86], out[598], _35303_);
  xor g_45654_(out[90], out[602], _35304_);
  xor g_45655_(out[85], out[597], _35305_);
  xor g_45656_(out[95], out[607], _35306_);
  xor g_45657_(out[88], out[600], _35307_);
  or g_45658_(_35300_, _35307_, _35308_);
  xor g_45659_(out[82], out[594], _35309_);
  or g_45660_(_35304_, _35309_, _35310_);
  or g_45661_(_35308_, _35310_, _35311_);
  or g_45662_(_35295_, _35301_, _35312_);
  or g_45663_(_35305_, _35312_, _35313_);
  or g_45664_(_35311_, _35313_, _35314_);
  or g_45665_(_35299_, _35314_, _35315_);
  xor g_45666_(out[92], out[604], _35316_);
  or g_45667_(_35302_, _35316_, _35317_);
  xor g_45668_(out[87], out[599], _35318_);
  or g_45669_(_35303_, _35318_, _35319_);
  or g_45670_(_35317_, _35319_, _35320_);
  or g_45671_(_35293_, _35294_, _35321_);
  or g_45672_(_35306_, _35321_, _35322_);
  or g_45673_(_35320_, _35322_, _35323_);
  or g_45674_(_35296_, _35323_, _35324_);
  or g_45675_(_35315_, _35324_, _35325_);
  xor g_45676_(out[71], out[599], _35326_);
  and g_45677_(_39548_, out[603], _35327_);
  xor g_45678_(out[78], out[606], _35328_);
  xor g_45679_(out[72], out[600], _35329_);
  xor g_45680_(out[65], out[593], _35330_);
  xor g_45681_(out[77], out[605], _35331_);
  xor g_45682_(out[73], out[601], _35332_);
  xor g_45683_(out[68], out[596], _35333_);
  xor g_45684_(out[66], out[594], _35334_);
  and g_45685_(out[75], _39911_, _35335_);
  xor g_45686_(out[67], out[595], _35336_);
  xor g_45687_(out[70], out[598], _35337_);
  xor g_45688_(out[79], out[607], _35338_);
  xor g_45689_(out[74], out[602], _35339_);
  xor g_45690_(out[69], out[597], _35340_);
  xor g_45691_(out[64], out[592], _35341_);
  or g_45692_(_35328_, _35333_, _35342_);
  or g_45693_(_35329_, _35331_, _35343_);
  or g_45694_(_35334_, _35339_, _35344_);
  or g_45695_(_35343_, _35344_, _35345_);
  or g_45696_(_35332_, _35336_, _35346_);
  or g_45697_(_35340_, _35341_, _35347_);
  or g_45698_(_35346_, _35347_, _35348_);
  or g_45699_(_35345_, _35348_, _35349_);
  xor g_45700_(out[76], out[604], _35350_);
  or g_45701_(_35327_, _35350_, _35351_);
  or g_45702_(_35326_, _35337_, _35352_);
  or g_45703_(_35351_, _35352_, _35353_);
  or g_45704_(_35330_, _35335_, _35354_);
  or g_45705_(_35338_, _35354_, _35355_);
  or g_45706_(_35353_, _35355_, _35356_);
  or g_45707_(_35349_, _35356_, _35357_);
  or g_45708_(_35342_, _35357_, _35358_);
  xor g_45709_(out[58], out[602], _35359_);
  xor g_45710_(out[50], out[594], _35360_);
  xor g_45711_(out[49], out[593], _35361_);
  and g_45712_(_39537_, out[603], _35362_);
  and g_45713_(out[59], _39911_, _35363_);
  xor g_45714_(out[61], out[605], _35364_);
  xor g_45715_(out[51], out[595], _35365_);
  xor g_45716_(out[62], out[606], _35366_);
  xor g_45717_(out[60], out[604], _35367_);
  xor g_45718_(out[56], out[600], _35368_);
  xor g_45719_(out[63], out[607], _35369_);
  xor g_45720_(out[53], out[597], _35370_);
  xor g_45721_(out[54], out[598], _35371_);
  xor g_45722_(out[48], out[592], _35372_);
  xor g_45723_(out[52], out[596], _35373_);
  or g_45724_(_35364_, _35368_, _35374_);
  xor g_45725_(out[57], out[601], _35375_);
  or g_45726_(_35359_, _35360_, _35376_);
  or g_45727_(_35374_, _35376_, _35377_);
  or g_45728_(_35365_, _35375_, _35378_);
  or g_45729_(_35370_, _35378_, _35379_);
  or g_45730_(_35377_, _35379_, _35380_);
  or g_45731_(_35366_, _35373_, _35381_);
  or g_45732_(_35380_, _35381_, _35382_);
  or g_45733_(_35362_, _35367_, _35383_);
  xor g_45734_(out[55], out[599], _35384_);
  or g_45735_(_35371_, _35384_, _35385_);
  or g_45736_(_35383_, _35385_, _35386_);
  or g_45737_(_35361_, _35363_, _35387_);
  or g_45738_(_35369_, _35387_, _35388_);
  or g_45739_(_35386_, _35388_, _35389_);
  or g_45740_(_35372_, _35389_, _35390_);
  or g_45741_(_35382_, _35390_, _35391_);
  not g_45742_(_35391_, _35392_);
  xor g_45743_(out[39], out[599], _35393_);
  and g_45744_(_39526_, out[603], _35394_);
  xor g_45745_(out[46], out[606], _35395_);
  xor g_45746_(out[40], out[600], _35396_);
  xor g_45747_(out[33], out[593], _35397_);
  xor g_45748_(out[45], out[605], _35398_);
  xor g_45749_(out[41], out[601], _35399_);
  xor g_45750_(out[36], out[596], _35400_);
  xor g_45751_(out[34], out[594], _35401_);
  and g_45752_(out[43], _39911_, _35402_);
  xor g_45753_(out[35], out[595], _35403_);
  xor g_45754_(out[38], out[598], _35404_);
  xor g_45755_(out[47], out[607], _35405_);
  xor g_45756_(out[42], out[602], _35406_);
  xor g_45757_(out[37], out[597], _35407_);
  xor g_45758_(out[32], out[592], _35408_);
  or g_45759_(_35395_, _35400_, _35409_);
  or g_45760_(_35396_, _35398_, _35410_);
  or g_45761_(_35401_, _35406_, _35411_);
  or g_45762_(_35410_, _35411_, _35412_);
  or g_45763_(_35399_, _35403_, _35413_);
  or g_45764_(_35407_, _35408_, _35414_);
  or g_45765_(_35413_, _35414_, _35415_);
  or g_45766_(_35412_, _35415_, _35416_);
  xor g_45767_(out[44], out[604], _35417_);
  or g_45768_(_35394_, _35417_, _35418_);
  or g_45769_(_35393_, _35404_, _35419_);
  or g_45770_(_35418_, _35419_, _35420_);
  or g_45771_(_35397_, _35402_, _35421_);
  or g_45772_(_35405_, _35421_, _35422_);
  or g_45773_(_35420_, _35422_, _35423_);
  or g_45774_(_35416_, _35423_, _35424_);
  or g_45775_(_35409_, _35424_, _35425_);
  not g_45776_(_35425_, _35426_);
  xor g_45777_(out[28], out[604], _35427_);
  and g_45778_(_39493_, out[603], _35428_);
  xor g_45779_(out[24], out[600], _35429_);
  xor g_45780_(out[22], out[598], _35430_);
  xor g_45781_(out[29], out[605], _35431_);
  xor g_45782_(out[30], out[606], _35432_);
  xor g_45783_(out[18], out[594], _35433_);
  xor g_45784_(out[25], out[601], _35434_);
  xor g_45785_(out[21], out[597], _35435_);
  xor g_45786_(out[17], out[593], _35436_);
  and g_45787_(out[27], _39911_, _35437_);
  or g_45788_(_35429_, _35431_, _35438_);
  xor g_45789_(out[31], out[607], _35439_);
  xor g_45790_(out[26], out[602], _35440_);
  xor g_45791_(out[20], out[596], _35441_);
  xor g_45792_(out[19], out[595], _35442_);
  xor g_45793_(out[16], out[592], _35443_);
  or g_45794_(_35433_, _35440_, _35444_);
  or g_45795_(_35438_, _35444_, _35445_);
  or g_45796_(_35434_, _35442_, _35446_);
  or g_45797_(_35435_, _35446_, _35447_);
  or g_45798_(_35445_, _35447_, _35448_);
  or g_45799_(_35432_, _35441_, _35449_);
  or g_45800_(_35448_, _35449_, _35450_);
  or g_45801_(_35427_, _35428_, _35451_);
  xor g_45802_(out[23], out[599], _35452_);
  or g_45803_(_35430_, _35452_, _35453_);
  or g_45804_(_35451_, _35453_, _35454_);
  or g_45805_(_35436_, _35437_, _35455_);
  or g_45806_(_35439_, _35455_, _35456_);
  or g_45807_(_35454_, _35456_, _35457_);
  or g_45808_(_35443_, _35457_, _35458_);
  or g_45809_(_35450_, _35458_, _35459_);
  not g_45810_(_35459_, _35460_);
  xor g_45811_(out[1], out[593], _35461_);
  and g_45812_(_39438_, out[603], _35462_);
  and g_45813_(out[11], _39911_, _35463_);
  xor g_45814_(out[9], out[601], _35464_);
  xor g_45815_(out[0], out[592], _35465_);
  xor g_45816_(out[14], out[606], _35466_);
  xor g_45817_(out[4], out[596], _35467_);
  or g_45818_(_35466_, _35467_, _35468_);
  xor g_45819_(out[13], out[605], _35469_);
  xor g_45820_(out[3], out[595], _35470_);
  xor g_45821_(out[12], out[604], _35471_);
  xor g_45822_(out[6], out[598], _35472_);
  xor g_45823_(out[10], out[602], _35473_);
  xor g_45824_(out[5], out[597], _35474_);
  xor g_45825_(out[15], out[607], _35475_);
  xor g_45826_(out[8], out[600], _35476_);
  or g_45827_(_35469_, _35476_, _35477_);
  xor g_45828_(out[2], out[594], _35478_);
  or g_45829_(_35473_, _35478_, _35479_);
  or g_45830_(_35477_, _35479_, _35480_);
  or g_45831_(_35464_, _35470_, _35481_);
  or g_45832_(_35474_, _35481_, _35482_);
  or g_45833_(_35480_, _35482_, _35483_);
  or g_45834_(_35468_, _35483_, _35484_);
  or g_45835_(_35462_, _35471_, _35485_);
  xor g_45836_(out[7], out[599], _35486_);
  or g_45837_(_35472_, _35486_, _35487_);
  or g_45838_(_35485_, _35487_, _35488_);
  or g_45839_(_35461_, _35463_, _35489_);
  or g_45840_(_35475_, _35489_, _35490_);
  or g_45841_(_35488_, _35490_, _35491_);
  or g_45842_(_35465_, _35491_, _35492_);
  or g_45843_(_35484_, _35492_, _35493_);
  xor g_45844_(out[311], out[583], _35494_);
  and g_45845_(_39724_, out[587], _35495_);
  xor g_45846_(out[318], out[590], _35496_);
  xor g_45847_(out[312], out[584], _35497_);
  xor g_45848_(out[305], out[577], _35498_);
  xor g_45849_(out[317], out[589], _35499_);
  xor g_45850_(out[313], out[585], _35500_);
  xor g_45851_(out[308], out[580], _35501_);
  xor g_45852_(out[306], out[578], _35502_);
  and g_45853_(out[315], _39900_, _35503_);
  xor g_45854_(out[307], out[579], _35504_);
  xor g_45855_(out[310], out[582], _35505_);
  xor g_45856_(out[319], out[591], _35506_);
  xor g_45857_(out[314], out[586], _35507_);
  xor g_45858_(out[309], out[581], _35508_);
  xor g_45859_(out[304], out[576], _35509_);
  or g_45860_(_35496_, _35501_, _35510_);
  or g_45861_(_35497_, _35499_, _35511_);
  or g_45862_(_35502_, _35507_, _35512_);
  or g_45863_(_35511_, _35512_, _35513_);
  or g_45864_(_35500_, _35504_, _35514_);
  or g_45865_(_35508_, _35509_, _35515_);
  or g_45866_(_35514_, _35515_, _35516_);
  or g_45867_(_35513_, _35516_, _35517_);
  xor g_45868_(out[316], out[588], _35518_);
  or g_45869_(_35495_, _35518_, _35519_);
  or g_45870_(_35494_, _35505_, _35520_);
  or g_45871_(_35519_, _35520_, _35521_);
  or g_45872_(_35498_, _35503_, _35522_);
  or g_45873_(_35506_, _35522_, _35523_);
  or g_45874_(_35521_, _35523_, _35524_);
  or g_45875_(_35517_, _35524_, _35525_);
  or g_45876_(_35510_, _35525_, _35526_);
  and g_45877_(out[299], _39900_, _35527_);
  xor g_45878_(out[292], out[580], _35528_);
  xor g_45879_(out[302], out[590], _35529_);
  or g_45880_(_35528_, _35529_, _35530_);
  xor g_45881_(out[301], out[589], _35531_);
  xor g_45882_(out[291], out[579], _35532_);
  xor g_45883_(out[288], out[576], _35533_);
  and g_45884_(_39702_, out[587], _35534_);
  xor g_45885_(out[298], out[586], _35535_);
  xor g_45886_(out[303], out[591], _35536_);
  xor g_45887_(out[294], out[582], _35537_);
  xor g_45888_(out[293], out[581], _35538_);
  xor g_45889_(out[296], out[584], _35539_);
  or g_45890_(_35531_, _35539_, _35540_);
  xor g_45891_(out[290], out[578], _35541_);
  xor g_45892_(out[297], out[585], _35542_);
  xor g_45893_(out[289], out[577], _35543_);
  or g_45894_(_35535_, _35541_, _35544_);
  or g_45895_(_35540_, _35544_, _35545_);
  or g_45896_(_35532_, _35542_, _35546_);
  or g_45897_(_35538_, _35546_, _35547_);
  or g_45898_(_35545_, _35547_, _35548_);
  or g_45899_(_35530_, _35548_, _35549_);
  xor g_45900_(out[300], out[588], _35550_);
  or g_45901_(_35534_, _35550_, _35551_);
  xor g_45902_(out[295], out[583], _35552_);
  or g_45903_(_35537_, _35552_, _35553_);
  or g_45904_(_35551_, _35553_, _35554_);
  or g_45905_(_35527_, _35543_, _35555_);
  or g_45906_(_35536_, _35555_, _35556_);
  or g_45907_(_35554_, _35556_, _35557_);
  or g_45908_(_35533_, _35557_, _35558_);
  or g_45909_(_35549_, _35558_, _35559_);
  xor g_45910_(out[279], out[583], _35560_);
  and g_45911_(_39691_, out[587], _35561_);
  xor g_45912_(out[286], out[590], _35562_);
  xor g_45913_(out[280], out[584], _35563_);
  xor g_45914_(out[273], out[577], _35564_);
  xor g_45915_(out[285], out[589], _35565_);
  xor g_45916_(out[281], out[585], _35566_);
  xor g_45917_(out[276], out[580], _35567_);
  xor g_45918_(out[274], out[578], _35568_);
  and g_45919_(out[283], _39900_, _35569_);
  xor g_45920_(out[275], out[579], _35570_);
  xor g_45921_(out[278], out[582], _35571_);
  xor g_45922_(out[287], out[591], _35572_);
  xor g_45923_(out[282], out[586], _35573_);
  xor g_45924_(out[277], out[581], _35574_);
  xor g_45925_(out[272], out[576], _35575_);
  or g_45926_(_35562_, _35567_, _35576_);
  or g_45927_(_35563_, _35565_, _35577_);
  or g_45928_(_35568_, _35573_, _35578_);
  or g_45929_(_35577_, _35578_, _35579_);
  or g_45930_(_35566_, _35570_, _35580_);
  or g_45931_(_35574_, _35575_, _35581_);
  or g_45932_(_35580_, _35581_, _35582_);
  or g_45933_(_35579_, _35582_, _35583_);
  xor g_45934_(out[284], out[588], _35584_);
  or g_45935_(_35561_, _35584_, _35585_);
  or g_45936_(_35560_, _35571_, _35586_);
  or g_45937_(_35585_, _35586_, _35587_);
  or g_45938_(_35564_, _35569_, _35588_);
  or g_45939_(_35572_, _35588_, _35589_);
  or g_45940_(_35587_, _35589_, _35590_);
  or g_45941_(_35583_, _35590_, _35591_);
  or g_45942_(_35576_, _35591_, _35592_);
  not g_45943_(_35592_, _35593_);
  xor g_45944_(out[257], out[577], _35594_);
  and g_45945_(_39680_, out[587], _35595_);
  and g_45946_(out[267], _39900_, _35596_);
  xor g_45947_(out[265], out[585], _35597_);
  xor g_45948_(out[256], out[576], _35598_);
  xor g_45949_(out[270], out[590], _35599_);
  xor g_45950_(out[260], out[580], _35600_);
  or g_45951_(_35599_, _35600_, _35601_);
  xor g_45952_(out[269], out[589], _35602_);
  xor g_45953_(out[259], out[579], _35603_);
  xor g_45954_(out[268], out[588], _35604_);
  xor g_45955_(out[262], out[582], _35605_);
  xor g_45956_(out[266], out[586], _35606_);
  xor g_45957_(out[261], out[581], _35607_);
  xor g_45958_(out[271], out[591], _35608_);
  xor g_45959_(out[264], out[584], _35609_);
  or g_45960_(_35602_, _35609_, _35610_);
  xor g_45961_(out[258], out[578], _35611_);
  or g_45962_(_35606_, _35611_, _35612_);
  or g_45963_(_35610_, _35612_, _35613_);
  or g_45964_(_35597_, _35603_, _35614_);
  or g_45965_(_35607_, _35614_, _35615_);
  or g_45966_(_35613_, _35615_, _35616_);
  or g_45967_(_35601_, _35616_, _35617_);
  or g_45968_(_35595_, _35604_, _35618_);
  xor g_45969_(out[263], out[583], _35619_);
  or g_45970_(_35605_, _35619_, _35620_);
  or g_45971_(_35618_, _35620_, _35621_);
  or g_45972_(_35594_, _35596_, _35622_);
  or g_45973_(_35608_, _35622_, _35623_);
  or g_45974_(_35621_, _35623_, _35624_);
  or g_45975_(_35598_, _35624_, _35625_);
  or g_45976_(_35617_, _35625_, _35626_);
  not g_45977_(_35626_, _35627_);
  xor g_45978_(out[247], out[583], _35628_);
  and g_45979_(_39669_, out[587], _35629_);
  xor g_45980_(out[254], out[590], _35630_);
  xor g_45981_(out[248], out[584], _35631_);
  xor g_45982_(out[241], out[577], _35632_);
  xor g_45983_(out[253], out[589], _35633_);
  xor g_45984_(out[249], out[585], _35634_);
  xor g_45985_(out[244], out[580], _35635_);
  xor g_45986_(out[242], out[578], _35636_);
  and g_45987_(out[251], _39900_, _35637_);
  xor g_45988_(out[243], out[579], _35638_);
  xor g_45989_(out[246], out[582], _35639_);
  xor g_45990_(out[255], out[591], _35640_);
  xor g_45991_(out[250], out[586], _35641_);
  xor g_45992_(out[245], out[581], _35642_);
  xor g_45993_(out[240], out[576], _35643_);
  or g_45994_(_35630_, _35635_, _35644_);
  or g_45995_(_35631_, _35633_, _35645_);
  or g_45996_(_35636_, _35641_, _35646_);
  or g_45997_(_35645_, _35646_, _35647_);
  or g_45998_(_35634_, _35638_, _35648_);
  or g_45999_(_35642_, _35643_, _35649_);
  or g_46000_(_35648_, _35649_, _35650_);
  or g_46001_(_35647_, _35650_, _35651_);
  xor g_46002_(out[252], out[588], _35652_);
  or g_46003_(_35629_, _35652_, _35653_);
  or g_46004_(_35628_, _35639_, _35654_);
  or g_46005_(_35653_, _35654_, _35655_);
  or g_46006_(_35632_, _35637_, _35656_);
  or g_46007_(_35640_, _35656_, _35657_);
  or g_46008_(_35655_, _35657_, _35658_);
  or g_46009_(_35651_, _35658_, _35659_);
  or g_46010_(_35644_, _35659_, _35660_);
  not g_46011_(_35660_, _35661_);
  xor g_46012_(out[225], out[577], _35662_);
  and g_46013_(out[235], _39900_, _35663_);
  xor g_46014_(out[233], out[585], _35664_);
  xor g_46015_(out[224], out[576], _35665_);
  xor g_46016_(out[238], out[590], _35666_);
  xor g_46017_(out[228], out[580], _35667_);
  or g_46018_(_35666_, _35667_, _35668_);
  xor g_46019_(out[237], out[589], _35669_);
  xor g_46020_(out[227], out[579], _35670_);
  and g_46021_(_39658_, out[587], _35671_);
  xor g_46022_(out[230], out[582], _35672_);
  xor g_46023_(out[234], out[586], _35673_);
  xor g_46024_(out[229], out[581], _35674_);
  xor g_46025_(out[239], out[591], _35675_);
  xor g_46026_(out[232], out[584], _35676_);
  or g_46027_(_35669_, _35676_, _35677_);
  xor g_46028_(out[226], out[578], _35678_);
  or g_46029_(_35673_, _35678_, _35679_);
  or g_46030_(_35677_, _35679_, _35680_);
  or g_46031_(_35664_, _35670_, _35681_);
  or g_46032_(_35674_, _35681_, _35682_);
  or g_46033_(_35680_, _35682_, _35683_);
  or g_46034_(_35668_, _35683_, _35684_);
  xor g_46035_(out[236], out[588], _35685_);
  or g_46036_(_35671_, _35685_, _35686_);
  xor g_46037_(out[231], out[583], _35687_);
  or g_46038_(_35672_, _35687_, _35688_);
  or g_46039_(_35686_, _35688_, _35689_);
  or g_46040_(_35662_, _35663_, _35690_);
  or g_46041_(_35675_, _35690_, _35691_);
  or g_46042_(_35689_, _35691_, _35692_);
  or g_46043_(_35665_, _35692_, _35693_);
  or g_46044_(_35684_, _35693_, _35694_);
  xor g_46045_(out[215], out[583], _35695_);
  and g_46046_(_39647_, out[587], _35696_);
  xor g_46047_(out[222], out[590], _35697_);
  xor g_46048_(out[216], out[584], _35698_);
  xor g_46049_(out[209], out[577], _35699_);
  xor g_46050_(out[221], out[589], _35700_);
  xor g_46051_(out[217], out[585], _35701_);
  xor g_46052_(out[212], out[580], _35702_);
  xor g_46053_(out[210], out[578], _35703_);
  and g_46054_(out[219], _39900_, _35704_);
  xor g_46055_(out[211], out[579], _35705_);
  xor g_46056_(out[214], out[582], _35706_);
  xor g_46057_(out[223], out[591], _35707_);
  xor g_46058_(out[218], out[586], _35708_);
  xor g_46059_(out[213], out[581], _35709_);
  xor g_46060_(out[208], out[576], _35710_);
  or g_46061_(_35697_, _35702_, _35711_);
  or g_46062_(_35698_, _35700_, _35712_);
  or g_46063_(_35703_, _35708_, _35713_);
  or g_46064_(_35712_, _35713_, _35714_);
  or g_46065_(_35701_, _35705_, _35715_);
  or g_46066_(_35709_, _35710_, _35716_);
  or g_46067_(_35715_, _35716_, _35717_);
  or g_46068_(_35714_, _35717_, _35718_);
  xor g_46069_(out[220], out[588], _35719_);
  or g_46070_(_35696_, _35719_, _35720_);
  or g_46071_(_35695_, _35706_, _35721_);
  or g_46072_(_35720_, _35721_, _35722_);
  or g_46073_(_35699_, _35704_, _35723_);
  or g_46074_(_35707_, _35723_, _35724_);
  or g_46075_(_35722_, _35724_, _35725_);
  or g_46076_(_35718_, _35725_, _35726_);
  or g_46077_(_35711_, _35726_, _35727_);
  xor g_46078_(out[202], out[586], _35728_);
  xor g_46079_(out[194], out[578], _35729_);
  xor g_46080_(out[193], out[577], _35730_);
  and g_46081_(_39636_, out[587], _35731_);
  and g_46082_(out[203], _39900_, _35732_);
  xor g_46083_(out[205], out[589], _35733_);
  xor g_46084_(out[195], out[579], _35734_);
  xor g_46085_(out[206], out[590], _35735_);
  xor g_46086_(out[204], out[588], _35736_);
  xor g_46087_(out[200], out[584], _35737_);
  xor g_46088_(out[207], out[591], _35738_);
  xor g_46089_(out[197], out[581], _35739_);
  xor g_46090_(out[198], out[582], _35740_);
  xor g_46091_(out[192], out[576], _35741_);
  xor g_46092_(out[196], out[580], _35742_);
  or g_46093_(_35733_, _35737_, _35743_);
  xor g_46094_(out[201], out[585], _35744_);
  or g_46095_(_35728_, _35729_, _35745_);
  or g_46096_(_35743_, _35745_, _35746_);
  or g_46097_(_35734_, _35744_, _35747_);
  or g_46098_(_35739_, _35747_, _35748_);
  or g_46099_(_35746_, _35748_, _35749_);
  or g_46100_(_35735_, _35742_, _35750_);
  or g_46101_(_35749_, _35750_, _35751_);
  or g_46102_(_35731_, _35736_, _35752_);
  xor g_46103_(out[199], out[583], _35753_);
  or g_46104_(_35740_, _35753_, _35754_);
  or g_46105_(_35752_, _35754_, _35755_);
  or g_46106_(_35730_, _35732_, _35756_);
  or g_46107_(_35738_, _35756_, _35757_);
  or g_46108_(_35755_, _35757_, _35758_);
  or g_46109_(_35741_, _35758_, _35759_);
  or g_46110_(_35751_, _35759_, _35760_);
  not g_46111_(_35760_, _35761_);
  xor g_46112_(out[183], out[583], _35762_);
  and g_46113_(_39625_, out[587], _35763_);
  xor g_46114_(out[190], out[590], _35764_);
  xor g_46115_(out[184], out[584], _35765_);
  xor g_46116_(out[177], out[577], _35766_);
  xor g_46117_(out[189], out[589], _35767_);
  xor g_46118_(out[185], out[585], _35768_);
  xor g_46119_(out[180], out[580], _35769_);
  xor g_46120_(out[178], out[578], _35770_);
  and g_46121_(out[187], _39900_, _35771_);
  xor g_46122_(out[179], out[579], _35772_);
  xor g_46123_(out[182], out[582], _35773_);
  xor g_46124_(out[191], out[591], _35774_);
  xor g_46125_(out[186], out[586], _35775_);
  xor g_46126_(out[181], out[581], _35776_);
  xor g_46127_(out[176], out[576], _35777_);
  or g_46128_(_35764_, _35769_, _35778_);
  or g_46129_(_35765_, _35767_, _35779_);
  or g_46130_(_35770_, _35775_, _35780_);
  or g_46131_(_35779_, _35780_, _35781_);
  or g_46132_(_35768_, _35772_, _35782_);
  or g_46133_(_35776_, _35777_, _35783_);
  or g_46134_(_35782_, _35783_, _35784_);
  or g_46135_(_35781_, _35784_, _35785_);
  xor g_46136_(out[188], out[588], _35786_);
  or g_46137_(_35763_, _35786_, _35787_);
  or g_46138_(_35762_, _35773_, _35788_);
  or g_46139_(_35787_, _35788_, _35789_);
  or g_46140_(_35766_, _35771_, _35790_);
  or g_46141_(_35774_, _35790_, _35791_);
  or g_46142_(_35789_, _35791_, _35792_);
  or g_46143_(_35785_, _35792_, _35793_);
  or g_46144_(_35778_, _35793_, _35794_);
  not g_46145_(_35794_, _35795_);
  xor g_46146_(out[161], out[577], _35796_);
  and g_46147_(out[171], _39900_, _35797_);
  xor g_46148_(out[169], out[585], _35798_);
  xor g_46149_(out[160], out[576], _35799_);
  xor g_46150_(out[174], out[590], _35800_);
  xor g_46151_(out[164], out[580], _35801_);
  or g_46152_(_35800_, _35801_, _35802_);
  xor g_46153_(out[173], out[589], _35803_);
  xor g_46154_(out[163], out[579], _35804_);
  and g_46155_(_39614_, out[587], _35805_);
  xor g_46156_(out[166], out[582], _35806_);
  xor g_46157_(out[170], out[586], _35807_);
  xor g_46158_(out[165], out[581], _35808_);
  xor g_46159_(out[175], out[591], _35809_);
  xor g_46160_(out[168], out[584], _35810_);
  or g_46161_(_35803_, _35810_, _35811_);
  xor g_46162_(out[162], out[578], _35812_);
  or g_46163_(_35807_, _35812_, _35813_);
  or g_46164_(_35811_, _35813_, _35814_);
  or g_46165_(_35798_, _35804_, _35815_);
  or g_46166_(_35808_, _35815_, _35816_);
  or g_46167_(_35814_, _35816_, _35817_);
  or g_46168_(_35802_, _35817_, _35818_);
  xor g_46169_(out[172], out[588], _35819_);
  or g_46170_(_35805_, _35819_, _35820_);
  xor g_46171_(out[167], out[583], _35821_);
  or g_46172_(_35806_, _35821_, _35822_);
  or g_46173_(_35820_, _35822_, _35823_);
  or g_46174_(_35796_, _35797_, _35824_);
  or g_46175_(_35809_, _35824_, _35825_);
  or g_46176_(_35823_, _35825_, _35826_);
  or g_46177_(_35799_, _35826_, _35827_);
  or g_46178_(_35818_, _35827_, _35828_);
  xor g_46179_(out[151], out[583], _35829_);
  and g_46180_(_39603_, out[587], _35830_);
  xor g_46181_(out[158], out[590], _35831_);
  xor g_46182_(out[152], out[584], _35832_);
  xor g_46183_(out[145], out[577], _35833_);
  xor g_46184_(out[157], out[589], _35834_);
  xor g_46185_(out[153], out[585], _35835_);
  xor g_46186_(out[148], out[580], _35836_);
  xor g_46187_(out[146], out[578], _35837_);
  and g_46188_(out[155], _39900_, _35838_);
  xor g_46189_(out[147], out[579], _35839_);
  xor g_46190_(out[150], out[582], _35840_);
  xor g_46191_(out[159], out[591], _35841_);
  xor g_46192_(out[154], out[586], _35842_);
  xor g_46193_(out[149], out[581], _35843_);
  xor g_46194_(out[144], out[576], _35844_);
  or g_46195_(_35831_, _35836_, _35845_);
  or g_46196_(_35832_, _35834_, _35846_);
  or g_46197_(_35837_, _35842_, _35847_);
  or g_46198_(_35846_, _35847_, _35848_);
  or g_46199_(_35835_, _35839_, _35849_);
  or g_46200_(_35843_, _35844_, _35850_);
  or g_46201_(_35849_, _35850_, _35851_);
  or g_46202_(_35848_, _35851_, _35852_);
  xor g_46203_(out[156], out[588], _35853_);
  or g_46204_(_35830_, _35853_, _35854_);
  or g_46205_(_35829_, _35840_, _35855_);
  or g_46206_(_35854_, _35855_, _35856_);
  or g_46207_(_35833_, _35838_, _35857_);
  or g_46208_(_35841_, _35857_, _35858_);
  or g_46209_(_35856_, _35858_, _35859_);
  or g_46210_(_35852_, _35859_, _35860_);
  or g_46211_(_35845_, _35860_, _35861_);
  not g_46212_(_35861_, _35862_);
  xor g_46213_(out[136], out[584], _35863_);
  xor g_46214_(out[133], out[581], _35864_);
  xor g_46215_(out[131], out[579], _35865_);
  xor g_46216_(out[142], out[590], _35866_);
  xor g_46217_(out[141], out[589], _35867_);
  xor g_46218_(out[130], out[578], _35868_);
  xor g_46219_(out[137], out[585], _35869_);
  xor g_46220_(out[134], out[582], _35870_);
  xor g_46221_(out[143], out[591], _35871_);
  xor g_46222_(out[138], out[586], _35872_);
  xor g_46223_(out[132], out[580], _35873_);
  xor g_46224_(out[128], out[576], _35874_);
  and g_46225_(_39592_, out[587], _35875_);
  and g_46226_(out[139], _39900_, _35876_);
  or g_46227_(_35863_, _35867_, _35877_);
  xor g_46228_(out[129], out[577], _35878_);
  or g_46229_(_35868_, _35872_, _35879_);
  or g_46230_(_35877_, _35879_, _35880_);
  or g_46231_(_35865_, _35869_, _35881_);
  or g_46232_(_35864_, _35881_, _35882_);
  or g_46233_(_35880_, _35882_, _35883_);
  or g_46234_(_35866_, _35873_, _35884_);
  or g_46235_(_35883_, _35884_, _35885_);
  xor g_46236_(out[140], out[588], _35886_);
  or g_46237_(_35875_, _35886_, _35887_);
  xor g_46238_(out[135], out[583], _35888_);
  or g_46239_(_35870_, _35888_, _35889_);
  or g_46240_(_35887_, _35889_, _35890_);
  or g_46241_(_35876_, _35878_, _35891_);
  or g_46242_(_35871_, _35891_, _35892_);
  or g_46243_(_35890_, _35892_, _35893_);
  or g_46244_(_35874_, _35893_, _35894_);
  or g_46245_(_35885_, _35894_, _35895_);
  xor g_46246_(out[119], out[583], _35896_);
  and g_46247_(_39581_, out[587], _35897_);
  xor g_46248_(out[126], out[590], _35898_);
  xor g_46249_(out[120], out[584], _35899_);
  xor g_46250_(out[113], out[577], _35900_);
  xor g_46251_(out[125], out[589], _35901_);
  xor g_46252_(out[121], out[585], _35902_);
  xor g_46253_(out[116], out[580], _35903_);
  xor g_46254_(out[114], out[578], _35904_);
  and g_46255_(out[123], _39900_, _35905_);
  xor g_46256_(out[115], out[579], _35906_);
  xor g_46257_(out[118], out[582], _35907_);
  xor g_46258_(out[127], out[591], _35908_);
  xor g_46259_(out[122], out[586], _35909_);
  xor g_46260_(out[117], out[581], _35910_);
  xor g_46261_(out[112], out[576], _35911_);
  or g_46262_(_35898_, _35903_, _35912_);
  or g_46263_(_35899_, _35901_, _35913_);
  or g_46264_(_35904_, _35909_, _35914_);
  or g_46265_(_35913_, _35914_, _35915_);
  or g_46266_(_35902_, _35906_, _35916_);
  or g_46267_(_35910_, _35911_, _35917_);
  or g_46268_(_35916_, _35917_, _35918_);
  or g_46269_(_35915_, _35918_, _35919_);
  xor g_46270_(out[124], out[588], _35920_);
  or g_46271_(_35897_, _35920_, _35921_);
  or g_46272_(_35896_, _35907_, _35922_);
  or g_46273_(_35921_, _35922_, _35923_);
  or g_46274_(_35900_, _35905_, _35924_);
  or g_46275_(_35908_, _35924_, _35925_);
  or g_46276_(_35923_, _35925_, _35926_);
  or g_46277_(_35919_, _35926_, _35927_);
  or g_46278_(_35912_, _35927_, _35928_);
  xor g_46279_(out[97], out[577], _35929_);
  and g_46280_(out[107], _39900_, _35930_);
  xor g_46281_(out[105], out[585], _35931_);
  xor g_46282_(out[96], out[576], _35932_);
  xor g_46283_(out[110], out[590], _35933_);
  xor g_46284_(out[100], out[580], _35934_);
  or g_46285_(_35933_, _35934_, _35935_);
  xor g_46286_(out[109], out[589], _35936_);
  xor g_46287_(out[99], out[579], _35937_);
  and g_46288_(_39570_, out[587], _35938_);
  xor g_46289_(out[102], out[582], _35939_);
  xor g_46290_(out[106], out[586], _35940_);
  xor g_46291_(out[101], out[581], _35941_);
  xor g_46292_(out[111], out[591], _35942_);
  xor g_46293_(out[104], out[584], _35943_);
  or g_46294_(_35936_, _35943_, _35944_);
  xor g_46295_(out[98], out[578], _35945_);
  or g_46296_(_35940_, _35945_, _35946_);
  or g_46297_(_35944_, _35946_, _35947_);
  or g_46298_(_35931_, _35937_, _35948_);
  or g_46299_(_35941_, _35948_, _35949_);
  or g_46300_(_35947_, _35949_, _35950_);
  or g_46301_(_35935_, _35950_, _35951_);
  xor g_46302_(out[108], out[588], _35952_);
  or g_46303_(_35938_, _35952_, _35953_);
  xor g_46304_(out[103], out[583], _35954_);
  or g_46305_(_35939_, _35954_, _35955_);
  or g_46306_(_35953_, _35955_, _35956_);
  or g_46307_(_35929_, _35930_, _35957_);
  or g_46308_(_35942_, _35957_, _35958_);
  or g_46309_(_35956_, _35958_, _35959_);
  or g_46310_(_35932_, _35959_, _35960_);
  or g_46311_(_35951_, _35960_, _35961_);
  xor g_46312_(out[87], out[583], _35962_);
  and g_46313_(_39559_, out[587], _35963_);
  xor g_46314_(out[94], out[590], _35964_);
  xor g_46315_(out[88], out[584], _35965_);
  xor g_46316_(out[81], out[577], _35966_);
  xor g_46317_(out[93], out[589], _35967_);
  xor g_46318_(out[89], out[585], _35968_);
  xor g_46319_(out[84], out[580], _35969_);
  xor g_46320_(out[82], out[578], _35970_);
  and g_46321_(out[91], _39900_, _35971_);
  xor g_46322_(out[83], out[579], _35972_);
  xor g_46323_(out[86], out[582], _35973_);
  xor g_46324_(out[95], out[591], _35974_);
  xor g_46325_(out[90], out[586], _35975_);
  xor g_46326_(out[85], out[581], _35976_);
  xor g_46327_(out[80], out[576], _35977_);
  or g_46328_(_35964_, _35969_, _35978_);
  or g_46329_(_35965_, _35967_, _35979_);
  or g_46330_(_35970_, _35975_, _35980_);
  or g_46331_(_35979_, _35980_, _35981_);
  or g_46332_(_35968_, _35972_, _35982_);
  or g_46333_(_35976_, _35977_, _35983_);
  or g_46334_(_35982_, _35983_, _35984_);
  or g_46335_(_35981_, _35984_, _35985_);
  xor g_46336_(out[92], out[588], _35986_);
  or g_46337_(_35963_, _35986_, _35987_);
  or g_46338_(_35962_, _35973_, _35988_);
  or g_46339_(_35987_, _35988_, _35989_);
  or g_46340_(_35966_, _35971_, _35990_);
  or g_46341_(_35974_, _35990_, _35991_);
  or g_46342_(_35989_, _35991_, _35992_);
  or g_46343_(_35985_, _35992_, _35993_);
  or g_46344_(_35978_, _35993_, _35994_);
  and g_46345_(out[75], _39900_, _35995_);
  and g_46346_(_39548_, out[587], _35996_);
  xor g_46347_(out[65], out[577], _35997_);
  xor g_46348_(out[67], out[579], _35998_);
  xor g_46349_(out[71], out[583], _35999_);
  xor g_46350_(out[73], out[585], _36000_);
  xor g_46351_(out[79], out[591], _36001_);
  xor g_46352_(out[66], out[578], _36002_);
  xor g_46353_(out[78], out[590], _36003_);
  xor g_46354_(out[77], out[589], _36004_);
  xor g_46355_(out[72], out[584], _36005_);
  or g_46356_(_36004_, _36005_, _36006_);
  xor g_46357_(out[68], out[580], _36007_);
  xor g_46358_(out[70], out[582], _36008_);
  xor g_46359_(out[74], out[586], _36009_);
  xor g_46360_(out[69], out[581], _36010_);
  xor g_46361_(out[64], out[576], _36011_);
  or g_46362_(_36002_, _36009_, _36012_);
  or g_46363_(_36006_, _36012_, _36013_);
  or g_46364_(_35998_, _36000_, _36014_);
  or g_46365_(_36010_, _36014_, _36015_);
  or g_46366_(_36013_, _36015_, _36016_);
  or g_46367_(_36003_, _36007_, _36017_);
  or g_46368_(_36016_, _36017_, _36018_);
  xor g_46369_(out[76], out[588], _36019_);
  or g_46370_(_35996_, _36019_, _36020_);
  or g_46371_(_35999_, _36008_, _36021_);
  or g_46372_(_36020_, _36021_, _36022_);
  or g_46373_(_35995_, _35997_, _36023_);
  or g_46374_(_36001_, _36023_, _36024_);
  or g_46375_(_36022_, _36024_, _36025_);
  or g_46376_(_36011_, _36025_, _36026_);
  or g_46377_(_36018_, _36026_, _36027_);
  xor g_46378_(out[55], out[583], _36028_);
  and g_46379_(_39537_, out[587], _36029_);
  xor g_46380_(out[62], out[590], _36030_);
  xor g_46381_(out[56], out[584], _36031_);
  xor g_46382_(out[49], out[577], _36032_);
  xor g_46383_(out[61], out[589], _36033_);
  xor g_46384_(out[57], out[585], _36034_);
  xor g_46385_(out[52], out[580], _36035_);
  xor g_46386_(out[50], out[578], _36036_);
  and g_46387_(out[59], _39900_, _36037_);
  xor g_46388_(out[51], out[579], _36038_);
  xor g_46389_(out[54], out[582], _36039_);
  xor g_46390_(out[63], out[591], _36040_);
  xor g_46391_(out[58], out[586], _36041_);
  xor g_46392_(out[53], out[581], _36042_);
  xor g_46393_(out[48], out[576], _36043_);
  or g_46394_(_36030_, _36035_, _36044_);
  or g_46395_(_36031_, _36033_, _36045_);
  or g_46396_(_36036_, _36041_, _36046_);
  or g_46397_(_36045_, _36046_, _36047_);
  or g_46398_(_36034_, _36038_, _36048_);
  or g_46399_(_36042_, _36043_, _36049_);
  or g_46400_(_36048_, _36049_, _36050_);
  or g_46401_(_36047_, _36050_, _36051_);
  xor g_46402_(out[60], out[588], _36052_);
  or g_46403_(_36029_, _36052_, _36053_);
  or g_46404_(_36028_, _36039_, _36054_);
  or g_46405_(_36053_, _36054_, _36055_);
  or g_46406_(_36032_, _36037_, _36056_);
  or g_46407_(_36040_, _36056_, _36057_);
  or g_46408_(_36055_, _36057_, _36058_);
  or g_46409_(_36051_, _36058_, _36059_);
  or g_46410_(_36044_, _36059_, _36060_);
  xor g_46411_(out[33], out[577], _36061_);
  and g_46412_(_39526_, out[587], _36062_);
  and g_46413_(out[43], _39900_, _36063_);
  xor g_46414_(out[46], out[590], _36064_);
  xor g_46415_(out[35], out[579], _36065_);
  xor g_46416_(out[36], out[580], _36066_);
  xor g_46417_(out[34], out[578], _36067_);
  xor g_46418_(out[41], out[585], _36068_);
  xor g_46419_(out[32], out[576], _36069_);
  xor g_46420_(out[44], out[588], _36070_);
  xor g_46421_(out[38], out[582], _36071_);
  xor g_46422_(out[42], out[586], _36072_);
  xor g_46423_(out[37], out[581], _36073_);
  xor g_46424_(out[47], out[591], _36074_);
  xor g_46425_(out[45], out[589], _36075_);
  xor g_46426_(out[40], out[584], _36076_);
  or g_46427_(_36064_, _36066_, _36077_);
  or g_46428_(_36075_, _36076_, _36078_);
  or g_46429_(_36067_, _36072_, _36079_);
  or g_46430_(_36078_, _36079_, _36080_);
  or g_46431_(_36065_, _36068_, _36081_);
  or g_46432_(_36069_, _36073_, _36082_);
  or g_46433_(_36081_, _36082_, _36083_);
  or g_46434_(_36080_, _36083_, _36084_);
  or g_46435_(_36062_, _36070_, _36085_);
  xor g_46436_(out[39], out[583], _36086_);
  or g_46437_(_36071_, _36086_, _36087_);
  or g_46438_(_36085_, _36087_, _36088_);
  or g_46439_(_36061_, _36063_, _36089_);
  or g_46440_(_36074_, _36089_, _36090_);
  or g_46441_(_36088_, _36090_, _36091_);
  or g_46442_(_36084_, _36091_, _36092_);
  or g_46443_(_36077_, _36092_, _36093_);
  not g_46444_(_36093_, _36094_);
  xor g_46445_(out[23], out[583], _36095_);
  and g_46446_(_39493_, out[587], _36096_);
  xor g_46447_(out[30], out[590], _36097_);
  xor g_46448_(out[24], out[584], _36098_);
  xor g_46449_(out[17], out[577], _36099_);
  xor g_46450_(out[29], out[589], _36100_);
  xor g_46451_(out[25], out[585], _36101_);
  xor g_46452_(out[20], out[580], _36102_);
  xor g_46453_(out[18], out[578], _36103_);
  and g_46454_(out[27], _39900_, _36104_);
  xor g_46455_(out[19], out[579], _36105_);
  xor g_46456_(out[22], out[582], _36106_);
  xor g_46457_(out[31], out[591], _36107_);
  xor g_46458_(out[26], out[586], _36108_);
  xor g_46459_(out[21], out[581], _36109_);
  xor g_46460_(out[16], out[576], _36110_);
  or g_46461_(_36097_, _36102_, _36111_);
  or g_46462_(_36098_, _36100_, _36112_);
  or g_46463_(_36103_, _36108_, _36113_);
  or g_46464_(_36112_, _36113_, _36114_);
  or g_46465_(_36101_, _36105_, _36115_);
  or g_46466_(_36109_, _36110_, _36116_);
  or g_46467_(_36115_, _36116_, _36117_);
  or g_46468_(_36114_, _36117_, _36118_);
  xor g_46469_(out[28], out[588], _36119_);
  or g_46470_(_36096_, _36119_, _36120_);
  or g_46471_(_36095_, _36106_, _36121_);
  or g_46472_(_36120_, _36121_, _36122_);
  or g_46473_(_36099_, _36104_, _36123_);
  or g_46474_(_36107_, _36123_, _36124_);
  or g_46475_(_36122_, _36124_, _36125_);
  or g_46476_(_36118_, _36125_, _36126_);
  or g_46477_(_36111_, _36126_, _36127_);
  xor g_46478_(out[4], out[580], _36128_);
  xor g_46479_(out[12], out[588], _36129_);
  and g_46480_(_39438_, out[587], _36130_);
  xor g_46481_(out[10], out[586], _36131_);
  xor g_46482_(out[6], out[582], _36132_);
  xor g_46483_(out[5], out[581], _36133_);
  xor g_46484_(out[3], out[579], _36134_);
  xor g_46485_(out[13], out[589], _36135_);
  xor g_46486_(out[14], out[590], _36136_);
  xor g_46487_(out[1], out[577], _36137_);
  xor g_46488_(out[2], out[578], _36138_);
  and g_46489_(out[11], _39900_, _36139_);
  xor g_46490_(out[0], out[576], _36140_);
  xor g_46491_(out[15], out[591], _36141_);
  xor g_46492_(out[8], out[584], _36142_);
  or g_46493_(_36135_, _36142_, _36143_);
  xor g_46494_(out[9], out[585], _36144_);
  or g_46495_(_36131_, _36138_, _36145_);
  or g_46496_(_36143_, _36145_, _36146_);
  or g_46497_(_36134_, _36144_, _36147_);
  or g_46498_(_36133_, _36147_, _36148_);
  or g_46499_(_36146_, _36148_, _36149_);
  or g_46500_(_36128_, _36136_, _36150_);
  or g_46501_(_36149_, _36150_, _36151_);
  or g_46502_(_36129_, _36130_, _36152_);
  xor g_46503_(out[7], out[583], _36153_);
  or g_46504_(_36132_, _36153_, _36154_);
  or g_46505_(_36152_, _36154_, _36155_);
  or g_46506_(_36137_, _36139_, _36156_);
  or g_46507_(_36141_, _36156_, _36157_);
  or g_46508_(_36155_, _36157_, _36158_);
  or g_46509_(_36140_, _36158_, _36159_);
  or g_46510_(_36151_, _36159_, _36160_);
  not g_46511_(_36160_, _36161_);
  xor g_46512_(out[314], out[570], _36162_);
  xor g_46513_(out[306], out[562], _36163_);
  xor g_46514_(out[305], out[561], _36164_);
  and g_46515_(_39724_, out[571], _36165_);
  and g_46516_(out[315], _39889_, _36166_);
  xor g_46517_(out[317], out[573], _36167_);
  xor g_46518_(out[307], out[563], _36168_);
  xor g_46519_(out[318], out[574], _36169_);
  xor g_46520_(out[316], out[572], _36170_);
  xor g_46521_(out[312], out[568], _36171_);
  xor g_46522_(out[319], out[575], _36172_);
  xor g_46523_(out[309], out[565], _36173_);
  xor g_46524_(out[310], out[566], _36174_);
  xor g_46525_(out[304], out[560], _36175_);
  xor g_46526_(out[308], out[564], _36176_);
  or g_46527_(_36167_, _36171_, _36177_);
  xor g_46528_(out[313], out[569], _36178_);
  or g_46529_(_36162_, _36163_, _36179_);
  or g_46530_(_36177_, _36179_, _36180_);
  or g_46531_(_36168_, _36178_, _36181_);
  or g_46532_(_36173_, _36181_, _36182_);
  or g_46533_(_36180_, _36182_, _36183_);
  or g_46534_(_36169_, _36176_, _36184_);
  or g_46535_(_36183_, _36184_, _36185_);
  or g_46536_(_36165_, _36170_, _36186_);
  xor g_46537_(out[311], out[567], _36187_);
  or g_46538_(_36174_, _36187_, _36188_);
  or g_46539_(_36186_, _36188_, _36189_);
  or g_46540_(_36164_, _36166_, _36190_);
  or g_46541_(_36172_, _36190_, _36191_);
  or g_46542_(_36189_, _36191_, _36192_);
  or g_46543_(_36175_, _36192_, _36193_);
  or g_46544_(_36185_, _36193_, _36194_);
  not g_46545_(_36194_, _36195_);
  xor g_46546_(out[295], out[567], _36196_);
  and g_46547_(_39702_, out[571], _36197_);
  xor g_46548_(out[302], out[574], _36198_);
  xor g_46549_(out[296], out[568], _36199_);
  xor g_46550_(out[289], out[561], _36200_);
  xor g_46551_(out[301], out[573], _36201_);
  xor g_46552_(out[297], out[569], _36202_);
  xor g_46553_(out[292], out[564], _36203_);
  xor g_46554_(out[290], out[562], _36204_);
  and g_46555_(out[299], _39889_, _36205_);
  xor g_46556_(out[291], out[563], _36206_);
  xor g_46557_(out[294], out[566], _36207_);
  xor g_46558_(out[303], out[575], _36208_);
  xor g_46559_(out[298], out[570], _36209_);
  xor g_46560_(out[293], out[565], _36210_);
  xor g_46561_(out[288], out[560], _36211_);
  or g_46562_(_36198_, _36203_, _36212_);
  or g_46563_(_36199_, _36201_, _36213_);
  or g_46564_(_36204_, _36209_, _36214_);
  or g_46565_(_36213_, _36214_, _36215_);
  or g_46566_(_36202_, _36206_, _36216_);
  or g_46567_(_36210_, _36211_, _36217_);
  or g_46568_(_36216_, _36217_, _36218_);
  or g_46569_(_36215_, _36218_, _36219_);
  xor g_46570_(out[300], out[572], _36220_);
  or g_46571_(_36197_, _36220_, _36221_);
  or g_46572_(_36196_, _36207_, _36222_);
  or g_46573_(_36221_, _36222_, _36223_);
  or g_46574_(_36200_, _36205_, _36224_);
  or g_46575_(_36208_, _36224_, _36225_);
  or g_46576_(_36223_, _36225_, _36226_);
  or g_46577_(_36219_, _36226_, _36227_);
  or g_46578_(_36212_, _36227_, _36228_);
  xor g_46579_(out[273], out[561], _36229_);
  and g_46580_(out[283], _39889_, _36230_);
  xor g_46581_(out[286], out[574], _36231_);
  xor g_46582_(out[275], out[563], _36232_);
  xor g_46583_(out[276], out[564], _36233_);
  xor g_46584_(out[274], out[562], _36234_);
  xor g_46585_(out[281], out[569], _36235_);
  xor g_46586_(out[272], out[560], _36236_);
  and g_46587_(_39691_, out[571], _36237_);
  xor g_46588_(out[278], out[566], _36238_);
  xor g_46589_(out[282], out[570], _36239_);
  xor g_46590_(out[277], out[565], _36240_);
  xor g_46591_(out[287], out[575], _36241_);
  xor g_46592_(out[285], out[573], _36242_);
  xor g_46593_(out[280], out[568], _36243_);
  or g_46594_(_36231_, _36233_, _36244_);
  or g_46595_(_36242_, _36243_, _36245_);
  or g_46596_(_36234_, _36239_, _36246_);
  or g_46597_(_36245_, _36246_, _36247_);
  or g_46598_(_36232_, _36235_, _36248_);
  or g_46599_(_36236_, _36240_, _36249_);
  or g_46600_(_36248_, _36249_, _36250_);
  or g_46601_(_36247_, _36250_, _36251_);
  xor g_46602_(out[284], out[572], _36252_);
  or g_46603_(_36237_, _36252_, _36253_);
  xor g_46604_(out[279], out[567], _36254_);
  or g_46605_(_36238_, _36254_, _36255_);
  or g_46606_(_36253_, _36255_, _36256_);
  or g_46607_(_36229_, _36230_, _36257_);
  or g_46608_(_36241_, _36257_, _36258_);
  or g_46609_(_36256_, _36258_, _36259_);
  or g_46610_(_36251_, _36259_, _36260_);
  or g_46611_(_36244_, _36260_, _36261_);
  xor g_46612_(out[263], out[567], _36262_);
  and g_46613_(_39680_, out[571], _36263_);
  xor g_46614_(out[270], out[574], _36264_);
  xor g_46615_(out[264], out[568], _36265_);
  xor g_46616_(out[257], out[561], _36266_);
  xor g_46617_(out[269], out[573], _36267_);
  xor g_46618_(out[265], out[569], _36268_);
  xor g_46619_(out[260], out[564], _36269_);
  xor g_46620_(out[258], out[562], _36270_);
  and g_46621_(out[267], _39889_, _36271_);
  xor g_46622_(out[259], out[563], _36272_);
  xor g_46623_(out[262], out[566], _36273_);
  xor g_46624_(out[271], out[575], _36274_);
  xor g_46625_(out[266], out[570], _36275_);
  xor g_46626_(out[261], out[565], _36276_);
  xor g_46627_(out[256], out[560], _36277_);
  or g_46628_(_36264_, _36269_, _36278_);
  or g_46629_(_36265_, _36267_, _36279_);
  or g_46630_(_36270_, _36275_, _36280_);
  or g_46631_(_36279_, _36280_, _36281_);
  or g_46632_(_36268_, _36272_, _36282_);
  or g_46633_(_36276_, _36277_, _36283_);
  or g_46634_(_36282_, _36283_, _36284_);
  or g_46635_(_36281_, _36284_, _36285_);
  xor g_46636_(out[268], out[572], _36286_);
  or g_46637_(_36263_, _36286_, _36287_);
  or g_46638_(_36262_, _36273_, _36288_);
  or g_46639_(_36287_, _36288_, _36289_);
  or g_46640_(_36266_, _36271_, _36290_);
  or g_46641_(_36274_, _36290_, _36291_);
  or g_46642_(_36289_, _36291_, _36292_);
  or g_46643_(_36285_, _36292_, _36293_);
  or g_46644_(_36278_, _36293_, _36294_);
  not g_46645_(_36294_, _36295_);
  xor g_46646_(out[241], out[561], _36296_);
  and g_46647_(out[251], _39889_, _36297_);
  xor g_46648_(out[249], out[569], _36298_);
  xor g_46649_(out[240], out[560], _36299_);
  xor g_46650_(out[254], out[574], _36300_);
  xor g_46651_(out[244], out[564], _36301_);
  or g_46652_(_36300_, _36301_, _36302_);
  xor g_46653_(out[253], out[573], _36303_);
  xor g_46654_(out[243], out[563], _36304_);
  and g_46655_(_39669_, out[571], _36305_);
  xor g_46656_(out[246], out[566], _36306_);
  xor g_46657_(out[250], out[570], _36307_);
  xor g_46658_(out[245], out[565], _36308_);
  xor g_46659_(out[255], out[575], _36309_);
  xor g_46660_(out[248], out[568], _36310_);
  or g_46661_(_36303_, _36310_, _36311_);
  xor g_46662_(out[242], out[562], _36312_);
  or g_46663_(_36307_, _36312_, _36313_);
  or g_46664_(_36311_, _36313_, _36314_);
  or g_46665_(_36298_, _36304_, _36315_);
  or g_46666_(_36308_, _36315_, _36316_);
  or g_46667_(_36314_, _36316_, _36317_);
  or g_46668_(_36302_, _36317_, _36318_);
  xor g_46669_(out[252], out[572], _36319_);
  or g_46670_(_36305_, _36319_, _36320_);
  xor g_46671_(out[247], out[567], _36321_);
  or g_46672_(_36306_, _36321_, _36322_);
  or g_46673_(_36320_, _36322_, _36323_);
  or g_46674_(_36296_, _36297_, _36324_);
  or g_46675_(_36309_, _36324_, _36325_);
  or g_46676_(_36323_, _36325_, _36326_);
  or g_46677_(_36299_, _36326_, _36327_);
  or g_46678_(_36318_, _36327_, _36328_);
  not g_46679_(_36328_, _36329_);
  xor g_46680_(out[231], out[567], _36330_);
  and g_46681_(_39658_, out[571], _36331_);
  xor g_46682_(out[238], out[574], _36332_);
  xor g_46683_(out[232], out[568], _36333_);
  xor g_46684_(out[225], out[561], _36334_);
  xor g_46685_(out[237], out[573], _36335_);
  xor g_46686_(out[233], out[569], _36336_);
  xor g_46687_(out[228], out[564], _36337_);
  xor g_46688_(out[226], out[562], _36338_);
  and g_46689_(out[235], _39889_, _36339_);
  xor g_46690_(out[227], out[563], _36340_);
  xor g_46691_(out[230], out[566], _36341_);
  xor g_46692_(out[239], out[575], _36342_);
  xor g_46693_(out[234], out[570], _36343_);
  xor g_46694_(out[229], out[565], _36344_);
  xor g_46695_(out[224], out[560], _36345_);
  or g_46696_(_36332_, _36337_, _36346_);
  or g_46697_(_36333_, _36335_, _36347_);
  or g_46698_(_36338_, _36343_, _36348_);
  or g_46699_(_36347_, _36348_, _36349_);
  or g_46700_(_36336_, _36340_, _36350_);
  or g_46701_(_36344_, _36345_, _36351_);
  or g_46702_(_36350_, _36351_, _36352_);
  or g_46703_(_36349_, _36352_, _36353_);
  xor g_46704_(out[236], out[572], _36354_);
  or g_46705_(_36331_, _36354_, _36355_);
  or g_46706_(_36330_, _36341_, _36356_);
  or g_46707_(_36355_, _36356_, _36357_);
  or g_46708_(_36334_, _36339_, _36358_);
  or g_46709_(_36342_, _36358_, _36359_);
  or g_46710_(_36357_, _36359_, _36360_);
  or g_46711_(_36353_, _36360_, _36361_);
  or g_46712_(_36346_, _36361_, _36362_);
  xor g_46713_(out[209], out[561], _36363_);
  and g_46714_(out[219], _39889_, _36364_);
  xor g_46715_(out[217], out[569], _36365_);
  xor g_46716_(out[208], out[560], _36366_);
  xor g_46717_(out[222], out[574], _36367_);
  xor g_46718_(out[212], out[564], _36368_);
  or g_46719_(_36367_, _36368_, _36369_);
  xor g_46720_(out[221], out[573], _36370_);
  xor g_46721_(out[211], out[563], _36371_);
  and g_46722_(_39647_, out[571], _36372_);
  xor g_46723_(out[214], out[566], _36373_);
  xor g_46724_(out[218], out[570], _36374_);
  xor g_46725_(out[213], out[565], _36375_);
  xor g_46726_(out[223], out[575], _36376_);
  xor g_46727_(out[216], out[568], _36377_);
  or g_46728_(_36370_, _36377_, _36378_);
  xor g_46729_(out[210], out[562], _36379_);
  or g_46730_(_36374_, _36379_, _36380_);
  or g_46731_(_36378_, _36380_, _36381_);
  or g_46732_(_36365_, _36371_, _36382_);
  or g_46733_(_36375_, _36382_, _36383_);
  or g_46734_(_36381_, _36383_, _36384_);
  or g_46735_(_36369_, _36384_, _36385_);
  xor g_46736_(out[220], out[572], _36386_);
  or g_46737_(_36372_, _36386_, _36387_);
  xor g_46738_(out[215], out[567], _36388_);
  or g_46739_(_36373_, _36388_, _36389_);
  or g_46740_(_36387_, _36389_, _36390_);
  or g_46741_(_36363_, _36364_, _36391_);
  or g_46742_(_36376_, _36391_, _36392_);
  or g_46743_(_36390_, _36392_, _36393_);
  or g_46744_(_36366_, _36393_, _36394_);
  or g_46745_(_36385_, _36394_, _36395_);
  xor g_46746_(out[199], out[567], _36396_);
  and g_46747_(_39636_, out[571], _36397_);
  xor g_46748_(out[206], out[574], _36398_);
  xor g_46749_(out[200], out[568], _36399_);
  xor g_46750_(out[193], out[561], _36400_);
  xor g_46751_(out[205], out[573], _36401_);
  xor g_46752_(out[201], out[569], _36402_);
  xor g_46753_(out[196], out[564], _36403_);
  xor g_46754_(out[194], out[562], _36404_);
  and g_46755_(out[203], _39889_, _36405_);
  xor g_46756_(out[195], out[563], _36406_);
  xor g_46757_(out[198], out[566], _36407_);
  xor g_46758_(out[207], out[575], _36408_);
  xor g_46759_(out[202], out[570], _36409_);
  xor g_46760_(out[197], out[565], _36410_);
  xor g_46761_(out[192], out[560], _36411_);
  or g_46762_(_36398_, _36403_, _36412_);
  or g_46763_(_36399_, _36401_, _36413_);
  or g_46764_(_36404_, _36409_, _36414_);
  or g_46765_(_36413_, _36414_, _36415_);
  or g_46766_(_36402_, _36406_, _36416_);
  or g_46767_(_36410_, _36411_, _36417_);
  or g_46768_(_36416_, _36417_, _36418_);
  or g_46769_(_36415_, _36418_, _36419_);
  xor g_46770_(out[204], out[572], _36420_);
  or g_46771_(_36397_, _36420_, _36421_);
  or g_46772_(_36396_, _36407_, _36422_);
  or g_46773_(_36421_, _36422_, _36423_);
  or g_46774_(_36400_, _36405_, _36424_);
  or g_46775_(_36408_, _36424_, _36425_);
  or g_46776_(_36423_, _36425_, _36426_);
  or g_46777_(_36419_, _36426_, _36427_);
  or g_46778_(_36412_, _36427_, _36428_);
  not g_46779_(_36428_, _36429_);
  xor g_46780_(out[177], out[561], _36430_);
  and g_46781_(out[187], _39889_, _36431_);
  xor g_46782_(out[185], out[569], _36432_);
  xor g_46783_(out[176], out[560], _36433_);
  xor g_46784_(out[190], out[574], _36434_);
  xor g_46785_(out[180], out[564], _36435_);
  or g_46786_(_36434_, _36435_, _36436_);
  xor g_46787_(out[189], out[573], _36437_);
  xor g_46788_(out[179], out[563], _36438_);
  and g_46789_(_39625_, out[571], _36439_);
  xor g_46790_(out[182], out[566], _36440_);
  xor g_46791_(out[186], out[570], _36441_);
  xor g_46792_(out[181], out[565], _36442_);
  xor g_46793_(out[191], out[575], _36443_);
  xor g_46794_(out[184], out[568], _36444_);
  or g_46795_(_36437_, _36444_, _36445_);
  xor g_46796_(out[178], out[562], _36446_);
  or g_46797_(_36441_, _36446_, _36447_);
  or g_46798_(_36445_, _36447_, _36448_);
  or g_46799_(_36432_, _36438_, _36449_);
  or g_46800_(_36442_, _36449_, _36450_);
  or g_46801_(_36448_, _36450_, _36451_);
  or g_46802_(_36436_, _36451_, _36452_);
  xor g_46803_(out[188], out[572], _36453_);
  or g_46804_(_36439_, _36453_, _36454_);
  xor g_46805_(out[183], out[567], _36455_);
  or g_46806_(_36440_, _36455_, _36456_);
  or g_46807_(_36454_, _36456_, _36457_);
  or g_46808_(_36430_, _36431_, _36458_);
  or g_46809_(_36443_, _36458_, _36459_);
  or g_46810_(_36457_, _36459_, _36460_);
  or g_46811_(_36433_, _36460_, _36461_);
  or g_46812_(_36452_, _36461_, _36462_);
  xor g_46813_(out[167], out[567], _36463_);
  and g_46814_(_39614_, out[571], _36464_);
  xor g_46815_(out[174], out[574], _36465_);
  xor g_46816_(out[168], out[568], _36466_);
  xor g_46817_(out[161], out[561], _36467_);
  xor g_46818_(out[173], out[573], _36468_);
  xor g_46819_(out[169], out[569], _36469_);
  xor g_46820_(out[164], out[564], _36470_);
  xor g_46821_(out[162], out[562], _36471_);
  and g_46822_(out[171], _39889_, _36472_);
  xor g_46823_(out[163], out[563], _36473_);
  xor g_46824_(out[166], out[566], _36474_);
  xor g_46825_(out[175], out[575], _36475_);
  xor g_46826_(out[170], out[570], _36476_);
  xor g_46827_(out[165], out[565], _36477_);
  xor g_46828_(out[160], out[560], _36478_);
  or g_46829_(_36465_, _36470_, _36479_);
  or g_46830_(_36466_, _36468_, _36480_);
  or g_46831_(_36471_, _36476_, _36481_);
  or g_46832_(_36480_, _36481_, _36482_);
  or g_46833_(_36469_, _36473_, _36483_);
  or g_46834_(_36477_, _36478_, _36484_);
  or g_46835_(_36483_, _36484_, _36485_);
  or g_46836_(_36482_, _36485_, _36486_);
  xor g_46837_(out[172], out[572], _36487_);
  or g_46838_(_36464_, _36487_, _36488_);
  or g_46839_(_36463_, _36474_, _36489_);
  or g_46840_(_36488_, _36489_, _36490_);
  or g_46841_(_36467_, _36472_, _36491_);
  or g_46842_(_36475_, _36491_, _36492_);
  or g_46843_(_36490_, _36492_, _36493_);
  or g_46844_(_36486_, _36493_, _36494_);
  or g_46845_(_36479_, _36494_, _36495_);
  xor g_46846_(out[148], out[564], _36496_);
  xor g_46847_(out[156], out[572], _36497_);
  and g_46848_(_39603_, out[571], _36498_);
  xor g_46849_(out[154], out[570], _36499_);
  xor g_46850_(out[150], out[566], _36500_);
  xor g_46851_(out[149], out[565], _36501_);
  xor g_46852_(out[147], out[563], _36502_);
  xor g_46853_(out[157], out[573], _36503_);
  xor g_46854_(out[158], out[574], _36504_);
  xor g_46855_(out[145], out[561], _36505_);
  xor g_46856_(out[146], out[562], _36506_);
  and g_46857_(out[155], _39889_, _36507_);
  xor g_46858_(out[144], out[560], _36508_);
  xor g_46859_(out[159], out[575], _36509_);
  xor g_46860_(out[152], out[568], _36510_);
  or g_46861_(_36503_, _36510_, _36511_);
  xor g_46862_(out[153], out[569], _36512_);
  or g_46863_(_36499_, _36506_, _36513_);
  or g_46864_(_36511_, _36513_, _36514_);
  or g_46865_(_36502_, _36512_, _36515_);
  or g_46866_(_36501_, _36515_, _36516_);
  or g_46867_(_36514_, _36516_, _36517_);
  or g_46868_(_36496_, _36504_, _36518_);
  or g_46869_(_36517_, _36518_, _36519_);
  or g_46870_(_36497_, _36498_, _36520_);
  xor g_46871_(out[151], out[567], _36521_);
  or g_46872_(_36500_, _36521_, _36522_);
  or g_46873_(_36520_, _36522_, _36523_);
  or g_46874_(_36505_, _36507_, _36524_);
  or g_46875_(_36509_, _36524_, _36525_);
  or g_46876_(_36523_, _36525_, _36526_);
  or g_46877_(_36508_, _36526_, _36527_);
  or g_46878_(_36519_, _36527_, _36528_);
  xor g_46879_(out[135], out[567], _36529_);
  and g_46880_(_39592_, out[571], _36530_);
  xor g_46881_(out[142], out[574], _36531_);
  xor g_46882_(out[136], out[568], _36532_);
  xor g_46883_(out[129], out[561], _36533_);
  xor g_46884_(out[141], out[573], _36534_);
  xor g_46885_(out[137], out[569], _36535_);
  xor g_46886_(out[132], out[564], _36536_);
  xor g_46887_(out[130], out[562], _36537_);
  and g_46888_(out[139], _39889_, _36538_);
  xor g_46889_(out[131], out[563], _36539_);
  xor g_46890_(out[134], out[566], _36540_);
  xor g_46891_(out[143], out[575], _36541_);
  xor g_46892_(out[138], out[570], _36542_);
  xor g_46893_(out[133], out[565], _36543_);
  xor g_46894_(out[128], out[560], _36544_);
  or g_46895_(_36531_, _36536_, _36545_);
  or g_46896_(_36532_, _36534_, _36546_);
  or g_46897_(_36537_, _36542_, _36547_);
  or g_46898_(_36546_, _36547_, _36548_);
  or g_46899_(_36535_, _36539_, _36549_);
  or g_46900_(_36543_, _36544_, _36550_);
  or g_46901_(_36549_, _36550_, _36551_);
  or g_46902_(_36548_, _36551_, _36552_);
  xor g_46903_(out[140], out[572], _36553_);
  or g_46904_(_36530_, _36553_, _36554_);
  or g_46905_(_36529_, _36540_, _36555_);
  or g_46906_(_36554_, _36555_, _36556_);
  or g_46907_(_36533_, _36538_, _36557_);
  or g_46908_(_36541_, _36557_, _36558_);
  or g_46909_(_36556_, _36558_, _36559_);
  or g_46910_(_36552_, _36559_, _36560_);
  or g_46911_(_36545_, _36560_, _36561_);
  xor g_46912_(out[115], out[563], _36562_);
  xor g_46913_(out[116], out[564], _36563_);
  xor g_46914_(out[126], out[574], _36564_);
  xor g_46915_(out[114], out[562], _36565_);
  xor g_46916_(out[117], out[565], _36566_);
  xor g_46917_(out[121], out[569], _36567_);
  xor g_46918_(out[120], out[568], _36568_);
  xor g_46919_(out[127], out[575], _36569_);
  xor g_46920_(out[122], out[570], _36570_);
  xor g_46921_(out[118], out[566], _36571_);
  xor g_46922_(out[112], out[560], _36572_);
  and g_46923_(_39581_, out[571], _36573_);
  and g_46924_(out[123], _39889_, _36574_);
  xor g_46925_(out[125], out[573], _36575_);
  or g_46926_(_36568_, _36575_, _36576_);
  xor g_46927_(out[113], out[561], _36577_);
  or g_46928_(_36565_, _36570_, _36578_);
  or g_46929_(_36576_, _36578_, _36579_);
  or g_46930_(_36562_, _36567_, _36580_);
  or g_46931_(_36566_, _36580_, _36581_);
  or g_46932_(_36579_, _36581_, _36582_);
  or g_46933_(_36563_, _36564_, _36583_);
  or g_46934_(_36582_, _36583_, _36584_);
  xor g_46935_(out[124], out[572], _36585_);
  or g_46936_(_36573_, _36585_, _36586_);
  xor g_46937_(out[119], out[567], _36587_);
  or g_46938_(_36571_, _36587_, _36588_);
  or g_46939_(_36586_, _36588_, _36589_);
  or g_46940_(_36574_, _36577_, _36590_);
  or g_46941_(_36569_, _36590_, _36591_);
  or g_46942_(_36589_, _36591_, _36592_);
  or g_46943_(_36572_, _36592_, _36593_);
  or g_46944_(_36584_, _36593_, _36594_);
  xor g_46945_(out[103], out[567], _36595_);
  and g_46946_(_39570_, out[571], _36596_);
  xor g_46947_(out[110], out[574], _36597_);
  xor g_46948_(out[104], out[568], _36598_);
  xor g_46949_(out[97], out[561], _36599_);
  xor g_46950_(out[109], out[573], _36600_);
  xor g_46951_(out[105], out[569], _36601_);
  xor g_46952_(out[100], out[564], _36602_);
  xor g_46953_(out[98], out[562], _36603_);
  and g_46954_(out[107], _39889_, _36604_);
  xor g_46955_(out[99], out[563], _36605_);
  xor g_46956_(out[102], out[566], _36606_);
  xor g_46957_(out[111], out[575], _36607_);
  xor g_46958_(out[106], out[570], _36608_);
  xor g_46959_(out[101], out[565], _36609_);
  xor g_46960_(out[96], out[560], _36610_);
  or g_46961_(_36597_, _36602_, _36611_);
  or g_46962_(_36598_, _36600_, _36612_);
  or g_46963_(_36603_, _36608_, _36613_);
  or g_46964_(_36612_, _36613_, _36614_);
  or g_46965_(_36601_, _36605_, _36615_);
  or g_46966_(_36609_, _36610_, _36616_);
  or g_46967_(_36615_, _36616_, _36617_);
  or g_46968_(_36614_, _36617_, _36618_);
  xor g_46969_(out[108], out[572], _36619_);
  or g_46970_(_36596_, _36619_, _36620_);
  or g_46971_(_36595_, _36606_, _36621_);
  or g_46972_(_36620_, _36621_, _36622_);
  or g_46973_(_36599_, _36604_, _36623_);
  or g_46974_(_36607_, _36623_, _36624_);
  or g_46975_(_36622_, _36624_, _36625_);
  or g_46976_(_36618_, _36625_, _36626_);
  or g_46977_(_36611_, _36626_, _36627_);
  xor g_46978_(out[90], out[570], _36628_);
  xor g_46979_(out[82], out[562], _36629_);
  xor g_46980_(out[81], out[561], _36630_);
  and g_46981_(_39559_, out[571], _36631_);
  and g_46982_(out[91], _39889_, _36632_);
  xor g_46983_(out[93], out[573], _36633_);
  xor g_46984_(out[83], out[563], _36634_);
  xor g_46985_(out[94], out[574], _36635_);
  xor g_46986_(out[92], out[572], _36636_);
  xor g_46987_(out[88], out[568], _36637_);
  xor g_46988_(out[95], out[575], _36638_);
  xor g_46989_(out[85], out[565], _36639_);
  xor g_46990_(out[86], out[566], _36640_);
  xor g_46991_(out[80], out[560], _36641_);
  xor g_46992_(out[84], out[564], _36642_);
  or g_46993_(_36633_, _36637_, _36643_);
  xor g_46994_(out[89], out[569], _36644_);
  or g_46995_(_36628_, _36629_, _36645_);
  or g_46996_(_36643_, _36645_, _36646_);
  or g_46997_(_36634_, _36644_, _36647_);
  or g_46998_(_36639_, _36647_, _36648_);
  or g_46999_(_36646_, _36648_, _36649_);
  or g_47000_(_36635_, _36642_, _36650_);
  or g_47001_(_36649_, _36650_, _36651_);
  or g_47002_(_36631_, _36636_, _36652_);
  xor g_47003_(out[87], out[567], _36653_);
  or g_47004_(_36640_, _36653_, _36654_);
  or g_47005_(_36652_, _36654_, _36655_);
  or g_47006_(_36630_, _36632_, _36656_);
  or g_47007_(_36638_, _36656_, _36657_);
  or g_47008_(_36655_, _36657_, _36658_);
  or g_47009_(_36641_, _36658_, _36659_);
  or g_47010_(_36651_, _36659_, _36660_);
  xor g_47011_(out[71], out[567], _36661_);
  and g_47012_(_39548_, out[571], _36662_);
  xor g_47013_(out[78], out[574], _36663_);
  xor g_47014_(out[72], out[568], _36664_);
  xor g_47015_(out[65], out[561], _36665_);
  xor g_47016_(out[77], out[573], _36666_);
  xor g_47017_(out[73], out[569], _36667_);
  xor g_47018_(out[68], out[564], _36668_);
  xor g_47019_(out[66], out[562], _36669_);
  and g_47020_(out[75], _39889_, _36670_);
  xor g_47021_(out[67], out[563], _36671_);
  xor g_47022_(out[70], out[566], _36672_);
  xor g_47023_(out[79], out[575], _36673_);
  xor g_47024_(out[74], out[570], _36674_);
  xor g_47025_(out[69], out[565], _36675_);
  xor g_47026_(out[64], out[560], _36676_);
  or g_47027_(_36663_, _36668_, _36677_);
  or g_47028_(_36664_, _36666_, _36678_);
  or g_47029_(_36669_, _36674_, _36679_);
  or g_47030_(_36678_, _36679_, _36680_);
  or g_47031_(_36667_, _36671_, _36681_);
  or g_47032_(_36675_, _36676_, _36682_);
  or g_47033_(_36681_, _36682_, _36683_);
  or g_47034_(_36680_, _36683_, _36684_);
  xor g_47035_(out[76], out[572], _36685_);
  or g_47036_(_36662_, _36685_, _36686_);
  or g_47037_(_36661_, _36672_, _36687_);
  or g_47038_(_36686_, _36687_, _36688_);
  or g_47039_(_36665_, _36670_, _36689_);
  or g_47040_(_36673_, _36689_, _36690_);
  or g_47041_(_36688_, _36690_, _36691_);
  or g_47042_(_36684_, _36691_, _36692_);
  or g_47043_(_36677_, _36692_, _36693_);
  xor g_47044_(out[49], out[561], _36694_);
  and g_47045_(_39537_, out[571], _36695_);
  and g_47046_(out[59], _39889_, _36696_);
  xor g_47047_(out[56], out[568], _36697_);
  xor g_47048_(out[58], out[570], _36698_);
  xor g_47049_(out[50], out[562], _36699_);
  xor g_47050_(out[52], out[564], _36700_);
  xor g_47051_(out[61], out[573], _36701_);
  xor g_47052_(out[57], out[569], _36702_);
  xor g_47053_(out[51], out[563], _36703_);
  xor g_47054_(out[53], out[565], _36704_);
  xor g_47055_(out[62], out[574], _36705_);
  xor g_47056_(out[48], out[560], _36706_);
  xor g_47057_(out[63], out[575], _36707_);
  or g_47058_(_36697_, _36701_, _36708_);
  xor g_47059_(out[54], out[566], _36709_);
  or g_47060_(_36698_, _36699_, _36710_);
  or g_47061_(_36708_, _36710_, _36711_);
  or g_47062_(_36702_, _36703_, _36712_);
  or g_47063_(_36704_, _36712_, _36713_);
  or g_47064_(_36711_, _36713_, _36714_);
  or g_47065_(_36700_, _36705_, _36715_);
  or g_47066_(_36714_, _36715_, _36716_);
  xor g_47067_(out[60], out[572], _36717_);
  or g_47068_(_36695_, _36717_, _36718_);
  xor g_47069_(out[55], out[567], _36719_);
  or g_47070_(_36709_, _36719_, _36720_);
  or g_47071_(_36718_, _36720_, _36721_);
  or g_47072_(_36694_, _36696_, _36722_);
  or g_47073_(_36707_, _36722_, _36723_);
  or g_47074_(_36721_, _36723_, _36724_);
  or g_47075_(_36706_, _36724_, _36725_);
  or g_47076_(_36716_, _36725_, _36726_);
  xor g_47077_(out[39], out[567], _36727_);
  and g_47078_(_39526_, out[571], _36728_);
  xor g_47079_(out[46], out[574], _36729_);
  xor g_47080_(out[40], out[568], _36730_);
  xor g_47081_(out[33], out[561], _36731_);
  xor g_47082_(out[45], out[573], _36732_);
  xor g_47083_(out[41], out[569], _36733_);
  xor g_47084_(out[36], out[564], _36734_);
  xor g_47085_(out[34], out[562], _36735_);
  and g_47086_(out[43], _39889_, _36736_);
  xor g_47087_(out[35], out[563], _36737_);
  xor g_47088_(out[38], out[566], _36738_);
  xor g_47089_(out[47], out[575], _36739_);
  xor g_47090_(out[42], out[570], _36740_);
  xor g_47091_(out[37], out[565], _36741_);
  xor g_47092_(out[32], out[560], _36742_);
  or g_47093_(_36729_, _36734_, _36743_);
  or g_47094_(_36730_, _36732_, _36744_);
  or g_47095_(_36735_, _36740_, _36745_);
  or g_47096_(_36744_, _36745_, _36746_);
  or g_47097_(_36733_, _36737_, _36747_);
  or g_47098_(_36741_, _36742_, _36748_);
  or g_47099_(_36747_, _36748_, _36749_);
  or g_47100_(_36746_, _36749_, _36750_);
  xor g_47101_(out[44], out[572], _36751_);
  or g_47102_(_36728_, _36751_, _36752_);
  or g_47103_(_36727_, _36738_, _36753_);
  or g_47104_(_36752_, _36753_, _36754_);
  or g_47105_(_36731_, _36736_, _36755_);
  or g_47106_(_36739_, _36755_, _36756_);
  or g_47107_(_36754_, _36756_, _36757_);
  or g_47108_(_36750_, _36757_, _36758_);
  or g_47109_(_36743_, _36758_, _36759_);
  xor g_47110_(out[17], out[561], _36760_);
  and g_47111_(out[27], _39889_, _36761_);
  xor g_47112_(out[30], out[574], _36762_);
  xor g_47113_(out[19], out[563], _36763_);
  xor g_47114_(out[20], out[564], _36764_);
  xor g_47115_(out[18], out[562], _36765_);
  xor g_47116_(out[25], out[569], _36766_);
  xor g_47117_(out[16], out[560], _36767_);
  and g_47118_(_39493_, out[571], _36768_);
  xor g_47119_(out[22], out[566], _36769_);
  xor g_47120_(out[26], out[570], _36770_);
  xor g_47121_(out[21], out[565], _36771_);
  xor g_47122_(out[31], out[575], _36772_);
  xor g_47123_(out[29], out[573], _36773_);
  xor g_47124_(out[24], out[568], _36774_);
  or g_47125_(_36762_, _36764_, _36775_);
  or g_47126_(_36773_, _36774_, _36776_);
  or g_47127_(_36765_, _36770_, _36777_);
  or g_47128_(_36776_, _36777_, _36778_);
  or g_47129_(_36763_, _36766_, _36779_);
  or g_47130_(_36767_, _36771_, _36780_);
  or g_47131_(_36779_, _36780_, _36781_);
  or g_47132_(_36778_, _36781_, _36782_);
  xor g_47133_(out[28], out[572], _36783_);
  or g_47134_(_36768_, _36783_, _36784_);
  xor g_47135_(out[23], out[567], _36785_);
  or g_47136_(_36769_, _36785_, _36786_);
  or g_47137_(_36784_, _36786_, _36787_);
  or g_47138_(_36760_, _36761_, _36788_);
  or g_47139_(_36772_, _36788_, _36789_);
  or g_47140_(_36787_, _36789_, _36790_);
  or g_47141_(_36782_, _36790_, _36791_);
  or g_47142_(_36775_, _36791_, _36792_);
  xor g_47143_(out[1], out[561], _36793_);
  and g_47144_(_39438_, out[571], _36794_);
  and g_47145_(out[11], _39889_, _36795_);
  xor g_47146_(out[8], out[568], _36796_);
  xor g_47147_(out[10], out[570], _36797_);
  xor g_47148_(out[2], out[562], _36798_);
  xor g_47149_(out[4], out[564], _36799_);
  xor g_47150_(out[5], out[565], _36800_);
  xor g_47151_(out[9], out[569], _36801_);
  xor g_47152_(out[3], out[563], _36802_);
  xor g_47153_(out[14], out[574], _36803_);
  xor g_47154_(out[0], out[560], _36804_);
  xor g_47155_(out[15], out[575], _36805_);
  xor g_47156_(out[13], out[573], _36806_);
  or g_47157_(_36796_, _36806_, _36807_);
  xor g_47158_(out[6], out[566], _36808_);
  or g_47159_(_36797_, _36798_, _36809_);
  or g_47160_(_36807_, _36809_, _36810_);
  or g_47161_(_36801_, _36802_, _36811_);
  or g_47162_(_36800_, _36811_, _36812_);
  or g_47163_(_36810_, _36812_, _36813_);
  or g_47164_(_36799_, _36803_, _36814_);
  or g_47165_(_36813_, _36814_, _36815_);
  xor g_47166_(out[12], out[572], _36816_);
  or g_47167_(_36794_, _36816_, _36817_);
  xor g_47168_(out[7], out[567], _36818_);
  or g_47169_(_36808_, _36818_, _36819_);
  or g_47170_(_36817_, _36819_, _36820_);
  or g_47171_(_36793_, _36795_, _36821_);
  or g_47172_(_36805_, _36821_, _36822_);
  or g_47173_(_36820_, _36822_, _36823_);
  or g_47174_(_36804_, _36823_, _36824_);
  or g_47175_(_36815_, _36824_, _36825_);
  xor g_47176_(out[311], out[551], _36826_);
  and g_47177_(_39724_, out[555], _36827_);
  xor g_47178_(out[318], out[558], _36828_);
  xor g_47179_(out[312], out[552], _36829_);
  xor g_47180_(out[305], out[545], _36830_);
  xor g_47181_(out[317], out[557], _36831_);
  xor g_47182_(out[313], out[553], _36832_);
  xor g_47183_(out[308], out[548], _36833_);
  xor g_47184_(out[306], out[546], _36834_);
  and g_47185_(out[315], _39878_, _36835_);
  xor g_47186_(out[307], out[547], _36836_);
  xor g_47187_(out[310], out[550], _36837_);
  xor g_47188_(out[319], out[559], _36838_);
  xor g_47189_(out[314], out[554], _36839_);
  xor g_47190_(out[309], out[549], _36840_);
  xor g_47191_(out[304], out[544], _36841_);
  or g_47192_(_36828_, _36833_, _36842_);
  or g_47193_(_36829_, _36831_, _36843_);
  or g_47194_(_36834_, _36839_, _36844_);
  or g_47195_(_36843_, _36844_, _36845_);
  or g_47196_(_36832_, _36836_, _36846_);
  or g_47197_(_36840_, _36841_, _36847_);
  or g_47198_(_36846_, _36847_, _36848_);
  or g_47199_(_36845_, _36848_, _36849_);
  xor g_47200_(out[316], out[556], _36850_);
  or g_47201_(_36827_, _36850_, _36851_);
  or g_47202_(_36826_, _36837_, _36852_);
  or g_47203_(_36851_, _36852_, _36853_);
  or g_47204_(_36830_, _36835_, _36854_);
  or g_47205_(_36838_, _36854_, _36855_);
  or g_47206_(_36853_, _36855_, _36856_);
  or g_47207_(_36849_, _36856_, _36857_);
  or g_47208_(_36842_, _36857_, _36858_);
  xor g_47209_(out[298], out[554], _36859_);
  xor g_47210_(out[290], out[546], _36860_);
  xor g_47211_(out[289], out[545], _36861_);
  and g_47212_(_39702_, out[555], _36862_);
  and g_47213_(out[299], _39878_, _36863_);
  xor g_47214_(out[301], out[557], _36864_);
  xor g_47215_(out[291], out[547], _36865_);
  xor g_47216_(out[302], out[558], _36866_);
  xor g_47217_(out[300], out[556], _36867_);
  xor g_47218_(out[296], out[552], _36868_);
  xor g_47219_(out[303], out[559], _36869_);
  xor g_47220_(out[293], out[549], _36870_);
  xor g_47221_(out[294], out[550], _36871_);
  xor g_47222_(out[288], out[544], _36872_);
  xor g_47223_(out[292], out[548], _36873_);
  or g_47224_(_36864_, _36868_, _36874_);
  xor g_47225_(out[297], out[553], _36875_);
  or g_47226_(_36859_, _36860_, _36876_);
  or g_47227_(_36874_, _36876_, _36877_);
  or g_47228_(_36865_, _36875_, _36878_);
  or g_47229_(_36870_, _36878_, _36879_);
  or g_47230_(_36877_, _36879_, _36880_);
  or g_47231_(_36866_, _36873_, _36881_);
  or g_47232_(_36880_, _36881_, _36882_);
  or g_47233_(_36862_, _36867_, _36883_);
  xor g_47234_(out[295], out[551], _36884_);
  or g_47235_(_36871_, _36884_, _36885_);
  or g_47236_(_36883_, _36885_, _36886_);
  or g_47237_(_36861_, _36863_, _36887_);
  or g_47238_(_36869_, _36887_, _36888_);
  or g_47239_(_36886_, _36888_, _36889_);
  or g_47240_(_36872_, _36889_, _36890_);
  or g_47241_(_36882_, _36890_, _36891_);
  xor g_47242_(out[279], out[551], _36892_);
  and g_47243_(_39691_, out[555], _36893_);
  xor g_47244_(out[286], out[558], _36894_);
  xor g_47245_(out[280], out[552], _36895_);
  xor g_47246_(out[273], out[545], _36896_);
  xor g_47247_(out[285], out[557], _36897_);
  xor g_47248_(out[281], out[553], _36898_);
  xor g_47249_(out[276], out[548], _36899_);
  xor g_47250_(out[274], out[546], _36900_);
  and g_47251_(out[283], _39878_, _36901_);
  xor g_47252_(out[275], out[547], _36902_);
  xor g_47253_(out[278], out[550], _36903_);
  xor g_47254_(out[287], out[559], _36904_);
  xor g_47255_(out[282], out[554], _36905_);
  xor g_47256_(out[277], out[549], _36906_);
  xor g_47257_(out[272], out[544], _36907_);
  or g_47258_(_36894_, _36899_, _36908_);
  or g_47259_(_36895_, _36897_, _36909_);
  or g_47260_(_36900_, _36905_, _36910_);
  or g_47261_(_36909_, _36910_, _36911_);
  or g_47262_(_36898_, _36902_, _36912_);
  or g_47263_(_36906_, _36907_, _36913_);
  or g_47264_(_36912_, _36913_, _36914_);
  or g_47265_(_36911_, _36914_, _36915_);
  xor g_47266_(out[284], out[556], _36916_);
  or g_47267_(_36893_, _36916_, _36917_);
  or g_47268_(_36892_, _36903_, _36918_);
  or g_47269_(_36917_, _36918_, _36919_);
  or g_47270_(_36896_, _36901_, _36920_);
  or g_47271_(_36904_, _36920_, _36921_);
  or g_47272_(_36919_, _36921_, _36922_);
  or g_47273_(_36915_, _36922_, _36923_);
  or g_47274_(_36908_, _36923_, _36924_);
  not g_47275_(_36924_, _36925_);
  and g_47276_(out[267], _39878_, _36926_);
  xor g_47277_(out[260], out[548], _36927_);
  xor g_47278_(out[270], out[558], _36928_);
  or g_47279_(_36927_, _36928_, _36929_);
  xor g_47280_(out[269], out[557], _36930_);
  xor g_47281_(out[259], out[547], _36931_);
  xor g_47282_(out[256], out[544], _36932_);
  and g_47283_(_39680_, out[555], _36933_);
  xor g_47284_(out[266], out[554], _36934_);
  xor g_47285_(out[271], out[559], _36935_);
  xor g_47286_(out[262], out[550], _36936_);
  xor g_47287_(out[261], out[549], _36937_);
  xor g_47288_(out[264], out[552], _36938_);
  or g_47289_(_36930_, _36938_, _36939_);
  xor g_47290_(out[258], out[546], _36940_);
  xor g_47291_(out[265], out[553], _36941_);
  xor g_47292_(out[257], out[545], _36942_);
  or g_47293_(_36934_, _36940_, _36943_);
  or g_47294_(_36939_, _36943_, _36944_);
  or g_47295_(_36931_, _36941_, _36945_);
  or g_47296_(_36937_, _36945_, _36946_);
  or g_47297_(_36944_, _36946_, _36947_);
  or g_47298_(_36929_, _36947_, _36948_);
  xor g_47299_(out[268], out[556], _36949_);
  or g_47300_(_36933_, _36949_, _36950_);
  xor g_47301_(out[263], out[551], _36951_);
  or g_47302_(_36936_, _36951_, _36952_);
  or g_47303_(_36950_, _36952_, _36953_);
  or g_47304_(_36926_, _36942_, _36954_);
  or g_47305_(_36935_, _36954_, _36955_);
  or g_47306_(_36953_, _36955_, _36956_);
  or g_47307_(_36932_, _36956_, _36957_);
  or g_47308_(_36948_, _36957_, _36958_);
  xor g_47309_(out[247], out[551], _36959_);
  and g_47310_(_39669_, out[555], _36960_);
  xor g_47311_(out[254], out[558], _36961_);
  xor g_47312_(out[248], out[552], _36962_);
  xor g_47313_(out[241], out[545], _36963_);
  xor g_47314_(out[253], out[557], _36964_);
  xor g_47315_(out[249], out[553], _36965_);
  xor g_47316_(out[244], out[548], _36966_);
  xor g_47317_(out[242], out[546], _36967_);
  and g_47318_(out[251], _39878_, _36968_);
  xor g_47319_(out[243], out[547], _36969_);
  xor g_47320_(out[246], out[550], _36970_);
  xor g_47321_(out[255], out[559], _36971_);
  xor g_47322_(out[250], out[554], _36972_);
  xor g_47323_(out[245], out[549], _36973_);
  xor g_47324_(out[240], out[544], _36974_);
  or g_47325_(_36961_, _36966_, _36975_);
  or g_47326_(_36962_, _36964_, _36976_);
  or g_47327_(_36967_, _36972_, _36977_);
  or g_47328_(_36976_, _36977_, _36978_);
  or g_47329_(_36965_, _36969_, _36979_);
  or g_47330_(_36973_, _36974_, _36980_);
  or g_47331_(_36979_, _36980_, _36981_);
  or g_47332_(_36978_, _36981_, _36982_);
  xor g_47333_(out[252], out[556], _36983_);
  or g_47334_(_36960_, _36983_, _36984_);
  or g_47335_(_36959_, _36970_, _36985_);
  or g_47336_(_36984_, _36985_, _36986_);
  or g_47337_(_36963_, _36968_, _36987_);
  or g_47338_(_36971_, _36987_, _36988_);
  or g_47339_(_36986_, _36988_, _36989_);
  or g_47340_(_36982_, _36989_, _36990_);
  or g_47341_(_36975_, _36990_, _36991_);
  xor g_47342_(out[225], out[545], _36992_);
  and g_47343_(out[235], _39878_, _36993_);
  xor g_47344_(out[233], out[553], _36994_);
  xor g_47345_(out[224], out[544], _36995_);
  xor g_47346_(out[238], out[558], _36996_);
  xor g_47347_(out[228], out[548], _36997_);
  or g_47348_(_36996_, _36997_, _36998_);
  xor g_47349_(out[237], out[557], _36999_);
  xor g_47350_(out[227], out[547], _37000_);
  and g_47351_(_39658_, out[555], _37001_);
  xor g_47352_(out[230], out[550], _37002_);
  xor g_47353_(out[234], out[554], _37003_);
  xor g_47354_(out[229], out[549], _37004_);
  xor g_47355_(out[239], out[559], _37005_);
  xor g_47356_(out[232], out[552], _37006_);
  or g_47357_(_36999_, _37006_, _37007_);
  xor g_47358_(out[226], out[546], _37008_);
  or g_47359_(_37003_, _37008_, _37009_);
  or g_47360_(_37007_, _37009_, _37010_);
  or g_47361_(_36994_, _37000_, _37011_);
  or g_47362_(_37004_, _37011_, _37012_);
  or g_47363_(_37010_, _37012_, _37013_);
  or g_47364_(_36998_, _37013_, _37014_);
  xor g_47365_(out[236], out[556], _37015_);
  or g_47366_(_37001_, _37015_, _37016_);
  xor g_47367_(out[231], out[551], _37017_);
  or g_47368_(_37002_, _37017_, _37018_);
  or g_47369_(_37016_, _37018_, _37019_);
  or g_47370_(_36992_, _36993_, _37020_);
  or g_47371_(_37005_, _37020_, _37021_);
  or g_47372_(_37019_, _37021_, _37022_);
  or g_47373_(_36995_, _37022_, _37023_);
  or g_47374_(_37014_, _37023_, _37024_);
  xor g_47375_(out[215], out[551], _37025_);
  and g_47376_(_39647_, out[555], _37026_);
  xor g_47377_(out[222], out[558], _37027_);
  xor g_47378_(out[216], out[552], _37028_);
  xor g_47379_(out[209], out[545], _37029_);
  xor g_47380_(out[221], out[557], _37030_);
  xor g_47381_(out[217], out[553], _37031_);
  xor g_47382_(out[212], out[548], _37032_);
  xor g_47383_(out[210], out[546], _37033_);
  and g_47384_(out[219], _39878_, _37034_);
  xor g_47385_(out[211], out[547], _37035_);
  xor g_47386_(out[214], out[550], _37036_);
  xor g_47387_(out[223], out[559], _37037_);
  xor g_47388_(out[218], out[554], _37038_);
  xor g_47389_(out[213], out[549], _37039_);
  xor g_47390_(out[208], out[544], _37040_);
  or g_47391_(_37027_, _37032_, _37041_);
  or g_47392_(_37028_, _37030_, _37042_);
  or g_47393_(_37033_, _37038_, _37043_);
  or g_47394_(_37042_, _37043_, _37044_);
  or g_47395_(_37031_, _37035_, _37045_);
  or g_47396_(_37039_, _37040_, _37046_);
  or g_47397_(_37045_, _37046_, _37047_);
  or g_47398_(_37044_, _37047_, _37048_);
  xor g_47399_(out[220], out[556], _37049_);
  or g_47400_(_37026_, _37049_, _37050_);
  or g_47401_(_37025_, _37036_, _37051_);
  or g_47402_(_37050_, _37051_, _37052_);
  or g_47403_(_37029_, _37034_, _37053_);
  or g_47404_(_37037_, _37053_, _37054_);
  or g_47405_(_37052_, _37054_, _37055_);
  or g_47406_(_37048_, _37055_, _37056_);
  or g_47407_(_37041_, _37056_, _37057_);
  not g_47408_(_37057_, _37058_);
  xor g_47409_(out[193], out[545], _37059_);
  and g_47410_(_39636_, out[555], _37060_);
  and g_47411_(out[203], _39878_, _37061_);
  xor g_47412_(out[206], out[558], _37062_);
  xor g_47413_(out[195], out[547], _37063_);
  xor g_47414_(out[196], out[548], _37064_);
  xor g_47415_(out[194], out[546], _37065_);
  xor g_47416_(out[201], out[553], _37066_);
  xor g_47417_(out[192], out[544], _37067_);
  xor g_47418_(out[204], out[556], _37068_);
  xor g_47419_(out[198], out[550], _37069_);
  xor g_47420_(out[202], out[554], _37070_);
  xor g_47421_(out[197], out[549], _37071_);
  xor g_47422_(out[207], out[559], _37072_);
  xor g_47423_(out[205], out[557], _37073_);
  xor g_47424_(out[200], out[552], _37074_);
  or g_47425_(_37062_, _37064_, _37075_);
  or g_47426_(_37073_, _37074_, _37076_);
  or g_47427_(_37065_, _37070_, _37077_);
  or g_47428_(_37076_, _37077_, _37078_);
  or g_47429_(_37063_, _37066_, _37079_);
  or g_47430_(_37067_, _37071_, _37080_);
  or g_47431_(_37079_, _37080_, _37081_);
  or g_47432_(_37078_, _37081_, _37082_);
  or g_47433_(_37060_, _37068_, _37083_);
  xor g_47434_(out[199], out[551], _37084_);
  or g_47435_(_37069_, _37084_, _37085_);
  or g_47436_(_37083_, _37085_, _37086_);
  or g_47437_(_37059_, _37061_, _37087_);
  or g_47438_(_37072_, _37087_, _37088_);
  or g_47439_(_37086_, _37088_, _37089_);
  or g_47440_(_37082_, _37089_, _37090_);
  or g_47441_(_37075_, _37090_, _37091_);
  not g_47442_(_37091_, _37092_);
  xor g_47443_(out[183], out[551], _37093_);
  and g_47444_(_39625_, out[555], _37094_);
  xor g_47445_(out[190], out[558], _37095_);
  xor g_47446_(out[184], out[552], _37096_);
  xor g_47447_(out[177], out[545], _37097_);
  xor g_47448_(out[189], out[557], _37098_);
  xor g_47449_(out[185], out[553], _37099_);
  xor g_47450_(out[180], out[548], _37100_);
  xor g_47451_(out[178], out[546], _37101_);
  and g_47452_(out[187], _39878_, _37102_);
  xor g_47453_(out[179], out[547], _37103_);
  xor g_47454_(out[182], out[550], _37104_);
  xor g_47455_(out[191], out[559], _37105_);
  xor g_47456_(out[186], out[554], _37106_);
  xor g_47457_(out[181], out[549], _37107_);
  xor g_47458_(out[176], out[544], _37108_);
  or g_47459_(_37095_, _37100_, _37109_);
  or g_47460_(_37096_, _37098_, _37110_);
  or g_47461_(_37101_, _37106_, _37111_);
  or g_47462_(_37110_, _37111_, _37112_);
  or g_47463_(_37099_, _37103_, _37113_);
  or g_47464_(_37107_, _37108_, _37114_);
  or g_47465_(_37113_, _37114_, _37115_);
  or g_47466_(_37112_, _37115_, _37116_);
  xor g_47467_(out[188], out[556], _37117_);
  or g_47468_(_37094_, _37117_, _37118_);
  or g_47469_(_37093_, _37104_, _37119_);
  or g_47470_(_37118_, _37119_, _37120_);
  or g_47471_(_37097_, _37102_, _37121_);
  or g_47472_(_37105_, _37121_, _37122_);
  or g_47473_(_37120_, _37122_, _37123_);
  or g_47474_(_37116_, _37123_, _37124_);
  or g_47475_(_37109_, _37124_, _37125_);
  not g_47476_(_37125_, _37126_);
  xor g_47477_(out[161], out[545], _37127_);
  and g_47478_(out[171], _39878_, _37128_);
  xor g_47479_(out[169], out[553], _37129_);
  xor g_47480_(out[160], out[544], _37130_);
  xor g_47481_(out[174], out[558], _37131_);
  xor g_47482_(out[164], out[548], _37132_);
  or g_47483_(_37131_, _37132_, _37133_);
  xor g_47484_(out[173], out[557], _37134_);
  xor g_47485_(out[163], out[547], _37135_);
  and g_47486_(_39614_, out[555], _37136_);
  xor g_47487_(out[166], out[550], _37137_);
  xor g_47488_(out[170], out[554], _37138_);
  xor g_47489_(out[165], out[549], _37139_);
  xor g_47490_(out[175], out[559], _37140_);
  xor g_47491_(out[168], out[552], _37141_);
  or g_47492_(_37134_, _37141_, _37142_);
  xor g_47493_(out[162], out[546], _37143_);
  or g_47494_(_37138_, _37143_, _37144_);
  or g_47495_(_37142_, _37144_, _37145_);
  or g_47496_(_37129_, _37135_, _37146_);
  or g_47497_(_37139_, _37146_, _37147_);
  or g_47498_(_37145_, _37147_, _37148_);
  or g_47499_(_37133_, _37148_, _37149_);
  xor g_47500_(out[172], out[556], _37150_);
  or g_47501_(_37136_, _37150_, _37151_);
  xor g_47502_(out[167], out[551], _37152_);
  or g_47503_(_37137_, _37152_, _37153_);
  or g_47504_(_37151_, _37153_, _37154_);
  or g_47505_(_37127_, _37128_, _37155_);
  or g_47506_(_37140_, _37155_, _37156_);
  or g_47507_(_37154_, _37156_, _37157_);
  or g_47508_(_37130_, _37157_, _37158_);
  or g_47509_(_37149_, _37158_, _37159_);
  xor g_47510_(out[151], out[551], _37160_);
  and g_47511_(_39603_, out[555], _37161_);
  xor g_47512_(out[158], out[558], _37162_);
  xor g_47513_(out[152], out[552], _37163_);
  xor g_47514_(out[145], out[545], _37164_);
  xor g_47515_(out[157], out[557], _37165_);
  xor g_47516_(out[153], out[553], _37166_);
  xor g_47517_(out[148], out[548], _37167_);
  xor g_47518_(out[146], out[546], _37168_);
  and g_47519_(out[155], _39878_, _37169_);
  xor g_47520_(out[147], out[547], _37170_);
  xor g_47521_(out[150], out[550], _37171_);
  xor g_47522_(out[159], out[559], _37172_);
  xor g_47523_(out[154], out[554], _37173_);
  xor g_47524_(out[149], out[549], _37174_);
  xor g_47525_(out[144], out[544], _37175_);
  or g_47526_(_37162_, _37167_, _37176_);
  or g_47527_(_37163_, _37165_, _37177_);
  or g_47528_(_37168_, _37173_, _37178_);
  or g_47529_(_37177_, _37178_, _37179_);
  or g_47530_(_37166_, _37170_, _37180_);
  or g_47531_(_37174_, _37175_, _37181_);
  or g_47532_(_37180_, _37181_, _37182_);
  or g_47533_(_37179_, _37182_, _37183_);
  xor g_47534_(out[156], out[556], _37184_);
  or g_47535_(_37161_, _37184_, _37185_);
  or g_47536_(_37160_, _37171_, _37186_);
  or g_47537_(_37185_, _37186_, _37187_);
  or g_47538_(_37164_, _37169_, _37188_);
  or g_47539_(_37172_, _37188_, _37189_);
  or g_47540_(_37187_, _37189_, _37190_);
  or g_47541_(_37183_, _37190_, _37191_);
  or g_47542_(_37176_, _37191_, _37192_);
  xor g_47543_(out[129], out[545], _37193_);
  and g_47544_(_39592_, out[555], _37194_);
  and g_47545_(out[139], _39878_, _37195_);
  xor g_47546_(out[136], out[552], _37196_);
  xor g_47547_(out[138], out[554], _37197_);
  xor g_47548_(out[130], out[546], _37198_);
  xor g_47549_(out[132], out[548], _37199_);
  xor g_47550_(out[133], out[549], _37200_);
  xor g_47551_(out[137], out[553], _37201_);
  xor g_47552_(out[131], out[547], _37202_);
  xor g_47553_(out[142], out[558], _37203_);
  xor g_47554_(out[128], out[544], _37204_);
  xor g_47555_(out[143], out[559], _37205_);
  xor g_47556_(out[141], out[557], _37206_);
  or g_47557_(_37196_, _37206_, _37207_);
  xor g_47558_(out[134], out[550], _37208_);
  or g_47559_(_37197_, _37198_, _37209_);
  or g_47560_(_37207_, _37209_, _37210_);
  or g_47561_(_37201_, _37202_, _37211_);
  or g_47562_(_37200_, _37211_, _37212_);
  or g_47563_(_37210_, _37212_, _37213_);
  or g_47564_(_37199_, _37203_, _37214_);
  or g_47565_(_37213_, _37214_, _37215_);
  xor g_47566_(out[140], out[556], _37216_);
  or g_47567_(_37194_, _37216_, _37217_);
  xor g_47568_(out[135], out[551], _37218_);
  or g_47569_(_37208_, _37218_, _37219_);
  or g_47570_(_37217_, _37219_, _37220_);
  or g_47571_(_37193_, _37195_, _37221_);
  or g_47572_(_37205_, _37221_, _37222_);
  or g_47573_(_37220_, _37222_, _37223_);
  or g_47574_(_37204_, _37223_, _37224_);
  or g_47575_(_37215_, _37224_, _37225_);
  not g_47576_(_37225_, _37226_);
  xor g_47577_(out[119], out[551], _37227_);
  and g_47578_(_39581_, out[555], _37228_);
  xor g_47579_(out[126], out[558], _37229_);
  xor g_47580_(out[120], out[552], _37230_);
  xor g_47581_(out[113], out[545], _37231_);
  xor g_47582_(out[125], out[557], _37232_);
  xor g_47583_(out[121], out[553], _37233_);
  xor g_47584_(out[116], out[548], _37234_);
  xor g_47585_(out[114], out[546], _37235_);
  and g_47586_(out[123], _39878_, _37236_);
  xor g_47587_(out[115], out[547], _37237_);
  xor g_47588_(out[118], out[550], _37238_);
  xor g_47589_(out[127], out[559], _37239_);
  xor g_47590_(out[122], out[554], _37240_);
  xor g_47591_(out[117], out[549], _37241_);
  xor g_47592_(out[112], out[544], _37242_);
  or g_47593_(_37229_, _37234_, _37243_);
  or g_47594_(_37230_, _37232_, _37244_);
  or g_47595_(_37235_, _37240_, _37245_);
  or g_47596_(_37244_, _37245_, _37246_);
  or g_47597_(_37233_, _37237_, _37247_);
  or g_47598_(_37241_, _37242_, _37248_);
  or g_47599_(_37247_, _37248_, _37249_);
  or g_47600_(_37246_, _37249_, _37250_);
  xor g_47601_(out[124], out[556], _37251_);
  or g_47602_(_37228_, _37251_, _37252_);
  or g_47603_(_37227_, _37238_, _37253_);
  or g_47604_(_37252_, _37253_, _37254_);
  or g_47605_(_37231_, _37236_, _37255_);
  or g_47606_(_37239_, _37255_, _37256_);
  or g_47607_(_37254_, _37256_, _37257_);
  or g_47608_(_37250_, _37257_, _37258_);
  or g_47609_(_37243_, _37258_, _37259_);
  xor g_47610_(out[108], out[556], _37260_);
  and g_47611_(_39570_, out[555], _37261_);
  xor g_47612_(out[104], out[552], _37262_);
  xor g_47613_(out[102], out[550], _37263_);
  xor g_47614_(out[109], out[557], _37264_);
  xor g_47615_(out[110], out[558], _37265_);
  xor g_47616_(out[98], out[546], _37266_);
  xor g_47617_(out[105], out[553], _37267_);
  xor g_47618_(out[101], out[549], _37268_);
  xor g_47619_(out[97], out[545], _37269_);
  and g_47620_(out[107], _39878_, _37270_);
  or g_47621_(_37262_, _37264_, _37271_);
  xor g_47622_(out[111], out[559], _37272_);
  xor g_47623_(out[106], out[554], _37273_);
  xor g_47624_(out[100], out[548], _37274_);
  xor g_47625_(out[99], out[547], _37275_);
  xor g_47626_(out[96], out[544], _37276_);
  or g_47627_(_37266_, _37273_, _37277_);
  or g_47628_(_37271_, _37277_, _37278_);
  or g_47629_(_37267_, _37275_, _37279_);
  or g_47630_(_37268_, _37279_, _37280_);
  or g_47631_(_37278_, _37280_, _37281_);
  or g_47632_(_37265_, _37274_, _37282_);
  or g_47633_(_37281_, _37282_, _37283_);
  or g_47634_(_37260_, _37261_, _37284_);
  xor g_47635_(out[103], out[551], _37285_);
  or g_47636_(_37263_, _37285_, _37286_);
  or g_47637_(_37284_, _37286_, _37287_);
  or g_47638_(_37269_, _37270_, _37288_);
  or g_47639_(_37272_, _37288_, _37289_);
  or g_47640_(_37287_, _37289_, _37290_);
  or g_47641_(_37276_, _37290_, _37291_);
  or g_47642_(_37283_, _37291_, _37292_);
  xor g_47643_(out[87], out[551], _37293_);
  and g_47644_(_39559_, out[555], _37294_);
  xor g_47645_(out[94], out[558], _37295_);
  xor g_47646_(out[88], out[552], _37296_);
  xor g_47647_(out[81], out[545], _37297_);
  xor g_47648_(out[93], out[557], _37298_);
  xor g_47649_(out[89], out[553], _37299_);
  xor g_47650_(out[84], out[548], _37300_);
  xor g_47651_(out[82], out[546], _37301_);
  and g_47652_(out[91], _39878_, _37302_);
  xor g_47653_(out[83], out[547], _37303_);
  xor g_47654_(out[86], out[550], _37304_);
  xor g_47655_(out[95], out[559], _37305_);
  xor g_47656_(out[90], out[554], _37306_);
  xor g_47657_(out[85], out[549], _37307_);
  xor g_47658_(out[80], out[544], _37308_);
  or g_47659_(_37295_, _37300_, _37309_);
  or g_47660_(_37296_, _37298_, _37310_);
  or g_47661_(_37301_, _37306_, _37311_);
  or g_47662_(_37310_, _37311_, _37312_);
  or g_47663_(_37299_, _37303_, _37313_);
  or g_47664_(_37307_, _37308_, _37314_);
  or g_47665_(_37313_, _37314_, _37315_);
  or g_47666_(_37312_, _37315_, _37316_);
  xor g_47667_(out[92], out[556], _37317_);
  or g_47668_(_37294_, _37317_, _37318_);
  or g_47669_(_37293_, _37304_, _37319_);
  or g_47670_(_37318_, _37319_, _37320_);
  or g_47671_(_37297_, _37302_, _37321_);
  or g_47672_(_37305_, _37321_, _37322_);
  or g_47673_(_37320_, _37322_, _37323_);
  or g_47674_(_37316_, _37323_, _37324_);
  or g_47675_(_37309_, _37324_, _37325_);
  not g_47676_(_37325_, _37326_);
  xor g_47677_(out[67], out[547], _37327_);
  xor g_47678_(out[68], out[548], _37328_);
  xor g_47679_(out[78], out[558], _37329_);
  xor g_47680_(out[66], out[546], _37330_);
  xor g_47681_(out[69], out[549], _37331_);
  xor g_47682_(out[73], out[553], _37332_);
  xor g_47683_(out[72], out[552], _37333_);
  xor g_47684_(out[79], out[559], _37334_);
  xor g_47685_(out[74], out[554], _37335_);
  xor g_47686_(out[70], out[550], _37336_);
  xor g_47687_(out[64], out[544], _37337_);
  and g_47688_(_39548_, out[555], _37338_);
  and g_47689_(out[75], _39878_, _37339_);
  xor g_47690_(out[77], out[557], _37340_);
  or g_47691_(_37333_, _37340_, _37341_);
  xor g_47692_(out[65], out[545], _37342_);
  or g_47693_(_37330_, _37335_, _37343_);
  or g_47694_(_37341_, _37343_, _37344_);
  or g_47695_(_37327_, _37332_, _37345_);
  or g_47696_(_37331_, _37345_, _37346_);
  or g_47697_(_37344_, _37346_, _37347_);
  or g_47698_(_37328_, _37329_, _37348_);
  or g_47699_(_37347_, _37348_, _37349_);
  xor g_47700_(out[76], out[556], _37350_);
  or g_47701_(_37338_, _37350_, _37351_);
  xor g_47702_(out[71], out[551], _37352_);
  or g_47703_(_37336_, _37352_, _37353_);
  or g_47704_(_37351_, _37353_, _37354_);
  or g_47705_(_37339_, _37342_, _37355_);
  or g_47706_(_37334_, _37355_, _37356_);
  or g_47707_(_37354_, _37356_, _37357_);
  or g_47708_(_37337_, _37357_, _37358_);
  or g_47709_(_37349_, _37358_, _37359_);
  not g_47710_(_37359_, _37360_);
  xor g_47711_(out[55], out[551], _37361_);
  and g_47712_(_39537_, out[555], _37362_);
  xor g_47713_(out[62], out[558], _37363_);
  xor g_47714_(out[56], out[552], _37364_);
  xor g_47715_(out[49], out[545], _37365_);
  xor g_47716_(out[61], out[557], _37366_);
  xor g_47717_(out[57], out[553], _37367_);
  xor g_47718_(out[52], out[548], _37368_);
  xor g_47719_(out[50], out[546], _37369_);
  and g_47720_(out[59], _39878_, _37370_);
  xor g_47721_(out[51], out[547], _37371_);
  xor g_47722_(out[54], out[550], _37372_);
  xor g_47723_(out[63], out[559], _37373_);
  xor g_47724_(out[58], out[554], _37374_);
  xor g_47725_(out[53], out[549], _37375_);
  xor g_47726_(out[48], out[544], _37376_);
  or g_47727_(_37363_, _37368_, _37377_);
  or g_47728_(_37364_, _37366_, _37378_);
  or g_47729_(_37369_, _37374_, _37379_);
  or g_47730_(_37378_, _37379_, _37380_);
  or g_47731_(_37367_, _37371_, _37381_);
  or g_47732_(_37375_, _37376_, _37382_);
  or g_47733_(_37381_, _37382_, _37383_);
  or g_47734_(_37380_, _37383_, _37384_);
  xor g_47735_(out[60], out[556], _37385_);
  or g_47736_(_37362_, _37385_, _37386_);
  or g_47737_(_37361_, _37372_, _37387_);
  or g_47738_(_37386_, _37387_, _37388_);
  or g_47739_(_37365_, _37370_, _37389_);
  or g_47740_(_37373_, _37389_, _37390_);
  or g_47741_(_37388_, _37390_, _37391_);
  or g_47742_(_37384_, _37391_, _37392_);
  or g_47743_(_37377_, _37392_, _37393_);
  and g_47744_(out[43], _39878_, _37394_);
  xor g_47745_(out[36], out[548], _37395_);
  xor g_47746_(out[46], out[558], _37396_);
  or g_47747_(_37395_, _37396_, _37397_);
  xor g_47748_(out[45], out[557], _37398_);
  xor g_47749_(out[35], out[547], _37399_);
  xor g_47750_(out[32], out[544], _37400_);
  and g_47751_(_39526_, out[555], _37401_);
  xor g_47752_(out[42], out[554], _37402_);
  xor g_47753_(out[47], out[559], _37403_);
  xor g_47754_(out[38], out[550], _37404_);
  xor g_47755_(out[37], out[549], _37405_);
  xor g_47756_(out[40], out[552], _37406_);
  or g_47757_(_37398_, _37406_, _37407_);
  xor g_47758_(out[34], out[546], _37408_);
  xor g_47759_(out[41], out[553], _37409_);
  xor g_47760_(out[33], out[545], _37410_);
  or g_47761_(_37402_, _37408_, _37411_);
  or g_47762_(_37407_, _37411_, _37412_);
  or g_47763_(_37399_, _37409_, _37413_);
  or g_47764_(_37405_, _37413_, _37414_);
  or g_47765_(_37412_, _37414_, _37415_);
  or g_47766_(_37397_, _37415_, _37416_);
  xor g_47767_(out[44], out[556], _37417_);
  or g_47768_(_37401_, _37417_, _37418_);
  xor g_47769_(out[39], out[551], _37419_);
  or g_47770_(_37404_, _37419_, _37420_);
  or g_47771_(_37418_, _37420_, _37421_);
  or g_47772_(_37394_, _37410_, _37422_);
  or g_47773_(_37403_, _37422_, _37423_);
  or g_47774_(_37421_, _37423_, _37424_);
  or g_47775_(_37400_, _37424_, _37425_);
  or g_47776_(_37416_, _37425_, _37426_);
  xor g_47777_(out[23], out[551], _37427_);
  and g_47778_(_39493_, out[555], _37428_);
  xor g_47779_(out[30], out[558], _37429_);
  xor g_47780_(out[24], out[552], _37430_);
  xor g_47781_(out[17], out[545], _37431_);
  xor g_47782_(out[29], out[557], _37432_);
  xor g_47783_(out[25], out[553], _37433_);
  xor g_47784_(out[20], out[548], _37434_);
  xor g_47785_(out[18], out[546], _37435_);
  and g_47786_(out[27], _39878_, _37436_);
  xor g_47787_(out[19], out[547], _37437_);
  xor g_47788_(out[22], out[550], _37438_);
  xor g_47789_(out[31], out[559], _37439_);
  xor g_47790_(out[26], out[554], _37440_);
  xor g_47791_(out[21], out[549], _37441_);
  xor g_47792_(out[16], out[544], _37442_);
  or g_47793_(_37429_, _37434_, _37443_);
  or g_47794_(_37430_, _37432_, _37444_);
  or g_47795_(_37435_, _37440_, _37445_);
  or g_47796_(_37444_, _37445_, _37446_);
  or g_47797_(_37433_, _37437_, _37447_);
  or g_47798_(_37441_, _37442_, _37448_);
  or g_47799_(_37447_, _37448_, _37449_);
  or g_47800_(_37446_, _37449_, _37450_);
  xor g_47801_(out[28], out[556], _37451_);
  or g_47802_(_37428_, _37451_, _37452_);
  or g_47803_(_37427_, _37438_, _37453_);
  or g_47804_(_37452_, _37453_, _37454_);
  or g_47805_(_37431_, _37436_, _37455_);
  or g_47806_(_37439_, _37455_, _37456_);
  or g_47807_(_37454_, _37456_, _37457_);
  or g_47808_(_37450_, _37457_, _37458_);
  or g_47809_(_37443_, _37458_, _37459_);
  and g_47810_(_39438_, out[555], _37460_);
  and g_47811_(out[11], _39878_, _37461_);
  xor g_47812_(out[10], out[554], _37462_);
  xor g_47813_(out[15], out[559], _37463_);
  xor g_47814_(out[14], out[558], _37464_);
  xor g_47815_(out[0], out[544], _37465_);
  xor g_47816_(out[2], out[546], _37466_);
  xor g_47817_(out[3], out[547], _37467_);
  xor g_47818_(out[9], out[553], _37468_);
  xor g_47819_(out[1], out[545], _37469_);
  xor g_47820_(out[5], out[549], _37470_);
  xor g_47821_(out[6], out[550], _37471_);
  xor g_47822_(out[4], out[548], _37472_);
  xor g_47823_(out[13], out[557], _37473_);
  xor g_47824_(out[8], out[552], _37474_);
  or g_47825_(_37473_, _37474_, _37475_);
  or g_47826_(_37462_, _37466_, _37476_);
  or g_47827_(_37475_, _37476_, _37477_);
  or g_47828_(_37467_, _37468_, _37478_);
  or g_47829_(_37470_, _37478_, _37479_);
  or g_47830_(_37477_, _37479_, _37480_);
  or g_47831_(_37464_, _37472_, _37481_);
  or g_47832_(_37480_, _37481_, _37482_);
  xor g_47833_(out[12], out[556], _37483_);
  or g_47834_(_37460_, _37483_, _37484_);
  xor g_47835_(out[7], out[551], _37485_);
  or g_47836_(_37471_, _37485_, _37486_);
  or g_47837_(_37484_, _37486_, _37487_);
  or g_47838_(_37461_, _37469_, _37488_);
  or g_47839_(_37463_, _37488_, _37489_);
  or g_47840_(_37487_, _37489_, _37490_);
  or g_47841_(_37465_, _37490_, _37491_);
  or g_47842_(_37482_, _37491_, _37492_);
  xor g_47843_(out[305], out[529], _37493_);
  and g_47844_(out[315], _39867_, _37494_);
  xor g_47845_(out[313], out[537], _37495_);
  xor g_47846_(out[304], out[528], _37496_);
  xor g_47847_(out[318], out[542], _37497_);
  xor g_47848_(out[308], out[532], _37498_);
  or g_47849_(_37497_, _37498_, _37499_);
  xor g_47850_(out[317], out[541], _37500_);
  xor g_47851_(out[307], out[531], _37501_);
  and g_47852_(_39724_, out[539], _37502_);
  xor g_47853_(out[310], out[534], _37503_);
  xor g_47854_(out[314], out[538], _37504_);
  xor g_47855_(out[309], out[533], _37505_);
  xor g_47856_(out[319], out[543], _37506_);
  xor g_47857_(out[312], out[536], _37507_);
  or g_47858_(_37500_, _37507_, _37508_);
  xor g_47859_(out[306], out[530], _37509_);
  or g_47860_(_37504_, _37509_, _37510_);
  or g_47861_(_37508_, _37510_, _37511_);
  or g_47862_(_37495_, _37501_, _37512_);
  or g_47863_(_37505_, _37512_, _37513_);
  or g_47864_(_37511_, _37513_, _37514_);
  or g_47865_(_37499_, _37514_, _37515_);
  xor g_47866_(out[316], out[540], _37516_);
  or g_47867_(_37502_, _37516_, _37517_);
  xor g_47868_(out[311], out[535], _37518_);
  or g_47869_(_37503_, _37518_, _37519_);
  or g_47870_(_37517_, _37519_, _37520_);
  or g_47871_(_37493_, _37494_, _37521_);
  or g_47872_(_37506_, _37521_, _37522_);
  or g_47873_(_37520_, _37522_, _37523_);
  or g_47874_(_37496_, _37523_, _37524_);
  or g_47875_(_37515_, _37524_, _37525_);
  xor g_47876_(out[295], out[535], _37526_);
  and g_47877_(_39702_, out[539], _37527_);
  xor g_47878_(out[302], out[542], _37528_);
  xor g_47879_(out[296], out[536], _37529_);
  xor g_47880_(out[289], out[529], _37530_);
  xor g_47881_(out[301], out[541], _37531_);
  xor g_47882_(out[297], out[537], _37532_);
  xor g_47883_(out[292], out[532], _37533_);
  xor g_47884_(out[290], out[530], _37534_);
  and g_47885_(out[299], _39867_, _37535_);
  xor g_47886_(out[291], out[531], _37536_);
  xor g_47887_(out[294], out[534], _37537_);
  xor g_47888_(out[303], out[543], _37538_);
  xor g_47889_(out[298], out[538], _37539_);
  xor g_47890_(out[293], out[533], _37540_);
  xor g_47891_(out[288], out[528], _37541_);
  or g_47892_(_37528_, _37533_, _37542_);
  or g_47893_(_37529_, _37531_, _37543_);
  or g_47894_(_37534_, _37539_, _37544_);
  or g_47895_(_37543_, _37544_, _37545_);
  or g_47896_(_37532_, _37536_, _37546_);
  or g_47897_(_37540_, _37541_, _37547_);
  or g_47898_(_37546_, _37547_, _37548_);
  or g_47899_(_37545_, _37548_, _37549_);
  xor g_47900_(out[300], out[540], _37550_);
  or g_47901_(_37527_, _37550_, _37551_);
  or g_47902_(_37526_, _37537_, _37552_);
  or g_47903_(_37551_, _37552_, _37553_);
  or g_47904_(_37530_, _37535_, _37554_);
  or g_47905_(_37538_, _37554_, _37555_);
  or g_47906_(_37553_, _37555_, _37556_);
  or g_47907_(_37549_, _37556_, _37557_);
  or g_47908_(_37542_, _37557_, _37558_);
  xor g_47909_(out[273], out[529], _37559_);
  and g_47910_(out[283], _39867_, _37560_);
  xor g_47911_(out[281], out[537], _37561_);
  xor g_47912_(out[272], out[528], _37562_);
  xor g_47913_(out[286], out[542], _37563_);
  xor g_47914_(out[276], out[532], _37564_);
  or g_47915_(_37563_, _37564_, _37565_);
  xor g_47916_(out[285], out[541], _37566_);
  xor g_47917_(out[275], out[531], _37567_);
  and g_47918_(_39691_, out[539], _37568_);
  xor g_47919_(out[278], out[534], _37569_);
  xor g_47920_(out[282], out[538], _37570_);
  xor g_47921_(out[277], out[533], _37571_);
  xor g_47922_(out[287], out[543], _37572_);
  xor g_47923_(out[280], out[536], _37573_);
  or g_47924_(_37566_, _37573_, _37574_);
  xor g_47925_(out[274], out[530], _37575_);
  or g_47926_(_37570_, _37575_, _37576_);
  or g_47927_(_37574_, _37576_, _37577_);
  or g_47928_(_37561_, _37567_, _37578_);
  or g_47929_(_37571_, _37578_, _37579_);
  or g_47930_(_37577_, _37579_, _37580_);
  or g_47931_(_37565_, _37580_, _37581_);
  xor g_47932_(out[284], out[540], _37582_);
  or g_47933_(_37568_, _37582_, _37583_);
  xor g_47934_(out[279], out[535], _37584_);
  or g_47935_(_37569_, _37584_, _37585_);
  or g_47936_(_37583_, _37585_, _37586_);
  or g_47937_(_37559_, _37560_, _37587_);
  or g_47938_(_37572_, _37587_, _37588_);
  or g_47939_(_37586_, _37588_, _37589_);
  or g_47940_(_37562_, _37589_, _37590_);
  or g_47941_(_37581_, _37590_, _37591_);
  xor g_47942_(out[263], out[535], _37592_);
  and g_47943_(_39680_, out[539], _37593_);
  xor g_47944_(out[270], out[542], _37594_);
  xor g_47945_(out[264], out[536], _37595_);
  xor g_47946_(out[257], out[529], _37596_);
  xor g_47947_(out[269], out[541], _37597_);
  xor g_47948_(out[265], out[537], _37598_);
  xor g_47949_(out[260], out[532], _37599_);
  xor g_47950_(out[258], out[530], _37600_);
  and g_47951_(out[267], _39867_, _37601_);
  xor g_47952_(out[259], out[531], _37602_);
  xor g_47953_(out[262], out[534], _37603_);
  xor g_47954_(out[271], out[543], _37604_);
  xor g_47955_(out[266], out[538], _37605_);
  xor g_47956_(out[261], out[533], _37606_);
  xor g_47957_(out[256], out[528], _37607_);
  or g_47958_(_37594_, _37599_, _37608_);
  or g_47959_(_37595_, _37597_, _37609_);
  or g_47960_(_37600_, _37605_, _37610_);
  or g_47961_(_37609_, _37610_, _37611_);
  or g_47962_(_37598_, _37602_, _37612_);
  or g_47963_(_37606_, _37607_, _37613_);
  or g_47964_(_37612_, _37613_, _37614_);
  or g_47965_(_37611_, _37614_, _37615_);
  xor g_47966_(out[268], out[540], _37616_);
  or g_47967_(_37593_, _37616_, _37617_);
  or g_47968_(_37592_, _37603_, _37618_);
  or g_47969_(_37617_, _37618_, _37619_);
  or g_47970_(_37596_, _37601_, _37620_);
  or g_47971_(_37604_, _37620_, _37621_);
  or g_47972_(_37619_, _37621_, _37622_);
  or g_47973_(_37615_, _37622_, _37623_);
  or g_47974_(_37608_, _37623_, _37624_);
  xor g_47975_(out[241], out[529], _37625_);
  and g_47976_(out[251], _39867_, _37626_);
  xor g_47977_(out[249], out[537], _37627_);
  xor g_47978_(out[240], out[528], _37628_);
  xor g_47979_(out[254], out[542], _37629_);
  xor g_47980_(out[244], out[532], _37630_);
  or g_47981_(_37629_, _37630_, _37631_);
  xor g_47982_(out[253], out[541], _37632_);
  xor g_47983_(out[243], out[531], _37633_);
  and g_47984_(_39669_, out[539], _37634_);
  xor g_47985_(out[246], out[534], _37635_);
  xor g_47986_(out[250], out[538], _37636_);
  xor g_47987_(out[245], out[533], _37637_);
  xor g_47988_(out[255], out[543], _37638_);
  xor g_47989_(out[248], out[536], _37639_);
  or g_47990_(_37632_, _37639_, _37640_);
  xor g_47991_(out[242], out[530], _37641_);
  or g_47992_(_37636_, _37641_, _37642_);
  or g_47993_(_37640_, _37642_, _37643_);
  or g_47994_(_37627_, _37633_, _37644_);
  or g_47995_(_37637_, _37644_, _37645_);
  or g_47996_(_37643_, _37645_, _37646_);
  or g_47997_(_37631_, _37646_, _37647_);
  xor g_47998_(out[252], out[540], _37648_);
  or g_47999_(_37634_, _37648_, _37649_);
  xor g_48000_(out[247], out[535], _37650_);
  or g_48001_(_37635_, _37650_, _37651_);
  or g_48002_(_37649_, _37651_, _37652_);
  or g_48003_(_37625_, _37626_, _37653_);
  or g_48004_(_37638_, _37653_, _37654_);
  or g_48005_(_37652_, _37654_, _37655_);
  or g_48006_(_37628_, _37655_, _37656_);
  or g_48007_(_37647_, _37656_, _37657_);
  xor g_48008_(out[231], out[535], _37658_);
  and g_48009_(_39658_, out[539], _37659_);
  xor g_48010_(out[238], out[542], _37660_);
  xor g_48011_(out[232], out[536], _37661_);
  xor g_48012_(out[225], out[529], _37662_);
  xor g_48013_(out[237], out[541], _37663_);
  xor g_48014_(out[233], out[537], _37664_);
  xor g_48015_(out[228], out[532], _37665_);
  xor g_48016_(out[226], out[530], _37666_);
  and g_48017_(out[235], _39867_, _37667_);
  xor g_48018_(out[227], out[531], _37668_);
  xor g_48019_(out[230], out[534], _37669_);
  xor g_48020_(out[239], out[543], _37670_);
  xor g_48021_(out[234], out[538], _37671_);
  xor g_48022_(out[229], out[533], _37672_);
  xor g_48023_(out[224], out[528], _37673_);
  or g_48024_(_37660_, _37665_, _37674_);
  or g_48025_(_37661_, _37663_, _37675_);
  or g_48026_(_37666_, _37671_, _37676_);
  or g_48027_(_37675_, _37676_, _37677_);
  or g_48028_(_37664_, _37668_, _37678_);
  or g_48029_(_37672_, _37673_, _37679_);
  or g_48030_(_37678_, _37679_, _37680_);
  or g_48031_(_37677_, _37680_, _37681_);
  xor g_48032_(out[236], out[540], _37682_);
  or g_48033_(_37659_, _37682_, _37683_);
  or g_48034_(_37658_, _37669_, _37684_);
  or g_48035_(_37683_, _37684_, _37685_);
  or g_48036_(_37662_, _37667_, _37686_);
  or g_48037_(_37670_, _37686_, _37687_);
  or g_48038_(_37685_, _37687_, _37688_);
  or g_48039_(_37681_, _37688_, _37689_);
  or g_48040_(_37674_, _37689_, _37690_);
  xor g_48041_(out[209], out[529], _37691_);
  and g_48042_(out[219], _39867_, _37692_);
  xor g_48043_(out[217], out[537], _37693_);
  xor g_48044_(out[208], out[528], _37694_);
  xor g_48045_(out[222], out[542], _37695_);
  xor g_48046_(out[212], out[532], _37696_);
  or g_48047_(_37695_, _37696_, _37697_);
  xor g_48048_(out[221], out[541], _37698_);
  xor g_48049_(out[211], out[531], _37699_);
  and g_48050_(_39647_, out[539], _37700_);
  xor g_48051_(out[214], out[534], _37701_);
  xor g_48052_(out[218], out[538], _37702_);
  xor g_48053_(out[213], out[533], _37703_);
  xor g_48054_(out[223], out[543], _37704_);
  xor g_48055_(out[216], out[536], _37705_);
  or g_48056_(_37698_, _37705_, _37706_);
  xor g_48057_(out[210], out[530], _37707_);
  or g_48058_(_37702_, _37707_, _37708_);
  or g_48059_(_37706_, _37708_, _37709_);
  or g_48060_(_37693_, _37699_, _37710_);
  or g_48061_(_37703_, _37710_, _37711_);
  or g_48062_(_37709_, _37711_, _37712_);
  or g_48063_(_37697_, _37712_, _37713_);
  xor g_48064_(out[220], out[540], _37714_);
  or g_48065_(_37700_, _37714_, _37715_);
  xor g_48066_(out[215], out[535], _37716_);
  or g_48067_(_37701_, _37716_, _37717_);
  or g_48068_(_37715_, _37717_, _37718_);
  or g_48069_(_37691_, _37692_, _37719_);
  or g_48070_(_37704_, _37719_, _37720_);
  or g_48071_(_37718_, _37720_, _37721_);
  or g_48072_(_37694_, _37721_, _37722_);
  or g_48073_(_37713_, _37722_, _37723_);
  xor g_48074_(out[199], out[535], _37724_);
  and g_48075_(_39636_, out[539], _37725_);
  xor g_48076_(out[206], out[542], _37726_);
  xor g_48077_(out[200], out[536], _37727_);
  xor g_48078_(out[193], out[529], _37728_);
  xor g_48079_(out[205], out[541], _37729_);
  xor g_48080_(out[201], out[537], _37730_);
  xor g_48081_(out[196], out[532], _37731_);
  xor g_48082_(out[194], out[530], _37732_);
  and g_48083_(out[203], _39867_, _37733_);
  xor g_48084_(out[195], out[531], _37734_);
  xor g_48085_(out[198], out[534], _37735_);
  xor g_48086_(out[207], out[543], _37736_);
  xor g_48087_(out[202], out[538], _37737_);
  xor g_48088_(out[197], out[533], _37738_);
  xor g_48089_(out[192], out[528], _37739_);
  or g_48090_(_37726_, _37731_, _37740_);
  or g_48091_(_37727_, _37729_, _37741_);
  or g_48092_(_37732_, _37737_, _37742_);
  or g_48093_(_37741_, _37742_, _37743_);
  or g_48094_(_37730_, _37734_, _37744_);
  or g_48095_(_37738_, _37739_, _37745_);
  or g_48096_(_37744_, _37745_, _37746_);
  or g_48097_(_37743_, _37746_, _37747_);
  xor g_48098_(out[204], out[540], _37748_);
  or g_48099_(_37725_, _37748_, _37749_);
  or g_48100_(_37724_, _37735_, _37750_);
  or g_48101_(_37749_, _37750_, _37751_);
  or g_48102_(_37728_, _37733_, _37752_);
  or g_48103_(_37736_, _37752_, _37753_);
  or g_48104_(_37751_, _37753_, _37754_);
  or g_48105_(_37747_, _37754_, _37755_);
  or g_48106_(_37740_, _37755_, _37756_);
  xor g_48107_(out[177], out[529], _37757_);
  and g_48108_(out[187], _39867_, _37758_);
  xor g_48109_(out[185], out[537], _37759_);
  xor g_48110_(out[176], out[528], _37760_);
  xor g_48111_(out[190], out[542], _37761_);
  xor g_48112_(out[180], out[532], _37762_);
  or g_48113_(_37761_, _37762_, _37763_);
  xor g_48114_(out[189], out[541], _37764_);
  xor g_48115_(out[179], out[531], _37765_);
  and g_48116_(_39625_, out[539], _37766_);
  xor g_48117_(out[182], out[534], _37767_);
  xor g_48118_(out[186], out[538], _37768_);
  xor g_48119_(out[181], out[533], _37769_);
  xor g_48120_(out[191], out[543], _37770_);
  xor g_48121_(out[184], out[536], _37771_);
  or g_48122_(_37764_, _37771_, _37772_);
  xor g_48123_(out[178], out[530], _37773_);
  or g_48124_(_37768_, _37773_, _37774_);
  or g_48125_(_37772_, _37774_, _37775_);
  or g_48126_(_37759_, _37765_, _37776_);
  or g_48127_(_37769_, _37776_, _37777_);
  or g_48128_(_37775_, _37777_, _37778_);
  or g_48129_(_37763_, _37778_, _37779_);
  xor g_48130_(out[188], out[540], _37780_);
  or g_48131_(_37766_, _37780_, _37781_);
  xor g_48132_(out[183], out[535], _37782_);
  or g_48133_(_37767_, _37782_, _37783_);
  or g_48134_(_37781_, _37783_, _37784_);
  or g_48135_(_37757_, _37758_, _37785_);
  or g_48136_(_37770_, _37785_, _37786_);
  or g_48137_(_37784_, _37786_, _37787_);
  or g_48138_(_37760_, _37787_, _37788_);
  or g_48139_(_37779_, _37788_, _37789_);
  xor g_48140_(out[167], out[535], _37790_);
  and g_48141_(_39614_, out[539], _37791_);
  xor g_48142_(out[174], out[542], _37792_);
  xor g_48143_(out[168], out[536], _37793_);
  xor g_48144_(out[161], out[529], _37794_);
  xor g_48145_(out[173], out[541], _37795_);
  xor g_48146_(out[169], out[537], _37796_);
  xor g_48147_(out[164], out[532], _37797_);
  xor g_48148_(out[162], out[530], _37798_);
  and g_48149_(out[171], _39867_, _37799_);
  xor g_48150_(out[163], out[531], _37800_);
  xor g_48151_(out[166], out[534], _37801_);
  xor g_48152_(out[175], out[543], _37802_);
  xor g_48153_(out[170], out[538], _37803_);
  xor g_48154_(out[165], out[533], _37804_);
  xor g_48155_(out[160], out[528], _37805_);
  or g_48156_(_37792_, _37797_, _37806_);
  or g_48157_(_37793_, _37795_, _37807_);
  or g_48158_(_37798_, _37803_, _37808_);
  or g_48159_(_37807_, _37808_, _37809_);
  or g_48160_(_37796_, _37800_, _37810_);
  or g_48161_(_37804_, _37805_, _37811_);
  or g_48162_(_37810_, _37811_, _37812_);
  or g_48163_(_37809_, _37812_, _37813_);
  xor g_48164_(out[172], out[540], _37814_);
  or g_48165_(_37791_, _37814_, _37815_);
  or g_48166_(_37790_, _37801_, _37816_);
  or g_48167_(_37815_, _37816_, _37817_);
  or g_48168_(_37794_, _37799_, _37818_);
  or g_48169_(_37802_, _37818_, _37819_);
  or g_48170_(_37817_, _37819_, _37820_);
  or g_48171_(_37813_, _37820_, _37821_);
  or g_48172_(_37806_, _37821_, _37822_);
  xor g_48173_(out[145], out[529], _37823_);
  and g_48174_(out[155], _39867_, _37824_);
  xor g_48175_(out[158], out[542], _37825_);
  xor g_48176_(out[147], out[531], _37826_);
  xor g_48177_(out[148], out[532], _37827_);
  xor g_48178_(out[146], out[530], _37828_);
  xor g_48179_(out[153], out[537], _37829_);
  xor g_48180_(out[144], out[528], _37830_);
  and g_48181_(_39603_, out[539], _37831_);
  xor g_48182_(out[150], out[534], _37832_);
  xor g_48183_(out[154], out[538], _37833_);
  xor g_48184_(out[149], out[533], _37834_);
  xor g_48185_(out[159], out[543], _37835_);
  xor g_48186_(out[157], out[541], _37836_);
  xor g_48187_(out[152], out[536], _37837_);
  or g_48188_(_37825_, _37827_, _37838_);
  or g_48189_(_37836_, _37837_, _37839_);
  or g_48190_(_37828_, _37833_, _37840_);
  or g_48191_(_37839_, _37840_, _37841_);
  or g_48192_(_37826_, _37829_, _37842_);
  or g_48193_(_37830_, _37834_, _37843_);
  or g_48194_(_37842_, _37843_, _37844_);
  or g_48195_(_37841_, _37844_, _37845_);
  xor g_48196_(out[156], out[540], _37846_);
  or g_48197_(_37831_, _37846_, _37847_);
  xor g_48198_(out[151], out[535], _37848_);
  or g_48199_(_37832_, _37848_, _37849_);
  or g_48200_(_37847_, _37849_, _37850_);
  or g_48201_(_37823_, _37824_, _37851_);
  or g_48202_(_37835_, _37851_, _37852_);
  or g_48203_(_37850_, _37852_, _37853_);
  or g_48204_(_37845_, _37853_, _37854_);
  or g_48205_(_37838_, _37854_, _37855_);
  xor g_48206_(out[135], out[535], _37856_);
  and g_48207_(_39592_, out[539], _37857_);
  xor g_48208_(out[142], out[542], _37858_);
  xor g_48209_(out[136], out[536], _37859_);
  xor g_48210_(out[129], out[529], _37860_);
  xor g_48211_(out[141], out[541], _37861_);
  xor g_48212_(out[137], out[537], _37862_);
  xor g_48213_(out[132], out[532], _37863_);
  xor g_48214_(out[130], out[530], _37864_);
  and g_48215_(out[139], _39867_, _37865_);
  xor g_48216_(out[131], out[531], _37866_);
  xor g_48217_(out[134], out[534], _37867_);
  xor g_48218_(out[143], out[543], _37868_);
  xor g_48219_(out[138], out[538], _37869_);
  xor g_48220_(out[133], out[533], _37870_);
  xor g_48221_(out[128], out[528], _37871_);
  or g_48222_(_37858_, _37863_, _37872_);
  or g_48223_(_37859_, _37861_, _37873_);
  or g_48224_(_37864_, _37869_, _37874_);
  or g_48225_(_37873_, _37874_, _37875_);
  or g_48226_(_37862_, _37866_, _37876_);
  or g_48227_(_37870_, _37871_, _37877_);
  or g_48228_(_37876_, _37877_, _37878_);
  or g_48229_(_37875_, _37878_, _37879_);
  xor g_48230_(out[140], out[540], _37880_);
  or g_48231_(_37857_, _37880_, _37881_);
  or g_48232_(_37856_, _37867_, _37882_);
  or g_48233_(_37881_, _37882_, _37883_);
  or g_48234_(_37860_, _37865_, _37884_);
  or g_48235_(_37868_, _37884_, _37885_);
  or g_48236_(_37883_, _37885_, _37886_);
  or g_48237_(_37879_, _37886_, _37887_);
  or g_48238_(_37872_, _37887_, _37888_);
  xor g_48239_(out[122], out[538], _37889_);
  xor g_48240_(out[114], out[530], _37890_);
  xor g_48241_(out[113], out[529], _37891_);
  and g_48242_(_39581_, out[539], _37892_);
  and g_48243_(out[123], _39867_, _37893_);
  xor g_48244_(out[125], out[541], _37894_);
  xor g_48245_(out[115], out[531], _37895_);
  xor g_48246_(out[126], out[542], _37896_);
  xor g_48247_(out[124], out[540], _37897_);
  xor g_48248_(out[120], out[536], _37898_);
  xor g_48249_(out[127], out[543], _37899_);
  xor g_48250_(out[117], out[533], _37900_);
  xor g_48251_(out[118], out[534], _37901_);
  xor g_48252_(out[112], out[528], _37902_);
  xor g_48253_(out[116], out[532], _37903_);
  or g_48254_(_37894_, _37898_, _37904_);
  xor g_48255_(out[121], out[537], _37905_);
  or g_48256_(_37889_, _37890_, _37906_);
  or g_48257_(_37904_, _37906_, _37907_);
  or g_48258_(_37895_, _37905_, _37908_);
  or g_48259_(_37900_, _37908_, _37909_);
  or g_48260_(_37907_, _37909_, _37910_);
  or g_48261_(_37896_, _37903_, _37911_);
  or g_48262_(_37910_, _37911_, _37912_);
  or g_48263_(_37892_, _37897_, _37913_);
  xor g_48264_(out[119], out[535], _37914_);
  or g_48265_(_37901_, _37914_, _37915_);
  or g_48266_(_37913_, _37915_, _37916_);
  or g_48267_(_37891_, _37893_, _37917_);
  or g_48268_(_37899_, _37917_, _37918_);
  or g_48269_(_37916_, _37918_, _37919_);
  or g_48270_(_37902_, _37919_, _37920_);
  or g_48271_(_37912_, _37920_, _37921_);
  xor g_48272_(out[103], out[535], _37922_);
  and g_48273_(_39570_, out[539], _37923_);
  xor g_48274_(out[110], out[542], _37924_);
  xor g_48275_(out[104], out[536], _37925_);
  xor g_48276_(out[97], out[529], _37926_);
  xor g_48277_(out[109], out[541], _37927_);
  xor g_48278_(out[105], out[537], _37928_);
  xor g_48279_(out[100], out[532], _37929_);
  xor g_48280_(out[98], out[530], _37930_);
  and g_48281_(out[107], _39867_, _37931_);
  xor g_48282_(out[99], out[531], _37932_);
  xor g_48283_(out[102], out[534], _37933_);
  xor g_48284_(out[111], out[543], _37934_);
  xor g_48285_(out[106], out[538], _37935_);
  xor g_48286_(out[101], out[533], _37936_);
  xor g_48287_(out[96], out[528], _37937_);
  or g_48288_(_37924_, _37929_, _37938_);
  or g_48289_(_37925_, _37927_, _37939_);
  or g_48290_(_37930_, _37935_, _37940_);
  or g_48291_(_37939_, _37940_, _37941_);
  or g_48292_(_37928_, _37932_, _37942_);
  or g_48293_(_37936_, _37937_, _37943_);
  or g_48294_(_37942_, _37943_, _37944_);
  or g_48295_(_37941_, _37944_, _37945_);
  xor g_48296_(out[108], out[540], _37946_);
  or g_48297_(_37923_, _37946_, _37947_);
  or g_48298_(_37922_, _37933_, _37948_);
  or g_48299_(_37947_, _37948_, _37949_);
  or g_48300_(_37926_, _37931_, _37950_);
  or g_48301_(_37934_, _37950_, _37951_);
  or g_48302_(_37949_, _37951_, _37952_);
  or g_48303_(_37945_, _37952_, _37953_);
  or g_48304_(_37938_, _37953_, _37954_);
  xor g_48305_(out[81], out[529], _37955_);
  and g_48306_(out[91], _39867_, _37956_);
  xor g_48307_(out[89], out[537], _37957_);
  xor g_48308_(out[80], out[528], _37958_);
  xor g_48309_(out[94], out[542], _37959_);
  xor g_48310_(out[84], out[532], _37960_);
  or g_48311_(_37959_, _37960_, _37961_);
  xor g_48312_(out[93], out[541], _37962_);
  xor g_48313_(out[83], out[531], _37963_);
  and g_48314_(_39559_, out[539], _37964_);
  xor g_48315_(out[86], out[534], _37965_);
  xor g_48316_(out[90], out[538], _37966_);
  xor g_48317_(out[85], out[533], _37967_);
  xor g_48318_(out[95], out[543], _37968_);
  xor g_48319_(out[88], out[536], _37969_);
  or g_48320_(_37962_, _37969_, _37970_);
  xor g_48321_(out[82], out[530], _37971_);
  or g_48322_(_37966_, _37971_, _37972_);
  or g_48323_(_37970_, _37972_, _37973_);
  or g_48324_(_37957_, _37963_, _37974_);
  or g_48325_(_37967_, _37974_, _37975_);
  or g_48326_(_37973_, _37975_, _37976_);
  or g_48327_(_37961_, _37976_, _37977_);
  xor g_48328_(out[92], out[540], _37978_);
  or g_48329_(_37964_, _37978_, _37979_);
  xor g_48330_(out[87], out[535], _37980_);
  or g_48331_(_37965_, _37980_, _37981_);
  or g_48332_(_37979_, _37981_, _37982_);
  or g_48333_(_37955_, _37956_, _37983_);
  or g_48334_(_37968_, _37983_, _37984_);
  or g_48335_(_37982_, _37984_, _37985_);
  or g_48336_(_37958_, _37985_, _37986_);
  or g_48337_(_37977_, _37986_, _37987_);
  xor g_48338_(out[71], out[535], _37988_);
  and g_48339_(_39548_, out[539], _37989_);
  xor g_48340_(out[78], out[542], _37990_);
  xor g_48341_(out[72], out[536], _37991_);
  xor g_48342_(out[65], out[529], _37992_);
  xor g_48343_(out[77], out[541], _37993_);
  xor g_48344_(out[73], out[537], _37994_);
  xor g_48345_(out[68], out[532], _37995_);
  xor g_48346_(out[66], out[530], _37996_);
  and g_48347_(out[75], _39867_, _37997_);
  xor g_48348_(out[67], out[531], _37998_);
  xor g_48349_(out[70], out[534], _37999_);
  xor g_48350_(out[79], out[543], _38000_);
  xor g_48351_(out[74], out[538], _38001_);
  xor g_48352_(out[69], out[533], _38002_);
  xor g_48353_(out[64], out[528], _38003_);
  or g_48354_(_37990_, _37995_, _38004_);
  or g_48355_(_37991_, _37993_, _38005_);
  or g_48356_(_37996_, _38001_, _38006_);
  or g_48357_(_38005_, _38006_, _38007_);
  or g_48358_(_37994_, _37998_, _38008_);
  or g_48359_(_38002_, _38003_, _38009_);
  or g_48360_(_38008_, _38009_, _38010_);
  or g_48361_(_38007_, _38010_, _38011_);
  xor g_48362_(out[76], out[540], _38012_);
  or g_48363_(_37989_, _38012_, _38013_);
  or g_48364_(_37988_, _37999_, _38014_);
  or g_48365_(_38013_, _38014_, _38015_);
  or g_48366_(_37992_, _37997_, _38016_);
  or g_48367_(_38000_, _38016_, _38017_);
  or g_48368_(_38015_, _38017_, _38018_);
  or g_48369_(_38011_, _38018_, _38019_);
  or g_48370_(_38004_, _38019_, _38020_);
  xor g_48371_(out[49], out[529], _38021_);
  and g_48372_(out[59], _39867_, _38022_);
  xor g_48373_(out[57], out[537], _38023_);
  xor g_48374_(out[48], out[528], _38024_);
  xor g_48375_(out[62], out[542], _38025_);
  xor g_48376_(out[52], out[532], _38026_);
  or g_48377_(_38025_, _38026_, _38027_);
  xor g_48378_(out[61], out[541], _38028_);
  xor g_48379_(out[51], out[531], _38029_);
  and g_48380_(_39537_, out[539], _38030_);
  xor g_48381_(out[54], out[534], _38031_);
  xor g_48382_(out[58], out[538], _38032_);
  xor g_48383_(out[53], out[533], _38033_);
  xor g_48384_(out[63], out[543], _38034_);
  xor g_48385_(out[56], out[536], _38035_);
  or g_48386_(_38028_, _38035_, _38036_);
  xor g_48387_(out[50], out[530], _38037_);
  or g_48388_(_38032_, _38037_, _38038_);
  or g_48389_(_38036_, _38038_, _38039_);
  or g_48390_(_38023_, _38029_, _38040_);
  or g_48391_(_38033_, _38040_, _38041_);
  or g_48392_(_38039_, _38041_, _38042_);
  or g_48393_(_38027_, _38042_, _38043_);
  xor g_48394_(out[60], out[540], _38044_);
  or g_48395_(_38030_, _38044_, _38045_);
  xor g_48396_(out[55], out[535], _38046_);
  or g_48397_(_38031_, _38046_, _38047_);
  or g_48398_(_38045_, _38047_, _38048_);
  or g_48399_(_38021_, _38022_, _38049_);
  or g_48400_(_38034_, _38049_, _38050_);
  or g_48401_(_38048_, _38050_, _38051_);
  or g_48402_(_38024_, _38051_, _38052_);
  or g_48403_(_38043_, _38052_, _38053_);
  xor g_48404_(out[39], out[535], _38054_);
  and g_48405_(_39526_, out[539], _38055_);
  xor g_48406_(out[46], out[542], _38056_);
  xor g_48407_(out[40], out[536], _38057_);
  xor g_48408_(out[33], out[529], _38058_);
  xor g_48409_(out[45], out[541], _38059_);
  xor g_48410_(out[41], out[537], _38060_);
  xor g_48411_(out[36], out[532], _38061_);
  xor g_48412_(out[34], out[530], _38062_);
  and g_48413_(out[43], _39867_, _38063_);
  xor g_48414_(out[35], out[531], _38064_);
  xor g_48415_(out[38], out[534], _38065_);
  xor g_48416_(out[47], out[543], _38066_);
  xor g_48417_(out[42], out[538], _38067_);
  xor g_48418_(out[37], out[533], _38068_);
  xor g_48419_(out[32], out[528], _38069_);
  or g_48420_(_38056_, _38061_, _38070_);
  or g_48421_(_38057_, _38059_, _38071_);
  or g_48422_(_38062_, _38067_, _38072_);
  or g_48423_(_38071_, _38072_, _38073_);
  or g_48424_(_38060_, _38064_, _38074_);
  or g_48425_(_38068_, _38069_, _38075_);
  or g_48426_(_38074_, _38075_, _38076_);
  or g_48427_(_38073_, _38076_, _38077_);
  xor g_48428_(out[44], out[540], _38078_);
  or g_48429_(_38055_, _38078_, _38079_);
  or g_48430_(_38054_, _38065_, _38080_);
  or g_48431_(_38079_, _38080_, _38081_);
  or g_48432_(_38058_, _38063_, _38082_);
  or g_48433_(_38066_, _38082_, _38083_);
  or g_48434_(_38081_, _38083_, _38084_);
  or g_48435_(_38077_, _38084_, _38085_);
  or g_48436_(_38070_, _38085_, _38086_);
  xor g_48437_(out[17], out[529], _38087_);
  and g_48438_(out[27], _39867_, _38088_);
  xor g_48439_(out[25], out[537], _38089_);
  xor g_48440_(out[16], out[528], _38090_);
  xor g_48441_(out[30], out[542], _38091_);
  xor g_48442_(out[20], out[532], _38092_);
  or g_48443_(_38091_, _38092_, _38093_);
  xor g_48444_(out[29], out[541], _38094_);
  xor g_48445_(out[19], out[531], _38095_);
  and g_48446_(_39493_, out[539], _38096_);
  xor g_48447_(out[22], out[534], _38097_);
  xor g_48448_(out[26], out[538], _38098_);
  xor g_48449_(out[21], out[533], _38099_);
  xor g_48450_(out[31], out[543], _38100_);
  xor g_48451_(out[24], out[536], _38101_);
  or g_48452_(_38094_, _38101_, _38102_);
  xor g_48453_(out[18], out[530], _38103_);
  or g_48454_(_38098_, _38103_, _38104_);
  or g_48455_(_38102_, _38104_, _38105_);
  or g_48456_(_38089_, _38095_, _38106_);
  or g_48457_(_38099_, _38106_, _38107_);
  or g_48458_(_38105_, _38107_, _38108_);
  or g_48459_(_38093_, _38108_, _38109_);
  xor g_48460_(out[28], out[540], _38110_);
  or g_48461_(_38096_, _38110_, _38111_);
  xor g_48462_(out[23], out[535], _38112_);
  or g_48463_(_38097_, _38112_, _38113_);
  or g_48464_(_38111_, _38113_, _38114_);
  or g_48465_(_38087_, _38088_, _38115_);
  or g_48466_(_38100_, _38115_, _38116_);
  or g_48467_(_38114_, _38116_, _38117_);
  or g_48468_(_38090_, _38117_, _38118_);
  or g_48469_(_38109_, _38118_, _38119_);
  xor g_48470_(out[1], out[529], _38120_);
  and g_48471_(_39438_, out[539], _38121_);
  and g_48472_(out[11], _39867_, _38122_);
  xor g_48473_(out[13], out[541], _38123_);
  xor g_48474_(out[10], out[538], _38124_);
  xor g_48475_(out[4], out[532], _38125_);
  xor g_48476_(out[14], out[542], _38126_);
  or g_48477_(_38125_, _38126_, _38127_);
  xor g_48478_(out[8], out[536], _38128_);
  xor g_48479_(out[0], out[528], _38129_);
  xor g_48480_(out[2], out[530], _38130_);
  xor g_48481_(out[9], out[537], _38131_);
  xor g_48482_(out[5], out[533], _38132_);
  xor g_48483_(out[3], out[531], _38133_);
  xor g_48484_(out[15], out[543], _38134_);
  xor g_48485_(out[6], out[534], _38135_);
  or g_48486_(_38123_, _38128_, _38136_);
  or g_48487_(_38124_, _38130_, _38137_);
  or g_48488_(_38136_, _38137_, _38138_);
  or g_48489_(_38131_, _38133_, _38139_);
  or g_48490_(_38129_, _38132_, _38140_);
  or g_48491_(_38139_, _38140_, _38141_);
  or g_48492_(_38138_, _38141_, _38142_);
  xor g_48493_(out[12], out[540], _38143_);
  or g_48494_(_38121_, _38143_, _38144_);
  xor g_48495_(out[7], out[535], _38145_);
  or g_48496_(_38135_, _38145_, _38146_);
  or g_48497_(_38144_, _38146_, _38147_);
  or g_48498_(_38120_, _38122_, _38148_);
  or g_48499_(_38134_, _38148_, _38149_);
  or g_48500_(_38147_, _38149_, _38150_);
  or g_48501_(_38142_, _38150_, _38151_);
  or g_48502_(_38127_, _38151_, _38152_);
  xor g_48503_(out[311], out[519], _38153_);
  and g_48504_(_39724_, out[523], _38154_);
  xor g_48505_(out[318], out[526], _38155_);
  xor g_48506_(out[312], out[520], _38156_);
  xor g_48507_(out[305], out[513], _38157_);
  xor g_48508_(out[317], out[525], _38158_);
  xor g_48509_(out[313], out[521], _38159_);
  xor g_48510_(out[308], out[516], _38160_);
  xor g_48511_(out[306], out[514], _38161_);
  and g_48512_(out[315], _39856_, _38162_);
  xor g_48513_(out[307], out[515], _38163_);
  xor g_48514_(out[310], out[518], _38164_);
  xor g_48515_(out[319], out[527], _38165_);
  xor g_48516_(out[314], out[522], _38166_);
  xor g_48517_(out[309], out[517], _38167_);
  xor g_48518_(out[304], out[512], _38168_);
  or g_48519_(_38155_, _38160_, _38169_);
  or g_48520_(_38156_, _38158_, _38170_);
  or g_48521_(_38161_, _38166_, _38171_);
  or g_48522_(_38170_, _38171_, _38172_);
  or g_48523_(_38159_, _38163_, _38173_);
  or g_48524_(_38167_, _38168_, _38174_);
  or g_48525_(_38173_, _38174_, _38175_);
  or g_48526_(_38172_, _38175_, _38176_);
  xor g_48527_(out[316], out[524], _38177_);
  or g_48528_(_38154_, _38177_, _38178_);
  or g_48529_(_38153_, _38164_, _38179_);
  or g_48530_(_38178_, _38179_, _38180_);
  or g_48531_(_38157_, _38162_, _38181_);
  or g_48532_(_38165_, _38181_, _38182_);
  or g_48533_(_38180_, _38182_, _38183_);
  or g_48534_(_38176_, _38183_, _38184_);
  or g_48535_(_38169_, _38184_, _38185_);
  xor g_48536_(out[300], out[524], _38186_);
  and g_48537_(_39702_, out[523], _38187_);
  xor g_48538_(out[301], out[525], _38188_);
  xor g_48539_(out[294], out[518], _38189_);
  xor g_48540_(out[296], out[520], _38190_);
  xor g_48541_(out[297], out[521], _38191_);
  xor g_48542_(out[302], out[526], _38192_);
  xor g_48543_(out[292], out[516], _38193_);
  or g_48544_(_38192_, _38193_, _38194_);
  xor g_48545_(out[293], out[517], _38195_);
  xor g_48546_(out[289], out[513], _38196_);
  and g_48547_(out[299], _39856_, _38197_);
  xor g_48548_(out[303], out[527], _38198_);
  xor g_48549_(out[298], out[522], _38199_);
  xor g_48550_(out[288], out[512], _38200_);
  xor g_48551_(out[290], out[514], _38201_);
  xor g_48552_(out[291], out[515], _38202_);
  or g_48553_(_38188_, _38190_, _38203_);
  or g_48554_(_38199_, _38201_, _38204_);
  or g_48555_(_38203_, _38204_, _38205_);
  or g_48556_(_38191_, _38202_, _38206_);
  or g_48557_(_38195_, _38200_, _38207_);
  or g_48558_(_38206_, _38207_, _38208_);
  or g_48559_(_38205_, _38208_, _38209_);
  or g_48560_(_38186_, _38187_, _38210_);
  xor g_48561_(out[295], out[519], _38211_);
  or g_48562_(_38189_, _38211_, _38212_);
  or g_48563_(_38210_, _38212_, _38213_);
  or g_48564_(_38196_, _38197_, _38214_);
  or g_48565_(_38198_, _38214_, _38215_);
  or g_48566_(_38213_, _38215_, _38216_);
  or g_48567_(_38209_, _38216_, _38217_);
  or g_48568_(_38194_, _38217_, _38218_);
  xor g_48569_(out[279], out[519], _38219_);
  and g_48570_(_39691_, out[523], _38220_);
  xor g_48571_(out[286], out[526], _38221_);
  xor g_48572_(out[280], out[520], _38222_);
  xor g_48573_(out[273], out[513], _38223_);
  xor g_48574_(out[285], out[525], _38224_);
  xor g_48575_(out[281], out[521], _38225_);
  xor g_48576_(out[276], out[516], _38226_);
  xor g_48577_(out[274], out[514], _38227_);
  and g_48578_(out[283], _39856_, _38228_);
  xor g_48579_(out[275], out[515], _38229_);
  xor g_48580_(out[278], out[518], _38230_);
  xor g_48581_(out[287], out[527], _38231_);
  xor g_48582_(out[282], out[522], _38232_);
  xor g_48583_(out[277], out[517], _38233_);
  xor g_48584_(out[272], out[512], _38234_);
  or g_48585_(_38221_, _38226_, _38235_);
  or g_48586_(_38222_, _38224_, _38236_);
  or g_48587_(_38227_, _38232_, _38237_);
  or g_48588_(_38236_, _38237_, _38238_);
  or g_48589_(_38225_, _38229_, _38239_);
  or g_48590_(_38233_, _38234_, _38240_);
  or g_48591_(_38239_, _38240_, _38241_);
  or g_48592_(_38238_, _38241_, _38242_);
  xor g_48593_(out[284], out[524], _38243_);
  or g_48594_(_38220_, _38243_, _38244_);
  or g_48595_(_38219_, _38230_, _38245_);
  or g_48596_(_38244_, _38245_, _38246_);
  or g_48597_(_38223_, _38228_, _38247_);
  or g_48598_(_38231_, _38247_, _38248_);
  or g_48599_(_38246_, _38248_, _38249_);
  or g_48600_(_38242_, _38249_, _38250_);
  or g_48601_(_38235_, _38250_, _38251_);
  xor g_48602_(out[257], out[513], _38252_);
  and g_48603_(_39680_, out[523], _38253_);
  and g_48604_(out[267], _39856_, _38254_);
  xor g_48605_(out[265], out[521], _38255_);
  xor g_48606_(out[256], out[512], _38256_);
  xor g_48607_(out[270], out[526], _38257_);
  xor g_48608_(out[260], out[516], _38258_);
  or g_48609_(_38257_, _38258_, _38259_);
  xor g_48610_(out[269], out[525], _38260_);
  xor g_48611_(out[259], out[515], _38261_);
  xor g_48612_(out[268], out[524], _38262_);
  xor g_48613_(out[262], out[518], _38263_);
  xor g_48614_(out[266], out[522], _38264_);
  xor g_48615_(out[261], out[517], _38265_);
  xor g_48616_(out[271], out[527], _38266_);
  xor g_48617_(out[264], out[520], _38267_);
  or g_48618_(_38260_, _38267_, _38268_);
  xor g_48619_(out[258], out[514], _38269_);
  or g_48620_(_38264_, _38269_, _38270_);
  or g_48621_(_38268_, _38270_, _38271_);
  or g_48622_(_38255_, _38261_, _38272_);
  or g_48623_(_38265_, _38272_, _38273_);
  or g_48624_(_38271_, _38273_, _38274_);
  or g_48625_(_38259_, _38274_, _38275_);
  or g_48626_(_38253_, _38262_, _38276_);
  xor g_48627_(out[263], out[519], _38277_);
  or g_48628_(_38263_, _38277_, _38278_);
  or g_48629_(_38276_, _38278_, _38279_);
  or g_48630_(_38252_, _38254_, _38280_);
  or g_48631_(_38266_, _38280_, _38281_);
  or g_48632_(_38279_, _38281_, _38282_);
  or g_48633_(_38256_, _38282_, _38283_);
  or g_48634_(_38275_, _38283_, _38284_);
  xor g_48635_(out[247], out[519], _38285_);
  and g_48636_(_39669_, out[523], _38286_);
  xor g_48637_(out[254], out[526], _38287_);
  xor g_48638_(out[248], out[520], _38288_);
  xor g_48639_(out[241], out[513], _38289_);
  xor g_48640_(out[253], out[525], _38290_);
  xor g_48641_(out[249], out[521], _38291_);
  xor g_48642_(out[244], out[516], _38292_);
  xor g_48643_(out[242], out[514], _38293_);
  and g_48644_(out[251], _39856_, _38294_);
  xor g_48645_(out[243], out[515], _38295_);
  xor g_48646_(out[246], out[518], _38296_);
  xor g_48647_(out[255], out[527], _38297_);
  xor g_48648_(out[250], out[522], _38298_);
  xor g_48649_(out[245], out[517], _38299_);
  xor g_48650_(out[240], out[512], _38300_);
  or g_48651_(_38287_, _38292_, _38301_);
  or g_48652_(_38288_, _38290_, _38302_);
  or g_48653_(_38293_, _38298_, _38303_);
  or g_48654_(_38302_, _38303_, _38304_);
  or g_48655_(_38291_, _38295_, _38305_);
  or g_48656_(_38299_, _38300_, _38306_);
  or g_48657_(_38305_, _38306_, _38307_);
  or g_48658_(_38304_, _38307_, _38308_);
  xor g_48659_(out[252], out[524], _38309_);
  or g_48660_(_38286_, _38309_, _38310_);
  or g_48661_(_38285_, _38296_, _38311_);
  or g_48662_(_38310_, _38311_, _38312_);
  or g_48663_(_38289_, _38294_, _38313_);
  or g_48664_(_38297_, _38313_, _38314_);
  or g_48665_(_38312_, _38314_, _38315_);
  or g_48666_(_38308_, _38315_, _38316_);
  or g_48667_(_38301_, _38316_, _38317_);
  xor g_48668_(out[226], out[514], _38318_);
  xor g_48669_(out[224], out[512], _38319_);
  xor g_48670_(out[233], out[521], _38320_);
  xor g_48671_(out[232], out[520], _38321_);
  xor g_48672_(out[229], out[517], _38322_);
  xor g_48673_(out[238], out[526], _38323_);
  xor g_48674_(out[237], out[525], _38324_);
  xor g_48675_(out[239], out[527], _38325_);
  xor g_48676_(out[234], out[522], _38326_);
  xor g_48677_(out[230], out[518], _38327_);
  xor g_48678_(out[227], out[515], _38328_);
  and g_48679_(_39658_, out[523], _38329_);
  and g_48680_(out[235], _39856_, _38330_);
  xor g_48681_(out[228], out[516], _38331_);
  xor g_48682_(out[225], out[513], _38332_);
  or g_48683_(_38323_, _38331_, _38333_);
  or g_48684_(_38321_, _38324_, _38334_);
  or g_48685_(_38318_, _38326_, _38335_);
  or g_48686_(_38334_, _38335_, _38336_);
  or g_48687_(_38320_, _38328_, _38337_);
  or g_48688_(_38319_, _38322_, _38338_);
  or g_48689_(_38337_, _38338_, _38339_);
  or g_48690_(_38336_, _38339_, _38340_);
  xor g_48691_(out[236], out[524], _38341_);
  or g_48692_(_38329_, _38341_, _38342_);
  xor g_48693_(out[231], out[519], _38343_);
  or g_48694_(_38327_, _38343_, _38344_);
  or g_48695_(_38342_, _38344_, _38345_);
  or g_48696_(_38330_, _38332_, _38346_);
  or g_48697_(_38325_, _38346_, _38347_);
  or g_48698_(_38345_, _38347_, _38348_);
  or g_48699_(_38340_, _38348_, _38349_);
  or g_48700_(_38333_, _38349_, _38350_);
  xor g_48701_(out[215], out[519], _38351_);
  and g_48702_(_39647_, out[523], _38352_);
  xor g_48703_(out[222], out[526], _38353_);
  xor g_48704_(out[216], out[520], _38354_);
  xor g_48705_(out[209], out[513], _38355_);
  xor g_48706_(out[221], out[525], _38356_);
  xor g_48707_(out[217], out[521], _38357_);
  xor g_48708_(out[212], out[516], _38358_);
  xor g_48709_(out[210], out[514], _38359_);
  and g_48710_(out[219], _39856_, _38360_);
  xor g_48711_(out[211], out[515], _38361_);
  xor g_48712_(out[214], out[518], _38362_);
  xor g_48713_(out[223], out[527], _38363_);
  xor g_48714_(out[218], out[522], _38364_);
  xor g_48715_(out[213], out[517], _38365_);
  xor g_48716_(out[208], out[512], _38366_);
  or g_48717_(_38353_, _38358_, _38367_);
  or g_48718_(_38354_, _38356_, _38368_);
  or g_48719_(_38359_, _38364_, _38369_);
  or g_48720_(_38368_, _38369_, _38370_);
  or g_48721_(_38357_, _38361_, _38371_);
  or g_48722_(_38365_, _38366_, _38372_);
  or g_48723_(_38371_, _38372_, _38373_);
  or g_48724_(_38370_, _38373_, _38374_);
  xor g_48725_(out[220], out[524], _38375_);
  or g_48726_(_38352_, _38375_, _38376_);
  or g_48727_(_38351_, _38362_, _38377_);
  or g_48728_(_38376_, _38377_, _38378_);
  or g_48729_(_38355_, _38360_, _38379_);
  or g_48730_(_38363_, _38379_, _38380_);
  or g_48731_(_38378_, _38380_, _38381_);
  or g_48732_(_38374_, _38381_, _38382_);
  or g_48733_(_38367_, _38382_, _38383_);
  xor g_48734_(out[204], out[524], _38384_);
  and g_48735_(_39636_, out[523], _38385_);
  xor g_48736_(out[200], out[520], _38386_);
  xor g_48737_(out[198], out[518], _38387_);
  xor g_48738_(out[205], out[525], _38388_);
  xor g_48739_(out[206], out[526], _38389_);
  xor g_48740_(out[194], out[514], _38390_);
  xor g_48741_(out[201], out[521], _38391_);
  xor g_48742_(out[197], out[517], _38392_);
  xor g_48743_(out[193], out[513], _38393_);
  and g_48744_(out[203], _39856_, _38394_);
  or g_48745_(_38386_, _38388_, _38395_);
  xor g_48746_(out[207], out[527], _38396_);
  xor g_48747_(out[202], out[522], _38397_);
  xor g_48748_(out[196], out[516], _38398_);
  xor g_48749_(out[195], out[515], _38399_);
  xor g_48750_(out[192], out[512], _38400_);
  or g_48751_(_38390_, _38397_, _38401_);
  or g_48752_(_38395_, _38401_, _38402_);
  or g_48753_(_38391_, _38399_, _38403_);
  or g_48754_(_38392_, _38403_, _38404_);
  or g_48755_(_38402_, _38404_, _38405_);
  or g_48756_(_38389_, _38398_, _38406_);
  or g_48757_(_38405_, _38406_, _38407_);
  or g_48758_(_38384_, _38385_, _38408_);
  xor g_48759_(out[199], out[519], _38409_);
  or g_48760_(_38387_, _38409_, _38410_);
  or g_48761_(_38408_, _38410_, _38411_);
  or g_48762_(_38393_, _38394_, _38412_);
  or g_48763_(_38396_, _38412_, _38413_);
  or g_48764_(_38411_, _38413_, _38414_);
  or g_48765_(_38400_, _38414_, _38415_);
  or g_48766_(_38407_, _38415_, _38416_);
  xor g_48767_(out[183], out[519], _38417_);
  and g_48768_(_39625_, out[523], _38418_);
  xor g_48769_(out[190], out[526], _38419_);
  xor g_48770_(out[184], out[520], _38420_);
  xor g_48771_(out[177], out[513], _38421_);
  xor g_48772_(out[189], out[525], _38422_);
  xor g_48773_(out[185], out[521], _38423_);
  xor g_48774_(out[180], out[516], _38424_);
  xor g_48775_(out[178], out[514], _38425_);
  and g_48776_(out[187], _39856_, _38426_);
  xor g_48777_(out[179], out[515], _38427_);
  xor g_48778_(out[182], out[518], _38428_);
  xor g_48779_(out[191], out[527], _38429_);
  xor g_48780_(out[186], out[522], _38430_);
  xor g_48781_(out[181], out[517], _38431_);
  xor g_48782_(out[176], out[512], _38432_);
  or g_48783_(_38419_, _38424_, _38433_);
  or g_48784_(_38420_, _38422_, _38434_);
  or g_48785_(_38425_, _38430_, _38435_);
  or g_48786_(_38434_, _38435_, _38436_);
  or g_48787_(_38423_, _38427_, _38437_);
  or g_48788_(_38431_, _38432_, _38438_);
  or g_48789_(_38437_, _38438_, _38439_);
  or g_48790_(_38436_, _38439_, _38440_);
  xor g_48791_(out[188], out[524], _38441_);
  or g_48792_(_38418_, _38441_, _38442_);
  or g_48793_(_38417_, _38428_, _38443_);
  or g_48794_(_38442_, _38443_, _38444_);
  or g_48795_(_38421_, _38426_, _38445_);
  or g_48796_(_38429_, _38445_, _38446_);
  or g_48797_(_38444_, _38446_, _38447_);
  or g_48798_(_38440_, _38447_, _38448_);
  or g_48799_(_38433_, _38448_, _38449_);
  not g_48800_(_38449_, _38450_);
  xor g_48801_(out[161], out[513], _38451_);
  and g_48802_(_39614_, out[523], _38452_);
  and g_48803_(out[171], _39856_, _38453_);
  xor g_48804_(out[168], out[520], _38454_);
  xor g_48805_(out[170], out[522], _38455_);
  xor g_48806_(out[162], out[514], _38456_);
  xor g_48807_(out[164], out[516], _38457_);
  xor g_48808_(out[173], out[525], _38458_);
  xor g_48809_(out[169], out[521], _38459_);
  xor g_48810_(out[163], out[515], _38460_);
  xor g_48811_(out[165], out[517], _38461_);
  xor g_48812_(out[174], out[526], _38462_);
  xor g_48813_(out[160], out[512], _38463_);
  xor g_48814_(out[175], out[527], _38464_);
  or g_48815_(_38454_, _38458_, _38465_);
  xor g_48816_(out[166], out[518], _38466_);
  or g_48817_(_38455_, _38456_, _38467_);
  or g_48818_(_38465_, _38467_, _38468_);
  or g_48819_(_38459_, _38460_, _38469_);
  or g_48820_(_38461_, _38469_, _38470_);
  or g_48821_(_38468_, _38470_, _38471_);
  or g_48822_(_38457_, _38462_, _38472_);
  or g_48823_(_38471_, _38472_, _38473_);
  xor g_48824_(out[172], out[524], _38474_);
  or g_48825_(_38452_, _38474_, _38475_);
  xor g_48826_(out[167], out[519], _38476_);
  or g_48827_(_38466_, _38476_, _38477_);
  or g_48828_(_38475_, _38477_, _38478_);
  or g_48829_(_38451_, _38453_, _38479_);
  or g_48830_(_38464_, _38479_, _38480_);
  or g_48831_(_38478_, _38480_, _38481_);
  or g_48832_(_38463_, _38481_, _38482_);
  or g_48833_(_38473_, _38482_, _38483_);
  not g_48834_(_38483_, _38484_);
  xor g_48835_(out[151], out[519], _38485_);
  and g_48836_(_39603_, out[523], _38486_);
  xor g_48837_(out[158], out[526], _38487_);
  xor g_48838_(out[152], out[520], _38488_);
  xor g_48839_(out[145], out[513], _38489_);
  xor g_48840_(out[157], out[525], _38490_);
  xor g_48841_(out[153], out[521], _38491_);
  xor g_48842_(out[148], out[516], _38492_);
  xor g_48843_(out[146], out[514], _38493_);
  and g_48844_(out[155], _39856_, _38494_);
  xor g_48845_(out[147], out[515], _38495_);
  xor g_48846_(out[150], out[518], _38496_);
  xor g_48847_(out[159], out[527], _38497_);
  xor g_48848_(out[154], out[522], _38498_);
  xor g_48849_(out[149], out[517], _38499_);
  xor g_48850_(out[144], out[512], _38500_);
  or g_48851_(_38487_, _38492_, _38501_);
  or g_48852_(_38488_, _38490_, _38502_);
  or g_48853_(_38493_, _38498_, _38503_);
  or g_48854_(_38502_, _38503_, _38504_);
  or g_48855_(_38491_, _38495_, _38505_);
  or g_48856_(_38499_, _38500_, _38506_);
  or g_48857_(_38505_, _38506_, _38507_);
  or g_48858_(_38504_, _38507_, _38508_);
  xor g_48859_(out[156], out[524], _38509_);
  or g_48860_(_38486_, _38509_, _38510_);
  or g_48861_(_38485_, _38496_, _38511_);
  or g_48862_(_38510_, _38511_, _38512_);
  or g_48863_(_38489_, _38494_, _38513_);
  or g_48864_(_38497_, _38513_, _38514_);
  or g_48865_(_38512_, _38514_, _38515_);
  or g_48866_(_38508_, _38515_, _38516_);
  or g_48867_(_38501_, _38516_, _38517_);
  and g_48868_(out[139], _39856_, _38518_);
  xor g_48869_(out[132], out[516], _38519_);
  xor g_48870_(out[142], out[526], _38520_);
  or g_48871_(_38519_, _38520_, _38521_);
  xor g_48872_(out[141], out[525], _38522_);
  xor g_48873_(out[131], out[515], _38523_);
  xor g_48874_(out[128], out[512], _38524_);
  and g_48875_(_39592_, out[523], _38525_);
  xor g_48876_(out[138], out[522], _38526_);
  xor g_48877_(out[143], out[527], _38527_);
  xor g_48878_(out[134], out[518], _38528_);
  xor g_48879_(out[133], out[517], _38529_);
  xor g_48880_(out[136], out[520], _38530_);
  or g_48881_(_38522_, _38530_, _38531_);
  xor g_48882_(out[130], out[514], _38532_);
  xor g_48883_(out[137], out[521], _38533_);
  xor g_48884_(out[129], out[513], _38534_);
  or g_48885_(_38526_, _38532_, _38535_);
  or g_48886_(_38531_, _38535_, _38536_);
  or g_48887_(_38523_, _38533_, _38537_);
  or g_48888_(_38529_, _38537_, _38538_);
  or g_48889_(_38536_, _38538_, _38539_);
  or g_48890_(_38521_, _38539_, _38540_);
  xor g_48891_(out[140], out[524], _38541_);
  or g_48892_(_38525_, _38541_, _38542_);
  xor g_48893_(out[135], out[519], _38543_);
  or g_48894_(_38528_, _38543_, _38544_);
  or g_48895_(_38542_, _38544_, _38545_);
  or g_48896_(_38518_, _38534_, _38546_);
  or g_48897_(_38527_, _38546_, _38547_);
  or g_48898_(_38545_, _38547_, _38548_);
  or g_48899_(_38524_, _38548_, _38549_);
  or g_48900_(_38540_, _38549_, _38550_);
  xor g_48901_(out[119], out[519], _38551_);
  and g_48902_(_39581_, out[523], _38552_);
  xor g_48903_(out[126], out[526], _38553_);
  xor g_48904_(out[120], out[520], _38554_);
  xor g_48905_(out[113], out[513], _38555_);
  xor g_48906_(out[125], out[525], _38556_);
  xor g_48907_(out[121], out[521], _38557_);
  xor g_48908_(out[116], out[516], _38558_);
  xor g_48909_(out[114], out[514], _38559_);
  and g_48910_(out[123], _39856_, _38560_);
  xor g_48911_(out[115], out[515], _38561_);
  xor g_48912_(out[118], out[518], _38562_);
  xor g_48913_(out[127], out[527], _38563_);
  xor g_48914_(out[122], out[522], _38564_);
  xor g_48915_(out[117], out[517], _38565_);
  xor g_48916_(out[112], out[512], _38566_);
  or g_48917_(_38553_, _38558_, _38567_);
  or g_48918_(_38554_, _38556_, _38568_);
  or g_48919_(_38559_, _38564_, _38569_);
  or g_48920_(_38568_, _38569_, _38570_);
  or g_48921_(_38557_, _38561_, _38571_);
  or g_48922_(_38565_, _38566_, _38572_);
  or g_48923_(_38571_, _38572_, _38573_);
  or g_48924_(_38570_, _38573_, _38574_);
  xor g_48925_(out[124], out[524], _38575_);
  or g_48926_(_38552_, _38575_, _38576_);
  or g_48927_(_38551_, _38562_, _38577_);
  or g_48928_(_38576_, _38577_, _38578_);
  or g_48929_(_38555_, _38560_, _38579_);
  or g_48930_(_38563_, _38579_, _38580_);
  or g_48931_(_38578_, _38580_, _38581_);
  or g_48932_(_38574_, _38581_, _38582_);
  or g_48933_(_38567_, _38582_, _38583_);
  xor g_48934_(out[109], out[525], _38584_);
  xor g_48935_(out[98], out[514], _38585_);
  xor g_48936_(out[101], out[517], _38586_);
  xor g_48937_(out[105], out[521], _38587_);
  xor g_48938_(out[100], out[516], _38588_);
  xor g_48939_(out[104], out[520], _38589_);
  xor g_48940_(out[110], out[526], _38590_);
  xor g_48941_(out[102], out[518], _38591_);
  xor g_48942_(out[111], out[527], _38592_);
  xor g_48943_(out[106], out[522], _38593_);
  xor g_48944_(out[96], out[512], _38594_);
  xor g_48945_(out[99], out[515], _38595_);
  and g_48946_(_39570_, out[523], _38596_);
  and g_48947_(out[107], _39856_, _38597_);
  xor g_48948_(out[97], out[513], _38598_);
  or g_48949_(_38588_, _38590_, _38599_);
  or g_48950_(_38584_, _38589_, _38600_);
  or g_48951_(_38585_, _38593_, _38601_);
  or g_48952_(_38600_, _38601_, _38602_);
  or g_48953_(_38587_, _38595_, _38603_);
  or g_48954_(_38586_, _38594_, _38604_);
  or g_48955_(_38603_, _38604_, _38605_);
  or g_48956_(_38602_, _38605_, _38606_);
  xor g_48957_(out[108], out[524], _38607_);
  or g_48958_(_38596_, _38607_, _38608_);
  xor g_48959_(out[103], out[519], _38609_);
  or g_48960_(_38591_, _38609_, _38610_);
  or g_48961_(_38608_, _38610_, _38611_);
  or g_48962_(_38597_, _38598_, _38612_);
  or g_48963_(_38592_, _38612_, _38613_);
  or g_48964_(_38611_, _38613_, _38614_);
  or g_48965_(_38606_, _38614_, _38615_);
  or g_48966_(_38599_, _38615_, _38616_);
  not g_48967_(_38616_, _38617_);
  xor g_48968_(out[87], out[519], _38618_);
  and g_48969_(_39559_, out[523], _38619_);
  xor g_48970_(out[94], out[526], _38620_);
  xor g_48971_(out[88], out[520], _38621_);
  xor g_48972_(out[81], out[513], _38622_);
  xor g_48973_(out[93], out[525], _38623_);
  xor g_48974_(out[89], out[521], _38624_);
  xor g_48975_(out[84], out[516], _38625_);
  xor g_48976_(out[82], out[514], _38626_);
  and g_48977_(out[91], _39856_, _38627_);
  xor g_48978_(out[83], out[515], _38628_);
  xor g_48979_(out[86], out[518], _38629_);
  xor g_48980_(out[95], out[527], _38630_);
  xor g_48981_(out[90], out[522], _38631_);
  xor g_48982_(out[85], out[517], _38632_);
  xor g_48983_(out[80], out[512], _38633_);
  or g_48984_(_38620_, _38625_, _38634_);
  or g_48985_(_38621_, _38623_, _38635_);
  or g_48986_(_38626_, _38631_, _38636_);
  or g_48987_(_38635_, _38636_, _38637_);
  or g_48988_(_38624_, _38628_, _38638_);
  or g_48989_(_38632_, _38633_, _38639_);
  or g_48990_(_38638_, _38639_, _38640_);
  or g_48991_(_38637_, _38640_, _38641_);
  xor g_48992_(out[92], out[524], _38642_);
  or g_48993_(_38619_, _38642_, _38643_);
  or g_48994_(_38618_, _38629_, _38644_);
  or g_48995_(_38643_, _38644_, _38645_);
  or g_48996_(_38622_, _38627_, _38646_);
  or g_48997_(_38630_, _38646_, _38647_);
  or g_48998_(_38645_, _38647_, _38648_);
  or g_48999_(_38641_, _38648_, _38649_);
  or g_49000_(_38634_, _38649_, _38650_);
  not g_49001_(_38650_, _38651_);
  xor g_49002_(out[77], out[525], _38652_);
  xor g_49003_(out[74], out[522], _38653_);
  xor g_49004_(out[69], out[517], _38654_);
  and g_49005_(_39548_, out[523], _38655_);
  xor g_49006_(out[64], out[512], _38656_);
  and g_49007_(out[75], _39856_, _38657_);
  xor g_49008_(out[66], out[514], _38658_);
  xor g_49009_(out[67], out[515], _38659_);
  xor g_49010_(out[73], out[521], _38660_);
  xor g_49011_(out[65], out[513], _38661_);
  xor g_49012_(out[79], out[527], _38662_);
  xor g_49013_(out[78], out[526], _38663_);
  xor g_49014_(out[70], out[518], _38664_);
  xor g_49015_(out[68], out[516], _38665_);
  xor g_49016_(out[72], out[520], _38666_);
  or g_49017_(_38652_, _38666_, _38667_);
  or g_49018_(_38653_, _38658_, _38668_);
  or g_49019_(_38667_, _38668_, _38669_);
  or g_49020_(_38659_, _38660_, _38670_);
  or g_49021_(_38654_, _38670_, _38671_);
  or g_49022_(_38669_, _38671_, _38672_);
  or g_49023_(_38663_, _38665_, _38673_);
  or g_49024_(_38672_, _38673_, _38674_);
  xor g_49025_(out[76], out[524], _38675_);
  or g_49026_(_38655_, _38675_, _38676_);
  xor g_49027_(out[71], out[519], _38677_);
  or g_49028_(_38664_, _38677_, _38678_);
  or g_49029_(_38676_, _38678_, _38679_);
  or g_49030_(_38657_, _38661_, _38680_);
  or g_49031_(_38662_, _38680_, _38681_);
  or g_49032_(_38679_, _38681_, _38682_);
  or g_49033_(_38656_, _38682_, _38683_);
  or g_49034_(_38674_, _38683_, _38684_);
  xor g_49035_(out[55], out[519], _38685_);
  and g_49036_(_39537_, out[523], _38686_);
  xor g_49037_(out[62], out[526], _38687_);
  xor g_49038_(out[56], out[520], _38688_);
  xor g_49039_(out[49], out[513], _38689_);
  xor g_49040_(out[61], out[525], _38690_);
  xor g_49041_(out[57], out[521], _38691_);
  xor g_49042_(out[52], out[516], _38692_);
  xor g_49043_(out[50], out[514], _38693_);
  and g_49044_(out[59], _39856_, _38694_);
  xor g_49045_(out[51], out[515], _38695_);
  xor g_49046_(out[54], out[518], _38696_);
  xor g_49047_(out[63], out[527], _38697_);
  xor g_49048_(out[58], out[522], _38698_);
  xor g_49049_(out[53], out[517], _38699_);
  xor g_49050_(out[48], out[512], _38700_);
  or g_49051_(_38687_, _38692_, _38701_);
  or g_49052_(_38688_, _38690_, _38702_);
  or g_49053_(_38693_, _38698_, _38703_);
  or g_49054_(_38702_, _38703_, _38704_);
  or g_49055_(_38691_, _38695_, _38705_);
  or g_49056_(_38699_, _38700_, _38706_);
  or g_49057_(_38705_, _38706_, _38707_);
  or g_49058_(_38704_, _38707_, _38708_);
  xor g_49059_(out[60], out[524], _38709_);
  or g_49060_(_38686_, _38709_, _38710_);
  or g_49061_(_38685_, _38696_, _38711_);
  or g_49062_(_38710_, _38711_, _38712_);
  or g_49063_(_38689_, _38694_, _38713_);
  or g_49064_(_38697_, _38713_, _38714_);
  or g_49065_(_38712_, _38714_, _38715_);
  or g_49066_(_38708_, _38715_, _38716_);
  or g_49067_(_38701_, _38716_, _38717_);
  xor g_49068_(out[33], out[513], _38718_);
  and g_49069_(out[43], _39856_, _38719_);
  xor g_49070_(out[41], out[521], _38720_);
  xor g_49071_(out[32], out[512], _38721_);
  xor g_49072_(out[46], out[526], _38722_);
  xor g_49073_(out[36], out[516], _38723_);
  or g_49074_(_38722_, _38723_, _38724_);
  xor g_49075_(out[45], out[525], _38725_);
  xor g_49076_(out[35], out[515], _38726_);
  and g_49077_(_39526_, out[523], _38727_);
  xor g_49078_(out[38], out[518], _38728_);
  xor g_49079_(out[42], out[522], _38729_);
  xor g_49080_(out[37], out[517], _38730_);
  xor g_49081_(out[47], out[527], _38731_);
  xor g_49082_(out[40], out[520], _38732_);
  or g_49083_(_38725_, _38732_, _38733_);
  xor g_49084_(out[34], out[514], _38734_);
  or g_49085_(_38729_, _38734_, _38735_);
  or g_49086_(_38733_, _38735_, _38736_);
  or g_49087_(_38720_, _38726_, _38737_);
  or g_49088_(_38730_, _38737_, _38738_);
  or g_49089_(_38736_, _38738_, _38739_);
  or g_49090_(_38724_, _38739_, _38740_);
  xor g_49091_(out[44], out[524], _38741_);
  or g_49092_(_38727_, _38741_, _38742_);
  xor g_49093_(out[39], out[519], _38743_);
  or g_49094_(_38728_, _38743_, _38744_);
  or g_49095_(_38742_, _38744_, _38745_);
  or g_49096_(_38718_, _38719_, _38746_);
  or g_49097_(_38731_, _38746_, _38747_);
  or g_49098_(_38745_, _38747_, _38748_);
  or g_49099_(_38721_, _38748_, _38749_);
  or g_49100_(_38740_, _38749_, _38750_);
  xor g_49101_(out[23], out[519], _38751_);
  and g_49102_(_39493_, out[523], _38752_);
  xor g_49103_(out[30], out[526], _38753_);
  xor g_49104_(out[24], out[520], _38754_);
  xor g_49105_(out[17], out[513], _38755_);
  xor g_49106_(out[29], out[525], _38756_);
  xor g_49107_(out[25], out[521], _38757_);
  xor g_49108_(out[20], out[516], _38758_);
  xor g_49109_(out[18], out[514], _38759_);
  and g_49110_(out[27], _39856_, _38760_);
  xor g_49111_(out[19], out[515], _38761_);
  xor g_49112_(out[22], out[518], _38762_);
  xor g_49113_(out[31], out[527], _38763_);
  xor g_49114_(out[26], out[522], _38764_);
  xor g_49115_(out[21], out[517], _38765_);
  xor g_49116_(out[16], out[512], _38766_);
  or g_49117_(_38753_, _38758_, _38767_);
  or g_49118_(_38754_, _38756_, _38768_);
  or g_49119_(_38759_, _38764_, _38769_);
  or g_49120_(_38768_, _38769_, _38770_);
  or g_49121_(_38757_, _38761_, _38771_);
  or g_49122_(_38765_, _38766_, _38772_);
  or g_49123_(_38771_, _38772_, _38773_);
  or g_49124_(_38770_, _38773_, _38774_);
  xor g_49125_(out[28], out[524], _38775_);
  or g_49126_(_38752_, _38775_, _38776_);
  or g_49127_(_38751_, _38762_, _38777_);
  or g_49128_(_38776_, _38777_, _38778_);
  or g_49129_(_38755_, _38760_, _38779_);
  or g_49130_(_38763_, _38779_, _38780_);
  or g_49131_(_38778_, _38780_, _38781_);
  or g_49132_(_38774_, _38781_, _38782_);
  or g_49133_(_38767_, _38782_, _38783_);
  xor g_49134_(out[10], out[522], _38784_);
  xor g_49135_(out[2], out[514], _38785_);
  xor g_49136_(out[1], out[513], _38786_);
  and g_49137_(_39438_, out[523], _38787_);
  and g_49138_(out[11], _39856_, _38788_);
  xor g_49139_(out[13], out[525], _38789_);
  xor g_49140_(out[3], out[515], _38790_);
  xor g_49141_(out[14], out[526], _38791_);
  xor g_49142_(out[12], out[524], _38792_);
  xor g_49143_(out[8], out[520], _38793_);
  xor g_49144_(out[15], out[527], _38794_);
  xor g_49145_(out[5], out[517], _38795_);
  xor g_49146_(out[6], out[518], _38796_);
  xor g_49147_(out[0], out[512], _38797_);
  xor g_49148_(out[4], out[516], _38798_);
  or g_49149_(_38789_, _38793_, _38799_);
  xor g_49150_(out[9], out[521], _38800_);
  or g_49151_(_38784_, _38785_, _38801_);
  or g_49152_(_38799_, _38801_, _38802_);
  or g_49153_(_38790_, _38800_, _38803_);
  or g_49154_(_38795_, _38803_, _38804_);
  or g_49155_(_38802_, _38804_, _38805_);
  or g_49156_(_38791_, _38798_, _38806_);
  or g_49157_(_38805_, _38806_, _38807_);
  or g_49158_(_38787_, _38792_, _38808_);
  xor g_49159_(out[7], out[519], _38809_);
  or g_49160_(_38796_, _38809_, _38810_);
  or g_49161_(_38808_, _38810_, _38811_);
  or g_49162_(_38786_, _38788_, _38812_);
  or g_49163_(_38794_, _38812_, _38813_);
  or g_49164_(_38811_, _38813_, _38814_);
  or g_49165_(_38797_, _38814_, _38815_);
  or g_49166_(_38807_, _38815_, _38816_);
  not g_49167_(_38816_, _38817_);
  xor g_49168_(out[305], out[497], _38818_);
  and g_49169_(out[315], _39845_, _38819_);
  xor g_49170_(out[313], out[505], _38820_);
  xor g_49171_(out[304], out[496], _38821_);
  xor g_49172_(out[318], out[510], _38822_);
  xor g_49173_(out[308], out[500], _38823_);
  or g_49174_(_38822_, _38823_, _38824_);
  xor g_49175_(out[317], out[509], _38825_);
  xor g_49176_(out[307], out[499], _38826_);
  and g_49177_(_39724_, out[507], _38827_);
  xor g_49178_(out[310], out[502], _38828_);
  xor g_49179_(out[314], out[506], _38829_);
  xor g_49180_(out[309], out[501], _38830_);
  xor g_49181_(out[319], out[511], _38831_);
  xor g_49182_(out[312], out[504], _38832_);
  or g_49183_(_38825_, _38832_, _38833_);
  xor g_49184_(out[306], out[498], _38834_);
  or g_49185_(_38829_, _38834_, _38835_);
  or g_49186_(_38833_, _38835_, _38836_);
  or g_49187_(_38820_, _38826_, _38837_);
  or g_49188_(_38830_, _38837_, _38838_);
  or g_49189_(_38836_, _38838_, _38839_);
  or g_49190_(_38824_, _38839_, _38840_);
  xor g_49191_(out[316], out[508], _38841_);
  or g_49192_(_38827_, _38841_, _38842_);
  xor g_49193_(out[311], out[503], _38843_);
  or g_49194_(_38828_, _38843_, _38844_);
  or g_49195_(_38842_, _38844_, _38845_);
  or g_49196_(_38818_, _38819_, _38846_);
  or g_49197_(_38831_, _38846_, _38847_);
  or g_49198_(_38845_, _38847_, _38848_);
  or g_49199_(_38821_, _38848_, _38849_);
  or g_49200_(_38840_, _38849_, _38850_);
  xor g_49201_(out[295], out[503], _38851_);
  and g_49202_(_39702_, out[507], _38852_);
  xor g_49203_(out[302], out[510], _38853_);
  xor g_49204_(out[296], out[504], _38854_);
  xor g_49205_(out[289], out[497], _38855_);
  xor g_49206_(out[301], out[509], _38856_);
  xor g_49207_(out[297], out[505], _38857_);
  xor g_49208_(out[292], out[500], _38858_);
  xor g_49209_(out[290], out[498], _38859_);
  and g_49210_(out[299], _39845_, _38860_);
  xor g_49211_(out[291], out[499], _38861_);
  xor g_49212_(out[294], out[502], _38862_);
  xor g_49213_(out[303], out[511], _38863_);
  xor g_49214_(out[298], out[506], _38864_);
  xor g_49215_(out[293], out[501], _38865_);
  xor g_49216_(out[288], out[496], _38866_);
  or g_49217_(_38853_, _38858_, _38867_);
  or g_49218_(_38854_, _38856_, _38868_);
  or g_49219_(_38859_, _38864_, _38869_);
  or g_49220_(_38868_, _38869_, _38870_);
  or g_49221_(_38857_, _38861_, _38871_);
  or g_49222_(_38865_, _38866_, _38872_);
  or g_49223_(_38871_, _38872_, _38873_);
  or g_49224_(_38870_, _38873_, _38874_);
  xor g_49225_(out[300], out[508], _38875_);
  or g_49226_(_38852_, _38875_, _38876_);
  or g_49227_(_38851_, _38862_, _38877_);
  or g_49228_(_38876_, _38877_, _38878_);
  or g_49229_(_38855_, _38860_, _38879_);
  or g_49230_(_38863_, _38879_, _38880_);
  or g_49231_(_38878_, _38880_, _38881_);
  or g_49232_(_38874_, _38881_, _38882_);
  or g_49233_(_38867_, _38882_, _38883_);
  xor g_49234_(out[273], out[497], _38884_);
  and g_49235_(out[283], _39845_, _38885_);
  xor g_49236_(out[286], out[510], _38886_);
  xor g_49237_(out[275], out[499], _38887_);
  xor g_49238_(out[276], out[500], _38888_);
  xor g_49239_(out[274], out[498], _38889_);
  xor g_49240_(out[281], out[505], _38890_);
  xor g_49241_(out[272], out[496], _38891_);
  and g_49242_(_39691_, out[507], _38892_);
  xor g_49243_(out[278], out[502], _38893_);
  xor g_49244_(out[282], out[506], _38894_);
  xor g_49245_(out[277], out[501], _38895_);
  xor g_49246_(out[287], out[511], _38896_);
  xor g_49247_(out[285], out[509], _38897_);
  xor g_49248_(out[280], out[504], _38898_);
  or g_49249_(_38886_, _38888_, _38899_);
  or g_49250_(_38897_, _38898_, _38900_);
  or g_49251_(_38889_, _38894_, _38901_);
  or g_49252_(_38900_, _38901_, _38902_);
  or g_49253_(_38887_, _38890_, _38903_);
  or g_49254_(_38891_, _38895_, _38904_);
  or g_49255_(_38903_, _38904_, _38905_);
  or g_49256_(_38902_, _38905_, _38906_);
  xor g_49257_(out[284], out[508], _38907_);
  or g_49258_(_38892_, _38907_, _38908_);
  xor g_49259_(out[279], out[503], _38909_);
  or g_49260_(_38893_, _38909_, _38910_);
  or g_49261_(_38908_, _38910_, _38911_);
  or g_49262_(_38884_, _38885_, _38912_);
  or g_49263_(_38896_, _38912_, _38913_);
  or g_49264_(_38911_, _38913_, _38914_);
  or g_49265_(_38906_, _38914_, _38915_);
  or g_49266_(_38899_, _38915_, _38916_);
  not g_49267_(_38916_, _38917_);
  xor g_49268_(out[263], out[503], _38918_);
  and g_49269_(_39680_, out[507], _38919_);
  xor g_49270_(out[270], out[510], _38920_);
  xor g_49271_(out[264], out[504], _38921_);
  xor g_49272_(out[257], out[497], _38922_);
  xor g_49273_(out[269], out[509], _38923_);
  xor g_49274_(out[265], out[505], _38924_);
  xor g_49275_(out[260], out[500], _38925_);
  xor g_49276_(out[258], out[498], _38926_);
  and g_49277_(out[267], _39845_, _38927_);
  xor g_49278_(out[259], out[499], _38928_);
  xor g_49279_(out[262], out[502], _38929_);
  xor g_49280_(out[271], out[511], _38930_);
  xor g_49281_(out[266], out[506], _38931_);
  xor g_49282_(out[261], out[501], _38932_);
  xor g_49283_(out[256], out[496], _38933_);
  or g_49284_(_38920_, _38925_, _38934_);
  or g_49285_(_38921_, _38923_, _38935_);
  or g_49286_(_38926_, _38931_, _38936_);
  or g_49287_(_38935_, _38936_, _38937_);
  or g_49288_(_38924_, _38928_, _38938_);
  or g_49289_(_38932_, _38933_, _38939_);
  or g_49290_(_38938_, _38939_, _38940_);
  or g_49291_(_38937_, _38940_, _38941_);
  xor g_49292_(out[268], out[508], _38942_);
  or g_49293_(_38919_, _38942_, _38943_);
  or g_49294_(_38918_, _38929_, _38944_);
  or g_49295_(_38943_, _38944_, _38945_);
  or g_49296_(_38922_, _38927_, _38946_);
  or g_49297_(_38930_, _38946_, _38947_);
  or g_49298_(_38945_, _38947_, _38948_);
  or g_49299_(_38941_, _38948_, _38949_);
  or g_49300_(_38934_, _38949_, _38950_);
  xor g_49301_(out[248], out[504], _38951_);
  xor g_49302_(out[245], out[501], _38952_);
  xor g_49303_(out[243], out[499], _38953_);
  xor g_49304_(out[254], out[510], _38954_);
  xor g_49305_(out[253], out[509], _38955_);
  xor g_49306_(out[242], out[498], _38956_);
  xor g_49307_(out[249], out[505], _38957_);
  xor g_49308_(out[246], out[502], _38958_);
  xor g_49309_(out[255], out[511], _38959_);
  xor g_49310_(out[250], out[506], _38960_);
  xor g_49311_(out[244], out[500], _38961_);
  xor g_49312_(out[240], out[496], _38962_);
  and g_49313_(_39669_, out[507], _38963_);
  and g_49314_(out[251], _39845_, _38964_);
  or g_49315_(_38951_, _38955_, _38965_);
  xor g_49316_(out[241], out[497], _38966_);
  or g_49317_(_38956_, _38960_, _38967_);
  or g_49318_(_38965_, _38967_, _38968_);
  or g_49319_(_38953_, _38957_, _38969_);
  or g_49320_(_38952_, _38969_, _38970_);
  or g_49321_(_38968_, _38970_, _38971_);
  or g_49322_(_38954_, _38961_, _38972_);
  or g_49323_(_38971_, _38972_, _38973_);
  xor g_49324_(out[252], out[508], _38974_);
  or g_49325_(_38963_, _38974_, _38975_);
  xor g_49326_(out[247], out[503], _38976_);
  or g_49327_(_38958_, _38976_, _38977_);
  or g_49328_(_38975_, _38977_, _38978_);
  or g_49329_(_38964_, _38966_, _38979_);
  or g_49330_(_38959_, _38979_, _38980_);
  or g_49331_(_38978_, _38980_, _38981_);
  or g_49332_(_38962_, _38981_, _38982_);
  or g_49333_(_38973_, _38982_, _38983_);
  not g_49334_(_38983_, _38984_);
  xor g_49335_(out[231], out[503], _38985_);
  and g_49336_(_39658_, out[507], _38986_);
  xor g_49337_(out[238], out[510], _38987_);
  xor g_49338_(out[232], out[504], _38988_);
  xor g_49339_(out[225], out[497], _38989_);
  xor g_49340_(out[237], out[509], _38990_);
  xor g_49341_(out[233], out[505], _38991_);
  xor g_49342_(out[228], out[500], _38992_);
  xor g_49343_(out[226], out[498], _38993_);
  and g_49344_(out[235], _39845_, _38994_);
  xor g_49345_(out[227], out[499], _38995_);
  xor g_49346_(out[230], out[502], _38996_);
  xor g_49347_(out[239], out[511], _38997_);
  xor g_49348_(out[234], out[506], _38998_);
  xor g_49349_(out[229], out[501], _38999_);
  xor g_49350_(out[224], out[496], _39000_);
  or g_49351_(_38987_, _38992_, _39001_);
  or g_49352_(_38988_, _38990_, _39002_);
  or g_49353_(_38993_, _38998_, _39003_);
  or g_49354_(_39002_, _39003_, _39004_);
  or g_49355_(_38991_, _38995_, _39005_);
  or g_49356_(_38999_, _39000_, _39006_);
  or g_49357_(_39005_, _39006_, _39007_);
  or g_49358_(_39004_, _39007_, _39008_);
  xor g_49359_(out[236], out[508], _39009_);
  or g_49360_(_38986_, _39009_, _39010_);
  or g_49361_(_38985_, _38996_, _39011_);
  or g_49362_(_39010_, _39011_, _39012_);
  or g_49363_(_38989_, _38994_, _39013_);
  or g_49364_(_38997_, _39013_, _39014_);
  or g_49365_(_39012_, _39014_, _39015_);
  or g_49366_(_39008_, _39015_, _39016_);
  or g_49367_(_39001_, _39016_, _39017_);
  xor g_49368_(out[209], out[497], _39018_);
  and g_49369_(out[219], _39845_, _39019_);
  xor g_49370_(out[217], out[505], _39020_);
  xor g_49371_(out[208], out[496], _39021_);
  xor g_49372_(out[222], out[510], _39022_);
  xor g_49373_(out[212], out[500], _39023_);
  or g_49374_(_39022_, _39023_, _39024_);
  xor g_49375_(out[221], out[509], _39025_);
  xor g_49376_(out[211], out[499], _39026_);
  and g_49377_(_39647_, out[507], _39027_);
  xor g_49378_(out[214], out[502], _39028_);
  xor g_49379_(out[218], out[506], _39029_);
  xor g_49380_(out[213], out[501], _39030_);
  xor g_49381_(out[223], out[511], _39031_);
  xor g_49382_(out[216], out[504], _39032_);
  or g_49383_(_39025_, _39032_, _39033_);
  xor g_49384_(out[210], out[498], _39034_);
  or g_49385_(_39029_, _39034_, _39035_);
  or g_49386_(_39033_, _39035_, _39036_);
  or g_49387_(_39020_, _39026_, _39037_);
  or g_49388_(_39030_, _39037_, _39038_);
  or g_49389_(_39036_, _39038_, _39039_);
  or g_49390_(_39024_, _39039_, _39040_);
  xor g_49391_(out[220], out[508], _39041_);
  or g_49392_(_39027_, _39041_, _39042_);
  xor g_49393_(out[215], out[503], _39043_);
  or g_49394_(_39028_, _39043_, _39044_);
  or g_49395_(_39042_, _39044_, _39045_);
  or g_49396_(_39018_, _39019_, _39046_);
  or g_49397_(_39031_, _39046_, _39047_);
  or g_49398_(_39045_, _39047_, _39048_);
  or g_49399_(_39021_, _39048_, _39049_);
  or g_49400_(_39040_, _39049_, _39050_);
  xor g_49401_(out[199], out[503], _39051_);
  and g_49402_(_39636_, out[507], _39052_);
  xor g_49403_(out[206], out[510], _39053_);
  xor g_49404_(out[200], out[504], _39054_);
  xor g_49405_(out[193], out[497], _39055_);
  xor g_49406_(out[205], out[509], _39056_);
  xor g_49407_(out[201], out[505], _39057_);
  xor g_49408_(out[196], out[500], _39058_);
  xor g_49409_(out[194], out[498], _39059_);
  and g_49410_(out[203], _39845_, _39060_);
  xor g_49411_(out[195], out[499], _39061_);
  xor g_49412_(out[198], out[502], _39062_);
  xor g_49413_(out[207], out[511], _39063_);
  xor g_49414_(out[202], out[506], _39064_);
  xor g_49415_(out[197], out[501], _39065_);
  xor g_49416_(out[192], out[496], _39066_);
  or g_49417_(_39053_, _39058_, _39067_);
  or g_49418_(_39054_, _39056_, _39068_);
  or g_49419_(_39059_, _39064_, _39069_);
  or g_49420_(_39068_, _39069_, _39070_);
  or g_49421_(_39057_, _39061_, _39071_);
  or g_49422_(_39065_, _39066_, _39072_);
  or g_49423_(_39071_, _39072_, _39073_);
  or g_49424_(_39070_, _39073_, _39074_);
  xor g_49425_(out[204], out[508], _39075_);
  or g_49426_(_39052_, _39075_, _39076_);
  or g_49427_(_39051_, _39062_, _39077_);
  or g_49428_(_39076_, _39077_, _39078_);
  or g_49429_(_39055_, _39060_, _39079_);
  or g_49430_(_39063_, _39079_, _39080_);
  or g_49431_(_39078_, _39080_, _39081_);
  or g_49432_(_39074_, _39081_, _39082_);
  or g_49433_(_39067_, _39082_, _39083_);
  not g_49434_(_39083_, _39084_);
  xor g_49435_(out[184], out[504], _39085_);
  xor g_49436_(out[181], out[501], _39086_);
  xor g_49437_(out[179], out[499], _39087_);
  xor g_49438_(out[190], out[510], _39088_);
  xor g_49439_(out[189], out[509], _39089_);
  xor g_49440_(out[178], out[498], _39090_);
  xor g_49441_(out[185], out[505], _39091_);
  xor g_49442_(out[182], out[502], _39092_);
  xor g_49443_(out[191], out[511], _39093_);
  xor g_49444_(out[186], out[506], _39094_);
  xor g_49445_(out[180], out[500], _39095_);
  xor g_49446_(out[176], out[496], _39096_);
  and g_49447_(_39625_, out[507], _39097_);
  and g_49448_(out[187], _39845_, _39098_);
  or g_49449_(_39085_, _39089_, _39099_);
  xor g_49450_(out[177], out[497], _39100_);
  or g_49451_(_39090_, _39094_, _39101_);
  or g_49452_(_39099_, _39101_, _39102_);
  or g_49453_(_39087_, _39091_, _39103_);
  or g_49454_(_39086_, _39103_, _39104_);
  or g_49455_(_39102_, _39104_, _39105_);
  or g_49456_(_39088_, _39095_, _39106_);
  or g_49457_(_39105_, _39106_, _39107_);
  xor g_49458_(out[188], out[508], _39108_);
  or g_49459_(_39097_, _39108_, _39109_);
  xor g_49460_(out[183], out[503], _39110_);
  or g_49461_(_39092_, _39110_, _39111_);
  or g_49462_(_39109_, _39111_, _39112_);
  or g_49463_(_39098_, _39100_, _39113_);
  or g_49464_(_39093_, _39113_, _39114_);
  or g_49465_(_39112_, _39114_, _39115_);
  or g_49466_(_39096_, _39115_, _39116_);
  or g_49467_(_39107_, _39116_, _39117_);
  not g_49468_(_39117_, _39118_);
  xor g_49469_(out[167], out[503], _39119_);
  and g_49470_(_39614_, out[507], _39120_);
  xor g_49471_(out[174], out[510], _39121_);
  xor g_49472_(out[168], out[504], _39122_);
  xor g_49473_(out[161], out[497], _39123_);
  xor g_49474_(out[173], out[509], _39124_);
  xor g_49475_(out[169], out[505], _39125_);
  xor g_49476_(out[164], out[500], _39126_);
  xor g_49477_(out[162], out[498], _39127_);
  and g_49478_(out[171], _39845_, _39128_);
  xor g_49479_(out[163], out[499], _39129_);
  xor g_49480_(out[166], out[502], _39130_);
  xor g_49481_(out[175], out[511], _39131_);
  xor g_49482_(out[170], out[506], _39132_);
  xor g_49483_(out[165], out[501], _39133_);
  xor g_49484_(out[160], out[496], _39134_);
  or g_49485_(_39121_, _39126_, _39135_);
  or g_49486_(_39122_, _39124_, _39136_);
  or g_49487_(_39127_, _39132_, _39137_);
  or g_49488_(_39136_, _39137_, _39138_);
  or g_49489_(_39125_, _39129_, _39139_);
  or g_49490_(_39133_, _39134_, _39140_);
  or g_49491_(_39139_, _39140_, _39141_);
  or g_49492_(_39138_, _39141_, _39142_);
  xor g_49493_(out[172], out[508], _39143_);
  or g_49494_(_39120_, _39143_, _39144_);
  or g_49495_(_39119_, _39130_, _39145_);
  or g_49496_(_39144_, _39145_, _39146_);
  or g_49497_(_39123_, _39128_, _39147_);
  or g_49498_(_39131_, _39147_, _39148_);
  or g_49499_(_39146_, _39148_, _39149_);
  or g_49500_(_39142_, _39149_, _39150_);
  or g_49501_(_39135_, _39150_, _39151_);
  xor g_49502_(out[156], out[508], _39152_);
  and g_49503_(_39603_, out[507], _39153_);
  xor g_49504_(out[157], out[509], _39154_);
  xor g_49505_(out[150], out[502], _39155_);
  xor g_49506_(out[152], out[504], _39156_);
  xor g_49507_(out[153], out[505], _39157_);
  xor g_49508_(out[158], out[510], _39158_);
  xor g_49509_(out[148], out[500], _39159_);
  or g_49510_(_39158_, _39159_, _39160_);
  xor g_49511_(out[149], out[501], _39161_);
  xor g_49512_(out[145], out[497], _39162_);
  and g_49513_(out[155], _39845_, _39163_);
  xor g_49514_(out[159], out[511], _39164_);
  xor g_49515_(out[154], out[506], _39165_);
  xor g_49516_(out[144], out[496], _39166_);
  xor g_49517_(out[146], out[498], _39167_);
  xor g_49518_(out[147], out[499], _39168_);
  or g_49519_(_39154_, _39156_, _39169_);
  or g_49520_(_39165_, _39167_, _39170_);
  or g_49521_(_39169_, _39170_, _39171_);
  or g_49522_(_39157_, _39168_, _39172_);
  or g_49523_(_39161_, _39166_, _39173_);
  or g_49524_(_39172_, _39173_, _39174_);
  or g_49525_(_39171_, _39174_, _39175_);
  or g_49526_(_39152_, _39153_, _39176_);
  xor g_49527_(out[151], out[503], _39177_);
  or g_49528_(_39155_, _39177_, _39178_);
  or g_49529_(_39176_, _39178_, _39179_);
  or g_49530_(_39162_, _39163_, _39180_);
  or g_49531_(_39164_, _39180_, _39181_);
  or g_49532_(_39179_, _39181_, _39182_);
  or g_49533_(_39175_, _39182_, _39183_);
  or g_49534_(_39160_, _39183_, _39184_);
  not g_49535_(_39184_, _39185_);
  xor g_49536_(out[135], out[503], _39186_);
  and g_49537_(_39592_, out[507], _39187_);
  xor g_49538_(out[142], out[510], _39188_);
  xor g_49539_(out[136], out[504], _39189_);
  xor g_49540_(out[129], out[497], _39190_);
  xor g_49541_(out[141], out[509], _39191_);
  xor g_49542_(out[137], out[505], _39192_);
  xor g_49543_(out[132], out[500], _39193_);
  xor g_49544_(out[130], out[498], _39194_);
  and g_49545_(out[139], _39845_, _39195_);
  xor g_49546_(out[131], out[499], _39196_);
  xor g_49547_(out[134], out[502], _39197_);
  xor g_49548_(out[143], out[511], _39198_);
  xor g_49549_(out[138], out[506], _39199_);
  xor g_49550_(out[133], out[501], _39200_);
  xor g_49551_(out[128], out[496], _39201_);
  or g_49552_(_39188_, _39193_, _39202_);
  or g_49553_(_39189_, _39191_, _39203_);
  or g_49554_(_39194_, _39199_, _39204_);
  or g_49555_(_39203_, _39204_, _39205_);
  or g_49556_(_39192_, _39196_, _39206_);
  or g_49557_(_39200_, _39201_, _39207_);
  or g_49558_(_39206_, _39207_, _39208_);
  or g_49559_(_39205_, _39208_, _39209_);
  xor g_49560_(out[140], out[508], _39210_);
  or g_49561_(_39187_, _39210_, _39211_);
  or g_49562_(_39186_, _39197_, _39212_);
  or g_49563_(_39211_, _39212_, _39213_);
  or g_49564_(_39190_, _39195_, _39214_);
  or g_49565_(_39198_, _39214_, _39215_);
  or g_49566_(_39213_, _39215_, _39216_);
  or g_49567_(_39209_, _39216_, _39217_);
  or g_49568_(_39202_, _39217_, _39218_);
  not g_49569_(_39218_, _39219_);
  xor g_49570_(out[113], out[497], _39220_);
  and g_49571_(out[123], _39845_, _39221_);
  xor g_49572_(out[126], out[510], _39222_);
  xor g_49573_(out[115], out[499], _39223_);
  xor g_49574_(out[116], out[500], _39224_);
  xor g_49575_(out[114], out[498], _39225_);
  xor g_49576_(out[121], out[505], _39226_);
  xor g_49577_(out[112], out[496], _39227_);
  and g_49578_(_39581_, out[507], _39228_);
  xor g_49579_(out[118], out[502], _39229_);
  xor g_49580_(out[122], out[506], _39230_);
  xor g_49581_(out[117], out[501], _39231_);
  xor g_49582_(out[127], out[511], _39232_);
  xor g_49583_(out[125], out[509], _39233_);
  xor g_49584_(out[120], out[504], _39234_);
  or g_49585_(_39222_, _39224_, _39235_);
  or g_49586_(_39233_, _39234_, _39236_);
  or g_49587_(_39225_, _39230_, _39237_);
  or g_49588_(_39236_, _39237_, _39238_);
  or g_49589_(_39223_, _39226_, _39239_);
  or g_49590_(_39227_, _39231_, _39240_);
  or g_49591_(_39239_, _39240_, _39241_);
  or g_49592_(_39238_, _39241_, _39242_);
  xor g_49593_(out[124], out[508], _39243_);
  or g_49594_(_39228_, _39243_, _39244_);
  xor g_49595_(out[119], out[503], _39245_);
  or g_49596_(_39229_, _39245_, _39246_);
  or g_49597_(_39244_, _39246_, _39247_);
  or g_49598_(_39220_, _39221_, _39248_);
  or g_49599_(_39232_, _39248_, _39249_);
  or g_49600_(_39247_, _39249_, _39250_);
  or g_49601_(_39242_, _39250_, _39251_);
  or g_49602_(_39235_, _39251_, _39252_);
  not g_49603_(_39252_, _39253_);
  xor g_49604_(out[103], out[503], _39254_);
  and g_49605_(_39570_, out[507], _39255_);
  xor g_49606_(out[110], out[510], _39256_);
  xor g_49607_(out[104], out[504], _39257_);
  xor g_49608_(out[97], out[497], _39258_);
  xor g_49609_(out[109], out[509], _39259_);
  xor g_49610_(out[105], out[505], _39260_);
  xor g_49611_(out[100], out[500], _39261_);
  xor g_49612_(out[98], out[498], _39262_);
  and g_49613_(out[107], _39845_, _39263_);
  xor g_49614_(out[99], out[499], _39264_);
  xor g_49615_(out[102], out[502], _39265_);
  xor g_49616_(out[111], out[511], _39266_);
  xor g_49617_(out[106], out[506], _39267_);
  xor g_49618_(out[101], out[501], _39268_);
  xor g_49619_(out[96], out[496], _39269_);
  or g_49620_(_39256_, _39261_, _39270_);
  or g_49621_(_39257_, _39259_, _39271_);
  or g_49622_(_39262_, _39267_, _39272_);
  or g_49623_(_39271_, _39272_, _39273_);
  or g_49624_(_39260_, _39264_, _39274_);
  or g_49625_(_39268_, _39269_, _39275_);
  or g_49626_(_39274_, _39275_, _39276_);
  or g_49627_(_39273_, _39276_, _39277_);
  xor g_49628_(out[108], out[508], _39278_);
  or g_49629_(_39255_, _39278_, _39279_);
  or g_49630_(_39254_, _39265_, _39280_);
  or g_49631_(_39279_, _39280_, _39281_);
  or g_49632_(_39258_, _39263_, _39282_);
  or g_49633_(_39266_, _39282_, _39283_);
  or g_49634_(_39281_, _39283_, _39284_);
  or g_49635_(_39277_, _39284_, _39285_);
  or g_49636_(_39270_, _39285_, _39286_);
  xor g_49637_(out[83], out[499], _39287_);
  xor g_49638_(out[84], out[500], _39288_);
  xor g_49639_(out[94], out[510], _39289_);
  xor g_49640_(out[82], out[498], _39290_);
  xor g_49641_(out[85], out[501], _39291_);
  xor g_49642_(out[89], out[505], _39292_);
  xor g_49643_(out[88], out[504], _39293_);
  xor g_49644_(out[95], out[511], _39294_);
  xor g_49645_(out[90], out[506], _39296_);
  xor g_49646_(out[86], out[502], _39297_);
  xor g_49647_(out[80], out[496], _39298_);
  and g_49648_(_39559_, out[507], _39299_);
  and g_49649_(out[91], _39845_, _39300_);
  xor g_49650_(out[93], out[509], _39301_);
  or g_49651_(_39293_, _39301_, _39302_);
  xor g_49652_(out[81], out[497], _39303_);
  or g_49653_(_39290_, _39296_, _39304_);
  or g_49654_(_39302_, _39304_, _39305_);
  or g_49655_(_39287_, _39292_, _39307_);
  or g_49656_(_39291_, _39307_, _39308_);
  or g_49657_(_39305_, _39308_, _39309_);
  or g_49658_(_39288_, _39289_, _39310_);
  or g_49659_(_39309_, _39310_, _39311_);
  xor g_49660_(out[92], out[508], _39312_);
  or g_49661_(_39299_, _39312_, _39313_);
  xor g_49662_(out[87], out[503], _39314_);
  or g_49663_(_39297_, _39314_, _39315_);
  or g_49664_(_39313_, _39315_, _39316_);
  or g_49665_(_39300_, _39303_, _39318_);
  or g_49666_(_39294_, _39318_, _39319_);
  or g_49667_(_39316_, _39319_, _39320_);
  or g_49668_(_39298_, _39320_, _39321_);
  or g_49669_(_39311_, _39321_, _39322_);
  not g_49670_(_39322_, _39323_);
  xor g_49671_(out[71], out[503], _39324_);
  and g_49672_(_39548_, out[507], _39325_);
  xor g_49673_(out[78], out[510], _39326_);
  xor g_49674_(out[72], out[504], _39327_);
  xor g_49675_(out[65], out[497], _39329_);
  xor g_49676_(out[77], out[509], _39330_);
  xor g_49677_(out[73], out[505], _39331_);
  xor g_49678_(out[68], out[500], _39332_);
  xor g_49679_(out[66], out[498], _39333_);
  and g_49680_(out[75], _39845_, _39334_);
  xor g_49681_(out[67], out[499], _39335_);
  xor g_49682_(out[70], out[502], _39336_);
  xor g_49683_(out[79], out[511], _39337_);
  xor g_49684_(out[74], out[506], _39338_);
  xor g_49685_(out[69], out[501], _39340_);
  xor g_49686_(out[64], out[496], _39341_);
  or g_49687_(_39326_, _39332_, _39342_);
  or g_49688_(_39327_, _39330_, _39343_);
  or g_49689_(_39333_, _39338_, _39344_);
  or g_49690_(_39343_, _39344_, _39345_);
  or g_49691_(_39331_, _39335_, _39346_);
  or g_49692_(_39340_, _39341_, _39347_);
  or g_49693_(_39346_, _39347_, _39348_);
  or g_49694_(_39345_, _39348_, _39349_);
  xor g_49695_(out[76], out[508], _39351_);
  or g_49696_(_39325_, _39351_, _39352_);
  or g_49697_(_39324_, _39336_, _39353_);
  or g_49698_(_39352_, _39353_, _39354_);
  or g_49699_(_39329_, _39334_, _39355_);
  or g_49700_(_39337_, _39355_, _39356_);
  or g_49701_(_39354_, _39356_, _39357_);
  or g_49702_(_39349_, _39357_, _39358_);
  or g_49703_(_39342_, _39358_, _39359_);
  not g_49704_(_39359_, _39360_);
  xor g_49705_(out[60], out[508], _39362_);
  and g_49706_(_39537_, out[507], _39363_);
  xor g_49707_(out[56], out[504], _39364_);
  xor g_49708_(out[54], out[502], _39365_);
  xor g_49709_(out[61], out[509], _39366_);
  xor g_49710_(out[62], out[510], _39367_);
  xor g_49711_(out[50], out[498], _39368_);
  xor g_49712_(out[57], out[505], _39369_);
  xor g_49713_(out[53], out[501], _39370_);
  xor g_49714_(out[49], out[497], _39371_);
  and g_49715_(out[59], _39845_, _39373_);
  or g_49716_(_39364_, _39366_, _39374_);
  xor g_49717_(out[63], out[511], _39375_);
  xor g_49718_(out[58], out[506], _39376_);
  xor g_49719_(out[52], out[500], _39377_);
  xor g_49720_(out[51], out[499], _39378_);
  xor g_49721_(out[48], out[496], _39379_);
  or g_49722_(_39368_, _39376_, _39380_);
  or g_49723_(_39374_, _39380_, _39381_);
  or g_49724_(_39369_, _39378_, _39382_);
  or g_49725_(_39370_, _39382_, _39384_);
  or g_49726_(_39381_, _39384_, _39385_);
  or g_49727_(_39367_, _39377_, _39386_);
  or g_49728_(_39385_, _39386_, _39387_);
  or g_49729_(_39362_, _39363_, _39388_);
  xor g_49730_(out[55], out[503], _39389_);
  or g_49731_(_39365_, _39389_, _39390_);
  or g_49732_(_39388_, _39390_, _39391_);
  or g_49733_(_39371_, _39373_, _39392_);
  or g_49734_(_39375_, _39392_, _39393_);
  or g_49735_(_39391_, _39393_, _39395_);
  or g_49736_(_39379_, _39395_, _39396_);
  or g_49737_(_39387_, _39396_, _39397_);
  not g_49738_(_39397_, _39398_);
  xor g_49739_(out[39], out[503], _39399_);
  and g_49740_(_39526_, out[507], _39400_);
  xor g_49741_(out[46], out[510], _39401_);
  xor g_49742_(out[40], out[504], _39402_);
  xor g_49743_(out[33], out[497], _39403_);
  xor g_49744_(out[45], out[509], _39404_);
  xor g_49745_(out[41], out[505], _39406_);
  xor g_49746_(out[36], out[500], _39407_);
  xor g_49747_(out[34], out[498], _39408_);
  and g_49748_(out[43], _39845_, _39409_);
  xor g_49749_(out[35], out[499], _39410_);
  xor g_49750_(out[38], out[502], _39411_);
  xor g_49751_(out[47], out[511], _39412_);
  xor g_49752_(out[42], out[506], _39413_);
  xor g_49753_(out[37], out[501], _39414_);
  xor g_49754_(out[32], out[496], _39415_);
  or g_49755_(_39401_, _39407_, _39417_);
  or g_49756_(_39402_, _39404_, _39418_);
  or g_49757_(_39408_, _39413_, _39419_);
  or g_49758_(_39418_, _39419_, _39420_);
  or g_49759_(_39406_, _39410_, _39421_);
  or g_49760_(_39414_, _39415_, _39422_);
  or g_49761_(_39421_, _39422_, _39423_);
  or g_49762_(_39420_, _39423_, _39424_);
  xor g_49763_(out[44], out[508], _39425_);
  or g_49764_(_39400_, _39425_, _39426_);
  or g_49765_(_39399_, _39411_, _39428_);
  or g_49766_(_39426_, _39428_, _39429_);
  or g_49767_(_39403_, _39409_, _39430_);
  or g_49768_(_39412_, _39430_, _39431_);
  or g_49769_(_39429_, _39431_, _39432_);
  or g_49770_(_39424_, _39432_, _39433_);
  or g_49771_(_39417_, _39433_, _39434_);
  xor g_49772_(out[29], out[509], _39435_);
  xor g_49773_(out[18], out[498], _39436_);
  xor g_49774_(out[21], out[501], _39437_);
  xor g_49775_(out[25], out[505], _39439_);
  xor g_49776_(out[20], out[500], _39440_);
  xor g_49777_(out[24], out[504], _39441_);
  xor g_49778_(out[30], out[510], _39442_);
  xor g_49779_(out[22], out[502], _39443_);
  xor g_49780_(out[31], out[511], _39444_);
  xor g_49781_(out[26], out[506], _39445_);
  xor g_49782_(out[16], out[496], _39446_);
  xor g_49783_(out[19], out[499], _39447_);
  and g_49784_(_39493_, out[507], _39448_);
  and g_49785_(out[27], _39845_, _39450_);
  xor g_49786_(out[17], out[497], _39451_);
  or g_49787_(_39440_, _39442_, _39452_);
  or g_49788_(_39435_, _39441_, _39453_);
  or g_49789_(_39436_, _39445_, _39454_);
  or g_49790_(_39453_, _39454_, _39455_);
  or g_49791_(_39439_, _39447_, _39456_);
  or g_49792_(_39437_, _39446_, _39457_);
  or g_49793_(_39456_, _39457_, _39458_);
  or g_49794_(_39455_, _39458_, _39459_);
  xor g_49795_(out[28], out[508], _39461_);
  or g_49796_(_39448_, _39461_, _39462_);
  xor g_49797_(out[23], out[503], _39463_);
  or g_49798_(_39443_, _39463_, _39464_);
  or g_49799_(_39462_, _39464_, _39465_);
  or g_49800_(_39450_, _39451_, _39466_);
  or g_49801_(_39444_, _39466_, _39467_);
  or g_49802_(_39465_, _39467_, _39468_);
  or g_49803_(_39459_, _39468_, _39469_);
  or g_49804_(_39452_, _39469_, _39470_);
  xor g_49805_(out[1], out[497], _39472_);
  and g_49806_(out[11], _39845_, _39473_);
  xor g_49807_(out[9], out[505], _39474_);
  xor g_49808_(out[0], out[496], _39475_);
  xor g_49809_(out[14], out[510], _39476_);
  xor g_49810_(out[4], out[500], _39477_);
  or g_49811_(_39476_, _39477_, _39478_);
  xor g_49812_(out[13], out[509], _39479_);
  xor g_49813_(out[3], out[499], _39480_);
  and g_49814_(_39438_, out[507], _39481_);
  xor g_49815_(out[6], out[502], _39483_);
  xor g_49816_(out[10], out[506], _39484_);
  xor g_49817_(out[5], out[501], _39485_);
  xor g_49818_(out[15], out[511], _39486_);
  xor g_49819_(out[8], out[504], _39487_);
  or g_49820_(_39479_, _39487_, _39488_);
  xor g_49821_(out[2], out[498], _39489_);
  or g_49822_(_39484_, _39489_, _39490_);
  or g_49823_(_39488_, _39490_, _39491_);
  or g_49824_(_39474_, _39480_, _39492_);
  or g_49825_(_39485_, _39492_, _39494_);
  or g_49826_(_39491_, _39494_, _39495_);
  or g_49827_(_39478_, _39495_, _39496_);
  xor g_49828_(out[12], out[508], _39497_);
  or g_49829_(_39481_, _39497_, _39498_);
  xor g_49830_(out[7], out[503], _39499_);
  or g_49831_(_39483_, _39499_, _39500_);
  or g_49832_(_39498_, _39500_, _39501_);
  or g_49833_(_39472_, _39473_, _39502_);
  or g_49834_(_39486_, _39502_, _39503_);
  or g_49835_(_39501_, _39503_, _39505_);
  or g_49836_(_39475_, _39505_, _39506_);
  or g_49837_(_39496_, _39506_, _39507_);
  xor g_49838_(out[311], out[487], _39508_);
  and g_49839_(_39724_, out[491], _39509_);
  xor g_49840_(out[318], out[494], _39510_);
  xor g_49841_(out[312], out[488], _39511_);
  xor g_49842_(out[305], out[481], _39512_);
  xor g_49843_(out[317], out[493], _39513_);
  xor g_49844_(out[313], out[489], _39514_);
  xor g_49845_(out[308], out[484], _39516_);
  xor g_49846_(out[306], out[482], _39517_);
  and g_49847_(out[315], _39834_, _39518_);
  xor g_49848_(out[307], out[483], _39519_);
  xor g_49849_(out[310], out[486], _39520_);
  xor g_49850_(out[319], out[495], _39521_);
  xor g_49851_(out[314], out[490], _39522_);
  xor g_49852_(out[309], out[485], _39523_);
  xor g_49853_(out[304], out[480], _39524_);
  or g_49854_(_39510_, _39516_, _39525_);
  or g_49855_(_39511_, _39513_, _39527_);
  or g_49856_(_39517_, _39522_, _39528_);
  or g_49857_(_39527_, _39528_, _39529_);
  or g_49858_(_39514_, _39519_, _39530_);
  or g_49859_(_39523_, _39524_, _39531_);
  or g_49860_(_39530_, _39531_, _39532_);
  or g_49861_(_39529_, _39532_, _39533_);
  xor g_49862_(out[316], out[492], _39534_);
  or g_49863_(_39509_, _39534_, _39535_);
  or g_49864_(_39508_, _39520_, _39536_);
  or g_49865_(_39535_, _39536_, _39538_);
  or g_49866_(_39512_, _39518_, _39539_);
  or g_49867_(_39521_, _39539_, _39540_);
  or g_49868_(_39538_, _39540_, _39541_);
  or g_49869_(_39533_, _39541_, _39542_);
  or g_49870_(_39525_, _39542_, _39543_);
  xor g_49871_(out[296], out[488], _39544_);
  xor g_49872_(out[293], out[485], _39545_);
  xor g_49873_(out[291], out[483], _39546_);
  xor g_49874_(out[302], out[494], _39547_);
  xor g_49875_(out[301], out[493], _39549_);
  xor g_49876_(out[290], out[482], _39550_);
  xor g_49877_(out[297], out[489], _39551_);
  xor g_49878_(out[294], out[486], _39552_);
  xor g_49879_(out[303], out[495], _39553_);
  xor g_49880_(out[298], out[490], _39554_);
  xor g_49881_(out[292], out[484], _39555_);
  xor g_49882_(out[288], out[480], _39556_);
  and g_49883_(_39702_, out[491], _39557_);
  and g_49884_(out[299], _39834_, _39558_);
  or g_49885_(_39544_, _39549_, _39560_);
  xor g_49886_(out[289], out[481], _39561_);
  or g_49887_(_39550_, _39554_, _39562_);
  or g_49888_(_39560_, _39562_, _39563_);
  or g_49889_(_39546_, _39551_, _39564_);
  or g_49890_(_39545_, _39564_, _39565_);
  or g_49891_(_39563_, _39565_, _39566_);
  or g_49892_(_39547_, _39555_, _39567_);
  or g_49893_(_39566_, _39567_, _39568_);
  xor g_49894_(out[300], out[492], _39569_);
  or g_49895_(_39557_, _39569_, _39571_);
  xor g_49896_(out[295], out[487], _39572_);
  or g_49897_(_39552_, _39572_, _39573_);
  or g_49898_(_39571_, _39573_, _39574_);
  or g_49899_(_39558_, _39561_, _39575_);
  or g_49900_(_39553_, _39575_, _39576_);
  or g_49901_(_39574_, _39576_, _39577_);
  or g_49902_(_39556_, _39577_, _39578_);
  or g_49903_(_39568_, _39578_, _39579_);
  not g_49904_(_39579_, _39580_);
  xor g_49905_(out[279], out[487], _39582_);
  and g_49906_(_39691_, out[491], _39583_);
  xor g_49907_(out[286], out[494], _39584_);
  xor g_49908_(out[280], out[488], _39585_);
  xor g_49909_(out[273], out[481], _39586_);
  xor g_49910_(out[285], out[493], _39587_);
  xor g_49911_(out[281], out[489], _39588_);
  xor g_49912_(out[276], out[484], _39589_);
  xor g_49913_(out[274], out[482], _39590_);
  and g_49914_(out[283], _39834_, _39591_);
  xor g_49915_(out[275], out[483], _39593_);
  xor g_49916_(out[278], out[486], _39594_);
  xor g_49917_(out[287], out[495], _39595_);
  xor g_49918_(out[282], out[490], _39596_);
  xor g_49919_(out[277], out[485], _39597_);
  xor g_49920_(out[272], out[480], _39598_);
  or g_49921_(_39584_, _39589_, _39599_);
  or g_49922_(_39585_, _39587_, _39600_);
  or g_49923_(_39590_, _39596_, _39601_);
  or g_49924_(_39600_, _39601_, _39602_);
  or g_49925_(_39588_, _39593_, _39604_);
  or g_49926_(_39597_, _39598_, _39605_);
  or g_49927_(_39604_, _39605_, _39606_);
  or g_49928_(_39602_, _39606_, _39607_);
  xor g_49929_(out[284], out[492], _39608_);
  or g_49930_(_39583_, _39608_, _39609_);
  or g_49931_(_39582_, _39594_, _39610_);
  or g_49932_(_39609_, _39610_, _39611_);
  or g_49933_(_39586_, _39591_, _39612_);
  or g_49934_(_39595_, _39612_, _39613_);
  or g_49935_(_39611_, _39613_, _39615_);
  or g_49936_(_39607_, _39615_, _39616_);
  or g_49937_(_39599_, _39616_, _39617_);
  xor g_49938_(out[268], out[492], _39618_);
  and g_49939_(_39680_, out[491], _39619_);
  xor g_49940_(out[264], out[488], _39620_);
  xor g_49941_(out[262], out[486], _39621_);
  xor g_49942_(out[269], out[493], _39622_);
  xor g_49943_(out[270], out[494], _39623_);
  xor g_49944_(out[258], out[482], _39624_);
  xor g_49945_(out[265], out[489], _39626_);
  xor g_49946_(out[261], out[485], _39627_);
  xor g_49947_(out[257], out[481], _39628_);
  and g_49948_(out[267], _39834_, _39629_);
  or g_49949_(_39620_, _39622_, _39630_);
  xor g_49950_(out[271], out[495], _39631_);
  xor g_49951_(out[266], out[490], _39632_);
  xor g_49952_(out[260], out[484], _39633_);
  xor g_49953_(out[259], out[483], _39634_);
  xor g_49954_(out[256], out[480], _39635_);
  or g_49955_(_39624_, _39632_, _39637_);
  or g_49956_(_39630_, _39637_, _39638_);
  or g_49957_(_39626_, _39634_, _39639_);
  or g_49958_(_39627_, _39639_, _39640_);
  or g_49959_(_39638_, _39640_, _39641_);
  or g_49960_(_39623_, _39633_, _39642_);
  or g_49961_(_39641_, _39642_, _39643_);
  or g_49962_(_39618_, _39619_, _39644_);
  xor g_49963_(out[263], out[487], _39645_);
  or g_49964_(_39621_, _39645_, _39646_);
  or g_49965_(_39644_, _39646_, _39648_);
  or g_49966_(_39628_, _39629_, _39649_);
  or g_49967_(_39631_, _39649_, _39650_);
  or g_49968_(_39648_, _39650_, _39651_);
  or g_49969_(_39635_, _39651_, _39652_);
  or g_49970_(_39643_, _39652_, _39653_);
  xor g_49971_(out[247], out[487], _39654_);
  and g_49972_(_39669_, out[491], _39655_);
  xor g_49973_(out[254], out[494], _39656_);
  xor g_49974_(out[248], out[488], _39657_);
  xor g_49975_(out[241], out[481], _39659_);
  xor g_49976_(out[253], out[493], _39660_);
  xor g_49977_(out[249], out[489], _39661_);
  xor g_49978_(out[244], out[484], _39662_);
  xor g_49979_(out[242], out[482], _39663_);
  and g_49980_(out[251], _39834_, _39664_);
  xor g_49981_(out[243], out[483], _39665_);
  xor g_49982_(out[246], out[486], _39666_);
  xor g_49983_(out[255], out[495], _39667_);
  xor g_49984_(out[250], out[490], _39668_);
  xor g_49985_(out[245], out[485], _39670_);
  xor g_49986_(out[240], out[480], _39671_);
  or g_49987_(_39656_, _39662_, _39672_);
  or g_49988_(_39657_, _39660_, _39673_);
  or g_49989_(_39663_, _39668_, _39674_);
  or g_49990_(_39673_, _39674_, _39675_);
  or g_49991_(_39661_, _39665_, _39676_);
  or g_49992_(_39670_, _39671_, _39677_);
  or g_49993_(_39676_, _39677_, _39678_);
  or g_49994_(_39675_, _39678_, _39679_);
  xor g_49995_(out[252], out[492], _39681_);
  or g_49996_(_39655_, _39681_, _39682_);
  or g_49997_(_39654_, _39666_, _39683_);
  or g_49998_(_39682_, _39683_, _39684_);
  or g_49999_(_39659_, _39664_, _39685_);
  or g_50000_(_39667_, _39685_, _39686_);
  or g_50001_(_39684_, _39686_, _39687_);
  or g_50002_(_39679_, _39687_, _39688_);
  or g_50003_(_39672_, _39688_, _39689_);
  not g_50004_(_39689_, _39690_);
  and g_50005_(out[235], _39834_, _39692_);
  and g_50006_(_39658_, out[491], _39693_);
  xor g_50007_(out[232], out[488], _39694_);
  xor g_50008_(out[239], out[495], _39695_);
  xor g_50009_(out[225], out[481], _39696_);
  xor g_50010_(out[226], out[482], _39697_);
  xor g_50011_(out[228], out[484], _39698_);
  xor g_50012_(out[237], out[493], _39699_);
  xor g_50013_(out[233], out[489], _39700_);
  xor g_50014_(out[227], out[483], _39701_);
  xor g_50015_(out[229], out[485], _39703_);
  xor g_50016_(out[238], out[494], _39704_);
  xor g_50017_(out[224], out[480], _39705_);
  xor g_50018_(out[234], out[490], _39706_);
  or g_50019_(_39694_, _39699_, _39707_);
  xor g_50020_(out[230], out[486], _39708_);
  or g_50021_(_39697_, _39706_, _39709_);
  or g_50022_(_39707_, _39709_, _39710_);
  or g_50023_(_39700_, _39701_, _39711_);
  or g_50024_(_39703_, _39711_, _39712_);
  or g_50025_(_39710_, _39712_, _39714_);
  or g_50026_(_39698_, _39704_, _39715_);
  or g_50027_(_39714_, _39715_, _39716_);
  xor g_50028_(out[236], out[492], _39717_);
  or g_50029_(_39693_, _39717_, _39718_);
  xor g_50030_(out[231], out[487], _39719_);
  or g_50031_(_39708_, _39719_, _39720_);
  or g_50032_(_39718_, _39720_, _39721_);
  or g_50033_(_39692_, _39696_, _39722_);
  or g_50034_(_39695_, _39722_, _39723_);
  or g_50035_(_39721_, _39723_, _39725_);
  or g_50036_(_39705_, _39725_, _39726_);
  or g_50037_(_39716_, _39726_, _39727_);
  not g_50038_(_39727_, _39728_);
  xor g_50039_(out[215], out[487], _39729_);
  and g_50040_(_39647_, out[491], _39730_);
  xor g_50041_(out[222], out[494], _39731_);
  xor g_50042_(out[216], out[488], _39732_);
  xor g_50043_(out[209], out[481], _39733_);
  xor g_50044_(out[221], out[493], _39734_);
  xor g_50045_(out[217], out[489], _39736_);
  xor g_50046_(out[212], out[484], _39737_);
  xor g_50047_(out[210], out[482], _39738_);
  and g_50048_(out[219], _39834_, _39739_);
  xor g_50049_(out[211], out[483], _39740_);
  xor g_50050_(out[214], out[486], _39741_);
  xor g_50051_(out[223], out[495], _39742_);
  xor g_50052_(out[218], out[490], _39743_);
  xor g_50053_(out[213], out[485], _39744_);
  xor g_50054_(out[208], out[480], _39745_);
  or g_50055_(_39731_, _39737_, _39747_);
  or g_50056_(_39732_, _39734_, _39748_);
  or g_50057_(_39738_, _39743_, _39749_);
  or g_50058_(_39748_, _39749_, _39750_);
  or g_50059_(_39736_, _39740_, _39751_);
  or g_50060_(_39744_, _39745_, _39752_);
  or g_50061_(_39751_, _39752_, _39753_);
  or g_50062_(_39750_, _39753_, _39754_);
  xor g_50063_(out[220], out[492], _39755_);
  or g_50064_(_39730_, _39755_, _39756_);
  or g_50065_(_39729_, _39741_, _39758_);
  or g_50066_(_39756_, _39758_, _39759_);
  or g_50067_(_39733_, _39739_, _39760_);
  or g_50068_(_39742_, _39760_, _39761_);
  or g_50069_(_39759_, _39761_, _39762_);
  or g_50070_(_39754_, _39762_, _39763_);
  or g_50071_(_39747_, _39763_, _39764_);
  xor g_50072_(out[204], out[492], _39765_);
  and g_50073_(_39636_, out[491], _39766_);
  xor g_50074_(out[205], out[493], _39767_);
  xor g_50075_(out[198], out[486], _39769_);
  xor g_50076_(out[200], out[488], _39770_);
  xor g_50077_(out[201], out[489], _39771_);
  xor g_50078_(out[206], out[494], _39772_);
  xor g_50079_(out[196], out[484], _39773_);
  or g_50080_(_39772_, _39773_, _39774_);
  xor g_50081_(out[197], out[485], _39775_);
  xor g_50082_(out[193], out[481], _39776_);
  and g_50083_(out[203], _39834_, _39777_);
  xor g_50084_(out[207], out[495], _39778_);
  xor g_50085_(out[202], out[490], _39780_);
  xor g_50086_(out[192], out[480], _39781_);
  xor g_50087_(out[194], out[482], _39782_);
  xor g_50088_(out[195], out[483], _39783_);
  or g_50089_(_39767_, _39770_, _39784_);
  or g_50090_(_39780_, _39782_, _39785_);
  or g_50091_(_39784_, _39785_, _39786_);
  or g_50092_(_39771_, _39783_, _39787_);
  or g_50093_(_39775_, _39781_, _39788_);
  or g_50094_(_39787_, _39788_, _39789_);
  or g_50095_(_39786_, _39789_, _39791_);
  or g_50096_(_39765_, _39766_, _39792_);
  xor g_50097_(out[199], out[487], _39793_);
  or g_50098_(_39769_, _39793_, _39794_);
  or g_50099_(_39792_, _39794_, _39795_);
  or g_50100_(_39776_, _39777_, _39796_);
  or g_50101_(_39778_, _39796_, _39797_);
  or g_50102_(_39795_, _39797_, _39798_);
  or g_50103_(_39791_, _39798_, _39799_);
  or g_50104_(_39774_, _39799_, _39800_);
  xor g_50105_(out[183], out[487], _39802_);
  and g_50106_(_39625_, out[491], _39803_);
  xor g_50107_(out[190], out[494], _39804_);
  xor g_50108_(out[184], out[488], _39805_);
  xor g_50109_(out[177], out[481], _39806_);
  xor g_50110_(out[189], out[493], _39807_);
  xor g_50111_(out[185], out[489], _39808_);
  xor g_50112_(out[180], out[484], _39809_);
  xor g_50113_(out[178], out[482], _39810_);
  and g_50114_(out[187], _39834_, _39811_);
  xor g_50115_(out[179], out[483], _39813_);
  xor g_50116_(out[182], out[486], _39814_);
  xor g_50117_(out[191], out[495], _39815_);
  xor g_50118_(out[186], out[490], _39816_);
  xor g_50119_(out[181], out[485], _39817_);
  xor g_50120_(out[176], out[480], _39818_);
  or g_50121_(_39804_, _39809_, _39819_);
  or g_50122_(_39805_, _39807_, _39820_);
  or g_50123_(_39810_, _39816_, _39821_);
  or g_50124_(_39820_, _39821_, _39822_);
  or g_50125_(_39808_, _39813_, _39824_);
  or g_50126_(_39817_, _39818_, _39825_);
  or g_50127_(_39824_, _39825_, _39826_);
  or g_50128_(_39822_, _39826_, _39827_);
  xor g_50129_(out[188], out[492], _39828_);
  or g_50130_(_39803_, _39828_, _39829_);
  or g_50131_(_39802_, _39814_, _39830_);
  or g_50132_(_39829_, _39830_, _39831_);
  or g_50133_(_39806_, _39811_, _39832_);
  or g_50134_(_39815_, _39832_, _39833_);
  or g_50135_(_39831_, _39833_, _39835_);
  or g_50136_(_39827_, _39835_, _39836_);
  or g_50137_(_39819_, _39836_, _39837_);
  not g_50138_(_39837_, _39838_);
  xor g_50139_(out[161], out[481], _39839_);
  and g_50140_(out[171], _39834_, _39840_);
  xor g_50141_(out[169], out[489], _39841_);
  xor g_50142_(out[160], out[480], _39842_);
  xor g_50143_(out[174], out[494], _39843_);
  xor g_50144_(out[164], out[484], _39844_);
  or g_50145_(_39843_, _39844_, _39846_);
  xor g_50146_(out[173], out[493], _39847_);
  xor g_50147_(out[163], out[483], _39848_);
  and g_50148_(_39614_, out[491], _39849_);
  xor g_50149_(out[166], out[486], _39850_);
  xor g_50150_(out[170], out[490], _39851_);
  xor g_50151_(out[165], out[485], _39852_);
  xor g_50152_(out[175], out[495], _39853_);
  xor g_50153_(out[168], out[488], _39854_);
  or g_50154_(_39847_, _39854_, _39855_);
  xor g_50155_(out[162], out[482], _39857_);
  or g_50156_(_39851_, _39857_, _39858_);
  or g_50157_(_39855_, _39858_, _39859_);
  or g_50158_(_39841_, _39848_, _39860_);
  or g_50159_(_39852_, _39860_, _39861_);
  or g_50160_(_39859_, _39861_, _39862_);
  or g_50161_(_39846_, _39862_, _39863_);
  xor g_50162_(out[172], out[492], _39864_);
  or g_50163_(_39849_, _39864_, _39865_);
  xor g_50164_(out[167], out[487], _39866_);
  or g_50165_(_39850_, _39866_, _39868_);
  or g_50166_(_39865_, _39868_, _39869_);
  or g_50167_(_39839_, _39840_, _39870_);
  or g_50168_(_39853_, _39870_, _39871_);
  or g_50169_(_39869_, _39871_, _39872_);
  or g_50170_(_39842_, _39872_, _39873_);
  or g_50171_(_39863_, _39873_, _39874_);
  xor g_50172_(out[151], out[487], _39875_);
  and g_50173_(_39603_, out[491], _39876_);
  xor g_50174_(out[158], out[494], _39877_);
  xor g_50175_(out[152], out[488], _39879_);
  xor g_50176_(out[145], out[481], _39880_);
  xor g_50177_(out[157], out[493], _39881_);
  xor g_50178_(out[153], out[489], _39882_);
  xor g_50179_(out[148], out[484], _39883_);
  xor g_50180_(out[146], out[482], _39884_);
  and g_50181_(out[155], _39834_, _39885_);
  xor g_50182_(out[147], out[483], _39886_);
  xor g_50183_(out[150], out[486], _39887_);
  xor g_50184_(out[159], out[495], _39888_);
  xor g_50185_(out[154], out[490], _39890_);
  xor g_50186_(out[149], out[485], _39891_);
  xor g_50187_(out[144], out[480], _39892_);
  or g_50188_(_39877_, _39883_, _39893_);
  or g_50189_(_39879_, _39881_, _39894_);
  or g_50190_(_39884_, _39890_, _39895_);
  or g_50191_(_39894_, _39895_, _39896_);
  or g_50192_(_39882_, _39886_, _39897_);
  or g_50193_(_39891_, _39892_, _39898_);
  or g_50194_(_39897_, _39898_, _39899_);
  or g_50195_(_39896_, _39899_, _39901_);
  xor g_50196_(out[156], out[492], _39902_);
  or g_50197_(_39876_, _39902_, _39903_);
  or g_50198_(_39875_, _39887_, _39904_);
  or g_50199_(_39903_, _39904_, _39905_);
  or g_50200_(_39880_, _39885_, _39906_);
  or g_50201_(_39888_, _39906_, _39907_);
  or g_50202_(_39905_, _39907_, _39908_);
  or g_50203_(_39901_, _39908_, _39909_);
  or g_50204_(_39893_, _39909_, _39910_);
  xor g_50205_(out[129], out[481], _39912_);
  and g_50206_(out[139], _39834_, _39913_);
  xor g_50207_(out[137], out[489], _39914_);
  xor g_50208_(out[128], out[480], _39915_);
  xor g_50209_(out[142], out[494], _39916_);
  xor g_50210_(out[132], out[484], _39917_);
  or g_50211_(_39916_, _39917_, _39918_);
  xor g_50212_(out[141], out[493], _39919_);
  xor g_50213_(out[131], out[483], _39920_);
  and g_50214_(_39592_, out[491], _39921_);
  xor g_50215_(out[134], out[486], _39923_);
  xor g_50216_(out[138], out[490], _39924_);
  xor g_50217_(out[133], out[485], _39925_);
  xor g_50218_(out[143], out[495], _39926_);
  xor g_50219_(out[136], out[488], _39927_);
  or g_50220_(_39919_, _39927_, _39928_);
  xor g_50221_(out[130], out[482], _39929_);
  or g_50222_(_39924_, _39929_, _39930_);
  or g_50223_(_39928_, _39930_, _39931_);
  or g_50224_(_39914_, _39920_, _39932_);
  or g_50225_(_39925_, _39932_, _39934_);
  or g_50226_(_39931_, _39934_, _39935_);
  or g_50227_(_39918_, _39935_, _39936_);
  xor g_50228_(out[140], out[492], _39937_);
  or g_50229_(_39921_, _39937_, _39938_);
  xor g_50230_(out[135], out[487], _39939_);
  or g_50231_(_39923_, _39939_, _39940_);
  or g_50232_(_39938_, _39940_, _39941_);
  or g_50233_(_39912_, _39913_, _39942_);
  or g_50234_(_39926_, _39942_, _39943_);
  or g_50235_(_39941_, _39943_, _39945_);
  or g_50236_(_39915_, _39945_, _39946_);
  or g_50237_(_39936_, _39946_, _39947_);
  not g_50238_(_39947_, _39948_);
  xor g_50239_(out[119], out[487], _39949_);
  and g_50240_(_39581_, out[491], _39950_);
  xor g_50241_(out[126], out[494], _39951_);
  xor g_50242_(out[120], out[488], _39952_);
  xor g_50243_(out[113], out[481], _39953_);
  xor g_50244_(out[125], out[493], _39954_);
  xor g_50245_(out[121], out[489], _39956_);
  xor g_50246_(out[116], out[484], _39957_);
  xor g_50247_(out[114], out[482], _39958_);
  and g_50248_(out[123], _39834_, _39959_);
  xor g_50249_(out[115], out[483], _39960_);
  xor g_50250_(out[118], out[486], _39961_);
  xor g_50251_(out[127], out[495], _39962_);
  xor g_50252_(out[122], out[490], _39963_);
  xor g_50253_(out[117], out[485], _39964_);
  xor g_50254_(out[112], out[480], _39965_);
  or g_50255_(_39951_, _39957_, _39967_);
  or g_50256_(_39952_, _39954_, _39968_);
  or g_50257_(_39958_, _39963_, _39969_);
  or g_50258_(_39968_, _39969_, _39970_);
  or g_50259_(_39956_, _39960_, _39971_);
  or g_50260_(_39964_, _39965_, _39972_);
  or g_50261_(_39971_, _39972_, _39973_);
  or g_50262_(_39970_, _39973_, _39974_);
  xor g_50263_(out[124], out[492], _39975_);
  or g_50264_(_39950_, _39975_, _39976_);
  or g_50265_(_39949_, _39961_, _39978_);
  or g_50266_(_39976_, _39978_, _39979_);
  or g_50267_(_39953_, _39959_, _39980_);
  or g_50268_(_39962_, _39980_, _39981_);
  or g_50269_(_39979_, _39981_, _39982_);
  or g_50270_(_39974_, _39982_, _39983_);
  or g_50271_(_39967_, _39983_, _39984_);
  xor g_50272_(out[97], out[481], _39985_);
  and g_50273_(out[107], _39834_, _39986_);
  xor g_50274_(out[105], out[489], _39987_);
  xor g_50275_(out[96], out[480], _39989_);
  xor g_50276_(out[110], out[494], _39990_);
  xor g_50277_(out[100], out[484], _39991_);
  or g_50278_(_39990_, _39991_, _39992_);
  xor g_50279_(out[109], out[493], _39993_);
  xor g_50280_(out[99], out[483], _39994_);
  and g_50281_(_39570_, out[491], _39995_);
  xor g_50282_(out[102], out[486], _39996_);
  xor g_50283_(out[106], out[490], _39997_);
  xor g_50284_(out[101], out[485], _39998_);
  xor g_50285_(out[111], out[495], _40000_);
  xor g_50286_(out[104], out[488], _40001_);
  or g_50287_(_39993_, _40001_, _40002_);
  xor g_50288_(out[98], out[482], _40003_);
  or g_50289_(_39997_, _40003_, _40004_);
  or g_50290_(_40002_, _40004_, _40005_);
  or g_50291_(_39987_, _39994_, _40006_);
  or g_50292_(_39998_, _40006_, _40007_);
  or g_50293_(_40005_, _40007_, _40008_);
  or g_50294_(_39992_, _40008_, _40009_);
  xor g_50295_(out[108], out[492], _40011_);
  or g_50296_(_39995_, _40011_, _40012_);
  xor g_50297_(out[103], out[487], _40013_);
  or g_50298_(_39996_, _40013_, _40014_);
  or g_50299_(_40012_, _40014_, _40015_);
  or g_50300_(_39985_, _39986_, _40016_);
  or g_50301_(_40000_, _40016_, _40017_);
  or g_50302_(_40015_, _40017_, _40018_);
  or g_50303_(_39989_, _40018_, _40019_);
  or g_50304_(_40009_, _40019_, _40020_);
  not g_50305_(_40020_, _40022_);
  xor g_50306_(out[87], out[487], _40023_);
  and g_50307_(_39559_, out[491], _40024_);
  xor g_50308_(out[94], out[494], _40025_);
  xor g_50309_(out[88], out[488], _40026_);
  xor g_50310_(out[81], out[481], _40027_);
  xor g_50311_(out[93], out[493], _40028_);
  xor g_50312_(out[89], out[489], _40029_);
  xor g_50313_(out[84], out[484], _40030_);
  xor g_50314_(out[82], out[482], _40031_);
  and g_50315_(out[91], _39834_, _40033_);
  xor g_50316_(out[83], out[483], _40034_);
  xor g_50317_(out[86], out[486], _40035_);
  xor g_50318_(out[95], out[495], _40036_);
  xor g_50319_(out[90], out[490], _40037_);
  xor g_50320_(out[85], out[485], _40038_);
  xor g_50321_(out[80], out[480], _40039_);
  or g_50322_(_40025_, _40030_, _40040_);
  or g_50323_(_40026_, _40028_, _40041_);
  or g_50324_(_40031_, _40037_, _40042_);
  or g_50325_(_40041_, _40042_, _40044_);
  or g_50326_(_40029_, _40034_, _40045_);
  or g_50327_(_40038_, _40039_, _40046_);
  or g_50328_(_40045_, _40046_, _40047_);
  or g_50329_(_40044_, _40047_, _40048_);
  xor g_50330_(out[92], out[492], _40049_);
  or g_50331_(_40024_, _40049_, _40050_);
  or g_50332_(_40023_, _40035_, _40051_);
  or g_50333_(_40050_, _40051_, _40052_);
  or g_50334_(_40027_, _40033_, _40053_);
  or g_50335_(_40036_, _40053_, _40055_);
  or g_50336_(_40052_, _40055_, _40056_);
  or g_50337_(_40048_, _40056_, _40057_);
  or g_50338_(_40040_, _40057_, _40058_);
  not g_50339_(_40058_, _40059_);
  xor g_50340_(out[67], out[483], _40060_);
  xor g_50341_(out[68], out[484], _40061_);
  xor g_50342_(out[78], out[494], _40062_);
  xor g_50343_(out[66], out[482], _40063_);
  xor g_50344_(out[69], out[485], _40064_);
  xor g_50345_(out[73], out[489], _40066_);
  xor g_50346_(out[72], out[488], _40067_);
  xor g_50347_(out[79], out[495], _40068_);
  xor g_50348_(out[74], out[490], _40069_);
  xor g_50349_(out[70], out[486], _40070_);
  xor g_50350_(out[64], out[480], _40071_);
  and g_50351_(_39548_, out[491], _40072_);
  and g_50352_(out[75], _39834_, _40073_);
  xor g_50353_(out[77], out[493], _40074_);
  or g_50354_(_40067_, _40074_, _40075_);
  xor g_50355_(out[65], out[481], _40077_);
  or g_50356_(_40063_, _40069_, _40078_);
  or g_50357_(_40075_, _40078_, _40079_);
  or g_50358_(_40060_, _40066_, _40080_);
  or g_50359_(_40064_, _40080_, _40081_);
  or g_50360_(_40079_, _40081_, _40082_);
  or g_50361_(_40061_, _40062_, _40083_);
  or g_50362_(_40082_, _40083_, _40084_);
  xor g_50363_(out[76], out[492], _40085_);
  or g_50364_(_40072_, _40085_, _40086_);
  xor g_50365_(out[71], out[487], _40088_);
  or g_50366_(_40070_, _40088_, _40089_);
  or g_50367_(_40086_, _40089_, _40090_);
  or g_50368_(_40073_, _40077_, _40091_);
  or g_50369_(_40068_, _40091_, _40092_);
  or g_50370_(_40090_, _40092_, _40093_);
  or g_50371_(_40071_, _40093_, _40094_);
  or g_50372_(_40084_, _40094_, _40095_);
  not g_50373_(_40095_, _40096_);
  xor g_50374_(out[55], out[487], _40097_);
  and g_50375_(_39537_, out[491], _40099_);
  xor g_50376_(out[62], out[494], _40100_);
  xor g_50377_(out[56], out[488], _40101_);
  xor g_50378_(out[49], out[481], _40102_);
  xor g_50379_(out[61], out[493], _40103_);
  xor g_50380_(out[57], out[489], _40104_);
  xor g_50381_(out[52], out[484], _40105_);
  xor g_50382_(out[50], out[482], _40106_);
  and g_50383_(out[59], _39834_, _40107_);
  xor g_50384_(out[51], out[483], _40108_);
  xor g_50385_(out[54], out[486], _40110_);
  xor g_50386_(out[63], out[495], _40111_);
  xor g_50387_(out[58], out[490], _40112_);
  xor g_50388_(out[53], out[485], _40113_);
  xor g_50389_(out[48], out[480], _40114_);
  or g_50390_(_40100_, _40105_, _40115_);
  or g_50391_(_40101_, _40103_, _40116_);
  or g_50392_(_40106_, _40112_, _40117_);
  or g_50393_(_40116_, _40117_, _40118_);
  or g_50394_(_40104_, _40108_, _40119_);
  or g_50395_(_40113_, _40114_, _40121_);
  or g_50396_(_40119_, _40121_, _40122_);
  or g_50397_(_40118_, _40122_, _40123_);
  xor g_50398_(out[60], out[492], _40124_);
  or g_50399_(_40099_, _40124_, _40125_);
  or g_50400_(_40097_, _40110_, _40126_);
  or g_50401_(_40125_, _40126_, _40127_);
  or g_50402_(_40102_, _40107_, _40128_);
  or g_50403_(_40111_, _40128_, _40129_);
  or g_50404_(_40127_, _40129_, _40130_);
  or g_50405_(_40123_, _40130_, _40132_);
  or g_50406_(_40115_, _40132_, _40133_);
  not g_50407_(_40133_, _40134_);
  xor g_50408_(out[42], out[490], _40135_);
  xor g_50409_(out[34], out[482], _40136_);
  xor g_50410_(out[33], out[481], _40137_);
  and g_50411_(_39526_, out[491], _40138_);
  and g_50412_(out[43], _39834_, _40139_);
  xor g_50413_(out[45], out[493], _40140_);
  xor g_50414_(out[35], out[483], _40141_);
  xor g_50415_(out[46], out[494], _40143_);
  xor g_50416_(out[44], out[492], _40144_);
  xor g_50417_(out[40], out[488], _40145_);
  xor g_50418_(out[47], out[495], _40146_);
  xor g_50419_(out[37], out[485], _40147_);
  xor g_50420_(out[38], out[486], _40148_);
  xor g_50421_(out[32], out[480], _40149_);
  xor g_50422_(out[36], out[484], _40150_);
  or g_50423_(_40140_, _40145_, _40151_);
  xor g_50424_(out[41], out[489], _40152_);
  or g_50425_(_40135_, _40136_, _40154_);
  or g_50426_(_40151_, _40154_, _40155_);
  or g_50427_(_40141_, _40152_, _40156_);
  or g_50428_(_40147_, _40156_, _40157_);
  or g_50429_(_40155_, _40157_, _40158_);
  or g_50430_(_40143_, _40150_, _40159_);
  or g_50431_(_40158_, _40159_, _40160_);
  or g_50432_(_40138_, _40144_, _40161_);
  xor g_50433_(out[39], out[487], _40162_);
  or g_50434_(_40148_, _40162_, _40163_);
  or g_50435_(_40161_, _40163_, _40165_);
  or g_50436_(_40137_, _40139_, _40166_);
  or g_50437_(_40146_, _40166_, _40167_);
  or g_50438_(_40165_, _40167_, _40168_);
  or g_50439_(_40149_, _40168_, _40169_);
  or g_50440_(_40160_, _40169_, _40170_);
  not g_50441_(_40170_, _40171_);
  xor g_50442_(out[23], out[487], _40172_);
  and g_50443_(_39493_, out[491], _40173_);
  xor g_50444_(out[30], out[494], _40174_);
  xor g_50445_(out[24], out[488], _40176_);
  xor g_50446_(out[17], out[481], _40177_);
  xor g_50447_(out[29], out[493], _40178_);
  xor g_50448_(out[25], out[489], _40179_);
  xor g_50449_(out[20], out[484], _40180_);
  xor g_50450_(out[18], out[482], _40181_);
  and g_50451_(out[27], _39834_, _40182_);
  xor g_50452_(out[19], out[483], _40183_);
  xor g_50453_(out[22], out[486], _40184_);
  xor g_50454_(out[31], out[495], _40185_);
  xor g_50455_(out[26], out[490], _40187_);
  xor g_50456_(out[21], out[485], _40188_);
  xor g_50457_(out[16], out[480], _40189_);
  or g_50458_(_40174_, _40180_, _40190_);
  or g_50459_(_40176_, _40178_, _40191_);
  or g_50460_(_40181_, _40187_, _40192_);
  or g_50461_(_40191_, _40192_, _40193_);
  or g_50462_(_40179_, _40183_, _40194_);
  or g_50463_(_40188_, _40189_, _40195_);
  or g_50464_(_40194_, _40195_, _40196_);
  or g_50465_(_40193_, _40196_, _40198_);
  xor g_50466_(out[28], out[492], _40199_);
  or g_50467_(_40173_, _40199_, _40200_);
  or g_50468_(_40172_, _40184_, _40201_);
  or g_50469_(_40200_, _40201_, _40202_);
  or g_50470_(_40177_, _40182_, _40203_);
  or g_50471_(_40185_, _40203_, _40204_);
  or g_50472_(_40202_, _40204_, _40205_);
  or g_50473_(_40198_, _40205_, _40206_);
  or g_50474_(_40190_, _40206_, _40207_);
  not g_50475_(_40207_, _40209_);
  and g_50476_(_39438_, out[491], _40210_);
  and g_50477_(out[11], _39834_, _40211_);
  xor g_50478_(out[4], out[484], _40212_);
  xor g_50479_(out[14], out[494], _40213_);
  or g_50480_(_40212_, _40213_, _40214_);
  xor g_50481_(out[13], out[493], _40215_);
  xor g_50482_(out[3], out[483], _40216_);
  xor g_50483_(out[0], out[480], _40217_);
  xor g_50484_(out[10], out[490], _40218_);
  xor g_50485_(out[15], out[495], _40220_);
  xor g_50486_(out[6], out[486], _40221_);
  xor g_50487_(out[5], out[485], _40222_);
  xor g_50488_(out[8], out[488], _40223_);
  or g_50489_(_40215_, _40223_, _40224_);
  xor g_50490_(out[2], out[482], _40225_);
  xor g_50491_(out[9], out[489], _40226_);
  xor g_50492_(out[1], out[481], _40227_);
  or g_50493_(_40218_, _40225_, _40228_);
  or g_50494_(_40224_, _40228_, _40229_);
  or g_50495_(_40216_, _40226_, _40231_);
  or g_50496_(_40222_, _40231_, _40232_);
  or g_50497_(_40229_, _40232_, _40233_);
  or g_50498_(_40214_, _40233_, _40234_);
  xor g_50499_(out[12], out[492], _40235_);
  or g_50500_(_40210_, _40235_, _40236_);
  xor g_50501_(out[7], out[487], _40237_);
  or g_50502_(_40221_, _40237_, _40238_);
  or g_50503_(_40236_, _40238_, _40239_);
  or g_50504_(_40211_, _40227_, _40240_);
  or g_50505_(_40220_, _40240_, _40242_);
  or g_50506_(_40239_, _40242_, _40243_);
  or g_50507_(_40217_, _40243_, _40244_);
  or g_50508_(_40234_, _40244_, _40245_);
  xor g_50509_(out[316], out[476], _40246_);
  and g_50510_(_39724_, out[475], _40247_);
  xor g_50511_(out[312], out[472], _40248_);
  xor g_50512_(out[310], out[470], _40249_);
  xor g_50513_(out[317], out[477], _40250_);
  xor g_50514_(out[318], out[478], _40251_);
  xor g_50515_(out[306], out[466], _40253_);
  xor g_50516_(out[313], out[473], _40254_);
  xor g_50517_(out[309], out[469], _40255_);
  xor g_50518_(out[305], out[465], _40256_);
  and g_50519_(out[315], _39823_, _40257_);
  or g_50520_(_40248_, _40250_, _40258_);
  xor g_50521_(out[319], out[479], _40259_);
  xor g_50522_(out[314], out[474], _40260_);
  xor g_50523_(out[308], out[468], _40261_);
  xor g_50524_(out[307], out[467], _40262_);
  xor g_50525_(out[304], out[464], _40264_);
  or g_50526_(_40253_, _40260_, _40265_);
  or g_50527_(_40258_, _40265_, _40266_);
  or g_50528_(_40254_, _40262_, _40267_);
  or g_50529_(_40255_, _40267_, _40268_);
  or g_50530_(_40266_, _40268_, _40269_);
  or g_50531_(_40251_, _40261_, _40270_);
  or g_50532_(_40269_, _40270_, _40271_);
  or g_50533_(_40246_, _40247_, _40272_);
  xor g_50534_(out[311], out[471], _40273_);
  or g_50535_(_40249_, _40273_, _40275_);
  or g_50536_(_40272_, _40275_, _40276_);
  or g_50537_(_40256_, _40257_, _40277_);
  or g_50538_(_40259_, _40277_, _40278_);
  or g_50539_(_40276_, _40278_, _40279_);
  or g_50540_(_40264_, _40279_, _40280_);
  or g_50541_(_40271_, _40280_, _40281_);
  xor g_50542_(out[295], out[471], _40282_);
  and g_50543_(_39702_, out[475], _40283_);
  xor g_50544_(out[302], out[478], _40284_);
  xor g_50545_(out[296], out[472], _40286_);
  xor g_50546_(out[289], out[465], _40287_);
  xor g_50547_(out[301], out[477], _40288_);
  xor g_50548_(out[297], out[473], _40289_);
  xor g_50549_(out[292], out[468], _40290_);
  xor g_50550_(out[290], out[466], _40291_);
  and g_50551_(out[299], _39823_, _40292_);
  xor g_50552_(out[291], out[467], _40293_);
  xor g_50553_(out[294], out[470], _40294_);
  xor g_50554_(out[303], out[479], _40295_);
  xor g_50555_(out[298], out[474], _40297_);
  xor g_50556_(out[293], out[469], _40298_);
  xor g_50557_(out[288], out[464], _40299_);
  or g_50558_(_40284_, _40290_, _40300_);
  or g_50559_(_40286_, _40288_, _40301_);
  or g_50560_(_40291_, _40297_, _40302_);
  or g_50561_(_40301_, _40302_, _40303_);
  or g_50562_(_40289_, _40293_, _40304_);
  or g_50563_(_40298_, _40299_, _40305_);
  or g_50564_(_40304_, _40305_, _40306_);
  or g_50565_(_40303_, _40306_, _40308_);
  xor g_50566_(out[300], out[476], _40309_);
  or g_50567_(_40283_, _40309_, _40310_);
  or g_50568_(_40282_, _40294_, _40311_);
  or g_50569_(_40310_, _40311_, _40312_);
  or g_50570_(_40287_, _40292_, _40313_);
  or g_50571_(_40295_, _40313_, _40314_);
  or g_50572_(_40312_, _40314_, _40315_);
  or g_50573_(_40308_, _40315_, _40316_);
  or g_50574_(_40300_, _40316_, _40317_);
  not g_50575_(_40317_, _40319_);
  and g_50576_(out[283], _39823_, _40320_);
  xor g_50577_(out[276], out[468], _40321_);
  xor g_50578_(out[286], out[478], _40322_);
  or g_50579_(_40321_, _40322_, _40323_);
  xor g_50580_(out[285], out[477], _40324_);
  xor g_50581_(out[275], out[467], _40325_);
  xor g_50582_(out[272], out[464], _40326_);
  and g_50583_(_39691_, out[475], _40327_);
  xor g_50584_(out[282], out[474], _40328_);
  xor g_50585_(out[287], out[479], _40330_);
  xor g_50586_(out[278], out[470], _40331_);
  xor g_50587_(out[277], out[469], _40332_);
  xor g_50588_(out[280], out[472], _40333_);
  or g_50589_(_40324_, _40333_, _40334_);
  xor g_50590_(out[274], out[466], _40335_);
  xor g_50591_(out[281], out[473], _40336_);
  xor g_50592_(out[273], out[465], _40337_);
  or g_50593_(_40328_, _40335_, _40338_);
  or g_50594_(_40334_, _40338_, _40339_);
  or g_50595_(_40325_, _40336_, _40341_);
  or g_50596_(_40332_, _40341_, _40342_);
  or g_50597_(_40339_, _40342_, _40343_);
  or g_50598_(_40323_, _40343_, _40344_);
  xor g_50599_(out[284], out[476], _40345_);
  or g_50600_(_40327_, _40345_, _40346_);
  xor g_50601_(out[279], out[471], _40347_);
  or g_50602_(_40331_, _40347_, _40348_);
  or g_50603_(_40346_, _40348_, _40349_);
  or g_50604_(_40320_, _40337_, _40350_);
  or g_50605_(_40330_, _40350_, _40352_);
  or g_50606_(_40349_, _40352_, _40353_);
  or g_50607_(_40326_, _40353_, _40354_);
  or g_50608_(_40344_, _40354_, _40355_);
  xor g_50609_(out[263], out[471], _40356_);
  and g_50610_(_39680_, out[475], _40357_);
  xor g_50611_(out[270], out[478], _40358_);
  xor g_50612_(out[264], out[472], _40359_);
  xor g_50613_(out[257], out[465], _40360_);
  xor g_50614_(out[269], out[477], _40361_);
  xor g_50615_(out[265], out[473], _40363_);
  xor g_50616_(out[260], out[468], _40364_);
  xor g_50617_(out[258], out[466], _40365_);
  and g_50618_(out[267], _39823_, _40366_);
  xor g_50619_(out[259], out[467], _40367_);
  xor g_50620_(out[262], out[470], _40368_);
  xor g_50621_(out[271], out[479], _40369_);
  xor g_50622_(out[266], out[474], _40370_);
  xor g_50623_(out[261], out[469], _40371_);
  xor g_50624_(out[256], out[464], _40372_);
  or g_50625_(_40358_, _40364_, _40374_);
  or g_50626_(_40359_, _40361_, _40375_);
  or g_50627_(_40365_, _40370_, _40376_);
  or g_50628_(_40375_, _40376_, _40377_);
  or g_50629_(_40363_, _40367_, _40378_);
  or g_50630_(_40371_, _40372_, _40379_);
  or g_50631_(_40378_, _40379_, _40380_);
  or g_50632_(_40377_, _40380_, _40381_);
  xor g_50633_(out[268], out[476], _40382_);
  or g_50634_(_40357_, _40382_, _40383_);
  or g_50635_(_40356_, _40368_, _40385_);
  or g_50636_(_40383_, _40385_, _40386_);
  or g_50637_(_40360_, _40366_, _40387_);
  or g_50638_(_40369_, _40387_, _40388_);
  or g_50639_(_40386_, _40388_, _40389_);
  or g_50640_(_40381_, _40389_, _40390_);
  or g_50641_(_40374_, _40390_, _40391_);
  xor g_50642_(out[252], out[476], _40392_);
  and g_50643_(_39669_, out[475], _40393_);
  xor g_50644_(out[248], out[472], _40394_);
  xor g_50645_(out[246], out[470], _40396_);
  xor g_50646_(out[253], out[477], _40397_);
  xor g_50647_(out[254], out[478], _40398_);
  xor g_50648_(out[242], out[466], _40399_);
  xor g_50649_(out[249], out[473], _40400_);
  xor g_50650_(out[245], out[469], _40401_);
  xor g_50651_(out[241], out[465], _40402_);
  and g_50652_(out[251], _39823_, _40403_);
  or g_50653_(_40394_, _40397_, _40404_);
  xor g_50654_(out[255], out[479], _40405_);
  xor g_50655_(out[250], out[474], _40407_);
  xor g_50656_(out[244], out[468], _40408_);
  xor g_50657_(out[243], out[467], _40409_);
  xor g_50658_(out[240], out[464], _40410_);
  or g_50659_(_40399_, _40407_, _40411_);
  or g_50660_(_40404_, _40411_, _40412_);
  or g_50661_(_40400_, _40409_, _40413_);
  or g_50662_(_40401_, _40413_, _40414_);
  or g_50663_(_40412_, _40414_, _40415_);
  or g_50664_(_40398_, _40408_, _40416_);
  or g_50665_(_40415_, _40416_, _40418_);
  or g_50666_(_40392_, _40393_, _40419_);
  xor g_50667_(out[247], out[471], _40420_);
  or g_50668_(_40396_, _40420_, _40421_);
  or g_50669_(_40419_, _40421_, _40422_);
  or g_50670_(_40402_, _40403_, _40423_);
  or g_50671_(_40405_, _40423_, _40424_);
  or g_50672_(_40422_, _40424_, _40425_);
  or g_50673_(_40410_, _40425_, _40426_);
  or g_50674_(_40418_, _40426_, _40427_);
  xor g_50675_(out[231], out[471], _40429_);
  and g_50676_(_39658_, out[475], _40430_);
  xor g_50677_(out[238], out[478], _40431_);
  xor g_50678_(out[232], out[472], _40432_);
  xor g_50679_(out[225], out[465], _40433_);
  xor g_50680_(out[237], out[477], _40434_);
  xor g_50681_(out[233], out[473], _40435_);
  xor g_50682_(out[228], out[468], _40436_);
  xor g_50683_(out[226], out[466], _40437_);
  and g_50684_(out[235], _39823_, _40438_);
  xor g_50685_(out[227], out[467], _40440_);
  xor g_50686_(out[230], out[470], _40441_);
  xor g_50687_(out[239], out[479], _40442_);
  xor g_50688_(out[234], out[474], _40443_);
  xor g_50689_(out[229], out[469], _40444_);
  xor g_50690_(out[224], out[464], _40445_);
  or g_50691_(_40431_, _40436_, _40446_);
  or g_50692_(_40432_, _40434_, _40447_);
  or g_50693_(_40437_, _40443_, _40448_);
  or g_50694_(_40447_, _40448_, _40449_);
  or g_50695_(_40435_, _40440_, _40451_);
  or g_50696_(_40444_, _40445_, _40452_);
  or g_50697_(_40451_, _40452_, _40453_);
  or g_50698_(_40449_, _40453_, _40454_);
  xor g_50699_(out[236], out[476], _40455_);
  or g_50700_(_40430_, _40455_, _40456_);
  or g_50701_(_40429_, _40441_, _40457_);
  or g_50702_(_40456_, _40457_, _40458_);
  or g_50703_(_40433_, _40438_, _40459_);
  or g_50704_(_40442_, _40459_, _40460_);
  or g_50705_(_40458_, _40460_, _40462_);
  or g_50706_(_40454_, _40462_, _40463_);
  or g_50707_(_40446_, _40463_, _40464_);
  xor g_50708_(out[209], out[465], _40465_);
  and g_50709_(out[219], _39823_, _40466_);
  xor g_50710_(out[217], out[473], _40467_);
  xor g_50711_(out[208], out[464], _40468_);
  xor g_50712_(out[222], out[478], _40469_);
  xor g_50713_(out[212], out[468], _40470_);
  or g_50714_(_40469_, _40470_, _40471_);
  xor g_50715_(out[221], out[477], _40473_);
  xor g_50716_(out[211], out[467], _40474_);
  and g_50717_(_39647_, out[475], _40475_);
  xor g_50718_(out[214], out[470], _40476_);
  xor g_50719_(out[218], out[474], _40477_);
  xor g_50720_(out[213], out[469], _40478_);
  xor g_50721_(out[223], out[479], _40479_);
  xor g_50722_(out[216], out[472], _40480_);
  or g_50723_(_40473_, _40480_, _40481_);
  xor g_50724_(out[210], out[466], _40482_);
  or g_50725_(_40477_, _40482_, _40484_);
  or g_50726_(_40481_, _40484_, _40485_);
  or g_50727_(_40467_, _40474_, _40486_);
  or g_50728_(_40478_, _40486_, _40487_);
  or g_50729_(_40485_, _40487_, _40488_);
  or g_50730_(_40471_, _40488_, _40489_);
  xor g_50731_(out[220], out[476], _40490_);
  or g_50732_(_40475_, _40490_, _40491_);
  xor g_50733_(out[215], out[471], _40492_);
  or g_50734_(_40476_, _40492_, _40493_);
  or g_50735_(_40491_, _40493_, _40495_);
  or g_50736_(_40465_, _40466_, _40496_);
  or g_50737_(_40479_, _40496_, _40497_);
  or g_50738_(_40495_, _40497_, _40498_);
  or g_50739_(_40468_, _40498_, _40499_);
  or g_50740_(_40489_, _40499_, _40500_);
  xor g_50741_(out[199], out[471], _40501_);
  and g_50742_(_39636_, out[475], _40502_);
  xor g_50743_(out[206], out[478], _40503_);
  xor g_50744_(out[200], out[472], _40504_);
  xor g_50745_(out[193], out[465], _40506_);
  xor g_50746_(out[205], out[477], _40507_);
  xor g_50747_(out[201], out[473], _40508_);
  xor g_50748_(out[196], out[468], _40509_);
  xor g_50749_(out[194], out[466], _40510_);
  and g_50750_(out[203], _39823_, _40511_);
  xor g_50751_(out[195], out[467], _40512_);
  xor g_50752_(out[198], out[470], _40513_);
  xor g_50753_(out[207], out[479], _40514_);
  xor g_50754_(out[202], out[474], _40515_);
  xor g_50755_(out[197], out[469], _40517_);
  xor g_50756_(out[192], out[464], _40518_);
  or g_50757_(_40503_, _40509_, _40519_);
  or g_50758_(_40504_, _40507_, _40520_);
  or g_50759_(_40510_, _40515_, _40521_);
  or g_50760_(_40520_, _40521_, _40522_);
  or g_50761_(_40508_, _40512_, _40523_);
  or g_50762_(_40517_, _40518_, _40524_);
  or g_50763_(_40523_, _40524_, _40525_);
  or g_50764_(_40522_, _40525_, _40526_);
  xor g_50765_(out[204], out[476], _40528_);
  or g_50766_(_40502_, _40528_, _40529_);
  or g_50767_(_40501_, _40513_, _40530_);
  or g_50768_(_40529_, _40530_, _40531_);
  or g_50769_(_40506_, _40511_, _40532_);
  or g_50770_(_40514_, _40532_, _40533_);
  or g_50771_(_40531_, _40533_, _40534_);
  or g_50772_(_40526_, _40534_, _40535_);
  or g_50773_(_40519_, _40535_, _40536_);
  and g_50774_(out[187], _39823_, _40537_);
  xor g_50775_(out[180], out[468], _40539_);
  xor g_50776_(out[190], out[478], _40540_);
  or g_50777_(_40539_, _40540_, _40541_);
  xor g_50778_(out[189], out[477], _40542_);
  xor g_50779_(out[179], out[467], _40543_);
  xor g_50780_(out[176], out[464], _40544_);
  and g_50781_(_39625_, out[475], _40545_);
  xor g_50782_(out[186], out[474], _40546_);
  xor g_50783_(out[191], out[479], _40547_);
  xor g_50784_(out[182], out[470], _40548_);
  xor g_50785_(out[181], out[469], _40550_);
  xor g_50786_(out[184], out[472], _40551_);
  or g_50787_(_40542_, _40551_, _40552_);
  xor g_50788_(out[178], out[466], _40553_);
  xor g_50789_(out[185], out[473], _40554_);
  xor g_50790_(out[177], out[465], _40555_);
  or g_50791_(_40546_, _40553_, _40556_);
  or g_50792_(_40552_, _40556_, _40557_);
  or g_50793_(_40543_, _40554_, _40558_);
  or g_50794_(_40550_, _40558_, _40559_);
  or g_50795_(_40557_, _40559_, _40561_);
  or g_50796_(_40541_, _40561_, _40562_);
  xor g_50797_(out[188], out[476], _40563_);
  or g_50798_(_40545_, _40563_, _40564_);
  xor g_50799_(out[183], out[471], _40565_);
  or g_50800_(_40548_, _40565_, _40566_);
  or g_50801_(_40564_, _40566_, _40567_);
  or g_50802_(_40537_, _40555_, _40568_);
  or g_50803_(_40547_, _40568_, _40569_);
  or g_50804_(_40567_, _40569_, _40570_);
  or g_50805_(_40544_, _40570_, _40572_);
  or g_50806_(_40562_, _40572_, _40573_);
  not g_50807_(_40573_, _40574_);
  xor g_50808_(out[167], out[471], _40575_);
  and g_50809_(_39614_, out[475], _40576_);
  xor g_50810_(out[174], out[478], _40577_);
  xor g_50811_(out[168], out[472], _40578_);
  xor g_50812_(out[161], out[465], _40579_);
  xor g_50813_(out[173], out[477], _40580_);
  xor g_50814_(out[169], out[473], _40581_);
  xor g_50815_(out[164], out[468], _40583_);
  xor g_50816_(out[162], out[466], _40584_);
  and g_50817_(out[171], _39823_, _40585_);
  xor g_50818_(out[163], out[467], _40586_);
  xor g_50819_(out[166], out[470], _40587_);
  xor g_50820_(out[175], out[479], _40588_);
  xor g_50821_(out[170], out[474], _40589_);
  xor g_50822_(out[165], out[469], _40590_);
  xor g_50823_(out[160], out[464], _40591_);
  or g_50824_(_40577_, _40583_, _40592_);
  or g_50825_(_40578_, _40580_, _40594_);
  or g_50826_(_40584_, _40589_, _40595_);
  or g_50827_(_40594_, _40595_, _40596_);
  or g_50828_(_40581_, _40586_, _40597_);
  or g_50829_(_40590_, _40591_, _40598_);
  or g_50830_(_40597_, _40598_, _40599_);
  or g_50831_(_40596_, _40599_, _40600_);
  xor g_50832_(out[172], out[476], _40601_);
  or g_50833_(_40576_, _40601_, _40602_);
  or g_50834_(_40575_, _40587_, _40603_);
  or g_50835_(_40602_, _40603_, _40605_);
  or g_50836_(_40579_, _40585_, _40606_);
  or g_50837_(_40588_, _40606_, _40607_);
  or g_50838_(_40605_, _40607_, _40608_);
  or g_50839_(_40600_, _40608_, _40609_);
  or g_50840_(_40592_, _40609_, _40610_);
  not g_50841_(_40610_, _40611_);
  xor g_50842_(out[145], out[465], _40612_);
  and g_50843_(out[155], _39823_, _40613_);
  xor g_50844_(out[158], out[478], _40614_);
  xor g_50845_(out[147], out[467], _40616_);
  xor g_50846_(out[148], out[468], _40617_);
  xor g_50847_(out[146], out[466], _40618_);
  xor g_50848_(out[153], out[473], _40619_);
  xor g_50849_(out[144], out[464], _40620_);
  and g_50850_(_39603_, out[475], _40621_);
  xor g_50851_(out[150], out[470], _40622_);
  xor g_50852_(out[154], out[474], _40623_);
  xor g_50853_(out[149], out[469], _40624_);
  xor g_50854_(out[159], out[479], _40625_);
  xor g_50855_(out[157], out[477], _40627_);
  xor g_50856_(out[152], out[472], _40628_);
  or g_50857_(_40614_, _40617_, _40629_);
  or g_50858_(_40627_, _40628_, _40630_);
  or g_50859_(_40618_, _40623_, _40631_);
  or g_50860_(_40630_, _40631_, _40632_);
  or g_50861_(_40616_, _40619_, _40633_);
  or g_50862_(_40620_, _40624_, _40634_);
  or g_50863_(_40633_, _40634_, _40635_);
  or g_50864_(_40632_, _40635_, _40636_);
  xor g_50865_(out[156], out[476], _40638_);
  or g_50866_(_40621_, _40638_, _40639_);
  xor g_50867_(out[151], out[471], _40640_);
  or g_50868_(_40622_, _40640_, _40641_);
  or g_50869_(_40639_, _40641_, _40642_);
  or g_50870_(_40612_, _40613_, _40643_);
  or g_50871_(_40625_, _40643_, _40644_);
  or g_50872_(_40642_, _40644_, _40645_);
  or g_50873_(_40636_, _40645_, _40646_);
  or g_50874_(_40629_, _40646_, _40647_);
  xor g_50875_(out[135], out[471], _40649_);
  and g_50876_(_39592_, out[475], _40650_);
  xor g_50877_(out[142], out[478], _40651_);
  xor g_50878_(out[136], out[472], _40652_);
  xor g_50879_(out[129], out[465], _40653_);
  xor g_50880_(out[141], out[477], _40654_);
  xor g_50881_(out[137], out[473], _40655_);
  xor g_50882_(out[132], out[468], _40656_);
  xor g_50883_(out[130], out[466], _40657_);
  and g_50884_(out[139], _39823_, _40658_);
  xor g_50885_(out[131], out[467], _40660_);
  xor g_50886_(out[134], out[470], _40661_);
  xor g_50887_(out[143], out[479], _40662_);
  xor g_50888_(out[138], out[474], _40663_);
  xor g_50889_(out[133], out[469], _40664_);
  xor g_50890_(out[128], out[464], _40665_);
  or g_50891_(_40651_, _40656_, _40666_);
  or g_50892_(_40652_, _40654_, _40667_);
  or g_50893_(_40657_, _40663_, _40668_);
  or g_50894_(_40667_, _40668_, _40669_);
  or g_50895_(_40655_, _40660_, _40671_);
  or g_50896_(_40664_, _40665_, _40672_);
  or g_50897_(_40671_, _40672_, _40673_);
  or g_50898_(_40669_, _40673_, _40674_);
  xor g_50899_(out[140], out[476], _40675_);
  or g_50900_(_40650_, _40675_, _40676_);
  or g_50901_(_40649_, _40661_, _40677_);
  or g_50902_(_40676_, _40677_, _40678_);
  or g_50903_(_40653_, _40658_, _40679_);
  or g_50904_(_40662_, _40679_, _40680_);
  or g_50905_(_40678_, _40680_, _40682_);
  or g_50906_(_40674_, _40682_, _40683_);
  or g_50907_(_40666_, _40683_, _40684_);
  xor g_50908_(out[120], out[472], _40685_);
  xor g_50909_(out[117], out[469], _40686_);
  xor g_50910_(out[115], out[467], _40687_);
  xor g_50911_(out[126], out[478], _40688_);
  xor g_50912_(out[125], out[477], _40689_);
  xor g_50913_(out[114], out[466], _40690_);
  xor g_50914_(out[121], out[473], _40691_);
  xor g_50915_(out[118], out[470], _40693_);
  xor g_50916_(out[127], out[479], _40694_);
  xor g_50917_(out[122], out[474], _40695_);
  xor g_50918_(out[116], out[468], _40696_);
  xor g_50919_(out[112], out[464], _40697_);
  and g_50920_(_39581_, out[475], _40698_);
  and g_50921_(out[123], _39823_, _40699_);
  or g_50922_(_40685_, _40689_, _40700_);
  xor g_50923_(out[113], out[465], _40701_);
  or g_50924_(_40690_, _40695_, _40702_);
  or g_50925_(_40700_, _40702_, _40704_);
  or g_50926_(_40687_, _40691_, _40705_);
  or g_50927_(_40686_, _40705_, _40706_);
  or g_50928_(_40704_, _40706_, _40707_);
  or g_50929_(_40688_, _40696_, _40708_);
  or g_50930_(_40707_, _40708_, _40709_);
  xor g_50931_(out[124], out[476], _40710_);
  or g_50932_(_40698_, _40710_, _40711_);
  xor g_50933_(out[119], out[471], _40712_);
  or g_50934_(_40693_, _40712_, _40713_);
  or g_50935_(_40711_, _40713_, _40715_);
  or g_50936_(_40699_, _40701_, _40716_);
  or g_50937_(_40694_, _40716_, _40717_);
  or g_50938_(_40715_, _40717_, _40718_);
  or g_50939_(_40697_, _40718_, _40719_);
  or g_50940_(_40709_, _40719_, _40720_);
  not g_50941_(_40720_, _40721_);
  xor g_50942_(out[103], out[471], _40722_);
  and g_50943_(_39570_, out[475], _40723_);
  xor g_50944_(out[110], out[478], _40724_);
  xor g_50945_(out[104], out[472], _40726_);
  xor g_50946_(out[97], out[465], _40727_);
  xor g_50947_(out[109], out[477], _40728_);
  xor g_50948_(out[105], out[473], _40729_);
  xor g_50949_(out[100], out[468], _40730_);
  xor g_50950_(out[98], out[466], _40731_);
  and g_50951_(out[107], _39823_, _40732_);
  xor g_50952_(out[99], out[467], _40733_);
  xor g_50953_(out[102], out[470], _40734_);
  xor g_50954_(out[111], out[479], _40735_);
  xor g_50955_(out[106], out[474], _40737_);
  xor g_50956_(out[101], out[469], _40738_);
  xor g_50957_(out[96], out[464], _40739_);
  or g_50958_(_40724_, _40730_, _40740_);
  or g_50959_(_40726_, _40728_, _40741_);
  or g_50960_(_40731_, _40737_, _40742_);
  or g_50961_(_40741_, _40742_, _40743_);
  or g_50962_(_40729_, _40733_, _40744_);
  or g_50963_(_40738_, _40739_, _40745_);
  or g_50964_(_40744_, _40745_, _40746_);
  or g_50965_(_40743_, _40746_, _40748_);
  xor g_50966_(out[108], out[476], _40749_);
  or g_50967_(_40723_, _40749_, _40750_);
  or g_50968_(_40722_, _40734_, _40751_);
  or g_50969_(_40750_, _40751_, _40752_);
  or g_50970_(_40727_, _40732_, _40753_);
  or g_50971_(_40735_, _40753_, _40754_);
  or g_50972_(_40752_, _40754_, _40755_);
  or g_50973_(_40748_, _40755_, _40756_);
  or g_50974_(_40740_, _40756_, _40757_);
  not g_50975_(_40757_, _40759_);
  xor g_50976_(out[81], out[465], _40760_);
  and g_50977_(out[91], _39823_, _40761_);
  xor g_50978_(out[89], out[473], _40762_);
  xor g_50979_(out[80], out[464], _40763_);
  xor g_50980_(out[94], out[478], _40764_);
  xor g_50981_(out[84], out[468], _40765_);
  or g_50982_(_40764_, _40765_, _40766_);
  xor g_50983_(out[93], out[477], _40767_);
  xor g_50984_(out[83], out[467], _40768_);
  and g_50985_(_39559_, out[475], _40770_);
  xor g_50986_(out[86], out[470], _40771_);
  xor g_50987_(out[90], out[474], _40772_);
  xor g_50988_(out[85], out[469], _40773_);
  xor g_50989_(out[95], out[479], _40774_);
  xor g_50990_(out[88], out[472], _40775_);
  or g_50991_(_40767_, _40775_, _40776_);
  xor g_50992_(out[82], out[466], _40777_);
  or g_50993_(_40772_, _40777_, _40778_);
  or g_50994_(_40776_, _40778_, _40779_);
  or g_50995_(_40762_, _40768_, _40781_);
  or g_50996_(_40773_, _40781_, _40782_);
  or g_50997_(_40779_, _40782_, _40783_);
  or g_50998_(_40766_, _40783_, _40784_);
  xor g_50999_(out[92], out[476], _40785_);
  or g_51000_(_40770_, _40785_, _40786_);
  xor g_51001_(out[87], out[471], _40787_);
  or g_51002_(_40771_, _40787_, _40788_);
  or g_51003_(_40786_, _40788_, _40789_);
  or g_51004_(_40760_, _40761_, _40790_);
  or g_51005_(_40774_, _40790_, _40792_);
  or g_51006_(_40789_, _40792_, _40793_);
  or g_51007_(_40763_, _40793_, _40794_);
  or g_51008_(_40784_, _40794_, _40795_);
  xor g_51009_(out[71], out[471], _40796_);
  and g_51010_(_39548_, out[475], _40797_);
  xor g_51011_(out[78], out[478], _40798_);
  xor g_51012_(out[72], out[472], _40799_);
  xor g_51013_(out[65], out[465], _40800_);
  xor g_51014_(out[77], out[477], _40801_);
  xor g_51015_(out[73], out[473], _40803_);
  xor g_51016_(out[68], out[468], _40804_);
  xor g_51017_(out[66], out[466], _40805_);
  and g_51018_(out[75], _39823_, _40806_);
  xor g_51019_(out[67], out[467], _40807_);
  xor g_51020_(out[70], out[470], _40808_);
  xor g_51021_(out[79], out[479], _40809_);
  xor g_51022_(out[74], out[474], _40810_);
  xor g_51023_(out[69], out[469], _40811_);
  xor g_51024_(out[64], out[464], _40812_);
  or g_51025_(_40798_, _40804_, _40814_);
  or g_51026_(_40799_, _40801_, _40815_);
  or g_51027_(_40805_, _40810_, _40816_);
  or g_51028_(_40815_, _40816_, _40817_);
  or g_51029_(_40803_, _40807_, _40818_);
  or g_51030_(_40811_, _40812_, _40819_);
  or g_51031_(_40818_, _40819_, _40820_);
  or g_51032_(_40817_, _40820_, _40821_);
  xor g_51033_(out[76], out[476], _40822_);
  or g_51034_(_40797_, _40822_, _40823_);
  or g_51035_(_40796_, _40808_, _40825_);
  or g_51036_(_40823_, _40825_, _40826_);
  or g_51037_(_40800_, _40806_, _40827_);
  or g_51038_(_40809_, _40827_, _40828_);
  or g_51039_(_40826_, _40828_, _40829_);
  or g_51040_(_40821_, _40829_, _40830_);
  or g_51041_(_40814_, _40830_, _40831_);
  xor g_51042_(out[49], out[465], _40832_);
  and g_51043_(_39537_, out[475], _40833_);
  and g_51044_(out[59], _39823_, _40834_);
  xor g_51045_(out[56], out[472], _40836_);
  xor g_51046_(out[58], out[474], _40837_);
  xor g_51047_(out[50], out[466], _40838_);
  xor g_51048_(out[52], out[468], _40839_);
  xor g_51049_(out[61], out[477], _40840_);
  xor g_51050_(out[57], out[473], _40841_);
  xor g_51051_(out[51], out[467], _40842_);
  xor g_51052_(out[53], out[469], _40843_);
  xor g_51053_(out[62], out[478], _40844_);
  xor g_51054_(out[48], out[464], _40845_);
  xor g_51055_(out[63], out[479], _40847_);
  or g_51056_(_40836_, _40840_, _40848_);
  xor g_51057_(out[54], out[470], _40849_);
  or g_51058_(_40837_, _40838_, _40850_);
  or g_51059_(_40848_, _40850_, _40851_);
  or g_51060_(_40841_, _40842_, _40852_);
  or g_51061_(_40843_, _40852_, _40853_);
  or g_51062_(_40851_, _40853_, _40854_);
  or g_51063_(_40839_, _40844_, _40855_);
  or g_51064_(_40854_, _40855_, _40856_);
  xor g_51065_(out[60], out[476], _40858_);
  or g_51066_(_40833_, _40858_, _40859_);
  xor g_51067_(out[55], out[471], _40860_);
  or g_51068_(_40849_, _40860_, _40861_);
  or g_51069_(_40859_, _40861_, _40862_);
  or g_51070_(_40832_, _40834_, _40863_);
  or g_51071_(_40847_, _40863_, _40864_);
  or g_51072_(_40862_, _40864_, _40865_);
  or g_51073_(_40845_, _40865_, _40866_);
  or g_51074_(_40856_, _40866_, _40867_);
  not g_51075_(_40867_, _40869_);
  xor g_51076_(out[39], out[471], _40870_);
  and g_51077_(_39526_, out[475], _40871_);
  xor g_51078_(out[46], out[478], _40872_);
  xor g_51079_(out[40], out[472], _40873_);
  xor g_51080_(out[33], out[465], _40874_);
  xor g_51081_(out[45], out[477], _40875_);
  xor g_51082_(out[41], out[473], _40876_);
  xor g_51083_(out[36], out[468], _40877_);
  xor g_51084_(out[34], out[466], _40878_);
  and g_51085_(out[43], _39823_, _40880_);
  xor g_51086_(out[35], out[467], _40881_);
  xor g_51087_(out[38], out[470], _40882_);
  xor g_51088_(out[47], out[479], _40883_);
  xor g_51089_(out[42], out[474], _40884_);
  xor g_51090_(out[37], out[469], _40885_);
  xor g_51091_(out[32], out[464], _40886_);
  or g_51092_(_40872_, _40877_, _40887_);
  or g_51093_(_40873_, _40875_, _40888_);
  or g_51094_(_40878_, _40884_, _40889_);
  or g_51095_(_40888_, _40889_, _40891_);
  or g_51096_(_40876_, _40881_, _40892_);
  or g_51097_(_40885_, _40886_, _40893_);
  or g_51098_(_40892_, _40893_, _40894_);
  or g_51099_(_40891_, _40894_, _40895_);
  xor g_51100_(out[44], out[476], _40896_);
  or g_51101_(_40871_, _40896_, _40897_);
  or g_51102_(_40870_, _40882_, _40898_);
  or g_51103_(_40897_, _40898_, _40899_);
  or g_51104_(_40874_, _40880_, _40900_);
  or g_51105_(_40883_, _40900_, _40902_);
  or g_51106_(_40899_, _40902_, _40903_);
  or g_51107_(_40895_, _40903_, _40904_);
  or g_51108_(_40887_, _40904_, _40905_);
  not g_51109_(_40905_, _40906_);
  and g_51110_(out[27], _39823_, _40907_);
  xor g_51111_(out[20], out[468], _40908_);
  xor g_51112_(out[30], out[478], _40909_);
  or g_51113_(_40908_, _40909_, _40910_);
  xor g_51114_(out[29], out[477], _40911_);
  xor g_51115_(out[19], out[467], _40913_);
  xor g_51116_(out[16], out[464], _40914_);
  and g_51117_(_39493_, out[475], _40915_);
  xor g_51118_(out[26], out[474], _40916_);
  xor g_51119_(out[31], out[479], _40917_);
  xor g_51120_(out[22], out[470], _40918_);
  xor g_51121_(out[21], out[469], _40919_);
  xor g_51122_(out[24], out[472], _40920_);
  or g_51123_(_40911_, _40920_, _40921_);
  xor g_51124_(out[18], out[466], _40922_);
  xor g_51125_(out[25], out[473], _40924_);
  xor g_51126_(out[17], out[465], _40925_);
  or g_51127_(_40916_, _40922_, _40926_);
  or g_51128_(_40921_, _40926_, _40927_);
  or g_51129_(_40913_, _40924_, _40928_);
  or g_51130_(_40919_, _40928_, _40929_);
  or g_51131_(_40927_, _40929_, _40930_);
  or g_51132_(_40910_, _40930_, _40931_);
  xor g_51133_(out[28], out[476], _40932_);
  or g_51134_(_40915_, _40932_, _40933_);
  xor g_51135_(out[23], out[471], _40935_);
  or g_51136_(_40918_, _40935_, _40936_);
  or g_51137_(_40933_, _40936_, _40937_);
  or g_51138_(_40907_, _40925_, _40938_);
  or g_51139_(_40917_, _40938_, _40939_);
  or g_51140_(_40937_, _40939_, _40940_);
  or g_51141_(_40914_, _40940_, _40941_);
  or g_51142_(_40931_, _40941_, _40942_);
  xor g_51143_(out[12], out[476], _40943_);
  and g_51144_(_39438_, out[475], _40944_);
  xor g_51145_(out[8], out[472], _40946_);
  xor g_51146_(out[6], out[470], _40947_);
  xor g_51147_(out[13], out[477], _40948_);
  xor g_51148_(out[14], out[478], _40949_);
  xor g_51149_(out[2], out[466], _40950_);
  xor g_51150_(out[9], out[473], _40951_);
  xor g_51151_(out[5], out[469], _40952_);
  xor g_51152_(out[1], out[465], _40953_);
  and g_51153_(out[11], _39823_, _40954_);
  or g_51154_(_40946_, _40948_, _40955_);
  xor g_51155_(out[15], out[479], _40957_);
  xor g_51156_(out[10], out[474], _40958_);
  xor g_51157_(out[4], out[468], _40959_);
  xor g_51158_(out[3], out[467], _40960_);
  xor g_51159_(out[0], out[464], _40961_);
  or g_51160_(_40950_, _40958_, _40962_);
  or g_51161_(_40955_, _40962_, _40963_);
  or g_51162_(_40951_, _40960_, _40964_);
  or g_51163_(_40952_, _40964_, _40965_);
  or g_51164_(_40963_, _40965_, _40966_);
  or g_51165_(_40949_, _40959_, _40968_);
  or g_51166_(_40966_, _40968_, _40969_);
  or g_51167_(_40943_, _40944_, _40970_);
  xor g_51168_(out[7], out[471], _40971_);
  or g_51169_(_40947_, _40971_, _40972_);
  or g_51170_(_40970_, _40972_, _40973_);
  or g_51171_(_40953_, _40954_, _40974_);
  or g_51172_(_40957_, _40974_, _40975_);
  or g_51173_(_40973_, _40975_, _40976_);
  or g_51174_(_40961_, _40976_, _40977_);
  or g_51175_(_40969_, _40977_, _40979_);
  xor g_51176_(out[311], out[455], _40980_);
  and g_51177_(_39724_, out[459], _40981_);
  xor g_51178_(out[318], out[462], _40982_);
  xor g_51179_(out[312], out[456], _40983_);
  xor g_51180_(out[305], out[449], _40984_);
  xor g_51181_(out[317], out[461], _40985_);
  xor g_51182_(out[313], out[457], _40986_);
  xor g_51183_(out[308], out[452], _40987_);
  xor g_51184_(out[306], out[450], _40988_);
  and g_51185_(out[315], _39812_, _40990_);
  xor g_51186_(out[307], out[451], _40991_);
  xor g_51187_(out[310], out[454], _40992_);
  xor g_51188_(out[319], out[463], _40993_);
  xor g_51189_(out[314], out[458], _40994_);
  xor g_51190_(out[309], out[453], _40995_);
  xor g_51191_(out[304], out[448], _40996_);
  or g_51192_(_40982_, _40987_, _40997_);
  or g_51193_(_40983_, _40985_, _40998_);
  or g_51194_(_40988_, _40994_, _40999_);
  or g_51195_(_40998_, _40999_, _41001_);
  or g_51196_(_40986_, _40991_, _41002_);
  or g_51197_(_40995_, _40996_, _41003_);
  or g_51198_(_41002_, _41003_, _41004_);
  or g_51199_(_41001_, _41004_, _41005_);
  xor g_51200_(out[316], out[460], _41006_);
  or g_51201_(_40981_, _41006_, _41007_);
  or g_51202_(_40980_, _40992_, _41008_);
  or g_51203_(_41007_, _41008_, _41009_);
  or g_51204_(_40984_, _40990_, _41010_);
  or g_51205_(_40993_, _41010_, _41012_);
  or g_51206_(_41009_, _41012_, _41013_);
  or g_51207_(_41005_, _41013_, _41014_);
  or g_51208_(_40997_, _41014_, _41015_);
  not g_51209_(_41015_, _41016_);
  xor g_51210_(out[289], out[449], _41017_);
  and g_51211_(out[299], _39812_, _41018_);
  xor g_51212_(out[297], out[457], _41019_);
  xor g_51213_(out[288], out[448], _41020_);
  xor g_51214_(out[302], out[462], _41021_);
  xor g_51215_(out[292], out[452], _41023_);
  or g_51216_(_41021_, _41023_, _41024_);
  xor g_51217_(out[301], out[461], _41025_);
  xor g_51218_(out[291], out[451], _41026_);
  and g_51219_(_39702_, out[459], _41027_);
  xor g_51220_(out[294], out[454], _41028_);
  xor g_51221_(out[298], out[458], _41029_);
  xor g_51222_(out[293], out[453], _41030_);
  xor g_51223_(out[303], out[463], _41031_);
  xor g_51224_(out[296], out[456], _41032_);
  or g_51225_(_41025_, _41032_, _41034_);
  xor g_51226_(out[290], out[450], _41035_);
  or g_51227_(_41029_, _41035_, _41036_);
  or g_51228_(_41034_, _41036_, _41037_);
  or g_51229_(_41019_, _41026_, _41038_);
  or g_51230_(_41030_, _41038_, _41039_);
  or g_51231_(_41037_, _41039_, _41040_);
  or g_51232_(_41024_, _41040_, _41041_);
  xor g_51233_(out[300], out[460], _41042_);
  or g_51234_(_41027_, _41042_, _41043_);
  xor g_51235_(out[295], out[455], _41045_);
  or g_51236_(_41028_, _41045_, _41046_);
  or g_51237_(_41043_, _41046_, _41047_);
  or g_51238_(_41017_, _41018_, _41048_);
  or g_51239_(_41031_, _41048_, _41049_);
  or g_51240_(_41047_, _41049_, _41050_);
  or g_51241_(_41020_, _41050_, _41051_);
  or g_51242_(_41041_, _41051_, _41052_);
  xor g_51243_(out[279], out[455], _41053_);
  and g_51244_(_39691_, out[459], _41054_);
  xor g_51245_(out[286], out[462], _41056_);
  xor g_51246_(out[280], out[456], _41057_);
  xor g_51247_(out[273], out[449], _41058_);
  xor g_51248_(out[285], out[461], _41059_);
  xor g_51249_(out[281], out[457], _41060_);
  xor g_51250_(out[276], out[452], _41061_);
  xor g_51251_(out[274], out[450], _41062_);
  and g_51252_(out[283], _39812_, _41063_);
  xor g_51253_(out[275], out[451], _41064_);
  xor g_51254_(out[278], out[454], _41065_);
  xor g_51255_(out[287], out[463], _41067_);
  xor g_51256_(out[282], out[458], _41068_);
  xor g_51257_(out[277], out[453], _41069_);
  xor g_51258_(out[272], out[448], _41070_);
  or g_51259_(_41056_, _41061_, _41071_);
  or g_51260_(_41057_, _41059_, _41072_);
  or g_51261_(_41062_, _41068_, _41073_);
  or g_51262_(_41072_, _41073_, _41074_);
  or g_51263_(_41060_, _41064_, _41075_);
  or g_51264_(_41069_, _41070_, _41076_);
  or g_51265_(_41075_, _41076_, _41078_);
  or g_51266_(_41074_, _41078_, _41079_);
  xor g_51267_(out[284], out[460], _41080_);
  or g_51268_(_41054_, _41080_, _41081_);
  or g_51269_(_41053_, _41065_, _41082_);
  or g_51270_(_41081_, _41082_, _41083_);
  or g_51271_(_41058_, _41063_, _41084_);
  or g_51272_(_41067_, _41084_, _41085_);
  or g_51273_(_41083_, _41085_, _41086_);
  or g_51274_(_41079_, _41086_, _41087_);
  or g_51275_(_41071_, _41087_, _41089_);
  and g_51276_(out[267], _39812_, _41090_);
  xor g_51277_(out[260], out[452], _41091_);
  xor g_51278_(out[270], out[462], _41092_);
  or g_51279_(_41091_, _41092_, _41093_);
  xor g_51280_(out[269], out[461], _41094_);
  xor g_51281_(out[259], out[451], _41095_);
  xor g_51282_(out[256], out[448], _41096_);
  and g_51283_(_39680_, out[459], _41097_);
  xor g_51284_(out[266], out[458], _41098_);
  xor g_51285_(out[271], out[463], _41100_);
  xor g_51286_(out[262], out[454], _41101_);
  xor g_51287_(out[261], out[453], _41102_);
  xor g_51288_(out[264], out[456], _41103_);
  or g_51289_(_41094_, _41103_, _41104_);
  xor g_51290_(out[258], out[450], _41105_);
  xor g_51291_(out[265], out[457], _41106_);
  xor g_51292_(out[257], out[449], _41107_);
  or g_51293_(_41098_, _41105_, _41108_);
  or g_51294_(_41104_, _41108_, _41109_);
  or g_51295_(_41095_, _41106_, _41111_);
  or g_51296_(_41102_, _41111_, _41112_);
  or g_51297_(_41109_, _41112_, _41113_);
  or g_51298_(_41093_, _41113_, _41114_);
  xor g_51299_(out[268], out[460], _41115_);
  or g_51300_(_41097_, _41115_, _41116_);
  xor g_51301_(out[263], out[455], _41117_);
  or g_51302_(_41101_, _41117_, _41118_);
  or g_51303_(_41116_, _41118_, _41119_);
  or g_51304_(_41090_, _41107_, _41120_);
  or g_51305_(_41100_, _41120_, _41122_);
  or g_51306_(_41119_, _41122_, _41123_);
  or g_51307_(_41096_, _41123_, _41124_);
  or g_51308_(_41114_, _41124_, _41125_);
  xor g_51309_(out[247], out[455], _41126_);
  and g_51310_(_39669_, out[459], _41127_);
  xor g_51311_(out[254], out[462], _41128_);
  xor g_51312_(out[248], out[456], _41129_);
  xor g_51313_(out[241], out[449], _41130_);
  xor g_51314_(out[253], out[461], _41131_);
  xor g_51315_(out[249], out[457], _41133_);
  xor g_51316_(out[244], out[452], _41134_);
  xor g_51317_(out[242], out[450], _41135_);
  and g_51318_(out[251], _39812_, _41136_);
  xor g_51319_(out[243], out[451], _41137_);
  xor g_51320_(out[246], out[454], _41138_);
  xor g_51321_(out[255], out[463], _41139_);
  xor g_51322_(out[250], out[458], _41140_);
  xor g_51323_(out[245], out[453], _41141_);
  xor g_51324_(out[240], out[448], _41142_);
  or g_51325_(_41128_, _41134_, _41144_);
  or g_51326_(_41129_, _41131_, _41145_);
  or g_51327_(_41135_, _41140_, _41146_);
  or g_51328_(_41145_, _41146_, _41147_);
  or g_51329_(_41133_, _41137_, _41148_);
  or g_51330_(_41141_, _41142_, _41149_);
  or g_51331_(_41148_, _41149_, _41150_);
  or g_51332_(_41147_, _41150_, _41151_);
  xor g_51333_(out[252], out[460], _41152_);
  or g_51334_(_41127_, _41152_, _41153_);
  or g_51335_(_41126_, _41138_, _41155_);
  or g_51336_(_41153_, _41155_, _41156_);
  or g_51337_(_41130_, _41136_, _41157_);
  or g_51338_(_41139_, _41157_, _41158_);
  or g_51339_(_41156_, _41158_, _41159_);
  or g_51340_(_41151_, _41159_, _41160_);
  or g_51341_(_41144_, _41160_, _41161_);
  xor g_51342_(out[225], out[449], _41162_);
  and g_51343_(_39658_, out[459], _41163_);
  and g_51344_(out[235], _39812_, _41164_);
  xor g_51345_(out[233], out[457], _41166_);
  xor g_51346_(out[224], out[448], _41167_);
  xor g_51347_(out[238], out[462], _41168_);
  xor g_51348_(out[228], out[452], _41169_);
  or g_51349_(_41168_, _41169_, _41170_);
  xor g_51350_(out[237], out[461], _41171_);
  xor g_51351_(out[227], out[451], _41172_);
  xor g_51352_(out[236], out[460], _41173_);
  xor g_51353_(out[230], out[454], _41174_);
  xor g_51354_(out[234], out[458], _41175_);
  xor g_51355_(out[229], out[453], _41177_);
  xor g_51356_(out[239], out[463], _41178_);
  xor g_51357_(out[232], out[456], _41179_);
  or g_51358_(_41171_, _41179_, _41180_);
  xor g_51359_(out[226], out[450], _41181_);
  or g_51360_(_41175_, _41181_, _41182_);
  or g_51361_(_41180_, _41182_, _41183_);
  or g_51362_(_41166_, _41172_, _41184_);
  or g_51363_(_41177_, _41184_, _41185_);
  or g_51364_(_41183_, _41185_, _41186_);
  or g_51365_(_41170_, _41186_, _41188_);
  or g_51366_(_41163_, _41173_, _41189_);
  xor g_51367_(out[231], out[455], _41190_);
  or g_51368_(_41174_, _41190_, _41191_);
  or g_51369_(_41189_, _41191_, _41192_);
  or g_51370_(_41162_, _41164_, _41193_);
  or g_51371_(_41178_, _41193_, _41194_);
  or g_51372_(_41192_, _41194_, _41195_);
  or g_51373_(_41167_, _41195_, _41196_);
  or g_51374_(_41188_, _41196_, _41197_);
  not g_51375_(_41197_, _41199_);
  xor g_51376_(out[215], out[455], _41200_);
  and g_51377_(_39647_, out[459], _41201_);
  xor g_51378_(out[222], out[462], _41202_);
  xor g_51379_(out[216], out[456], _41203_);
  xor g_51380_(out[209], out[449], _41204_);
  xor g_51381_(out[221], out[461], _41205_);
  xor g_51382_(out[217], out[457], _41206_);
  xor g_51383_(out[212], out[452], _41207_);
  xor g_51384_(out[210], out[450], _41208_);
  and g_51385_(out[219], _39812_, _41210_);
  xor g_51386_(out[211], out[451], _41211_);
  xor g_51387_(out[214], out[454], _41212_);
  xor g_51388_(out[223], out[463], _41213_);
  xor g_51389_(out[218], out[458], _41214_);
  xor g_51390_(out[213], out[453], _41215_);
  xor g_51391_(out[208], out[448], _41216_);
  or g_51392_(_41202_, _41207_, _41217_);
  or g_51393_(_41203_, _41205_, _41218_);
  or g_51394_(_41208_, _41214_, _41219_);
  or g_51395_(_41218_, _41219_, _41221_);
  or g_51396_(_41206_, _41211_, _41222_);
  or g_51397_(_41215_, _41216_, _41223_);
  or g_51398_(_41222_, _41223_, _41224_);
  or g_51399_(_41221_, _41224_, _41225_);
  xor g_51400_(out[220], out[460], _41226_);
  or g_51401_(_41201_, _41226_, _41227_);
  or g_51402_(_41200_, _41212_, _41228_);
  or g_51403_(_41227_, _41228_, _41229_);
  or g_51404_(_41204_, _41210_, _41230_);
  or g_51405_(_41213_, _41230_, _41232_);
  or g_51406_(_41229_, _41232_, _41233_);
  or g_51407_(_41225_, _41233_, _41234_);
  or g_51408_(_41217_, _41234_, _41235_);
  not g_51409_(_41235_, _41236_);
  xor g_51410_(out[193], out[449], _41237_);
  and g_51411_(out[203], _39812_, _41238_);
  xor g_51412_(out[201], out[457], _41239_);
  xor g_51413_(out[192], out[448], _41240_);
  xor g_51414_(out[206], out[462], _41241_);
  xor g_51415_(out[196], out[452], _41243_);
  or g_51416_(_41241_, _41243_, _41244_);
  xor g_51417_(out[205], out[461], _41245_);
  xor g_51418_(out[195], out[451], _41246_);
  and g_51419_(_39636_, out[459], _41247_);
  xor g_51420_(out[198], out[454], _41248_);
  xor g_51421_(out[202], out[458], _41249_);
  xor g_51422_(out[197], out[453], _41250_);
  xor g_51423_(out[207], out[463], _41251_);
  xor g_51424_(out[200], out[456], _41252_);
  or g_51425_(_41245_, _41252_, _41254_);
  xor g_51426_(out[194], out[450], _41255_);
  or g_51427_(_41249_, _41255_, _41256_);
  or g_51428_(_41254_, _41256_, _41257_);
  or g_51429_(_41239_, _41246_, _41258_);
  or g_51430_(_41250_, _41258_, _41259_);
  or g_51431_(_41257_, _41259_, _41260_);
  or g_51432_(_41244_, _41260_, _41261_);
  xor g_51433_(out[204], out[460], _41262_);
  or g_51434_(_41247_, _41262_, _41263_);
  xor g_51435_(out[199], out[455], _41265_);
  or g_51436_(_41248_, _41265_, _41266_);
  or g_51437_(_41263_, _41266_, _41267_);
  or g_51438_(_41237_, _41238_, _41268_);
  or g_51439_(_41251_, _41268_, _41269_);
  or g_51440_(_41267_, _41269_, _41270_);
  or g_51441_(_41240_, _41270_, _41271_);
  or g_51442_(_41261_, _41271_, _41272_);
  xor g_51443_(out[183], out[455], _41273_);
  and g_51444_(_39625_, out[459], _41274_);
  xor g_51445_(out[190], out[462], _41276_);
  xor g_51446_(out[184], out[456], _41277_);
  xor g_51447_(out[177], out[449], _41278_);
  xor g_51448_(out[189], out[461], _41279_);
  xor g_51449_(out[185], out[457], _41280_);
  xor g_51450_(out[180], out[452], _41281_);
  xor g_51451_(out[178], out[450], _41282_);
  and g_51452_(out[187], _39812_, _41283_);
  xor g_51453_(out[179], out[451], _41284_);
  xor g_51454_(out[182], out[454], _41285_);
  xor g_51455_(out[191], out[463], _41287_);
  xor g_51456_(out[186], out[458], _41288_);
  xor g_51457_(out[181], out[453], _41289_);
  xor g_51458_(out[176], out[448], _41290_);
  or g_51459_(_41276_, _41281_, _41291_);
  or g_51460_(_41277_, _41279_, _41292_);
  or g_51461_(_41282_, _41288_, _41293_);
  or g_51462_(_41292_, _41293_, _41294_);
  or g_51463_(_41280_, _41284_, _41295_);
  or g_51464_(_41289_, _41290_, _41296_);
  or g_51465_(_41295_, _41296_, _41298_);
  or g_51466_(_41294_, _41298_, _41299_);
  xor g_51467_(out[188], out[460], _41300_);
  or g_51468_(_41274_, _41300_, _41301_);
  or g_51469_(_41273_, _41285_, _41302_);
  or g_51470_(_41301_, _41302_, _41303_);
  or g_51471_(_41278_, _41283_, _41304_);
  or g_51472_(_41287_, _41304_, _41305_);
  or g_51473_(_41303_, _41305_, _41306_);
  or g_51474_(_41299_, _41306_, _41307_);
  or g_51475_(_41291_, _41307_, _41309_);
  xor g_51476_(out[161], out[449], _41310_);
  and g_51477_(_39614_, out[459], _41311_);
  and g_51478_(out[171], _39812_, _41312_);
  xor g_51479_(out[169], out[457], _41313_);
  xor g_51480_(out[160], out[448], _41314_);
  xor g_51481_(out[174], out[462], _41315_);
  xor g_51482_(out[164], out[452], _41316_);
  or g_51483_(_41315_, _41316_, _41317_);
  xor g_51484_(out[173], out[461], _41318_);
  xor g_51485_(out[163], out[451], _41320_);
  xor g_51486_(out[172], out[460], _41321_);
  xor g_51487_(out[166], out[454], _41322_);
  xor g_51488_(out[170], out[458], _41323_);
  xor g_51489_(out[165], out[453], _41324_);
  xor g_51490_(out[175], out[463], _41325_);
  xor g_51491_(out[168], out[456], _41326_);
  or g_51492_(_41318_, _41326_, _41327_);
  xor g_51493_(out[162], out[450], _41328_);
  or g_51494_(_41323_, _41328_, _41329_);
  or g_51495_(_41327_, _41329_, _41331_);
  or g_51496_(_41313_, _41320_, _41332_);
  or g_51497_(_41324_, _41332_, _41333_);
  or g_51498_(_41331_, _41333_, _41334_);
  or g_51499_(_41317_, _41334_, _41335_);
  or g_51500_(_41311_, _41321_, _41336_);
  xor g_51501_(out[167], out[455], _41337_);
  or g_51502_(_41322_, _41337_, _41338_);
  or g_51503_(_41336_, _41338_, _41339_);
  or g_51504_(_41310_, _41312_, _41340_);
  or g_51505_(_41325_, _41340_, _41342_);
  or g_51506_(_41339_, _41342_, _41343_);
  or g_51507_(_41314_, _41343_, _41344_);
  or g_51508_(_41335_, _41344_, _41345_);
  not g_51509_(_41345_, _41346_);
  xor g_51510_(out[151], out[455], _41347_);
  and g_51511_(_39603_, out[459], _41348_);
  xor g_51512_(out[158], out[462], _41349_);
  xor g_51513_(out[152], out[456], _41350_);
  xor g_51514_(out[145], out[449], _41351_);
  xor g_51515_(out[157], out[461], _41353_);
  xor g_51516_(out[153], out[457], _41354_);
  xor g_51517_(out[148], out[452], _41355_);
  xor g_51518_(out[146], out[450], _41356_);
  and g_51519_(out[155], _39812_, _41357_);
  xor g_51520_(out[147], out[451], _41358_);
  xor g_51521_(out[150], out[454], _41359_);
  xor g_51522_(out[159], out[463], _41360_);
  xor g_51523_(out[154], out[458], _41361_);
  xor g_51524_(out[149], out[453], _41362_);
  xor g_51525_(out[144], out[448], _41364_);
  or g_51526_(_41349_, _41355_, _41365_);
  or g_51527_(_41350_, _41353_, _41366_);
  or g_51528_(_41356_, _41361_, _41367_);
  or g_51529_(_41366_, _41367_, _41368_);
  or g_51530_(_41354_, _41358_, _41369_);
  or g_51531_(_41362_, _41364_, _41370_);
  or g_51532_(_41369_, _41370_, _41371_);
  or g_51533_(_41368_, _41371_, _41372_);
  xor g_51534_(out[156], out[460], _41373_);
  or g_51535_(_41348_, _41373_, _41375_);
  or g_51536_(_41347_, _41359_, _41376_);
  or g_51537_(_41375_, _41376_, _41377_);
  or g_51538_(_41351_, _41357_, _41378_);
  or g_51539_(_41360_, _41378_, _41379_);
  or g_51540_(_41377_, _41379_, _41380_);
  or g_51541_(_41372_, _41380_, _41381_);
  or g_51542_(_41365_, _41381_, _41382_);
  not g_51543_(_41382_, _41383_);
  and g_51544_(out[139], _39812_, _41384_);
  xor g_51545_(out[132], out[452], _41386_);
  xor g_51546_(out[142], out[462], _41387_);
  or g_51547_(_41386_, _41387_, _41388_);
  xor g_51548_(out[141], out[461], _41389_);
  xor g_51549_(out[131], out[451], _41390_);
  xor g_51550_(out[128], out[448], _41391_);
  and g_51551_(_39592_, out[459], _41392_);
  xor g_51552_(out[138], out[458], _41393_);
  xor g_51553_(out[143], out[463], _41394_);
  xor g_51554_(out[134], out[454], _41395_);
  xor g_51555_(out[133], out[453], _41397_);
  xor g_51556_(out[136], out[456], _41398_);
  or g_51557_(_41389_, _41398_, _41399_);
  xor g_51558_(out[130], out[450], _41400_);
  xor g_51559_(out[137], out[457], _41401_);
  xor g_51560_(out[129], out[449], _41402_);
  or g_51561_(_41393_, _41400_, _41403_);
  or g_51562_(_41399_, _41403_, _41404_);
  or g_51563_(_41390_, _41401_, _41405_);
  or g_51564_(_41397_, _41405_, _41406_);
  or g_51565_(_41404_, _41406_, _41408_);
  or g_51566_(_41388_, _41408_, _41409_);
  xor g_51567_(out[140], out[460], _41410_);
  or g_51568_(_41392_, _41410_, _41411_);
  xor g_51569_(out[135], out[455], _41412_);
  or g_51570_(_41395_, _41412_, _41413_);
  or g_51571_(_41411_, _41413_, _41414_);
  or g_51572_(_41384_, _41402_, _41415_);
  or g_51573_(_41394_, _41415_, _41416_);
  or g_51574_(_41414_, _41416_, _41417_);
  or g_51575_(_41391_, _41417_, _41419_);
  or g_51576_(_41409_, _41419_, _41420_);
  xor g_51577_(out[119], out[455], _41421_);
  and g_51578_(_39581_, out[459], _41422_);
  xor g_51579_(out[126], out[462], _41423_);
  xor g_51580_(out[120], out[456], _41424_);
  xor g_51581_(out[113], out[449], _41425_);
  xor g_51582_(out[125], out[461], _41426_);
  xor g_51583_(out[121], out[457], _41427_);
  xor g_51584_(out[116], out[452], _41428_);
  xor g_51585_(out[114], out[450], _41430_);
  and g_51586_(out[123], _39812_, _41431_);
  xor g_51587_(out[115], out[451], _41432_);
  xor g_51588_(out[118], out[454], _41433_);
  xor g_51589_(out[127], out[463], _41434_);
  xor g_51590_(out[122], out[458], _41435_);
  xor g_51591_(out[117], out[453], _41436_);
  xor g_51592_(out[112], out[448], _41437_);
  or g_51593_(_41423_, _41428_, _41438_);
  or g_51594_(_41424_, _41426_, _41439_);
  or g_51595_(_41430_, _41435_, _41441_);
  or g_51596_(_41439_, _41441_, _41442_);
  or g_51597_(_41427_, _41432_, _41443_);
  or g_51598_(_41436_, _41437_, _41444_);
  or g_51599_(_41443_, _41444_, _41445_);
  or g_51600_(_41442_, _41445_, _41446_);
  xor g_51601_(out[124], out[460], _41447_);
  or g_51602_(_41422_, _41447_, _41448_);
  or g_51603_(_41421_, _41433_, _41449_);
  or g_51604_(_41448_, _41449_, _41450_);
  or g_51605_(_41425_, _41431_, _41452_);
  or g_51606_(_41434_, _41452_, _41453_);
  or g_51607_(_41450_, _41453_, _41454_);
  or g_51608_(_41446_, _41454_, _41455_);
  or g_51609_(_41438_, _41455_, _41456_);
  and g_51610_(out[107], _39812_, _41457_);
  xor g_51611_(out[100], out[452], _41458_);
  xor g_51612_(out[110], out[462], _41459_);
  or g_51613_(_41458_, _41459_, _41460_);
  xor g_51614_(out[109], out[461], _41461_);
  xor g_51615_(out[99], out[451], _41463_);
  xor g_51616_(out[96], out[448], _41464_);
  and g_51617_(_39570_, out[459], _41465_);
  xor g_51618_(out[106], out[458], _41466_);
  xor g_51619_(out[111], out[463], _41467_);
  xor g_51620_(out[102], out[454], _41468_);
  xor g_51621_(out[101], out[453], _41469_);
  xor g_51622_(out[104], out[456], _41470_);
  or g_51623_(_41461_, _41470_, _41471_);
  xor g_51624_(out[98], out[450], _41472_);
  xor g_51625_(out[105], out[457], _41474_);
  xor g_51626_(out[97], out[449], _41475_);
  or g_51627_(_41466_, _41472_, _41476_);
  or g_51628_(_41471_, _41476_, _41477_);
  or g_51629_(_41463_, _41474_, _41478_);
  or g_51630_(_41469_, _41478_, _41479_);
  or g_51631_(_41477_, _41479_, _41480_);
  or g_51632_(_41460_, _41480_, _41481_);
  xor g_51633_(out[108], out[460], _41482_);
  or g_51634_(_41465_, _41482_, _41483_);
  xor g_51635_(out[103], out[455], _41485_);
  or g_51636_(_41468_, _41485_, _41486_);
  or g_51637_(_41483_, _41486_, _41487_);
  or g_51638_(_41457_, _41475_, _41488_);
  or g_51639_(_41467_, _41488_, _41489_);
  or g_51640_(_41487_, _41489_, _41490_);
  or g_51641_(_41464_, _41490_, _41491_);
  or g_51642_(_41481_, _41491_, _41492_);
  xor g_51643_(out[87], out[455], _41493_);
  and g_51644_(_39559_, out[459], _41494_);
  xor g_51645_(out[94], out[462], _41496_);
  xor g_51646_(out[88], out[456], _41497_);
  xor g_51647_(out[81], out[449], _41498_);
  xor g_51648_(out[93], out[461], _41499_);
  xor g_51649_(out[89], out[457], _41500_);
  xor g_51650_(out[84], out[452], _41501_);
  xor g_51651_(out[82], out[450], _41502_);
  and g_51652_(out[91], _39812_, _41503_);
  xor g_51653_(out[83], out[451], _41504_);
  xor g_51654_(out[86], out[454], _41505_);
  xor g_51655_(out[95], out[463], _41507_);
  xor g_51656_(out[90], out[458], _41508_);
  xor g_51657_(out[85], out[453], _41509_);
  xor g_51658_(out[80], out[448], _41510_);
  or g_51659_(_41496_, _41501_, _41511_);
  or g_51660_(_41497_, _41499_, _41512_);
  or g_51661_(_41502_, _41508_, _41513_);
  or g_51662_(_41512_, _41513_, _41514_);
  or g_51663_(_41500_, _41504_, _41515_);
  or g_51664_(_41509_, _41510_, _41516_);
  or g_51665_(_41515_, _41516_, _41518_);
  or g_51666_(_41514_, _41518_, _41519_);
  xor g_51667_(out[92], out[460], _41520_);
  or g_51668_(_41494_, _41520_, _41521_);
  or g_51669_(_41493_, _41505_, _41522_);
  or g_51670_(_41521_, _41522_, _41523_);
  or g_51671_(_41498_, _41503_, _41524_);
  or g_51672_(_41507_, _41524_, _41525_);
  or g_51673_(_41523_, _41525_, _41526_);
  or g_51674_(_41519_, _41526_, _41527_);
  or g_51675_(_41511_, _41527_, _41529_);
  xor g_51676_(out[65], out[449], _41530_);
  and g_51677_(_39548_, out[459], _41531_);
  and g_51678_(out[75], _39812_, _41532_);
  xor g_51679_(out[73], out[457], _41533_);
  xor g_51680_(out[64], out[448], _41534_);
  xor g_51681_(out[78], out[462], _41535_);
  xor g_51682_(out[68], out[452], _41536_);
  or g_51683_(_41535_, _41536_, _41537_);
  xor g_51684_(out[77], out[461], _41538_);
  xor g_51685_(out[67], out[451], _41540_);
  xor g_51686_(out[76], out[460], _41541_);
  xor g_51687_(out[70], out[454], _41542_);
  xor g_51688_(out[74], out[458], _41543_);
  xor g_51689_(out[69], out[453], _41544_);
  xor g_51690_(out[79], out[463], _41545_);
  xor g_51691_(out[72], out[456], _41546_);
  or g_51692_(_41538_, _41546_, _41547_);
  xor g_51693_(out[66], out[450], _41548_);
  or g_51694_(_41543_, _41548_, _41549_);
  or g_51695_(_41547_, _41549_, _41551_);
  or g_51696_(_41533_, _41540_, _41552_);
  or g_51697_(_41544_, _41552_, _41553_);
  or g_51698_(_41551_, _41553_, _41554_);
  or g_51699_(_41537_, _41554_, _41555_);
  or g_51700_(_41531_, _41541_, _41556_);
  xor g_51701_(out[71], out[455], _41557_);
  or g_51702_(_41542_, _41557_, _41558_);
  or g_51703_(_41556_, _41558_, _41559_);
  or g_51704_(_41530_, _41532_, _41560_);
  or g_51705_(_41545_, _41560_, _41562_);
  or g_51706_(_41559_, _41562_, _41563_);
  or g_51707_(_41534_, _41563_, _41564_);
  or g_51708_(_41555_, _41564_, _41565_);
  not g_51709_(_41565_, _41566_);
  xor g_51710_(out[55], out[455], _41567_);
  and g_51711_(_39537_, out[459], _41568_);
  xor g_51712_(out[62], out[462], _41569_);
  xor g_51713_(out[56], out[456], _41570_);
  xor g_51714_(out[49], out[449], _41571_);
  xor g_51715_(out[61], out[461], _41573_);
  xor g_51716_(out[57], out[457], _41574_);
  xor g_51717_(out[52], out[452], _41575_);
  xor g_51718_(out[50], out[450], _41576_);
  and g_51719_(out[59], _39812_, _41577_);
  xor g_51720_(out[51], out[451], _41578_);
  xor g_51721_(out[54], out[454], _41579_);
  xor g_51722_(out[63], out[463], _41580_);
  xor g_51723_(out[58], out[458], _41581_);
  xor g_51724_(out[53], out[453], _41582_);
  xor g_51725_(out[48], out[448], _41584_);
  or g_51726_(_41569_, _41575_, _41585_);
  or g_51727_(_41570_, _41573_, _41586_);
  or g_51728_(_41576_, _41581_, _41587_);
  or g_51729_(_41586_, _41587_, _41588_);
  or g_51730_(_41574_, _41578_, _41589_);
  or g_51731_(_41582_, _41584_, _41590_);
  or g_51732_(_41589_, _41590_, _41591_);
  or g_51733_(_41588_, _41591_, _41592_);
  xor g_51734_(out[60], out[460], _41593_);
  or g_51735_(_41568_, _41593_, _41595_);
  or g_51736_(_41567_, _41579_, _41596_);
  or g_51737_(_41595_, _41596_, _41597_);
  or g_51738_(_41571_, _41577_, _41598_);
  or g_51739_(_41580_, _41598_, _41599_);
  or g_51740_(_41597_, _41599_, _41600_);
  or g_51741_(_41592_, _41600_, _41601_);
  or g_51742_(_41585_, _41601_, _41602_);
  not g_51743_(_41602_, _41603_);
  and g_51744_(out[43], _39812_, _41604_);
  and g_51745_(_39526_, out[459], _41606_);
  xor g_51746_(out[35], out[451], _41607_);
  xor g_51747_(out[33], out[449], _41608_);
  xor g_51748_(out[46], out[462], _41609_);
  xor g_51749_(out[37], out[453], _41610_);
  xor g_51750_(out[40], out[456], _41611_);
  xor g_51751_(out[42], out[458], _41612_);
  xor g_51752_(out[38], out[454], _41613_);
  xor g_51753_(out[36], out[452], _41614_);
  xor g_51754_(out[45], out[461], _41615_);
  xor g_51755_(out[47], out[463], _41617_);
  xor g_51756_(out[32], out[448], _41618_);
  xor g_51757_(out[34], out[450], _41619_);
  xor g_51758_(out[41], out[457], _41620_);
  or g_51759_(_41609_, _41614_, _41621_);
  or g_51760_(_41611_, _41615_, _41622_);
  or g_51761_(_41612_, _41619_, _41623_);
  or g_51762_(_41622_, _41623_, _41624_);
  or g_51763_(_41607_, _41620_, _41625_);
  or g_51764_(_41610_, _41618_, _41626_);
  or g_51765_(_41625_, _41626_, _41628_);
  or g_51766_(_41624_, _41628_, _41629_);
  xor g_51767_(out[44], out[460], _41630_);
  or g_51768_(_41606_, _41630_, _41631_);
  xor g_51769_(out[39], out[455], _41632_);
  or g_51770_(_41613_, _41632_, _41633_);
  or g_51771_(_41631_, _41633_, _41634_);
  or g_51772_(_41604_, _41608_, _41635_);
  or g_51773_(_41617_, _41635_, _41636_);
  or g_51774_(_41634_, _41636_, _41637_);
  or g_51775_(_41629_, _41637_, _41639_);
  or g_51776_(_41621_, _41639_, _41640_);
  xor g_51777_(out[23], out[455], _41641_);
  and g_51778_(_39493_, out[459], _41642_);
  xor g_51779_(out[30], out[462], _41643_);
  xor g_51780_(out[24], out[456], _41644_);
  xor g_51781_(out[17], out[449], _41645_);
  xor g_51782_(out[29], out[461], _41646_);
  xor g_51783_(out[25], out[457], _41647_);
  xor g_51784_(out[20], out[452], _41648_);
  xor g_51785_(out[18], out[450], _41650_);
  and g_51786_(out[27], _39812_, _41651_);
  xor g_51787_(out[19], out[451], _41652_);
  xor g_51788_(out[22], out[454], _41653_);
  xor g_51789_(out[31], out[463], _41654_);
  xor g_51790_(out[26], out[458], _41655_);
  xor g_51791_(out[21], out[453], _41656_);
  xor g_51792_(out[16], out[448], _41657_);
  or g_51793_(_41643_, _41648_, _41658_);
  or g_51794_(_41644_, _41646_, _41659_);
  or g_51795_(_41650_, _41655_, _41661_);
  or g_51796_(_41659_, _41661_, _41662_);
  or g_51797_(_41647_, _41652_, _41663_);
  or g_51798_(_41656_, _41657_, _41664_);
  or g_51799_(_41663_, _41664_, _41665_);
  or g_51800_(_41662_, _41665_, _41666_);
  xor g_51801_(out[28], out[460], _41667_);
  or g_51802_(_41642_, _41667_, _41668_);
  or g_51803_(_41641_, _41653_, _41669_);
  or g_51804_(_41668_, _41669_, _41670_);
  or g_51805_(_41645_, _41651_, _41672_);
  or g_51806_(_41654_, _41672_, _41673_);
  or g_51807_(_41670_, _41673_, _41674_);
  or g_51808_(_41666_, _41674_, _41675_);
  or g_51809_(_41658_, _41675_, _41676_);
  xor g_51810_(out[12], out[460], _41677_);
  and g_51811_(_39438_, out[459], _41678_);
  xor g_51812_(out[8], out[456], _41679_);
  xor g_51813_(out[6], out[454], _41680_);
  xor g_51814_(out[13], out[461], _41681_);
  xor g_51815_(out[14], out[462], _41683_);
  xor g_51816_(out[2], out[450], _41684_);
  xor g_51817_(out[9], out[457], _41685_);
  xor g_51818_(out[5], out[453], _41686_);
  xor g_51819_(out[1], out[449], _41687_);
  and g_51820_(out[11], _39812_, _41688_);
  or g_51821_(_41679_, _41681_, _41689_);
  xor g_51822_(out[15], out[463], _41690_);
  xor g_51823_(out[10], out[458], _41691_);
  xor g_51824_(out[4], out[452], _41692_);
  xor g_51825_(out[3], out[451], _41694_);
  xor g_51826_(out[0], out[448], _41695_);
  or g_51827_(_41684_, _41691_, _41696_);
  or g_51828_(_41689_, _41696_, _41697_);
  or g_51829_(_41685_, _41694_, _41698_);
  or g_51830_(_41686_, _41698_, _41699_);
  or g_51831_(_41697_, _41699_, _41700_);
  or g_51832_(_41683_, _41692_, _41701_);
  or g_51833_(_41700_, _41701_, _41702_);
  or g_51834_(_41677_, _41678_, _41703_);
  xor g_51835_(out[7], out[455], _41705_);
  or g_51836_(_41680_, _41705_, _41706_);
  or g_51837_(_41703_, _41706_, _41707_);
  or g_51838_(_41687_, _41688_, _41708_);
  or g_51839_(_41690_, _41708_, _41709_);
  or g_51840_(_41707_, _41709_, _41710_);
  or g_51841_(_41695_, _41710_, _41711_);
  or g_51842_(_41702_, _41711_, _41712_);
  xor g_51843_(out[307], out[435], _41713_);
  xor g_51844_(out[308], out[436], _41714_);
  xor g_51845_(out[318], out[446], _41716_);
  xor g_51846_(out[306], out[434], _41717_);
  xor g_51847_(out[309], out[437], _41718_);
  xor g_51848_(out[313], out[441], _41719_);
  xor g_51849_(out[312], out[440], _41720_);
  xor g_51850_(out[319], out[447], _41721_);
  xor g_51851_(out[314], out[442], _41722_);
  xor g_51852_(out[310], out[438], _41723_);
  xor g_51853_(out[304], out[432], _41724_);
  and g_51854_(_39724_, out[443], _41725_);
  and g_51855_(out[315], _39801_, _41727_);
  xor g_51856_(out[317], out[445], _41728_);
  or g_51857_(_41720_, _41728_, _41729_);
  xor g_51858_(out[305], out[433], _41730_);
  or g_51859_(_41717_, _41722_, _41731_);
  or g_51860_(_41729_, _41731_, _41732_);
  or g_51861_(_41713_, _41719_, _41733_);
  or g_51862_(_41718_, _41733_, _41734_);
  or g_51863_(_41732_, _41734_, _41735_);
  or g_51864_(_41714_, _41716_, _41736_);
  or g_51865_(_41735_, _41736_, _41738_);
  xor g_51866_(out[316], out[444], _41739_);
  or g_51867_(_41725_, _41739_, _41740_);
  xor g_51868_(out[311], out[439], _41741_);
  or g_51869_(_41723_, _41741_, _41742_);
  or g_51870_(_41740_, _41742_, _41743_);
  or g_51871_(_41727_, _41730_, _41744_);
  or g_51872_(_41721_, _41744_, _41745_);
  or g_51873_(_41743_, _41745_, _41746_);
  or g_51874_(_41724_, _41746_, _41747_);
  or g_51875_(_41738_, _41747_, _41749_);
  xor g_51876_(out[295], out[439], _41750_);
  and g_51877_(_39702_, out[443], _41751_);
  xor g_51878_(out[302], out[446], _41752_);
  xor g_51879_(out[296], out[440], _41753_);
  xor g_51880_(out[289], out[433], _41754_);
  xor g_51881_(out[301], out[445], _41755_);
  xor g_51882_(out[297], out[441], _41756_);
  xor g_51883_(out[292], out[436], _41757_);
  xor g_51884_(out[290], out[434], _41758_);
  and g_51885_(out[299], _39801_, _41760_);
  xor g_51886_(out[291], out[435], _41761_);
  xor g_51887_(out[294], out[438], _41762_);
  xor g_51888_(out[303], out[447], _41763_);
  xor g_51889_(out[298], out[442], _41764_);
  xor g_51890_(out[293], out[437], _41765_);
  xor g_51891_(out[288], out[432], _41766_);
  or g_51892_(_41752_, _41757_, _41767_);
  or g_51893_(_41753_, _41755_, _41768_);
  or g_51894_(_41758_, _41764_, _41769_);
  or g_51895_(_41768_, _41769_, _41771_);
  or g_51896_(_41756_, _41761_, _41772_);
  or g_51897_(_41765_, _41766_, _41773_);
  or g_51898_(_41772_, _41773_, _41774_);
  or g_51899_(_41771_, _41774_, _41775_);
  xor g_51900_(out[300], out[444], _41776_);
  or g_51901_(_41751_, _41776_, _41777_);
  or g_51902_(_41750_, _41762_, _41778_);
  or g_51903_(_41777_, _41778_, _41779_);
  or g_51904_(_41754_, _41760_, _41780_);
  or g_51905_(_41763_, _41780_, _41782_);
  or g_51906_(_41779_, _41782_, _41783_);
  or g_51907_(_41775_, _41783_, _41784_);
  or g_51908_(_41767_, _41784_, _41785_);
  not g_51909_(_41785_, _41786_);
  and g_51910_(out[283], _39801_, _41787_);
  xor g_51911_(out[276], out[436], _41788_);
  xor g_51912_(out[274], out[434], _41789_);
  xor g_51913_(out[281], out[441], _41790_);
  xor g_51914_(out[272], out[432], _41791_);
  xor g_51915_(out[275], out[435], _41793_);
  and g_51916_(_39691_, out[443], _41794_);
  xor g_51917_(out[282], out[442], _41795_);
  xor g_51918_(out[287], out[447], _41796_);
  xor g_51919_(out[278], out[438], _41797_);
  xor g_51920_(out[277], out[437], _41798_);
  xor g_51921_(out[285], out[445], _41799_);
  xor g_51922_(out[286], out[446], _41800_);
  xor g_51923_(out[280], out[440], _41801_);
  xor g_51924_(out[273], out[433], _41802_);
  or g_51925_(_41788_, _41800_, _41804_);
  or g_51926_(_41799_, _41801_, _41805_);
  or g_51927_(_41789_, _41795_, _41806_);
  or g_51928_(_41805_, _41806_, _41807_);
  or g_51929_(_41790_, _41793_, _41808_);
  or g_51930_(_41791_, _41798_, _41809_);
  or g_51931_(_41808_, _41809_, _41810_);
  or g_51932_(_41807_, _41810_, _41811_);
  xor g_51933_(out[284], out[444], _41812_);
  or g_51934_(_41794_, _41812_, _41813_);
  xor g_51935_(out[279], out[439], _41815_);
  or g_51936_(_41797_, _41815_, _41816_);
  or g_51937_(_41813_, _41816_, _41817_);
  or g_51938_(_41787_, _41802_, _41818_);
  or g_51939_(_41796_, _41818_, _41819_);
  or g_51940_(_41817_, _41819_, _41820_);
  or g_51941_(_41811_, _41820_, _41821_);
  or g_51942_(_41804_, _41821_, _41822_);
  xor g_51943_(out[263], out[439], _41823_);
  and g_51944_(_39680_, out[443], _41824_);
  xor g_51945_(out[270], out[446], _41826_);
  xor g_51946_(out[264], out[440], _41827_);
  xor g_51947_(out[257], out[433], _41828_);
  xor g_51948_(out[269], out[445], _41829_);
  xor g_51949_(out[265], out[441], _41830_);
  xor g_51950_(out[260], out[436], _41831_);
  xor g_51951_(out[258], out[434], _41832_);
  and g_51952_(out[267], _39801_, _41833_);
  xor g_51953_(out[259], out[435], _41834_);
  xor g_51954_(out[262], out[438], _41835_);
  xor g_51955_(out[271], out[447], _41837_);
  xor g_51956_(out[266], out[442], _41838_);
  xor g_51957_(out[261], out[437], _41839_);
  xor g_51958_(out[256], out[432], _41840_);
  or g_51959_(_41826_, _41831_, _41841_);
  or g_51960_(_41827_, _41829_, _41842_);
  or g_51961_(_41832_, _41838_, _41843_);
  or g_51962_(_41842_, _41843_, _41844_);
  or g_51963_(_41830_, _41834_, _41845_);
  or g_51964_(_41839_, _41840_, _41846_);
  or g_51965_(_41845_, _41846_, _41848_);
  or g_51966_(_41844_, _41848_, _41849_);
  xor g_51967_(out[268], out[444], _41850_);
  or g_51968_(_41824_, _41850_, _41851_);
  or g_51969_(_41823_, _41835_, _41852_);
  or g_51970_(_41851_, _41852_, _41853_);
  or g_51971_(_41828_, _41833_, _41854_);
  or g_51972_(_41837_, _41854_, _41855_);
  or g_51973_(_41853_, _41855_, _41856_);
  or g_51974_(_41849_, _41856_, _41857_);
  or g_51975_(_41841_, _41857_, _41859_);
  xor g_51976_(out[241], out[433], _41860_);
  and g_51977_(out[251], _39801_, _41861_);
  xor g_51978_(out[249], out[441], _41862_);
  xor g_51979_(out[240], out[432], _41863_);
  xor g_51980_(out[254], out[446], _41864_);
  xor g_51981_(out[244], out[436], _41865_);
  or g_51982_(_41864_, _41865_, _41866_);
  xor g_51983_(out[253], out[445], _41867_);
  xor g_51984_(out[243], out[435], _41868_);
  and g_51985_(_39669_, out[443], _41870_);
  xor g_51986_(out[246], out[438], _41871_);
  xor g_51987_(out[250], out[442], _41872_);
  xor g_51988_(out[245], out[437], _41873_);
  xor g_51989_(out[255], out[447], _41874_);
  xor g_51990_(out[248], out[440], _41875_);
  or g_51991_(_41867_, _41875_, _41876_);
  xor g_51992_(out[242], out[434], _41877_);
  or g_51993_(_41872_, _41877_, _41878_);
  or g_51994_(_41876_, _41878_, _41879_);
  or g_51995_(_41862_, _41868_, _41881_);
  or g_51996_(_41873_, _41881_, _41882_);
  or g_51997_(_41879_, _41882_, _41883_);
  or g_51998_(_41866_, _41883_, _41884_);
  xor g_51999_(out[252], out[444], _41885_);
  or g_52000_(_41870_, _41885_, _41886_);
  xor g_52001_(out[247], out[439], _41887_);
  or g_52002_(_41871_, _41887_, _41888_);
  or g_52003_(_41886_, _41888_, _41889_);
  or g_52004_(_41860_, _41861_, _41890_);
  or g_52005_(_41874_, _41890_, _41892_);
  or g_52006_(_41889_, _41892_, _41893_);
  or g_52007_(_41863_, _41893_, _41894_);
  or g_52008_(_41884_, _41894_, _41895_);
  xor g_52009_(out[231], out[439], _41896_);
  and g_52010_(_39658_, out[443], _41897_);
  xor g_52011_(out[238], out[446], _41898_);
  xor g_52012_(out[232], out[440], _41899_);
  xor g_52013_(out[225], out[433], _41900_);
  xor g_52014_(out[237], out[445], _41901_);
  xor g_52015_(out[233], out[441], _41903_);
  xor g_52016_(out[228], out[436], _41904_);
  xor g_52017_(out[226], out[434], _41905_);
  and g_52018_(out[235], _39801_, _41906_);
  xor g_52019_(out[227], out[435], _41907_);
  xor g_52020_(out[230], out[438], _41908_);
  xor g_52021_(out[239], out[447], _41909_);
  xor g_52022_(out[234], out[442], _41910_);
  xor g_52023_(out[229], out[437], _41911_);
  xor g_52024_(out[224], out[432], _41912_);
  or g_52025_(_41898_, _41904_, _41914_);
  or g_52026_(_41899_, _41901_, _41915_);
  or g_52027_(_41905_, _41910_, _41916_);
  or g_52028_(_41915_, _41916_, _41917_);
  or g_52029_(_41903_, _41907_, _41918_);
  or g_52030_(_41911_, _41912_, _41919_);
  or g_52031_(_41918_, _41919_, _41920_);
  or g_52032_(_41917_, _41920_, _41921_);
  xor g_52033_(out[236], out[444], _41922_);
  or g_52034_(_41897_, _41922_, _41923_);
  or g_52035_(_41896_, _41908_, _41925_);
  or g_52036_(_41923_, _41925_, _41926_);
  or g_52037_(_41900_, _41906_, _41927_);
  or g_52038_(_41909_, _41927_, _41928_);
  or g_52039_(_41926_, _41928_, _41929_);
  or g_52040_(_41921_, _41929_, _41930_);
  or g_52041_(_41914_, _41930_, _41931_);
  xor g_52042_(out[209], out[433], _41932_);
  and g_52043_(out[219], _39801_, _41933_);
  xor g_52044_(out[217], out[441], _41934_);
  xor g_52045_(out[208], out[432], _41936_);
  xor g_52046_(out[222], out[446], _41937_);
  xor g_52047_(out[212], out[436], _41938_);
  or g_52048_(_41937_, _41938_, _41939_);
  xor g_52049_(out[221], out[445], _41940_);
  xor g_52050_(out[211], out[435], _41941_);
  and g_52051_(_39647_, out[443], _41942_);
  xor g_52052_(out[214], out[438], _41943_);
  xor g_52053_(out[218], out[442], _41944_);
  xor g_52054_(out[213], out[437], _41945_);
  xor g_52055_(out[223], out[447], _41947_);
  xor g_52056_(out[216], out[440], _41948_);
  or g_52057_(_41940_, _41948_, _41949_);
  xor g_52058_(out[210], out[434], _41950_);
  or g_52059_(_41944_, _41950_, _41951_);
  or g_52060_(_41949_, _41951_, _41952_);
  or g_52061_(_41934_, _41941_, _41953_);
  or g_52062_(_41945_, _41953_, _41954_);
  or g_52063_(_41952_, _41954_, _41955_);
  or g_52064_(_41939_, _41955_, _41956_);
  xor g_52065_(out[220], out[444], _41958_);
  or g_52066_(_41942_, _41958_, _41959_);
  xor g_52067_(out[215], out[439], _41960_);
  or g_52068_(_41943_, _41960_, _41961_);
  or g_52069_(_41959_, _41961_, _41962_);
  or g_52070_(_41932_, _41933_, _41963_);
  or g_52071_(_41947_, _41963_, _41964_);
  or g_52072_(_41962_, _41964_, _41965_);
  or g_52073_(_41936_, _41965_, _41966_);
  or g_52074_(_41956_, _41966_, _41967_);
  xor g_52075_(out[199], out[439], _41969_);
  and g_52076_(_39636_, out[443], _41970_);
  xor g_52077_(out[206], out[446], _41971_);
  xor g_52078_(out[200], out[440], _41972_);
  xor g_52079_(out[193], out[433], _41973_);
  xor g_52080_(out[205], out[445], _41974_);
  xor g_52081_(out[201], out[441], _41975_);
  xor g_52082_(out[196], out[436], _41976_);
  xor g_52083_(out[194], out[434], _41977_);
  and g_52084_(out[203], _39801_, _41978_);
  xor g_52085_(out[195], out[435], _41980_);
  xor g_52086_(out[198], out[438], _41981_);
  xor g_52087_(out[207], out[447], _41982_);
  xor g_52088_(out[202], out[442], _41983_);
  xor g_52089_(out[197], out[437], _41984_);
  xor g_52090_(out[192], out[432], _41985_);
  or g_52091_(_41971_, _41976_, _41986_);
  or g_52092_(_41972_, _41974_, _41987_);
  or g_52093_(_41977_, _41983_, _41988_);
  or g_52094_(_41987_, _41988_, _41989_);
  or g_52095_(_41975_, _41980_, _41991_);
  or g_52096_(_41984_, _41985_, _41992_);
  or g_52097_(_41991_, _41992_, _41993_);
  or g_52098_(_41989_, _41993_, _41994_);
  xor g_52099_(out[204], out[444], _41995_);
  or g_52100_(_41970_, _41995_, _41996_);
  or g_52101_(_41969_, _41981_, _41997_);
  or g_52102_(_41996_, _41997_, _41998_);
  or g_52103_(_41973_, _41978_, _41999_);
  or g_52104_(_41982_, _41999_, _42000_);
  or g_52105_(_41998_, _42000_, _42002_);
  or g_52106_(_41994_, _42002_, _42003_);
  or g_52107_(_41986_, _42003_, _42004_);
  xor g_52108_(out[177], out[433], _42005_);
  and g_52109_(out[187], _39801_, _42006_);
  xor g_52110_(out[185], out[441], _42007_);
  xor g_52111_(out[176], out[432], _42008_);
  xor g_52112_(out[190], out[446], _42009_);
  xor g_52113_(out[180], out[436], _42010_);
  or g_52114_(_42009_, _42010_, _42011_);
  xor g_52115_(out[189], out[445], _42013_);
  xor g_52116_(out[179], out[435], _42014_);
  and g_52117_(_39625_, out[443], _42015_);
  xor g_52118_(out[182], out[438], _42016_);
  xor g_52119_(out[186], out[442], _42017_);
  xor g_52120_(out[181], out[437], _42018_);
  xor g_52121_(out[191], out[447], _42019_);
  xor g_52122_(out[184], out[440], _42020_);
  or g_52123_(_42013_, _42020_, _42021_);
  xor g_52124_(out[178], out[434], _42022_);
  or g_52125_(_42017_, _42022_, _42024_);
  or g_52126_(_42021_, _42024_, _42025_);
  or g_52127_(_42007_, _42014_, _42026_);
  or g_52128_(_42018_, _42026_, _42027_);
  or g_52129_(_42025_, _42027_, _42028_);
  or g_52130_(_42011_, _42028_, _42029_);
  xor g_52131_(out[188], out[444], _42030_);
  or g_52132_(_42015_, _42030_, _42031_);
  xor g_52133_(out[183], out[439], _42032_);
  or g_52134_(_42016_, _42032_, _42033_);
  or g_52135_(_42031_, _42033_, _42035_);
  or g_52136_(_42005_, _42006_, _42036_);
  or g_52137_(_42019_, _42036_, _42037_);
  or g_52138_(_42035_, _42037_, _42038_);
  or g_52139_(_42008_, _42038_, _42039_);
  or g_52140_(_42029_, _42039_, _42040_);
  xor g_52141_(out[167], out[439], _42041_);
  and g_52142_(_39614_, out[443], _42042_);
  xor g_52143_(out[174], out[446], _42043_);
  xor g_52144_(out[168], out[440], _42044_);
  xor g_52145_(out[161], out[433], _42046_);
  xor g_52146_(out[173], out[445], _42047_);
  xor g_52147_(out[169], out[441], _42048_);
  xor g_52148_(out[164], out[436], _42049_);
  xor g_52149_(out[162], out[434], _42050_);
  and g_52150_(out[171], _39801_, _42051_);
  xor g_52151_(out[163], out[435], _42052_);
  xor g_52152_(out[166], out[438], _42053_);
  xor g_52153_(out[175], out[447], _42054_);
  xor g_52154_(out[170], out[442], _42055_);
  xor g_52155_(out[165], out[437], _42057_);
  xor g_52156_(out[160], out[432], _42058_);
  or g_52157_(_42043_, _42049_, _42059_);
  or g_52158_(_42044_, _42047_, _42060_);
  or g_52159_(_42050_, _42055_, _42061_);
  or g_52160_(_42060_, _42061_, _42062_);
  or g_52161_(_42048_, _42052_, _42063_);
  or g_52162_(_42057_, _42058_, _42064_);
  or g_52163_(_42063_, _42064_, _42065_);
  or g_52164_(_42062_, _42065_, _42066_);
  xor g_52165_(out[172], out[444], _42068_);
  or g_52166_(_42042_, _42068_, _42069_);
  or g_52167_(_42041_, _42053_, _42070_);
  or g_52168_(_42069_, _42070_, _42071_);
  or g_52169_(_42046_, _42051_, _42072_);
  or g_52170_(_42054_, _42072_, _42073_);
  or g_52171_(_42071_, _42073_, _42074_);
  or g_52172_(_42066_, _42074_, _42075_);
  or g_52173_(_42059_, _42075_, _42076_);
  xor g_52174_(out[148], out[436], _42077_);
  xor g_52175_(out[156], out[444], _42079_);
  and g_52176_(_39603_, out[443], _42080_);
  xor g_52177_(out[154], out[442], _42081_);
  xor g_52178_(out[150], out[438], _42082_);
  xor g_52179_(out[149], out[437], _42083_);
  xor g_52180_(out[147], out[435], _42084_);
  xor g_52181_(out[157], out[445], _42085_);
  xor g_52182_(out[158], out[446], _42086_);
  xor g_52183_(out[145], out[433], _42087_);
  xor g_52184_(out[146], out[434], _42088_);
  and g_52185_(out[155], _39801_, _42090_);
  xor g_52186_(out[144], out[432], _42091_);
  xor g_52187_(out[159], out[447], _42092_);
  xor g_52188_(out[152], out[440], _42093_);
  or g_52189_(_42085_, _42093_, _42094_);
  xor g_52190_(out[153], out[441], _42095_);
  or g_52191_(_42081_, _42088_, _42096_);
  or g_52192_(_42094_, _42096_, _42097_);
  or g_52193_(_42084_, _42095_, _42098_);
  or g_52194_(_42083_, _42098_, _42099_);
  or g_52195_(_42097_, _42099_, _42101_);
  or g_52196_(_42077_, _42086_, _42102_);
  or g_52197_(_42101_, _42102_, _42103_);
  or g_52198_(_42079_, _42080_, _42104_);
  xor g_52199_(out[151], out[439], _42105_);
  or g_52200_(_42082_, _42105_, _42106_);
  or g_52201_(_42104_, _42106_, _42107_);
  or g_52202_(_42087_, _42090_, _42108_);
  or g_52203_(_42092_, _42108_, _42109_);
  or g_52204_(_42107_, _42109_, _42110_);
  or g_52205_(_42091_, _42110_, _42112_);
  or g_52206_(_42103_, _42112_, _42113_);
  not g_52207_(_42113_, _42114_);
  xor g_52208_(out[135], out[439], _42115_);
  and g_52209_(_39592_, out[443], _42116_);
  xor g_52210_(out[142], out[446], _42117_);
  xor g_52211_(out[136], out[440], _42118_);
  xor g_52212_(out[129], out[433], _42119_);
  xor g_52213_(out[141], out[445], _42120_);
  xor g_52214_(out[137], out[441], _42121_);
  xor g_52215_(out[132], out[436], _42123_);
  xor g_52216_(out[130], out[434], _42124_);
  and g_52217_(out[139], _39801_, _42125_);
  xor g_52218_(out[131], out[435], _42126_);
  xor g_52219_(out[134], out[438], _42127_);
  xor g_52220_(out[143], out[447], _42128_);
  xor g_52221_(out[138], out[442], _42129_);
  xor g_52222_(out[133], out[437], _42130_);
  xor g_52223_(out[128], out[432], _42131_);
  or g_52224_(_42117_, _42123_, _42132_);
  or g_52225_(_42118_, _42120_, _42134_);
  or g_52226_(_42124_, _42129_, _42135_);
  or g_52227_(_42134_, _42135_, _42136_);
  or g_52228_(_42121_, _42126_, _42137_);
  or g_52229_(_42130_, _42131_, _42138_);
  or g_52230_(_42137_, _42138_, _42139_);
  or g_52231_(_42136_, _42139_, _42140_);
  xor g_52232_(out[140], out[444], _42141_);
  or g_52233_(_42116_, _42141_, _42142_);
  or g_52234_(_42115_, _42127_, _42143_);
  or g_52235_(_42142_, _42143_, _42145_);
  or g_52236_(_42119_, _42125_, _42146_);
  or g_52237_(_42128_, _42146_, _42147_);
  or g_52238_(_42145_, _42147_, _42148_);
  or g_52239_(_42140_, _42148_, _42149_);
  or g_52240_(_42132_, _42149_, _42150_);
  xor g_52241_(out[113], out[433], _42151_);
  and g_52242_(out[123], _39801_, _42152_);
  xor g_52243_(out[116], out[436], _42153_);
  xor g_52244_(out[118], out[438], _42154_);
  xor g_52245_(out[115], out[435], _42156_);
  xor g_52246_(out[119], out[439], _42157_);
  and g_52247_(_39581_, out[443], _42158_);
  xor g_52248_(out[122], out[442], _42159_);
  xor g_52249_(out[114], out[434], _42160_);
  or g_52250_(_42159_, _42160_, _42161_);
  xor g_52251_(out[126], out[446], _42162_);
  xor g_52252_(out[112], out[432], _42163_);
  xor g_52253_(out[125], out[445], _42164_);
  xor g_52254_(out[120], out[440], _42165_);
  or g_52255_(_42164_, _42165_, _42167_);
  xor g_52256_(out[121], out[441], _42168_);
  xor g_52257_(out[127], out[447], _42169_);
  xor g_52258_(out[117], out[437], _42170_);
  or g_52259_(_42161_, _42167_, _42171_);
  or g_52260_(_42156_, _42168_, _42172_);
  or g_52261_(_42170_, _42172_, _42173_);
  or g_52262_(_42171_, _42173_, _42174_);
  or g_52263_(_42153_, _42162_, _42175_);
  or g_52264_(_42174_, _42175_, _42176_);
  xor g_52265_(out[124], out[444], _42178_);
  or g_52266_(_42158_, _42178_, _42179_);
  or g_52267_(_42154_, _42157_, _42180_);
  or g_52268_(_42179_, _42180_, _42181_);
  or g_52269_(_42151_, _42152_, _42182_);
  or g_52270_(_42169_, _42182_, _42183_);
  or g_52271_(_42181_, _42183_, _42184_);
  or g_52272_(_42163_, _42184_, _42185_);
  or g_52273_(_42176_, _42185_, _42186_);
  xor g_52274_(out[103], out[439], _42187_);
  and g_52275_(_39570_, out[443], _42189_);
  xor g_52276_(out[110], out[446], _42190_);
  xor g_52277_(out[104], out[440], _42191_);
  xor g_52278_(out[97], out[433], _42192_);
  xor g_52279_(out[109], out[445], _42193_);
  xor g_52280_(out[105], out[441], _42194_);
  xor g_52281_(out[100], out[436], _42195_);
  xor g_52282_(out[98], out[434], _42196_);
  and g_52283_(out[107], _39801_, _42197_);
  xor g_52284_(out[99], out[435], _42198_);
  xor g_52285_(out[102], out[438], _42200_);
  xor g_52286_(out[111], out[447], _42201_);
  xor g_52287_(out[106], out[442], _42202_);
  xor g_52288_(out[101], out[437], _42203_);
  xor g_52289_(out[96], out[432], _42204_);
  or g_52290_(_42190_, _42195_, _42205_);
  or g_52291_(_42191_, _42193_, _42206_);
  or g_52292_(_42196_, _42202_, _42207_);
  or g_52293_(_42206_, _42207_, _42208_);
  or g_52294_(_42194_, _42198_, _42209_);
  or g_52295_(_42203_, _42204_, _42211_);
  or g_52296_(_42209_, _42211_, _42212_);
  or g_52297_(_42208_, _42212_, _42213_);
  xor g_52298_(out[108], out[444], _42214_);
  or g_52299_(_42189_, _42214_, _42215_);
  or g_52300_(_42187_, _42200_, _42216_);
  or g_52301_(_42215_, _42216_, _42217_);
  or g_52302_(_42192_, _42197_, _42218_);
  or g_52303_(_42201_, _42218_, _42219_);
  or g_52304_(_42217_, _42219_, _42220_);
  or g_52305_(_42213_, _42220_, _42222_);
  or g_52306_(_42205_, _42222_, _42223_);
  xor g_52307_(out[92], out[444], _42224_);
  and g_52308_(_39559_, out[443], _42225_);
  xor g_52309_(out[88], out[440], _42226_);
  xor g_52310_(out[86], out[438], _42227_);
  xor g_52311_(out[93], out[445], _42228_);
  xor g_52312_(out[94], out[446], _42229_);
  xor g_52313_(out[82], out[434], _42230_);
  xor g_52314_(out[89], out[441], _42231_);
  xor g_52315_(out[85], out[437], _42233_);
  xor g_52316_(out[81], out[433], _42234_);
  and g_52317_(out[91], _39801_, _42235_);
  or g_52318_(_42226_, _42228_, _42236_);
  xor g_52319_(out[95], out[447], _42237_);
  xor g_52320_(out[90], out[442], _42238_);
  xor g_52321_(out[84], out[436], _42239_);
  xor g_52322_(out[83], out[435], _42240_);
  xor g_52323_(out[80], out[432], _42241_);
  or g_52324_(_42230_, _42238_, _42242_);
  or g_52325_(_42236_, _42242_, _42244_);
  or g_52326_(_42231_, _42240_, _42245_);
  or g_52327_(_42233_, _42245_, _42246_);
  or g_52328_(_42244_, _42246_, _42247_);
  or g_52329_(_42229_, _42239_, _42248_);
  or g_52330_(_42247_, _42248_, _42249_);
  or g_52331_(_42224_, _42225_, _42250_);
  xor g_52332_(out[87], out[439], _42251_);
  or g_52333_(_42227_, _42251_, _42252_);
  or g_52334_(_42250_, _42252_, _42253_);
  or g_52335_(_42234_, _42235_, _42255_);
  or g_52336_(_42237_, _42255_, _42256_);
  or g_52337_(_42253_, _42256_, _42257_);
  or g_52338_(_42241_, _42257_, _42258_);
  or g_52339_(_42249_, _42258_, _42259_);
  xor g_52340_(out[71], out[439], _42260_);
  and g_52341_(_39548_, out[443], _42261_);
  xor g_52342_(out[78], out[446], _42262_);
  xor g_52343_(out[72], out[440], _42263_);
  xor g_52344_(out[65], out[433], _42264_);
  xor g_52345_(out[77], out[445], _42266_);
  xor g_52346_(out[73], out[441], _42267_);
  xor g_52347_(out[68], out[436], _42268_);
  xor g_52348_(out[66], out[434], _42269_);
  and g_52349_(out[75], _39801_, _42270_);
  xor g_52350_(out[67], out[435], _42271_);
  xor g_52351_(out[70], out[438], _42272_);
  xor g_52352_(out[79], out[447], _42273_);
  xor g_52353_(out[74], out[442], _42274_);
  xor g_52354_(out[69], out[437], _42275_);
  xor g_52355_(out[64], out[432], _42277_);
  or g_52356_(_42262_, _42268_, _42278_);
  or g_52357_(_42263_, _42266_, _42279_);
  or g_52358_(_42269_, _42274_, _42280_);
  or g_52359_(_42279_, _42280_, _42281_);
  or g_52360_(_42267_, _42271_, _42282_);
  or g_52361_(_42275_, _42277_, _42283_);
  or g_52362_(_42282_, _42283_, _42284_);
  or g_52363_(_42281_, _42284_, _42285_);
  xor g_52364_(out[76], out[444], _42286_);
  or g_52365_(_42261_, _42286_, _42288_);
  or g_52366_(_42260_, _42272_, _42289_);
  or g_52367_(_42288_, _42289_, _42290_);
  or g_52368_(_42264_, _42270_, _42291_);
  or g_52369_(_42273_, _42291_, _42292_);
  or g_52370_(_42290_, _42292_, _42293_);
  or g_52371_(_42285_, _42293_, _42294_);
  or g_52372_(_42278_, _42294_, _42295_);
  not g_52373_(_42295_, _42296_);
  xor g_52374_(out[51], out[435], _42297_);
  xor g_52375_(out[52], out[436], _42299_);
  xor g_52376_(out[62], out[446], _42300_);
  xor g_52377_(out[50], out[434], _42301_);
  xor g_52378_(out[53], out[437], _42302_);
  xor g_52379_(out[57], out[441], _42303_);
  xor g_52380_(out[56], out[440], _42304_);
  xor g_52381_(out[63], out[447], _42305_);
  xor g_52382_(out[58], out[442], _42306_);
  xor g_52383_(out[54], out[438], _42307_);
  xor g_52384_(out[48], out[432], _42308_);
  and g_52385_(_39537_, out[443], _42310_);
  and g_52386_(out[59], _39801_, _42311_);
  xor g_52387_(out[61], out[445], _42312_);
  or g_52388_(_42304_, _42312_, _42313_);
  xor g_52389_(out[49], out[433], _42314_);
  or g_52390_(_42301_, _42306_, _42315_);
  or g_52391_(_42313_, _42315_, _42316_);
  or g_52392_(_42297_, _42303_, _42317_);
  or g_52393_(_42302_, _42317_, _42318_);
  or g_52394_(_42316_, _42318_, _42319_);
  or g_52395_(_42299_, _42300_, _42321_);
  or g_52396_(_42319_, _42321_, _42322_);
  xor g_52397_(out[60], out[444], _42323_);
  or g_52398_(_42310_, _42323_, _42324_);
  xor g_52399_(out[55], out[439], _42325_);
  or g_52400_(_42307_, _42325_, _42326_);
  or g_52401_(_42324_, _42326_, _42327_);
  or g_52402_(_42311_, _42314_, _42328_);
  or g_52403_(_42305_, _42328_, _42329_);
  or g_52404_(_42327_, _42329_, _42330_);
  or g_52405_(_42308_, _42330_, _42332_);
  or g_52406_(_42322_, _42332_, _42333_);
  not g_52407_(_42333_, _42334_);
  xor g_52408_(out[39], out[439], _42335_);
  and g_52409_(_39526_, out[443], _42336_);
  xor g_52410_(out[46], out[446], _42337_);
  xor g_52411_(out[40], out[440], _42338_);
  xor g_52412_(out[33], out[433], _42339_);
  xor g_52413_(out[45], out[445], _42340_);
  xor g_52414_(out[41], out[441], _42341_);
  xor g_52415_(out[36], out[436], _42343_);
  xor g_52416_(out[34], out[434], _42344_);
  and g_52417_(out[43], _39801_, _42345_);
  xor g_52418_(out[35], out[435], _42346_);
  xor g_52419_(out[38], out[438], _42347_);
  xor g_52420_(out[47], out[447], _42348_);
  xor g_52421_(out[42], out[442], _42349_);
  xor g_52422_(out[37], out[437], _42350_);
  xor g_52423_(out[32], out[432], _42351_);
  or g_52424_(_42337_, _42343_, _42352_);
  or g_52425_(_42338_, _42340_, _42354_);
  or g_52426_(_42344_, _42349_, _42355_);
  or g_52427_(_42354_, _42355_, _42356_);
  or g_52428_(_42341_, _42346_, _42357_);
  or g_52429_(_42350_, _42351_, _42358_);
  or g_52430_(_42357_, _42358_, _42359_);
  or g_52431_(_42356_, _42359_, _42360_);
  xor g_52432_(out[44], out[444], _42361_);
  or g_52433_(_42336_, _42361_, _42362_);
  or g_52434_(_42335_, _42347_, _42363_);
  or g_52435_(_42362_, _42363_, _42365_);
  or g_52436_(_42339_, _42345_, _42366_);
  or g_52437_(_42348_, _42366_, _42367_);
  or g_52438_(_42365_, _42367_, _42368_);
  or g_52439_(_42360_, _42368_, _42369_);
  or g_52440_(_42352_, _42369_, _42370_);
  xor g_52441_(out[28], out[444], _42371_);
  and g_52442_(_39493_, out[443], _42372_);
  xor g_52443_(out[29], out[445], _42373_);
  xor g_52444_(out[22], out[438], _42374_);
  xor g_52445_(out[24], out[440], _42376_);
  xor g_52446_(out[25], out[441], _42377_);
  xor g_52447_(out[30], out[446], _42378_);
  xor g_52448_(out[20], out[436], _42379_);
  or g_52449_(_42378_, _42379_, _42380_);
  xor g_52450_(out[21], out[437], _42381_);
  xor g_52451_(out[17], out[433], _42382_);
  and g_52452_(out[27], _39801_, _42383_);
  xor g_52453_(out[31], out[447], _42384_);
  xor g_52454_(out[26], out[442], _42385_);
  xor g_52455_(out[16], out[432], _42387_);
  xor g_52456_(out[18], out[434], _42388_);
  xor g_52457_(out[19], out[435], _42389_);
  or g_52458_(_42373_, _42376_, _42390_);
  or g_52459_(_42385_, _42388_, _42391_);
  or g_52460_(_42390_, _42391_, _42392_);
  or g_52461_(_42377_, _42389_, _42393_);
  or g_52462_(_42381_, _42387_, _42394_);
  or g_52463_(_42393_, _42394_, _42395_);
  or g_52464_(_42392_, _42395_, _42396_);
  or g_52465_(_42371_, _42372_, _42398_);
  xor g_52466_(out[23], out[439], _42399_);
  or g_52467_(_42374_, _42399_, _42400_);
  or g_52468_(_42398_, _42400_, _42401_);
  or g_52469_(_42382_, _42383_, _42402_);
  or g_52470_(_42384_, _42402_, _42403_);
  or g_52471_(_42401_, _42403_, _42404_);
  or g_52472_(_42396_, _42404_, _42405_);
  or g_52473_(_42380_, _42405_, _42406_);
  xor g_52474_(out[1], out[433], _42407_);
  and g_52475_(out[11], _39801_, _42409_);
  xor g_52476_(out[14], out[446], _42410_);
  xor g_52477_(out[3], out[435], _42411_);
  xor g_52478_(out[4], out[436], _42412_);
  xor g_52479_(out[2], out[434], _42413_);
  xor g_52480_(out[9], out[441], _42414_);
  xor g_52481_(out[0], out[432], _42415_);
  and g_52482_(_39438_, out[443], _42416_);
  xor g_52483_(out[6], out[438], _42417_);
  xor g_52484_(out[10], out[442], _42418_);
  xor g_52485_(out[5], out[437], _42420_);
  xor g_52486_(out[15], out[447], _42421_);
  xor g_52487_(out[13], out[445], _42422_);
  xor g_52488_(out[8], out[440], _42423_);
  or g_52489_(_42410_, _42412_, _42424_);
  or g_52490_(_42422_, _42423_, _42425_);
  or g_52491_(_42413_, _42418_, _42426_);
  or g_52492_(_42425_, _42426_, _42427_);
  or g_52493_(_42411_, _42414_, _42428_);
  or g_52494_(_42415_, _42420_, _42429_);
  or g_52495_(_42428_, _42429_, _42431_);
  or g_52496_(_42427_, _42431_, _42432_);
  xor g_52497_(out[12], out[444], _42433_);
  or g_52498_(_42416_, _42433_, _42434_);
  xor g_52499_(out[7], out[439], _42435_);
  or g_52500_(_42417_, _42435_, _42436_);
  or g_52501_(_42434_, _42436_, _42437_);
  or g_52502_(_42407_, _42409_, _42438_);
  or g_52503_(_42421_, _42438_, _42439_);
  or g_52504_(_42437_, _42439_, _42440_);
  or g_52505_(_42432_, _42440_, _42442_);
  or g_52506_(_42424_, _42442_, _42443_);
  xor g_52507_(out[311], out[423], _42444_);
  and g_52508_(_39724_, out[427], _42445_);
  xor g_52509_(out[318], out[430], _42446_);
  xor g_52510_(out[312], out[424], _42447_);
  xor g_52511_(out[305], out[417], _42448_);
  xor g_52512_(out[317], out[429], _42449_);
  xor g_52513_(out[313], out[425], _42450_);
  xor g_52514_(out[308], out[420], _42451_);
  xor g_52515_(out[306], out[418], _42453_);
  and g_52516_(out[315], _39790_, _42454_);
  xor g_52517_(out[307], out[419], _42455_);
  xor g_52518_(out[310], out[422], _42456_);
  xor g_52519_(out[319], out[431], _42457_);
  xor g_52520_(out[314], out[426], _42458_);
  xor g_52521_(out[309], out[421], _42459_);
  xor g_52522_(out[304], out[416], _42460_);
  or g_52523_(_42446_, _42451_, _42461_);
  or g_52524_(_42447_, _42449_, _42462_);
  or g_52525_(_42453_, _42458_, _42464_);
  or g_52526_(_42462_, _42464_, _42465_);
  or g_52527_(_42450_, _42455_, _42466_);
  or g_52528_(_42459_, _42460_, _42467_);
  or g_52529_(_42466_, _42467_, _42468_);
  or g_52530_(_42465_, _42468_, _42469_);
  xor g_52531_(out[316], out[428], _42470_);
  or g_52532_(_42445_, _42470_, _42471_);
  or g_52533_(_42444_, _42456_, _42472_);
  or g_52534_(_42471_, _42472_, _42473_);
  or g_52535_(_42448_, _42454_, _42475_);
  or g_52536_(_42457_, _42475_, _42476_);
  or g_52537_(_42473_, _42476_, _42477_);
  or g_52538_(_42469_, _42477_, _42478_);
  or g_52539_(_42461_, _42478_, _42479_);
  xor g_52540_(out[298], out[426], _42480_);
  xor g_52541_(out[290], out[418], _42481_);
  xor g_52542_(out[289], out[417], _42482_);
  and g_52543_(_39702_, out[427], _42483_);
  and g_52544_(out[299], _39790_, _42484_);
  xor g_52545_(out[301], out[429], _42486_);
  xor g_52546_(out[291], out[419], _42487_);
  xor g_52547_(out[302], out[430], _42488_);
  xor g_52548_(out[300], out[428], _42489_);
  xor g_52549_(out[296], out[424], _42490_);
  xor g_52550_(out[303], out[431], _42491_);
  xor g_52551_(out[293], out[421], _42492_);
  xor g_52552_(out[294], out[422], _42493_);
  xor g_52553_(out[288], out[416], _42494_);
  xor g_52554_(out[292], out[420], _42495_);
  or g_52555_(_42486_, _42490_, _42497_);
  xor g_52556_(out[297], out[425], _42498_);
  or g_52557_(_42480_, _42481_, _42499_);
  or g_52558_(_42497_, _42499_, _42500_);
  or g_52559_(_42487_, _42498_, _42501_);
  or g_52560_(_42492_, _42501_, _42502_);
  or g_52561_(_42500_, _42502_, _42503_);
  or g_52562_(_42488_, _42495_, _42504_);
  or g_52563_(_42503_, _42504_, _42505_);
  or g_52564_(_42483_, _42489_, _42506_);
  xor g_52565_(out[295], out[423], _42508_);
  or g_52566_(_42493_, _42508_, _42509_);
  or g_52567_(_42506_, _42509_, _42510_);
  or g_52568_(_42482_, _42484_, _42511_);
  or g_52569_(_42491_, _42511_, _42512_);
  or g_52570_(_42510_, _42512_, _42513_);
  or g_52571_(_42494_, _42513_, _42514_);
  or g_52572_(_42505_, _42514_, _42515_);
  not g_52573_(_42515_, _42516_);
  xor g_52574_(out[279], out[423], _42517_);
  and g_52575_(_39691_, out[427], _42519_);
  xor g_52576_(out[286], out[430], _42520_);
  xor g_52577_(out[280], out[424], _42521_);
  xor g_52578_(out[273], out[417], _42522_);
  xor g_52579_(out[285], out[429], _42523_);
  xor g_52580_(out[281], out[425], _42524_);
  xor g_52581_(out[276], out[420], _42525_);
  xor g_52582_(out[274], out[418], _42526_);
  and g_52583_(out[283], _39790_, _42527_);
  xor g_52584_(out[275], out[419], _42528_);
  xor g_52585_(out[278], out[422], _42530_);
  xor g_52586_(out[287], out[431], _42531_);
  xor g_52587_(out[282], out[426], _42532_);
  xor g_52588_(out[277], out[421], _42533_);
  xor g_52589_(out[272], out[416], _42534_);
  or g_52590_(_42520_, _42525_, _42535_);
  or g_52591_(_42521_, _42523_, _42536_);
  or g_52592_(_42526_, _42532_, _42537_);
  or g_52593_(_42536_, _42537_, _42538_);
  or g_52594_(_42524_, _42528_, _42539_);
  or g_52595_(_42533_, _42534_, _42541_);
  or g_52596_(_42539_, _42541_, _42542_);
  or g_52597_(_42538_, _42542_, _42543_);
  xor g_52598_(out[284], out[428], _42544_);
  or g_52599_(_42519_, _42544_, _42545_);
  or g_52600_(_42517_, _42530_, _42546_);
  or g_52601_(_42545_, _42546_, _42547_);
  or g_52602_(_42522_, _42527_, _42548_);
  or g_52603_(_42531_, _42548_, _42549_);
  or g_52604_(_42547_, _42549_, _42550_);
  or g_52605_(_42543_, _42550_, _42552_);
  or g_52606_(_42535_, _42552_, _42553_);
  xor g_52607_(out[259], out[419], _42554_);
  xor g_52608_(out[260], out[420], _42555_);
  xor g_52609_(out[270], out[430], _42556_);
  xor g_52610_(out[258], out[418], _42557_);
  xor g_52611_(out[261], out[421], _42558_);
  xor g_52612_(out[265], out[425], _42559_);
  xor g_52613_(out[264], out[424], _42560_);
  xor g_52614_(out[271], out[431], _42561_);
  xor g_52615_(out[266], out[426], _42563_);
  xor g_52616_(out[262], out[422], _42564_);
  xor g_52617_(out[256], out[416], _42565_);
  and g_52618_(_39680_, out[427], _42566_);
  and g_52619_(out[267], _39790_, _42567_);
  xor g_52620_(out[269], out[429], _42568_);
  or g_52621_(_42560_, _42568_, _42569_);
  xor g_52622_(out[257], out[417], _42570_);
  or g_52623_(_42557_, _42563_, _42571_);
  or g_52624_(_42569_, _42571_, _42572_);
  or g_52625_(_42554_, _42559_, _42574_);
  or g_52626_(_42558_, _42574_, _42575_);
  or g_52627_(_42572_, _42575_, _42576_);
  or g_52628_(_42555_, _42556_, _42577_);
  or g_52629_(_42576_, _42577_, _42578_);
  xor g_52630_(out[268], out[428], _42579_);
  or g_52631_(_42566_, _42579_, _42580_);
  xor g_52632_(out[263], out[423], _42581_);
  or g_52633_(_42564_, _42581_, _42582_);
  or g_52634_(_42580_, _42582_, _42583_);
  or g_52635_(_42567_, _42570_, _42585_);
  or g_52636_(_42561_, _42585_, _42586_);
  or g_52637_(_42583_, _42586_, _42587_);
  or g_52638_(_42565_, _42587_, _42588_);
  or g_52639_(_42578_, _42588_, _42589_);
  xor g_52640_(out[247], out[423], _42590_);
  and g_52641_(_39669_, out[427], _42591_);
  xor g_52642_(out[254], out[430], _42592_);
  xor g_52643_(out[248], out[424], _42593_);
  xor g_52644_(out[241], out[417], _42594_);
  xor g_52645_(out[253], out[429], _42596_);
  xor g_52646_(out[249], out[425], _42597_);
  xor g_52647_(out[244], out[420], _42598_);
  xor g_52648_(out[242], out[418], _42599_);
  and g_52649_(out[251], _39790_, _42600_);
  xor g_52650_(out[243], out[419], _42601_);
  xor g_52651_(out[246], out[422], _42602_);
  xor g_52652_(out[255], out[431], _42603_);
  xor g_52653_(out[250], out[426], _42604_);
  xor g_52654_(out[245], out[421], _42605_);
  xor g_52655_(out[240], out[416], _42607_);
  or g_52656_(_42592_, _42598_, _42608_);
  or g_52657_(_42593_, _42596_, _42609_);
  or g_52658_(_42599_, _42604_, _42610_);
  or g_52659_(_42609_, _42610_, _42611_);
  or g_52660_(_42597_, _42601_, _42612_);
  or g_52661_(_42605_, _42607_, _42613_);
  or g_52662_(_42612_, _42613_, _42614_);
  or g_52663_(_42611_, _42614_, _42615_);
  xor g_52664_(out[252], out[428], _42616_);
  or g_52665_(_42591_, _42616_, _42618_);
  or g_52666_(_42590_, _42602_, _42619_);
  or g_52667_(_42618_, _42619_, _42620_);
  or g_52668_(_42594_, _42600_, _42621_);
  or g_52669_(_42603_, _42621_, _42622_);
  or g_52670_(_42620_, _42622_, _42623_);
  or g_52671_(_42615_, _42623_, _42624_);
  or g_52672_(_42608_, _42624_, _42625_);
  not g_52673_(_42625_, _42626_);
  xor g_52674_(out[225], out[417], _42627_);
  and g_52675_(out[235], _39790_, _42629_);
  xor g_52676_(out[238], out[430], _42630_);
  xor g_52677_(out[227], out[419], _42631_);
  xor g_52678_(out[228], out[420], _42632_);
  xor g_52679_(out[226], out[418], _42633_);
  xor g_52680_(out[233], out[425], _42634_);
  xor g_52681_(out[224], out[416], _42635_);
  and g_52682_(_39658_, out[427], _42636_);
  xor g_52683_(out[230], out[422], _42637_);
  xor g_52684_(out[234], out[426], _42638_);
  xor g_52685_(out[229], out[421], _42640_);
  xor g_52686_(out[239], out[431], _42641_);
  xor g_52687_(out[237], out[429], _42642_);
  xor g_52688_(out[232], out[424], _42643_);
  or g_52689_(_42630_, _42632_, _42644_);
  or g_52690_(_42642_, _42643_, _42645_);
  or g_52691_(_42633_, _42638_, _42646_);
  or g_52692_(_42645_, _42646_, _42647_);
  or g_52693_(_42631_, _42634_, _42648_);
  or g_52694_(_42635_, _42640_, _42649_);
  or g_52695_(_42648_, _42649_, _42651_);
  or g_52696_(_42647_, _42651_, _42652_);
  xor g_52697_(out[236], out[428], _42653_);
  or g_52698_(_42636_, _42653_, _42654_);
  xor g_52699_(out[231], out[423], _42655_);
  or g_52700_(_42637_, _42655_, _42656_);
  or g_52701_(_42654_, _42656_, _42657_);
  or g_52702_(_42627_, _42629_, _42658_);
  or g_52703_(_42641_, _42658_, _42659_);
  or g_52704_(_42657_, _42659_, _42660_);
  or g_52705_(_42652_, _42660_, _42662_);
  or g_52706_(_42644_, _42662_, _42663_);
  not g_52707_(_42663_, _42664_);
  xor g_52708_(out[215], out[423], _42665_);
  and g_52709_(_39647_, out[427], _42666_);
  xor g_52710_(out[222], out[430], _42667_);
  xor g_52711_(out[216], out[424], _42668_);
  xor g_52712_(out[209], out[417], _42669_);
  xor g_52713_(out[221], out[429], _42670_);
  xor g_52714_(out[217], out[425], _42671_);
  xor g_52715_(out[212], out[420], _42673_);
  xor g_52716_(out[210], out[418], _42674_);
  and g_52717_(out[219], _39790_, _42675_);
  xor g_52718_(out[211], out[419], _42676_);
  xor g_52719_(out[214], out[422], _42677_);
  xor g_52720_(out[223], out[431], _42678_);
  xor g_52721_(out[218], out[426], _42679_);
  xor g_52722_(out[213], out[421], _42680_);
  xor g_52723_(out[208], out[416], _42681_);
  or g_52724_(_42667_, _42673_, _42682_);
  or g_52725_(_42668_, _42670_, _42684_);
  or g_52726_(_42674_, _42679_, _42685_);
  or g_52727_(_42684_, _42685_, _42686_);
  or g_52728_(_42671_, _42676_, _42687_);
  or g_52729_(_42680_, _42681_, _42688_);
  or g_52730_(_42687_, _42688_, _42689_);
  or g_52731_(_42686_, _42689_, _42690_);
  xor g_52732_(out[220], out[428], _42691_);
  or g_52733_(_42666_, _42691_, _42692_);
  or g_52734_(_42665_, _42677_, _42693_);
  or g_52735_(_42692_, _42693_, _42695_);
  or g_52736_(_42669_, _42675_, _42696_);
  or g_52737_(_42678_, _42696_, _42697_);
  or g_52738_(_42695_, _42697_, _42698_);
  or g_52739_(_42690_, _42698_, _42699_);
  or g_52740_(_42682_, _42699_, _42700_);
  xor g_52741_(out[193], out[417], _42701_);
  and g_52742_(_39636_, out[427], _42702_);
  and g_52743_(out[203], _39790_, _42703_);
  xor g_52744_(out[201], out[425], _42704_);
  xor g_52745_(out[192], out[416], _42706_);
  xor g_52746_(out[206], out[430], _42707_);
  xor g_52747_(out[196], out[420], _42708_);
  or g_52748_(_42707_, _42708_, _42709_);
  xor g_52749_(out[205], out[429], _42710_);
  xor g_52750_(out[195], out[419], _42711_);
  xor g_52751_(out[204], out[428], _42712_);
  xor g_52752_(out[198], out[422], _42713_);
  xor g_52753_(out[202], out[426], _42714_);
  xor g_52754_(out[197], out[421], _42715_);
  xor g_52755_(out[207], out[431], _42717_);
  xor g_52756_(out[200], out[424], _42718_);
  or g_52757_(_42710_, _42718_, _42719_);
  xor g_52758_(out[194], out[418], _42720_);
  or g_52759_(_42714_, _42720_, _42721_);
  or g_52760_(_42719_, _42721_, _42722_);
  or g_52761_(_42704_, _42711_, _42723_);
  or g_52762_(_42715_, _42723_, _42724_);
  or g_52763_(_42722_, _42724_, _42725_);
  or g_52764_(_42709_, _42725_, _42726_);
  or g_52765_(_42702_, _42712_, _42728_);
  xor g_52766_(out[199], out[423], _42729_);
  or g_52767_(_42713_, _42729_, _42730_);
  or g_52768_(_42728_, _42730_, _42731_);
  or g_52769_(_42701_, _42703_, _42732_);
  or g_52770_(_42717_, _42732_, _42733_);
  or g_52771_(_42731_, _42733_, _42734_);
  or g_52772_(_42706_, _42734_, _42735_);
  or g_52773_(_42726_, _42735_, _42736_);
  not g_52774_(_42736_, _42737_);
  xor g_52775_(out[183], out[423], _42739_);
  and g_52776_(_39625_, out[427], _42740_);
  xor g_52777_(out[190], out[430], _42741_);
  xor g_52778_(out[184], out[424], _42742_);
  xor g_52779_(out[177], out[417], _42743_);
  xor g_52780_(out[189], out[429], _42744_);
  xor g_52781_(out[185], out[425], _42745_);
  xor g_52782_(out[180], out[420], _42746_);
  xor g_52783_(out[178], out[418], _42747_);
  and g_52784_(out[187], _39790_, _42748_);
  xor g_52785_(out[179], out[419], _42750_);
  xor g_52786_(out[182], out[422], _42751_);
  xor g_52787_(out[191], out[431], _42752_);
  xor g_52788_(out[186], out[426], _42753_);
  xor g_52789_(out[181], out[421], _42754_);
  xor g_52790_(out[176], out[416], _42755_);
  or g_52791_(_42741_, _42746_, _42756_);
  or g_52792_(_42742_, _42744_, _42757_);
  or g_52793_(_42747_, _42753_, _42758_);
  or g_52794_(_42757_, _42758_, _42759_);
  or g_52795_(_42745_, _42750_, _42761_);
  or g_52796_(_42754_, _42755_, _42762_);
  or g_52797_(_42761_, _42762_, _42763_);
  or g_52798_(_42759_, _42763_, _42764_);
  xor g_52799_(out[188], out[428], _42765_);
  or g_52800_(_42740_, _42765_, _42766_);
  or g_52801_(_42739_, _42751_, _42767_);
  or g_52802_(_42766_, _42767_, _42768_);
  or g_52803_(_42743_, _42748_, _42769_);
  or g_52804_(_42752_, _42769_, _42770_);
  or g_52805_(_42768_, _42770_, _42772_);
  or g_52806_(_42764_, _42772_, _42773_);
  or g_52807_(_42756_, _42773_, _42774_);
  not g_52808_(_42774_, _42775_);
  xor g_52809_(out[161], out[417], _42776_);
  and g_52810_(out[171], _39790_, _42777_);
  xor g_52811_(out[169], out[425], _42778_);
  xor g_52812_(out[160], out[416], _42779_);
  xor g_52813_(out[174], out[430], _42780_);
  xor g_52814_(out[164], out[420], _42781_);
  or g_52815_(_42780_, _42781_, _42783_);
  xor g_52816_(out[173], out[429], _42784_);
  xor g_52817_(out[163], out[419], _42785_);
  and g_52818_(_39614_, out[427], _42786_);
  xor g_52819_(out[166], out[422], _42787_);
  xor g_52820_(out[170], out[426], _42788_);
  xor g_52821_(out[165], out[421], _42789_);
  xor g_52822_(out[175], out[431], _42790_);
  xor g_52823_(out[168], out[424], _42791_);
  or g_52824_(_42784_, _42791_, _42792_);
  xor g_52825_(out[162], out[418], _42794_);
  or g_52826_(_42788_, _42794_, _42795_);
  or g_52827_(_42792_, _42795_, _42796_);
  or g_52828_(_42778_, _42785_, _42797_);
  or g_52829_(_42789_, _42797_, _42798_);
  or g_52830_(_42796_, _42798_, _42799_);
  or g_52831_(_42783_, _42799_, _42800_);
  xor g_52832_(out[172], out[428], _42801_);
  or g_52833_(_42786_, _42801_, _42802_);
  xor g_52834_(out[167], out[423], _42803_);
  or g_52835_(_42787_, _42803_, _42805_);
  or g_52836_(_42802_, _42805_, _42806_);
  or g_52837_(_42776_, _42777_, _42807_);
  or g_52838_(_42790_, _42807_, _42808_);
  or g_52839_(_42806_, _42808_, _42809_);
  or g_52840_(_42779_, _42809_, _42810_);
  or g_52841_(_42800_, _42810_, _42811_);
  xor g_52842_(out[151], out[423], _42812_);
  and g_52843_(_39603_, out[427], _42813_);
  xor g_52844_(out[158], out[430], _42814_);
  xor g_52845_(out[152], out[424], _42816_);
  xor g_52846_(out[145], out[417], _42817_);
  xor g_52847_(out[157], out[429], _42818_);
  xor g_52848_(out[153], out[425], _42819_);
  xor g_52849_(out[148], out[420], _42820_);
  xor g_52850_(out[146], out[418], _42821_);
  and g_52851_(out[155], _39790_, _42822_);
  xor g_52852_(out[147], out[419], _42823_);
  xor g_52853_(out[150], out[422], _42824_);
  xor g_52854_(out[159], out[431], _42825_);
  xor g_52855_(out[154], out[426], _42827_);
  xor g_52856_(out[149], out[421], _42828_);
  xor g_52857_(out[144], out[416], _42829_);
  or g_52858_(_42814_, _42820_, _42830_);
  or g_52859_(_42816_, _42818_, _42831_);
  or g_52860_(_42821_, _42827_, _42832_);
  or g_52861_(_42831_, _42832_, _42833_);
  or g_52862_(_42819_, _42823_, _42834_);
  or g_52863_(_42828_, _42829_, _42835_);
  or g_52864_(_42834_, _42835_, _42836_);
  or g_52865_(_42833_, _42836_, _42838_);
  xor g_52866_(out[156], out[428], _42839_);
  or g_52867_(_42813_, _42839_, _42840_);
  or g_52868_(_42812_, _42824_, _42841_);
  or g_52869_(_42840_, _42841_, _42842_);
  or g_52870_(_42817_, _42822_, _42843_);
  or g_52871_(_42825_, _42843_, _42844_);
  or g_52872_(_42842_, _42844_, _42845_);
  or g_52873_(_42838_, _42845_, _42846_);
  or g_52874_(_42830_, _42846_, _42847_);
  xor g_52875_(out[129], out[417], _42849_);
  and g_52876_(out[139], _39790_, _42850_);
  xor g_52877_(out[142], out[430], _42851_);
  xor g_52878_(out[131], out[419], _42852_);
  xor g_52879_(out[132], out[420], _42853_);
  xor g_52880_(out[130], out[418], _42854_);
  xor g_52881_(out[137], out[425], _42855_);
  xor g_52882_(out[128], out[416], _42856_);
  and g_52883_(_39592_, out[427], _42857_);
  xor g_52884_(out[134], out[422], _42858_);
  xor g_52885_(out[138], out[426], _42860_);
  xor g_52886_(out[133], out[421], _42861_);
  xor g_52887_(out[143], out[431], _42862_);
  xor g_52888_(out[141], out[429], _42863_);
  xor g_52889_(out[136], out[424], _42864_);
  or g_52890_(_42851_, _42853_, _42865_);
  or g_52891_(_42863_, _42864_, _42866_);
  or g_52892_(_42854_, _42860_, _42867_);
  or g_52893_(_42866_, _42867_, _42868_);
  or g_52894_(_42852_, _42855_, _42869_);
  or g_52895_(_42856_, _42861_, _42871_);
  or g_52896_(_42869_, _42871_, _42872_);
  or g_52897_(_42868_, _42872_, _42873_);
  xor g_52898_(out[140], out[428], _42874_);
  or g_52899_(_42857_, _42874_, _42875_);
  xor g_52900_(out[135], out[423], _42876_);
  or g_52901_(_42858_, _42876_, _42877_);
  or g_52902_(_42875_, _42877_, _42878_);
  or g_52903_(_42849_, _42850_, _42879_);
  or g_52904_(_42862_, _42879_, _42880_);
  or g_52905_(_42878_, _42880_, _42882_);
  or g_52906_(_42873_, _42882_, _42883_);
  or g_52907_(_42865_, _42883_, _42884_);
  xor g_52908_(out[119], out[423], _42885_);
  and g_52909_(_39581_, out[427], _42886_);
  xor g_52910_(out[126], out[430], _42887_);
  xor g_52911_(out[120], out[424], _42888_);
  xor g_52912_(out[113], out[417], _42889_);
  xor g_52913_(out[125], out[429], _42890_);
  xor g_52914_(out[121], out[425], _42891_);
  xor g_52915_(out[116], out[420], _42893_);
  xor g_52916_(out[114], out[418], _42894_);
  and g_52917_(out[123], _39790_, _42895_);
  xor g_52918_(out[115], out[419], _42896_);
  xor g_52919_(out[118], out[422], _42897_);
  xor g_52920_(out[127], out[431], _42898_);
  xor g_52921_(out[122], out[426], _42899_);
  xor g_52922_(out[117], out[421], _42900_);
  xor g_52923_(out[112], out[416], _42901_);
  or g_52924_(_42887_, _42893_, _42902_);
  or g_52925_(_42888_, _42890_, _42904_);
  or g_52926_(_42894_, _42899_, _42905_);
  or g_52927_(_42904_, _42905_, _42906_);
  or g_52928_(_42891_, _42896_, _42907_);
  or g_52929_(_42900_, _42901_, _42908_);
  or g_52930_(_42907_, _42908_, _42909_);
  or g_52931_(_42906_, _42909_, _42910_);
  xor g_52932_(out[124], out[428], _42911_);
  or g_52933_(_42886_, _42911_, _42912_);
  or g_52934_(_42885_, _42897_, _42913_);
  or g_52935_(_42912_, _42913_, _42915_);
  or g_52936_(_42889_, _42895_, _42916_);
  or g_52937_(_42898_, _42916_, _42917_);
  or g_52938_(_42915_, _42917_, _42918_);
  or g_52939_(_42910_, _42918_, _42919_);
  or g_52940_(_42902_, _42919_, _42920_);
  xor g_52941_(out[104], out[424], _42921_);
  xor g_52942_(out[101], out[421], _42922_);
  xor g_52943_(out[99], out[419], _42923_);
  xor g_52944_(out[110], out[430], _42924_);
  xor g_52945_(out[109], out[429], _42926_);
  xor g_52946_(out[98], out[418], _42927_);
  xor g_52947_(out[105], out[425], _42928_);
  xor g_52948_(out[102], out[422], _42929_);
  xor g_52949_(out[111], out[431], _42930_);
  xor g_52950_(out[106], out[426], _42931_);
  xor g_52951_(out[100], out[420], _42932_);
  xor g_52952_(out[96], out[416], _42933_);
  and g_52953_(_39570_, out[427], _42934_);
  and g_52954_(out[107], _39790_, _42935_);
  or g_52955_(_42921_, _42926_, _42937_);
  xor g_52956_(out[97], out[417], _42938_);
  or g_52957_(_42927_, _42931_, _42939_);
  or g_52958_(_42937_, _42939_, _42940_);
  or g_52959_(_42923_, _42928_, _42941_);
  or g_52960_(_42922_, _42941_, _42942_);
  or g_52961_(_42940_, _42942_, _42943_);
  or g_52962_(_42924_, _42932_, _42944_);
  or g_52963_(_42943_, _42944_, _42945_);
  xor g_52964_(out[108], out[428], _42946_);
  or g_52965_(_42934_, _42946_, _42948_);
  xor g_52966_(out[103], out[423], _42949_);
  or g_52967_(_42929_, _42949_, _42950_);
  or g_52968_(_42948_, _42950_, _42951_);
  or g_52969_(_42935_, _42938_, _42952_);
  or g_52970_(_42930_, _42952_, _42953_);
  or g_52971_(_42951_, _42953_, _42954_);
  or g_52972_(_42933_, _42954_, _42955_);
  or g_52973_(_42945_, _42955_, _42956_);
  not g_52974_(_42956_, _42957_);
  xor g_52975_(out[87], out[423], _42959_);
  and g_52976_(_39559_, out[427], _42960_);
  xor g_52977_(out[94], out[430], _42961_);
  xor g_52978_(out[88], out[424], _42962_);
  xor g_52979_(out[81], out[417], _42963_);
  xor g_52980_(out[93], out[429], _42964_);
  xor g_52981_(out[89], out[425], _42965_);
  xor g_52982_(out[84], out[420], _42966_);
  xor g_52983_(out[82], out[418], _42967_);
  and g_52984_(out[91], _39790_, _42968_);
  xor g_52985_(out[83], out[419], _42970_);
  xor g_52986_(out[86], out[422], _42971_);
  xor g_52987_(out[95], out[431], _42972_);
  xor g_52988_(out[90], out[426], _42973_);
  xor g_52989_(out[85], out[421], _42974_);
  xor g_52990_(out[80], out[416], _42975_);
  or g_52991_(_42961_, _42966_, _42976_);
  or g_52992_(_42962_, _42964_, _42977_);
  or g_52993_(_42967_, _42973_, _42978_);
  or g_52994_(_42977_, _42978_, _42979_);
  or g_52995_(_42965_, _42970_, _42981_);
  or g_52996_(_42974_, _42975_, _42982_);
  or g_52997_(_42981_, _42982_, _42983_);
  or g_52998_(_42979_, _42983_, _42984_);
  xor g_52999_(out[92], out[428], _42985_);
  or g_53000_(_42960_, _42985_, _42986_);
  or g_53001_(_42959_, _42971_, _42987_);
  or g_53002_(_42986_, _42987_, _42988_);
  or g_53003_(_42963_, _42968_, _42989_);
  or g_53004_(_42972_, _42989_, _42990_);
  or g_53005_(_42988_, _42990_, _42992_);
  or g_53006_(_42984_, _42992_, _42993_);
  or g_53007_(_42976_, _42993_, _42994_);
  not g_53008_(_42994_, _42995_);
  xor g_53009_(out[65], out[417], _42996_);
  and g_53010_(out[75], _39790_, _42997_);
  xor g_53011_(out[73], out[425], _42998_);
  xor g_53012_(out[64], out[416], _42999_);
  xor g_53013_(out[78], out[430], _43000_);
  xor g_53014_(out[68], out[420], _43001_);
  or g_53015_(_43000_, _43001_, _43003_);
  xor g_53016_(out[77], out[429], _43004_);
  xor g_53017_(out[67], out[419], _43005_);
  and g_53018_(_39548_, out[427], _43006_);
  xor g_53019_(out[70], out[422], _43007_);
  xor g_53020_(out[74], out[426], _43008_);
  xor g_53021_(out[69], out[421], _43009_);
  xor g_53022_(out[79], out[431], _43010_);
  xor g_53023_(out[72], out[424], _43011_);
  or g_53024_(_43004_, _43011_, _43012_);
  xor g_53025_(out[66], out[418], _43014_);
  or g_53026_(_43008_, _43014_, _43015_);
  or g_53027_(_43012_, _43015_, _43016_);
  or g_53028_(_42998_, _43005_, _43017_);
  or g_53029_(_43009_, _43017_, _43018_);
  or g_53030_(_43016_, _43018_, _43019_);
  or g_53031_(_43003_, _43019_, _43020_);
  xor g_53032_(out[76], out[428], _43021_);
  or g_53033_(_43006_, _43021_, _43022_);
  xor g_53034_(out[71], out[423], _43023_);
  or g_53035_(_43007_, _43023_, _43025_);
  or g_53036_(_43022_, _43025_, _43026_);
  or g_53037_(_42996_, _42997_, _43027_);
  or g_53038_(_43010_, _43027_, _43028_);
  or g_53039_(_43026_, _43028_, _43029_);
  or g_53040_(_42999_, _43029_, _43030_);
  or g_53041_(_43020_, _43030_, _43031_);
  xor g_53042_(out[55], out[423], _43032_);
  and g_53043_(_39537_, out[427], _43033_);
  xor g_53044_(out[62], out[430], _43034_);
  xor g_53045_(out[56], out[424], _43036_);
  xor g_53046_(out[49], out[417], _43037_);
  xor g_53047_(out[61], out[429], _43038_);
  xor g_53048_(out[57], out[425], _43039_);
  xor g_53049_(out[52], out[420], _43040_);
  xor g_53050_(out[50], out[418], _43041_);
  and g_53051_(out[59], _39790_, _43042_);
  xor g_53052_(out[51], out[419], _43043_);
  xor g_53053_(out[54], out[422], _43044_);
  xor g_53054_(out[63], out[431], _43045_);
  xor g_53055_(out[58], out[426], _43047_);
  xor g_53056_(out[53], out[421], _43048_);
  xor g_53057_(out[48], out[416], _43049_);
  or g_53058_(_43034_, _43040_, _43050_);
  or g_53059_(_43036_, _43038_, _43051_);
  or g_53060_(_43041_, _43047_, _43052_);
  or g_53061_(_43051_, _43052_, _43053_);
  or g_53062_(_43039_, _43043_, _43054_);
  or g_53063_(_43048_, _43049_, _43055_);
  or g_53064_(_43054_, _43055_, _43056_);
  or g_53065_(_43053_, _43056_, _43058_);
  xor g_53066_(out[60], out[428], _43059_);
  or g_53067_(_43033_, _43059_, _43060_);
  or g_53068_(_43032_, _43044_, _43061_);
  or g_53069_(_43060_, _43061_, _43062_);
  or g_53070_(_43037_, _43042_, _43063_);
  or g_53071_(_43045_, _43063_, _43064_);
  or g_53072_(_43062_, _43064_, _43065_);
  or g_53073_(_43058_, _43065_, _43066_);
  or g_53074_(_43050_, _43066_, _43067_);
  xor g_53075_(out[45], out[429], _43069_);
  xor g_53076_(out[34], out[418], _43070_);
  xor g_53077_(out[37], out[421], _43071_);
  xor g_53078_(out[41], out[425], _43072_);
  xor g_53079_(out[36], out[420], _43073_);
  xor g_53080_(out[40], out[424], _43074_);
  xor g_53081_(out[46], out[430], _43075_);
  xor g_53082_(out[38], out[422], _43076_);
  xor g_53083_(out[47], out[431], _43077_);
  xor g_53084_(out[42], out[426], _43078_);
  xor g_53085_(out[32], out[416], _43080_);
  xor g_53086_(out[35], out[419], _43081_);
  and g_53087_(_39526_, out[427], _43082_);
  and g_53088_(out[43], _39790_, _43083_);
  xor g_53089_(out[33], out[417], _43084_);
  or g_53090_(_43073_, _43075_, _43085_);
  or g_53091_(_43069_, _43074_, _43086_);
  or g_53092_(_43070_, _43078_, _43087_);
  or g_53093_(_43086_, _43087_, _43088_);
  or g_53094_(_43072_, _43081_, _43089_);
  or g_53095_(_43071_, _43080_, _43091_);
  or g_53096_(_43089_, _43091_, _43092_);
  or g_53097_(_43088_, _43092_, _43093_);
  xor g_53098_(out[44], out[428], _43094_);
  or g_53099_(_43082_, _43094_, _43095_);
  xor g_53100_(out[39], out[423], _43096_);
  or g_53101_(_43076_, _43096_, _43097_);
  or g_53102_(_43095_, _43097_, _43098_);
  or g_53103_(_43083_, _43084_, _43099_);
  or g_53104_(_43077_, _43099_, _43100_);
  or g_53105_(_43098_, _43100_, _43102_);
  or g_53106_(_43093_, _43102_, _43103_);
  or g_53107_(_43085_, _43103_, _43104_);
  not g_53108_(_43104_, _43105_);
  xor g_53109_(out[23], out[423], _43106_);
  and g_53110_(_39493_, out[427], _43107_);
  xor g_53111_(out[30], out[430], _43108_);
  xor g_53112_(out[24], out[424], _43109_);
  xor g_53113_(out[17], out[417], _43110_);
  xor g_53114_(out[29], out[429], _43111_);
  xor g_53115_(out[25], out[425], _43113_);
  xor g_53116_(out[20], out[420], _43114_);
  xor g_53117_(out[18], out[418], _43115_);
  and g_53118_(out[27], _39790_, _43116_);
  xor g_53119_(out[19], out[419], _43117_);
  xor g_53120_(out[22], out[422], _43118_);
  xor g_53121_(out[31], out[431], _43119_);
  xor g_53122_(out[26], out[426], _43120_);
  xor g_53123_(out[21], out[421], _43121_);
  xor g_53124_(out[16], out[416], _43122_);
  or g_53125_(_43108_, _43114_, _43124_);
  or g_53126_(_43109_, _43111_, _43125_);
  or g_53127_(_43115_, _43120_, _43126_);
  or g_53128_(_43125_, _43126_, _43127_);
  or g_53129_(_43113_, _43117_, _43128_);
  or g_53130_(_43121_, _43122_, _43129_);
  or g_53131_(_43128_, _43129_, _43130_);
  or g_53132_(_43127_, _43130_, _43131_);
  xor g_53133_(out[28], out[428], _43132_);
  or g_53134_(_43107_, _43132_, _43133_);
  or g_53135_(_43106_, _43118_, _43135_);
  or g_53136_(_43133_, _43135_, _43136_);
  or g_53137_(_43110_, _43116_, _43137_);
  or g_53138_(_43119_, _43137_, _43138_);
  or g_53139_(_43136_, _43138_, _43139_);
  or g_53140_(_43131_, _43139_, _43140_);
  or g_53141_(_43124_, _43140_, _43141_);
  xor g_53142_(out[12], out[428], _43142_);
  and g_53143_(_39438_, out[427], _43143_);
  xor g_53144_(out[8], out[424], _43144_);
  xor g_53145_(out[6], out[422], _21890_);
  xor g_53146_(out[13], out[429], _21891_);
  xor g_53147_(out[14], out[430], _21892_);
  xor g_53148_(out[2], out[418], _21893_);
  xor g_53149_(out[9], out[425], _21894_);
  xor g_53150_(out[5], out[421], _21895_);
  xor g_53151_(out[1], out[417], _21896_);
  and g_53152_(out[11], _39790_, _21897_);
  or g_53153_(_43144_, _21891_, _21898_);
  xor g_53154_(out[15], out[431], _21899_);
  xor g_53155_(out[10], out[426], _21901_);
  xor g_53156_(out[4], out[420], _21902_);
  xor g_53157_(out[3], out[419], _21903_);
  xor g_53158_(out[0], out[416], _21904_);
  or g_53159_(_21893_, _21901_, _21905_);
  or g_53160_(_21898_, _21905_, _21906_);
  or g_53161_(_21894_, _21903_, _21907_);
  or g_53162_(_21895_, _21907_, _21908_);
  or g_53163_(_21906_, _21908_, _21909_);
  or g_53164_(_21892_, _21902_, _21910_);
  or g_53165_(_21909_, _21910_, _21912_);
  or g_53166_(_43142_, _43143_, _21913_);
  xor g_53167_(out[7], out[423], _21914_);
  or g_53168_(_21890_, _21914_, _21915_);
  or g_53169_(_21913_, _21915_, _21916_);
  or g_53170_(_21896_, _21897_, _21917_);
  or g_53171_(_21899_, _21917_, _21918_);
  or g_53172_(_21916_, _21918_, _21919_);
  or g_53173_(_21904_, _21919_, _21920_);
  or g_53174_(_21912_, _21920_, _21921_);
  xor g_53175_(out[307], out[403], _21923_);
  xor g_53176_(out[308], out[404], _21924_);
  xor g_53177_(out[318], out[414], _21925_);
  xor g_53178_(out[306], out[402], _21926_);
  xor g_53179_(out[309], out[405], _21927_);
  xor g_53180_(out[313], out[409], _21928_);
  xor g_53181_(out[312], out[408], _21929_);
  xor g_53182_(out[319], out[415], _21930_);
  xor g_53183_(out[314], out[410], _21931_);
  xor g_53184_(out[310], out[406], _21932_);
  xor g_53185_(out[304], out[400], _21934_);
  and g_53186_(_39724_, out[411], _21935_);
  and g_53187_(out[315], _39779_, _21936_);
  xor g_53188_(out[317], out[413], _21937_);
  or g_53189_(_21929_, _21937_, _21938_);
  xor g_53190_(out[305], out[401], _21939_);
  or g_53191_(_21926_, _21931_, _21940_);
  or g_53192_(_21938_, _21940_, _21941_);
  or g_53193_(_21923_, _21928_, _21942_);
  or g_53194_(_21927_, _21942_, _21943_);
  or g_53195_(_21941_, _21943_, _21945_);
  or g_53196_(_21924_, _21925_, _21946_);
  or g_53197_(_21945_, _21946_, _21947_);
  xor g_53198_(out[316], out[412], _21948_);
  or g_53199_(_21935_, _21948_, _21949_);
  xor g_53200_(out[311], out[407], _21950_);
  or g_53201_(_21932_, _21950_, _21951_);
  or g_53202_(_21949_, _21951_, _21952_);
  or g_53203_(_21936_, _21939_, _21953_);
  or g_53204_(_21930_, _21953_, _21954_);
  or g_53205_(_21952_, _21954_, _21956_);
  or g_53206_(_21934_, _21956_, _21957_);
  or g_53207_(_21947_, _21957_, _21958_);
  not g_53208_(_21958_, _21959_);
  xor g_53209_(out[295], out[407], _21960_);
  and g_53210_(_39702_, out[411], _21961_);
  xor g_53211_(out[302], out[414], _21962_);
  xor g_53212_(out[296], out[408], _21963_);
  xor g_53213_(out[289], out[401], _21964_);
  xor g_53214_(out[301], out[413], _21965_);
  xor g_53215_(out[297], out[409], _21967_);
  xor g_53216_(out[292], out[404], _21968_);
  xor g_53217_(out[290], out[402], _21969_);
  and g_53218_(out[299], _39779_, _21970_);
  xor g_53219_(out[291], out[403], _21971_);
  xor g_53220_(out[294], out[406], _21972_);
  xor g_53221_(out[303], out[415], _21973_);
  xor g_53222_(out[298], out[410], _21974_);
  xor g_53223_(out[293], out[405], _21975_);
  xor g_53224_(out[288], out[400], _21976_);
  or g_53225_(_21962_, _21968_, _21978_);
  or g_53226_(_21963_, _21965_, _21979_);
  or g_53227_(_21969_, _21974_, _21980_);
  or g_53228_(_21979_, _21980_, _21981_);
  or g_53229_(_21967_, _21971_, _21982_);
  or g_53230_(_21975_, _21976_, _21983_);
  or g_53231_(_21982_, _21983_, _21984_);
  or g_53232_(_21981_, _21984_, _21985_);
  xor g_53233_(out[300], out[412], _21986_);
  or g_53234_(_21961_, _21986_, _21987_);
  or g_53235_(_21960_, _21972_, _21989_);
  or g_53236_(_21987_, _21989_, _21990_);
  or g_53237_(_21964_, _21970_, _21991_);
  or g_53238_(_21973_, _21991_, _21992_);
  or g_53239_(_21990_, _21992_, _21993_);
  or g_53240_(_21985_, _21993_, _21994_);
  or g_53241_(_21978_, _21994_, _21995_);
  not g_53242_(_21995_, _21996_);
  xor g_53243_(out[273], out[401], _21997_);
  and g_53244_(out[283], _39779_, _21998_);
  xor g_53245_(out[281], out[409], _22000_);
  xor g_53246_(out[272], out[400], _22001_);
  xor g_53247_(out[286], out[414], _22002_);
  xor g_53248_(out[276], out[404], _22003_);
  or g_53249_(_22002_, _22003_, _22004_);
  xor g_53250_(out[285], out[413], _22005_);
  xor g_53251_(out[275], out[403], _22006_);
  and g_53252_(_39691_, out[411], _22007_);
  xor g_53253_(out[278], out[406], _22008_);
  xor g_53254_(out[282], out[410], _22009_);
  xor g_53255_(out[277], out[405], _22011_);
  xor g_53256_(out[287], out[415], _22012_);
  xor g_53257_(out[280], out[408], _22013_);
  or g_53258_(_22005_, _22013_, _22014_);
  xor g_53259_(out[274], out[402], _22015_);
  or g_53260_(_22009_, _22015_, _22016_);
  or g_53261_(_22014_, _22016_, _22017_);
  or g_53262_(_22000_, _22006_, _22018_);
  or g_53263_(_22011_, _22018_, _22019_);
  or g_53264_(_22017_, _22019_, _22020_);
  or g_53265_(_22004_, _22020_, _22022_);
  xor g_53266_(out[284], out[412], _22023_);
  or g_53267_(_22007_, _22023_, _22024_);
  xor g_53268_(out[279], out[407], _22025_);
  or g_53269_(_22008_, _22025_, _22026_);
  or g_53270_(_22024_, _22026_, _22027_);
  or g_53271_(_21997_, _21998_, _22028_);
  or g_53272_(_22012_, _22028_, _22029_);
  or g_53273_(_22027_, _22029_, _22030_);
  or g_53274_(_22001_, _22030_, _22031_);
  or g_53275_(_22022_, _22031_, _22033_);
  not g_53276_(_22033_, _22034_);
  xor g_53277_(out[263], out[407], _22035_);
  and g_53278_(_39680_, out[411], _22036_);
  xor g_53279_(out[270], out[414], _22037_);
  xor g_53280_(out[264], out[408], _22038_);
  xor g_53281_(out[257], out[401], _22039_);
  xor g_53282_(out[269], out[413], _22040_);
  xor g_53283_(out[265], out[409], _22041_);
  xor g_53284_(out[260], out[404], _22042_);
  xor g_53285_(out[258], out[402], _22044_);
  and g_53286_(out[267], _39779_, _22045_);
  xor g_53287_(out[259], out[403], _22046_);
  xor g_53288_(out[262], out[406], _22047_);
  xor g_53289_(out[271], out[415], _22048_);
  xor g_53290_(out[266], out[410], _22049_);
  xor g_53291_(out[261], out[405], _22050_);
  xor g_53292_(out[256], out[400], _22051_);
  or g_53293_(_22037_, _22042_, _22052_);
  or g_53294_(_22038_, _22040_, _22053_);
  or g_53295_(_22044_, _22049_, _22055_);
  or g_53296_(_22053_, _22055_, _22056_);
  or g_53297_(_22041_, _22046_, _22057_);
  or g_53298_(_22050_, _22051_, _22058_);
  or g_53299_(_22057_, _22058_, _22059_);
  or g_53300_(_22056_, _22059_, _22060_);
  xor g_53301_(out[268], out[412], _22061_);
  or g_53302_(_22036_, _22061_, _22062_);
  or g_53303_(_22035_, _22047_, _22063_);
  or g_53304_(_22062_, _22063_, _22064_);
  or g_53305_(_22039_, _22045_, _22066_);
  or g_53306_(_22048_, _22066_, _22067_);
  or g_53307_(_22064_, _22067_, _22068_);
  or g_53308_(_22060_, _22068_, _22069_);
  or g_53309_(_22052_, _22069_, _22070_);
  and g_53310_(out[251], _39779_, _22071_);
  and g_53311_(_39669_, out[411], _22072_);
  xor g_53312_(out[241], out[401], _22073_);
  xor g_53313_(out[243], out[403], _22074_);
  xor g_53314_(out[247], out[407], _22075_);
  xor g_53315_(out[249], out[409], _22077_);
  xor g_53316_(out[255], out[415], _22078_);
  xor g_53317_(out[242], out[402], _22079_);
  xor g_53318_(out[254], out[414], _22080_);
  xor g_53319_(out[253], out[413], _22081_);
  xor g_53320_(out[248], out[408], _22082_);
  or g_53321_(_22081_, _22082_, _22083_);
  xor g_53322_(out[244], out[404], _22084_);
  xor g_53323_(out[246], out[406], _22085_);
  xor g_53324_(out[250], out[410], _22086_);
  xor g_53325_(out[245], out[405], _22088_);
  xor g_53326_(out[240], out[400], _22089_);
  or g_53327_(_22079_, _22086_, _22090_);
  or g_53328_(_22083_, _22090_, _22091_);
  or g_53329_(_22074_, _22077_, _22092_);
  or g_53330_(_22088_, _22092_, _22093_);
  or g_53331_(_22091_, _22093_, _22094_);
  or g_53332_(_22080_, _22084_, _22095_);
  or g_53333_(_22094_, _22095_, _22096_);
  xor g_53334_(out[252], out[412], _22097_);
  or g_53335_(_22072_, _22097_, _22099_);
  or g_53336_(_22075_, _22085_, _22100_);
  or g_53337_(_22099_, _22100_, _22101_);
  or g_53338_(_22071_, _22073_, _22102_);
  or g_53339_(_22078_, _22102_, _22103_);
  or g_53340_(_22101_, _22103_, _22104_);
  or g_53341_(_22089_, _22104_, _22105_);
  or g_53342_(_22096_, _22105_, _22106_);
  not g_53343_(_22106_, _22107_);
  xor g_53344_(out[231], out[407], _22108_);
  and g_53345_(_39658_, out[411], _22110_);
  xor g_53346_(out[238], out[414], _22111_);
  xor g_53347_(out[232], out[408], _22112_);
  xor g_53348_(out[225], out[401], _22113_);
  xor g_53349_(out[237], out[413], _22114_);
  xor g_53350_(out[233], out[409], _22115_);
  xor g_53351_(out[228], out[404], _22116_);
  xor g_53352_(out[226], out[402], _22117_);
  and g_53353_(out[235], _39779_, _22118_);
  xor g_53354_(out[227], out[403], _22119_);
  xor g_53355_(out[230], out[406], _22121_);
  xor g_53356_(out[239], out[415], _22122_);
  xor g_53357_(out[234], out[410], _22123_);
  xor g_53358_(out[229], out[405], _22124_);
  xor g_53359_(out[224], out[400], _22125_);
  or g_53360_(_22111_, _22116_, _22126_);
  or g_53361_(_22112_, _22114_, _22127_);
  or g_53362_(_22117_, _22123_, _22128_);
  or g_53363_(_22127_, _22128_, _22129_);
  or g_53364_(_22115_, _22119_, _22130_);
  or g_53365_(_22124_, _22125_, _22132_);
  or g_53366_(_22130_, _22132_, _22133_);
  or g_53367_(_22129_, _22133_, _22134_);
  xor g_53368_(out[236], out[412], _22135_);
  or g_53369_(_22110_, _22135_, _22136_);
  or g_53370_(_22108_, _22121_, _22137_);
  or g_53371_(_22136_, _22137_, _22138_);
  or g_53372_(_22113_, _22118_, _22139_);
  or g_53373_(_22122_, _22139_, _22140_);
  or g_53374_(_22138_, _22140_, _22141_);
  or g_53375_(_22134_, _22141_, _22143_);
  or g_53376_(_22126_, _22143_, _22144_);
  xor g_53377_(out[218], out[410], _22145_);
  xor g_53378_(out[210], out[402], _22146_);
  xor g_53379_(out[209], out[401], _22147_);
  and g_53380_(_39647_, out[411], _22148_);
  and g_53381_(out[219], _39779_, _22149_);
  xor g_53382_(out[221], out[413], _22150_);
  xor g_53383_(out[211], out[403], _22151_);
  xor g_53384_(out[222], out[414], _22152_);
  xor g_53385_(out[220], out[412], _22154_);
  xor g_53386_(out[216], out[408], _22155_);
  xor g_53387_(out[223], out[415], _22156_);
  xor g_53388_(out[213], out[405], _22157_);
  xor g_53389_(out[214], out[406], _22158_);
  xor g_53390_(out[208], out[400], _22159_);
  xor g_53391_(out[212], out[404], _22160_);
  or g_53392_(_22150_, _22155_, _22161_);
  xor g_53393_(out[217], out[409], _22162_);
  or g_53394_(_22145_, _22146_, _22163_);
  or g_53395_(_22161_, _22163_, _22165_);
  or g_53396_(_22151_, _22162_, _22166_);
  or g_53397_(_22157_, _22166_, _22167_);
  or g_53398_(_22165_, _22167_, _22168_);
  or g_53399_(_22152_, _22160_, _22169_);
  or g_53400_(_22168_, _22169_, _22170_);
  or g_53401_(_22148_, _22154_, _22171_);
  xor g_53402_(out[215], out[407], _22172_);
  or g_53403_(_22158_, _22172_, _22173_);
  or g_53404_(_22171_, _22173_, _22174_);
  or g_53405_(_22147_, _22149_, _22176_);
  or g_53406_(_22156_, _22176_, _22177_);
  or g_53407_(_22174_, _22177_, _22178_);
  or g_53408_(_22159_, _22178_, _22179_);
  or g_53409_(_22170_, _22179_, _22180_);
  xor g_53410_(out[199], out[407], _22181_);
  and g_53411_(_39636_, out[411], _22182_);
  xor g_53412_(out[206], out[414], _22183_);
  xor g_53413_(out[200], out[408], _22184_);
  xor g_53414_(out[193], out[401], _22185_);
  xor g_53415_(out[205], out[413], _22187_);
  xor g_53416_(out[201], out[409], _22188_);
  xor g_53417_(out[196], out[404], _22189_);
  xor g_53418_(out[194], out[402], _22190_);
  and g_53419_(out[203], _39779_, _22191_);
  xor g_53420_(out[195], out[403], _22192_);
  xor g_53421_(out[198], out[406], _22193_);
  xor g_53422_(out[207], out[415], _22194_);
  xor g_53423_(out[202], out[410], _22195_);
  xor g_53424_(out[197], out[405], _22196_);
  xor g_53425_(out[192], out[400], _22198_);
  or g_53426_(_22183_, _22189_, _22199_);
  or g_53427_(_22184_, _22187_, _22200_);
  or g_53428_(_22190_, _22195_, _22201_);
  or g_53429_(_22200_, _22201_, _22202_);
  or g_53430_(_22188_, _22192_, _22203_);
  or g_53431_(_22196_, _22198_, _22204_);
  or g_53432_(_22203_, _22204_, _22205_);
  or g_53433_(_22202_, _22205_, _22206_);
  xor g_53434_(out[204], out[412], _22207_);
  or g_53435_(_22182_, _22207_, _22209_);
  or g_53436_(_22181_, _22193_, _22210_);
  or g_53437_(_22209_, _22210_, _22211_);
  or g_53438_(_22185_, _22191_, _22212_);
  or g_53439_(_22194_, _22212_, _22213_);
  or g_53440_(_22211_, _22213_, _22214_);
  or g_53441_(_22206_, _22214_, _22215_);
  or g_53442_(_22199_, _22215_, _22216_);
  not g_53443_(_22216_, _22217_);
  xor g_53444_(out[177], out[401], _22218_);
  and g_53445_(_39625_, out[411], _22220_);
  and g_53446_(out[187], _39779_, _22221_);
  xor g_53447_(out[189], out[413], _22222_);
  xor g_53448_(out[186], out[410], _22223_);
  xor g_53449_(out[184], out[408], _22224_);
  xor g_53450_(out[176], out[400], _22225_);
  xor g_53451_(out[190], out[414], _22226_);
  xor g_53452_(out[181], out[405], _22227_);
  xor g_53453_(out[178], out[402], _22228_);
  xor g_53454_(out[185], out[409], _22229_);
  xor g_53455_(out[179], out[403], _22231_);
  xor g_53456_(out[191], out[415], _22232_);
  xor g_53457_(out[180], out[404], _22233_);
  xor g_53458_(out[182], out[406], _22234_);
  or g_53459_(_22226_, _22233_, _22235_);
  or g_53460_(_22222_, _22224_, _22236_);
  or g_53461_(_22223_, _22228_, _22237_);
  or g_53462_(_22236_, _22237_, _22238_);
  or g_53463_(_22229_, _22231_, _22239_);
  or g_53464_(_22225_, _22227_, _22240_);
  or g_53465_(_22239_, _22240_, _22242_);
  or g_53466_(_22238_, _22242_, _22243_);
  xor g_53467_(out[188], out[412], _22244_);
  or g_53468_(_22220_, _22244_, _22245_);
  xor g_53469_(out[183], out[407], _22246_);
  or g_53470_(_22234_, _22246_, _22247_);
  or g_53471_(_22245_, _22247_, _22248_);
  or g_53472_(_22218_, _22221_, _22249_);
  or g_53473_(_22232_, _22249_, _22250_);
  or g_53474_(_22248_, _22250_, _22251_);
  or g_53475_(_22243_, _22251_, _22253_);
  or g_53476_(_22235_, _22253_, _22254_);
  xor g_53477_(out[167], out[407], _22255_);
  and g_53478_(_39614_, out[411], _22256_);
  xor g_53479_(out[174], out[414], _22257_);
  xor g_53480_(out[168], out[408], _22258_);
  xor g_53481_(out[161], out[401], _22259_);
  xor g_53482_(out[173], out[413], _22260_);
  xor g_53483_(out[169], out[409], _22261_);
  xor g_53484_(out[164], out[404], _22262_);
  xor g_53485_(out[162], out[402], _22264_);
  and g_53486_(out[171], _39779_, _22265_);
  xor g_53487_(out[163], out[403], _22266_);
  xor g_53488_(out[166], out[406], _22267_);
  xor g_53489_(out[175], out[415], _22268_);
  xor g_53490_(out[170], out[410], _22269_);
  xor g_53491_(out[165], out[405], _22270_);
  xor g_53492_(out[160], out[400], _22271_);
  or g_53493_(_22257_, _22262_, _22272_);
  or g_53494_(_22258_, _22260_, _22273_);
  or g_53495_(_22264_, _22269_, _22275_);
  or g_53496_(_22273_, _22275_, _22276_);
  or g_53497_(_22261_, _22266_, _22277_);
  or g_53498_(_22270_, _22271_, _22278_);
  or g_53499_(_22277_, _22278_, _22279_);
  or g_53500_(_22276_, _22279_, _22280_);
  xor g_53501_(out[172], out[412], _22281_);
  or g_53502_(_22256_, _22281_, _22282_);
  or g_53503_(_22255_, _22267_, _22283_);
  or g_53504_(_22282_, _22283_, _22284_);
  or g_53505_(_22259_, _22265_, _22286_);
  or g_53506_(_22268_, _22286_, _22287_);
  or g_53507_(_22284_, _22287_, _22288_);
  or g_53508_(_22280_, _22288_, _22289_);
  or g_53509_(_22272_, _22289_, _22290_);
  xor g_53510_(out[145], out[401], _22291_);
  and g_53511_(out[155], _39779_, _22292_);
  xor g_53512_(out[158], out[414], _22293_);
  xor g_53513_(out[147], out[403], _22294_);
  xor g_53514_(out[148], out[404], _22295_);
  xor g_53515_(out[146], out[402], _22297_);
  xor g_53516_(out[153], out[409], _22298_);
  xor g_53517_(out[144], out[400], _22299_);
  and g_53518_(_39603_, out[411], _22300_);
  xor g_53519_(out[150], out[406], _22301_);
  xor g_53520_(out[154], out[410], _22302_);
  xor g_53521_(out[149], out[405], _22303_);
  xor g_53522_(out[159], out[415], _22304_);
  xor g_53523_(out[157], out[413], _22305_);
  xor g_53524_(out[152], out[408], _22306_);
  or g_53525_(_22293_, _22295_, _22308_);
  or g_53526_(_22305_, _22306_, _22309_);
  or g_53527_(_22297_, _22302_, _22310_);
  or g_53528_(_22309_, _22310_, _22311_);
  or g_53529_(_22294_, _22298_, _22312_);
  or g_53530_(_22299_, _22303_, _22313_);
  or g_53531_(_22312_, _22313_, _22314_);
  or g_53532_(_22311_, _22314_, _22315_);
  xor g_53533_(out[156], out[412], _22316_);
  or g_53534_(_22300_, _22316_, _22317_);
  xor g_53535_(out[151], out[407], _22319_);
  or g_53536_(_22301_, _22319_, _22320_);
  or g_53537_(_22317_, _22320_, _22321_);
  or g_53538_(_22291_, _22292_, _22322_);
  or g_53539_(_22304_, _22322_, _22323_);
  or g_53540_(_22321_, _22323_, _22324_);
  or g_53541_(_22315_, _22324_, _22325_);
  or g_53542_(_22308_, _22325_, _22326_);
  xor g_53543_(out[135], out[407], _22327_);
  and g_53544_(_39592_, out[411], _22328_);
  xor g_53545_(out[142], out[414], _22330_);
  xor g_53546_(out[136], out[408], _22331_);
  xor g_53547_(out[129], out[401], _22332_);
  xor g_53548_(out[141], out[413], _22333_);
  xor g_53549_(out[137], out[409], _22334_);
  xor g_53550_(out[132], out[404], _22335_);
  xor g_53551_(out[130], out[402], _22336_);
  and g_53552_(out[139], _39779_, _22337_);
  xor g_53553_(out[131], out[403], _22338_);
  xor g_53554_(out[134], out[406], _22339_);
  xor g_53555_(out[143], out[415], _22341_);
  xor g_53556_(out[138], out[410], _22342_);
  xor g_53557_(out[133], out[405], _22343_);
  xor g_53558_(out[128], out[400], _22344_);
  or g_53559_(_22330_, _22335_, _22345_);
  or g_53560_(_22331_, _22333_, _22346_);
  or g_53561_(_22336_, _22342_, _22347_);
  or g_53562_(_22346_, _22347_, _22348_);
  or g_53563_(_22334_, _22338_, _22349_);
  or g_53564_(_22343_, _22344_, _22350_);
  or g_53565_(_22349_, _22350_, _22352_);
  or g_53566_(_22348_, _22352_, _22353_);
  xor g_53567_(out[140], out[412], _22354_);
  or g_53568_(_22328_, _22354_, _22355_);
  or g_53569_(_22327_, _22339_, _22356_);
  or g_53570_(_22355_, _22356_, _22357_);
  or g_53571_(_22332_, _22337_, _22358_);
  or g_53572_(_22341_, _22358_, _22359_);
  or g_53573_(_22357_, _22359_, _22360_);
  or g_53574_(_22353_, _22360_, _22361_);
  or g_53575_(_22345_, _22361_, _22363_);
  xor g_53576_(out[113], out[401], _22364_);
  and g_53577_(out[123], _39779_, _22365_);
  xor g_53578_(out[121], out[409], _22366_);
  xor g_53579_(out[112], out[400], _22367_);
  xor g_53580_(out[126], out[414], _22368_);
  xor g_53581_(out[116], out[404], _22369_);
  or g_53582_(_22368_, _22369_, _22370_);
  xor g_53583_(out[125], out[413], _22371_);
  xor g_53584_(out[115], out[403], _22372_);
  and g_53585_(_39581_, out[411], _22374_);
  xor g_53586_(out[118], out[406], _22375_);
  xor g_53587_(out[122], out[410], _22376_);
  xor g_53588_(out[117], out[405], _22377_);
  xor g_53589_(out[127], out[415], _22378_);
  xor g_53590_(out[120], out[408], _22379_);
  or g_53591_(_22371_, _22379_, _22380_);
  xor g_53592_(out[114], out[402], _22381_);
  or g_53593_(_22376_, _22381_, _22382_);
  or g_53594_(_22380_, _22382_, _22383_);
  or g_53595_(_22366_, _22372_, _22385_);
  or g_53596_(_22377_, _22385_, _22386_);
  or g_53597_(_22383_, _22386_, _22387_);
  or g_53598_(_22370_, _22387_, _22388_);
  xor g_53599_(out[124], out[412], _22389_);
  or g_53600_(_22374_, _22389_, _22390_);
  xor g_53601_(out[119], out[407], _22391_);
  or g_53602_(_22375_, _22391_, _22392_);
  or g_53603_(_22390_, _22392_, _22393_);
  or g_53604_(_22364_, _22365_, _22394_);
  or g_53605_(_22378_, _22394_, _22396_);
  or g_53606_(_22393_, _22396_, _22397_);
  or g_53607_(_22367_, _22397_, _22398_);
  or g_53608_(_22388_, _22398_, _22399_);
  xor g_53609_(out[103], out[407], _22400_);
  and g_53610_(_39570_, out[411], _22401_);
  xor g_53611_(out[110], out[414], _22402_);
  xor g_53612_(out[104], out[408], _22403_);
  xor g_53613_(out[97], out[401], _22404_);
  xor g_53614_(out[109], out[413], _22405_);
  xor g_53615_(out[105], out[409], _22407_);
  xor g_53616_(out[100], out[404], _22408_);
  xor g_53617_(out[98], out[402], _22409_);
  and g_53618_(out[107], _39779_, _22410_);
  xor g_53619_(out[99], out[403], _22411_);
  xor g_53620_(out[102], out[406], _22412_);
  xor g_53621_(out[111], out[415], _22413_);
  xor g_53622_(out[106], out[410], _22414_);
  xor g_53623_(out[101], out[405], _22415_);
  xor g_53624_(out[96], out[400], _22416_);
  or g_53625_(_22402_, _22408_, _22418_);
  or g_53626_(_22403_, _22405_, _22419_);
  or g_53627_(_22409_, _22414_, _22420_);
  or g_53628_(_22419_, _22420_, _22421_);
  or g_53629_(_22407_, _22411_, _22422_);
  or g_53630_(_22415_, _22416_, _22423_);
  or g_53631_(_22422_, _22423_, _22424_);
  or g_53632_(_22421_, _22424_, _22425_);
  xor g_53633_(out[108], out[412], _22426_);
  or g_53634_(_22401_, _22426_, _22427_);
  or g_53635_(_22400_, _22412_, _22429_);
  or g_53636_(_22427_, _22429_, _22430_);
  or g_53637_(_22404_, _22410_, _22431_);
  or g_53638_(_22413_, _22431_, _22432_);
  or g_53639_(_22430_, _22432_, _22433_);
  or g_53640_(_22425_, _22433_, _22434_);
  or g_53641_(_22418_, _22434_, _22435_);
  and g_53642_(out[91], _39779_, _22436_);
  and g_53643_(_39559_, out[411], _22437_);
  xor g_53644_(out[88], out[408], _22438_);
  xor g_53645_(out[95], out[415], _22440_);
  xor g_53646_(out[81], out[401], _22441_);
  xor g_53647_(out[82], out[402], _22442_);
  xor g_53648_(out[84], out[404], _22443_);
  xor g_53649_(out[85], out[405], _22444_);
  xor g_53650_(out[89], out[409], _22445_);
  xor g_53651_(out[83], out[403], _22446_);
  xor g_53652_(out[94], out[414], _22447_);
  xor g_53653_(out[80], out[400], _22448_);
  xor g_53654_(out[90], out[410], _22449_);
  xor g_53655_(out[93], out[413], _22451_);
  or g_53656_(_22438_, _22451_, _22452_);
  xor g_53657_(out[86], out[406], _22453_);
  or g_53658_(_22442_, _22449_, _22454_);
  or g_53659_(_22452_, _22454_, _22455_);
  or g_53660_(_22445_, _22446_, _22456_);
  or g_53661_(_22444_, _22456_, _22457_);
  or g_53662_(_22455_, _22457_, _22458_);
  or g_53663_(_22443_, _22447_, _22459_);
  or g_53664_(_22458_, _22459_, _22460_);
  xor g_53665_(out[92], out[412], _22462_);
  or g_53666_(_22437_, _22462_, _22463_);
  xor g_53667_(out[87], out[407], _22464_);
  or g_53668_(_22453_, _22464_, _22465_);
  or g_53669_(_22463_, _22465_, _22466_);
  or g_53670_(_22436_, _22441_, _22467_);
  or g_53671_(_22440_, _22467_, _22468_);
  or g_53672_(_22466_, _22468_, _22469_);
  or g_53673_(_22448_, _22469_, _22470_);
  or g_53674_(_22460_, _22470_, _22471_);
  xor g_53675_(out[71], out[407], _22473_);
  and g_53676_(_39548_, out[411], _22474_);
  xor g_53677_(out[78], out[414], _22475_);
  xor g_53678_(out[72], out[408], _22476_);
  xor g_53679_(out[65], out[401], _22477_);
  xor g_53680_(out[77], out[413], _22478_);
  xor g_53681_(out[73], out[409], _22479_);
  xor g_53682_(out[68], out[404], _22480_);
  xor g_53683_(out[66], out[402], _22481_);
  and g_53684_(out[75], _39779_, _22482_);
  xor g_53685_(out[67], out[403], _22484_);
  xor g_53686_(out[70], out[406], _22485_);
  xor g_53687_(out[79], out[415], _22486_);
  xor g_53688_(out[74], out[410], _22487_);
  xor g_53689_(out[69], out[405], _22488_);
  xor g_53690_(out[64], out[400], _22489_);
  or g_53691_(_22475_, _22480_, _22490_);
  or g_53692_(_22476_, _22478_, _22491_);
  or g_53693_(_22481_, _22487_, _22492_);
  or g_53694_(_22491_, _22492_, _22493_);
  or g_53695_(_22479_, _22484_, _22495_);
  or g_53696_(_22488_, _22489_, _22496_);
  or g_53697_(_22495_, _22496_, _22497_);
  or g_53698_(_22493_, _22497_, _22498_);
  xor g_53699_(out[76], out[412], _22499_);
  or g_53700_(_22474_, _22499_, _22500_);
  or g_53701_(_22473_, _22485_, _22501_);
  or g_53702_(_22500_, _22501_, _22502_);
  or g_53703_(_22477_, _22482_, _22503_);
  or g_53704_(_22486_, _22503_, _22504_);
  or g_53705_(_22502_, _22504_, _22506_);
  or g_53706_(_22498_, _22506_, _22507_);
  or g_53707_(_22490_, _22507_, _22508_);
  xor g_53708_(out[49], out[401], _22509_);
  and g_53709_(out[59], _39779_, _22510_);
  xor g_53710_(out[57], out[409], _22511_);
  xor g_53711_(out[48], out[400], _22512_);
  xor g_53712_(out[62], out[414], _22513_);
  xor g_53713_(out[52], out[404], _22514_);
  or g_53714_(_22513_, _22514_, _22515_);
  xor g_53715_(out[61], out[413], _22517_);
  xor g_53716_(out[51], out[403], _22518_);
  and g_53717_(_39537_, out[411], _22519_);
  xor g_53718_(out[54], out[406], _22520_);
  xor g_53719_(out[58], out[410], _22521_);
  xor g_53720_(out[53], out[405], _22522_);
  xor g_53721_(out[63], out[415], _22523_);
  xor g_53722_(out[56], out[408], _22524_);
  or g_53723_(_22517_, _22524_, _22525_);
  xor g_53724_(out[50], out[402], _22526_);
  or g_53725_(_22521_, _22526_, _22528_);
  or g_53726_(_22525_, _22528_, _22529_);
  or g_53727_(_22511_, _22518_, _22530_);
  or g_53728_(_22522_, _22530_, _22531_);
  or g_53729_(_22529_, _22531_, _22532_);
  or g_53730_(_22515_, _22532_, _22533_);
  xor g_53731_(out[60], out[412], _22534_);
  or g_53732_(_22519_, _22534_, _22535_);
  xor g_53733_(out[55], out[407], _22536_);
  or g_53734_(_22520_, _22536_, _22537_);
  or g_53735_(_22535_, _22537_, _22539_);
  or g_53736_(_22509_, _22510_, _22540_);
  or g_53737_(_22523_, _22540_, _22541_);
  or g_53738_(_22539_, _22541_, _22542_);
  or g_53739_(_22512_, _22542_, _22543_);
  or g_53740_(_22533_, _22543_, _22544_);
  xor g_53741_(out[39], out[407], _22545_);
  and g_53742_(_39526_, out[411], _22546_);
  xor g_53743_(out[46], out[414], _22547_);
  xor g_53744_(out[40], out[408], _22548_);
  xor g_53745_(out[33], out[401], _22550_);
  xor g_53746_(out[45], out[413], _22551_);
  xor g_53747_(out[41], out[409], _22552_);
  xor g_53748_(out[36], out[404], _22553_);
  xor g_53749_(out[34], out[402], _22554_);
  and g_53750_(out[43], _39779_, _22555_);
  xor g_53751_(out[35], out[403], _22556_);
  xor g_53752_(out[38], out[406], _22557_);
  xor g_53753_(out[47], out[415], _22558_);
  xor g_53754_(out[42], out[410], _22559_);
  xor g_53755_(out[37], out[405], _22561_);
  xor g_53756_(out[32], out[400], _22562_);
  or g_53757_(_22547_, _22553_, _22563_);
  or g_53758_(_22548_, _22551_, _22564_);
  or g_53759_(_22554_, _22559_, _22565_);
  or g_53760_(_22564_, _22565_, _22566_);
  or g_53761_(_22552_, _22556_, _22567_);
  or g_53762_(_22561_, _22562_, _22568_);
  or g_53763_(_22567_, _22568_, _22569_);
  or g_53764_(_22566_, _22569_, _22570_);
  xor g_53765_(out[44], out[412], _22572_);
  or g_53766_(_22546_, _22572_, _22573_);
  or g_53767_(_22545_, _22557_, _22574_);
  or g_53768_(_22573_, _22574_, _22575_);
  or g_53769_(_22550_, _22555_, _22576_);
  or g_53770_(_22558_, _22576_, _22577_);
  or g_53771_(_22575_, _22577_, _22578_);
  or g_53772_(_22570_, _22578_, _22579_);
  or g_53773_(_22563_, _22579_, _22580_);
  xor g_53774_(out[24], out[408], _22581_);
  xor g_53775_(out[21], out[405], _22583_);
  xor g_53776_(out[19], out[403], _22584_);
  xor g_53777_(out[30], out[414], _22585_);
  xor g_53778_(out[29], out[413], _22586_);
  xor g_53779_(out[18], out[402], _22587_);
  xor g_53780_(out[25], out[409], _22588_);
  xor g_53781_(out[22], out[406], _22589_);
  xor g_53782_(out[31], out[415], _22590_);
  xor g_53783_(out[26], out[410], _22591_);
  xor g_53784_(out[20], out[404], _22592_);
  xor g_53785_(out[16], out[400], _22594_);
  and g_53786_(_39493_, out[411], _22595_);
  and g_53787_(out[27], _39779_, _22596_);
  or g_53788_(_22581_, _22586_, _22597_);
  xor g_53789_(out[17], out[401], _22598_);
  or g_53790_(_22587_, _22591_, _22599_);
  or g_53791_(_22597_, _22599_, _22600_);
  or g_53792_(_22584_, _22588_, _22601_);
  or g_53793_(_22583_, _22601_, _22602_);
  or g_53794_(_22600_, _22602_, _22603_);
  or g_53795_(_22585_, _22592_, _22605_);
  or g_53796_(_22603_, _22605_, _22606_);
  xor g_53797_(out[28], out[412], _22607_);
  or g_53798_(_22595_, _22607_, _22608_);
  xor g_53799_(out[23], out[407], _22609_);
  or g_53800_(_22589_, _22609_, _22610_);
  or g_53801_(_22608_, _22610_, _22611_);
  or g_53802_(_22596_, _22598_, _22612_);
  or g_53803_(_22590_, _22612_, _22613_);
  or g_53804_(_22611_, _22613_, _22614_);
  or g_53805_(_22594_, _22614_, _22616_);
  or g_53806_(_22606_, _22616_, _22617_);
  not g_53807_(_22617_, _22618_);
  xor g_53808_(out[1], out[401], _22619_);
  and g_53809_(_39438_, out[411], _22620_);
  and g_53810_(out[11], _39779_, _22621_);
  xor g_53811_(out[14], out[414], _22622_);
  xor g_53812_(out[3], out[403], _22623_);
  xor g_53813_(out[4], out[404], _22624_);
  xor g_53814_(out[2], out[402], _22625_);
  xor g_53815_(out[9], out[409], _22627_);
  xor g_53816_(out[0], out[400], _22628_);
  xor g_53817_(out[12], out[412], _22629_);
  xor g_53818_(out[6], out[406], _22630_);
  xor g_53819_(out[10], out[410], _22631_);
  xor g_53820_(out[5], out[405], _22632_);
  xor g_53821_(out[15], out[415], _22633_);
  xor g_53822_(out[13], out[413], _22634_);
  xor g_53823_(out[8], out[408], _22635_);
  or g_53824_(_22622_, _22624_, _22636_);
  or g_53825_(_22634_, _22635_, _22638_);
  or g_53826_(_22625_, _22631_, _22639_);
  or g_53827_(_22638_, _22639_, _22640_);
  or g_53828_(_22623_, _22627_, _22641_);
  or g_53829_(_22628_, _22632_, _22642_);
  or g_53830_(_22641_, _22642_, _22643_);
  or g_53831_(_22640_, _22643_, _22644_);
  or g_53832_(_22620_, _22629_, _22645_);
  xor g_53833_(out[7], out[407], _22646_);
  or g_53834_(_22630_, _22646_, _22647_);
  or g_53835_(_22645_, _22647_, _22649_);
  or g_53836_(_22619_, _22621_, _22650_);
  or g_53837_(_22633_, _22650_, _22651_);
  or g_53838_(_22649_, _22651_, _22652_);
  or g_53839_(_22644_, _22652_, _22653_);
  or g_53840_(_22636_, _22653_, _22654_);
  xor g_53841_(out[311], out[391], _22655_);
  and g_53842_(_39724_, out[395], _22656_);
  xor g_53843_(out[318], out[398], _22657_);
  xor g_53844_(out[312], out[392], _22658_);
  xor g_53845_(out[305], out[385], _22660_);
  xor g_53846_(out[317], out[397], _22661_);
  xor g_53847_(out[313], out[393], _22662_);
  xor g_53848_(out[308], out[388], _22663_);
  xor g_53849_(out[306], out[386], _22664_);
  and g_53850_(out[315], _39768_, _22665_);
  xor g_53851_(out[307], out[387], _22666_);
  xor g_53852_(out[310], out[390], _22667_);
  xor g_53853_(out[319], out[399], _22668_);
  xor g_53854_(out[314], out[394], _22669_);
  xor g_53855_(out[309], out[389], _22671_);
  xor g_53856_(out[304], out[384], _22672_);
  or g_53857_(_22657_, _22663_, _22673_);
  or g_53858_(_22658_, _22661_, _22674_);
  or g_53859_(_22664_, _22669_, _22675_);
  or g_53860_(_22674_, _22675_, _22676_);
  or g_53861_(_22662_, _22666_, _22677_);
  or g_53862_(_22671_, _22672_, _22678_);
  or g_53863_(_22677_, _22678_, _22679_);
  or g_53864_(_22676_, _22679_, _22680_);
  xor g_53865_(out[316], out[396], _22682_);
  or g_53866_(_22656_, _22682_, _22683_);
  or g_53867_(_22655_, _22667_, _22684_);
  or g_53868_(_22683_, _22684_, _22685_);
  or g_53869_(_22660_, _22665_, _22686_);
  or g_53870_(_22668_, _22686_, _22687_);
  or g_53871_(_22685_, _22687_, _22688_);
  or g_53872_(_22680_, _22688_, _22689_);
  or g_53873_(_22673_, _22689_, _22690_);
  xor g_53874_(out[296], out[392], _22691_);
  xor g_53875_(out[293], out[389], _22693_);
  xor g_53876_(out[291], out[387], _22694_);
  xor g_53877_(out[302], out[398], _22695_);
  xor g_53878_(out[301], out[397], _22696_);
  xor g_53879_(out[290], out[386], _22697_);
  xor g_53880_(out[297], out[393], _22698_);
  xor g_53881_(out[294], out[390], _22699_);
  xor g_53882_(out[303], out[399], _22700_);
  xor g_53883_(out[298], out[394], _22701_);
  xor g_53884_(out[292], out[388], _22702_);
  xor g_53885_(out[288], out[384], _22704_);
  and g_53886_(_39702_, out[395], _22705_);
  and g_53887_(out[299], _39768_, _22706_);
  or g_53888_(_22691_, _22696_, _22707_);
  xor g_53889_(out[289], out[385], _22708_);
  or g_53890_(_22697_, _22701_, _22709_);
  or g_53891_(_22707_, _22709_, _22710_);
  or g_53892_(_22694_, _22698_, _22711_);
  or g_53893_(_22693_, _22711_, _22712_);
  or g_53894_(_22710_, _22712_, _22713_);
  or g_53895_(_22695_, _22702_, _22715_);
  or g_53896_(_22713_, _22715_, _22716_);
  xor g_53897_(out[300], out[396], _22717_);
  or g_53898_(_22705_, _22717_, _22718_);
  xor g_53899_(out[295], out[391], _22719_);
  or g_53900_(_22699_, _22719_, _22720_);
  or g_53901_(_22718_, _22720_, _22721_);
  or g_53902_(_22706_, _22708_, _22722_);
  or g_53903_(_22700_, _22722_, _22723_);
  or g_53904_(_22721_, _22723_, _22724_);
  or g_53905_(_22704_, _22724_, _22726_);
  or g_53906_(_22716_, _22726_, _22727_);
  xor g_53907_(out[279], out[391], _22728_);
  and g_53908_(_39691_, out[395], _22729_);
  xor g_53909_(out[286], out[398], _22730_);
  xor g_53910_(out[280], out[392], _22731_);
  xor g_53911_(out[273], out[385], _22732_);
  xor g_53912_(out[285], out[397], _22733_);
  xor g_53913_(out[281], out[393], _22734_);
  xor g_53914_(out[276], out[388], _22735_);
  xor g_53915_(out[274], out[386], _22737_);
  and g_53916_(out[283], _39768_, _22738_);
  xor g_53917_(out[275], out[387], _22739_);
  xor g_53918_(out[278], out[390], _22740_);
  xor g_53919_(out[287], out[399], _22741_);
  xor g_53920_(out[282], out[394], _22742_);
  xor g_53921_(out[277], out[389], _22743_);
  xor g_53922_(out[272], out[384], _22744_);
  or g_53923_(_22730_, _22735_, _22745_);
  or g_53924_(_22731_, _22733_, _22746_);
  or g_53925_(_22737_, _22742_, _22748_);
  or g_53926_(_22746_, _22748_, _22749_);
  or g_53927_(_22734_, _22739_, _22750_);
  or g_53928_(_22743_, _22744_, _22751_);
  or g_53929_(_22750_, _22751_, _22752_);
  or g_53930_(_22749_, _22752_, _22753_);
  xor g_53931_(out[284], out[396], _22754_);
  or g_53932_(_22729_, _22754_, _22755_);
  or g_53933_(_22728_, _22740_, _22756_);
  or g_53934_(_22755_, _22756_, _22757_);
  or g_53935_(_22732_, _22738_, _22759_);
  or g_53936_(_22741_, _22759_, _22760_);
  or g_53937_(_22757_, _22760_, _22761_);
  or g_53938_(_22753_, _22761_, _22762_);
  or g_53939_(_22745_, _22762_, _22763_);
  xor g_53940_(out[268], out[396], _22764_);
  and g_53941_(_39680_, out[395], _22765_);
  xor g_53942_(out[264], out[392], _22766_);
  xor g_53943_(out[262], out[390], _22767_);
  xor g_53944_(out[269], out[397], _22768_);
  xor g_53945_(out[270], out[398], _22770_);
  xor g_53946_(out[258], out[386], _22771_);
  xor g_53947_(out[265], out[393], _22772_);
  xor g_53948_(out[261], out[389], _22773_);
  xor g_53949_(out[257], out[385], _22774_);
  and g_53950_(out[267], _39768_, _22775_);
  or g_53951_(_22766_, _22768_, _22776_);
  xor g_53952_(out[271], out[399], _22777_);
  xor g_53953_(out[266], out[394], _22778_);
  xor g_53954_(out[260], out[388], _22779_);
  xor g_53955_(out[259], out[387], _22781_);
  xor g_53956_(out[256], out[384], _22782_);
  or g_53957_(_22771_, _22778_, _22783_);
  or g_53958_(_22776_, _22783_, _22784_);
  or g_53959_(_22772_, _22781_, _22785_);
  or g_53960_(_22773_, _22785_, _22786_);
  or g_53961_(_22784_, _22786_, _22787_);
  or g_53962_(_22770_, _22779_, _22788_);
  or g_53963_(_22787_, _22788_, _22789_);
  or g_53964_(_22764_, _22765_, _22790_);
  xor g_53965_(out[263], out[391], _22792_);
  or g_53966_(_22767_, _22792_, _22793_);
  or g_53967_(_22790_, _22793_, _22794_);
  or g_53968_(_22774_, _22775_, _22795_);
  or g_53969_(_22777_, _22795_, _22796_);
  or g_53970_(_22794_, _22796_, _22797_);
  or g_53971_(_22782_, _22797_, _22798_);
  or g_53972_(_22789_, _22798_, _22799_);
  xor g_53973_(out[247], out[391], _22800_);
  and g_53974_(_39669_, out[395], _22801_);
  xor g_53975_(out[254], out[398], _22803_);
  xor g_53976_(out[248], out[392], _22804_);
  xor g_53977_(out[241], out[385], _22805_);
  xor g_53978_(out[253], out[397], _22806_);
  xor g_53979_(out[249], out[393], _22807_);
  xor g_53980_(out[244], out[388], _22808_);
  xor g_53981_(out[242], out[386], _22809_);
  and g_53982_(out[251], _39768_, _22810_);
  xor g_53983_(out[243], out[387], _22811_);
  xor g_53984_(out[246], out[390], _22812_);
  xor g_53985_(out[255], out[399], _22814_);
  xor g_53986_(out[250], out[394], _22815_);
  xor g_53987_(out[245], out[389], _22816_);
  xor g_53988_(out[240], out[384], _22817_);
  or g_53989_(_22803_, _22808_, _22818_);
  or g_53990_(_22804_, _22806_, _22819_);
  or g_53991_(_22809_, _22815_, _22820_);
  or g_53992_(_22819_, _22820_, _22821_);
  or g_53993_(_22807_, _22811_, _22822_);
  or g_53994_(_22816_, _22817_, _22823_);
  or g_53995_(_22822_, _22823_, _22825_);
  or g_53996_(_22821_, _22825_, _22826_);
  xor g_53997_(out[252], out[396], _22827_);
  or g_53998_(_22801_, _22827_, _22828_);
  or g_53999_(_22800_, _22812_, _22829_);
  or g_54000_(_22828_, _22829_, _22830_);
  or g_54001_(_22805_, _22810_, _22831_);
  or g_54002_(_22814_, _22831_, _22832_);
  or g_54003_(_22830_, _22832_, _22833_);
  or g_54004_(_22826_, _22833_, _22834_);
  or g_54005_(_22818_, _22834_, _22836_);
  not g_54006_(_22836_, _22837_);
  xor g_54007_(out[232], out[392], _22838_);
  xor g_54008_(out[229], out[389], _22839_);
  xor g_54009_(out[227], out[387], _22840_);
  xor g_54010_(out[238], out[398], _22841_);
  xor g_54011_(out[237], out[397], _22842_);
  xor g_54012_(out[226], out[386], _22843_);
  xor g_54013_(out[233], out[393], _22844_);
  xor g_54014_(out[230], out[390], _22845_);
  xor g_54015_(out[239], out[399], _22847_);
  xor g_54016_(out[234], out[394], _22848_);
  xor g_54017_(out[228], out[388], _22849_);
  xor g_54018_(out[224], out[384], _22850_);
  and g_54019_(_39658_, out[395], _22851_);
  and g_54020_(out[235], _39768_, _22852_);
  or g_54021_(_22838_, _22842_, _22853_);
  xor g_54022_(out[225], out[385], _22854_);
  or g_54023_(_22843_, _22848_, _22855_);
  or g_54024_(_22853_, _22855_, _22856_);
  or g_54025_(_22840_, _22844_, _22858_);
  or g_54026_(_22839_, _22858_, _22859_);
  or g_54027_(_22856_, _22859_, _22860_);
  or g_54028_(_22841_, _22849_, _22861_);
  or g_54029_(_22860_, _22861_, _22862_);
  xor g_54030_(out[236], out[396], _22863_);
  or g_54031_(_22851_, _22863_, _22864_);
  xor g_54032_(out[231], out[391], _22865_);
  or g_54033_(_22845_, _22865_, _22866_);
  or g_54034_(_22864_, _22866_, _22867_);
  or g_54035_(_22852_, _22854_, _22869_);
  or g_54036_(_22847_, _22869_, _22870_);
  or g_54037_(_22867_, _22870_, _22871_);
  or g_54038_(_22850_, _22871_, _22872_);
  or g_54039_(_22862_, _22872_, _22873_);
  xor g_54040_(out[215], out[391], _22874_);
  and g_54041_(_39647_, out[395], _22875_);
  xor g_54042_(out[222], out[398], _22876_);
  xor g_54043_(out[216], out[392], _22877_);
  xor g_54044_(out[209], out[385], _22878_);
  xor g_54045_(out[221], out[397], _22880_);
  xor g_54046_(out[217], out[393], _22881_);
  xor g_54047_(out[212], out[388], _22882_);
  xor g_54048_(out[210], out[386], _22883_);
  and g_54049_(out[219], _39768_, _22884_);
  xor g_54050_(out[211], out[387], _22885_);
  xor g_54051_(out[214], out[390], _22886_);
  xor g_54052_(out[223], out[399], _22887_);
  xor g_54053_(out[218], out[394], _22888_);
  xor g_54054_(out[213], out[389], _22889_);
  xor g_54055_(out[208], out[384], _22891_);
  or g_54056_(_22876_, _22882_, _22892_);
  or g_54057_(_22877_, _22880_, _22893_);
  or g_54058_(_22883_, _22888_, _22894_);
  or g_54059_(_22893_, _22894_, _22895_);
  or g_54060_(_22881_, _22885_, _22896_);
  or g_54061_(_22889_, _22891_, _22897_);
  or g_54062_(_22896_, _22897_, _22898_);
  or g_54063_(_22895_, _22898_, _22899_);
  xor g_54064_(out[220], out[396], _22900_);
  or g_54065_(_22875_, _22900_, _22902_);
  or g_54066_(_22874_, _22886_, _22903_);
  or g_54067_(_22902_, _22903_, _22904_);
  or g_54068_(_22878_, _22884_, _22905_);
  or g_54069_(_22887_, _22905_, _22906_);
  or g_54070_(_22904_, _22906_, _22907_);
  or g_54071_(_22899_, _22907_, _22908_);
  or g_54072_(_22892_, _22908_, _22909_);
  xor g_54073_(out[193], out[385], _22910_);
  and g_54074_(_39636_, out[395], _22911_);
  and g_54075_(out[203], _39768_, _22913_);
  xor g_54076_(out[201], out[393], _22914_);
  xor g_54077_(out[192], out[384], _22915_);
  xor g_54078_(out[206], out[398], _22916_);
  xor g_54079_(out[196], out[388], _22917_);
  or g_54080_(_22916_, _22917_, _22918_);
  xor g_54081_(out[205], out[397], _22919_);
  xor g_54082_(out[195], out[387], _22920_);
  xor g_54083_(out[204], out[396], _22921_);
  xor g_54084_(out[198], out[390], _22922_);
  xor g_54085_(out[202], out[394], _22924_);
  xor g_54086_(out[197], out[389], _22925_);
  xor g_54087_(out[207], out[399], _22926_);
  xor g_54088_(out[200], out[392], _22927_);
  or g_54089_(_22919_, _22927_, _22928_);
  xor g_54090_(out[194], out[386], _22929_);
  or g_54091_(_22924_, _22929_, _22930_);
  or g_54092_(_22928_, _22930_, _22931_);
  or g_54093_(_22914_, _22920_, _22932_);
  or g_54094_(_22925_, _22932_, _22933_);
  or g_54095_(_22931_, _22933_, _22935_);
  or g_54096_(_22918_, _22935_, _22936_);
  or g_54097_(_22911_, _22921_, _22937_);
  xor g_54098_(out[199], out[391], _22938_);
  or g_54099_(_22922_, _22938_, _22939_);
  or g_54100_(_22937_, _22939_, _22940_);
  or g_54101_(_22910_, _22913_, _22941_);
  or g_54102_(_22926_, _22941_, _22942_);
  or g_54103_(_22940_, _22942_, _22943_);
  or g_54104_(_22915_, _22943_, _22944_);
  or g_54105_(_22936_, _22944_, _22946_);
  xor g_54106_(out[183], out[391], _22947_);
  and g_54107_(_39625_, out[395], _22948_);
  xor g_54108_(out[190], out[398], _22949_);
  xor g_54109_(out[184], out[392], _22950_);
  xor g_54110_(out[177], out[385], _22951_);
  xor g_54111_(out[189], out[397], _22952_);
  xor g_54112_(out[185], out[393], _22953_);
  xor g_54113_(out[180], out[388], _22954_);
  xor g_54114_(out[178], out[386], _22955_);
  and g_54115_(out[187], _39768_, _22957_);
  xor g_54116_(out[179], out[387], _22958_);
  xor g_54117_(out[182], out[390], _22959_);
  xor g_54118_(out[191], out[399], _22960_);
  xor g_54119_(out[186], out[394], _22961_);
  xor g_54120_(out[181], out[389], _22962_);
  xor g_54121_(out[176], out[384], _22963_);
  or g_54122_(_22949_, _22954_, _22964_);
  or g_54123_(_22950_, _22952_, _22965_);
  or g_54124_(_22955_, _22961_, _22966_);
  or g_54125_(_22965_, _22966_, _22968_);
  or g_54126_(_22953_, _22958_, _22969_);
  or g_54127_(_22962_, _22963_, _22970_);
  or g_54128_(_22969_, _22970_, _22971_);
  or g_54129_(_22968_, _22971_, _22972_);
  xor g_54130_(out[188], out[396], _22973_);
  or g_54131_(_22948_, _22973_, _22974_);
  or g_54132_(_22947_, _22959_, _22975_);
  or g_54133_(_22974_, _22975_, _22976_);
  or g_54134_(_22951_, _22957_, _22977_);
  or g_54135_(_22960_, _22977_, _22979_);
  or g_54136_(_22976_, _22979_, _22980_);
  or g_54137_(_22972_, _22980_, _22981_);
  or g_54138_(_22964_, _22981_, _22982_);
  not g_54139_(_22982_, _22983_);
  xor g_54140_(out[161], out[385], _22984_);
  and g_54141_(out[171], _39768_, _22985_);
  xor g_54142_(out[169], out[393], _22986_);
  xor g_54143_(out[160], out[384], _22987_);
  xor g_54144_(out[174], out[398], _22988_);
  xor g_54145_(out[164], out[388], _22990_);
  or g_54146_(_22988_, _22990_, _22991_);
  xor g_54147_(out[173], out[397], _22992_);
  xor g_54148_(out[163], out[387], _22993_);
  and g_54149_(_39614_, out[395], _22994_);
  xor g_54150_(out[166], out[390], _22995_);
  xor g_54151_(out[170], out[394], _22996_);
  xor g_54152_(out[165], out[389], _22997_);
  xor g_54153_(out[175], out[399], _22998_);
  xor g_54154_(out[168], out[392], _22999_);
  or g_54155_(_22992_, _22999_, _23001_);
  xor g_54156_(out[162], out[386], _23002_);
  or g_54157_(_22996_, _23002_, _23003_);
  or g_54158_(_23001_, _23003_, _23004_);
  or g_54159_(_22986_, _22993_, _23005_);
  or g_54160_(_22997_, _23005_, _23006_);
  or g_54161_(_23004_, _23006_, _23007_);
  or g_54162_(_22991_, _23007_, _23008_);
  xor g_54163_(out[172], out[396], _23009_);
  or g_54164_(_22994_, _23009_, _23010_);
  xor g_54165_(out[167], out[391], _23012_);
  or g_54166_(_22995_, _23012_, _23013_);
  or g_54167_(_23010_, _23013_, _23014_);
  or g_54168_(_22984_, _22985_, _23015_);
  or g_54169_(_22998_, _23015_, _23016_);
  or g_54170_(_23014_, _23016_, _23017_);
  or g_54171_(_22987_, _23017_, _23018_);
  or g_54172_(_23008_, _23018_, _23019_);
  xor g_54173_(out[151], out[391], _23020_);
  and g_54174_(_39603_, out[395], _23021_);
  xor g_54175_(out[158], out[398], _23023_);
  xor g_54176_(out[152], out[392], _23024_);
  xor g_54177_(out[145], out[385], _23025_);
  xor g_54178_(out[157], out[397], _23026_);
  xor g_54179_(out[153], out[393], _23027_);
  xor g_54180_(out[148], out[388], _23028_);
  xor g_54181_(out[146], out[386], _23029_);
  and g_54182_(out[155], _39768_, _23030_);
  xor g_54183_(out[147], out[387], _23031_);
  xor g_54184_(out[150], out[390], _23032_);
  xor g_54185_(out[159], out[399], _23034_);
  xor g_54186_(out[154], out[394], _23035_);
  xor g_54187_(out[149], out[389], _23036_);
  xor g_54188_(out[144], out[384], _23037_);
  or g_54189_(_23023_, _23028_, _23038_);
  or g_54190_(_23024_, _23026_, _23039_);
  or g_54191_(_23029_, _23035_, _23040_);
  or g_54192_(_23039_, _23040_, _23041_);
  or g_54193_(_23027_, _23031_, _23042_);
  or g_54194_(_23036_, _23037_, _23043_);
  or g_54195_(_23042_, _23043_, _23045_);
  or g_54196_(_23041_, _23045_, _23046_);
  xor g_54197_(out[156], out[396], _23047_);
  or g_54198_(_23021_, _23047_, _23048_);
  or g_54199_(_23020_, _23032_, _23049_);
  or g_54200_(_23048_, _23049_, _23050_);
  or g_54201_(_23025_, _23030_, _23051_);
  or g_54202_(_23034_, _23051_, _23052_);
  or g_54203_(_23050_, _23052_, _23053_);
  or g_54204_(_23046_, _23053_, _23054_);
  or g_54205_(_23038_, _23054_, _23056_);
  and g_54206_(out[139], _39768_, _23057_);
  xor g_54207_(out[132], out[388], _23058_);
  xor g_54208_(out[142], out[398], _23059_);
  or g_54209_(_23058_, _23059_, _23060_);
  xor g_54210_(out[141], out[397], _23061_);
  xor g_54211_(out[131], out[387], _23062_);
  xor g_54212_(out[128], out[384], _23063_);
  and g_54213_(_39592_, out[395], _23064_);
  xor g_54214_(out[138], out[394], _23065_);
  xor g_54215_(out[143], out[399], _23067_);
  xor g_54216_(out[134], out[390], _23068_);
  xor g_54217_(out[133], out[389], _23069_);
  xor g_54218_(out[136], out[392], _23070_);
  or g_54219_(_23061_, _23070_, _23071_);
  xor g_54220_(out[130], out[386], _23072_);
  xor g_54221_(out[137], out[393], _23073_);
  xor g_54222_(out[129], out[385], _23074_);
  or g_54223_(_23065_, _23072_, _23075_);
  or g_54224_(_23071_, _23075_, _23076_);
  or g_54225_(_23062_, _23073_, _23078_);
  or g_54226_(_23069_, _23078_, _23079_);
  or g_54227_(_23076_, _23079_, _23080_);
  or g_54228_(_23060_, _23080_, _23081_);
  xor g_54229_(out[140], out[396], _23082_);
  or g_54230_(_23064_, _23082_, _23083_);
  xor g_54231_(out[135], out[391], _23084_);
  or g_54232_(_23068_, _23084_, _23085_);
  or g_54233_(_23083_, _23085_, _23086_);
  or g_54234_(_23057_, _23074_, _23087_);
  or g_54235_(_23067_, _23087_, _23089_);
  or g_54236_(_23086_, _23089_, _23090_);
  or g_54237_(_23063_, _23090_, _23091_);
  or g_54238_(_23081_, _23091_, _23092_);
  xor g_54239_(out[119], out[391], _23093_);
  and g_54240_(_39581_, out[395], _23094_);
  xor g_54241_(out[126], out[398], _23095_);
  xor g_54242_(out[120], out[392], _23096_);
  xor g_54243_(out[113], out[385], _23097_);
  xor g_54244_(out[125], out[397], _23098_);
  xor g_54245_(out[121], out[393], _23100_);
  xor g_54246_(out[116], out[388], _23101_);
  xor g_54247_(out[114], out[386], _23102_);
  and g_54248_(out[123], _39768_, _23103_);
  xor g_54249_(out[115], out[387], _23104_);
  xor g_54250_(out[118], out[390], _23105_);
  xor g_54251_(out[127], out[399], _23106_);
  xor g_54252_(out[122], out[394], _23107_);
  xor g_54253_(out[117], out[389], _23108_);
  xor g_54254_(out[112], out[384], _23109_);
  or g_54255_(_23095_, _23101_, _23111_);
  or g_54256_(_23096_, _23098_, _23112_);
  or g_54257_(_23102_, _23107_, _23113_);
  or g_54258_(_23112_, _23113_, _23114_);
  or g_54259_(_23100_, _23104_, _23115_);
  or g_54260_(_23108_, _23109_, _23116_);
  or g_54261_(_23115_, _23116_, _23117_);
  or g_54262_(_23114_, _23117_, _23118_);
  xor g_54263_(out[124], out[396], _23119_);
  or g_54264_(_23094_, _23119_, _23120_);
  or g_54265_(_23093_, _23105_, _23122_);
  or g_54266_(_23120_, _23122_, _23123_);
  or g_54267_(_23097_, _23103_, _23124_);
  or g_54268_(_23106_, _23124_, _23125_);
  or g_54269_(_23123_, _23125_, _23126_);
  or g_54270_(_23118_, _23126_, _23127_);
  or g_54271_(_23111_, _23127_, _23128_);
  xor g_54272_(out[97], out[385], _23129_);
  and g_54273_(out[107], _39768_, _23130_);
  xor g_54274_(out[105], out[393], _23131_);
  xor g_54275_(out[96], out[384], _23133_);
  xor g_54276_(out[110], out[398], _23134_);
  xor g_54277_(out[100], out[388], _23135_);
  or g_54278_(_23134_, _23135_, _23136_);
  xor g_54279_(out[109], out[397], _23137_);
  xor g_54280_(out[99], out[387], _23138_);
  and g_54281_(_39570_, out[395], _23139_);
  xor g_54282_(out[102], out[390], _23140_);
  xor g_54283_(out[106], out[394], _23141_);
  xor g_54284_(out[101], out[389], _23142_);
  xor g_54285_(out[111], out[399], _23144_);
  xor g_54286_(out[104], out[392], _23145_);
  or g_54287_(_23137_, _23145_, _23146_);
  xor g_54288_(out[98], out[386], _23147_);
  or g_54289_(_23141_, _23147_, _23148_);
  or g_54290_(_23146_, _23148_, _23149_);
  or g_54291_(_23131_, _23138_, _23150_);
  or g_54292_(_23142_, _23150_, _23151_);
  or g_54293_(_23149_, _23151_, _23152_);
  or g_54294_(_23136_, _23152_, _23153_);
  xor g_54295_(out[108], out[396], _23155_);
  or g_54296_(_23139_, _23155_, _23156_);
  xor g_54297_(out[103], out[391], _23157_);
  or g_54298_(_23140_, _23157_, _23158_);
  or g_54299_(_23156_, _23158_, _23159_);
  or g_54300_(_23129_, _23130_, _23160_);
  or g_54301_(_23144_, _23160_, _23161_);
  or g_54302_(_23159_, _23161_, _23162_);
  or g_54303_(_23133_, _23162_, _23163_);
  or g_54304_(_23153_, _23163_, _23164_);
  xor g_54305_(out[87], out[391], _23166_);
  and g_54306_(_39559_, out[395], _23167_);
  xor g_54307_(out[94], out[398], _23168_);
  xor g_54308_(out[88], out[392], _23169_);
  xor g_54309_(out[81], out[385], _23170_);
  xor g_54310_(out[93], out[397], _23171_);
  xor g_54311_(out[89], out[393], _23172_);
  xor g_54312_(out[84], out[388], _23173_);
  xor g_54313_(out[82], out[386], _23174_);
  and g_54314_(out[91], _39768_, _23175_);
  xor g_54315_(out[83], out[387], _23177_);
  xor g_54316_(out[86], out[390], _23178_);
  xor g_54317_(out[95], out[399], _23179_);
  xor g_54318_(out[90], out[394], _23180_);
  xor g_54319_(out[85], out[389], _23181_);
  xor g_54320_(out[80], out[384], _23182_);
  or g_54321_(_23168_, _23173_, _23183_);
  or g_54322_(_23169_, _23171_, _23184_);
  or g_54323_(_23174_, _23180_, _23185_);
  or g_54324_(_23184_, _23185_, _23186_);
  or g_54325_(_23172_, _23177_, _23188_);
  or g_54326_(_23181_, _23182_, _23189_);
  or g_54327_(_23188_, _23189_, _23190_);
  or g_54328_(_23186_, _23190_, _23191_);
  xor g_54329_(out[92], out[396], _23192_);
  or g_54330_(_23167_, _23192_, _23193_);
  or g_54331_(_23166_, _23178_, _23194_);
  or g_54332_(_23193_, _23194_, _23195_);
  or g_54333_(_23170_, _23175_, _23196_);
  or g_54334_(_23179_, _23196_, _23197_);
  or g_54335_(_23195_, _23197_, _23199_);
  or g_54336_(_23191_, _23199_, _23200_);
  or g_54337_(_23183_, _23200_, _23201_);
  xor g_54338_(out[74], out[394], _23202_);
  xor g_54339_(out[66], out[386], _23203_);
  xor g_54340_(out[65], out[385], _23204_);
  and g_54341_(_39548_, out[395], _23205_);
  and g_54342_(out[75], _39768_, _23206_);
  xor g_54343_(out[77], out[397], _23207_);
  xor g_54344_(out[67], out[387], _23208_);
  xor g_54345_(out[78], out[398], _23210_);
  xor g_54346_(out[76], out[396], _23211_);
  xor g_54347_(out[72], out[392], _23212_);
  xor g_54348_(out[79], out[399], _23213_);
  xor g_54349_(out[69], out[389], _23214_);
  xor g_54350_(out[70], out[390], _23215_);
  xor g_54351_(out[64], out[384], _23216_);
  xor g_54352_(out[68], out[388], _23217_);
  or g_54353_(_23207_, _23212_, _23218_);
  xor g_54354_(out[73], out[393], _23219_);
  or g_54355_(_23202_, _23203_, _23221_);
  or g_54356_(_23218_, _23221_, _23222_);
  or g_54357_(_23208_, _23219_, _23223_);
  or g_54358_(_23214_, _23223_, _23224_);
  or g_54359_(_23222_, _23224_, _23225_);
  or g_54360_(_23210_, _23217_, _23226_);
  or g_54361_(_23225_, _23226_, _23227_);
  or g_54362_(_23205_, _23211_, _23228_);
  xor g_54363_(out[71], out[391], _23229_);
  or g_54364_(_23215_, _23229_, _23230_);
  or g_54365_(_23228_, _23230_, _23232_);
  or g_54366_(_23204_, _23206_, _23233_);
  or g_54367_(_23213_, _23233_, _23234_);
  or g_54368_(_23232_, _23234_, _23235_);
  or g_54369_(_23216_, _23235_, _23236_);
  or g_54370_(_23227_, _23236_, _23237_);
  not g_54371_(_23237_, _23238_);
  xor g_54372_(out[55], out[391], _23239_);
  and g_54373_(_39537_, out[395], _23240_);
  xor g_54374_(out[62], out[398], _23241_);
  xor g_54375_(out[56], out[392], _23243_);
  xor g_54376_(out[49], out[385], _23244_);
  xor g_54377_(out[61], out[397], _23245_);
  xor g_54378_(out[57], out[393], _23246_);
  xor g_54379_(out[52], out[388], _23247_);
  xor g_54380_(out[50], out[386], _23248_);
  and g_54381_(out[59], _39768_, _23249_);
  xor g_54382_(out[51], out[387], _23250_);
  xor g_54383_(out[54], out[390], _23251_);
  xor g_54384_(out[63], out[399], _23252_);
  xor g_54385_(out[58], out[394], _23254_);
  xor g_54386_(out[53], out[389], _23255_);
  xor g_54387_(out[48], out[384], _23256_);
  or g_54388_(_23241_, _23247_, _23257_);
  or g_54389_(_23243_, _23245_, _23258_);
  or g_54390_(_23248_, _23254_, _23259_);
  or g_54391_(_23258_, _23259_, _23260_);
  or g_54392_(_23246_, _23250_, _23261_);
  or g_54393_(_23255_, _23256_, _23262_);
  or g_54394_(_23261_, _23262_, _23263_);
  or g_54395_(_23260_, _23263_, _23265_);
  xor g_54396_(out[60], out[396], _23266_);
  or g_54397_(_23240_, _23266_, _23267_);
  or g_54398_(_23239_, _23251_, _23268_);
  or g_54399_(_23267_, _23268_, _23269_);
  or g_54400_(_23244_, _23249_, _23270_);
  or g_54401_(_23252_, _23270_, _23271_);
  or g_54402_(_23269_, _23271_, _23272_);
  or g_54403_(_23265_, _23272_, _23273_);
  or g_54404_(_23257_, _23273_, _23274_);
  not g_54405_(_23274_, _23276_);
  xor g_54406_(out[32], out[384], _23277_);
  xor g_54407_(out[37], out[389], _23278_);
  xor g_54408_(out[47], out[399], _23279_);
  xor g_54409_(out[42], out[394], _23280_);
  xor g_54410_(out[35], out[387], _23281_);
  xor g_54411_(out[34], out[386], _23282_);
  and g_54412_(_39526_, out[395], _23283_);
  and g_54413_(out[43], _39768_, _23284_);
  xor g_54414_(out[36], out[388], _23285_);
  xor g_54415_(out[41], out[393], _23287_);
  xor g_54416_(out[40], out[392], _23288_);
  xor g_54417_(out[38], out[390], _23289_);
  xor g_54418_(out[33], out[385], _23290_);
  xor g_54419_(out[45], out[397], _23291_);
  xor g_54420_(out[46], out[398], _23292_);
  or g_54421_(_23285_, _23292_, _23293_);
  or g_54422_(_23288_, _23291_, _23294_);
  or g_54423_(_23280_, _23282_, _23295_);
  or g_54424_(_23294_, _23295_, _23296_);
  or g_54425_(_23281_, _23287_, _23298_);
  or g_54426_(_23277_, _23278_, _23299_);
  or g_54427_(_23298_, _23299_, _23300_);
  or g_54428_(_23296_, _23300_, _23301_);
  xor g_54429_(out[44], out[396], _23302_);
  or g_54430_(_23283_, _23302_, _23303_);
  xor g_54431_(out[39], out[391], _23304_);
  or g_54432_(_23289_, _23304_, _23305_);
  or g_54433_(_23303_, _23305_, _23306_);
  or g_54434_(_23284_, _23290_, _23307_);
  or g_54435_(_23279_, _23307_, _23309_);
  or g_54436_(_23306_, _23309_, _23310_);
  or g_54437_(_23301_, _23310_, _23311_);
  or g_54438_(_23293_, _23311_, _23312_);
  xor g_54439_(out[23], out[391], _23313_);
  and g_54440_(_39493_, out[395], _23314_);
  xor g_54441_(out[30], out[398], _23315_);
  xor g_54442_(out[24], out[392], _23316_);
  xor g_54443_(out[17], out[385], _23317_);
  xor g_54444_(out[29], out[397], _23318_);
  xor g_54445_(out[25], out[393], _23320_);
  xor g_54446_(out[20], out[388], _23321_);
  xor g_54447_(out[18], out[386], _23322_);
  and g_54448_(out[27], _39768_, _23323_);
  xor g_54449_(out[19], out[387], _23324_);
  xor g_54450_(out[22], out[390], _23325_);
  xor g_54451_(out[31], out[399], _23326_);
  xor g_54452_(out[26], out[394], _23327_);
  xor g_54453_(out[21], out[389], _23328_);
  xor g_54454_(out[16], out[384], _23329_);
  or g_54455_(_23315_, _23321_, _23331_);
  or g_54456_(_23316_, _23318_, _23332_);
  or g_54457_(_23322_, _23327_, _23333_);
  or g_54458_(_23332_, _23333_, _23334_);
  or g_54459_(_23320_, _23324_, _23335_);
  or g_54460_(_23328_, _23329_, _23336_);
  or g_54461_(_23335_, _23336_, _23337_);
  or g_54462_(_23334_, _23337_, _23338_);
  xor g_54463_(out[28], out[396], _23339_);
  or g_54464_(_23314_, _23339_, _23340_);
  or g_54465_(_23313_, _23325_, _23342_);
  or g_54466_(_23340_, _23342_, _23343_);
  or g_54467_(_23317_, _23323_, _23344_);
  or g_54468_(_23326_, _23344_, _23345_);
  or g_54469_(_23343_, _23345_, _23346_);
  or g_54470_(_23338_, _23346_, _23347_);
  or g_54471_(_23331_, _23347_, _23348_);
  xor g_54472_(out[1], out[385], _23349_);
  and g_54473_(out[11], _39768_, _23350_);
  xor g_54474_(out[9], out[393], _23351_);
  xor g_54475_(out[0], out[384], _23353_);
  xor g_54476_(out[14], out[398], _23354_);
  xor g_54477_(out[4], out[388], _23355_);
  or g_54478_(_23354_, _23355_, _23356_);
  xor g_54479_(out[13], out[397], _23357_);
  xor g_54480_(out[3], out[387], _23358_);
  and g_54481_(_39438_, out[395], _23359_);
  xor g_54482_(out[6], out[390], _23360_);
  xor g_54483_(out[10], out[394], _23361_);
  xor g_54484_(out[5], out[389], _23362_);
  xor g_54485_(out[15], out[399], _23364_);
  xor g_54486_(out[8], out[392], _23365_);
  or g_54487_(_23357_, _23365_, _23366_);
  xor g_54488_(out[2], out[386], _23367_);
  or g_54489_(_23361_, _23367_, _23368_);
  or g_54490_(_23366_, _23368_, _23369_);
  or g_54491_(_23351_, _23358_, _23370_);
  or g_54492_(_23362_, _23370_, _23371_);
  or g_54493_(_23369_, _23371_, _23372_);
  or g_54494_(_23356_, _23372_, _23373_);
  xor g_54495_(out[12], out[396], _23375_);
  or g_54496_(_23359_, _23375_, _23376_);
  xor g_54497_(out[7], out[391], _23377_);
  or g_54498_(_23360_, _23377_, _23378_);
  or g_54499_(_23376_, _23378_, _23379_);
  or g_54500_(_23349_, _23350_, _23380_);
  or g_54501_(_23364_, _23380_, _23381_);
  or g_54502_(_23379_, _23381_, _23382_);
  or g_54503_(_23353_, _23382_, _23383_);
  or g_54504_(_23373_, _23383_, _23384_);
  xor g_54505_(out[316], out[380], _23386_);
  and g_54506_(_39724_, out[379], _23387_);
  xor g_54507_(out[312], out[376], _23388_);
  xor g_54508_(out[310], out[374], _23389_);
  xor g_54509_(out[317], out[381], _23390_);
  xor g_54510_(out[318], out[382], _23391_);
  xor g_54511_(out[306], out[370], _23392_);
  xor g_54512_(out[313], out[377], _23393_);
  xor g_54513_(out[309], out[373], _23394_);
  xor g_54514_(out[305], out[369], _23395_);
  and g_54515_(out[315], _39757_, _23397_);
  or g_54516_(_23388_, _23390_, _23398_);
  xor g_54517_(out[319], out[383], _23399_);
  xor g_54518_(out[314], out[378], _23400_);
  xor g_54519_(out[308], out[372], _23401_);
  xor g_54520_(out[307], out[371], _23402_);
  xor g_54521_(out[304], out[368], _23403_);
  or g_54522_(_23392_, _23400_, _23404_);
  or g_54523_(_23398_, _23404_, _23405_);
  or g_54524_(_23393_, _23402_, _23406_);
  or g_54525_(_23394_, _23406_, _23408_);
  or g_54526_(_23405_, _23408_, _23409_);
  or g_54527_(_23391_, _23401_, _23410_);
  or g_54528_(_23409_, _23410_, _23411_);
  or g_54529_(_23386_, _23387_, _23412_);
  xor g_54530_(out[311], out[375], _23413_);
  or g_54531_(_23389_, _23413_, _23414_);
  or g_54532_(_23412_, _23414_, _23415_);
  or g_54533_(_23395_, _23397_, _23416_);
  or g_54534_(_23399_, _23416_, _23417_);
  or g_54535_(_23415_, _23417_, _23419_);
  or g_54536_(_23403_, _23419_, _23420_);
  or g_54537_(_23411_, _23420_, _23421_);
  xor g_54538_(out[295], out[375], _23422_);
  and g_54539_(_39702_, out[379], _23423_);
  xor g_54540_(out[302], out[382], _23424_);
  xor g_54541_(out[296], out[376], _23425_);
  xor g_54542_(out[289], out[369], _23426_);
  xor g_54543_(out[301], out[381], _23427_);
  xor g_54544_(out[297], out[377], _23428_);
  xor g_54545_(out[292], out[372], _23430_);
  xor g_54546_(out[290], out[370], _23431_);
  and g_54547_(out[299], _39757_, _23432_);
  xor g_54548_(out[291], out[371], _23433_);
  xor g_54549_(out[294], out[374], _23434_);
  xor g_54550_(out[303], out[383], _23435_);
  xor g_54551_(out[298], out[378], _23436_);
  xor g_54552_(out[293], out[373], _23437_);
  xor g_54553_(out[288], out[368], _23438_);
  or g_54554_(_23424_, _23430_, _23439_);
  or g_54555_(_23425_, _23427_, _23441_);
  or g_54556_(_23431_, _23436_, _23442_);
  or g_54557_(_23441_, _23442_, _23443_);
  or g_54558_(_23428_, _23433_, _23444_);
  or g_54559_(_23437_, _23438_, _23445_);
  or g_54560_(_23444_, _23445_, _23446_);
  or g_54561_(_23443_, _23446_, _23447_);
  xor g_54562_(out[300], out[380], _23448_);
  or g_54563_(_23423_, _23448_, _23449_);
  or g_54564_(_23422_, _23434_, _23450_);
  or g_54565_(_23449_, _23450_, _23452_);
  or g_54566_(_23426_, _23432_, _23453_);
  or g_54567_(_23435_, _23453_, _23454_);
  or g_54568_(_23452_, _23454_, _23455_);
  or g_54569_(_23447_, _23455_, _23456_);
  or g_54570_(_23439_, _23456_, _23457_);
  not g_54571_(_23457_, _23458_);
  xor g_54572_(out[273], out[369], _23459_);
  and g_54573_(out[283], _39757_, _23460_);
  xor g_54574_(out[286], out[382], _23461_);
  xor g_54575_(out[275], out[371], _23463_);
  xor g_54576_(out[276], out[372], _23464_);
  xor g_54577_(out[274], out[370], _23465_);
  xor g_54578_(out[281], out[377], _23466_);
  xor g_54579_(out[272], out[368], _23467_);
  and g_54580_(_39691_, out[379], _23468_);
  xor g_54581_(out[278], out[374], _23469_);
  xor g_54582_(out[282], out[378], _23470_);
  xor g_54583_(out[277], out[373], _23471_);
  xor g_54584_(out[287], out[383], _23472_);
  xor g_54585_(out[285], out[381], _23474_);
  xor g_54586_(out[280], out[376], _23475_);
  or g_54587_(_23461_, _23464_, _23476_);
  or g_54588_(_23474_, _23475_, _23477_);
  or g_54589_(_23465_, _23470_, _23478_);
  or g_54590_(_23477_, _23478_, _23479_);
  or g_54591_(_23463_, _23466_, _23480_);
  or g_54592_(_23467_, _23471_, _23481_);
  or g_54593_(_23480_, _23481_, _23482_);
  or g_54594_(_23479_, _23482_, _23483_);
  xor g_54595_(out[284], out[380], _23485_);
  or g_54596_(_23468_, _23485_, _23486_);
  xor g_54597_(out[279], out[375], _23487_);
  or g_54598_(_23469_, _23487_, _23488_);
  or g_54599_(_23486_, _23488_, _23489_);
  or g_54600_(_23459_, _23460_, _23490_);
  or g_54601_(_23472_, _23490_, _23491_);
  or g_54602_(_23489_, _23491_, _23492_);
  or g_54603_(_23483_, _23492_, _23493_);
  or g_54604_(_23476_, _23493_, _23494_);
  xor g_54605_(out[263], out[375], _23496_);
  and g_54606_(_39680_, out[379], _23497_);
  xor g_54607_(out[270], out[382], _23498_);
  xor g_54608_(out[264], out[376], _23499_);
  xor g_54609_(out[257], out[369], _23500_);
  xor g_54610_(out[269], out[381], _23501_);
  xor g_54611_(out[265], out[377], _23502_);
  xor g_54612_(out[260], out[372], _23503_);
  xor g_54613_(out[258], out[370], _23504_);
  and g_54614_(out[267], _39757_, _23505_);
  xor g_54615_(out[259], out[371], _23507_);
  xor g_54616_(out[262], out[374], _23508_);
  xor g_54617_(out[271], out[383], _23509_);
  xor g_54618_(out[266], out[378], _23510_);
  xor g_54619_(out[261], out[373], _23511_);
  xor g_54620_(out[256], out[368], _23512_);
  or g_54621_(_23498_, _23503_, _23513_);
  or g_54622_(_23499_, _23501_, _23514_);
  or g_54623_(_23504_, _23510_, _23515_);
  or g_54624_(_23514_, _23515_, _23516_);
  or g_54625_(_23502_, _23507_, _23518_);
  or g_54626_(_23511_, _23512_, _23519_);
  or g_54627_(_23518_, _23519_, _23520_);
  or g_54628_(_23516_, _23520_, _23521_);
  xor g_54629_(out[268], out[380], _23522_);
  or g_54630_(_23497_, _23522_, _23523_);
  or g_54631_(_23496_, _23508_, _23524_);
  or g_54632_(_23523_, _23524_, _23525_);
  or g_54633_(_23500_, _23505_, _23526_);
  or g_54634_(_23509_, _23526_, _23527_);
  or g_54635_(_23525_, _23527_, _23529_);
  or g_54636_(_23521_, _23529_, _23530_);
  or g_54637_(_23513_, _23530_, _23531_);
  xor g_54638_(out[248], out[376], _23532_);
  xor g_54639_(out[245], out[373], _23533_);
  xor g_54640_(out[243], out[371], _23534_);
  xor g_54641_(out[254], out[382], _23535_);
  xor g_54642_(out[253], out[381], _23536_);
  xor g_54643_(out[242], out[370], _23537_);
  xor g_54644_(out[249], out[377], _23538_);
  xor g_54645_(out[246], out[374], _23540_);
  xor g_54646_(out[255], out[383], _23541_);
  xor g_54647_(out[250], out[378], _23542_);
  xor g_54648_(out[244], out[372], _23543_);
  xor g_54649_(out[240], out[368], _23544_);
  and g_54650_(_39669_, out[379], _23545_);
  and g_54651_(out[251], _39757_, _23546_);
  or g_54652_(_23532_, _23536_, _23547_);
  xor g_54653_(out[241], out[369], _23548_);
  or g_54654_(_23537_, _23542_, _23549_);
  or g_54655_(_23547_, _23549_, _23551_);
  or g_54656_(_23534_, _23538_, _23552_);
  or g_54657_(_23533_, _23552_, _23553_);
  or g_54658_(_23551_, _23553_, _23554_);
  or g_54659_(_23535_, _23543_, _23555_);
  or g_54660_(_23554_, _23555_, _23556_);
  xor g_54661_(out[252], out[380], _23557_);
  or g_54662_(_23545_, _23557_, _23558_);
  xor g_54663_(out[247], out[375], _23559_);
  or g_54664_(_23540_, _23559_, _23560_);
  or g_54665_(_23558_, _23560_, _23562_);
  or g_54666_(_23546_, _23548_, _23563_);
  or g_54667_(_23541_, _23563_, _23564_);
  or g_54668_(_23562_, _23564_, _23565_);
  or g_54669_(_23544_, _23565_, _23566_);
  or g_54670_(_23556_, _23566_, _23567_);
  not g_54671_(_23567_, _23568_);
  xor g_54672_(out[231], out[375], _23569_);
  and g_54673_(_39658_, out[379], _23570_);
  xor g_54674_(out[238], out[382], _23571_);
  xor g_54675_(out[232], out[376], _23573_);
  xor g_54676_(out[225], out[369], _23574_);
  xor g_54677_(out[237], out[381], _23575_);
  xor g_54678_(out[233], out[377], _23576_);
  xor g_54679_(out[228], out[372], _23577_);
  xor g_54680_(out[226], out[370], _23578_);
  and g_54681_(out[235], _39757_, _23579_);
  xor g_54682_(out[227], out[371], _23580_);
  xor g_54683_(out[230], out[374], _23581_);
  xor g_54684_(out[239], out[383], _23582_);
  xor g_54685_(out[234], out[378], _23584_);
  xor g_54686_(out[229], out[373], _23585_);
  xor g_54687_(out[224], out[368], _23586_);
  or g_54688_(_23571_, _23577_, _23587_);
  or g_54689_(_23573_, _23575_, _23588_);
  or g_54690_(_23578_, _23584_, _23589_);
  or g_54691_(_23588_, _23589_, _23590_);
  or g_54692_(_23576_, _23580_, _23591_);
  or g_54693_(_23585_, _23586_, _23592_);
  or g_54694_(_23591_, _23592_, _23593_);
  or g_54695_(_23590_, _23593_, _23595_);
  xor g_54696_(out[236], out[380], _23596_);
  or g_54697_(_23570_, _23596_, _23597_);
  or g_54698_(_23569_, _23581_, _23598_);
  or g_54699_(_23597_, _23598_, _23599_);
  or g_54700_(_23574_, _23579_, _23600_);
  or g_54701_(_23582_, _23600_, _23601_);
  or g_54702_(_23599_, _23601_, _23602_);
  or g_54703_(_23595_, _23602_, _23603_);
  or g_54704_(_23587_, _23603_, _23604_);
  xor g_54705_(out[218], out[378], _23606_);
  xor g_54706_(out[210], out[370], _23607_);
  xor g_54707_(out[209], out[369], _23608_);
  and g_54708_(_39647_, out[379], _23609_);
  and g_54709_(out[219], _39757_, _23610_);
  xor g_54710_(out[221], out[381], _23611_);
  xor g_54711_(out[211], out[371], _23612_);
  xor g_54712_(out[222], out[382], _23613_);
  xor g_54713_(out[220], out[380], _23614_);
  xor g_54714_(out[216], out[376], _23615_);
  xor g_54715_(out[223], out[383], _23617_);
  xor g_54716_(out[213], out[373], _23618_);
  xor g_54717_(out[214], out[374], _23619_);
  xor g_54718_(out[208], out[368], _23620_);
  xor g_54719_(out[212], out[372], _23621_);
  or g_54720_(_23611_, _23615_, _23622_);
  xor g_54721_(out[217], out[377], _23623_);
  or g_54722_(_23606_, _23607_, _23624_);
  or g_54723_(_23622_, _23624_, _23625_);
  or g_54724_(_23612_, _23623_, _23626_);
  or g_54725_(_23618_, _23626_, _23628_);
  or g_54726_(_23625_, _23628_, _23629_);
  or g_54727_(_23613_, _23621_, _23630_);
  or g_54728_(_23629_, _23630_, _23631_);
  or g_54729_(_23609_, _23614_, _23632_);
  xor g_54730_(out[215], out[375], _23633_);
  or g_54731_(_23619_, _23633_, _23634_);
  or g_54732_(_23632_, _23634_, _23635_);
  or g_54733_(_23608_, _23610_, _23636_);
  or g_54734_(_23617_, _23636_, _23637_);
  or g_54735_(_23635_, _23637_, _23639_);
  or g_54736_(_23620_, _23639_, _23640_);
  or g_54737_(_23631_, _23640_, _23641_);
  xor g_54738_(out[199], out[375], _23642_);
  and g_54739_(_39636_, out[379], _23643_);
  xor g_54740_(out[206], out[382], _23644_);
  xor g_54741_(out[200], out[376], _23645_);
  xor g_54742_(out[193], out[369], _23646_);
  xor g_54743_(out[205], out[381], _23647_);
  xor g_54744_(out[201], out[377], _23648_);
  xor g_54745_(out[196], out[372], _23650_);
  xor g_54746_(out[194], out[370], _23651_);
  and g_54747_(out[203], _39757_, _23652_);
  xor g_54748_(out[195], out[371], _23653_);
  xor g_54749_(out[198], out[374], _23654_);
  xor g_54750_(out[207], out[383], _23655_);
  xor g_54751_(out[202], out[378], _23656_);
  xor g_54752_(out[197], out[373], _23657_);
  xor g_54753_(out[192], out[368], _23658_);
  or g_54754_(_23644_, _23650_, _23659_);
  or g_54755_(_23645_, _23647_, _23661_);
  or g_54756_(_23651_, _23656_, _23662_);
  or g_54757_(_23661_, _23662_, _23663_);
  or g_54758_(_23648_, _23653_, _23664_);
  or g_54759_(_23657_, _23658_, _23665_);
  or g_54760_(_23664_, _23665_, _23666_);
  or g_54761_(_23663_, _23666_, _23667_);
  xor g_54762_(out[204], out[380], _23668_);
  or g_54763_(_23643_, _23668_, _23669_);
  or g_54764_(_23642_, _23654_, _23670_);
  or g_54765_(_23669_, _23670_, _23672_);
  or g_54766_(_23646_, _23652_, _23673_);
  or g_54767_(_23655_, _23673_, _23674_);
  or g_54768_(_23672_, _23674_, _23675_);
  or g_54769_(_23667_, _23675_, _23676_);
  or g_54770_(_23659_, _23676_, _23677_);
  xor g_54771_(out[184], out[376], _23678_);
  xor g_54772_(out[181], out[373], _23679_);
  xor g_54773_(out[179], out[371], _23680_);
  xor g_54774_(out[190], out[382], _23681_);
  xor g_54775_(out[189], out[381], _23683_);
  xor g_54776_(out[178], out[370], _23684_);
  xor g_54777_(out[185], out[377], _23685_);
  xor g_54778_(out[182], out[374], _23686_);
  xor g_54779_(out[191], out[383], _23687_);
  xor g_54780_(out[186], out[378], _23688_);
  xor g_54781_(out[180], out[372], _23689_);
  xor g_54782_(out[176], out[368], _23690_);
  and g_54783_(_39625_, out[379], _23691_);
  and g_54784_(out[187], _39757_, _23692_);
  or g_54785_(_23678_, _23683_, _23694_);
  xor g_54786_(out[177], out[369], _23695_);
  or g_54787_(_23684_, _23688_, _23696_);
  or g_54788_(_23694_, _23696_, _23697_);
  or g_54789_(_23680_, _23685_, _23698_);
  or g_54790_(_23679_, _23698_, _23699_);
  or g_54791_(_23697_, _23699_, _23700_);
  or g_54792_(_23681_, _23689_, _23701_);
  or g_54793_(_23700_, _23701_, _23702_);
  xor g_54794_(out[188], out[380], _23703_);
  or g_54795_(_23691_, _23703_, _23705_);
  xor g_54796_(out[183], out[375], _23706_);
  or g_54797_(_23686_, _23706_, _23707_);
  or g_54798_(_23705_, _23707_, _23708_);
  or g_54799_(_23692_, _23695_, _23709_);
  or g_54800_(_23687_, _23709_, _23710_);
  or g_54801_(_23708_, _23710_, _23711_);
  or g_54802_(_23690_, _23711_, _23712_);
  or g_54803_(_23702_, _23712_, _23713_);
  xor g_54804_(out[167], out[375], _23714_);
  and g_54805_(_39614_, out[379], _23716_);
  xor g_54806_(out[174], out[382], _23717_);
  xor g_54807_(out[168], out[376], _23718_);
  xor g_54808_(out[161], out[369], _23719_);
  xor g_54809_(out[173], out[381], _23720_);
  xor g_54810_(out[169], out[377], _23721_);
  xor g_54811_(out[164], out[372], _23722_);
  xor g_54812_(out[162], out[370], _23723_);
  and g_54813_(out[171], _39757_, _23724_);
  xor g_54814_(out[163], out[371], _23725_);
  xor g_54815_(out[166], out[374], _23727_);
  xor g_54816_(out[175], out[383], _23728_);
  xor g_54817_(out[170], out[378], _23729_);
  xor g_54818_(out[165], out[373], _23730_);
  xor g_54819_(out[160], out[368], _23731_);
  or g_54820_(_23717_, _23722_, _23732_);
  or g_54821_(_23718_, _23720_, _23733_);
  or g_54822_(_23723_, _23729_, _23734_);
  or g_54823_(_23733_, _23734_, _23735_);
  or g_54824_(_23721_, _23725_, _23736_);
  or g_54825_(_23730_, _23731_, _23738_);
  or g_54826_(_23736_, _23738_, _23739_);
  or g_54827_(_23735_, _23739_, _23740_);
  xor g_54828_(out[172], out[380], _23741_);
  or g_54829_(_23716_, _23741_, _23742_);
  or g_54830_(_23714_, _23727_, _23743_);
  or g_54831_(_23742_, _23743_, _23744_);
  or g_54832_(_23719_, _23724_, _23745_);
  or g_54833_(_23728_, _23745_, _23746_);
  or g_54834_(_23744_, _23746_, _23747_);
  or g_54835_(_23740_, _23747_, _23749_);
  or g_54836_(_23732_, _23749_, _23750_);
  not g_54837_(_23750_, _23751_);
  and g_54838_(out[155], _39757_, _23752_);
  xor g_54839_(out[148], out[372], _23753_);
  xor g_54840_(out[158], out[382], _23754_);
  or g_54841_(_23753_, _23754_, _23755_);
  xor g_54842_(out[157], out[381], _23756_);
  xor g_54843_(out[147], out[371], _23757_);
  xor g_54844_(out[144], out[368], _23758_);
  and g_54845_(_39603_, out[379], _23760_);
  xor g_54846_(out[154], out[378], _23761_);
  xor g_54847_(out[159], out[383], _23762_);
  xor g_54848_(out[150], out[374], _23763_);
  xor g_54849_(out[149], out[373], _23764_);
  xor g_54850_(out[152], out[376], _23765_);
  or g_54851_(_23756_, _23765_, _23766_);
  xor g_54852_(out[146], out[370], _23767_);
  xor g_54853_(out[153], out[377], _23768_);
  xor g_54854_(out[145], out[369], _23769_);
  or g_54855_(_23761_, _23767_, _23771_);
  or g_54856_(_23766_, _23771_, _23772_);
  or g_54857_(_23757_, _23768_, _23773_);
  or g_54858_(_23764_, _23773_, _23774_);
  or g_54859_(_23772_, _23774_, _23775_);
  or g_54860_(_23755_, _23775_, _23776_);
  xor g_54861_(out[156], out[380], _23777_);
  or g_54862_(_23760_, _23777_, _23778_);
  xor g_54863_(out[151], out[375], _23779_);
  or g_54864_(_23763_, _23779_, _23780_);
  or g_54865_(_23778_, _23780_, _23782_);
  or g_54866_(_23752_, _23769_, _23783_);
  or g_54867_(_23762_, _23783_, _23784_);
  or g_54868_(_23782_, _23784_, _23785_);
  or g_54869_(_23758_, _23785_, _23786_);
  or g_54870_(_23776_, _23786_, _23787_);
  xor g_54871_(out[135], out[375], _23788_);
  and g_54872_(_39592_, out[379], _23789_);
  xor g_54873_(out[142], out[382], _23790_);
  xor g_54874_(out[136], out[376], _23791_);
  xor g_54875_(out[129], out[369], _23793_);
  xor g_54876_(out[141], out[381], _23794_);
  xor g_54877_(out[137], out[377], _23795_);
  xor g_54878_(out[132], out[372], _23796_);
  xor g_54879_(out[130], out[370], _23797_);
  and g_54880_(out[139], _39757_, _23798_);
  xor g_54881_(out[131], out[371], _23799_);
  xor g_54882_(out[134], out[374], _23800_);
  xor g_54883_(out[143], out[383], _23801_);
  xor g_54884_(out[138], out[378], _23802_);
  xor g_54885_(out[133], out[373], _23804_);
  xor g_54886_(out[128], out[368], _23805_);
  or g_54887_(_23790_, _23796_, _23806_);
  or g_54888_(_23791_, _23794_, _23807_);
  or g_54889_(_23797_, _23802_, _23808_);
  or g_54890_(_23807_, _23808_, _23809_);
  or g_54891_(_23795_, _23799_, _23810_);
  or g_54892_(_23804_, _23805_, _23811_);
  or g_54893_(_23810_, _23811_, _23812_);
  or g_54894_(_23809_, _23812_, _23813_);
  xor g_54895_(out[140], out[380], _23815_);
  or g_54896_(_23789_, _23815_, _23816_);
  or g_54897_(_23788_, _23800_, _23817_);
  or g_54898_(_23816_, _23817_, _23818_);
  or g_54899_(_23793_, _23798_, _23819_);
  or g_54900_(_23801_, _23819_, _23820_);
  or g_54901_(_23818_, _23820_, _23821_);
  or g_54902_(_23813_, _23821_, _23822_);
  or g_54903_(_23806_, _23822_, _23823_);
  xor g_54904_(out[113], out[369], _23824_);
  and g_54905_(out[123], _39757_, _23826_);
  xor g_54906_(out[116], out[372], _23827_);
  xor g_54907_(out[118], out[374], _23828_);
  xor g_54908_(out[115], out[371], _23829_);
  xor g_54909_(out[119], out[375], _23830_);
  and g_54910_(_39581_, out[379], _23831_);
  xor g_54911_(out[122], out[378], _23832_);
  xor g_54912_(out[114], out[370], _23833_);
  or g_54913_(_23832_, _23833_, _23834_);
  xor g_54914_(out[126], out[382], _23835_);
  xor g_54915_(out[112], out[368], _23837_);
  xor g_54916_(out[125], out[381], _23838_);
  xor g_54917_(out[120], out[376], _23839_);
  or g_54918_(_23838_, _23839_, _23840_);
  xor g_54919_(out[121], out[377], _23841_);
  xor g_54920_(out[127], out[383], _23842_);
  xor g_54921_(out[117], out[373], _23843_);
  or g_54922_(_23834_, _23840_, _23844_);
  or g_54923_(_23829_, _23841_, _23845_);
  or g_54924_(_23843_, _23845_, _23846_);
  or g_54925_(_23844_, _23846_, _23848_);
  or g_54926_(_23827_, _23835_, _23849_);
  or g_54927_(_23848_, _23849_, _23850_);
  xor g_54928_(out[124], out[380], _23851_);
  or g_54929_(_23831_, _23851_, _23852_);
  or g_54930_(_23828_, _23830_, _23853_);
  or g_54931_(_23852_, _23853_, _23854_);
  or g_54932_(_23824_, _23826_, _23855_);
  or g_54933_(_23842_, _23855_, _23856_);
  or g_54934_(_23854_, _23856_, _23857_);
  or g_54935_(_23837_, _23857_, _23859_);
  or g_54936_(_23850_, _23859_, _23860_);
  not g_54937_(_23860_, _23861_);
  xor g_54938_(out[103], out[375], _23862_);
  and g_54939_(_39570_, out[379], _23863_);
  xor g_54940_(out[110], out[382], _23864_);
  xor g_54941_(out[104], out[376], _23865_);
  xor g_54942_(out[97], out[369], _23866_);
  xor g_54943_(out[109], out[381], _23867_);
  xor g_54944_(out[105], out[377], _23868_);
  xor g_54945_(out[100], out[372], _23870_);
  xor g_54946_(out[98], out[370], _23871_);
  and g_54947_(out[107], _39757_, _23872_);
  xor g_54948_(out[99], out[371], _23873_);
  xor g_54949_(out[102], out[374], _23874_);
  xor g_54950_(out[111], out[383], _23875_);
  xor g_54951_(out[106], out[378], _23876_);
  xor g_54952_(out[101], out[373], _23877_);
  xor g_54953_(out[96], out[368], _23878_);
  or g_54954_(_23864_, _23870_, _23879_);
  or g_54955_(_23865_, _23867_, _23881_);
  or g_54956_(_23871_, _23876_, _23882_);
  or g_54957_(_23881_, _23882_, _23883_);
  or g_54958_(_23868_, _23873_, _23884_);
  or g_54959_(_23877_, _23878_, _23885_);
  or g_54960_(_23884_, _23885_, _23886_);
  or g_54961_(_23883_, _23886_, _23887_);
  xor g_54962_(out[108], out[380], _23888_);
  or g_54963_(_23863_, _23888_, _23889_);
  or g_54964_(_23862_, _23874_, _23890_);
  or g_54965_(_23889_, _23890_, _23892_);
  or g_54966_(_23866_, _23872_, _23893_);
  or g_54967_(_23875_, _23893_, _23894_);
  or g_54968_(_23892_, _23894_, _23895_);
  or g_54969_(_23887_, _23895_, _23896_);
  or g_54970_(_23879_, _23896_, _23897_);
  xor g_54971_(out[84], out[372], _23898_);
  xor g_54972_(out[92], out[380], _23899_);
  and g_54973_(_39559_, out[379], _23900_);
  xor g_54974_(out[90], out[378], _23901_);
  xor g_54975_(out[86], out[374], _23903_);
  xor g_54976_(out[85], out[373], _23904_);
  xor g_54977_(out[83], out[371], _23905_);
  xor g_54978_(out[93], out[381], _23906_);
  xor g_54979_(out[94], out[382], _23907_);
  xor g_54980_(out[81], out[369], _23908_);
  xor g_54981_(out[82], out[370], _23909_);
  and g_54982_(out[91], _39757_, _23910_);
  xor g_54983_(out[80], out[368], _23911_);
  xor g_54984_(out[95], out[383], _23912_);
  xor g_54985_(out[88], out[376], _23914_);
  or g_54986_(_23906_, _23914_, _23915_);
  xor g_54987_(out[89], out[377], _23916_);
  or g_54988_(_23901_, _23909_, _23917_);
  or g_54989_(_23915_, _23917_, _23918_);
  or g_54990_(_23905_, _23916_, _23919_);
  or g_54991_(_23904_, _23919_, _23920_);
  or g_54992_(_23918_, _23920_, _23921_);
  or g_54993_(_23898_, _23907_, _23922_);
  or g_54994_(_23921_, _23922_, _23923_);
  or g_54995_(_23899_, _23900_, _23925_);
  xor g_54996_(out[87], out[375], _23926_);
  or g_54997_(_23903_, _23926_, _23927_);
  or g_54998_(_23925_, _23927_, _23928_);
  or g_54999_(_23908_, _23910_, _23929_);
  or g_55000_(_23912_, _23929_, _23930_);
  or g_55001_(_23928_, _23930_, _23931_);
  or g_55002_(_23911_, _23931_, _23932_);
  or g_55003_(_23923_, _23932_, _23933_);
  xor g_55004_(out[71], out[375], _23934_);
  and g_55005_(_39548_, out[379], _23936_);
  xor g_55006_(out[78], out[382], _23937_);
  xor g_55007_(out[72], out[376], _23938_);
  xor g_55008_(out[65], out[369], _23939_);
  xor g_55009_(out[77], out[381], _23940_);
  xor g_55010_(out[73], out[377], _23941_);
  xor g_55011_(out[68], out[372], _23942_);
  xor g_55012_(out[66], out[370], _23943_);
  and g_55013_(out[75], _39757_, _23944_);
  xor g_55014_(out[67], out[371], _23945_);
  xor g_55015_(out[70], out[374], _23947_);
  xor g_55016_(out[79], out[383], _23948_);
  xor g_55017_(out[74], out[378], _23949_);
  xor g_55018_(out[69], out[373], _23950_);
  xor g_55019_(out[64], out[368], _23951_);
  or g_55020_(_23937_, _23942_, _23952_);
  or g_55021_(_23938_, _23940_, _23953_);
  or g_55022_(_23943_, _23949_, _23954_);
  or g_55023_(_23953_, _23954_, _23955_);
  or g_55024_(_23941_, _23945_, _23956_);
  or g_55025_(_23950_, _23951_, _23958_);
  or g_55026_(_23956_, _23958_, _23959_);
  or g_55027_(_23955_, _23959_, _23960_);
  xor g_55028_(out[76], out[380], _23961_);
  or g_55029_(_23936_, _23961_, _23962_);
  or g_55030_(_23934_, _23947_, _23963_);
  or g_55031_(_23962_, _23963_, _23964_);
  or g_55032_(_23939_, _23944_, _23965_);
  or g_55033_(_23948_, _23965_, _23966_);
  or g_55034_(_23964_, _23966_, _23967_);
  or g_55035_(_23960_, _23967_, _23969_);
  or g_55036_(_23952_, _23969_, _23970_);
  xor g_55037_(out[51], out[371], _23971_);
  xor g_55038_(out[52], out[372], _23972_);
  xor g_55039_(out[62], out[382], _23973_);
  xor g_55040_(out[50], out[370], _23974_);
  xor g_55041_(out[53], out[373], _23975_);
  xor g_55042_(out[57], out[377], _23976_);
  xor g_55043_(out[56], out[376], _23977_);
  xor g_55044_(out[63], out[383], _23978_);
  xor g_55045_(out[58], out[378], _23980_);
  xor g_55046_(out[54], out[374], _23981_);
  xor g_55047_(out[48], out[368], _23982_);
  and g_55048_(_39537_, out[379], _23983_);
  and g_55049_(out[59], _39757_, _23984_);
  xor g_55050_(out[61], out[381], _23985_);
  or g_55051_(_23977_, _23985_, _23986_);
  xor g_55052_(out[49], out[369], _23987_);
  or g_55053_(_23974_, _23980_, _23988_);
  or g_55054_(_23986_, _23988_, _23989_);
  or g_55055_(_23971_, _23976_, _23991_);
  or g_55056_(_23975_, _23991_, _23992_);
  or g_55057_(_23989_, _23992_, _23993_);
  or g_55058_(_23972_, _23973_, _23994_);
  or g_55059_(_23993_, _23994_, _23995_);
  xor g_55060_(out[60], out[380], _23996_);
  or g_55061_(_23983_, _23996_, _23997_);
  xor g_55062_(out[55], out[375], _23998_);
  or g_55063_(_23981_, _23998_, _23999_);
  or g_55064_(_23997_, _23999_, _24000_);
  or g_55065_(_23984_, _23987_, _24002_);
  or g_55066_(_23978_, _24002_, _24003_);
  or g_55067_(_24000_, _24003_, _24004_);
  or g_55068_(_23982_, _24004_, _24005_);
  or g_55069_(_23995_, _24005_, _24006_);
  xor g_55070_(out[39], out[375], _24007_);
  and g_55071_(_39526_, out[379], _24008_);
  xor g_55072_(out[46], out[382], _24009_);
  xor g_55073_(out[40], out[376], _24010_);
  xor g_55074_(out[33], out[369], _24011_);
  xor g_55075_(out[45], out[381], _24013_);
  xor g_55076_(out[41], out[377], _24014_);
  xor g_55077_(out[36], out[372], _24015_);
  xor g_55078_(out[34], out[370], _24016_);
  and g_55079_(out[43], _39757_, _24017_);
  xor g_55080_(out[35], out[371], _24018_);
  xor g_55081_(out[38], out[374], _24019_);
  xor g_55082_(out[47], out[383], _24020_);
  xor g_55083_(out[42], out[378], _24021_);
  xor g_55084_(out[37], out[373], _24022_);
  xor g_55085_(out[32], out[368], _24024_);
  or g_55086_(_24009_, _24015_, _24025_);
  or g_55087_(_24010_, _24013_, _24026_);
  or g_55088_(_24016_, _24021_, _24027_);
  or g_55089_(_24026_, _24027_, _24028_);
  or g_55090_(_24014_, _24018_, _24029_);
  or g_55091_(_24022_, _24024_, _24030_);
  or g_55092_(_24029_, _24030_, _24031_);
  or g_55093_(_24028_, _24031_, _24032_);
  xor g_55094_(out[44], out[380], _24033_);
  or g_55095_(_24008_, _24033_, _24035_);
  or g_55096_(_24007_, _24019_, _24036_);
  or g_55097_(_24035_, _24036_, _24037_);
  or g_55098_(_24011_, _24017_, _24038_);
  or g_55099_(_24020_, _24038_, _24039_);
  or g_55100_(_24037_, _24039_, _24040_);
  or g_55101_(_24032_, _24040_, _24041_);
  or g_55102_(_24025_, _24041_, _24042_);
  not g_55103_(_24042_, _24043_);
  xor g_55104_(out[17], out[369], _24044_);
  and g_55105_(out[27], _39757_, _24046_);
  xor g_55106_(out[30], out[382], _24047_);
  xor g_55107_(out[19], out[371], _24048_);
  xor g_55108_(out[20], out[372], _24049_);
  xor g_55109_(out[18], out[370], _24050_);
  xor g_55110_(out[25], out[377], _24051_);
  xor g_55111_(out[16], out[368], _24052_);
  and g_55112_(_39493_, out[379], _24053_);
  xor g_55113_(out[22], out[374], _24054_);
  xor g_55114_(out[26], out[378], _24055_);
  xor g_55115_(out[21], out[373], _24057_);
  xor g_55116_(out[31], out[383], _24058_);
  xor g_55117_(out[29], out[381], _24059_);
  xor g_55118_(out[24], out[376], _24060_);
  or g_55119_(_24047_, _24049_, _24061_);
  or g_55120_(_24059_, _24060_, _24062_);
  or g_55121_(_24050_, _24055_, _24063_);
  or g_55122_(_24062_, _24063_, _24064_);
  or g_55123_(_24048_, _24051_, _24065_);
  or g_55124_(_24052_, _24057_, _24066_);
  or g_55125_(_24065_, _24066_, _24068_);
  or g_55126_(_24064_, _24068_, _24069_);
  xor g_55127_(out[28], out[380], _24070_);
  or g_55128_(_24053_, _24070_, _24071_);
  xor g_55129_(out[23], out[375], _24072_);
  or g_55130_(_24054_, _24072_, _24073_);
  or g_55131_(_24071_, _24073_, _24074_);
  or g_55132_(_24044_, _24046_, _24075_);
  or g_55133_(_24058_, _24075_, _24076_);
  or g_55134_(_24074_, _24076_, _24077_);
  or g_55135_(_24069_, _24077_, _24079_);
  or g_55136_(_24061_, _24079_, _24080_);
  xor g_55137_(out[1], out[369], _24081_);
  and g_55138_(_39438_, out[379], _24082_);
  and g_55139_(out[11], _39757_, _24083_);
  xor g_55140_(out[8], out[376], _24084_);
  xor g_55141_(out[10], out[378], _24085_);
  xor g_55142_(out[2], out[370], _24086_);
  xor g_55143_(out[4], out[372], _24087_);
  xor g_55144_(out[5], out[373], _24088_);
  xor g_55145_(out[9], out[377], _24090_);
  xor g_55146_(out[3], out[371], _24091_);
  xor g_55147_(out[14], out[382], _24092_);
  xor g_55148_(out[0], out[368], _24093_);
  xor g_55149_(out[15], out[383], _24094_);
  xor g_55150_(out[13], out[381], _24095_);
  or g_55151_(_24084_, _24095_, _24096_);
  xor g_55152_(out[6], out[374], _24097_);
  or g_55153_(_24085_, _24086_, _24098_);
  or g_55154_(_24096_, _24098_, _24099_);
  or g_55155_(_24090_, _24091_, _24101_);
  or g_55156_(_24088_, _24101_, _24102_);
  or g_55157_(_24099_, _24102_, _24103_);
  or g_55158_(_24087_, _24092_, _24104_);
  or g_55159_(_24103_, _24104_, _24105_);
  xor g_55160_(out[12], out[380], _24106_);
  or g_55161_(_24082_, _24106_, _24107_);
  xor g_55162_(out[7], out[375], _24108_);
  or g_55163_(_24097_, _24108_, _24109_);
  or g_55164_(_24107_, _24109_, _24110_);
  or g_55165_(_24081_, _24083_, _24112_);
  or g_55166_(_24094_, _24112_, _24113_);
  or g_55167_(_24110_, _24113_, _24114_);
  or g_55168_(_24093_, _24114_, _24115_);
  or g_55169_(_24105_, _24115_, _24116_);
  xor g_55170_(out[311], out[359], _24117_);
  and g_55171_(_39724_, out[363], _24118_);
  xor g_55172_(out[318], out[366], _24119_);
  xor g_55173_(out[312], out[360], _24120_);
  xor g_55174_(out[305], out[353], _24121_);
  xor g_55175_(out[317], out[365], _24123_);
  xor g_55176_(out[313], out[361], _24124_);
  xor g_55177_(out[308], out[356], _24125_);
  xor g_55178_(out[306], out[354], _24126_);
  and g_55179_(out[315], _39746_, _24127_);
  xor g_55180_(out[307], out[355], _24128_);
  xor g_55181_(out[310], out[358], _24129_);
  xor g_55182_(out[319], out[367], _24130_);
  xor g_55183_(out[314], out[362], _24131_);
  xor g_55184_(out[309], out[357], _24132_);
  xor g_55185_(out[304], out[352], _24134_);
  or g_55186_(_24119_, _24125_, _24135_);
  or g_55187_(_24120_, _24123_, _24136_);
  or g_55188_(_24126_, _24131_, _24137_);
  or g_55189_(_24136_, _24137_, _24138_);
  or g_55190_(_24124_, _24128_, _24139_);
  or g_55191_(_24132_, _24134_, _24140_);
  or g_55192_(_24139_, _24140_, _24141_);
  or g_55193_(_24138_, _24141_, _24142_);
  xor g_55194_(out[316], out[364], _24143_);
  or g_55195_(_24118_, _24143_, _24145_);
  or g_55196_(_24117_, _24129_, _24146_);
  or g_55197_(_24145_, _24146_, _24147_);
  or g_55198_(_24121_, _24127_, _24148_);
  or g_55199_(_24130_, _24148_, _24149_);
  or g_55200_(_24147_, _24149_, _24150_);
  or g_55201_(_24142_, _24150_, _24151_);
  or g_55202_(_24135_, _24151_, _24152_);
  not g_55203_(_24152_, _24153_);
  xor g_55204_(out[289], out[353], _24154_);
  and g_55205_(_39702_, out[363], _24156_);
  and g_55206_(out[299], _39746_, _24157_);
  xor g_55207_(out[297], out[361], _24158_);
  xor g_55208_(out[288], out[352], _24159_);
  xor g_55209_(out[302], out[366], _24160_);
  xor g_55210_(out[292], out[356], _24161_);
  or g_55211_(_24160_, _24161_, _24162_);
  xor g_55212_(out[301], out[365], _24163_);
  xor g_55213_(out[291], out[355], _24164_);
  xor g_55214_(out[300], out[364], _24165_);
  xor g_55215_(out[294], out[358], _24167_);
  xor g_55216_(out[298], out[362], _24168_);
  xor g_55217_(out[293], out[357], _24169_);
  xor g_55218_(out[303], out[367], _24170_);
  xor g_55219_(out[296], out[360], _24171_);
  or g_55220_(_24163_, _24171_, _24172_);
  xor g_55221_(out[290], out[354], _24173_);
  or g_55222_(_24168_, _24173_, _24174_);
  or g_55223_(_24172_, _24174_, _24175_);
  or g_55224_(_24158_, _24164_, _24176_);
  or g_55225_(_24169_, _24176_, _24178_);
  or g_55226_(_24175_, _24178_, _24179_);
  or g_55227_(_24162_, _24179_, _24180_);
  or g_55228_(_24156_, _24165_, _24181_);
  xor g_55229_(out[295], out[359], _24182_);
  or g_55230_(_24167_, _24182_, _24183_);
  or g_55231_(_24181_, _24183_, _24184_);
  or g_55232_(_24154_, _24157_, _24185_);
  or g_55233_(_24170_, _24185_, _24186_);
  or g_55234_(_24184_, _24186_, _24187_);
  or g_55235_(_24159_, _24187_, _24189_);
  or g_55236_(_24180_, _24189_, _24190_);
  not g_55237_(_24190_, _24191_);
  xor g_55238_(out[279], out[359], _24192_);
  and g_55239_(_39691_, out[363], _24193_);
  xor g_55240_(out[286], out[366], _24194_);
  xor g_55241_(out[280], out[360], _24195_);
  xor g_55242_(out[273], out[353], _24196_);
  xor g_55243_(out[285], out[365], _24197_);
  xor g_55244_(out[281], out[361], _24198_);
  xor g_55245_(out[276], out[356], _24200_);
  xor g_55246_(out[274], out[354], _24201_);
  and g_55247_(out[283], _39746_, _24202_);
  xor g_55248_(out[275], out[355], _24203_);
  xor g_55249_(out[278], out[358], _24204_);
  xor g_55250_(out[287], out[367], _24205_);
  xor g_55251_(out[282], out[362], _24206_);
  xor g_55252_(out[277], out[357], _24207_);
  xor g_55253_(out[272], out[352], _24208_);
  or g_55254_(_24194_, _24200_, _24209_);
  or g_55255_(_24195_, _24197_, _24211_);
  or g_55256_(_24201_, _24206_, _24212_);
  or g_55257_(_24211_, _24212_, _24213_);
  or g_55258_(_24198_, _24203_, _24214_);
  or g_55259_(_24207_, _24208_, _24215_);
  or g_55260_(_24214_, _24215_, _24216_);
  or g_55261_(_24213_, _24216_, _24217_);
  xor g_55262_(out[284], out[364], _24218_);
  or g_55263_(_24193_, _24218_, _24219_);
  or g_55264_(_24192_, _24204_, _24220_);
  or g_55265_(_24219_, _24220_, _24222_);
  or g_55266_(_24196_, _24202_, _24223_);
  or g_55267_(_24205_, _24223_, _24224_);
  or g_55268_(_24222_, _24224_, _24225_);
  or g_55269_(_24217_, _24225_, _24226_);
  or g_55270_(_24209_, _24226_, _24227_);
  xor g_55271_(out[264], out[360], _24228_);
  xor g_55272_(out[261], out[357], _24229_);
  xor g_55273_(out[259], out[355], _24230_);
  xor g_55274_(out[270], out[366], _24231_);
  xor g_55275_(out[269], out[365], _24233_);
  xor g_55276_(out[258], out[354], _24234_);
  xor g_55277_(out[265], out[361], _24235_);
  xor g_55278_(out[262], out[358], _24236_);
  xor g_55279_(out[271], out[367], _24237_);
  xor g_55280_(out[266], out[362], _24238_);
  xor g_55281_(out[260], out[356], _24239_);
  xor g_55282_(out[256], out[352], _24240_);
  and g_55283_(_39680_, out[363], _24241_);
  and g_55284_(out[267], _39746_, _24242_);
  or g_55285_(_24228_, _24233_, _24244_);
  xor g_55286_(out[257], out[353], _24245_);
  or g_55287_(_24234_, _24238_, _24246_);
  or g_55288_(_24244_, _24246_, _24247_);
  or g_55289_(_24230_, _24235_, _24248_);
  or g_55290_(_24229_, _24248_, _24249_);
  or g_55291_(_24247_, _24249_, _24250_);
  or g_55292_(_24231_, _24239_, _24251_);
  or g_55293_(_24250_, _24251_, _24252_);
  xor g_55294_(out[268], out[364], _24253_);
  or g_55295_(_24241_, _24253_, _24255_);
  xor g_55296_(out[263], out[359], _24256_);
  or g_55297_(_24236_, _24256_, _24257_);
  or g_55298_(_24255_, _24257_, _24258_);
  or g_55299_(_24242_, _24245_, _24259_);
  or g_55300_(_24237_, _24259_, _24260_);
  or g_55301_(_24258_, _24260_, _24261_);
  or g_55302_(_24240_, _24261_, _24262_);
  or g_55303_(_24252_, _24262_, _24263_);
  xor g_55304_(out[247], out[359], _24264_);
  and g_55305_(_39669_, out[363], _24266_);
  xor g_55306_(out[254], out[366], _24267_);
  xor g_55307_(out[248], out[360], _24268_);
  xor g_55308_(out[241], out[353], _24269_);
  xor g_55309_(out[253], out[365], _24270_);
  xor g_55310_(out[249], out[361], _24271_);
  xor g_55311_(out[244], out[356], _24272_);
  xor g_55312_(out[242], out[354], _24273_);
  and g_55313_(out[251], _39746_, _24274_);
  xor g_55314_(out[243], out[355], _24275_);
  xor g_55315_(out[246], out[358], _24277_);
  xor g_55316_(out[255], out[367], _24278_);
  xor g_55317_(out[250], out[362], _24279_);
  xor g_55318_(out[245], out[357], _24280_);
  xor g_55319_(out[240], out[352], _24281_);
  or g_55320_(_24267_, _24272_, _24282_);
  or g_55321_(_24268_, _24270_, _24283_);
  or g_55322_(_24273_, _24279_, _24284_);
  or g_55323_(_24283_, _24284_, _24285_);
  or g_55324_(_24271_, _24275_, _24286_);
  or g_55325_(_24280_, _24281_, _24288_);
  or g_55326_(_24286_, _24288_, _24289_);
  or g_55327_(_24285_, _24289_, _24290_);
  xor g_55328_(out[252], out[364], _24291_);
  or g_55329_(_24266_, _24291_, _24292_);
  or g_55330_(_24264_, _24277_, _24293_);
  or g_55331_(_24292_, _24293_, _24294_);
  or g_55332_(_24269_, _24274_, _24295_);
  or g_55333_(_24278_, _24295_, _24296_);
  or g_55334_(_24294_, _24296_, _24297_);
  or g_55335_(_24290_, _24297_, _24299_);
  or g_55336_(_24282_, _24299_, _24300_);
  xor g_55337_(out[236], out[364], _24301_);
  and g_55338_(_39658_, out[363], _24302_);
  xor g_55339_(out[232], out[360], _24303_);
  xor g_55340_(out[230], out[358], _24304_);
  xor g_55341_(out[237], out[365], _24305_);
  xor g_55342_(out[238], out[366], _24306_);
  xor g_55343_(out[226], out[354], _24307_);
  xor g_55344_(out[233], out[361], _24308_);
  xor g_55345_(out[229], out[357], _24310_);
  xor g_55346_(out[225], out[353], _24311_);
  and g_55347_(out[235], _39746_, _24312_);
  or g_55348_(_24303_, _24305_, _24313_);
  xor g_55349_(out[239], out[367], _24314_);
  xor g_55350_(out[234], out[362], _24315_);
  xor g_55351_(out[228], out[356], _24316_);
  xor g_55352_(out[227], out[355], _24317_);
  xor g_55353_(out[224], out[352], _24318_);
  or g_55354_(_24307_, _24315_, _24319_);
  or g_55355_(_24313_, _24319_, _24321_);
  or g_55356_(_24308_, _24317_, _24322_);
  or g_55357_(_24310_, _24322_, _24323_);
  or g_55358_(_24321_, _24323_, _24324_);
  or g_55359_(_24306_, _24316_, _24325_);
  or g_55360_(_24324_, _24325_, _24326_);
  or g_55361_(_24301_, _24302_, _24327_);
  xor g_55362_(out[231], out[359], _24328_);
  or g_55363_(_24304_, _24328_, _24329_);
  or g_55364_(_24327_, _24329_, _24330_);
  or g_55365_(_24311_, _24312_, _24332_);
  or g_55366_(_24314_, _24332_, _24333_);
  or g_55367_(_24330_, _24333_, _24334_);
  or g_55368_(_24318_, _24334_, _24335_);
  or g_55369_(_24326_, _24335_, _24336_);
  xor g_55370_(out[215], out[359], _24337_);
  and g_55371_(_39647_, out[363], _24338_);
  xor g_55372_(out[222], out[366], _24339_);
  xor g_55373_(out[216], out[360], _24340_);
  xor g_55374_(out[209], out[353], _24341_);
  xor g_55375_(out[221], out[365], _24343_);
  xor g_55376_(out[217], out[361], _24344_);
  xor g_55377_(out[212], out[356], _24345_);
  xor g_55378_(out[210], out[354], _24346_);
  and g_55379_(out[219], _39746_, _24347_);
  xor g_55380_(out[211], out[355], _24348_);
  xor g_55381_(out[214], out[358], _24349_);
  xor g_55382_(out[223], out[367], _24350_);
  xor g_55383_(out[218], out[362], _24351_);
  xor g_55384_(out[213], out[357], _24352_);
  xor g_55385_(out[208], out[352], _24354_);
  or g_55386_(_24339_, _24345_, _24355_);
  or g_55387_(_24340_, _24343_, _24356_);
  or g_55388_(_24346_, _24351_, _24357_);
  or g_55389_(_24356_, _24357_, _24358_);
  or g_55390_(_24344_, _24348_, _24359_);
  or g_55391_(_24352_, _24354_, _24360_);
  or g_55392_(_24359_, _24360_, _24361_);
  or g_55393_(_24358_, _24361_, _24362_);
  xor g_55394_(out[220], out[364], _24363_);
  or g_55395_(_24338_, _24363_, _24365_);
  or g_55396_(_24337_, _24349_, _24366_);
  or g_55397_(_24365_, _24366_, _24367_);
  or g_55398_(_24341_, _24347_, _24368_);
  or g_55399_(_24350_, _24368_, _24369_);
  or g_55400_(_24367_, _24369_, _24370_);
  or g_55401_(_24362_, _24370_, _24371_);
  or g_55402_(_24355_, _24371_, _24372_);
  xor g_55403_(out[200], out[360], _24373_);
  xor g_55404_(out[197], out[357], _24374_);
  xor g_55405_(out[195], out[355], _24376_);
  xor g_55406_(out[206], out[366], _24377_);
  xor g_55407_(out[205], out[365], _24378_);
  xor g_55408_(out[194], out[354], _24379_);
  xor g_55409_(out[201], out[361], _24380_);
  xor g_55410_(out[198], out[358], _24381_);
  xor g_55411_(out[207], out[367], _24382_);
  xor g_55412_(out[202], out[362], _24383_);
  xor g_55413_(out[196], out[356], _24384_);
  xor g_55414_(out[192], out[352], _24385_);
  and g_55415_(_39636_, out[363], _24387_);
  and g_55416_(out[203], _39746_, _24388_);
  or g_55417_(_24373_, _24378_, _24389_);
  xor g_55418_(out[193], out[353], _24390_);
  or g_55419_(_24379_, _24383_, _24391_);
  or g_55420_(_24389_, _24391_, _24392_);
  or g_55421_(_24376_, _24380_, _24393_);
  or g_55422_(_24374_, _24393_, _24394_);
  or g_55423_(_24392_, _24394_, _24395_);
  or g_55424_(_24377_, _24384_, _24396_);
  or g_55425_(_24395_, _24396_, _24398_);
  xor g_55426_(out[204], out[364], _24399_);
  or g_55427_(_24387_, _24399_, _24400_);
  xor g_55428_(out[199], out[359], _24401_);
  or g_55429_(_24381_, _24401_, _24402_);
  or g_55430_(_24400_, _24402_, _24403_);
  or g_55431_(_24388_, _24390_, _24404_);
  or g_55432_(_24382_, _24404_, _24405_);
  or g_55433_(_24403_, _24405_, _24406_);
  or g_55434_(_24385_, _24406_, _24407_);
  or g_55435_(_24398_, _24407_, _24409_);
  xor g_55436_(out[183], out[359], _24410_);
  and g_55437_(_39625_, out[363], _24411_);
  xor g_55438_(out[190], out[366], _24412_);
  xor g_55439_(out[184], out[360], _24413_);
  xor g_55440_(out[177], out[353], _24414_);
  xor g_55441_(out[189], out[365], _24415_);
  xor g_55442_(out[185], out[361], _24416_);
  xor g_55443_(out[180], out[356], _24417_);
  xor g_55444_(out[178], out[354], _24418_);
  and g_55445_(out[187], _39746_, _24420_);
  xor g_55446_(out[179], out[355], _24421_);
  xor g_55447_(out[182], out[358], _24422_);
  xor g_55448_(out[191], out[367], _24423_);
  xor g_55449_(out[186], out[362], _24424_);
  xor g_55450_(out[181], out[357], _24425_);
  xor g_55451_(out[176], out[352], _24426_);
  or g_55452_(_24412_, _24417_, _24427_);
  or g_55453_(_24413_, _24415_, _24428_);
  or g_55454_(_24418_, _24424_, _24429_);
  or g_55455_(_24428_, _24429_, _24431_);
  or g_55456_(_24416_, _24421_, _24432_);
  or g_55457_(_24425_, _24426_, _24433_);
  or g_55458_(_24432_, _24433_, _24434_);
  or g_55459_(_24431_, _24434_, _24435_);
  xor g_55460_(out[188], out[364], _24436_);
  or g_55461_(_24411_, _24436_, _24437_);
  or g_55462_(_24410_, _24422_, _24438_);
  or g_55463_(_24437_, _24438_, _24439_);
  or g_55464_(_24414_, _24420_, _24440_);
  or g_55465_(_24423_, _24440_, _24442_);
  or g_55466_(_24439_, _24442_, _24443_);
  or g_55467_(_24435_, _24443_, _24444_);
  or g_55468_(_24427_, _24444_, _24445_);
  not g_55469_(_24445_, _24446_);
  xor g_55470_(out[161], out[353], _24447_);
  and g_55471_(out[171], _39746_, _24448_);
  xor g_55472_(out[169], out[361], _24449_);
  xor g_55473_(out[160], out[352], _24450_);
  xor g_55474_(out[174], out[366], _24451_);
  xor g_55475_(out[164], out[356], _24453_);
  or g_55476_(_24451_, _24453_, _24454_);
  xor g_55477_(out[173], out[365], _24455_);
  xor g_55478_(out[163], out[355], _24456_);
  and g_55479_(_39614_, out[363], _24457_);
  xor g_55480_(out[166], out[358], _24458_);
  xor g_55481_(out[170], out[362], _24459_);
  xor g_55482_(out[165], out[357], _24460_);
  xor g_55483_(out[175], out[367], _24461_);
  xor g_55484_(out[168], out[360], _24462_);
  or g_55485_(_24455_, _24462_, _24464_);
  xor g_55486_(out[162], out[354], _24465_);
  or g_55487_(_24459_, _24465_, _24466_);
  or g_55488_(_24464_, _24466_, _24467_);
  or g_55489_(_24449_, _24456_, _24468_);
  or g_55490_(_24460_, _24468_, _24469_);
  or g_55491_(_24467_, _24469_, _24470_);
  or g_55492_(_24454_, _24470_, _24471_);
  xor g_55493_(out[172], out[364], _24472_);
  or g_55494_(_24457_, _24472_, _24473_);
  xor g_55495_(out[167], out[359], _24475_);
  or g_55496_(_24458_, _24475_, _24476_);
  or g_55497_(_24473_, _24476_, _24477_);
  or g_55498_(_24447_, _24448_, _24478_);
  or g_55499_(_24461_, _24478_, _24479_);
  or g_55500_(_24477_, _24479_, _24480_);
  or g_55501_(_24450_, _24480_, _24481_);
  or g_55502_(_24471_, _24481_, _24482_);
  xor g_55503_(out[151], out[359], _24483_);
  and g_55504_(_39603_, out[363], _24484_);
  xor g_55505_(out[158], out[366], _24486_);
  xor g_55506_(out[152], out[360], _24487_);
  xor g_55507_(out[145], out[353], _24488_);
  xor g_55508_(out[157], out[365], _24489_);
  xor g_55509_(out[153], out[361], _24490_);
  xor g_55510_(out[148], out[356], _24491_);
  xor g_55511_(out[146], out[354], _24492_);
  and g_55512_(out[155], _39746_, _24493_);
  xor g_55513_(out[147], out[355], _24494_);
  xor g_55514_(out[150], out[358], _24495_);
  xor g_55515_(out[159], out[367], _24497_);
  xor g_55516_(out[154], out[362], _24498_);
  xor g_55517_(out[149], out[357], _24499_);
  xor g_55518_(out[144], out[352], _24500_);
  or g_55519_(_24486_, _24491_, _24501_);
  or g_55520_(_24487_, _24489_, _24502_);
  or g_55521_(_24492_, _24498_, _24503_);
  or g_55522_(_24502_, _24503_, _24504_);
  or g_55523_(_24490_, _24494_, _24505_);
  or g_55524_(_24499_, _24500_, _24506_);
  or g_55525_(_24505_, _24506_, _24508_);
  or g_55526_(_24504_, _24508_, _24509_);
  xor g_55527_(out[156], out[364], _24510_);
  or g_55528_(_24484_, _24510_, _24511_);
  or g_55529_(_24483_, _24495_, _24512_);
  or g_55530_(_24511_, _24512_, _24513_);
  or g_55531_(_24488_, _24493_, _24514_);
  or g_55532_(_24497_, _24514_, _24515_);
  or g_55533_(_24513_, _24515_, _24516_);
  or g_55534_(_24509_, _24516_, _24517_);
  or g_55535_(_24501_, _24517_, _24519_);
  xor g_55536_(out[129], out[353], _24520_);
  and g_55537_(out[139], _39746_, _24521_);
  xor g_55538_(out[137], out[361], _24522_);
  xor g_55539_(out[128], out[352], _24523_);
  xor g_55540_(out[142], out[366], _24524_);
  xor g_55541_(out[132], out[356], _24525_);
  or g_55542_(_24524_, _24525_, _24526_);
  xor g_55543_(out[141], out[365], _24527_);
  xor g_55544_(out[131], out[355], _24528_);
  and g_55545_(_39592_, out[363], _24530_);
  xor g_55546_(out[134], out[358], _24531_);
  xor g_55547_(out[138], out[362], _24532_);
  xor g_55548_(out[133], out[357], _24533_);
  xor g_55549_(out[143], out[367], _24534_);
  xor g_55550_(out[136], out[360], _24535_);
  or g_55551_(_24527_, _24535_, _24536_);
  xor g_55552_(out[130], out[354], _24537_);
  or g_55553_(_24532_, _24537_, _24538_);
  or g_55554_(_24536_, _24538_, _24539_);
  or g_55555_(_24522_, _24528_, _24541_);
  or g_55556_(_24533_, _24541_, _24542_);
  or g_55557_(_24539_, _24542_, _24543_);
  or g_55558_(_24526_, _24543_, _24544_);
  xor g_55559_(out[140], out[364], _24545_);
  or g_55560_(_24530_, _24545_, _24546_);
  xor g_55561_(out[135], out[359], _24547_);
  or g_55562_(_24531_, _24547_, _24548_);
  or g_55563_(_24546_, _24548_, _24549_);
  or g_55564_(_24520_, _24521_, _24550_);
  or g_55565_(_24534_, _24550_, _24552_);
  or g_55566_(_24549_, _24552_, _24553_);
  or g_55567_(_24523_, _24553_, _24554_);
  or g_55568_(_24544_, _24554_, _24555_);
  xor g_55569_(out[119], out[359], _24556_);
  and g_55570_(_39581_, out[363], _24557_);
  xor g_55571_(out[126], out[366], _24558_);
  xor g_55572_(out[120], out[360], _24559_);
  xor g_55573_(out[113], out[353], _24560_);
  xor g_55574_(out[125], out[365], _24561_);
  xor g_55575_(out[121], out[361], _24563_);
  xor g_55576_(out[116], out[356], _24564_);
  xor g_55577_(out[114], out[354], _24565_);
  and g_55578_(out[123], _39746_, _24566_);
  xor g_55579_(out[115], out[355], _24567_);
  xor g_55580_(out[118], out[358], _24568_);
  xor g_55581_(out[127], out[367], _24569_);
  xor g_55582_(out[122], out[362], _24570_);
  xor g_55583_(out[117], out[357], _24571_);
  xor g_55584_(out[112], out[352], _24572_);
  or g_55585_(_24558_, _24564_, _24574_);
  or g_55586_(_24559_, _24561_, _24575_);
  or g_55587_(_24565_, _24570_, _24576_);
  or g_55588_(_24575_, _24576_, _24577_);
  or g_55589_(_24563_, _24567_, _24578_);
  or g_55590_(_24571_, _24572_, _24579_);
  or g_55591_(_24578_, _24579_, _24580_);
  or g_55592_(_24577_, _24580_, _24581_);
  xor g_55593_(out[124], out[364], _24582_);
  or g_55594_(_24557_, _24582_, _24583_);
  or g_55595_(_24556_, _24568_, _24585_);
  or g_55596_(_24583_, _24585_, _24586_);
  or g_55597_(_24560_, _24566_, _24587_);
  or g_55598_(_24569_, _24587_, _24588_);
  or g_55599_(_24586_, _24588_, _24589_);
  or g_55600_(_24581_, _24589_, _24590_);
  or g_55601_(_24574_, _24590_, _24591_);
  xor g_55602_(out[97], out[353], _24592_);
  and g_55603_(out[107], _39746_, _24593_);
  xor g_55604_(out[105], out[361], _24594_);
  xor g_55605_(out[96], out[352], _24596_);
  xor g_55606_(out[110], out[366], _24597_);
  xor g_55607_(out[100], out[356], _24598_);
  or g_55608_(_24597_, _24598_, _24599_);
  xor g_55609_(out[109], out[365], _24600_);
  xor g_55610_(out[99], out[355], _24601_);
  and g_55611_(_39570_, out[363], _24602_);
  xor g_55612_(out[102], out[358], _24603_);
  xor g_55613_(out[106], out[362], _24604_);
  xor g_55614_(out[101], out[357], _24605_);
  xor g_55615_(out[111], out[367], _24607_);
  xor g_55616_(out[104], out[360], _24608_);
  or g_55617_(_24600_, _24608_, _24609_);
  xor g_55618_(out[98], out[354], _24610_);
  or g_55619_(_24604_, _24610_, _24611_);
  or g_55620_(_24609_, _24611_, _24612_);
  or g_55621_(_24594_, _24601_, _24613_);
  or g_55622_(_24605_, _24613_, _24614_);
  or g_55623_(_24612_, _24614_, _24615_);
  or g_55624_(_24599_, _24615_, _24616_);
  xor g_55625_(out[108], out[364], _24618_);
  or g_55626_(_24602_, _24618_, _24619_);
  xor g_55627_(out[103], out[359], _24620_);
  or g_55628_(_24603_, _24620_, _24621_);
  or g_55629_(_24619_, _24621_, _24622_);
  or g_55630_(_24592_, _24593_, _24623_);
  or g_55631_(_24607_, _24623_, _24624_);
  or g_55632_(_24622_, _24624_, _24625_);
  or g_55633_(_24596_, _24625_, _24626_);
  or g_55634_(_24616_, _24626_, _24627_);
  xor g_55635_(out[87], out[359], _24629_);
  and g_55636_(_39559_, out[363], _24630_);
  xor g_55637_(out[94], out[366], _24631_);
  xor g_55638_(out[88], out[360], _24632_);
  xor g_55639_(out[81], out[353], _24633_);
  xor g_55640_(out[93], out[365], _24634_);
  xor g_55641_(out[89], out[361], _24635_);
  xor g_55642_(out[84], out[356], _24636_);
  xor g_55643_(out[82], out[354], _24637_);
  and g_55644_(out[91], _39746_, _24638_);
  xor g_55645_(out[83], out[355], _24640_);
  xor g_55646_(out[86], out[358], _24641_);
  xor g_55647_(out[95], out[367], _24642_);
  xor g_55648_(out[90], out[362], _24643_);
  xor g_55649_(out[85], out[357], _24644_);
  xor g_55650_(out[80], out[352], _24645_);
  or g_55651_(_24631_, _24636_, _24646_);
  or g_55652_(_24632_, _24634_, _24647_);
  or g_55653_(_24637_, _24643_, _24648_);
  or g_55654_(_24647_, _24648_, _24649_);
  or g_55655_(_24635_, _24640_, _24651_);
  or g_55656_(_24644_, _24645_, _24652_);
  or g_55657_(_24651_, _24652_, _24653_);
  or g_55658_(_24649_, _24653_, _24654_);
  xor g_55659_(out[92], out[364], _24655_);
  or g_55660_(_24630_, _24655_, _24656_);
  or g_55661_(_24629_, _24641_, _24657_);
  or g_55662_(_24656_, _24657_, _24658_);
  or g_55663_(_24633_, _24638_, _24659_);
  or g_55664_(_24642_, _24659_, _24660_);
  or g_55665_(_24658_, _24660_, _24662_);
  or g_55666_(_24654_, _24662_, _24663_);
  or g_55667_(_24646_, _24663_, _24664_);
  xor g_55668_(out[65], out[353], _24665_);
  and g_55669_(out[75], _39746_, _24666_);
  xor g_55670_(out[73], out[361], _24667_);
  xor g_55671_(out[64], out[352], _24668_);
  xor g_55672_(out[78], out[366], _24669_);
  xor g_55673_(out[68], out[356], _24670_);
  or g_55674_(_24669_, _24670_, _24671_);
  xor g_55675_(out[77], out[365], _24673_);
  xor g_55676_(out[67], out[355], _24674_);
  and g_55677_(_39548_, out[363], _24675_);
  xor g_55678_(out[70], out[358], _24676_);
  xor g_55679_(out[74], out[362], _24677_);
  xor g_55680_(out[69], out[357], _24678_);
  xor g_55681_(out[79], out[367], _24679_);
  xor g_55682_(out[72], out[360], _24680_);
  or g_55683_(_24673_, _24680_, _24681_);
  xor g_55684_(out[66], out[354], _24682_);
  or g_55685_(_24677_, _24682_, _24684_);
  or g_55686_(_24681_, _24684_, _24685_);
  or g_55687_(_24667_, _24674_, _24686_);
  or g_55688_(_24678_, _24686_, _24687_);
  or g_55689_(_24685_, _24687_, _24688_);
  or g_55690_(_24671_, _24688_, _24689_);
  xor g_55691_(out[76], out[364], _24690_);
  or g_55692_(_24675_, _24690_, _24691_);
  xor g_55693_(out[71], out[359], _24692_);
  or g_55694_(_24676_, _24692_, _24693_);
  or g_55695_(_24691_, _24693_, _24695_);
  or g_55696_(_24665_, _24666_, _24696_);
  or g_55697_(_24679_, _24696_, _24697_);
  or g_55698_(_24695_, _24697_, _24698_);
  or g_55699_(_24668_, _24698_, _24699_);
  or g_55700_(_24689_, _24699_, _24700_);
  xor g_55701_(out[55], out[359], _24701_);
  and g_55702_(_39537_, out[363], _24702_);
  xor g_55703_(out[62], out[366], _24703_);
  xor g_55704_(out[56], out[360], _24704_);
  xor g_55705_(out[49], out[353], _24706_);
  xor g_55706_(out[61], out[365], _24707_);
  xor g_55707_(out[57], out[361], _24708_);
  xor g_55708_(out[52], out[356], _24709_);
  xor g_55709_(out[50], out[354], _24710_);
  and g_55710_(out[59], _39746_, _24711_);
  xor g_55711_(out[51], out[355], _24712_);
  xor g_55712_(out[54], out[358], _24713_);
  xor g_55713_(out[63], out[367], _24714_);
  xor g_55714_(out[58], out[362], _24715_);
  xor g_55715_(out[53], out[357], _24717_);
  xor g_55716_(out[48], out[352], _24718_);
  or g_55717_(_24703_, _24709_, _24719_);
  or g_55718_(_24704_, _24707_, _24720_);
  or g_55719_(_24710_, _24715_, _24721_);
  or g_55720_(_24720_, _24721_, _24722_);
  or g_55721_(_24708_, _24712_, _24723_);
  or g_55722_(_24717_, _24718_, _24724_);
  or g_55723_(_24723_, _24724_, _24725_);
  or g_55724_(_24722_, _24725_, _24726_);
  xor g_55725_(out[60], out[364], _24728_);
  or g_55726_(_24702_, _24728_, _24729_);
  or g_55727_(_24701_, _24713_, _24730_);
  or g_55728_(_24729_, _24730_, _24731_);
  or g_55729_(_24706_, _24711_, _24732_);
  or g_55730_(_24714_, _24732_, _24733_);
  or g_55731_(_24731_, _24733_, _24734_);
  or g_55732_(_24726_, _24734_, _24735_);
  or g_55733_(_24719_, _24735_, _24736_);
  not g_55734_(_24736_, _24737_);
  xor g_55735_(out[33], out[353], _24739_);
  and g_55736_(out[43], _39746_, _24740_);
  xor g_55737_(out[41], out[361], _24741_);
  xor g_55738_(out[32], out[352], _24742_);
  xor g_55739_(out[46], out[366], _24743_);
  xor g_55740_(out[36], out[356], _24744_);
  or g_55741_(_24743_, _24744_, _24745_);
  xor g_55742_(out[45], out[365], _24746_);
  xor g_55743_(out[35], out[355], _24747_);
  and g_55744_(_39526_, out[363], _24748_);
  xor g_55745_(out[38], out[358], _24750_);
  xor g_55746_(out[42], out[362], _24751_);
  xor g_55747_(out[37], out[357], _24752_);
  xor g_55748_(out[47], out[367], _24753_);
  xor g_55749_(out[40], out[360], _24754_);
  or g_55750_(_24746_, _24754_, _24755_);
  xor g_55751_(out[34], out[354], _24756_);
  or g_55752_(_24751_, _24756_, _24757_);
  or g_55753_(_24755_, _24757_, _24758_);
  or g_55754_(_24741_, _24747_, _24759_);
  or g_55755_(_24752_, _24759_, _24761_);
  or g_55756_(_24758_, _24761_, _24762_);
  or g_55757_(_24745_, _24762_, _24763_);
  xor g_55758_(out[44], out[364], _24764_);
  or g_55759_(_24748_, _24764_, _24765_);
  xor g_55760_(out[39], out[359], _24766_);
  or g_55761_(_24750_, _24766_, _24767_);
  or g_55762_(_24765_, _24767_, _24768_);
  or g_55763_(_24739_, _24740_, _24769_);
  or g_55764_(_24753_, _24769_, _24770_);
  or g_55765_(_24768_, _24770_, _24772_);
  or g_55766_(_24742_, _24772_, _24773_);
  or g_55767_(_24763_, _24773_, _24774_);
  xor g_55768_(out[23], out[359], _24775_);
  and g_55769_(_39493_, out[363], _24776_);
  xor g_55770_(out[30], out[366], _24777_);
  xor g_55771_(out[24], out[360], _24778_);
  xor g_55772_(out[17], out[353], _24779_);
  xor g_55773_(out[29], out[365], _24780_);
  xor g_55774_(out[25], out[361], _24781_);
  xor g_55775_(out[20], out[356], _24783_);
  xor g_55776_(out[18], out[354], _24784_);
  and g_55777_(out[27], _39746_, _24785_);
  xor g_55778_(out[19], out[355], _24786_);
  xor g_55779_(out[22], out[358], _24787_);
  xor g_55780_(out[31], out[367], _24788_);
  xor g_55781_(out[26], out[362], _24789_);
  xor g_55782_(out[21], out[357], _24790_);
  xor g_55783_(out[16], out[352], _24791_);
  or g_55784_(_24777_, _24783_, _24792_);
  or g_55785_(_24778_, _24780_, _24794_);
  or g_55786_(_24784_, _24789_, _24795_);
  or g_55787_(_24794_, _24795_, _24796_);
  or g_55788_(_24781_, _24786_, _24797_);
  or g_55789_(_24790_, _24791_, _24798_);
  or g_55790_(_24797_, _24798_, _24799_);
  or g_55791_(_24796_, _24799_, _24800_);
  xor g_55792_(out[28], out[364], _24801_);
  or g_55793_(_24776_, _24801_, _24802_);
  or g_55794_(_24775_, _24787_, _24803_);
  or g_55795_(_24802_, _24803_, _24805_);
  or g_55796_(_24779_, _24785_, _24806_);
  or g_55797_(_24788_, _24806_, _24807_);
  or g_55798_(_24805_, _24807_, _24808_);
  or g_55799_(_24800_, _24808_, _24809_);
  or g_55800_(_24792_, _24809_, _24810_);
  and g_55801_(_39438_, out[363], _24811_);
  and g_55802_(out[11], _39746_, _24812_);
  xor g_55803_(out[2], out[354], _24813_);
  xor g_55804_(out[9], out[361], _24814_);
  xor g_55805_(out[8], out[360], _24816_);
  xor g_55806_(out[1], out[353], _24817_);
  xor g_55807_(out[5], out[357], _24818_);
  xor g_55808_(out[0], out[352], _24819_);
  xor g_55809_(out[6], out[358], _24820_);
  xor g_55810_(out[15], out[367], _24821_);
  xor g_55811_(out[10], out[362], _24822_);
  xor g_55812_(out[3], out[355], _24823_);
  xor g_55813_(out[14], out[366], _24824_);
  xor g_55814_(out[4], out[356], _24825_);
  xor g_55815_(out[13], out[365], _24827_);
  or g_55816_(_24816_, _24827_, _24828_);
  or g_55817_(_24813_, _24822_, _24829_);
  or g_55818_(_24828_, _24829_, _24830_);
  or g_55819_(_24814_, _24823_, _24831_);
  or g_55820_(_24818_, _24831_, _24832_);
  or g_55821_(_24830_, _24832_, _24833_);
  or g_55822_(_24824_, _24825_, _24834_);
  or g_55823_(_24833_, _24834_, _24835_);
  xor g_55824_(out[12], out[364], _24836_);
  or g_55825_(_24811_, _24836_, _24838_);
  xor g_55826_(out[7], out[359], _24839_);
  or g_55827_(_24820_, _24839_, _24840_);
  or g_55828_(_24838_, _24840_, _24841_);
  or g_55829_(_24812_, _24817_, _24842_);
  or g_55830_(_24821_, _24842_, _24843_);
  or g_55831_(_24841_, _24843_, _24844_);
  or g_55832_(_24819_, _24844_, _24845_);
  or g_55833_(_24835_, _24845_, _24846_);
  not g_55834_(_24846_, _24847_);
  xor g_55835_(out[305], out[337], _24849_);
  and g_55836_(out[315], _39735_, _24850_);
  xor g_55837_(out[313], out[345], _24851_);
  xor g_55838_(out[304], out[336], _24852_);
  xor g_55839_(out[318], out[350], _24853_);
  xor g_55840_(out[308], out[340], _24854_);
  or g_55841_(_24853_, _24854_, _24855_);
  xor g_55842_(out[317], out[349], _24856_);
  xor g_55843_(out[307], out[339], _24857_);
  and g_55844_(_39724_, out[347], _24858_);
  xor g_55845_(out[310], out[342], _24860_);
  xor g_55846_(out[314], out[346], _24861_);
  xor g_55847_(out[309], out[341], _24862_);
  xor g_55848_(out[319], out[351], _24863_);
  xor g_55849_(out[312], out[344], _24864_);
  or g_55850_(_24856_, _24864_, _24865_);
  xor g_55851_(out[306], out[338], _24866_);
  or g_55852_(_24861_, _24866_, _24867_);
  or g_55853_(_24865_, _24867_, _24868_);
  or g_55854_(_24851_, _24857_, _24869_);
  or g_55855_(_24862_, _24869_, _24871_);
  or g_55856_(_24868_, _24871_, _24872_);
  or g_55857_(_24855_, _24872_, _24873_);
  xor g_55858_(out[316], out[348], _24874_);
  or g_55859_(_24858_, _24874_, _24875_);
  xor g_55860_(out[311], out[343], _24876_);
  or g_55861_(_24860_, _24876_, _24877_);
  or g_55862_(_24875_, _24877_, _24878_);
  or g_55863_(_24849_, _24850_, _24879_);
  or g_55864_(_24863_, _24879_, _24880_);
  or g_55865_(_24878_, _24880_, _24882_);
  or g_55866_(_24852_, _24882_, _24883_);
  or g_55867_(_24873_, _24883_, _24884_);
  xor g_55868_(out[295], out[343], _24885_);
  and g_55869_(_39702_, out[347], _24886_);
  xor g_55870_(out[302], out[350], _24887_);
  xor g_55871_(out[296], out[344], _24888_);
  xor g_55872_(out[289], out[337], _24889_);
  xor g_55873_(out[301], out[349], _24890_);
  xor g_55874_(out[297], out[345], _24891_);
  xor g_55875_(out[292], out[340], _24893_);
  xor g_55876_(out[290], out[338], _24894_);
  and g_55877_(out[299], _39735_, _24895_);
  xor g_55878_(out[291], out[339], _24896_);
  xor g_55879_(out[294], out[342], _24897_);
  xor g_55880_(out[303], out[351], _24898_);
  xor g_55881_(out[298], out[346], _24899_);
  xor g_55882_(out[293], out[341], _24900_);
  xor g_55883_(out[288], out[336], _24901_);
  or g_55884_(_24887_, _24893_, _24902_);
  or g_55885_(_24888_, _24890_, _24904_);
  or g_55886_(_24894_, _24899_, _24905_);
  or g_55887_(_24904_, _24905_, _24906_);
  or g_55888_(_24891_, _24896_, _24907_);
  or g_55889_(_24900_, _24901_, _24908_);
  or g_55890_(_24907_, _24908_, _24909_);
  or g_55891_(_24906_, _24909_, _24910_);
  xor g_55892_(out[300], out[348], _24911_);
  or g_55893_(_24886_, _24911_, _24912_);
  or g_55894_(_24885_, _24897_, _24913_);
  or g_55895_(_24912_, _24913_, _24915_);
  or g_55896_(_24889_, _24895_, _24916_);
  or g_55897_(_24898_, _24916_, _24917_);
  or g_55898_(_24915_, _24917_, _24918_);
  or g_55899_(_24910_, _24918_, _24919_);
  or g_55900_(_24902_, _24919_, _24920_);
  not g_55901_(_24920_, _24921_);
  xor g_55902_(out[273], out[337], _24922_);
  and g_55903_(out[283], _39735_, _24923_);
  xor g_55904_(out[281], out[345], _24924_);
  xor g_55905_(out[272], out[336], _24926_);
  xor g_55906_(out[286], out[350], _24927_);
  xor g_55907_(out[276], out[340], _24928_);
  or g_55908_(_24927_, _24928_, _24929_);
  xor g_55909_(out[285], out[349], _24930_);
  xor g_55910_(out[275], out[339], _24931_);
  and g_55911_(_39691_, out[347], _24932_);
  xor g_55912_(out[278], out[342], _24933_);
  xor g_55913_(out[282], out[346], _24934_);
  xor g_55914_(out[277], out[341], _24935_);
  xor g_55915_(out[287], out[351], _24937_);
  xor g_55916_(out[280], out[344], _24938_);
  or g_55917_(_24930_, _24938_, _24939_);
  xor g_55918_(out[274], out[338], _24940_);
  or g_55919_(_24934_, _24940_, _24941_);
  or g_55920_(_24939_, _24941_, _24942_);
  or g_55921_(_24924_, _24931_, _24943_);
  or g_55922_(_24935_, _24943_, _24944_);
  or g_55923_(_24942_, _24944_, _24945_);
  or g_55924_(_24929_, _24945_, _24946_);
  xor g_55925_(out[284], out[348], _24948_);
  or g_55926_(_24932_, _24948_, _24949_);
  xor g_55927_(out[279], out[343], _24950_);
  or g_55928_(_24933_, _24950_, _24951_);
  or g_55929_(_24949_, _24951_, _24952_);
  or g_55930_(_24922_, _24923_, _24953_);
  or g_55931_(_24937_, _24953_, _24954_);
  or g_55932_(_24952_, _24954_, _24955_);
  or g_55933_(_24926_, _24955_, _24956_);
  or g_55934_(_24946_, _24956_, _24957_);
  xor g_55935_(out[263], out[343], _24959_);
  and g_55936_(_39680_, out[347], _24960_);
  xor g_55937_(out[270], out[350], _24961_);
  xor g_55938_(out[264], out[344], _24962_);
  xor g_55939_(out[257], out[337], _24963_);
  xor g_55940_(out[269], out[349], _24964_);
  xor g_55941_(out[265], out[345], _24965_);
  xor g_55942_(out[260], out[340], _24966_);
  xor g_55943_(out[258], out[338], _24967_);
  and g_55944_(out[267], _39735_, _24968_);
  xor g_55945_(out[259], out[339], _24970_);
  xor g_55946_(out[262], out[342], _24971_);
  xor g_55947_(out[271], out[351], _24972_);
  xor g_55948_(out[266], out[346], _24973_);
  xor g_55949_(out[261], out[341], _24974_);
  xor g_55950_(out[256], out[336], _24975_);
  or g_55951_(_24961_, _24966_, _24976_);
  or g_55952_(_24962_, _24964_, _24977_);
  or g_55953_(_24967_, _24973_, _24978_);
  or g_55954_(_24977_, _24978_, _24979_);
  or g_55955_(_24965_, _24970_, _24981_);
  or g_55956_(_24974_, _24975_, _24982_);
  or g_55957_(_24981_, _24982_, _24983_);
  or g_55958_(_24979_, _24983_, _24984_);
  xor g_55959_(out[268], out[348], _24985_);
  or g_55960_(_24960_, _24985_, _24986_);
  or g_55961_(_24959_, _24971_, _24987_);
  or g_55962_(_24986_, _24987_, _24988_);
  or g_55963_(_24963_, _24968_, _24989_);
  or g_55964_(_24972_, _24989_, _24990_);
  or g_55965_(_24988_, _24990_, _24992_);
  or g_55966_(_24984_, _24992_, _24993_);
  or g_55967_(_24976_, _24993_, _24994_);
  xor g_55968_(out[241], out[337], _24995_);
  and g_55969_(out[251], _39735_, _24996_);
  xor g_55970_(out[254], out[350], _24997_);
  xor g_55971_(out[243], out[339], _24998_);
  xor g_55972_(out[244], out[340], _24999_);
  xor g_55973_(out[242], out[338], _25000_);
  xor g_55974_(out[249], out[345], _25001_);
  xor g_55975_(out[240], out[336], _25003_);
  and g_55976_(_39669_, out[347], _25004_);
  xor g_55977_(out[246], out[342], _25005_);
  xor g_55978_(out[250], out[346], _25006_);
  xor g_55979_(out[245], out[341], _25007_);
  xor g_55980_(out[255], out[351], _25008_);
  xor g_55981_(out[253], out[349], _25009_);
  xor g_55982_(out[248], out[344], _25010_);
  or g_55983_(_24997_, _24999_, _25011_);
  or g_55984_(_25009_, _25010_, _25012_);
  or g_55985_(_25000_, _25006_, _25014_);
  or g_55986_(_25012_, _25014_, _25015_);
  or g_55987_(_24998_, _25001_, _25016_);
  or g_55988_(_25003_, _25007_, _25017_);
  or g_55989_(_25016_, _25017_, _25018_);
  or g_55990_(_25015_, _25018_, _25019_);
  xor g_55991_(out[252], out[348], _25020_);
  or g_55992_(_25004_, _25020_, _25021_);
  xor g_55993_(out[247], out[343], _25022_);
  or g_55994_(_25005_, _25022_, _25023_);
  or g_55995_(_25021_, _25023_, _25025_);
  or g_55996_(_24995_, _24996_, _25026_);
  or g_55997_(_25008_, _25026_, _25027_);
  or g_55998_(_25025_, _25027_, _25028_);
  or g_55999_(_25019_, _25028_, _25029_);
  or g_56000_(_25011_, _25029_, _25030_);
  xor g_56001_(out[231], out[343], _25031_);
  and g_56002_(_39658_, out[347], _25032_);
  xor g_56003_(out[238], out[350], _25033_);
  xor g_56004_(out[232], out[344], _25034_);
  xor g_56005_(out[225], out[337], _25036_);
  xor g_56006_(out[237], out[349], _25037_);
  xor g_56007_(out[233], out[345], _25038_);
  xor g_56008_(out[228], out[340], _25039_);
  xor g_56009_(out[226], out[338], _25040_);
  and g_56010_(out[235], _39735_, _25041_);
  xor g_56011_(out[227], out[339], _25042_);
  xor g_56012_(out[230], out[342], _25043_);
  xor g_56013_(out[239], out[351], _25044_);
  xor g_56014_(out[234], out[346], _25045_);
  xor g_56015_(out[229], out[341], _25047_);
  xor g_56016_(out[224], out[336], _25048_);
  or g_56017_(_25033_, _25039_, _25049_);
  or g_56018_(_25034_, _25037_, _25050_);
  or g_56019_(_25040_, _25045_, _25051_);
  or g_56020_(_25050_, _25051_, _25052_);
  or g_56021_(_25038_, _25042_, _25053_);
  or g_56022_(_25047_, _25048_, _25054_);
  or g_56023_(_25053_, _25054_, _25055_);
  or g_56024_(_25052_, _25055_, _25056_);
  xor g_56025_(out[236], out[348], _25058_);
  or g_56026_(_25032_, _25058_, _25059_);
  or g_56027_(_25031_, _25043_, _25060_);
  or g_56028_(_25059_, _25060_, _25061_);
  or g_56029_(_25036_, _25041_, _25062_);
  or g_56030_(_25044_, _25062_, _25063_);
  or g_56031_(_25061_, _25063_, _25064_);
  or g_56032_(_25056_, _25064_, _25065_);
  or g_56033_(_25049_, _25065_, _25066_);
  and g_56034_(out[219], _39735_, _25067_);
  and g_56035_(_39647_, out[347], _25069_);
  xor g_56036_(out[216], out[344], _25070_);
  xor g_56037_(out[223], out[351], _25071_);
  xor g_56038_(out[209], out[337], _25072_);
  xor g_56039_(out[210], out[338], _25073_);
  xor g_56040_(out[212], out[340], _25074_);
  xor g_56041_(out[221], out[349], _25075_);
  xor g_56042_(out[217], out[345], _25076_);
  xor g_56043_(out[211], out[339], _25077_);
  xor g_56044_(out[213], out[341], _25078_);
  xor g_56045_(out[222], out[350], _25080_);
  xor g_56046_(out[208], out[336], _25081_);
  xor g_56047_(out[218], out[346], _25082_);
  or g_56048_(_25070_, _25075_, _25083_);
  xor g_56049_(out[214], out[342], _25084_);
  or g_56050_(_25073_, _25082_, _25085_);
  or g_56051_(_25083_, _25085_, _25086_);
  or g_56052_(_25076_, _25077_, _25087_);
  or g_56053_(_25078_, _25087_, _25088_);
  or g_56054_(_25086_, _25088_, _25089_);
  or g_56055_(_25074_, _25080_, _25091_);
  or g_56056_(_25089_, _25091_, _25092_);
  xor g_56057_(out[220], out[348], _25093_);
  or g_56058_(_25069_, _25093_, _25094_);
  xor g_56059_(out[215], out[343], _25095_);
  or g_56060_(_25084_, _25095_, _25096_);
  or g_56061_(_25094_, _25096_, _25097_);
  or g_56062_(_25067_, _25072_, _25098_);
  or g_56063_(_25071_, _25098_, _25099_);
  or g_56064_(_25097_, _25099_, _25100_);
  or g_56065_(_25081_, _25100_, _25102_);
  or g_56066_(_25092_, _25102_, _25103_);
  not g_56067_(_25103_, _25104_);
  xor g_56068_(out[199], out[343], _25105_);
  and g_56069_(_39636_, out[347], _25106_);
  xor g_56070_(out[206], out[350], _25107_);
  xor g_56071_(out[200], out[344], _25108_);
  xor g_56072_(out[193], out[337], _25109_);
  xor g_56073_(out[205], out[349], _25110_);
  xor g_56074_(out[201], out[345], _25111_);
  xor g_56075_(out[196], out[340], _25113_);
  xor g_56076_(out[194], out[338], _25114_);
  and g_56077_(out[203], _39735_, _25115_);
  xor g_56078_(out[195], out[339], _25116_);
  xor g_56079_(out[198], out[342], _25117_);
  xor g_56080_(out[207], out[351], _25118_);
  xor g_56081_(out[202], out[346], _25119_);
  xor g_56082_(out[197], out[341], _25120_);
  xor g_56083_(out[192], out[336], _25121_);
  or g_56084_(_25107_, _25113_, _25122_);
  or g_56085_(_25108_, _25110_, _25124_);
  or g_56086_(_25114_, _25119_, _25125_);
  or g_56087_(_25124_, _25125_, _25126_);
  or g_56088_(_25111_, _25116_, _25127_);
  or g_56089_(_25120_, _25121_, _25128_);
  or g_56090_(_25127_, _25128_, _25129_);
  or g_56091_(_25126_, _25129_, _25130_);
  xor g_56092_(out[204], out[348], _25131_);
  or g_56093_(_25106_, _25131_, _25132_);
  or g_56094_(_25105_, _25117_, _25133_);
  or g_56095_(_25132_, _25133_, _25135_);
  or g_56096_(_25109_, _25115_, _25136_);
  or g_56097_(_25118_, _25136_, _25137_);
  or g_56098_(_25135_, _25137_, _25138_);
  or g_56099_(_25130_, _25138_, _25139_);
  or g_56100_(_25122_, _25139_, _25140_);
  not g_56101_(_25140_, _25141_);
  xor g_56102_(out[177], out[337], _25142_);
  and g_56103_(out[187], _39735_, _25143_);
  xor g_56104_(out[185], out[345], _25144_);
  xor g_56105_(out[176], out[336], _25146_);
  xor g_56106_(out[190], out[350], _25147_);
  xor g_56107_(out[180], out[340], _25148_);
  or g_56108_(_25147_, _25148_, _25149_);
  xor g_56109_(out[189], out[349], _25150_);
  xor g_56110_(out[179], out[339], _25151_);
  and g_56111_(_39625_, out[347], _25152_);
  xor g_56112_(out[182], out[342], _25153_);
  xor g_56113_(out[186], out[346], _25154_);
  xor g_56114_(out[181], out[341], _25155_);
  xor g_56115_(out[191], out[351], _25157_);
  xor g_56116_(out[184], out[344], _25158_);
  or g_56117_(_25150_, _25158_, _25159_);
  xor g_56118_(out[178], out[338], _25160_);
  or g_56119_(_25154_, _25160_, _25161_);
  or g_56120_(_25159_, _25161_, _25162_);
  or g_56121_(_25144_, _25151_, _25163_);
  or g_56122_(_25155_, _25163_, _25164_);
  or g_56123_(_25162_, _25164_, _25165_);
  or g_56124_(_25149_, _25165_, _25166_);
  xor g_56125_(out[188], out[348], _25168_);
  or g_56126_(_25152_, _25168_, _25169_);
  xor g_56127_(out[183], out[343], _25170_);
  or g_56128_(_25153_, _25170_, _25171_);
  or g_56129_(_25169_, _25171_, _25172_);
  or g_56130_(_25142_, _25143_, _25173_);
  or g_56131_(_25157_, _25173_, _25174_);
  or g_56132_(_25172_, _25174_, _25175_);
  or g_56133_(_25146_, _25175_, _25176_);
  or g_56134_(_25166_, _25176_, _25177_);
  xor g_56135_(out[167], out[343], _25179_);
  and g_56136_(_39614_, out[347], _25180_);
  xor g_56137_(out[174], out[350], _25181_);
  xor g_56138_(out[168], out[344], _25182_);
  xor g_56139_(out[161], out[337], _25183_);
  xor g_56140_(out[173], out[349], _25184_);
  xor g_56141_(out[169], out[345], _25185_);
  xor g_56142_(out[164], out[340], _25186_);
  xor g_56143_(out[162], out[338], _25187_);
  and g_56144_(out[171], _39735_, _25188_);
  xor g_56145_(out[163], out[339], _25190_);
  xor g_56146_(out[166], out[342], _25191_);
  xor g_56147_(out[175], out[351], _25192_);
  xor g_56148_(out[170], out[346], _25193_);
  xor g_56149_(out[165], out[341], _25194_);
  xor g_56150_(out[160], out[336], _25195_);
  or g_56151_(_25181_, _25186_, _25196_);
  or g_56152_(_25182_, _25184_, _25197_);
  or g_56153_(_25187_, _25193_, _25198_);
  or g_56154_(_25197_, _25198_, _25199_);
  or g_56155_(_25185_, _25190_, _25201_);
  or g_56156_(_25194_, _25195_, _25202_);
  or g_56157_(_25201_, _25202_, _25203_);
  or g_56158_(_25199_, _25203_, _25204_);
  xor g_56159_(out[172], out[348], _25205_);
  or g_56160_(_25180_, _25205_, _25206_);
  or g_56161_(_25179_, _25191_, _25207_);
  or g_56162_(_25206_, _25207_, _25208_);
  or g_56163_(_25183_, _25188_, _25209_);
  or g_56164_(_25192_, _25209_, _25210_);
  or g_56165_(_25208_, _25210_, _25212_);
  or g_56166_(_25204_, _25212_, _25213_);
  or g_56167_(_25196_, _25213_, _25214_);
  xor g_56168_(out[157], out[349], _25215_);
  xor g_56169_(out[146], out[338], _25216_);
  xor g_56170_(out[149], out[341], _25217_);
  xor g_56171_(out[153], out[345], _25218_);
  xor g_56172_(out[148], out[340], _25219_);
  xor g_56173_(out[152], out[344], _25220_);
  xor g_56174_(out[158], out[350], _25221_);
  xor g_56175_(out[150], out[342], _25223_);
  xor g_56176_(out[159], out[351], _25224_);
  xor g_56177_(out[154], out[346], _25225_);
  xor g_56178_(out[144], out[336], _25226_);
  xor g_56179_(out[147], out[339], _25227_);
  and g_56180_(_39603_, out[347], _25228_);
  and g_56181_(out[155], _39735_, _25229_);
  xor g_56182_(out[145], out[337], _25230_);
  or g_56183_(_25219_, _25221_, _25231_);
  or g_56184_(_25215_, _25220_, _25232_);
  or g_56185_(_25216_, _25225_, _25234_);
  or g_56186_(_25232_, _25234_, _25235_);
  or g_56187_(_25218_, _25227_, _25236_);
  or g_56188_(_25217_, _25226_, _25237_);
  or g_56189_(_25236_, _25237_, _25238_);
  or g_56190_(_25235_, _25238_, _25239_);
  xor g_56191_(out[156], out[348], _25240_);
  or g_56192_(_25228_, _25240_, _25241_);
  xor g_56193_(out[151], out[343], _25242_);
  or g_56194_(_25223_, _25242_, _25243_);
  or g_56195_(_25241_, _25243_, _25245_);
  or g_56196_(_25229_, _25230_, _25246_);
  or g_56197_(_25224_, _25246_, _25247_);
  or g_56198_(_25245_, _25247_, _25248_);
  or g_56199_(_25239_, _25248_, _25249_);
  or g_56200_(_25231_, _25249_, _25250_);
  not g_56201_(_25250_, _25251_);
  xor g_56202_(out[135], out[343], _25252_);
  and g_56203_(_39592_, out[347], _25253_);
  xor g_56204_(out[142], out[350], _25254_);
  xor g_56205_(out[136], out[344], _25256_);
  xor g_56206_(out[129], out[337], _25257_);
  xor g_56207_(out[141], out[349], _25258_);
  xor g_56208_(out[137], out[345], _25259_);
  xor g_56209_(out[132], out[340], _25260_);
  xor g_56210_(out[130], out[338], _25261_);
  and g_56211_(out[139], _39735_, _25262_);
  xor g_56212_(out[131], out[339], _25263_);
  xor g_56213_(out[134], out[342], _25264_);
  xor g_56214_(out[143], out[351], _25265_);
  xor g_56215_(out[138], out[346], _25267_);
  xor g_56216_(out[133], out[341], _25268_);
  xor g_56217_(out[128], out[336], _25269_);
  or g_56218_(_25254_, _25260_, _25270_);
  or g_56219_(_25256_, _25258_, _25271_);
  or g_56220_(_25261_, _25267_, _25272_);
  or g_56221_(_25271_, _25272_, _25273_);
  or g_56222_(_25259_, _25263_, _25274_);
  or g_56223_(_25268_, _25269_, _25275_);
  or g_56224_(_25274_, _25275_, _25276_);
  or g_56225_(_25273_, _25276_, _25278_);
  xor g_56226_(out[140], out[348], _25279_);
  or g_56227_(_25253_, _25279_, _25280_);
  or g_56228_(_25252_, _25264_, _25281_);
  or g_56229_(_25280_, _25281_, _25282_);
  or g_56230_(_25257_, _25262_, _25283_);
  or g_56231_(_25265_, _25283_, _25284_);
  or g_56232_(_25282_, _25284_, _25285_);
  or g_56233_(_25278_, _25285_, _25286_);
  or g_56234_(_25270_, _25286_, _25287_);
  xor g_56235_(out[124], out[348], _25289_);
  and g_56236_(_39581_, out[347], _25290_);
  xor g_56237_(out[120], out[344], _25291_);
  xor g_56238_(out[118], out[342], _25292_);
  xor g_56239_(out[125], out[349], _25293_);
  xor g_56240_(out[126], out[350], _25294_);
  xor g_56241_(out[114], out[338], _25295_);
  xor g_56242_(out[121], out[345], _25296_);
  xor g_56243_(out[117], out[341], _25297_);
  xor g_56244_(out[113], out[337], _25298_);
  and g_56245_(out[123], _39735_, _25300_);
  or g_56246_(_25291_, _25293_, _25301_);
  xor g_56247_(out[127], out[351], _25302_);
  xor g_56248_(out[122], out[346], _25303_);
  xor g_56249_(out[116], out[340], _25304_);
  xor g_56250_(out[115], out[339], _25305_);
  xor g_56251_(out[112], out[336], _25306_);
  or g_56252_(_25295_, _25303_, _25307_);
  or g_56253_(_25301_, _25307_, _25308_);
  or g_56254_(_25296_, _25305_, _25309_);
  or g_56255_(_25297_, _25309_, _25311_);
  or g_56256_(_25308_, _25311_, _25312_);
  or g_56257_(_25294_, _25304_, _25313_);
  or g_56258_(_25312_, _25313_, _25314_);
  or g_56259_(_25289_, _25290_, _25315_);
  xor g_56260_(out[119], out[343], _25316_);
  or g_56261_(_25292_, _25316_, _25317_);
  or g_56262_(_25315_, _25317_, _25318_);
  or g_56263_(_25298_, _25300_, _25319_);
  or g_56264_(_25302_, _25319_, _25320_);
  or g_56265_(_25318_, _25320_, _25322_);
  or g_56266_(_25306_, _25322_, _25323_);
  or g_56267_(_25314_, _25323_, _25324_);
  xor g_56268_(out[103], out[343], _25325_);
  and g_56269_(_39570_, out[347], _25326_);
  xor g_56270_(out[110], out[350], _25327_);
  xor g_56271_(out[104], out[344], _25328_);
  xor g_56272_(out[97], out[337], _25329_);
  xor g_56273_(out[109], out[349], _25330_);
  xor g_56274_(out[105], out[345], _25331_);
  xor g_56275_(out[100], out[340], _25333_);
  xor g_56276_(out[98], out[338], _25334_);
  and g_56277_(out[107], _39735_, _25335_);
  xor g_56278_(out[99], out[339], _25336_);
  xor g_56279_(out[102], out[342], _25337_);
  xor g_56280_(out[111], out[351], _25338_);
  xor g_56281_(out[106], out[346], _25339_);
  xor g_56282_(out[101], out[341], _25340_);
  xor g_56283_(out[96], out[336], _25341_);
  or g_56284_(_25327_, _25333_, _25342_);
  or g_56285_(_25328_, _25330_, _25344_);
  or g_56286_(_25334_, _25339_, _25345_);
  or g_56287_(_25344_, _25345_, _25346_);
  or g_56288_(_25331_, _25336_, _25347_);
  or g_56289_(_25340_, _25341_, _25348_);
  or g_56290_(_25347_, _25348_, _25349_);
  or g_56291_(_25346_, _25349_, _25350_);
  xor g_56292_(out[108], out[348], _25351_);
  or g_56293_(_25326_, _25351_, _25352_);
  or g_56294_(_25325_, _25337_, _25353_);
  or g_56295_(_25352_, _25353_, _25355_);
  or g_56296_(_25329_, _25335_, _25356_);
  or g_56297_(_25338_, _25356_, _25357_);
  or g_56298_(_25355_, _25357_, _25358_);
  or g_56299_(_25350_, _25358_, _25359_);
  or g_56300_(_25342_, _25359_, _25360_);
  not g_56301_(_25360_, _25361_);
  xor g_56302_(out[81], out[337], _25362_);
  and g_56303_(out[91], _39735_, _25363_);
  xor g_56304_(out[89], out[345], _25364_);
  xor g_56305_(out[80], out[336], _25366_);
  xor g_56306_(out[94], out[350], _25367_);
  xor g_56307_(out[84], out[340], _25368_);
  or g_56308_(_25367_, _25368_, _25369_);
  xor g_56309_(out[93], out[349], _25370_);
  xor g_56310_(out[83], out[339], _25371_);
  and g_56311_(_39559_, out[347], _25372_);
  xor g_56312_(out[86], out[342], _25373_);
  xor g_56313_(out[90], out[346], _25374_);
  xor g_56314_(out[85], out[341], _25375_);
  xor g_56315_(out[95], out[351], _25377_);
  xor g_56316_(out[88], out[344], _25378_);
  or g_56317_(_25370_, _25378_, _25379_);
  xor g_56318_(out[82], out[338], _25380_);
  or g_56319_(_25374_, _25380_, _25381_);
  or g_56320_(_25379_, _25381_, _25382_);
  or g_56321_(_25364_, _25371_, _25383_);
  or g_56322_(_25375_, _25383_, _25384_);
  or g_56323_(_25382_, _25384_, _25385_);
  or g_56324_(_25369_, _25385_, _25386_);
  xor g_56325_(out[92], out[348], _25388_);
  or g_56326_(_25372_, _25388_, _25389_);
  xor g_56327_(out[87], out[343], _25390_);
  or g_56328_(_25373_, _25390_, _25391_);
  or g_56329_(_25389_, _25391_, _25392_);
  or g_56330_(_25362_, _25363_, _25393_);
  or g_56331_(_25377_, _25393_, _25394_);
  or g_56332_(_25392_, _25394_, _25395_);
  or g_56333_(_25366_, _25395_, _25396_);
  or g_56334_(_25386_, _25396_, _25397_);
  xor g_56335_(out[71], out[343], _25399_);
  and g_56336_(_39548_, out[347], _25400_);
  xor g_56337_(out[78], out[350], _25401_);
  xor g_56338_(out[72], out[344], _25402_);
  xor g_56339_(out[65], out[337], _25403_);
  xor g_56340_(out[77], out[349], _25404_);
  xor g_56341_(out[73], out[345], _25405_);
  xor g_56342_(out[68], out[340], _25406_);
  xor g_56343_(out[66], out[338], _25407_);
  and g_56344_(out[75], _39735_, _25408_);
  xor g_56345_(out[67], out[339], _25410_);
  xor g_56346_(out[70], out[342], _25411_);
  xor g_56347_(out[79], out[351], _25412_);
  xor g_56348_(out[74], out[346], _25413_);
  xor g_56349_(out[69], out[341], _25414_);
  xor g_56350_(out[64], out[336], _25415_);
  or g_56351_(_25401_, _25406_, _25416_);
  or g_56352_(_25402_, _25404_, _25417_);
  or g_56353_(_25407_, _25413_, _25418_);
  or g_56354_(_25417_, _25418_, _25419_);
  or g_56355_(_25405_, _25410_, _25421_);
  or g_56356_(_25414_, _25415_, _25422_);
  or g_56357_(_25421_, _25422_, _25423_);
  or g_56358_(_25419_, _25423_, _25424_);
  xor g_56359_(out[76], out[348], _25425_);
  or g_56360_(_25400_, _25425_, _25426_);
  or g_56361_(_25399_, _25411_, _25427_);
  or g_56362_(_25426_, _25427_, _25428_);
  or g_56363_(_25403_, _25408_, _25429_);
  or g_56364_(_25412_, _25429_, _25430_);
  or g_56365_(_25428_, _25430_, _25432_);
  or g_56366_(_25424_, _25432_, _25433_);
  or g_56367_(_25416_, _25433_, _25434_);
  xor g_56368_(out[49], out[337], _25435_);
  and g_56369_(out[59], _39735_, _25436_);
  xor g_56370_(out[57], out[345], _25437_);
  xor g_56371_(out[48], out[336], _25438_);
  xor g_56372_(out[62], out[350], _25439_);
  xor g_56373_(out[52], out[340], _25440_);
  or g_56374_(_25439_, _25440_, _25441_);
  xor g_56375_(out[61], out[349], _25443_);
  xor g_56376_(out[51], out[339], _25444_);
  and g_56377_(_39537_, out[347], _25445_);
  xor g_56378_(out[54], out[342], _25446_);
  xor g_56379_(out[58], out[346], _25447_);
  xor g_56380_(out[53], out[341], _25448_);
  xor g_56381_(out[63], out[351], _25449_);
  xor g_56382_(out[56], out[344], _25450_);
  or g_56383_(_25443_, _25450_, _25451_);
  xor g_56384_(out[50], out[338], _25452_);
  or g_56385_(_25447_, _25452_, _25454_);
  or g_56386_(_25451_, _25454_, _25455_);
  or g_56387_(_25437_, _25444_, _25456_);
  or g_56388_(_25448_, _25456_, _25457_);
  or g_56389_(_25455_, _25457_, _25458_);
  or g_56390_(_25441_, _25458_, _25459_);
  xor g_56391_(out[60], out[348], _25460_);
  or g_56392_(_25445_, _25460_, _25461_);
  xor g_56393_(out[55], out[343], _25462_);
  or g_56394_(_25446_, _25462_, _25463_);
  or g_56395_(_25461_, _25463_, _25465_);
  or g_56396_(_25435_, _25436_, _25466_);
  or g_56397_(_25449_, _25466_, _25467_);
  or g_56398_(_25465_, _25467_, _25468_);
  or g_56399_(_25438_, _25468_, _25469_);
  or g_56400_(_25459_, _25469_, _25470_);
  xor g_56401_(out[39], out[343], _25471_);
  and g_56402_(_39526_, out[347], _25472_);
  xor g_56403_(out[46], out[350], _25473_);
  xor g_56404_(out[40], out[344], _25474_);
  xor g_56405_(out[33], out[337], _25476_);
  xor g_56406_(out[45], out[349], _25477_);
  xor g_56407_(out[41], out[345], _25478_);
  xor g_56408_(out[36], out[340], _25479_);
  xor g_56409_(out[34], out[338], _25480_);
  and g_56410_(out[43], _39735_, _25481_);
  xor g_56411_(out[35], out[339], _25482_);
  xor g_56412_(out[38], out[342], _25483_);
  xor g_56413_(out[47], out[351], _25484_);
  xor g_56414_(out[42], out[346], _25485_);
  xor g_56415_(out[37], out[341], _25487_);
  xor g_56416_(out[32], out[336], _25488_);
  or g_56417_(_25473_, _25479_, _25489_);
  or g_56418_(_25474_, _25477_, _25490_);
  or g_56419_(_25480_, _25485_, _25491_);
  or g_56420_(_25490_, _25491_, _25492_);
  or g_56421_(_25478_, _25482_, _25493_);
  or g_56422_(_25487_, _25488_, _25494_);
  or g_56423_(_25493_, _25494_, _25495_);
  or g_56424_(_25492_, _25495_, _25496_);
  xor g_56425_(out[44], out[348], _25498_);
  or g_56426_(_25472_, _25498_, _25499_);
  or g_56427_(_25471_, _25483_, _25500_);
  or g_56428_(_25499_, _25500_, _25501_);
  or g_56429_(_25476_, _25481_, _25502_);
  or g_56430_(_25484_, _25502_, _25503_);
  or g_56431_(_25501_, _25503_, _25504_);
  or g_56432_(_25496_, _25504_, _25505_);
  or g_56433_(_25489_, _25505_, _25506_);
  xor g_56434_(out[17], out[337], _25507_);
  and g_56435_(out[27], _39735_, _25509_);
  xor g_56436_(out[25], out[345], _25510_);
  xor g_56437_(out[16], out[336], _25511_);
  xor g_56438_(out[30], out[350], _25512_);
  xor g_56439_(out[20], out[340], _25513_);
  or g_56440_(_25512_, _25513_, _25514_);
  xor g_56441_(out[29], out[349], _25515_);
  xor g_56442_(out[19], out[339], _25516_);
  and g_56443_(_39493_, out[347], _25517_);
  xor g_56444_(out[22], out[342], _25518_);
  xor g_56445_(out[26], out[346], _25520_);
  xor g_56446_(out[21], out[341], _25521_);
  xor g_56447_(out[31], out[351], _25522_);
  xor g_56448_(out[24], out[344], _25523_);
  or g_56449_(_25515_, _25523_, _25524_);
  xor g_56450_(out[18], out[338], _25525_);
  or g_56451_(_25520_, _25525_, _25526_);
  or g_56452_(_25524_, _25526_, _25527_);
  or g_56453_(_25510_, _25516_, _25528_);
  or g_56454_(_25521_, _25528_, _25529_);
  or g_56455_(_25527_, _25529_, _25531_);
  or g_56456_(_25514_, _25531_, _25532_);
  xor g_56457_(out[28], out[348], _25533_);
  or g_56458_(_25517_, _25533_, _25534_);
  xor g_56459_(out[23], out[343], _25535_);
  or g_56460_(_25518_, _25535_, _25536_);
  or g_56461_(_25534_, _25536_, _25537_);
  or g_56462_(_25507_, _25509_, _25538_);
  or g_56463_(_25522_, _25538_, _25539_);
  or g_56464_(_25537_, _25539_, _25540_);
  or g_56465_(_25511_, _25540_, _25542_);
  or g_56466_(_25532_, _25542_, _25543_);
  not g_56467_(_25543_, _25544_);
  and g_56468_(out[11], _39735_, _25545_);
  and g_56469_(_39438_, out[347], _25546_);
  xor g_56470_(out[8], out[344], _25547_);
  xor g_56471_(out[15], out[351], _25548_);
  xor g_56472_(out[1], out[337], _25549_);
  xor g_56473_(out[2], out[338], _25550_);
  xor g_56474_(out[4], out[340], _25551_);
  xor g_56475_(out[5], out[341], _25553_);
  xor g_56476_(out[9], out[345], _25554_);
  xor g_56477_(out[3], out[339], _25555_);
  xor g_56478_(out[14], out[350], _25556_);
  xor g_56479_(out[0], out[336], _25557_);
  xor g_56480_(out[10], out[346], _25558_);
  xor g_56481_(out[13], out[349], _25559_);
  or g_56482_(_25547_, _25559_, _25560_);
  xor g_56483_(out[6], out[342], _25561_);
  or g_56484_(_25550_, _25558_, _25562_);
  or g_56485_(_25560_, _25562_, _25564_);
  or g_56486_(_25554_, _25555_, _25565_);
  or g_56487_(_25553_, _25565_, _25566_);
  or g_56488_(_25564_, _25566_, _25567_);
  or g_56489_(_25551_, _25556_, _25568_);
  or g_56490_(_25567_, _25568_, _25569_);
  xor g_56491_(out[12], out[348], _25570_);
  or g_56492_(_25546_, _25570_, _25571_);
  xor g_56493_(out[7], out[343], _25572_);
  or g_56494_(_25561_, _25572_, _25573_);
  or g_56495_(_25571_, _25573_, _25575_);
  or g_56496_(_25545_, _25549_, _25576_);
  or g_56497_(_25548_, _25576_, _25577_);
  or g_56498_(_25575_, _25577_, _25578_);
  or g_56499_(_25557_, _25578_, _25579_);
  or g_56500_(_25569_, _25579_, _25580_);
  xor g_56501_(out[330], out[314], _25581_);
  xor g_56502_(out[322], out[306], _25582_);
  xor g_56503_(out[321], out[305], _25583_);
  and g_56504_(_39427_, out[315], _25584_);
  and g_56505_(out[331], _39724_, _25586_);
  xor g_56506_(out[333], out[317], _25587_);
  xor g_56507_(out[323], out[307], _25588_);
  xor g_56508_(out[334], out[318], _25589_);
  xor g_56509_(out[332], out[316], _25590_);
  xor g_56510_(out[328], out[312], _25591_);
  xor g_56511_(out[335], out[319], _25592_);
  xor g_56512_(out[325], out[309], _25593_);
  xor g_56513_(out[326], out[310], _25594_);
  xor g_56514_(out[320], out[304], _25595_);
  xor g_56515_(out[324], out[308], _25597_);
  or g_56516_(_25587_, _25591_, _25598_);
  xor g_56517_(out[329], out[313], _25599_);
  or g_56518_(_25581_, _25582_, _25600_);
  or g_56519_(_25598_, _25600_, _25601_);
  or g_56520_(_25588_, _25599_, _25602_);
  or g_56521_(_25593_, _25602_, _25603_);
  or g_56522_(_25601_, _25603_, _25604_);
  or g_56523_(_25589_, _25597_, _25605_);
  or g_56524_(_25604_, _25605_, _25606_);
  or g_56525_(_25584_, _25590_, _25608_);
  xor g_56526_(out[327], out[311], _25609_);
  or g_56527_(_25594_, _25609_, _25610_);
  or g_56528_(_25608_, _25610_, _25611_);
  or g_56529_(_25583_, _25586_, _25612_);
  or g_56530_(_25592_, _25612_, _25613_);
  or g_56531_(_25611_, _25613_, _25614_);
  or g_56532_(_25595_, _25614_, _25615_);
  or g_56533_(_25606_, _25615_, _25616_);
  xor g_56534_(out[332], out[300], _25617_);
  and g_56535_(_39427_, out[299], _25619_);
  xor g_56536_(out[328], out[296], _25620_);
  xor g_56537_(out[326], out[294], _25621_);
  xor g_56538_(out[333], out[301], _25622_);
  xor g_56539_(out[334], out[302], _25623_);
  xor g_56540_(out[322], out[290], _25624_);
  xor g_56541_(out[329], out[297], _25625_);
  xor g_56542_(out[325], out[293], _25626_);
  xor g_56543_(out[321], out[289], _25627_);
  and g_56544_(out[331], _39702_, _25628_);
  or g_56545_(_25620_, _25622_, _25630_);
  xor g_56546_(out[335], out[303], _25631_);
  xor g_56547_(out[330], out[298], _25632_);
  xor g_56548_(out[324], out[292], _25633_);
  xor g_56549_(out[323], out[291], _25634_);
  xor g_56550_(out[320], out[288], _25635_);
  or g_56551_(_25624_, _25632_, _25636_);
  or g_56552_(_25630_, _25636_, _25637_);
  or g_56553_(_25625_, _25634_, _25638_);
  or g_56554_(_25626_, _25638_, _25639_);
  or g_56555_(_25637_, _25639_, _25641_);
  or g_56556_(_25623_, _25633_, _25642_);
  or g_56557_(_25641_, _25642_, _25643_);
  or g_56558_(_25617_, _25619_, _25644_);
  xor g_56559_(out[327], out[295], _25645_);
  or g_56560_(_25621_, _25645_, _25646_);
  or g_56561_(_25644_, _25646_, _25647_);
  or g_56562_(_25627_, _25628_, _25648_);
  or g_56563_(_25631_, _25648_, _25649_);
  or g_56564_(_25647_, _25649_, _25650_);
  or g_56565_(_25635_, _25650_, _25652_);
  or g_56566_(_25643_, _25652_, _25653_);
  xor g_56567_(out[321], out[273], _25654_);
  and g_56568_(_39427_, out[283], _25655_);
  and g_56569_(out[331], _39691_, _25656_);
  xor g_56570_(out[329], out[281], _25657_);
  xor g_56571_(out[320], out[272], _25658_);
  xor g_56572_(out[334], out[286], _25659_);
  xor g_56573_(out[324], out[276], _25660_);
  or g_56574_(_25659_, _25660_, _25661_);
  xor g_56575_(out[333], out[285], _25663_);
  xor g_56576_(out[323], out[275], _25664_);
  xor g_56577_(out[332], out[284], _25665_);
  xor g_56578_(out[326], out[278], _25666_);
  xor g_56579_(out[330], out[282], _25667_);
  xor g_56580_(out[325], out[277], _25668_);
  xor g_56581_(out[335], out[287], _25669_);
  xor g_56582_(out[328], out[280], _25670_);
  or g_56583_(_25663_, _25670_, _25671_);
  xor g_56584_(out[322], out[274], _25672_);
  or g_56585_(_25667_, _25672_, _25674_);
  or g_56586_(_25671_, _25674_, _25675_);
  or g_56587_(_25657_, _25664_, _25676_);
  or g_56588_(_25668_, _25676_, _25677_);
  or g_56589_(_25675_, _25677_, _25678_);
  or g_56590_(_25661_, _25678_, _25679_);
  or g_56591_(_25655_, _25665_, _25680_);
  xor g_56592_(out[327], out[279], _25681_);
  or g_56593_(_25666_, _25681_, _25682_);
  or g_56594_(_25680_, _25682_, _25683_);
  or g_56595_(_25654_, _25656_, _25685_);
  or g_56596_(_25669_, _25685_, _25686_);
  or g_56597_(_25683_, _25686_, _25687_);
  or g_56598_(_25658_, _25687_, _25688_);
  or g_56599_(_25679_, _25688_, _25689_);
  xor g_56600_(out[321], out[257], _25690_);
  and g_56601_(out[331], _39680_, _25691_);
  xor g_56602_(out[329], out[265], _25692_);
  xor g_56603_(out[320], out[256], _25693_);
  xor g_56604_(out[334], out[270], _25694_);
  xor g_56605_(out[324], out[260], _25696_);
  or g_56606_(_25694_, _25696_, _25697_);
  xor g_56607_(out[333], out[269], _25698_);
  xor g_56608_(out[323], out[259], _25699_);
  and g_56609_(_39427_, out[267], _25700_);
  xor g_56610_(out[326], out[262], _25701_);
  xor g_56611_(out[330], out[266], _25702_);
  xor g_56612_(out[325], out[261], _25703_);
  xor g_56613_(out[335], out[271], _25704_);
  xor g_56614_(out[328], out[264], _25705_);
  or g_56615_(_25698_, _25705_, _25707_);
  xor g_56616_(out[322], out[258], _25708_);
  or g_56617_(_25702_, _25708_, _25709_);
  or g_56618_(_25707_, _25709_, _25710_);
  or g_56619_(_25692_, _25699_, _25711_);
  or g_56620_(_25703_, _25711_, _25712_);
  or g_56621_(_25710_, _25712_, _25713_);
  or g_56622_(_25697_, _25713_, _25714_);
  xor g_56623_(out[332], out[268], _25715_);
  or g_56624_(_25700_, _25715_, _25716_);
  xor g_56625_(out[327], out[263], _25718_);
  or g_56626_(_25701_, _25718_, _25719_);
  or g_56627_(_25716_, _25719_, _25720_);
  or g_56628_(_25690_, _25691_, _25721_);
  or g_56629_(_25704_, _25721_, _25722_);
  or g_56630_(_25720_, _25722_, _25723_);
  or g_56631_(_25693_, _25723_, _25724_);
  or g_56632_(_25714_, _25724_, _25725_);
  not g_56633_(_25725_, _25726_);
  and g_56634_(out[331], _39669_, _25727_);
  and g_56635_(_39427_, out[251], _25729_);
  xor g_56636_(out[328], out[248], _25730_);
  xor g_56637_(out[335], out[255], _25731_);
  xor g_56638_(out[321], out[241], _25732_);
  xor g_56639_(out[322], out[242], _25733_);
  xor g_56640_(out[324], out[244], _25734_);
  xor g_56641_(out[325], out[245], _25735_);
  xor g_56642_(out[329], out[249], _25736_);
  xor g_56643_(out[323], out[243], _25737_);
  xor g_56644_(out[334], out[254], _25738_);
  xor g_56645_(out[320], out[240], _25740_);
  xor g_56646_(out[330], out[250], _25741_);
  xor g_56647_(out[333], out[253], _25742_);
  or g_56648_(_25730_, _25742_, _25743_);
  xor g_56649_(out[326], out[246], _25744_);
  or g_56650_(_25733_, _25741_, _25745_);
  or g_56651_(_25743_, _25745_, _25746_);
  or g_56652_(_25736_, _25737_, _25747_);
  or g_56653_(_25735_, _25747_, _25748_);
  or g_56654_(_25746_, _25748_, _25749_);
  or g_56655_(_25734_, _25738_, _25751_);
  or g_56656_(_25749_, _25751_, _25752_);
  xor g_56657_(out[332], out[252], _25753_);
  or g_56658_(_25729_, _25753_, _25754_);
  xor g_56659_(out[327], out[247], _25755_);
  or g_56660_(_25744_, _25755_, _25756_);
  or g_56661_(_25754_, _25756_, _25757_);
  or g_56662_(_25727_, _25732_, _25758_);
  or g_56663_(_25731_, _25758_, _25759_);
  or g_56664_(_25757_, _25759_, _25760_);
  or g_56665_(_25740_, _25760_, _25762_);
  or g_56666_(_25752_, _25762_, _25763_);
  xor g_56667_(out[321], out[225], _25764_);
  and g_56668_(_39427_, out[235], _25765_);
  and g_56669_(out[331], _39658_, _25766_);
  xor g_56670_(out[334], out[238], _25767_);
  xor g_56671_(out[323], out[227], _25768_);
  xor g_56672_(out[324], out[228], _25769_);
  xor g_56673_(out[322], out[226], _25770_);
  xor g_56674_(out[329], out[233], _25771_);
  xor g_56675_(out[320], out[224], _25773_);
  xor g_56676_(out[332], out[236], _25774_);
  xor g_56677_(out[326], out[230], _25775_);
  xor g_56678_(out[330], out[234], _25776_);
  xor g_56679_(out[325], out[229], _25777_);
  xor g_56680_(out[335], out[239], _25778_);
  xor g_56681_(out[333], out[237], _25779_);
  xor g_56682_(out[328], out[232], _25780_);
  or g_56683_(_25767_, _25769_, _25781_);
  or g_56684_(_25779_, _25780_, _25782_);
  or g_56685_(_25770_, _25776_, _25784_);
  or g_56686_(_25782_, _25784_, _25785_);
  or g_56687_(_25768_, _25771_, _25786_);
  or g_56688_(_25773_, _25777_, _25787_);
  or g_56689_(_25786_, _25787_, _25788_);
  or g_56690_(_25785_, _25788_, _25789_);
  or g_56691_(_25765_, _25774_, _25790_);
  xor g_56692_(out[327], out[231], _25791_);
  or g_56693_(_25775_, _25791_, _25792_);
  or g_56694_(_25790_, _25792_, _25793_);
  or g_56695_(_25764_, _25766_, _25795_);
  or g_56696_(_25778_, _25795_, _25796_);
  or g_56697_(_25793_, _25796_, _25797_);
  or g_56698_(_25789_, _25797_, _25798_);
  or g_56699_(_25781_, _25798_, _25799_);
  xor g_56700_(out[328], out[216], _25800_);
  xor g_56701_(out[325], out[213], _25801_);
  xor g_56702_(out[323], out[211], _25802_);
  xor g_56703_(out[334], out[222], _25803_);
  xor g_56704_(out[333], out[221], _25804_);
  xor g_56705_(out[322], out[210], _25806_);
  xor g_56706_(out[329], out[217], _25807_);
  xor g_56707_(out[326], out[214], _25808_);
  xor g_56708_(out[335], out[223], _25809_);
  xor g_56709_(out[330], out[218], _25810_);
  xor g_56710_(out[324], out[212], _25811_);
  xor g_56711_(out[320], out[208], _25812_);
  and g_56712_(_39427_, out[219], _25813_);
  and g_56713_(out[331], _39647_, _25814_);
  or g_56714_(_25800_, _25804_, _25815_);
  xor g_56715_(out[321], out[209], _25817_);
  or g_56716_(_25806_, _25810_, _25818_);
  or g_56717_(_25815_, _25818_, _25819_);
  or g_56718_(_25802_, _25807_, _25820_);
  or g_56719_(_25801_, _25820_, _25821_);
  or g_56720_(_25819_, _25821_, _25822_);
  or g_56721_(_25803_, _25811_, _25823_);
  or g_56722_(_25822_, _25823_, _25824_);
  xor g_56723_(out[332], out[220], _25825_);
  or g_56724_(_25813_, _25825_, _25826_);
  xor g_56725_(out[327], out[215], _25828_);
  or g_56726_(_25808_, _25828_, _25829_);
  or g_56727_(_25826_, _25829_, _25830_);
  or g_56728_(_25814_, _25817_, _25831_);
  or g_56729_(_25809_, _25831_, _25832_);
  or g_56730_(_25830_, _25832_, _25833_);
  or g_56731_(_25812_, _25833_, _25834_);
  or g_56732_(_25824_, _25834_, _25835_);
  not g_56733_(_25835_, _25836_);
  xor g_56734_(out[330], out[202], _25837_);
  xor g_56735_(out[322], out[194], _25839_);
  xor g_56736_(out[321], out[193], _25840_);
  and g_56737_(_39427_, out[203], _25841_);
  and g_56738_(out[331], _39636_, _25842_);
  xor g_56739_(out[333], out[205], _25843_);
  xor g_56740_(out[323], out[195], _25844_);
  xor g_56741_(out[334], out[206], _25845_);
  xor g_56742_(out[332], out[204], _25846_);
  xor g_56743_(out[328], out[200], _25847_);
  xor g_56744_(out[335], out[207], _25848_);
  xor g_56745_(out[325], out[197], _25850_);
  xor g_56746_(out[326], out[198], _25851_);
  xor g_56747_(out[320], out[192], _25852_);
  xor g_56748_(out[324], out[196], _25853_);
  or g_56749_(_25843_, _25847_, _25854_);
  xor g_56750_(out[329], out[201], _25855_);
  or g_56751_(_25837_, _25839_, _25856_);
  or g_56752_(_25854_, _25856_, _25857_);
  or g_56753_(_25844_, _25855_, _25858_);
  or g_56754_(_25850_, _25858_, _25859_);
  or g_56755_(_25857_, _25859_, _25861_);
  or g_56756_(_25845_, _25853_, _25862_);
  or g_56757_(_25861_, _25862_, _25863_);
  or g_56758_(_25841_, _25846_, _25864_);
  xor g_56759_(out[327], out[199], _25865_);
  or g_56760_(_25851_, _25865_, _25866_);
  or g_56761_(_25864_, _25866_, _25867_);
  or g_56762_(_25840_, _25842_, _25868_);
  or g_56763_(_25848_, _25868_, _25869_);
  or g_56764_(_25867_, _25869_, _25870_);
  or g_56765_(_25852_, _25870_, _25872_);
  or g_56766_(_25863_, _25872_, _25873_);
  not g_56767_(_25873_, _25874_);
  xor g_56768_(out[321], out[177], _25875_);
  and g_56769_(out[331], _39625_, _25876_);
  xor g_56770_(out[329], out[185], _25877_);
  xor g_56771_(out[320], out[176], _25878_);
  xor g_56772_(out[334], out[190], _25879_);
  xor g_56773_(out[324], out[180], _25880_);
  or g_56774_(_25879_, _25880_, _25881_);
  xor g_56775_(out[333], out[189], _25883_);
  xor g_56776_(out[323], out[179], _25884_);
  and g_56777_(_39427_, out[187], _25885_);
  xor g_56778_(out[326], out[182], _25886_);
  xor g_56779_(out[330], out[186], _25887_);
  xor g_56780_(out[325], out[181], _25888_);
  xor g_56781_(out[335], out[191], _25889_);
  xor g_56782_(out[328], out[184], _25890_);
  or g_56783_(_25883_, _25890_, _25891_);
  xor g_56784_(out[322], out[178], _25892_);
  or g_56785_(_25887_, _25892_, _25894_);
  or g_56786_(_25891_, _25894_, _25895_);
  or g_56787_(_25877_, _25884_, _25896_);
  or g_56788_(_25888_, _25896_, _25897_);
  or g_56789_(_25895_, _25897_, _25898_);
  or g_56790_(_25881_, _25898_, _25899_);
  xor g_56791_(out[332], out[188], _25900_);
  or g_56792_(_25885_, _25900_, _25901_);
  xor g_56793_(out[327], out[183], _25902_);
  or g_56794_(_25886_, _25902_, _25903_);
  or g_56795_(_25901_, _25903_, _25905_);
  or g_56796_(_25875_, _25876_, _25906_);
  or g_56797_(_25889_, _25906_, _25907_);
  or g_56798_(_25905_, _25907_, _25908_);
  or g_56799_(_25878_, _25908_, _25909_);
  or g_56800_(_25899_, _25909_, _25910_);
  xor g_56801_(out[321], out[161], _25911_);
  and g_56802_(_39427_, out[171], _25912_);
  and g_56803_(out[331], _39614_, _25913_);
  xor g_56804_(out[329], out[169], _25914_);
  xor g_56805_(out[320], out[160], _25916_);
  xor g_56806_(out[334], out[174], _25917_);
  xor g_56807_(out[324], out[164], _25918_);
  or g_56808_(_25917_, _25918_, _25919_);
  xor g_56809_(out[333], out[173], _25920_);
  xor g_56810_(out[323], out[163], _25921_);
  xor g_56811_(out[332], out[172], _25922_);
  xor g_56812_(out[326], out[166], _25923_);
  xor g_56813_(out[330], out[170], _25924_);
  xor g_56814_(out[325], out[165], _25925_);
  xor g_56815_(out[335], out[175], _25927_);
  xor g_56816_(out[328], out[168], _25928_);
  or g_56817_(_25920_, _25928_, _25929_);
  xor g_56818_(out[322], out[162], _25930_);
  or g_56819_(_25924_, _25930_, _25931_);
  or g_56820_(_25929_, _25931_, _25932_);
  or g_56821_(_25914_, _25921_, _25933_);
  or g_56822_(_25925_, _25933_, _25934_);
  or g_56823_(_25932_, _25934_, _25935_);
  or g_56824_(_25919_, _25935_, _25936_);
  or g_56825_(_25912_, _25922_, _25938_);
  xor g_56826_(out[327], out[167], _25939_);
  or g_56827_(_25923_, _25939_, _25940_);
  or g_56828_(_25938_, _25940_, _25941_);
  or g_56829_(_25911_, _25913_, _25942_);
  or g_56830_(_25927_, _25942_, _25943_);
  or g_56831_(_25941_, _25943_, _25944_);
  or g_56832_(_25916_, _25944_, _25945_);
  or g_56833_(_25936_, _25945_, _25946_);
  xor g_56834_(out[333], out[157], _25947_);
  xor g_56835_(out[322], out[146], _25949_);
  xor g_56836_(out[325], out[149], _25950_);
  xor g_56837_(out[329], out[153], _25951_);
  xor g_56838_(out[324], out[148], _25952_);
  xor g_56839_(out[328], out[152], _25953_);
  xor g_56840_(out[334], out[158], _25954_);
  xor g_56841_(out[326], out[150], _25955_);
  xor g_56842_(out[335], out[159], _25956_);
  xor g_56843_(out[330], out[154], _25957_);
  xor g_56844_(out[320], out[144], _25958_);
  xor g_56845_(out[323], out[147], _25960_);
  and g_56846_(_39427_, out[155], _25961_);
  and g_56847_(out[331], _39603_, _25962_);
  xor g_56848_(out[321], out[145], _25963_);
  or g_56849_(_25952_, _25954_, _25964_);
  or g_56850_(_25947_, _25953_, _25965_);
  or g_56851_(_25949_, _25957_, _25966_);
  or g_56852_(_25965_, _25966_, _25967_);
  or g_56853_(_25951_, _25960_, _25968_);
  or g_56854_(_25950_, _25958_, _25969_);
  or g_56855_(_25968_, _25969_, _25971_);
  or g_56856_(_25967_, _25971_, _25972_);
  xor g_56857_(out[332], out[156], _25973_);
  or g_56858_(_25961_, _25973_, _25974_);
  xor g_56859_(out[327], out[151], _25975_);
  or g_56860_(_25955_, _25975_, _25976_);
  or g_56861_(_25974_, _25976_, _25977_);
  or g_56862_(_25962_, _25963_, _25978_);
  or g_56863_(_25956_, _25978_, _25979_);
  or g_56864_(_25977_, _25979_, _25980_);
  or g_56865_(_25972_, _25980_, _25982_);
  or g_56866_(_25964_, _25982_, _25983_);
  not g_56867_(_25983_, _25984_);
  xor g_56868_(out[321], out[129], _25985_);
  and g_56869_(out[331], _39592_, _25986_);
  xor g_56870_(out[329], out[137], _25987_);
  xor g_56871_(out[320], out[128], _25988_);
  xor g_56872_(out[334], out[142], _25989_);
  xor g_56873_(out[324], out[132], _25990_);
  or g_56874_(_25989_, _25990_, _25991_);
  xor g_56875_(out[333], out[141], _25993_);
  xor g_56876_(out[323], out[131], _25994_);
  and g_56877_(_39427_, out[139], _25995_);
  xor g_56878_(out[326], out[134], _25996_);
  xor g_56879_(out[330], out[138], _25997_);
  xor g_56880_(out[325], out[133], _25998_);
  xor g_56881_(out[335], out[143], _25999_);
  xor g_56882_(out[328], out[136], _26000_);
  or g_56883_(_25993_, _26000_, _26001_);
  xor g_56884_(out[322], out[130], _26002_);
  or g_56885_(_25997_, _26002_, _26004_);
  or g_56886_(_26001_, _26004_, _26005_);
  or g_56887_(_25987_, _25994_, _26006_);
  or g_56888_(_25998_, _26006_, _26007_);
  or g_56889_(_26005_, _26007_, _26008_);
  or g_56890_(_25991_, _26008_, _26009_);
  xor g_56891_(out[332], out[140], _26010_);
  or g_56892_(_25995_, _26010_, _26011_);
  xor g_56893_(out[327], out[135], _26012_);
  or g_56894_(_25996_, _26012_, _26013_);
  or g_56895_(_26011_, _26013_, _26015_);
  or g_56896_(_25985_, _25986_, _26016_);
  or g_56897_(_25999_, _26016_, _26017_);
  or g_56898_(_26015_, _26017_, _26018_);
  or g_56899_(_25988_, _26018_, _26019_);
  or g_56900_(_26009_, _26019_, _26020_);
  xor g_56901_(out[321], out[113], _26021_);
  and g_56902_(_39427_, out[123], _26022_);
  and g_56903_(out[331], _39581_, _26023_);
  xor g_56904_(out[329], out[121], _26024_);
  xor g_56905_(out[320], out[112], _26026_);
  xor g_56906_(out[334], out[126], _26027_);
  xor g_56907_(out[324], out[116], _26028_);
  or g_56908_(_26027_, _26028_, _26029_);
  xor g_56909_(out[333], out[125], _26030_);
  xor g_56910_(out[323], out[115], _26031_);
  xor g_56911_(out[332], out[124], _26032_);
  xor g_56912_(out[326], out[118], _26033_);
  xor g_56913_(out[330], out[122], _26034_);
  xor g_56914_(out[325], out[117], _26035_);
  xor g_56915_(out[335], out[127], _26037_);
  xor g_56916_(out[328], out[120], _26038_);
  or g_56917_(_26030_, _26038_, _26039_);
  xor g_56918_(out[322], out[114], _26040_);
  or g_56919_(_26034_, _26040_, _26041_);
  or g_56920_(_26039_, _26041_, _26042_);
  or g_56921_(_26024_, _26031_, _26043_);
  or g_56922_(_26035_, _26043_, _26044_);
  or g_56923_(_26042_, _26044_, _26045_);
  or g_56924_(_26029_, _26045_, _26046_);
  or g_56925_(_26022_, _26032_, _26048_);
  xor g_56926_(out[327], out[119], _26049_);
  or g_56927_(_26033_, _26049_, _26050_);
  or g_56928_(_26048_, _26050_, _26051_);
  or g_56929_(_26021_, _26023_, _26052_);
  or g_56930_(_26037_, _26052_, _26053_);
  or g_56931_(_26051_, _26053_, _26054_);
  or g_56932_(_26026_, _26054_, _26055_);
  or g_56933_(_26046_, _26055_, _26056_);
  xor g_56934_(out[321], out[97], _26057_);
  and g_56935_(_39427_, out[107], _26059_);
  and g_56936_(out[331], _39570_, _26060_);
  xor g_56937_(out[334], out[110], _26061_);
  xor g_56938_(out[323], out[99], _26062_);
  xor g_56939_(out[324], out[100], _26063_);
  xor g_56940_(out[322], out[98], _26064_);
  xor g_56941_(out[329], out[105], _26065_);
  xor g_56942_(out[320], out[96], _26066_);
  xor g_56943_(out[332], out[108], _26067_);
  xor g_56944_(out[326], out[102], _26068_);
  xor g_56945_(out[330], out[106], _26070_);
  xor g_56946_(out[325], out[101], _26071_);
  xor g_56947_(out[335], out[111], _26072_);
  xor g_56948_(out[333], out[109], _26073_);
  xor g_56949_(out[328], out[104], _26074_);
  or g_56950_(_26061_, _26063_, _26075_);
  or g_56951_(_26073_, _26074_, _26076_);
  or g_56952_(_26064_, _26070_, _26077_);
  or g_56953_(_26076_, _26077_, _26078_);
  or g_56954_(_26062_, _26065_, _26079_);
  or g_56955_(_26066_, _26071_, _26081_);
  or g_56956_(_26079_, _26081_, _26082_);
  or g_56957_(_26078_, _26082_, _26083_);
  or g_56958_(_26059_, _26067_, _26084_);
  xor g_56959_(out[327], out[103], _26085_);
  or g_56960_(_26068_, _26085_, _26086_);
  or g_56961_(_26084_, _26086_, _26087_);
  or g_56962_(_26057_, _26060_, _26088_);
  or g_56963_(_26072_, _26088_, _26089_);
  or g_56964_(_26087_, _26089_, _26090_);
  or g_56965_(_26083_, _26090_, _26092_);
  or g_56966_(_26075_, _26092_, _26093_);
  xor g_56967_(out[328], out[88], _26094_);
  xor g_56968_(out[325], out[85], _26095_);
  xor g_56969_(out[323], out[83], _26096_);
  xor g_56970_(out[334], out[94], _26097_);
  xor g_56971_(out[333], out[93], _26098_);
  xor g_56972_(out[322], out[82], _26099_);
  xor g_56973_(out[329], out[89], _26100_);
  xor g_56974_(out[326], out[86], _26101_);
  xor g_56975_(out[335], out[95], _26103_);
  xor g_56976_(out[330], out[90], _26104_);
  xor g_56977_(out[324], out[84], _26105_);
  xor g_56978_(out[320], out[80], _26106_);
  and g_56979_(_39427_, out[91], _26107_);
  and g_56980_(out[331], _39559_, _26108_);
  or g_56981_(_26094_, _26098_, _26109_);
  xor g_56982_(out[321], out[81], _26110_);
  or g_56983_(_26099_, _26104_, _26111_);
  or g_56984_(_26109_, _26111_, _26112_);
  or g_56985_(_26096_, _26100_, _26114_);
  or g_56986_(_26095_, _26114_, _26115_);
  or g_56987_(_26112_, _26115_, _26116_);
  or g_56988_(_26097_, _26105_, _26117_);
  or g_56989_(_26116_, _26117_, _26118_);
  xor g_56990_(out[332], out[92], _26119_);
  or g_56991_(_26107_, _26119_, _26120_);
  xor g_56992_(out[327], out[87], _26121_);
  or g_56993_(_26101_, _26121_, _26122_);
  or g_56994_(_26120_, _26122_, _26123_);
  or g_56995_(_26108_, _26110_, _26125_);
  or g_56996_(_26103_, _26125_, _26126_);
  or g_56997_(_26123_, _26126_, _26127_);
  or g_56998_(_26106_, _26127_, _26128_);
  or g_56999_(_26118_, _26128_, _26129_);
  xor g_57000_(out[321], out[65], _26130_);
  and g_57001_(_39427_, out[75], _26131_);
  and g_57002_(out[331], _39548_, _26132_);
  xor g_57003_(out[329], out[73], _26133_);
  xor g_57004_(out[320], out[64], _26134_);
  xor g_57005_(out[334], out[78], _26136_);
  xor g_57006_(out[324], out[68], _26137_);
  or g_57007_(_26136_, _26137_, _26138_);
  xor g_57008_(out[333], out[77], _26139_);
  xor g_57009_(out[323], out[67], _26140_);
  xor g_57010_(out[332], out[76], _26141_);
  xor g_57011_(out[326], out[70], _26142_);
  xor g_57012_(out[330], out[74], _26143_);
  xor g_57013_(out[325], out[69], _26144_);
  xor g_57014_(out[335], out[79], _26145_);
  xor g_57015_(out[328], out[72], _26147_);
  or g_57016_(_26139_, _26147_, _26148_);
  xor g_57017_(out[322], out[66], _26149_);
  or g_57018_(_26143_, _26149_, _26150_);
  or g_57019_(_26148_, _26150_, _26151_);
  or g_57020_(_26133_, _26140_, _26152_);
  or g_57021_(_26144_, _26152_, _26153_);
  or g_57022_(_26151_, _26153_, _26154_);
  or g_57023_(_26138_, _26154_, _26155_);
  or g_57024_(_26131_, _26141_, _26156_);
  xor g_57025_(out[327], out[71], _26158_);
  or g_57026_(_26142_, _26158_, _26159_);
  or g_57027_(_26156_, _26159_, _26160_);
  or g_57028_(_26130_, _26132_, _26161_);
  or g_57029_(_26145_, _26161_, _26162_);
  or g_57030_(_26160_, _26162_, _26163_);
  or g_57031_(_26134_, _26163_, _26164_);
  or g_57032_(_26155_, _26164_, _26165_);
  not g_57033_(_26165_, _26166_);
  and g_57034_(out[331], _39537_, _26167_);
  xor g_57035_(out[324], out[52], _26169_);
  xor g_57036_(out[334], out[62], _26170_);
  or g_57037_(_26169_, _26170_, _26171_);
  xor g_57038_(out[333], out[61], _26172_);
  xor g_57039_(out[323], out[51], _26173_);
  xor g_57040_(out[320], out[48], _26174_);
  and g_57041_(_39427_, out[59], _26175_);
  xor g_57042_(out[330], out[58], _26176_);
  xor g_57043_(out[335], out[63], _26177_);
  xor g_57044_(out[326], out[54], _26178_);
  xor g_57045_(out[325], out[53], _26180_);
  xor g_57046_(out[328], out[56], _26181_);
  or g_57047_(_26172_, _26181_, _26182_);
  xor g_57048_(out[322], out[50], _26183_);
  xor g_57049_(out[329], out[57], _26184_);
  xor g_57050_(out[321], out[49], _26185_);
  or g_57051_(_26176_, _26183_, _26186_);
  or g_57052_(_26182_, _26186_, _26187_);
  or g_57053_(_26173_, _26184_, _26188_);
  or g_57054_(_26180_, _26188_, _26189_);
  or g_57055_(_26187_, _26189_, _26191_);
  or g_57056_(_26171_, _26191_, _26192_);
  xor g_57057_(out[332], out[60], _26193_);
  or g_57058_(_26175_, _26193_, _26194_);
  xor g_57059_(out[327], out[55], _26195_);
  or g_57060_(_26178_, _26195_, _26196_);
  or g_57061_(_26194_, _26196_, _26197_);
  or g_57062_(_26167_, _26185_, _26198_);
  or g_57063_(_26177_, _26198_, _26199_);
  or g_57064_(_26197_, _26199_, _26200_);
  or g_57065_(_26174_, _26200_, _26202_);
  or g_57066_(_26192_, _26202_, _26203_);
  xor g_57067_(out[329], out[41], _26204_);
  and g_57068_(out[327], _39515_, _26205_);
  xor g_57069_(out[330], out[42], _26206_);
  xor g_57070_(out[328], out[40], _26207_);
  xor g_57071_(out[324], out[36], _26208_);
  xor g_57072_(out[320], out[32], _26209_);
  xor g_57073_(out[331], out[43], _26210_);
  xor g_57074_(out[321], out[33], _26211_);
  and g_57075_(_39372_, out[39], _26213_);
  xor g_57076_(out[334], out[46], _26214_);
  xor g_57077_(out[326], out[38], _26215_);
  xor g_57078_(out[333], out[45], _26216_);
  xor g_57079_(out[332], out[44], _26217_);
  xor g_57080_(out[323], out[35], _26218_);
  or g_57081_(_26208_, _26218_, _26219_);
  xor g_57082_(out[325], out[37], _26220_);
  or g_57083_(_26206_, _26215_, _26221_);
  or g_57084_(_26219_, _26221_, _26222_);
  or g_57085_(_26210_, _26220_, _26224_);
  or g_57086_(_26216_, _26224_, _26225_);
  or g_57087_(_26222_, _26225_, _26226_);
  or g_57088_(_26209_, _26217_, _26227_);
  or g_57089_(_26226_, _26227_, _26228_);
  xor g_57090_(out[322], out[34], _26229_);
  or g_57091_(_26213_, _26229_, _26230_);
  xor g_57092_(out[335], out[47], _26231_);
  or g_57093_(_26214_, _26231_, _26232_);
  or g_57094_(_26230_, _26232_, _26233_);
  or g_57095_(_26204_, _26205_, _26235_);
  or g_57096_(_26211_, _26235_, _26236_);
  or g_57097_(_26233_, _26236_, _26237_);
  or g_57098_(_26207_, _26237_, _26238_);
  or g_57099_(_26228_, _26238_, _26239_);
  xor g_57100_(out[320], out[16], _26240_);
  xor g_57101_(out[329], out[25], _26241_);
  xor g_57102_(out[325], out[21], _26242_);
  and g_57103_(out[332], _39504_, _26243_);
  xor g_57104_(out[321], out[17], _26244_);
  xor g_57105_(out[327], out[23], _26246_);
  xor g_57106_(out[335], out[31], _26247_);
  xor g_57107_(out[326], out[22], _26248_);
  xor g_57108_(out[330], out[26], _26249_);
  xor g_57109_(out[322], out[18], _26250_);
  xor g_57110_(out[324], out[20], _26251_);
  xor g_57111_(out[334], out[30], _26252_);
  xor g_57112_(out[331], out[27], _26253_);
  xor g_57113_(out[323], out[19], _26254_);
  and g_57114_(_39449_, out[28], _26255_);
  or g_57115_(_26240_, _26250_, _26257_);
  or g_57116_(_26241_, _26252_, _26258_);
  or g_57117_(_26248_, _26253_, _26259_);
  or g_57118_(_26258_, _26259_, _26260_);
  or g_57119_(_26246_, _26249_, _26261_);
  or g_57120_(_26251_, _26254_, _26262_);
  or g_57121_(_26261_, _26262_, _26263_);
  or g_57122_(_26260_, _26263_, _26264_);
  xor g_57123_(out[333], out[29], _26265_);
  or g_57124_(_26255_, _26265_, _26266_);
  xor g_57125_(out[328], out[24], _26268_);
  or g_57126_(_26244_, _26268_, _26269_);
  or g_57127_(_26266_, _26269_, _26270_);
  or g_57128_(_26242_, _26243_, _26271_);
  or g_57129_(_26247_, _26271_, _26272_);
  or g_57130_(_26270_, _26272_, _26273_);
  or g_57131_(_26264_, _26273_, _26274_);
  or g_57132_(_26257_, _26274_, _26275_);
  xor g_57133_(_39295_, out[0], _26276_);
  xor g_57134_(_39328_, out[3], _26277_);
  xor g_57135_(_39405_, out[9], _26279_);
  or g_57136_(_39372_, out[7], _26280_);
  xor g_57137_(_39471_, out[14], _26281_);
  xor g_57138_(_39427_, out[11], _26282_);
  xor g_57139_(_39394_, out[8], _26283_);
  xor g_57140_(_39416_, out[10], _26284_);
  xor g_57141_(_39350_, out[5], _26285_);
  xor g_57142_(_39339_, out[4], _26286_);
  xor g_57143_(_39361_, out[6], _26287_);
  xor g_57144_(_39449_, out[12], _26288_);
  xor g_57145_(_39460_, out[13], _26290_);
  xor g_57146_(_39306_, out[1], _26291_);
  or g_57147_(out[327], _39383_, _26292_);
  and g_57148_(_26276_, _26288_, _26293_);
  and g_57149_(_26277_, _26286_, _26294_);
  and g_57150_(_26284_, _26287_, _26295_);
  and g_57151_(_26294_, _26295_, _26296_);
  and g_57152_(_26282_, _26285_, _26297_);
  and g_57153_(_26283_, _26290_, _26298_);
  and g_57154_(_26297_, _26298_, _26299_);
  and g_57155_(_26296_, _26299_, _26301_);
  xor g_57156_(_39317_, out[2], _26302_);
  and g_57157_(_26292_, _26302_, _26303_);
  xor g_57158_(_39482_, out[15], _26304_);
  and g_57159_(_26281_, _26304_, _26305_);
  and g_57160_(_26303_, _26305_, _26306_);
  and g_57161_(_26279_, _26280_, _26307_);
  and g_57162_(_26291_, _26307_, _26308_);
  and g_57163_(_26306_, _26308_, _26309_);
  and g_57164_(_26301_, _26309_, _26310_);
  and g_57165_(_26293_, _26310_, _26312_);
  not g_57166_(_26312_, _26313_);
  or g_57167_(_26275_, _26313_, _26314_);
  and g_57168_(_26275_, _26313_, _26315_);
  xor g_57169_(_26275_, _26312_, _26316_);
  xor g_57170_(_26239_, _26316_, _26317_);
  not g_57171_(_26317_, _26318_);
  or g_57172_(_26203_, _26318_, _26319_);
  xor g_57173_(_26203_, _26317_, _26320_);
  or g_57174_(_26165_, _26320_, _26321_);
  xor g_57175_(_26166_, _26320_, _26323_);
  not g_57176_(_26323_, _26324_);
  or g_57177_(_26129_, _26323_, _26325_);
  xor g_57178_(_26129_, _26323_, _26326_);
  xor g_57179_(_26129_, _26324_, _26327_);
  or g_57180_(_26093_, _26327_, _26328_);
  xor g_57181_(_26093_, _26326_, _26329_);
  not g_57182_(_26329_, _26330_);
  or g_57183_(_26056_, _26329_, _26331_);
  xor g_57184_(_26056_, _26329_, _26332_);
  xor g_57185_(_26056_, _26330_, _26334_);
  or g_57186_(_26020_, _26334_, _26335_);
  xor g_57187_(_26020_, _26332_, _26336_);
  or g_57188_(_25983_, _26336_, _26337_);
  not g_57189_(_26337_, _26338_);
  xor g_57190_(_25984_, _26336_, _26339_);
  not g_57191_(_26339_, _26340_);
  or g_57192_(_25946_, _26339_, _26341_);
  xor g_57193_(_25946_, _26339_, _26342_);
  xor g_57194_(_25946_, _26340_, _26343_);
  or g_57195_(_25910_, _26343_, _26345_);
  xor g_57196_(_25910_, _26342_, _26346_);
  or g_57197_(_25873_, _26346_, _26347_);
  xor g_57198_(_25874_, _26346_, _26348_);
  or g_57199_(_25835_, _26348_, _26349_);
  xor g_57200_(_25836_, _26348_, _26350_);
  not g_57201_(_26350_, _26351_);
  or g_57202_(_25799_, _26350_, _26352_);
  xor g_57203_(_25799_, _26350_, _26353_);
  xor g_57204_(_25799_, _26351_, _26354_);
  or g_57205_(_25763_, _26354_, _26356_);
  xor g_57206_(_25763_, _26353_, _26357_);
  or g_57207_(_25725_, _26357_, _26358_);
  xor g_57208_(_25726_, _26357_, _26359_);
  not g_57209_(_26359_, _26360_);
  or g_57210_(_25689_, _26359_, _26361_);
  xor g_57211_(_25689_, _26359_, _26362_);
  xor g_57212_(_25689_, _26360_, _26363_);
  or g_57213_(_25653_, _26363_, _26364_);
  xor g_57214_(_25653_, _26362_, _26365_);
  not g_57215_(_26365_, _26367_);
  or g_57216_(_25616_, _26365_, _26368_);
  xor g_57217_(_25616_, _26365_, _26369_);
  xor g_57218_(_25616_, _26367_, _26370_);
  or g_57219_(_25580_, _26370_, _26371_);
  xor g_57220_(_25580_, _26369_, _26372_);
  or g_57221_(_25543_, _26372_, _26373_);
  xor g_57222_(_25544_, _26372_, _26374_);
  not g_57223_(_26374_, _26375_);
  or g_57224_(_25506_, _26374_, _26376_);
  xor g_57225_(_25506_, _26374_, _26378_);
  xor g_57226_(_25506_, _26375_, _26379_);
  or g_57227_(_25470_, _26379_, _26380_);
  xor g_57228_(_25470_, _26378_, _26381_);
  not g_57229_(_26381_, _26382_);
  or g_57230_(_25434_, _26381_, _26383_);
  xor g_57231_(_25434_, _26381_, _26384_);
  xor g_57232_(_25434_, _26382_, _26385_);
  or g_57233_(_25397_, _26385_, _26386_);
  xor g_57234_(_25397_, _26384_, _26387_);
  or g_57235_(_25360_, _26387_, _26389_);
  xor g_57236_(_25361_, _26387_, _26390_);
  not g_57237_(_26390_, _26391_);
  or g_57238_(_25324_, _26390_, _26392_);
  xor g_57239_(_25324_, _26390_, _26393_);
  xor g_57240_(_25324_, _26391_, _26394_);
  or g_57241_(_25287_, _26394_, _26395_);
  xor g_57242_(_25287_, _26393_, _26396_);
  or g_57243_(_25250_, _26396_, _26397_);
  not g_57244_(_26397_, _26398_);
  xor g_57245_(_25251_, _26396_, _26400_);
  not g_57246_(_26400_, _26401_);
  or g_57247_(_25214_, _26400_, _26402_);
  not g_57248_(_26402_, _26403_);
  xor g_57249_(_25214_, _26400_, _26404_);
  xor g_57250_(_25214_, _26401_, _26405_);
  or g_57251_(_25177_, _26405_, _26406_);
  xor g_57252_(_25177_, _26404_, _26407_);
  or g_57253_(_25140_, _26407_, _26408_);
  xor g_57254_(_25141_, _26407_, _26409_);
  or g_57255_(_25103_, _26409_, _26411_);
  xor g_57256_(_25104_, _26409_, _26412_);
  not g_57257_(_26412_, _26413_);
  or g_57258_(_25066_, _26412_, _26414_);
  xor g_57259_(_25066_, _26412_, _26415_);
  xor g_57260_(_25066_, _26413_, _26416_);
  or g_57261_(_25030_, _26416_, _26417_);
  not g_57262_(_26417_, _26418_);
  xor g_57263_(_25030_, _26415_, _26419_);
  not g_57264_(_26419_, _26420_);
  or g_57265_(_24994_, _26419_, _26422_);
  xor g_57266_(_24994_, _26419_, _26423_);
  xor g_57267_(_24994_, _26420_, _26424_);
  or g_57268_(_24957_, _26424_, _26425_);
  xor g_57269_(_24957_, _26423_, _26426_);
  or g_57270_(_24920_, _26426_, _26427_);
  xor g_57271_(_24921_, _26426_, _26428_);
  or g_57272_(_24884_, _26428_, _26429_);
  xor g_57273_(_24884_, _26428_, _26430_);
  and g_57274_(_24847_, _26430_, _26431_);
  not g_57275_(_26431_, _26433_);
  xor g_57276_(_24846_, _26430_, _26434_);
  not g_57277_(_26434_, _26435_);
  or g_57278_(_24810_, _26434_, _26436_);
  xor g_57279_(_24810_, _26434_, _26437_);
  xor g_57280_(_24810_, _26435_, _26438_);
  or g_57281_(_24774_, _26438_, _26439_);
  xor g_57282_(_24774_, _26437_, _26440_);
  or g_57283_(_24736_, _26440_, _26441_);
  xor g_57284_(_24736_, _26440_, _26442_);
  xor g_57285_(_24737_, _26440_, _26444_);
  or g_57286_(_24700_, _26444_, _26445_);
  xor g_57287_(_24700_, _26442_, _26446_);
  not g_57288_(_26446_, _26447_);
  or g_57289_(_24664_, _26446_, _26448_);
  not g_57290_(_26448_, _26449_);
  xor g_57291_(_24664_, _26446_, _26450_);
  xor g_57292_(_24664_, _26447_, _26451_);
  or g_57293_(_24627_, _26451_, _26452_);
  xor g_57294_(_24627_, _26450_, _26453_);
  not g_57295_(_26453_, _26455_);
  or g_57296_(_24591_, _26453_, _26456_);
  xor g_57297_(_24591_, _26453_, _26457_);
  xor g_57298_(_24591_, _26455_, _26458_);
  or g_57299_(_24555_, _26458_, _26459_);
  xor g_57300_(_24555_, _26457_, _26460_);
  not g_57301_(_26460_, _26461_);
  or g_57302_(_24519_, _26460_, _26462_);
  xor g_57303_(_24519_, _26460_, _26463_);
  xor g_57304_(_24519_, _26461_, _26464_);
  or g_57305_(_24482_, _26464_, _26466_);
  xor g_57306_(_24482_, _26463_, _26467_);
  or g_57307_(_24445_, _26467_, _26468_);
  xor g_57308_(_24446_, _26467_, _26469_);
  not g_57309_(_26469_, _26470_);
  or g_57310_(_24409_, _26469_, _26471_);
  not g_57311_(_26471_, _26472_);
  xor g_57312_(_24409_, _26469_, _26473_);
  xor g_57313_(_24409_, _26470_, _26474_);
  or g_57314_(_24372_, _26474_, _26475_);
  not g_57315_(_26475_, _26477_);
  xor g_57316_(_24372_, _26473_, _26478_);
  or g_57317_(_24336_, _26478_, _26479_);
  xor g_57318_(_24336_, _26478_, _26480_);
  not g_57319_(_26480_, _26481_);
  or g_57320_(_24300_, _26481_, _26482_);
  xor g_57321_(_24300_, _26480_, _26483_);
  or g_57322_(_24263_, _26483_, _26484_);
  not g_57323_(_26484_, _26485_);
  and g_57324_(_24263_, _26483_, _26486_);
  xor g_57325_(_24263_, _26483_, _26488_);
  or g_57326_(_26485_, _26486_, _26489_);
  or g_57327_(_24227_, _26489_, _26490_);
  xor g_57328_(_24227_, _26488_, _26491_);
  or g_57329_(_24190_, _26491_, _26492_);
  xor g_57330_(_24191_, _26491_, _26493_);
  or g_57331_(_24152_, _26493_, _26494_);
  not g_57332_(_26494_, _26495_);
  xor g_57333_(_24153_, _26493_, _26496_);
  or g_57334_(_24116_, _26496_, _26497_);
  not g_57335_(_26497_, _26499_);
  and g_57336_(_24116_, _26496_, _26500_);
  xor g_57337_(_24116_, _26496_, _26501_);
  or g_57338_(_26499_, _26500_, _26502_);
  or g_57339_(_24080_, _26502_, _26503_);
  xor g_57340_(_24080_, _26501_, _26504_);
  or g_57341_(_24042_, _26504_, _26505_);
  xor g_57342_(_24043_, _26504_, _26506_);
  not g_57343_(_26506_, _26507_);
  or g_57344_(_24006_, _26506_, _26508_);
  xor g_57345_(_24006_, _26506_, _26510_);
  xor g_57346_(_24006_, _26507_, _26511_);
  or g_57347_(_23970_, _26511_, _26512_);
  xor g_57348_(_23970_, _26510_, _26513_);
  not g_57349_(_26513_, _26514_);
  or g_57350_(_23933_, _26513_, _26515_);
  xor g_57351_(_23933_, _26513_, _26516_);
  xor g_57352_(_23933_, _26514_, _26517_);
  or g_57353_(_23897_, _26517_, _26518_);
  xor g_57354_(_23897_, _26516_, _26519_);
  or g_57355_(_23860_, _26519_, _26521_);
  not g_57356_(_26521_, _26522_);
  xor g_57357_(_23861_, _26519_, _26523_);
  not g_57358_(_26523_, _26524_);
  or g_57359_(_23823_, _26523_, _26525_);
  xor g_57360_(_23823_, _26523_, _26526_);
  xor g_57361_(_23823_, _26524_, _26527_);
  or g_57362_(_23787_, _26527_, _26528_);
  xor g_57363_(_23787_, _26526_, _26529_);
  or g_57364_(_23750_, _26529_, _26530_);
  xor g_57365_(_23751_, _26529_, _26532_);
  not g_57366_(_26532_, _26533_);
  or g_57367_(_23713_, _26532_, _26534_);
  xor g_57368_(_23713_, _26532_, _26535_);
  xor g_57369_(_23713_, _26533_, _26536_);
  or g_57370_(_23677_, _26536_, _26537_);
  not g_57371_(_26537_, _26538_);
  xor g_57372_(_23677_, _26535_, _26539_);
  not g_57373_(_26539_, _26540_);
  or g_57374_(_23641_, _26539_, _26541_);
  xor g_57375_(_23641_, _26539_, _26543_);
  xor g_57376_(_23641_, _26540_, _26544_);
  or g_57377_(_23604_, _26544_, _26545_);
  xor g_57378_(_23604_, _26543_, _26546_);
  or g_57379_(_23567_, _26546_, _26547_);
  xor g_57380_(_23568_, _26546_, _26548_);
  not g_57381_(_26548_, _26549_);
  or g_57382_(_23531_, _26548_, _26550_);
  xor g_57383_(_23531_, _26548_, _26551_);
  xor g_57384_(_23531_, _26549_, _26552_);
  or g_57385_(_23494_, _26552_, _26554_);
  xor g_57386_(_23494_, _26551_, _26555_);
  or g_57387_(_23457_, _26555_, _26556_);
  xor g_57388_(_23458_, _26555_, _26557_);
  or g_57389_(_23421_, _26557_, _26558_);
  not g_57390_(_26558_, _26559_);
  xor g_57391_(_23421_, _26557_, _26560_);
  not g_57392_(_26560_, _26561_);
  or g_57393_(_23384_, _26561_, _26562_);
  xor g_57394_(_23384_, _26560_, _26563_);
  or g_57395_(_23348_, _26563_, _26565_);
  xor g_57396_(_23348_, _26563_, _26566_);
  not g_57397_(_26566_, _26567_);
  or g_57398_(_23312_, _26567_, _26568_);
  not g_57399_(_26568_, _26569_);
  xor g_57400_(_23312_, _26566_, _26570_);
  or g_57401_(_23274_, _26570_, _26571_);
  xor g_57402_(_23276_, _26570_, _26572_);
  or g_57403_(_23237_, _26572_, _26573_);
  not g_57404_(_26573_, _26574_);
  xor g_57405_(_23238_, _26572_, _26576_);
  not g_57406_(_26576_, _26577_);
  or g_57407_(_23201_, _26576_, _26578_);
  not g_57408_(_26578_, _26579_);
  xor g_57409_(_23201_, _26576_, _26580_);
  xor g_57410_(_23201_, _26577_, _26581_);
  or g_57411_(_23164_, _26581_, _26582_);
  xor g_57412_(_23164_, _26580_, _26583_);
  or g_57413_(_23128_, _26583_, _26584_);
  xor g_57414_(_23128_, _26583_, _26585_);
  not g_57415_(_26585_, _26587_);
  or g_57416_(_23092_, _26587_, _26588_);
  xor g_57417_(_23092_, _26585_, _26589_);
  not g_57418_(_26589_, _26590_);
  or g_57419_(_23056_, _26589_, _26591_);
  xor g_57420_(_23056_, _26589_, _26592_);
  xor g_57421_(_23056_, _26590_, _26593_);
  or g_57422_(_23019_, _26593_, _26594_);
  xor g_57423_(_23019_, _26592_, _26595_);
  or g_57424_(_22982_, _26595_, _26596_);
  xor g_57425_(_22983_, _26595_, _26598_);
  not g_57426_(_26598_, _26599_);
  or g_57427_(_22946_, _26598_, _26600_);
  xor g_57428_(_22946_, _26598_, _26601_);
  xor g_57429_(_22946_, _26599_, _26602_);
  or g_57430_(_22909_, _26602_, _26603_);
  xor g_57431_(_22909_, _26601_, _26604_);
  or g_57432_(_22873_, _26604_, _26605_);
  xor g_57433_(_22873_, _26604_, _26606_);
  not g_57434_(_26606_, _26607_);
  and g_57435_(_22837_, _26606_, _26609_);
  or g_57436_(_22836_, _26607_, _26610_);
  xor g_57437_(_22836_, _26606_, _26611_);
  or g_57438_(_22799_, _26611_, _26612_);
  xor g_57439_(_22799_, _26611_, _26613_);
  not g_57440_(_26613_, _26614_);
  or g_57441_(_22763_, _26614_, _26615_);
  xor g_57442_(_22763_, _26613_, _26616_);
  not g_57443_(_26616_, _26617_);
  or g_57444_(_22727_, _26616_, _26618_);
  xor g_57445_(_22727_, _26617_, _26620_);
  not g_57446_(_26620_, _26621_);
  or g_57447_(_22690_, _26620_, _26622_);
  xor g_57448_(_22690_, _26620_, _26623_);
  xor g_57449_(_22690_, _26621_, _26624_);
  or g_57450_(_22654_, _26624_, _26625_);
  not g_57451_(_26625_, _26626_);
  xor g_57452_(_22654_, _26623_, _26627_);
  or g_57453_(_22617_, _26627_, _26628_);
  xor g_57454_(_22618_, _26627_, _26629_);
  not g_57455_(_26629_, _26631_);
  or g_57456_(_22580_, _26629_, _26632_);
  xor g_57457_(_22580_, _26629_, _26633_);
  xor g_57458_(_22580_, _26631_, _26634_);
  or g_57459_(_22544_, _26634_, _26635_);
  not g_57460_(_26635_, _26636_);
  xor g_57461_(_22544_, _26633_, _26637_);
  not g_57462_(_26637_, _26638_);
  or g_57463_(_22508_, _26637_, _26639_);
  xor g_57464_(_22508_, _26637_, _26640_);
  xor g_57465_(_22508_, _26638_, _26642_);
  or g_57466_(_22471_, _26642_, _26643_);
  xor g_57467_(_22471_, _26640_, _26644_);
  not g_57468_(_26644_, _26645_);
  or g_57469_(_22435_, _26644_, _26646_);
  xor g_57470_(_22435_, _26644_, _26647_);
  xor g_57471_(_22435_, _26645_, _26648_);
  or g_57472_(_22399_, _26648_, _26649_);
  xor g_57473_(_22399_, _26647_, _26650_);
  or g_57474_(_22363_, _26650_, _26651_);
  xor g_57475_(_22363_, _26650_, _26653_);
  not g_57476_(_26653_, _26654_);
  or g_57477_(_22326_, _26654_, _26655_);
  xor g_57478_(_22326_, _26653_, _26656_);
  or g_57479_(_22290_, _26656_, _26657_);
  xor g_57480_(_22290_, _26656_, _26658_);
  not g_57481_(_26658_, _26659_);
  or g_57482_(_22254_, _26659_, _26660_);
  xor g_57483_(_22254_, _26658_, _26661_);
  or g_57484_(_22216_, _26661_, _26662_);
  xor g_57485_(_22217_, _26661_, _26664_);
  not g_57486_(_26664_, _26665_);
  or g_57487_(_22180_, _26664_, _26666_);
  xor g_57488_(_22180_, _26664_, _26667_);
  xor g_57489_(_22180_, _26665_, _26668_);
  or g_57490_(_22144_, _26668_, _26669_);
  xor g_57491_(_22144_, _26667_, _26670_);
  or g_57492_(_22106_, _26670_, _26671_);
  xor g_57493_(_22107_, _26670_, _26672_);
  or g_57494_(_22070_, _26672_, _26673_);
  xor g_57495_(_22070_, _26672_, _26675_);
  not g_57496_(_26675_, _26676_);
  and g_57497_(_22034_, _26675_, _26677_);
  or g_57498_(_22033_, _26676_, _26678_);
  xor g_57499_(_22033_, _26675_, _26679_);
  or g_57500_(_21995_, _26679_, _26680_);
  not g_57501_(_26680_, _26681_);
  xor g_57502_(_21996_, _26679_, _26682_);
  or g_57503_(_21958_, _26682_, _26683_);
  xor g_57504_(_21959_, _26682_, _26684_);
  not g_57505_(_26684_, _26686_);
  or g_57506_(_21921_, _26684_, _26687_);
  xor g_57507_(_21921_, _26684_, _26688_);
  xor g_57508_(_21921_, _26686_, _26689_);
  or g_57509_(_43141_, _26689_, _26690_);
  xor g_57510_(_43141_, _26688_, _26691_);
  or g_57511_(_43104_, _26691_, _26692_);
  xor g_57512_(_43105_, _26691_, _26693_);
  not g_57513_(_26693_, _26694_);
  or g_57514_(_43067_, _26693_, _26695_);
  xor g_57515_(_43067_, _26693_, _26697_);
  xor g_57516_(_43067_, _26694_, _26698_);
  or g_57517_(_43031_, _26698_, _26699_);
  not g_57518_(_26699_, _26700_);
  xor g_57519_(_43031_, _26697_, _26701_);
  or g_57520_(_42994_, _26701_, _26702_);
  not g_57521_(_26702_, _26703_);
  xor g_57522_(_42995_, _26701_, _26704_);
  or g_57523_(_42956_, _26704_, _26705_);
  xor g_57524_(_42957_, _26704_, _26706_);
  not g_57525_(_26706_, _26708_);
  or g_57526_(_42920_, _26706_, _26709_);
  xor g_57527_(_42920_, _26706_, _26710_);
  xor g_57528_(_42920_, _26708_, _26711_);
  or g_57529_(_42884_, _26711_, _26712_);
  xor g_57530_(_42884_, _26710_, _26713_);
  not g_57531_(_26713_, _26714_);
  or g_57532_(_42847_, _26713_, _26715_);
  xor g_57533_(_42847_, _26713_, _26716_);
  xor g_57534_(_42847_, _26714_, _26717_);
  or g_57535_(_42811_, _26717_, _26719_);
  xor g_57536_(_42811_, _26716_, _26720_);
  or g_57537_(_42774_, _26720_, _26721_);
  xor g_57538_(_42775_, _26720_, _26722_);
  or g_57539_(_42736_, _26722_, _26723_);
  xor g_57540_(_42736_, _26722_, _26724_);
  xor g_57541_(_42737_, _26722_, _26725_);
  or g_57542_(_42700_, _26725_, _26726_);
  xor g_57543_(_42700_, _26724_, _26727_);
  or g_57544_(_42663_, _26727_, _26728_);
  xor g_57545_(_42664_, _26727_, _26730_);
  or g_57546_(_42625_, _26730_, _26731_);
  xor g_57547_(_42626_, _26730_, _26732_);
  or g_57548_(_42589_, _26732_, _26733_);
  xor g_57549_(_42589_, _26732_, _26734_);
  not g_57550_(_26734_, _26735_);
  or g_57551_(_42553_, _26735_, _26736_);
  not g_57552_(_26736_, _26737_);
  xor g_57553_(_42553_, _26734_, _26738_);
  or g_57554_(_42515_, _26738_, _26739_);
  not g_57555_(_26739_, _26741_);
  xor g_57556_(_42516_, _26738_, _26742_);
  not g_57557_(_26742_, _26743_);
  or g_57558_(_42479_, _26742_, _26744_);
  xor g_57559_(_42479_, _26742_, _26745_);
  xor g_57560_(_42479_, _26743_, _26746_);
  or g_57561_(_42443_, _26746_, _26747_);
  xor g_57562_(_42443_, _26745_, _26748_);
  or g_57563_(_42406_, _26748_, _26749_);
  not g_57564_(_26749_, _26750_);
  and g_57565_(_42406_, _26748_, _26752_);
  xor g_57566_(_42406_, _26748_, _26753_);
  or g_57567_(_26750_, _26752_, _26754_);
  or g_57568_(_42370_, _26754_, _26755_);
  not g_57569_(_26755_, _26756_);
  xor g_57570_(_42370_, _26753_, _26757_);
  or g_57571_(_42333_, _26757_, _26758_);
  not g_57572_(_26758_, _26759_);
  xor g_57573_(_42334_, _26757_, _26760_);
  or g_57574_(_42295_, _26760_, _26761_);
  xor g_57575_(_42296_, _26760_, _26763_);
  not g_57576_(_26763_, _26764_);
  or g_57577_(_42259_, _26763_, _26765_);
  xor g_57578_(_42259_, _26763_, _26766_);
  xor g_57579_(_42259_, _26764_, _26767_);
  or g_57580_(_42223_, _26767_, _26768_);
  xor g_57581_(_42223_, _26766_, _26769_);
  or g_57582_(_42186_, _26769_, _26770_);
  xor g_57583_(_42186_, _26769_, _26771_);
  not g_57584_(_26771_, _26772_);
  or g_57585_(_42150_, _26772_, _26774_);
  xor g_57586_(_42150_, _26771_, _26775_);
  or g_57587_(_42113_, _26775_, _26776_);
  xor g_57588_(_42114_, _26775_, _26777_);
  not g_57589_(_26777_, _26778_);
  or g_57590_(_42076_, _26777_, _26779_);
  xor g_57591_(_42076_, _26777_, _26780_);
  xor g_57592_(_42076_, _26778_, _26781_);
  or g_57593_(_42040_, _26781_, _26782_);
  not g_57594_(_26782_, _26783_);
  xor g_57595_(_42040_, _26780_, _26785_);
  or g_57596_(_42004_, _26785_, _26786_);
  not g_57597_(_26786_, _26787_);
  and g_57598_(_42004_, _26785_, _26788_);
  xor g_57599_(_42004_, _26785_, _26789_);
  or g_57600_(_26787_, _26788_, _26790_);
  or g_57601_(_41967_, _26790_, _26791_);
  xor g_57602_(_41967_, _26789_, _26792_);
  not g_57603_(_26792_, _26793_);
  or g_57604_(_41931_, _26792_, _26794_);
  xor g_57605_(_41931_, _26792_, _26796_);
  xor g_57606_(_41931_, _26793_, _26797_);
  or g_57607_(_41895_, _26797_, _26798_);
  xor g_57608_(_41895_, _26796_, _26799_);
  not g_57609_(_26799_, _26800_);
  or g_57610_(_41859_, _26799_, _26801_);
  xor g_57611_(_41859_, _26799_, _26802_);
  xor g_57612_(_41859_, _26800_, _26803_);
  or g_57613_(_41822_, _26803_, _26804_);
  xor g_57614_(_41822_, _26802_, _26805_);
  or g_57615_(_41785_, _26805_, _26807_);
  xor g_57616_(_41786_, _26805_, _26808_);
  not g_57617_(_26808_, _26809_);
  or g_57618_(_41749_, _26808_, _26810_);
  xor g_57619_(_41749_, _26808_, _26811_);
  xor g_57620_(_41749_, _26809_, _26812_);
  or g_57621_(_41712_, _26812_, _26813_);
  xor g_57622_(_41712_, _26811_, _26814_);
  or g_57623_(_41676_, _26814_, _26815_);
  xor g_57624_(_41676_, _26814_, _26816_);
  not g_57625_(_26816_, _26818_);
  or g_57626_(_41640_, _26818_, _26819_);
  xor g_57627_(_41640_, _26816_, _26820_);
  or g_57628_(_41602_, _26820_, _26821_);
  xor g_57629_(_41603_, _26820_, _26822_);
  or g_57630_(_41565_, _26822_, _26823_);
  xor g_57631_(_41566_, _26822_, _26824_);
  not g_57632_(_26824_, _26825_);
  or g_57633_(_41529_, _26824_, _26826_);
  xor g_57634_(_41529_, _26824_, _26827_);
  xor g_57635_(_41529_, _26825_, _26829_);
  or g_57636_(_41492_, _26829_, _26830_);
  xor g_57637_(_41492_, _26827_, _26831_);
  not g_57638_(_26831_, _26832_);
  or g_57639_(_41456_, _26831_, _26833_);
  xor g_57640_(_41456_, _26831_, _26834_);
  xor g_57641_(_41456_, _26832_, _26835_);
  or g_57642_(_41420_, _26835_, _26836_);
  xor g_57643_(_41420_, _26834_, _26837_);
  or g_57644_(_41382_, _26837_, _26838_);
  xor g_57645_(_41383_, _26837_, _26840_);
  or g_57646_(_41345_, _26840_, _26841_);
  not g_57647_(_26841_, _26842_);
  xor g_57648_(_41346_, _26840_, _26843_);
  or g_57649_(_41309_, _26843_, _26844_);
  not g_57650_(_26844_, _26845_);
  and g_57651_(_41309_, _26843_, _26846_);
  xor g_57652_(_41309_, _26843_, _26847_);
  or g_57653_(_26845_, _26846_, _26848_);
  or g_57654_(_41272_, _26848_, _26849_);
  xor g_57655_(_41272_, _26847_, _26851_);
  or g_57656_(_41235_, _26851_, _26852_);
  xor g_57657_(_41236_, _26851_, _26853_);
  or g_57658_(_41197_, _26853_, _26854_);
  not g_57659_(_26854_, _26855_);
  xor g_57660_(_41199_, _26853_, _26856_);
  not g_57661_(_26856_, _26857_);
  or g_57662_(_41161_, _26856_, _26858_);
  xor g_57663_(_41161_, _26856_, _26859_);
  xor g_57664_(_41161_, _26857_, _26860_);
  or g_57665_(_41125_, _26860_, _26862_);
  xor g_57666_(_41125_, _26859_, _26863_);
  not g_57667_(_26863_, _26864_);
  or g_57668_(_41089_, _26863_, _26865_);
  xor g_57669_(_41089_, _26863_, _26866_);
  xor g_57670_(_41089_, _26864_, _26867_);
  or g_57671_(_41052_, _26867_, _26868_);
  xor g_57672_(_41052_, _26866_, _26869_);
  or g_57673_(_41015_, _26869_, _26870_);
  xor g_57674_(_41016_, _26869_, _26871_);
  or g_57675_(_40979_, _26871_, _26873_);
  not g_57676_(_26873_, _26874_);
  and g_57677_(_40979_, _26871_, _26875_);
  xor g_57678_(_40979_, _26871_, _26876_);
  or g_57679_(_26874_, _26875_, _26877_);
  or g_57680_(_40942_, _26877_, _26878_);
  xor g_57681_(_40942_, _26876_, _26879_);
  or g_57682_(_40905_, _26879_, _26880_);
  xor g_57683_(_40906_, _26879_, _26881_);
  or g_57684_(_40867_, _26881_, _26882_);
  xor g_57685_(_40869_, _26881_, _26884_);
  not g_57686_(_26884_, _26885_);
  or g_57687_(_40831_, _26884_, _26886_);
  xor g_57688_(_40831_, _26884_, _26887_);
  xor g_57689_(_40831_, _26885_, _26888_);
  or g_57690_(_40795_, _26888_, _26889_);
  xor g_57691_(_40795_, _26887_, _26890_);
  or g_57692_(_40757_, _26890_, _26891_);
  xor g_57693_(_40759_, _26890_, _26892_);
  or g_57694_(_40720_, _26892_, _26893_);
  xor g_57695_(_40721_, _26892_, _26895_);
  not g_57696_(_26895_, _26896_);
  or g_57697_(_40684_, _26895_, _26897_);
  xor g_57698_(_40684_, _26895_, _26898_);
  xor g_57699_(_40684_, _26896_, _26899_);
  or g_57700_(_40647_, _26899_, _26900_);
  xor g_57701_(_40647_, _26898_, _26901_);
  or g_57702_(_40610_, _26901_, _26902_);
  xor g_57703_(_40611_, _26901_, _26903_);
  or g_57704_(_40573_, _26903_, _26904_);
  xor g_57705_(_40574_, _26903_, _26906_);
  not g_57706_(_26906_, _26907_);
  or g_57707_(_40536_, _26906_, _26908_);
  xor g_57708_(_40536_, _26906_, _26909_);
  xor g_57709_(_40536_, _26907_, _26910_);
  or g_57710_(_40500_, _26910_, _26911_);
  xor g_57711_(_40500_, _26909_, _26912_);
  not g_57712_(_26912_, _26913_);
  or g_57713_(_40464_, _26912_, _26914_);
  xor g_57714_(_40464_, _26912_, _26915_);
  xor g_57715_(_40464_, _26913_, _26917_);
  or g_57716_(_40427_, _26917_, _26918_);
  xor g_57717_(_40427_, _26915_, _26919_);
  or g_57718_(_40391_, _26919_, _26920_);
  xor g_57719_(_40391_, _26919_, _26921_);
  not g_57720_(_26921_, _26922_);
  or g_57721_(_40355_, _26922_, _26923_);
  not g_57722_(_26923_, _26924_);
  xor g_57723_(_40355_, _26921_, _26925_);
  or g_57724_(_40317_, _26925_, _26926_);
  xor g_57725_(_40319_, _26925_, _26928_);
  not g_57726_(_26928_, _26929_);
  or g_57727_(_40281_, _26928_, _26930_);
  xor g_57728_(_40281_, _26928_, _26931_);
  xor g_57729_(_40281_, _26929_, _26932_);
  or g_57730_(_40245_, _26932_, _26933_);
  xor g_57731_(_40245_, _26931_, _26934_);
  or g_57732_(_40207_, _26934_, _26935_);
  xor g_57733_(_40209_, _26934_, _26936_);
  or g_57734_(_40170_, _26936_, _26937_);
  xor g_57735_(_40171_, _26936_, _26939_);
  or g_57736_(_40133_, _26939_, _26940_);
  not g_57737_(_26940_, _26941_);
  xor g_57738_(_40134_, _26939_, _26942_);
  or g_57739_(_40095_, _26942_, _26943_);
  xor g_57740_(_40096_, _26942_, _26944_);
  or g_57741_(_40058_, _26944_, _26945_);
  xor g_57742_(_40059_, _26944_, _26946_);
  or g_57743_(_40020_, _26946_, _26947_);
  xor g_57744_(_40022_, _26946_, _26948_);
  or g_57745_(_39984_, _26948_, _26950_);
  xor g_57746_(_39984_, _26948_, _26951_);
  and g_57747_(_39948_, _26951_, _26952_);
  not g_57748_(_26952_, _26953_);
  xor g_57749_(_39947_, _26951_, _26954_);
  not g_57750_(_26954_, _26955_);
  or g_57751_(_39910_, _26954_, _26956_);
  xor g_57752_(_39910_, _26954_, _26957_);
  xor g_57753_(_39910_, _26955_, _26958_);
  or g_57754_(_39874_, _26958_, _26959_);
  xor g_57755_(_39874_, _26957_, _26961_);
  or g_57756_(_39837_, _26961_, _26962_);
  xor g_57757_(_39838_, _26961_, _26963_);
  not g_57758_(_26963_, _26964_);
  or g_57759_(_39800_, _26963_, _26965_);
  xor g_57760_(_39800_, _26963_, _26966_);
  xor g_57761_(_39800_, _26964_, _26967_);
  or g_57762_(_39764_, _26967_, _26968_);
  xor g_57763_(_39764_, _26966_, _26969_);
  or g_57764_(_39727_, _26969_, _26970_);
  xor g_57765_(_39728_, _26969_, _26972_);
  or g_57766_(_39689_, _26972_, _26973_);
  xor g_57767_(_39690_, _26972_, _26974_);
  not g_57768_(_26974_, _26975_);
  or g_57769_(_39653_, _26974_, _26976_);
  xor g_57770_(_39653_, _26974_, _26977_);
  xor g_57771_(_39653_, _26975_, _26978_);
  or g_57772_(_39617_, _26978_, _26979_);
  xor g_57773_(_39617_, _26977_, _26980_);
  or g_57774_(_39579_, _26980_, _26981_);
  xor g_57775_(_39580_, _26980_, _26983_);
  not g_57776_(_26983_, _26984_);
  or g_57777_(_39543_, _26983_, _26985_);
  xor g_57778_(_39543_, _26983_, _26986_);
  xor g_57779_(_39543_, _26984_, _26987_);
  or g_57780_(_39507_, _26987_, _26988_);
  xor g_57781_(_39507_, _26986_, _26989_);
  or g_57782_(_39470_, _26989_, _26990_);
  not g_57783_(_26990_, _26991_);
  and g_57784_(_39470_, _26989_, _26992_);
  xor g_57785_(_39470_, _26989_, _26994_);
  or g_57786_(_26991_, _26992_, _26995_);
  or g_57787_(_39434_, _26995_, _26996_);
  xor g_57788_(_39434_, _26994_, _26997_);
  or g_57789_(_39397_, _26997_, _26998_);
  xor g_57790_(_39398_, _26997_, _26999_);
  or g_57791_(_39359_, _26999_, _27000_);
  xor g_57792_(_39360_, _26999_, _27001_);
  or g_57793_(_39322_, _27001_, _27002_);
  xor g_57794_(_39322_, _27001_, _27003_);
  xor g_57795_(_39323_, _27001_, _27005_);
  or g_57796_(_39286_, _27005_, _27006_);
  xor g_57797_(_39286_, _27003_, _27007_);
  or g_57798_(_39252_, _27007_, _27008_);
  xor g_57799_(_39253_, _27007_, _27009_);
  or g_57800_(_39218_, _27009_, _27010_);
  not g_57801_(_27010_, _27011_);
  xor g_57802_(_39219_, _27009_, _27012_);
  or g_57803_(_39184_, _27012_, _27013_);
  xor g_57804_(_39184_, _27012_, _27014_);
  xor g_57805_(_39185_, _27012_, _27016_);
  or g_57806_(_39151_, _27016_, _27017_);
  xor g_57807_(_39151_, _27014_, _27018_);
  or g_57808_(_39117_, _27018_, _27019_);
  not g_57809_(_27019_, _27020_);
  xor g_57810_(_39118_, _27018_, _27021_);
  or g_57811_(_39083_, _27021_, _27022_);
  xor g_57812_(_39083_, _27021_, _27023_);
  xor g_57813_(_39084_, _27021_, _27024_);
  or g_57814_(_39050_, _27024_, _27025_);
  xor g_57815_(_39050_, _27023_, _27027_);
  not g_57816_(_27027_, _27028_);
  or g_57817_(_39017_, _27027_, _27029_);
  xor g_57818_(_39017_, _27028_, _27030_);
  or g_57819_(_38983_, _27030_, _27031_);
  not g_57820_(_27031_, _27032_);
  xor g_57821_(_38984_, _27030_, _27033_);
  or g_57822_(_38950_, _27033_, _27034_);
  not g_57823_(_27034_, _27035_);
  xor g_57824_(_38950_, _27033_, _27036_);
  not g_57825_(_27036_, _27038_);
  and g_57826_(_38917_, _27036_, _27039_);
  or g_57827_(_38916_, _27038_, _27040_);
  xor g_57828_(_38916_, _27036_, _27041_);
  not g_57829_(_27041_, _27042_);
  or g_57830_(_38883_, _27041_, _27043_);
  xor g_57831_(_38883_, _27041_, _27044_);
  xor g_57832_(_38883_, _27042_, _27045_);
  or g_57833_(_38850_, _27045_, _27046_);
  xor g_57834_(_38850_, _27044_, _27047_);
  or g_57835_(_38816_, _27047_, _27049_);
  xor g_57836_(_38817_, _27047_, _27050_);
  not g_57837_(_27050_, _27051_);
  or g_57838_(_38783_, _27050_, _27052_);
  xor g_57839_(_38783_, _27050_, _27053_);
  xor g_57840_(_38783_, _27051_, _27054_);
  or g_57841_(_38750_, _27054_, _27055_);
  xor g_57842_(_38750_, _27053_, _27056_);
  or g_57843_(_38717_, _27056_, _27057_);
  not g_57844_(_27057_, _27058_);
  and g_57845_(_38717_, _27056_, _27060_);
  xor g_57846_(_38717_, _27056_, _27061_);
  or g_57847_(_27058_, _27060_, _27062_);
  or g_57848_(_38684_, _27062_, _27063_);
  xor g_57849_(_38684_, _27061_, _27064_);
  or g_57850_(_38650_, _27064_, _27065_);
  xor g_57851_(_38651_, _27064_, _27066_);
  or g_57852_(_38616_, _27066_, _27067_);
  xor g_57853_(_38617_, _27066_, _27068_);
  or g_57854_(_38583_, _27068_, _27069_);
  not g_57855_(_27069_, _27071_);
  and g_57856_(_38583_, _27068_, _27072_);
  or g_57857_(_27071_, _27072_, _27073_);
  not g_57858_(_27073_, _27074_);
  or g_57859_(_38550_, _27073_, _27075_);
  or g_57860_(_38550_, _27072_, _27076_);
  xor g_57861_(_38550_, _27073_, _27077_);
  xor g_57862_(_38550_, _27074_, _27078_);
  or g_57863_(_38517_, _27078_, _27079_);
  xor g_57864_(_38517_, _27077_, _27080_);
  or g_57865_(_38483_, _27080_, _27082_);
  xor g_57866_(_38484_, _27080_, _27083_);
  or g_57867_(_38449_, _27083_, _27084_);
  xor g_57868_(_38450_, _27083_, _27085_);
  not g_57869_(_27085_, _27086_);
  or g_57870_(_38416_, _27085_, _27087_);
  xor g_57871_(_38416_, _27085_, _27088_);
  xor g_57872_(_38416_, _27086_, _27089_);
  or g_57873_(_38383_, _27089_, _27090_);
  xor g_57874_(_38383_, _27088_, _27091_);
  or g_57875_(_38350_, _27091_, _27093_);
  xor g_57876_(_38350_, _27091_, _27094_);
  not g_57877_(_27094_, _27095_);
  or g_57878_(_38317_, _27095_, _27096_);
  xor g_57879_(_38317_, _27094_, _27097_);
  or g_57880_(_38284_, _27097_, _27098_);
  not g_57881_(_27098_, _27099_);
  xor g_57882_(_38284_, _27097_, _27100_);
  not g_57883_(_27100_, _27101_);
  or g_57884_(_38251_, _27101_, _27102_);
  xor g_57885_(_38251_, _27100_, _27104_);
  not g_57886_(_27104_, _27105_);
  or g_57887_(_38218_, _27104_, _27106_);
  xor g_57888_(_38218_, _27104_, _27107_);
  xor g_57889_(_38218_, _27105_, _27108_);
  or g_57890_(_38185_, _27108_, _27109_);
  xor g_57891_(_38185_, _27107_, _27110_);
  not g_57892_(_27110_, _27111_);
  or g_57893_(_38152_, _27110_, _27112_);
  xor g_57894_(_38152_, _27110_, _27113_);
  xor g_57895_(_38152_, _27111_, _27115_);
  or g_57896_(_38119_, _27115_, _27116_);
  xor g_57897_(_38119_, _27113_, _27117_);
  not g_57898_(_27117_, _27118_);
  or g_57899_(_38086_, _27117_, _27119_);
  xor g_57900_(_38086_, _27117_, _27120_);
  xor g_57901_(_38086_, _27118_, _27121_);
  or g_57902_(_38053_, _27121_, _27122_);
  xor g_57903_(_38053_, _27120_, _27123_);
  not g_57904_(_27123_, _27124_);
  or g_57905_(_38020_, _27123_, _27126_);
  xor g_57906_(_38020_, _27123_, _27127_);
  xor g_57907_(_38020_, _27124_, _27128_);
  or g_57908_(_37987_, _27128_, _27129_);
  xor g_57909_(_37987_, _27127_, _27130_);
  not g_57910_(_27130_, _27131_);
  or g_57911_(_37954_, _27130_, _27132_);
  xor g_57912_(_37954_, _27131_, _27133_);
  not g_57913_(_27133_, _27134_);
  or g_57914_(_37921_, _27133_, _27135_);
  xor g_57915_(_37921_, _27134_, _27137_);
  or g_57916_(_37888_, _27137_, _27138_);
  xor g_57917_(_37888_, _27137_, _27139_);
  not g_57918_(_27139_, _27140_);
  or g_57919_(_37855_, _27140_, _27141_);
  xor g_57920_(_37855_, _27139_, _27142_);
  not g_57921_(_27142_, _27143_);
  or g_57922_(_37822_, _27142_, _27144_);
  xor g_57923_(_37822_, _27142_, _27145_);
  xor g_57924_(_37822_, _27143_, _27146_);
  or g_57925_(_37789_, _27146_, _27148_);
  xor g_57926_(_37789_, _27145_, _27149_);
  or g_57927_(_37756_, _27149_, _27150_);
  xor g_57928_(_37756_, _27149_, _27151_);
  not g_57929_(_27151_, _27152_);
  or g_57930_(_37723_, _27152_, _27153_);
  xor g_57931_(_37723_, _27151_, _27154_);
  not g_57932_(_27154_, _27155_);
  or g_57933_(_37690_, _27154_, _27156_);
  xor g_57934_(_37690_, _27154_, _27157_);
  xor g_57935_(_37690_, _27155_, _27159_);
  or g_57936_(_37657_, _27159_, _27160_);
  xor g_57937_(_37657_, _27157_, _27161_);
  or g_57938_(_37624_, _27161_, _27162_);
  xor g_57939_(_37624_, _27161_, _27163_);
  not g_57940_(_27163_, _27164_);
  or g_57941_(_37591_, _27164_, _27165_);
  xor g_57942_(_37591_, _27163_, _27166_);
  not g_57943_(_27166_, _27167_);
  or g_57944_(_37558_, _27166_, _27168_);
  xor g_57945_(_37558_, _27167_, _27170_);
  not g_57946_(_27170_, _27171_);
  or g_57947_(_37525_, _27170_, _27172_);
  not g_57948_(_27172_, _27173_);
  xor g_57949_(_37525_, _27170_, _27174_);
  xor g_57950_(_37525_, _27171_, _27175_);
  or g_57951_(_37492_, _27175_, _27176_);
  xor g_57952_(_37492_, _27174_, _27177_);
  not g_57953_(_27177_, _27178_);
  or g_57954_(_37459_, _27177_, _27179_);
  xor g_57955_(_37459_, _27177_, _27181_);
  xor g_57956_(_37459_, _27178_, _27182_);
  or g_57957_(_37426_, _27182_, _27183_);
  xor g_57958_(_37426_, _27181_, _27184_);
  not g_57959_(_27184_, _27185_);
  or g_57960_(_37393_, _27184_, _27186_);
  xor g_57961_(_37393_, _27185_, _27187_);
  or g_57962_(_37359_, _27187_, _27188_);
  not g_57963_(_27188_, _27189_);
  xor g_57964_(_37360_, _27187_, _27190_);
  or g_57965_(_37325_, _27190_, _27192_);
  xor g_57966_(_37325_, _27190_, _27193_);
  xor g_57967_(_37326_, _27190_, _27194_);
  or g_57968_(_37292_, _27194_, _27195_);
  not g_57969_(_27195_, _27196_);
  xor g_57970_(_37292_, _27193_, _27197_);
  not g_57971_(_27197_, _27198_);
  or g_57972_(_37259_, _27197_, _27199_);
  xor g_57973_(_37259_, _27198_, _27200_);
  or g_57974_(_37225_, _27200_, _27201_);
  xor g_57975_(_37226_, _27200_, _27203_);
  not g_57976_(_27203_, _27204_);
  or g_57977_(_37192_, _27203_, _27205_);
  xor g_57978_(_37192_, _27203_, _27206_);
  xor g_57979_(_37192_, _27204_, _27207_);
  or g_57980_(_37159_, _27207_, _27208_);
  not g_57981_(_27208_, _27209_);
  xor g_57982_(_37159_, _27206_, _27210_);
  or g_57983_(_37125_, _27210_, _27211_);
  xor g_57984_(_37126_, _27210_, _27212_);
  or g_57985_(_37091_, _27212_, _27214_);
  xor g_57986_(_37091_, _27212_, _27215_);
  xor g_57987_(_37092_, _27212_, _27216_);
  and g_57988_(_37058_, _27215_, _27217_);
  or g_57989_(_37057_, _27216_, _27218_);
  xor g_57990_(_37058_, _27215_, _27219_);
  xor g_57991_(_37057_, _27215_, _27220_);
  or g_57992_(_37024_, _27220_, _27221_);
  xor g_57993_(_37024_, _27219_, _27222_);
  not g_57994_(_27222_, _27223_);
  or g_57995_(_36991_, _27222_, _27225_);
  xor g_57996_(_36991_, _27222_, _27226_);
  xor g_57997_(_36991_, _27223_, _27227_);
  or g_57998_(_36958_, _27227_, _27228_);
  xor g_57999_(_36958_, _27226_, _27229_);
  or g_58000_(_36924_, _27229_, _27230_);
  xor g_58001_(_36925_, _27229_, _27231_);
  not g_58002_(_27231_, _27232_);
  or g_58003_(_36891_, _27231_, _27233_);
  xor g_58004_(_36891_, _27231_, _27234_);
  xor g_58005_(_36891_, _27232_, _27236_);
  or g_58006_(_36858_, _27236_, _27237_);
  xor g_58007_(_36858_, _27234_, _27238_);
  or g_58008_(_36825_, _27238_, _27239_);
  xor g_58009_(_36825_, _27238_, _27240_);
  not g_58010_(_27240_, _27241_);
  or g_58011_(_36792_, _27241_, _27242_);
  xor g_58012_(_36792_, _27240_, _27243_);
  not g_58013_(_27243_, _27244_);
  or g_58014_(_36759_, _27243_, _27245_);
  xor g_58015_(_36759_, _27244_, _27247_);
  not g_58016_(_27247_, _27248_);
  or g_58017_(_36726_, _27247_, _27249_);
  xor g_58018_(_36726_, _27247_, _27250_);
  xor g_58019_(_36726_, _27248_, _27251_);
  or g_58020_(_36693_, _27251_, _27252_);
  not g_58021_(_27252_, _27253_);
  xor g_58022_(_36693_, _27250_, _27254_);
  or g_58023_(_36660_, _27254_, _27255_);
  xor g_58024_(_36660_, _27254_, _27256_);
  not g_58025_(_27256_, _27258_);
  or g_58026_(_36627_, _27258_, _27259_);
  xor g_58027_(_36627_, _27256_, _27260_);
  not g_58028_(_27260_, _27261_);
  or g_58029_(_36594_, _27260_, _27262_);
  xor g_58030_(_36594_, _27260_, _27263_);
  xor g_58031_(_36594_, _27261_, _27264_);
  or g_58032_(_36561_, _27264_, _27265_);
  xor g_58033_(_36561_, _27263_, _27266_);
  not g_58034_(_27266_, _27267_);
  or g_58035_(_36528_, _27266_, _27269_);
  xor g_58036_(_36528_, _27267_, _27270_);
  or g_58037_(_36495_, _27270_, _27271_);
  xor g_58038_(_36495_, _27270_, _27272_);
  not g_58039_(_27272_, _27273_);
  or g_58040_(_36462_, _27273_, _27274_);
  xor g_58041_(_36462_, _27272_, _27275_);
  or g_58042_(_36428_, _27275_, _27276_);
  xor g_58043_(_36428_, _27275_, _27277_);
  xor g_58044_(_36429_, _27275_, _27278_);
  or g_58045_(_36395_, _27278_, _27280_);
  xor g_58046_(_36395_, _27277_, _27281_);
  or g_58047_(_36362_, _27281_, _27282_);
  not g_58048_(_27282_, _27283_);
  xor g_58049_(_36362_, _27281_, _27284_);
  not g_58050_(_27284_, _27285_);
  and g_58051_(_36329_, _27284_, _27286_);
  or g_58052_(_36328_, _27285_, _27287_);
  xor g_58053_(_36328_, _27284_, _27288_);
  or g_58054_(_36294_, _27288_, _27289_);
  not g_58055_(_27289_, _27291_);
  xor g_58056_(_36294_, _27288_, _27292_);
  xor g_58057_(_36295_, _27288_, _27293_);
  or g_58058_(_36261_, _27293_, _27294_);
  xor g_58059_(_36261_, _27292_, _27295_);
  not g_58060_(_27295_, _27296_);
  or g_58061_(_36228_, _27295_, _27297_);
  xor g_58062_(_36228_, _27296_, _27298_);
  or g_58063_(_36194_, _27298_, _27299_);
  xor g_58064_(_36194_, _27298_, _27300_);
  xor g_58065_(_36195_, _27298_, _27302_);
  and g_58066_(_36161_, _27300_, _27303_);
  or g_58067_(_36160_, _27302_, _27304_);
  xor g_58068_(_36160_, _27300_, _27305_);
  or g_58069_(_36127_, _27305_, _27306_);
  not g_58070_(_27306_, _27307_);
  xor g_58071_(_36127_, _27305_, _27308_);
  and g_58072_(_36094_, _27308_, _27309_);
  not g_58073_(_27309_, _27310_);
  xor g_58074_(_36094_, _27308_, _27311_);
  xor g_58075_(_36093_, _27308_, _27313_);
  or g_58076_(_36060_, _27313_, _27314_);
  xor g_58077_(_36060_, _27311_, _27315_);
  not g_58078_(_27315_, _27316_);
  or g_58079_(_36027_, _27315_, _27317_);
  xor g_58080_(_36027_, _27316_, _27318_);
  or g_58081_(_35994_, _27318_, _27319_);
  not g_58082_(_27319_, _27320_);
  and g_58083_(_35994_, _27318_, _27321_);
  or g_58084_(_27320_, _27321_, _27322_);
  not g_58085_(_27322_, _27324_);
  or g_58086_(_35961_, _27322_, _27325_);
  or g_58087_(_35961_, _27321_, _27326_);
  xor g_58088_(_35961_, _27322_, _27327_);
  xor g_58089_(_35961_, _27324_, _27328_);
  or g_58090_(_35928_, _27328_, _27329_);
  not g_58091_(_27329_, _27330_);
  xor g_58092_(_35928_, _27327_, _27331_);
  not g_58093_(_27331_, _27332_);
  or g_58094_(_35895_, _27331_, _27333_);
  xor g_58095_(_35895_, _27332_, _27335_);
  or g_58096_(_35861_, _27335_, _27336_);
  xor g_58097_(_35861_, _27335_, _27337_);
  xor g_58098_(_35862_, _27335_, _27338_);
  or g_58099_(_35828_, _27338_, _27339_);
  xor g_58100_(_35828_, _27337_, _27340_);
  or g_58101_(_35794_, _27340_, _27341_);
  xor g_58102_(_35795_, _27340_, _27342_);
  or g_58103_(_35760_, _27342_, _27343_);
  xor g_58104_(_35761_, _27342_, _27344_);
  not g_58105_(_27344_, _27346_);
  or g_58106_(_35727_, _27344_, _27347_);
  not g_58107_(_27347_, _27348_);
  xor g_58108_(_35727_, _27344_, _27349_);
  xor g_58109_(_35727_, _27346_, _27350_);
  or g_58110_(_35694_, _27350_, _27351_);
  xor g_58111_(_35694_, _27349_, _27352_);
  or g_58112_(_35660_, _27352_, _27353_);
  xor g_58113_(_35661_, _27352_, _27354_);
  or g_58114_(_35626_, _27354_, _27355_);
  xor g_58115_(_35627_, _27354_, _27357_);
  or g_58116_(_35592_, _27357_, _27358_);
  xor g_58117_(_35592_, _27357_, _27359_);
  xor g_58118_(_35593_, _27357_, _27360_);
  or g_58119_(_35559_, _27360_, _27361_);
  xor g_58120_(_35559_, _27359_, _27362_);
  not g_58121_(_27362_, _27363_);
  or g_58122_(_35526_, _27362_, _27364_);
  xor g_58123_(_35526_, _27363_, _27365_);
  or g_58124_(_35493_, _27365_, _27366_);
  xor g_58125_(_35493_, _27365_, _27368_);
  not g_58126_(_27368_, _27369_);
  and g_58127_(_35460_, _27368_, _27370_);
  or g_58128_(_35459_, _27369_, _27371_);
  xor g_58129_(_35459_, _27368_, _27372_);
  or g_58130_(_35425_, _27372_, _27373_);
  xor g_58131_(_35426_, _27372_, _27374_);
  or g_58132_(_35391_, _27374_, _27375_);
  xor g_58133_(_35392_, _27374_, _27376_);
  not g_58134_(_27376_, _27377_);
  or g_58135_(_35358_, _27376_, _27379_);
  xor g_58136_(_35358_, _27376_, _27380_);
  xor g_58137_(_35358_, _27377_, _27381_);
  or g_58138_(_35325_, _27381_, _27382_);
  xor g_58139_(_35325_, _27380_, _27383_);
  not g_58140_(_27383_, _27384_);
  or g_58141_(_35292_, _27383_, _27385_);
  xor g_58142_(_35292_, _27384_, _27386_);
  not g_58143_(_27386_, _27387_);
  or g_58144_(_35259_, _27386_, _27388_);
  xor g_58145_(_35259_, _27386_, _27390_);
  xor g_58146_(_35259_, _27387_, _27391_);
  or g_58147_(_35226_, _27391_, _27392_);
  xor g_58148_(_35226_, _27390_, _27393_);
  or g_58149_(_35192_, _27393_, _27394_);
  xor g_58150_(_35193_, _27393_, _27395_);
  not g_58151_(_27395_, _27396_);
  or g_58152_(_35159_, _27395_, _27397_);
  xor g_58153_(_35159_, _27395_, _27398_);
  xor g_58154_(_35159_, _27396_, _27399_);
  or g_58155_(_35126_, _27399_, _27401_);
  xor g_58156_(_35126_, _27398_, _27402_);
  or g_58157_(_35093_, _27402_, _27403_);
  xor g_58158_(_35092_, _27402_, _27404_);
  or g_58159_(_35057_, _27404_, _27405_);
  xor g_58160_(_35057_, _27404_, _27406_);
  not g_58161_(_27406_, _27407_);
  or g_58162_(_35024_, _27407_, _27408_);
  xor g_58163_(_35024_, _27406_, _27409_);
  not g_58164_(_27409_, _27410_);
  or g_58165_(_34991_, _27409_, _27412_);
  xor g_58166_(_34991_, _27409_, _27413_);
  xor g_58167_(_34991_, _27410_, _27414_);
  or g_58168_(_34686_, _27414_, _27415_);
  xor g_58169_(_34686_, _27413_, _27416_);
  or g_58170_(_34313_, _27416_, _27417_);
  xor g_58171_(_34324_, _27416_, _27418_);
  not g_58172_(_27418_, _27419_);
  or g_58173_(_33950_, _27418_, _27420_);
  xor g_58174_(_33950_, _27418_, _27421_);
  xor g_58175_(_33950_, _27419_, _27423_);
  or g_58176_(_33588_, _27423_, _27424_);
  not g_58177_(_27424_, _27425_);
  xor g_58178_(_33588_, _27421_, _27426_);
  or g_58179_(_33214_, _27426_, _27427_);
  xor g_58180_(_33225_, _27426_, _27428_);
  not g_58181_(_27428_, _27429_);
  or g_58182_(_32851_, _27428_, _27430_);
  xor g_58183_(_32851_, _27428_, _27431_);
  xor g_58184_(_32851_, _27429_, _27432_);
  or g_58185_(_32488_, _27432_, _27434_);
  xor g_58186_(_32488_, _27431_, _27435_);
  not g_58187_(_27435_, _27436_);
  or g_58188_(_32126_, _27435_, _27437_);
  not g_58189_(_27437_, _27438_);
  xor g_58190_(_32126_, _27435_, _27439_);
  xor g_58191_(_32126_, _27436_, _27440_);
  or g_58192_(_31763_, _27440_, _27441_);
  xor g_58193_(_31763_, _27439_, _27442_);
  not g_58194_(_27442_, _27443_);
  or g_58195_(_31400_, _27442_, _27445_);
  xor g_58196_(_31400_, _27442_, _27446_);
  xor g_58197_(_31400_, _27443_, _27447_);
  or g_58198_(_31038_, _27447_, _27448_);
  xor g_58199_(_31038_, _27446_, _27449_);
  not g_58200_(_27449_, _27450_);
  or g_58201_(_30675_, _27449_, _27451_);
  xor g_58202_(_30675_, _27449_, _27452_);
  xor g_58203_(_30675_, _27450_, _27453_);
  or g_58204_(_30312_, _27453_, _27454_);
  xor g_58205_(_30312_, _27452_, _27456_);
  or g_58206_(_29949_, _27456_, _27457_);
  xor g_58207_(_29949_, _27456_, _27458_);
  not g_58208_(_27458_, _27459_);
  or g_58209_(_29587_, _27459_, _27460_);
  xor g_58210_(_29587_, _27458_, _27461_);
  not g_58211_(_27461_, _27462_);
  or g_58212_(_29224_, _27461_, _27463_);
  not g_58213_(_27463_, _27464_);
  xor g_58214_(_29224_, _27462_, _27465_);
  not g_58215_(_27465_, _27467_);
  or g_58216_(_28861_, _27465_, _27468_);
  xor g_58217_(_28861_, _27467_, _27469_);
  or g_58218_(_28499_, _27469_, _27470_);
  xor g_58219_(_28499_, _27469_, _27471_);
  not g_58220_(_27471_, _27472_);
  or g_58221_(_28136_, _27472_, _27473_);
  xor g_58222_(_28136_, _27471_, _27474_);
  or g_58223_(_27773_, _27474_, _27475_);
  xor g_58224_(_27773_, _27474_, _27476_);
  not g_58225_(_27476_, _27478_);
  or g_58226_(_27411_, _27478_, _27479_);
  xor g_58227_(_27411_, _27476_, _27480_);
  or g_58228_(_27048_, _27480_, _27481_);
  xor g_58229_(_27048_, _27480_, _27482_);
  not g_58230_(_27482_, _27483_);
  or g_58231_(_26685_, _27483_, _27484_);
  xor g_58232_(_26685_, _27482_, _27485_);
  not g_58233_(_27485_, _27486_);
  and g_58234_(_26322_, _27486_, _27487_);
  or g_58235_(_26311_, _27485_, _27489_);
  xor g_58236_(_26311_, _27485_, _27490_);
  not g_58237_(_27490_, _27491_);
  or g_58238_(_25948_, _27491_, _27492_);
  xor g_58239_(_25948_, _27490_, _27493_);
  not g_58240_(_27493_, _27494_);
  or g_58241_(_25585_, _27493_, _27495_);
  xor g_58242_(_25585_, _27494_, _27496_);
  not g_58243_(_27496_, _27497_);
  or g_58244_(_25222_, _27496_, _27498_);
  xor g_58245_(_25222_, _27496_, _27500_);
  xor g_58246_(_25222_, _27497_, _27501_);
  or g_58247_(_24859_, _27501_, _27502_);
  xor g_58248_(_24859_, _27500_, _27503_);
  not g_58249_(_27503_, _27504_);
  or g_58250_(_24496_, _27503_, _27505_);
  xor g_58251_(_24496_, _27504_, _27506_);
  not g_58252_(_27506_, _27507_);
  or g_58253_(_24133_, _27506_, _27508_);
  xor g_58254_(_24133_, _27506_, _27509_);
  xor g_58255_(_24133_, _27507_, _27511_);
  or g_58256_(_23770_, _27511_, _27512_);
  xor g_58257_(_23770_, _27509_, _27513_);
  not g_58258_(_27513_, _27514_);
  or g_58259_(_23407_, _27513_, _27515_);
  xor g_58260_(_23407_, _27514_, _27516_);
  not g_58261_(_27516_, _27517_);
  or g_58262_(_23044_, _27516_, _27518_);
  xor g_58263_(_23044_, _27517_, _27519_);
  not g_58264_(_27519_, _27520_);
  or g_58265_(_22681_, _27519_, _27522_);
  xor g_58266_(_22681_, _27520_, _27523_);
  or g_58267_(_22318_, _27523_, _27524_);
  not g_58268_(_27524_, _27525_);
  and g_58269_(_22318_, _27523_, _27526_);
  or g_58270_(_27525_, _27526_, _27527_);
  not g_58271_(_27527_, _27528_);
  or g_58272_(_21955_, _27527_, _27529_);
  xor g_58273_(_21955_, _27528_, _27530_);
  not g_58274_(_27530_, _27531_);
  or g_58275_(_42848_, _27530_, _27533_);
  xor g_58276_(_42848_, _27530_, _27534_);
  xor g_58277_(_42848_, _27531_, _27535_);
  or g_58278_(_42485_, _27535_, _27536_);
  xor g_58279_(_42485_, _27534_, _27537_);
  not g_58280_(_27537_, _27538_);
  or g_58281_(_42122_, _27537_, _27539_);
  xor g_58282_(_42122_, _27538_, _27540_);
  or g_58283_(_41759_, _27540_, _27541_);
  not g_58284_(_27541_, _27542_);
  and g_58285_(_41759_, _27540_, _27544_);
  or g_58286_(_27542_, _27544_, _27545_);
  or g_58287_(_41396_, _27545_, _27546_);
  xor g_58288_(_41396_, _27545_, _27547_);
  not g_58289_(_27547_, _27548_);
  or g_58290_(_41033_, _27548_, _27549_);
  not g_58291_(_27549_, _27550_);
  xor g_58292_(_41033_, _27547_, _27551_);
  not g_58293_(_27551_, _27552_);
  or g_58294_(_40670_, _27551_, _27553_);
  xor g_58295_(_40670_, _27552_, _27555_);
  or g_58296_(_40307_, _27555_, _27556_);
  xor g_58297_(_40307_, _27555_, out[640]);
  and g_58298_(_27536_, _27539_, _27557_);
  and g_58299_(_27518_, _27522_, _27558_);
  and g_58300_(_27512_, _27515_, _27559_);
  and g_58301_(_27505_, _27508_, _27560_);
  not g_58302_(_27560_, _27561_);
  and g_58303_(_27492_, _27495_, _27562_);
  not g_58304_(_27562_, _27563_);
  and g_58305_(_27412_, _27415_, _27565_);
  and g_58306_(_27364_, _27366_, _27566_);
  and g_58307_(_27353_, _27355_, _27567_);
  not g_58308_(_27567_, _27568_);
  and g_58309_(_27329_, _27333_, _27569_);
  and g_58310_(_27276_, _27280_, _27570_);
  and g_58311_(_27183_, _27186_, _27571_);
  and g_58312_(_27153_, _27156_, _27572_);
  and g_58313_(_27122_, _27126_, _27573_);
  and g_58314_(_27116_, _27119_, _27574_);
  not g_58315_(_27574_, _27576_);
  and g_58316_(_26897_, _26900_, _27577_);
  and g_58317_(_26791_, _26794_, _27578_);
  not g_58318_(_27578_, _27579_);
  and g_58319_(_26731_, _26733_, _27580_);
  and g_58320_(_26712_, _26715_, _27581_);
  not g_58321_(_27581_, _27582_);
  and g_58322_(_26687_, _26690_, _27583_);
  and g_58323_(_26669_, _26671_, _27584_);
  not g_58324_(_27584_, _27585_);
  and g_58325_(_26643_, _26646_, _27587_);
  not g_58326_(_27587_, _27588_);
  and g_58327_(_26596_, _26600_, _27589_);
  and g_58328_(_26547_, _26550_, _27590_);
  not g_58329_(_27590_, _27591_);
  and g_58330_(_26541_, _26545_, _27592_);
  and g_58331_(_26425_, _26427_, _27593_);
  and g_58332_(_26380_, _26383_, _27594_);
  not g_58333_(_27594_, _27595_);
  and g_58334_(_26373_, _26376_, _27596_);
  and g_58335_(_26368_, _26371_, _27598_);
  and g_58336_(_26356_, _26358_, _27599_);
  and g_58337_(_26349_, _26352_, _27600_);
  and g_58338_(_26345_, _26347_, _27601_);
  and g_58339_(_26337_, _26341_, _27602_);
  and g_58340_(_26331_, _26335_, _27603_);
  not g_58341_(_27603_, _27604_);
  and g_58342_(_26239_, _26314_, _27605_);
  or g_58343_(_26315_, _27605_, _27606_);
  not g_58344_(_27606_, _27607_);
  or g_58345_(_26319_, _27606_, _27609_);
  not g_58346_(_27609_, _27610_);
  or g_58347_(_26321_, _27606_, _27611_);
  xor g_58348_(_26321_, _27607_, _27612_);
  and g_58349_(_26319_, _27612_, _27613_);
  or g_58350_(_27610_, _27613_, _27614_);
  not g_58351_(_27614_, _27615_);
  and g_58352_(_26325_, _26328_, _27616_);
  xor g_58353_(_27615_, _27616_, _27617_);
  xor g_58354_(_27604_, _27617_, _27618_);
  xor g_58355_(_27603_, _27617_, _27620_);
  xor g_58356_(_27602_, _27620_, _27621_);
  not g_58357_(_27621_, _27622_);
  xor g_58358_(_27601_, _27622_, _27623_);
  xor g_58359_(_27600_, _27623_, _27624_);
  not g_58360_(_27624_, _27625_);
  xor g_58361_(_27599_, _27624_, _27626_);
  not g_58362_(_27626_, _27627_);
  or g_58363_(_26364_, _27626_, _27628_);
  not g_58364_(_27628_, _27629_);
  and g_58365_(_26361_, _26364_, _27631_);
  or g_58366_(_26361_, _27626_, _27632_);
  not g_58367_(_27632_, _27633_);
  xor g_58368_(_27627_, _27631_, _27634_);
  not g_58369_(_27634_, _27635_);
  xor g_58370_(_27598_, _27635_, _27636_);
  not g_58371_(_27636_, _27637_);
  xor g_58372_(_27598_, _27635_, _27638_);
  xor g_58373_(_27596_, _27637_, _27639_);
  or g_58374_(_27594_, _27639_, _27640_);
  xor g_58375_(_27594_, _27639_, _27642_);
  xor g_58376_(_27595_, _27639_, _27643_);
  and g_58377_(_26386_, _26389_, _27644_);
  or g_58378_(_26386_, _27643_, _27645_);
  xor g_58379_(_27642_, _27644_, _27646_);
  not g_58380_(_27646_, _27647_);
  or g_58381_(_26392_, _27646_, _27648_);
  xor g_58382_(_26392_, _27646_, _27649_);
  xor g_58383_(_26392_, _27647_, _27650_);
  or g_58384_(_26395_, _27650_, _27651_);
  not g_58385_(_27651_, _27653_);
  xor g_58386_(_26395_, _27649_, _27654_);
  or g_58387_(_26397_, _27654_, _27655_);
  xor g_58388_(_26398_, _27654_, _27656_);
  or g_58389_(_26402_, _27656_, _27657_);
  xor g_58390_(_26403_, _27656_, _27658_);
  not g_58391_(_27658_, _27659_);
  or g_58392_(_26406_, _27658_, _27660_);
  xor g_58393_(_26406_, _27658_, _27661_);
  xor g_58394_(_26406_, _27659_, _27662_);
  or g_58395_(_26408_, _27662_, _27664_);
  xor g_58396_(_26408_, _27661_, _27665_);
  not g_58397_(_27665_, _27666_);
  and g_58398_(_26411_, _26414_, _27667_);
  or g_58399_(_26411_, _27665_, _27668_);
  or g_58400_(_26414_, _27665_, _27669_);
  xor g_58401_(_27666_, _27667_, _27670_);
  not g_58402_(_27670_, _27671_);
  and g_58403_(_26417_, _26422_, _27672_);
  or g_58404_(_26422_, _27670_, _27673_);
  and g_58405_(_26418_, _27671_, _27675_);
  not g_58406_(_27675_, _27676_);
  xor g_58407_(_27671_, _27672_, _27677_);
  not g_58408_(_27677_, _27678_);
  or g_58409_(_26427_, _27677_, _27679_);
  or g_58410_(_26425_, _27677_, _27680_);
  not g_58411_(_27680_, _27681_);
  xor g_58412_(_27593_, _27678_, _27682_);
  or g_58413_(_26429_, _27682_, _27683_);
  xor g_58414_(_26429_, _27682_, _27684_);
  not g_58415_(_27684_, _27686_);
  or g_58416_(_26436_, _27686_, _27687_);
  xor g_58417_(_26436_, _27684_, _27688_);
  and g_58418_(_26433_, _27688_, _27689_);
  or g_58419_(_26433_, _27682_, _27690_);
  not g_58420_(_27690_, _27691_);
  or g_58421_(_27689_, _27691_, _27692_);
  or g_58422_(_26439_, _27692_, _27693_);
  xor g_58423_(_26439_, _27692_, _27694_);
  not g_58424_(_27694_, _27695_);
  and g_58425_(_26441_, _26445_, _27697_);
  xor g_58426_(_27694_, _27697_, _27698_);
  xor g_58427_(_27694_, _27697_, _27699_);
  or g_58428_(_26448_, _27698_, _27700_);
  xor g_58429_(_26448_, _27699_, _27701_);
  xor g_58430_(_26449_, _27699_, _27702_);
  or g_58431_(_26452_, _27702_, _27703_);
  xor g_58432_(_26452_, _27701_, _27704_);
  not g_58433_(_27704_, _27705_);
  or g_58434_(_26456_, _27704_, _27706_);
  xor g_58435_(_26456_, _27704_, _27708_);
  xor g_58436_(_26456_, _27705_, _27709_);
  or g_58437_(_26459_, _27709_, _27710_);
  xor g_58438_(_26459_, _27708_, _27711_);
  not g_58439_(_27711_, _27712_);
  or g_58440_(_26462_, _27711_, _27713_);
  xor g_58441_(_26462_, _27711_, _27714_);
  xor g_58442_(_26462_, _27712_, _27715_);
  or g_58443_(_26466_, _27715_, _27716_);
  xor g_58444_(_26466_, _27714_, _27717_);
  not g_58445_(_27717_, _27719_);
  or g_58446_(_26468_, _27717_, _27720_);
  xor g_58447_(_26468_, _27717_, _27721_);
  xor g_58448_(_26468_, _27719_, _27722_);
  and g_58449_(_26471_, _27722_, _27723_);
  or g_58450_(_26472_, _27721_, _27724_);
  or g_58451_(_26471_, _27717_, _27725_);
  not g_58452_(_27725_, _27726_);
  and g_58453_(_27724_, _27725_, _27727_);
  or g_58454_(_27723_, _27726_, _27728_);
  and g_58455_(_26475_, _27728_, _27730_);
  or g_58456_(_26477_, _27727_, _27731_);
  or g_58457_(_26475_, _27723_, _27732_);
  not g_58458_(_27732_, _27733_);
  and g_58459_(_27731_, _27732_, _27734_);
  or g_58460_(_27730_, _27733_, _27735_);
  or g_58461_(_26482_, _27735_, _27736_);
  not g_58462_(_27736_, _27737_);
  or g_58463_(_26479_, _27735_, _27738_);
  xor g_58464_(_26479_, _27734_, _27739_);
  or g_58465_(_26484_, _27739_, _27741_);
  xor g_58466_(_26485_, _27739_, _27742_);
  and g_58467_(_26482_, _27742_, _27743_);
  or g_58468_(_27737_, _27743_, _27744_);
  and g_58469_(_26490_, _26492_, _27745_);
  not g_58470_(_27745_, _27746_);
  or g_58471_(_26490_, _27744_, _27747_);
  or g_58472_(_26492_, _27744_, _27748_);
  xor g_58473_(_27744_, _27746_, _27749_);
  or g_58474_(_26494_, _27749_, _27750_);
  xor g_58475_(_26495_, _27749_, _27752_);
  or g_58476_(_26497_, _27752_, _27753_);
  xor g_58477_(_26499_, _27752_, _27754_);
  and g_58478_(_26503_, _27754_, _27755_);
  or g_58479_(_26503_, _27752_, _27756_);
  not g_58480_(_27756_, _27757_);
  or g_58481_(_27755_, _27757_, _27758_);
  and g_58482_(_26505_, _27758_, _27759_);
  or g_58483_(_26505_, _27754_, _27760_);
  not g_58484_(_27760_, _27761_);
  or g_58485_(_27759_, _27761_, _27763_);
  and g_58486_(_26508_, _26512_, _27764_);
  not g_58487_(_27764_, _27765_);
  or g_58488_(_27763_, _27764_, _27766_);
  xor g_58489_(_27763_, _27765_, _27767_);
  not g_58490_(_27767_, _27768_);
  or g_58491_(_26515_, _27767_, _27769_);
  xor g_58492_(_26515_, _27767_, _27770_);
  xor g_58493_(_26515_, _27768_, _27771_);
  or g_58494_(_26518_, _27771_, _27772_);
  xor g_58495_(_26518_, _27770_, _27774_);
  not g_58496_(_27774_, _27775_);
  or g_58497_(_26521_, _27774_, _27776_);
  not g_58498_(_27776_, _27777_);
  or g_58499_(_26525_, _27774_, _27778_);
  xor g_58500_(_26525_, _27774_, _27779_);
  xor g_58501_(_26525_, _27775_, _27780_);
  and g_58502_(_26521_, _27780_, _27781_);
  or g_58503_(_26522_, _27779_, _27782_);
  and g_58504_(_27776_, _27782_, _27783_);
  or g_58505_(_27777_, _27781_, _27785_);
  or g_58506_(_26528_, _27785_, _27786_);
  xor g_58507_(_26528_, _27783_, _27787_);
  not g_58508_(_27787_, _27788_);
  or g_58509_(_26534_, _27787_, _27789_);
  xor g_58510_(_26534_, _27788_, _27790_);
  and g_58511_(_26530_, _27790_, _27791_);
  or g_58512_(_26530_, _27785_, _27792_);
  not g_58513_(_27792_, _27793_);
  or g_58514_(_27791_, _27793_, _27794_);
  or g_58515_(_26537_, _27794_, _27796_);
  xor g_58516_(_26538_, _27794_, _27797_);
  and g_58517_(_26530_, _26534_, _27798_);
  xor g_58518_(_27787_, _27798_, _27799_);
  and g_58519_(_26538_, _27799_, _27800_);
  xor g_58520_(_26537_, _27799_, _27801_);
  xor g_58521_(_27592_, _27801_, _27802_);
  not g_58522_(_27802_, _27803_);
  xor g_58523_(_27590_, _27802_, _27804_);
  xor g_58524_(_27591_, _27802_, _27805_);
  and g_58525_(_26554_, _26556_, _27807_);
  or g_58526_(_26554_, _27804_, _27808_);
  not g_58527_(_27808_, _27809_);
  or g_58528_(_26556_, _27804_, _27810_);
  not g_58529_(_27810_, _27811_);
  or g_58530_(_27809_, _27811_, _27812_);
  xor g_58531_(_27805_, _27807_, _27813_);
  or g_58532_(_26558_, _27813_, _27814_);
  xor g_58533_(_26559_, _27813_, _27815_);
  not g_58534_(_27815_, _27816_);
  or g_58535_(_26562_, _27815_, _27818_);
  xor g_58536_(_26562_, _27815_, _27819_);
  xor g_58537_(_26562_, _27816_, _27820_);
  or g_58538_(_26565_, _27820_, _27821_);
  xor g_58539_(_26565_, _27819_, _27822_);
  or g_58540_(_26568_, _27822_, _27823_);
  xor g_58541_(_26568_, _27822_, _27824_);
  xor g_58542_(_26569_, _27822_, _27825_);
  or g_58543_(_26571_, _27825_, _27826_);
  xor g_58544_(_26571_, _27824_, _27827_);
  or g_58545_(_26573_, _27827_, _27829_);
  xor g_58546_(_26574_, _27827_, _27830_);
  or g_58547_(_26578_, _27830_, _27831_);
  xor g_58548_(_26578_, _27830_, _27832_);
  xor g_58549_(_26579_, _27830_, _27833_);
  or g_58550_(_26582_, _27833_, _27834_);
  xor g_58551_(_26582_, _27832_, _27835_);
  or g_58552_(_26588_, _27835_, _27836_);
  not g_58553_(_27836_, _27837_);
  and g_58554_(_26584_, _27835_, _27838_);
  or g_58555_(_26584_, _27833_, _27840_);
  not g_58556_(_27840_, _27841_);
  or g_58557_(_27838_, _27841_, _27842_);
  and g_58558_(_26588_, _27842_, _27843_);
  or g_58559_(_27837_, _27843_, _27844_);
  not g_58560_(_27844_, _27845_);
  and g_58561_(_26591_, _26594_, _27846_);
  or g_58562_(_26591_, _27844_, _27847_);
  xor g_58563_(_27844_, _27846_, _27848_);
  xor g_58564_(_27845_, _27846_, _27849_);
  xor g_58565_(_27589_, _27848_, _27851_);
  or g_58566_(_26603_, _27851_, _27852_);
  xor g_58567_(_26603_, _27851_, _27853_);
  not g_58568_(_27853_, _27854_);
  and g_58569_(_26609_, _27853_, _27855_);
  or g_58570_(_26610_, _27854_, _27856_);
  or g_58571_(_26605_, _27851_, _27857_);
  xor g_58572_(_26605_, _27853_, _27858_);
  and g_58573_(_26610_, _27858_, _27859_);
  or g_58574_(_27855_, _27859_, _27860_);
  and g_58575_(_26612_, _27860_, _27862_);
  or g_58576_(_26612_, _27858_, _27863_);
  not g_58577_(_27863_, _27864_);
  or g_58578_(_27862_, _27864_, _27865_);
  or g_58579_(_26618_, _27865_, _27866_);
  not g_58580_(_27866_, _27867_);
  and g_58581_(_26615_, _27865_, _27868_);
  or g_58582_(_26615_, _27860_, _27869_);
  not g_58583_(_27869_, _27870_);
  or g_58584_(_27868_, _27870_, _27871_);
  and g_58585_(_26618_, _27871_, _27873_);
  or g_58586_(_27867_, _27873_, _27874_);
  and g_58587_(_26622_, _27874_, _27875_);
  or g_58588_(_26622_, _27871_, _27876_);
  not g_58589_(_27876_, _27877_);
  or g_58590_(_27875_, _27877_, _27878_);
  or g_58591_(_26628_, _27878_, _27879_);
  not g_58592_(_27879_, _27880_);
  or g_58593_(_26625_, _27878_, _27881_);
  xor g_58594_(_26626_, _27878_, _27882_);
  and g_58595_(_26628_, _27882_, _27884_);
  or g_58596_(_27880_, _27884_, _27885_);
  and g_58597_(_26632_, _27885_, _27886_);
  or g_58598_(_26632_, _27882_, _27887_);
  not g_58599_(_27887_, _27888_);
  or g_58600_(_27886_, _27888_, _27889_);
  or g_58601_(_26639_, _27889_, _27890_);
  not g_58602_(_27890_, _27891_);
  xor g_58603_(_26636_, _27889_, _27892_);
  and g_58604_(_26639_, _27892_, _27893_);
  or g_58605_(_27891_, _27893_, _27895_);
  or g_58606_(_26635_, _27885_, _27896_);
  not g_58607_(_27896_, _27897_);
  xor g_58608_(_27587_, _27895_, _27898_);
  xor g_58609_(_27588_, _27895_, _27899_);
  or g_58610_(_26649_, _27899_, _27900_);
  xor g_58611_(_26649_, _27898_, _27901_);
  and g_58612_(_26651_, _27901_, _27902_);
  or g_58613_(_26651_, _27899_, _27903_);
  not g_58614_(_27903_, _27904_);
  or g_58615_(_27902_, _27904_, _27906_);
  or g_58616_(_26657_, _27906_, _27907_);
  not g_58617_(_27907_, _27908_);
  and g_58618_(_26655_, _27906_, _27909_);
  or g_58619_(_26655_, _27902_, _27910_);
  not g_58620_(_27910_, _27911_);
  or g_58621_(_27909_, _27911_, _27912_);
  and g_58622_(_26657_, _27912_, _27913_);
  or g_58623_(_27908_, _27913_, _27914_);
  and g_58624_(_26660_, _27914_, _27915_);
  or g_58625_(_26660_, _27912_, _27917_);
  not g_58626_(_27917_, _27918_);
  or g_58627_(_27915_, _27918_, _27919_);
  and g_58628_(_26662_, _26666_, _27920_);
  not g_58629_(_27920_, _27921_);
  xor g_58630_(_27919_, _27921_, _27922_);
  xor g_58631_(_27585_, _27922_, _27923_);
  or g_58632_(_26673_, _27923_, _27924_);
  xor g_58633_(_26673_, _27923_, _27925_);
  not g_58634_(_27925_, _27926_);
  and g_58635_(_26681_, _27925_, _27928_);
  or g_58636_(_26678_, _27926_, _27929_);
  xor g_58637_(_26677_, _27925_, _27930_);
  not g_58638_(_27930_, _27931_);
  or g_58639_(_26683_, _27931_, _27932_);
  xor g_58640_(_26683_, _27930_, _27933_);
  and g_58641_(_26680_, _27933_, _27934_);
  or g_58642_(_27928_, _27934_, _27935_);
  not g_58643_(_27935_, _27936_);
  xor g_58644_(_27583_, _27936_, _27937_);
  not g_58645_(_27937_, _27939_);
  and g_58646_(_26692_, _26695_, _27940_);
  or g_58647_(_27937_, _27940_, _27941_);
  not g_58648_(_27941_, _27942_);
  xor g_58649_(_27937_, _27940_, _27943_);
  xor g_58650_(_27939_, _27940_, _27944_);
  and g_58651_(_26700_, _27943_, _27945_);
  or g_58652_(_26699_, _27944_, _27946_);
  xor g_58653_(_26700_, _27943_, _27947_);
  xor g_58654_(_26699_, _27943_, _27948_);
  and g_58655_(_26703_, _27947_, _27950_);
  or g_58656_(_26702_, _27948_, _27951_);
  xor g_58657_(_26702_, _27947_, _27952_);
  not g_58658_(_27952_, _27953_);
  and g_58659_(_26705_, _26709_, _27954_);
  xor g_58660_(_27953_, _27954_, _27955_);
  xor g_58661_(_27582_, _27955_, _27956_);
  not g_58662_(_27956_, _27957_);
  or g_58663_(_26719_, _27956_, _27958_);
  or g_58664_(_26721_, _27956_, _27959_);
  and g_58665_(_26719_, _26721_, _27961_);
  or g_58666_(_27956_, _27961_, _27962_);
  xor g_58667_(_27956_, _27961_, _27963_);
  xor g_58668_(_27957_, _27961_, _27964_);
  or g_58669_(_26723_, _27964_, _27965_);
  xor g_58670_(_26723_, _27963_, _27966_);
  and g_58671_(_26726_, _26728_, _27967_);
  xor g_58672_(_27966_, _27967_, _27968_);
  not g_58673_(_27968_, _27969_);
  xor g_58674_(_27580_, _27968_, _27970_);
  or g_58675_(_26736_, _27970_, _27972_);
  xor g_58676_(_26737_, _27970_, _27973_);
  or g_58677_(_26739_, _27973_, _27974_);
  xor g_58678_(_26741_, _27973_, _27975_);
  and g_58679_(_26744_, _26747_, _27976_);
  xor g_58680_(_27975_, _27976_, _27977_);
  not g_58681_(_27977_, _27978_);
  and g_58682_(_26756_, _27977_, _27979_);
  or g_58683_(_26755_, _27978_, _27980_);
  and g_58684_(_26749_, _26755_, _27981_);
  and g_58685_(_26750_, _27977_, _27983_);
  or g_58686_(_26749_, _27978_, _27984_);
  xor g_58687_(_27977_, _27981_, _27985_);
  or g_58688_(_26758_, _27985_, _27986_);
  xor g_58689_(_26759_, _27985_, _27987_);
  or g_58690_(_26761_, _27987_, _27988_);
  or g_58691_(_26765_, _27987_, _27989_);
  and g_58692_(_26761_, _26765_, _27990_);
  not g_58693_(_27990_, _27991_);
  xor g_58694_(_27987_, _27990_, _27992_);
  xor g_58695_(_27987_, _27991_, _27994_);
  or g_58696_(_26768_, _27994_, _27995_);
  xor g_58697_(_26768_, _27992_, _27996_);
  and g_58698_(_26770_, _27996_, _27997_);
  or g_58699_(_26770_, _27994_, _27998_);
  not g_58700_(_27998_, _27999_);
  or g_58701_(_27997_, _27999_, _28000_);
  and g_58702_(_26774_, _28000_, _28001_);
  or g_58703_(_26774_, _27997_, _28002_);
  not g_58704_(_28002_, _28003_);
  or g_58705_(_28001_, _28003_, _28005_);
  and g_58706_(_26776_, _26779_, _28006_);
  xor g_58707_(_28005_, _28006_, _28007_);
  not g_58708_(_28007_, _28008_);
  and g_58709_(_26782_, _26786_, _28009_);
  xor g_58710_(_28007_, _28009_, _28010_);
  and g_58711_(_26787_, _28007_, _28011_);
  or g_58712_(_26786_, _28008_, _28012_);
  and g_58713_(_26783_, _28007_, _28013_);
  not g_58714_(_28013_, _28014_);
  xor g_58715_(_27578_, _28010_, _28016_);
  xor g_58716_(_27579_, _28010_, _28017_);
  or g_58717_(_26798_, _28017_, _28018_);
  xor g_58718_(_26798_, _28016_, _28019_);
  and g_58719_(_26801_, _28019_, _28020_);
  or g_58720_(_26801_, _28017_, _28021_);
  not g_58721_(_28021_, _28022_);
  or g_58722_(_28020_, _28022_, _28023_);
  or g_58723_(_26807_, _28023_, _28024_);
  not g_58724_(_28024_, _28025_);
  and g_58725_(_26804_, _28023_, _28027_);
  or g_58726_(_26804_, _28020_, _28028_);
  not g_58727_(_28028_, _28029_);
  or g_58728_(_28027_, _28029_, _28030_);
  and g_58729_(_26807_, _28030_, _28031_);
  or g_58730_(_28025_, _28031_, _28032_);
  not g_58731_(_28032_, _28033_);
  or g_58732_(_26810_, _28030_, _28034_);
  xor g_58733_(_26810_, _28032_, _28035_);
  xor g_58734_(_26810_, _28033_, _28036_);
  or g_58735_(_26815_, _28036_, _28038_);
  not g_58736_(_28038_, _28039_);
  or g_58737_(_26813_, _28036_, _28040_);
  xor g_58738_(_26813_, _28035_, _28041_);
  and g_58739_(_26815_, _28041_, _28042_);
  or g_58740_(_28039_, _28042_, _28043_);
  and g_58741_(_26819_, _28043_, _28044_);
  or g_58742_(_26819_, _28041_, _28045_);
  not g_58743_(_28045_, _28046_);
  or g_58744_(_28044_, _28046_, _28047_);
  not g_58745_(_28047_, _28049_);
  and g_58746_(_26821_, _26823_, _28050_);
  or g_58747_(_28047_, _28050_, _28051_);
  xor g_58748_(_28049_, _28050_, _28052_);
  or g_58749_(_26826_, _28052_, _28053_);
  not g_58750_(_28053_, _28054_);
  or g_58751_(_26830_, _28052_, _28055_);
  and g_58752_(_26826_, _26830_, _28056_);
  xor g_58753_(_28052_, _28056_, _28057_);
  not g_58754_(_28057_, _28058_);
  or g_58755_(_26833_, _28058_, _28060_);
  not g_58756_(_28060_, _28061_);
  or g_58757_(_26836_, _28058_, _28062_);
  xor g_58758_(_26836_, _28057_, _28063_);
  and g_58759_(_26833_, _28063_, _28064_);
  or g_58760_(_28061_, _28064_, _28065_);
  or g_58761_(_26838_, _28065_, _28066_);
  or g_58762_(_26841_, _28065_, _28067_);
  xor g_58763_(_26833_, _28057_, _28068_);
  xor g_58764_(_26836_, _28068_, _28069_);
  xor g_58765_(_26838_, _28069_, _28071_);
  xor g_58766_(_26842_, _28071_, _28072_);
  not g_58767_(_28072_, _28073_);
  or g_58768_(_26844_, _28072_, _28074_);
  not g_58769_(_28074_, _28075_);
  or g_58770_(_26849_, _28072_, _28076_);
  xor g_58771_(_26849_, _28072_, _28077_);
  xor g_58772_(_26849_, _28073_, _28078_);
  and g_58773_(_26844_, _28078_, _28079_);
  or g_58774_(_26845_, _28077_, _28080_);
  and g_58775_(_28074_, _28080_, _28082_);
  or g_58776_(_28075_, _28079_, _28083_);
  or g_58777_(_26852_, _28083_, _28084_);
  xor g_58778_(_26852_, _28082_, _28085_);
  and g_58779_(_26855_, _28082_, _28086_);
  or g_58780_(_26854_, _28083_, _28087_);
  xor g_58781_(_26855_, _28085_, _28088_);
  and g_58782_(_26858_, _26862_, _28089_);
  not g_58783_(_28089_, _28090_);
  xor g_58784_(_28088_, _28090_, _28091_);
  and g_58785_(_26865_, _26868_, _28093_);
  not g_58786_(_28093_, _28094_);
  xor g_58787_(_28091_, _28094_, _28095_);
  or g_58788_(_26870_, _28095_, _28096_);
  xor g_58789_(_26870_, _28095_, _28097_);
  not g_58790_(_28097_, _28098_);
  and g_58791_(_26874_, _28097_, _28099_);
  not g_58792_(_28099_, _28100_);
  xor g_58793_(_26873_, _28097_, _28101_);
  not g_58794_(_28101_, _28102_);
  and g_58795_(_26878_, _26880_, _28104_);
  xor g_58796_(_28101_, _28104_, _28105_);
  xor g_58797_(_28102_, _28104_, _28106_);
  or g_58798_(_26882_, _28106_, _28107_);
  xor g_58799_(_26882_, _28105_, _28108_);
  and g_58800_(_26886_, _26889_, _28109_);
  not g_58801_(_28109_, _28110_);
  xor g_58802_(_28108_, _28110_, _28111_);
  or g_58803_(_26893_, _28111_, _28112_);
  not g_58804_(_28112_, _28113_);
  and g_58805_(_26891_, _26893_, _28115_);
  and g_58806_(_28111_, _28115_, _28116_);
  or g_58807_(_26891_, _28111_, _28117_);
  not g_58808_(_28117_, _28118_);
  or g_58809_(_28116_, _28118_, _28119_);
  or g_58810_(_28113_, _28119_, _28120_);
  xor g_58811_(_28111_, _28115_, _28121_);
  xor g_58812_(_27577_, _28121_, _28122_);
  not g_58813_(_28122_, _28123_);
  or g_58814_(_26902_, _28122_, _28124_);
  not g_58815_(_28124_, _28126_);
  xor g_58816_(_26902_, _28123_, _28127_);
  not g_58817_(_28127_, _28128_);
  and g_58818_(_26904_, _26908_, _28129_);
  xor g_58819_(_28128_, _28129_, _28130_);
  xor g_58820_(_28127_, _28129_, _28131_);
  or g_58821_(_26911_, _28130_, _28132_);
  xor g_58822_(_26911_, _28131_, _28133_);
  not g_58823_(_28133_, _28134_);
  or g_58824_(_26914_, _28133_, _28135_);
  not g_58825_(_28135_, _28137_);
  xor g_58826_(_26914_, _28134_, _28138_);
  and g_58827_(_26918_, _28138_, _28139_);
  or g_58828_(_26918_, _28133_, _28140_);
  not g_58829_(_28140_, _28141_);
  or g_58830_(_28139_, _28141_, _28142_);
  not g_58831_(_28142_, _28143_);
  and g_58832_(_26924_, _28143_, _28144_);
  not g_58833_(_28144_, _28145_);
  and g_58834_(_26920_, _28142_, _28146_);
  or g_58835_(_26920_, _28139_, _28148_);
  not g_58836_(_28148_, _28149_);
  or g_58837_(_28146_, _28149_, _28150_);
  and g_58838_(_26923_, _28150_, _28151_);
  or g_58839_(_28144_, _28151_, _28152_);
  and g_58840_(_26926_, _28152_, _28153_);
  or g_58841_(_26926_, _28150_, _28154_);
  not g_58842_(_28154_, _28155_);
  or g_58843_(_28153_, _28155_, _28156_);
  not g_58844_(_28156_, _28157_);
  and g_58845_(_26930_, _26933_, _28159_);
  or g_58846_(_28156_, _28159_, _28160_);
  xor g_58847_(_28157_, _28159_, _28161_);
  not g_58848_(_28161_, _28162_);
  and g_58849_(_26935_, _26937_, _28163_);
  or g_58850_(_26937_, _28161_, _28164_);
  not g_58851_(_28164_, _28165_);
  or g_58852_(_26935_, _28161_, _28166_);
  xor g_58853_(_28162_, _28163_, _28167_);
  or g_58854_(_26940_, _28167_, _28168_);
  xor g_58855_(_26941_, _28167_, _28170_);
  not g_58856_(_28170_, _28171_);
  and g_58857_(_26943_, _26945_, _28172_);
  xor g_58858_(_28170_, _28172_, _28173_);
  xor g_58859_(_28171_, _28172_, _28174_);
  or g_58860_(_26947_, _28174_, _28175_);
  not g_58861_(_28175_, _28176_);
  xor g_58862_(_26947_, _28173_, _28177_);
  or g_58863_(_26953_, _28177_, _28178_);
  and g_58864_(_26952_, _28177_, _28179_);
  not g_58865_(_28179_, _28181_);
  and g_58866_(_26950_, _28177_, _28182_);
  not g_58867_(_28182_, _28183_);
  or g_58868_(_26950_, _28174_, _28184_);
  and g_58869_(_28178_, _28184_, _28185_);
  not g_58870_(_28185_, _28186_);
  and g_58871_(_28183_, _28185_, _28187_);
  or g_58872_(_28182_, _28186_, _28188_);
  and g_58873_(_28181_, _28188_, _28189_);
  or g_58874_(_28179_, _28187_, _28190_);
  and g_58875_(_26956_, _26959_, _28192_);
  xor g_58876_(_28190_, _28192_, _28193_);
  not g_58877_(_28193_, _28194_);
  and g_58878_(_26962_, _26965_, _28195_);
  xor g_58879_(_28194_, _28195_, _28196_);
  xor g_58880_(_28193_, _28195_, _28197_);
  or g_58881_(_26968_, _28196_, _28198_);
  xor g_58882_(_26968_, _28197_, _28199_);
  and g_58883_(_26970_, _26973_, _28200_);
  not g_58884_(_28200_, _28201_);
  or g_58885_(_26970_, _28199_, _28203_);
  or g_58886_(_28199_, _28200_, _28204_);
  xor g_58887_(_28199_, _28201_, _28205_);
  and g_58888_(_26976_, _26979_, _28206_);
  not g_58889_(_28206_, _28207_);
  or g_58890_(_26979_, _28205_, _28208_);
  or g_58891_(_26976_, _28205_, _28209_);
  xor g_58892_(_28205_, _28206_, _28210_);
  xor g_58893_(_28205_, _28207_, _28211_);
  or g_58894_(_26981_, _28211_, _28212_);
  xor g_58895_(_26981_, _28210_, _28214_);
  or g_58896_(_26985_, _28214_, _28215_);
  xor g_58897_(_26985_, _28214_, _28216_);
  and g_58898_(_26988_, _26990_, _28217_);
  xor g_58899_(_28216_, _28217_, _28218_);
  and g_58900_(_26996_, _26998_, _28219_);
  not g_58901_(_28219_, _28220_);
  or g_58902_(_26996_, _28218_, _28221_);
  not g_58903_(_28221_, _28222_);
  or g_58904_(_26998_, _28218_, _28223_);
  xor g_58905_(_28218_, _28220_, _28225_);
  not g_58906_(_28225_, _28226_);
  or g_58907_(_27000_, _28225_, _28227_);
  xor g_58908_(_27000_, _28225_, _28228_);
  xor g_58909_(_27000_, _28226_, _28229_);
  or g_58910_(_27006_, _28229_, _28230_);
  and g_58911_(_27002_, _27006_, _28231_);
  or g_58912_(_27002_, _28225_, _28232_);
  xor g_58913_(_28228_, _28231_, _28233_);
  or g_58914_(_27008_, _28233_, _28234_);
  xor g_58915_(_27008_, _28233_, _28236_);
  not g_58916_(_28236_, _28237_);
  or g_58917_(_27010_, _28237_, _28238_);
  xor g_58918_(_27011_, _28236_, _28239_);
  xor g_58919_(_27010_, _28236_, _28240_);
  and g_58920_(_27013_, _27017_, _28241_);
  or g_58921_(_27013_, _28240_, _28242_);
  or g_58922_(_27017_, _28240_, _28243_);
  and g_58923_(_28242_, _28243_, _28244_);
  xor g_58924_(_28239_, _28241_, _28245_);
  or g_58925_(_27019_, _28245_, _28247_);
  xor g_58926_(_27019_, _28245_, _28248_);
  xor g_58927_(_27020_, _28245_, _28249_);
  or g_58928_(_27022_, _28249_, _28250_);
  not g_58929_(_28250_, _28251_);
  or g_58930_(_27025_, _28249_, _28252_);
  xor g_58931_(_27025_, _28248_, _28253_);
  and g_58932_(_27022_, _28253_, _28254_);
  or g_58933_(_28251_, _28254_, _28255_);
  not g_58934_(_28255_, _28256_);
  or g_58935_(_27029_, _28255_, _28258_);
  xor g_58936_(_27029_, _28255_, _28259_);
  xor g_58937_(_27029_, _28256_, _28260_);
  and g_58938_(_27035_, _28259_, _28261_);
  not g_58939_(_28261_, _28262_);
  or g_58940_(_27031_, _28255_, _28263_);
  not g_58941_(_28263_, _28264_);
  and g_58942_(_27031_, _28260_, _28265_);
  or g_58943_(_27032_, _28259_, _28266_);
  and g_58944_(_28263_, _28266_, _28267_);
  or g_58945_(_28264_, _28265_, _28269_);
  and g_58946_(_27034_, _28269_, _28270_);
  or g_58947_(_28261_, _28270_, _28271_);
  or g_58948_(_27043_, _28271_, _28272_);
  not g_58949_(_28272_, _28273_);
  and g_58950_(_27040_, _28271_, _28274_);
  and g_58951_(_27039_, _28267_, _28275_);
  or g_58952_(_28274_, _28275_, _28276_);
  and g_58953_(_27043_, _28276_, _28277_);
  or g_58954_(_28273_, _28277_, _28278_);
  and g_58955_(_27046_, _27049_, _28280_);
  not g_58956_(_28280_, _28281_);
  xor g_58957_(_28278_, _28281_, _28282_);
  xor g_58958_(_28278_, _28280_, _28283_);
  or g_58959_(_27052_, _28282_, _28284_);
  xor g_58960_(_27052_, _28282_, _28285_);
  xor g_58961_(_27052_, _28283_, _28286_);
  or g_58962_(_27055_, _28286_, _28287_);
  xor g_58963_(_27055_, _28285_, _28288_);
  not g_58964_(_28288_, _28289_);
  or g_58965_(_27057_, _28288_, _28291_);
  not g_58966_(_28291_, _28292_);
  or g_58967_(_27063_, _28288_, _28293_);
  xor g_58968_(_27063_, _28288_, _28294_);
  xor g_58969_(_27063_, _28289_, _28295_);
  and g_58970_(_27057_, _28295_, _28296_);
  or g_58971_(_27058_, _28294_, _28297_);
  and g_58972_(_28291_, _28297_, _28298_);
  or g_58973_(_28292_, _28296_, _28299_);
  and g_58974_(_27065_, _27067_, _28300_);
  or g_58975_(_27065_, _28299_, _28302_);
  or g_58976_(_27067_, _28299_, _28303_);
  not g_58977_(_28303_, _28304_);
  xor g_58978_(_28298_, _28300_, _28305_);
  not g_58979_(_28305_, _28306_);
  and g_58980_(_27069_, _27076_, _28307_);
  or g_58981_(_28305_, _28307_, _28308_);
  xor g_58982_(_28306_, _28307_, _28309_);
  and g_58983_(_27079_, _27082_, _28310_);
  not g_58984_(_28310_, _28311_);
  or g_58985_(_27082_, _28309_, _28313_);
  or g_58986_(_27079_, _28309_, _28314_);
  xor g_58987_(_28309_, _28311_, _28315_);
  xor g_58988_(_28309_, _28310_, _28316_);
  or g_58989_(_27084_, _28315_, _28317_);
  xor g_58990_(_27084_, _28316_, _28318_);
  and g_58991_(_27087_, _28318_, _28319_);
  or g_58992_(_27087_, _28315_, _28320_);
  not g_58993_(_28320_, _28321_);
  or g_58994_(_28319_, _28321_, _28322_);
  and g_58995_(_27090_, _28322_, _28324_);
  or g_58996_(_27090_, _28319_, _28325_);
  not g_58997_(_28325_, _28326_);
  or g_58998_(_28324_, _28326_, _28327_);
  and g_58999_(_27093_, _28327_, _28328_);
  or g_59000_(_27093_, _28322_, _28329_);
  not g_59001_(_28329_, _28330_);
  or g_59002_(_28328_, _28330_, _28331_);
  and g_59003_(_27096_, _28331_, _28332_);
  or g_59004_(_27096_, _28327_, _28333_);
  not g_59005_(_28333_, _28335_);
  or g_59006_(_28332_, _28335_, _28336_);
  or g_59007_(_27102_, _28336_, _28337_);
  not g_59008_(_28337_, _28338_);
  or g_59009_(_27098_, _28336_, _28339_);
  xor g_59010_(_27099_, _28336_, _28340_);
  and g_59011_(_27102_, _28340_, _28341_);
  or g_59012_(_28338_, _28341_, _28342_);
  and g_59013_(_27106_, _28342_, _28343_);
  or g_59014_(_27106_, _28340_, _28344_);
  not g_59015_(_28344_, _28346_);
  or g_59016_(_28343_, _28346_, _28347_);
  and g_59017_(_27109_, _27112_, _28348_);
  xor g_59018_(_28347_, _28348_, _28349_);
  not g_59019_(_28349_, _28350_);
  and g_59020_(_27576_, _28349_, _28351_);
  xor g_59021_(_27574_, _28349_, _28352_);
  not g_59022_(_28352_, _28353_);
  xor g_59023_(_27573_, _28353_, _28354_);
  and g_59024_(_27129_, _27132_, _28355_);
  not g_59025_(_28355_, _28357_);
  or g_59026_(_27132_, _28354_, _28358_);
  not g_59027_(_28358_, _28359_);
  or g_59028_(_27129_, _28354_, _28360_);
  xor g_59029_(_28354_, _28357_, _28361_);
  not g_59030_(_28361_, _28362_);
  or g_59031_(_27135_, _28361_, _28363_);
  not g_59032_(_28363_, _28364_);
  xor g_59033_(_27135_, _28361_, _28365_);
  xor g_59034_(_27135_, _28362_, _28366_);
  and g_59035_(_27138_, _27141_, _28368_);
  or g_59036_(_27141_, _28366_, _28369_);
  or g_59037_(_27138_, _28361_, _28370_);
  and g_59038_(_28369_, _28370_, _28371_);
  xor g_59039_(_28365_, _28368_, _28372_);
  not g_59040_(_28372_, _28373_);
  and g_59041_(_27144_, _27148_, _28374_);
  or g_59042_(_28372_, _28374_, _28375_);
  xor g_59043_(_28372_, _28374_, _28376_);
  xor g_59044_(_28373_, _28374_, _28377_);
  or g_59045_(_27150_, _28377_, _28379_);
  not g_59046_(_28379_, _28380_);
  xor g_59047_(_27150_, _28377_, _28381_);
  xor g_59048_(_27150_, _28376_, _28382_);
  xor g_59049_(_27572_, _28382_, _28383_);
  xor g_59050_(_27572_, _28381_, _28384_);
  or g_59051_(_27160_, _28384_, _28385_);
  not g_59052_(_28385_, _28386_);
  xor g_59053_(_27160_, _28383_, _28387_);
  and g_59054_(_27162_, _28387_, _28388_);
  or g_59055_(_27162_, _28384_, _28390_);
  not g_59056_(_28390_, _28391_);
  or g_59057_(_28388_, _28391_, _28392_);
  and g_59058_(_27165_, _28392_, _28393_);
  or g_59059_(_27165_, _28387_, _28394_);
  not g_59060_(_28394_, _28395_);
  or g_59061_(_28393_, _28395_, _28396_);
  and g_59062_(_27168_, _28396_, _28397_);
  or g_59063_(_27168_, _28392_, _28398_);
  not g_59064_(_28398_, _28399_);
  or g_59065_(_28397_, _28399_, _28401_);
  or g_59066_(_27172_, _28401_, _28402_);
  xor g_59067_(_27173_, _28401_, _28403_);
  and g_59068_(_27176_, _27179_, _28404_);
  not g_59069_(_28404_, _28405_);
  xor g_59070_(_28403_, _28405_, _28406_);
  not g_59071_(_28406_, _28407_);
  xor g_59072_(_27571_, _28407_, _28408_);
  or g_59073_(_27188_, _28408_, _28409_);
  xor g_59074_(_27188_, _28408_, _28410_);
  xor g_59075_(_27189_, _28408_, _28412_);
  and g_59076_(_27196_, _28410_, _28413_);
  or g_59077_(_27195_, _28412_, _28414_);
  xor g_59078_(_27195_, _28410_, _28415_);
  and g_59079_(_27192_, _28415_, _28416_);
  or g_59080_(_27192_, _28412_, _28417_);
  not g_59081_(_28417_, _28418_);
  or g_59082_(_28416_, _28418_, _28419_);
  not g_59083_(_28419_, _28420_);
  or g_59084_(_27199_, _28419_, _28421_);
  xor g_59085_(_27199_, _28420_, _28423_);
  and g_59086_(_27201_, _27205_, _28424_);
  or g_59087_(_27205_, _28423_, _28425_);
  or g_59088_(_27201_, _28419_, _28426_);
  or g_59089_(_28423_, _28424_, _28427_);
  xor g_59090_(_28423_, _28424_, _28428_);
  not g_59091_(_28428_, _28429_);
  and g_59092_(_27209_, _28428_, _28430_);
  or g_59093_(_27208_, _28429_, _28431_);
  xor g_59094_(_27208_, _28428_, _28432_);
  not g_59095_(_28432_, _28434_);
  and g_59096_(_27211_, _27214_, _28435_);
  xor g_59097_(_28434_, _28435_, _28436_);
  or g_59098_(_27211_, _28432_, _28437_);
  or g_59099_(_27214_, _28432_, _28438_);
  or g_59100_(_27218_, _28436_, _28439_);
  xor g_59101_(_27217_, _28436_, _28440_);
  not g_59102_(_28440_, _28441_);
  and g_59103_(_27221_, _27225_, _28442_);
  xor g_59104_(_28441_, _28442_, _28443_);
  not g_59105_(_28443_, _28445_);
  or g_59106_(_27228_, _28443_, _28446_);
  xor g_59107_(_27228_, _28443_, _28447_);
  xor g_59108_(_27228_, _28445_, _28448_);
  or g_59109_(_27233_, _28448_, _28449_);
  or g_59110_(_27230_, _28448_, _28450_);
  and g_59111_(_27230_, _27233_, _28451_);
  xor g_59112_(_28447_, _28451_, _28452_);
  not g_59113_(_28452_, _28453_);
  or g_59114_(_27237_, _28452_, _28454_);
  xor g_59115_(_27237_, _28453_, _28456_);
  and g_59116_(_27239_, _28456_, _28457_);
  or g_59117_(_27239_, _28452_, _28458_);
  not g_59118_(_28458_, _28459_);
  or g_59119_(_28457_, _28459_, _28460_);
  and g_59120_(_27242_, _28460_, _28461_);
  or g_59121_(_27242_, _28456_, _28462_);
  not g_59122_(_28462_, _28463_);
  or g_59123_(_28461_, _28463_, _28464_);
  and g_59124_(_27245_, _27249_, _28465_);
  xor g_59125_(_28464_, _28465_, _28467_);
  not g_59126_(_28467_, _28468_);
  and g_59127_(_27252_, _27255_, _28469_);
  and g_59128_(_27253_, _28467_, _28470_);
  or g_59129_(_27252_, _28468_, _28471_);
  or g_59130_(_27255_, _28468_, _28472_);
  not g_59131_(_28472_, _28473_);
  xor g_59132_(_28467_, _28469_, _28474_);
  not g_59133_(_28474_, _28475_);
  and g_59134_(_27259_, _27262_, _28476_);
  xor g_59135_(_28475_, _28476_, _28478_);
  not g_59136_(_28478_, _28479_);
  or g_59137_(_27265_, _28478_, _28480_);
  not g_59138_(_28480_, _28481_);
  xor g_59139_(_27265_, _28479_, _28482_);
  or g_59140_(_27259_, _28474_, _28483_);
  or g_59141_(_27262_, _28474_, _28484_);
  and g_59142_(_27269_, _28482_, _28485_);
  or g_59143_(_27269_, _28478_, _28486_);
  not g_59144_(_28486_, _28487_);
  or g_59145_(_28485_, _28487_, _28489_);
  not g_59146_(_28489_, _28490_);
  and g_59147_(_27271_, _27274_, _28491_);
  xor g_59148_(_28490_, _28491_, _28492_);
  not g_59149_(_28492_, _28493_);
  xor g_59150_(_27570_, _28493_, _28494_);
  xor g_59151_(_27570_, _28492_, _28495_);
  or g_59152_(_27282_, _28494_, _28496_);
  xor g_59153_(_27283_, _28495_, _28497_);
  not g_59154_(_28497_, _28498_);
  and g_59155_(_27287_, _28498_, _28500_);
  or g_59156_(_27286_, _28497_, _28501_);
  or g_59157_(_27287_, _28494_, _28502_);
  not g_59158_(_28502_, _28503_);
  and g_59159_(_28501_, _28502_, _28504_);
  or g_59160_(_28500_, _28503_, _28505_);
  and g_59161_(_27289_, _27294_, _28506_);
  xor g_59162_(_28504_, _28506_, _28507_);
  not g_59163_(_28507_, _28508_);
  or g_59164_(_27297_, _28507_, _28509_);
  xor g_59165_(_27297_, _28507_, _28511_);
  xor g_59166_(_27297_, _28508_, _28512_);
  and g_59167_(_27303_, _28511_, _28513_);
  or g_59168_(_27304_, _28512_, _28514_);
  or g_59169_(_27299_, _28512_, _28515_);
  xor g_59170_(_27299_, _28511_, _28516_);
  and g_59171_(_27304_, _28516_, _28517_);
  not g_59172_(_28517_, _28518_);
  and g_59173_(_28514_, _28518_, _28519_);
  or g_59174_(_28513_, _28517_, _28520_);
  and g_59175_(_27306_, _28520_, _28522_);
  or g_59176_(_27307_, _28519_, _28523_);
  or g_59177_(_27306_, _28516_, _28524_);
  not g_59178_(_28524_, _28525_);
  and g_59179_(_28523_, _28524_, _28526_);
  or g_59180_(_28522_, _28525_, _28527_);
  and g_59181_(_27310_, _28527_, _28528_);
  or g_59182_(_27309_, _28526_, _28529_);
  and g_59183_(_27309_, _28519_, _28530_);
  not g_59184_(_28530_, _28531_);
  and g_59185_(_28529_, _28531_, _28533_);
  or g_59186_(_28528_, _28530_, _28534_);
  or g_59187_(_27314_, _28534_, _28535_);
  xor g_59188_(_27314_, _28533_, _28536_);
  not g_59189_(_28536_, _28537_);
  or g_59190_(_27317_, _28536_, _28538_);
  xor g_59191_(_27317_, _28537_, _28539_);
  not g_59192_(_28539_, _28540_);
  and g_59193_(_27319_, _27326_, _28541_);
  xor g_59194_(_28539_, _28541_, _28542_);
  xor g_59195_(_28540_, _28541_, _28544_);
  xor g_59196_(_27569_, _28542_, _28545_);
  xor g_59197_(_27569_, _28544_, _28546_);
  or g_59198_(_27336_, _28545_, _28547_);
  xor g_59199_(_27336_, _28546_, _28548_);
  not g_59200_(_28548_, _28549_);
  or g_59201_(_27339_, _28545_, _28550_);
  xor g_59202_(_27339_, _28549_, _28551_);
  not g_59203_(_28551_, _28552_);
  and g_59204_(_27341_, _27343_, _28553_);
  xor g_59205_(_28552_, _28553_, _28555_);
  xor g_59206_(_28551_, _28553_, _28556_);
  and g_59207_(_27347_, _27351_, _28557_);
  xor g_59208_(_28556_, _28557_, _28558_);
  xor g_59209_(_27567_, _28558_, _28559_);
  xor g_59210_(_27568_, _28558_, _28560_);
  or g_59211_(_27361_, _28560_, _28561_);
  and g_59212_(_27358_, _27361_, _28562_);
  or g_59213_(_27358_, _28560_, _28563_);
  xor g_59214_(_28559_, _28562_, _28564_);
  not g_59215_(_28564_, _28566_);
  xor g_59216_(_27566_, _28566_, _28567_);
  or g_59217_(_27371_, _28567_, _28568_);
  xor g_59218_(_27370_, _28567_, _28569_);
  and g_59219_(_27373_, _28569_, _28570_);
  or g_59220_(_27373_, _28567_, _28571_);
  not g_59221_(_28571_, _28572_);
  or g_59222_(_28570_, _28572_, _28573_);
  not g_59223_(_28573_, _28574_);
  and g_59224_(_27375_, _27379_, _28575_);
  xor g_59225_(_28574_, _28575_, _28577_);
  not g_59226_(_28577_, _28578_);
  or g_59227_(_27385_, _28577_, _28579_);
  and g_59228_(_27382_, _27385_, _28580_);
  or g_59229_(_27382_, _28577_, _28581_);
  xor g_59230_(_28577_, _28580_, _28582_);
  xor g_59231_(_28578_, _28580_, _28583_);
  or g_59232_(_27388_, _28583_, _28584_);
  xor g_59233_(_27388_, _28582_, _28585_);
  not g_59234_(_28585_, _28586_);
  or g_59235_(_27392_, _28585_, _28588_);
  or g_59236_(_27394_, _28585_, _28589_);
  not g_59237_(_28589_, _28590_);
  and g_59238_(_27392_, _27394_, _28591_);
  xor g_59239_(_28586_, _28591_, _28592_);
  not g_59240_(_28592_, _28593_);
  or g_59241_(_27397_, _28592_, _28594_);
  not g_59242_(_28594_, _28595_);
  xor g_59243_(_27397_, _28593_, _28596_);
  not g_59244_(_28596_, _28597_);
  and g_59245_(_27401_, _27403_, _28599_);
  or g_59246_(_27401_, _28596_, _28600_);
  or g_59247_(_27403_, _28596_, _28601_);
  xor g_59248_(_28597_, _28599_, _28602_);
  not g_59249_(_28602_, _28603_);
  and g_59250_(_27405_, _27408_, _28604_);
  xor g_59251_(_28603_, _28604_, _28605_);
  not g_59252_(_28605_, _28606_);
  xor g_59253_(_27565_, _28606_, _28607_);
  not g_59254_(_28607_, _28608_);
  or g_59255_(_27417_, _28607_, _28610_);
  xor g_59256_(_27417_, _28607_, _28611_);
  xor g_59257_(_27417_, _28608_, _28612_);
  and g_59258_(_27420_, _27424_, _28613_);
  xor g_59259_(_28612_, _28613_, _28614_);
  xor g_59260_(_28611_, _28613_, _28615_);
  and g_59261_(_27427_, _27430_, _28616_);
  or g_59262_(_27427_, _28615_, _28617_);
  not g_59263_(_28617_, _28618_);
  or g_59264_(_27430_, _28615_, _28619_);
  xor g_59265_(_28614_, _28616_, _28621_);
  not g_59266_(_28621_, _28622_);
  or g_59267_(_27434_, _28621_, _28623_);
  xor g_59268_(_27434_, _28621_, _28624_);
  xor g_59269_(_27434_, _28622_, _28625_);
  and g_59270_(_27437_, _28625_, _28626_);
  or g_59271_(_27438_, _28624_, _28627_);
  or g_59272_(_27437_, _28621_, _28628_);
  not g_59273_(_28628_, _28629_);
  and g_59274_(_28627_, _28628_, _28630_);
  or g_59275_(_28626_, _28629_, _28632_);
  and g_59276_(_27441_, _27445_, _28633_);
  xor g_59277_(_28630_, _28633_, _28634_);
  not g_59278_(_28634_, _28635_);
  and g_59279_(_27448_, _27451_, _28636_);
  xor g_59280_(_28635_, _28636_, _28637_);
  xor g_59281_(_28634_, _28636_, _28638_);
  or g_59282_(_27454_, _28637_, _28639_);
  xor g_59283_(_27454_, _28638_, _28640_);
  or g_59284_(_27448_, _28634_, _28641_);
  or g_59285_(_27451_, _28634_, _28643_);
  and g_59286_(_27457_, _28640_, _28644_);
  or g_59287_(_27457_, _28637_, _28645_);
  not g_59288_(_28645_, _28646_);
  or g_59289_(_28644_, _28646_, _28647_);
  and g_59290_(_27460_, _28647_, _28648_);
  or g_59291_(_27460_, _28640_, _28649_);
  not g_59292_(_28649_, _28650_);
  or g_59293_(_28648_, _28650_, _28651_);
  or g_59294_(_27463_, _28651_, _28652_);
  xor g_59295_(_27464_, _28651_, _28654_);
  and g_59296_(_27468_, _28654_, _28655_);
  or g_59297_(_27468_, _28651_, _28656_);
  not g_59298_(_28656_, _28657_);
  or g_59299_(_28655_, _28657_, _28658_);
  or g_59300_(_27473_, _28658_, _28659_);
  not g_59301_(_28659_, _28660_);
  and g_59302_(_27470_, _28658_, _28661_);
  or g_59303_(_27470_, _28654_, _28662_);
  not g_59304_(_28662_, _28663_);
  or g_59305_(_28661_, _28663_, _28665_);
  and g_59306_(_27473_, _28665_, _28666_);
  or g_59307_(_28660_, _28666_, _28667_);
  or g_59308_(_27479_, _28667_, _28668_);
  not g_59309_(_28668_, _28669_);
  and g_59310_(_27475_, _28667_, _28670_);
  or g_59311_(_27475_, _28665_, _28671_);
  not g_59312_(_28671_, _28672_);
  or g_59313_(_28670_, _28672_, _28673_);
  and g_59314_(_27479_, _28673_, _28674_);
  or g_59315_(_28669_, _28674_, _28676_);
  not g_59316_(_28676_, _28677_);
  or g_59317_(_27481_, _28676_, _28678_);
  xor g_59318_(_27481_, _28676_, _28679_);
  xor g_59319_(_27481_, _28677_, _28680_);
  and g_59320_(_27487_, _28679_, _28681_);
  or g_59321_(_27489_, _28680_, _28682_);
  or g_59322_(_27489_, _28679_, _28683_);
  and g_59323_(_27484_, _28680_, _28684_);
  or g_59324_(_27484_, _28676_, _28685_);
  not g_59325_(_28685_, _28687_);
  or g_59326_(_28681_, _28687_, _28688_);
  or g_59327_(_28684_, _28688_, _28689_);
  and g_59328_(_28683_, _28689_, _28690_);
  or g_59329_(_27495_, _28690_, _28691_);
  or g_59330_(_27492_, _28690_, _28692_);
  and g_59331_(_28691_, _28692_, _28693_);
  xor g_59332_(_27563_, _28690_, _28694_);
  not g_59333_(_28694_, _28695_);
  and g_59334_(_27498_, _27502_, _28696_);
  xor g_59335_(_28695_, _28696_, _28698_);
  or g_59336_(_27502_, _28694_, _28699_);
  not g_59337_(_28699_, _28700_);
  or g_59338_(_27498_, _28694_, _28701_);
  xor g_59339_(_27561_, _28698_, _28702_);
  not g_59340_(_28702_, _28703_);
  xor g_59341_(_27559_, _28703_, _28704_);
  xor g_59342_(_27558_, _28704_, _28705_);
  not g_59343_(_28705_, _28706_);
  and g_59344_(_27525_, _28705_, _28707_);
  or g_59345_(_27524_, _28706_, _28709_);
  xor g_59346_(_27524_, _28705_, _28710_);
  not g_59347_(_28710_, _28711_);
  and g_59348_(_27529_, _27533_, _28712_);
  xor g_59349_(_28711_, _28712_, _28713_);
  not g_59350_(_28713_, _28714_);
  xor g_59351_(_27557_, _28714_, _28715_);
  or g_59352_(_27541_, _28715_, _28716_);
  xor g_59353_(_27542_, _28715_, _28717_);
  and g_59354_(_27546_, _28717_, _28718_);
  not g_59355_(_28718_, _28720_);
  or g_59356_(_27546_, _28715_, _28721_);
  not g_59357_(_28721_, _28722_);
  and g_59358_(_28720_, _28721_, _28723_);
  or g_59359_(_28718_, _28722_, _28724_);
  and g_59360_(_27549_, _28724_, _28725_);
  or g_59361_(_27550_, _28723_, _28726_);
  or g_59362_(_27549_, _28718_, _28727_);
  not g_59363_(_28727_, _28728_);
  and g_59364_(_28726_, _28727_, _28729_);
  or g_59365_(_28725_, _28728_, _28731_);
  or g_59366_(_27553_, _28731_, _28732_);
  xor g_59367_(_27553_, _28729_, _28733_);
  or g_59368_(_27556_, _28733_, _28734_);
  xor g_59369_(_27556_, _28733_, out[641]);
  or g_59370_(_27539_, _28713_, _28735_);
  or g_59371_(_27536_, _28713_, _28736_);
  or g_59372_(_27533_, _28710_, _28737_);
  or g_59373_(_27518_, _28704_, _28738_);
  or g_59374_(_27515_, _28702_, _28739_);
  or g_59375_(_27512_, _28702_, _28741_);
  or g_59376_(_27508_, _28698_, _28742_);
  or g_59377_(_27505_, _28698_, _28743_);
  and g_59378_(_28693_, _28701_, _28744_);
  or g_59379_(_27445_, _28632_, _28745_);
  not g_59380_(_28745_, _28746_);
  or g_59381_(_27415_, _28605_, _28747_);
  not g_59382_(_28747_, _28748_);
  or g_59383_(_27408_, _28602_, _28749_);
  or g_59384_(_27405_, _28602_, _28750_);
  or g_59385_(_27379_, _28573_, _28752_);
  or g_59386_(_27366_, _28564_, _28753_);
  not g_59387_(_28753_, _28754_);
  or g_59388_(_27355_, _28558_, _28755_);
  or g_59389_(_27351_, _28555_, _28756_);
  not g_59390_(_28756_, _28757_);
  and g_59391_(_27348_, _28556_, _28758_);
  or g_59392_(_27347_, _28555_, _28759_);
  or g_59393_(_27341_, _28548_, _28760_);
  or g_59394_(_27333_, _28544_, _28761_);
  and g_59395_(_27330_, _28542_, _28763_);
  or g_59396_(_27329_, _28544_, _28764_);
  or g_59397_(_27325_, _28539_, _28765_);
  or g_59398_(_27294_, _28505_, _28766_);
  not g_59399_(_28766_, _28767_);
  or g_59400_(_27276_, _28492_, _28768_);
  or g_59401_(_27249_, _28464_, _28769_);
  or g_59402_(_27225_, _28440_, _28770_);
  or g_59403_(_27221_, _28436_, _28771_);
  or g_59404_(_27183_, _28406_, _28772_);
  not g_59405_(_28772_, _28774_);
  or g_59406_(_27156_, _28382_, _28775_);
  or g_59407_(_27153_, _28382_, _28776_);
  not g_59408_(_28776_, _28777_);
  or g_59409_(_27122_, _28352_, _28778_);
  or g_59410_(_27109_, _28342_, _28779_);
  and g_59411_(_28339_, _28344_, _28780_);
  not g_59412_(_28780_, _28781_);
  and g_59413_(_28313_, _28317_, _28782_);
  or g_59414_(_27049_, _28278_, _28783_);
  and g_59415_(_28244_, _28247_, _28785_);
  not g_59416_(_28785_, _28786_);
  and g_59417_(_26991_, _28216_, _28787_);
  not g_59418_(_28787_, _28788_);
  or g_59419_(_26988_, _28214_, _28789_);
  or g_59420_(_26965_, _28193_, _28790_);
  or g_59421_(_26962_, _28193_, _28791_);
  or g_59422_(_26959_, _28189_, _28792_);
  or g_59423_(_26956_, _28189_, _28793_);
  or g_59424_(_26943_, _28167_, _28794_);
  or g_59425_(_26908_, _28127_, _28796_);
  or g_59426_(_26904_, _28122_, _28797_);
  or g_59427_(_26900_, _28120_, _28798_);
  or g_59428_(_26868_, _28091_, _28799_);
  or g_59429_(_26865_, _28091_, _28800_);
  not g_59430_(_28800_, _28801_);
  or g_59431_(_26862_, _28088_, _28802_);
  not g_59432_(_28802_, _28803_);
  and g_59433_(_28045_, _28051_, _28804_);
  or g_59434_(_26794_, _28010_, _28805_);
  not g_59435_(_28805_, _28807_);
  or g_59436_(_26791_, _28010_, _28808_);
  or g_59437_(_26779_, _28005_, _28809_);
  not g_59438_(_28809_, _28810_);
  or g_59439_(_26776_, _28000_, _28811_);
  or g_59440_(_26747_, _27975_, _28812_);
  or g_59441_(_26744_, _27973_, _28813_);
  or g_59442_(_26731_, _27969_, _28814_);
  or g_59443_(_26728_, _27966_, _28815_);
  or g_59444_(_26715_, _27955_, _28816_);
  or g_59445_(_26712_, _27955_, _28818_);
  not g_59446_(_28818_, _28819_);
  or g_59447_(_26709_, _27952_, _28820_);
  or g_59448_(_26705_, _27952_, _28821_);
  not g_59449_(_28821_, _28822_);
  or g_59450_(_26690_, _27935_, _28823_);
  not g_59451_(_28823_, _28824_);
  or g_59452_(_26687_, _27935_, _28825_);
  not g_59453_(_28825_, _28826_);
  or g_59454_(_26671_, _27922_, _28827_);
  not g_59455_(_28827_, _28829_);
  or g_59456_(_26666_, _27919_, _28830_);
  or g_59457_(_26646_, _27895_, _28831_);
  and g_59458_(_27876_, _27881_, _28832_);
  or g_59459_(_26600_, _27849_, _28833_);
  or g_59460_(_26596_, _27849_, _28834_);
  or g_59461_(_26594_, _27844_, _28835_);
  and g_59462_(_28834_, _28835_, _28836_);
  and g_59463_(_27814_, _27818_, _28837_);
  or g_59464_(_26547_, _27803_, _28838_);
  not g_59465_(_28838_, _28840_);
  or g_59466_(_26545_, _27797_, _28841_);
  and g_59467_(_27769_, _27772_, _28842_);
  and g_59468_(_27716_, _27720_, _28843_);
  or g_59469_(_26371_, _27634_, _28844_);
  or g_59470_(_26368_, _27634_, _28845_);
  or g_59471_(_26358_, _27625_, _28846_);
  or g_59472_(_26356_, _27625_, _28847_);
  or g_59473_(_26347_, _27621_, _28848_);
  or g_59474_(_26345_, _27621_, _28849_);
  or g_59475_(_26341_, _27618_, _28851_);
  or g_59476_(_26335_, _27617_, _28852_);
  or g_59477_(_26331_, _27617_, _28853_);
  not g_59478_(_28853_, _28854_);
  or g_59479_(_26328_, _27613_, _28855_);
  and g_59480_(_27609_, _27611_, _28856_);
  or g_59481_(_26325_, _27614_, _28857_);
  and g_59482_(_28855_, _28857_, _28858_);
  and g_59483_(_28856_, _28858_, _28859_);
  or g_59484_(_28853_, _28859_, _28860_);
  xor g_59485_(_28853_, _28859_, _28862_);
  xor g_59486_(_28854_, _28859_, _28863_);
  or g_59487_(_28852_, _28863_, _28864_);
  xor g_59488_(_28852_, _28862_, _28865_);
  and g_59489_(_26338_, _27620_, _28866_);
  or g_59490_(_26337_, _27618_, _28867_);
  or g_59491_(_28865_, _28867_, _28868_);
  xor g_59492_(_28865_, _28866_, _28869_);
  not g_59493_(_28869_, _28870_);
  or g_59494_(_28851_, _28869_, _28871_);
  xor g_59495_(_28851_, _28870_, _28873_);
  not g_59496_(_28873_, _28874_);
  or g_59497_(_28849_, _28873_, _28875_);
  xor g_59498_(_28849_, _28874_, _28876_);
  not g_59499_(_28876_, _28877_);
  or g_59500_(_28848_, _28876_, _28878_);
  xor g_59501_(_28848_, _28877_, _28879_);
  or g_59502_(_26349_, _27623_, _28880_);
  not g_59503_(_28880_, _28881_);
  or g_59504_(_28879_, _28880_, _28882_);
  xor g_59505_(_28879_, _28881_, _28884_);
  or g_59506_(_26352_, _27623_, _28885_);
  not g_59507_(_28885_, _28886_);
  or g_59508_(_28884_, _28885_, _28887_);
  xor g_59509_(_28884_, _28886_, _28888_);
  and g_59510_(_28847_, _28888_, _28889_);
  or g_59511_(_28847_, _28888_, _28890_);
  not g_59512_(_28890_, _28891_);
  xor g_59513_(_28847_, _28888_, _28892_);
  or g_59514_(_28889_, _28891_, _28893_);
  or g_59515_(_28846_, _28893_, _28895_);
  xor g_59516_(_28846_, _28892_, _28896_);
  or g_59517_(_27632_, _28896_, _28897_);
  xor g_59518_(_27633_, _28896_, _28898_);
  or g_59519_(_27628_, _28898_, _28899_);
  xor g_59520_(_27629_, _28898_, _28900_);
  not g_59521_(_28900_, _28901_);
  or g_59522_(_28845_, _28900_, _28902_);
  xor g_59523_(_28845_, _28900_, _28903_);
  xor g_59524_(_28845_, _28901_, _28904_);
  or g_59525_(_28844_, _28904_, _28906_);
  xor g_59526_(_28844_, _28903_, _28907_);
  or g_59527_(_26373_, _27636_, _28908_);
  or g_59528_(_26373_, _27638_, _28909_);
  not g_59529_(_28909_, _28910_);
  or g_59530_(_28907_, _28908_, _28911_);
  xor g_59531_(_28907_, _28909_, _28912_);
  xor g_59532_(_28907_, _28910_, _28913_);
  or g_59533_(_26376_, _27636_, _28914_);
  or g_59534_(_28913_, _28914_, _28915_);
  xor g_59535_(_28912_, _28914_, _28917_);
  not g_59536_(_28917_, _28918_);
  and g_59537_(_27640_, _27645_, _28919_);
  xor g_59538_(_28918_, _28919_, _28920_);
  or g_59539_(_26389_, _27643_, _28921_);
  and g_59540_(_27648_, _28921_, _28922_);
  not g_59541_(_28922_, _28923_);
  xor g_59542_(_28920_, _28923_, _28924_);
  or g_59543_(_27651_, _28924_, _28925_);
  not g_59544_(_28925_, _28926_);
  xor g_59545_(_27653_, _28924_, _28928_);
  or g_59546_(_27655_, _28928_, _28929_);
  not g_59547_(_28929_, _28930_);
  xor g_59548_(_27655_, _28928_, _28931_);
  not g_59549_(_28931_, _28932_);
  and g_59550_(_27657_, _27660_, _28933_);
  xor g_59551_(_28931_, _28933_, _28934_);
  not g_59552_(_28934_, _28935_);
  and g_59553_(_27664_, _27668_, _28936_);
  xor g_59554_(_28935_, _28936_, _28937_);
  or g_59555_(_27669_, _28937_, _28939_);
  not g_59556_(_28939_, _28940_);
  xor g_59557_(_27669_, _28937_, _28941_);
  or g_59558_(_27657_, _28932_, _28942_);
  or g_59559_(_27660_, _28932_, _28943_);
  not g_59560_(_28943_, _28944_);
  and g_59561_(_27675_, _28941_, _28945_);
  not g_59562_(_28945_, _28946_);
  xor g_59563_(_27676_, _28941_, _28947_);
  not g_59564_(_28947_, _28948_);
  or g_59565_(_27673_, _28947_, _28950_);
  xor g_59566_(_27673_, _28948_, _28951_);
  or g_59567_(_27680_, _28951_, _28952_);
  xor g_59568_(_27681_, _28951_, _28953_);
  or g_59569_(_27679_, _28953_, _28954_);
  not g_59570_(_28954_, _28955_);
  xor g_59571_(_27679_, _28953_, _28956_);
  not g_59572_(_28956_, _28957_);
  or g_59573_(_27683_, _28957_, _28958_);
  not g_59574_(_28958_, _28959_);
  xor g_59575_(_27683_, _28956_, _28961_);
  or g_59576_(_27690_, _28961_, _28962_);
  xor g_59577_(_27691_, _28961_, _28963_);
  not g_59578_(_28963_, _28964_);
  or g_59579_(_27687_, _28963_, _28965_);
  xor g_59580_(_27687_, _28964_, _28966_);
  not g_59581_(_28966_, _28967_);
  or g_59582_(_27693_, _28966_, _28968_);
  xor g_59583_(_27693_, _28966_, _28969_);
  xor g_59584_(_27693_, _28967_, _28970_);
  or g_59585_(_26441_, _27692_, _28972_);
  not g_59586_(_28972_, _28973_);
  and g_59587_(_28969_, _28973_, _28974_);
  or g_59588_(_28970_, _28972_, _28975_);
  xor g_59589_(_28969_, _28972_, _28976_);
  not g_59590_(_28976_, _28977_);
  or g_59591_(_26445_, _27695_, _28978_);
  and g_59592_(_27700_, _28978_, _28979_);
  xor g_59593_(_28976_, _28979_, _28980_);
  xor g_59594_(_28977_, _28979_, _28981_);
  and g_59595_(_27703_, _27706_, _28983_);
  not g_59596_(_28983_, _28984_);
  or g_59597_(_27703_, _28981_, _28985_);
  and g_59598_(_28980_, _28984_, _28986_);
  xor g_59599_(_28980_, _28983_, _28987_);
  or g_59600_(_27713_, _28987_, _28988_);
  or g_59601_(_27710_, _28987_, _28989_);
  and g_59602_(_28988_, _28989_, _28990_);
  not g_59603_(_28990_, _28991_);
  and g_59604_(_27710_, _28987_, _28992_);
  and g_59605_(_27713_, _28992_, _28994_);
  or g_59606_(_28991_, _28994_, _28995_);
  not g_59607_(_28995_, _28996_);
  or g_59608_(_28843_, _28995_, _28997_);
  xor g_59609_(_28843_, _28996_, _28998_);
  or g_59610_(_27725_, _28998_, _28999_);
  and g_59611_(_27725_, _28998_, _29000_);
  xor g_59612_(_27726_, _28998_, _29001_);
  and g_59613_(_27732_, _27738_, _29002_);
  xor g_59614_(_29001_, _29002_, _29003_);
  and g_59615_(_27737_, _29003_, _29005_);
  xor g_59616_(_27737_, _29003_, _29006_);
  not g_59617_(_29006_, _29007_);
  or g_59618_(_27741_, _29007_, _29008_);
  xor g_59619_(_27741_, _29006_, _29009_);
  not g_59620_(_29009_, _29010_);
  or g_59621_(_27747_, _29009_, _29011_);
  xor g_59622_(_27747_, _29010_, _29012_);
  not g_59623_(_29012_, _29013_);
  and g_59624_(_27748_, _27750_, _29014_);
  xor g_59625_(_29013_, _29014_, _29016_);
  or g_59626_(_27753_, _29016_, _29017_);
  xor g_59627_(_27753_, _29016_, _29018_);
  not g_59628_(_29018_, _29019_);
  and g_59629_(_27757_, _29018_, _29020_);
  or g_59630_(_27756_, _29019_, _29021_);
  xor g_59631_(_27756_, _29018_, _29022_);
  or g_59632_(_27760_, _29022_, _29023_);
  xor g_59633_(_27761_, _29022_, _29024_);
  xor g_59634_(_27766_, _29024_, _29025_);
  not g_59635_(_29025_, _29027_);
  xor g_59636_(_28842_, _29025_, _29028_);
  or g_59637_(_27776_, _29028_, _29029_);
  xor g_59638_(_27777_, _29028_, _29030_);
  not g_59639_(_29030_, _29031_);
  or g_59640_(_27778_, _29030_, _29032_);
  xor g_59641_(_27778_, _29031_, _29033_);
  not g_59642_(_29033_, _29034_);
  or g_59643_(_27786_, _29033_, _29035_);
  xor g_59644_(_27786_, _29034_, _29036_);
  or g_59645_(_27792_, _29036_, _29038_);
  not g_59646_(_29038_, _29039_);
  xor g_59647_(_27792_, _29036_, _29040_);
  xor g_59648_(_27793_, _29036_, _29041_);
  or g_59649_(_27789_, _29041_, _29042_);
  xor g_59650_(_27789_, _29040_, _29043_);
  or g_59651_(_26541_, _27797_, _29044_);
  and g_59652_(_27796_, _29044_, _29045_);
  xor g_59653_(_29043_, _29045_, _29046_);
  not g_59654_(_29046_, _29047_);
  or g_59655_(_28841_, _29047_, _29049_);
  xor g_59656_(_28841_, _29046_, _29050_);
  xor g_59657_(_27800_, _29043_, _29051_);
  or g_59658_(_26541_, _27801_, _29052_);
  not g_59659_(_29052_, _29053_);
  or g_59660_(_29051_, _29052_, _29054_);
  xor g_59661_(_29051_, _29053_, _29055_);
  or g_59662_(_26545_, _27801_, _29056_);
  or g_59663_(_29055_, _29056_, _29057_);
  or g_59664_(_28838_, _29050_, _29058_);
  xor g_59665_(_28838_, _29050_, _29060_);
  xor g_59666_(_28840_, _29050_, _29061_);
  or g_59667_(_26550_, _27803_, _29062_);
  or g_59668_(_29061_, _29062_, _29063_);
  xor g_59669_(_29060_, _29062_, _29064_);
  not g_59670_(_29064_, _29065_);
  xor g_59671_(_27812_, _29064_, _29066_);
  xor g_59672_(_27812_, _29065_, _29067_);
  xor g_59673_(_28837_, _29067_, _29068_);
  not g_59674_(_29068_, _29069_);
  and g_59675_(_27821_, _27823_, _29071_);
  or g_59676_(_29068_, _29071_, _29072_);
  xor g_59677_(_29069_, _29071_, _29073_);
  not g_59678_(_29073_, _29074_);
  or g_59679_(_27826_, _29073_, _29075_);
  xor g_59680_(_27826_, _29074_, _29076_);
  and g_59681_(_27829_, _27831_, _29077_);
  xor g_59682_(_29076_, _29077_, _29078_);
  not g_59683_(_29078_, _29079_);
  or g_59684_(_27834_, _29079_, _29080_);
  not g_59685_(_29080_, _29082_);
  xor g_59686_(_27834_, _29078_, _29083_);
  or g_59687_(_27840_, _29083_, _29084_);
  xor g_59688_(_27841_, _29083_, _29085_);
  not g_59689_(_29085_, _29086_);
  and g_59690_(_27836_, _27847_, _29087_);
  xor g_59691_(_29086_, _29087_, _29088_);
  xor g_59692_(_28836_, _29088_, _29089_);
  not g_59693_(_29089_, _29090_);
  or g_59694_(_28833_, _29090_, _29091_);
  xor g_59695_(_28833_, _29089_, _29093_);
  not g_59696_(_29093_, _29094_);
  and g_59697_(_27852_, _27857_, _29095_);
  xor g_59698_(_29094_, _29095_, _29096_);
  or g_59699_(_27856_, _29096_, _29097_);
  xor g_59700_(_27855_, _29096_, _29098_);
  or g_59701_(_27863_, _29098_, _29099_);
  xor g_59702_(_27864_, _29098_, _29100_);
  or g_59703_(_27869_, _29100_, _29101_);
  xor g_59704_(_27870_, _29100_, _29102_);
  or g_59705_(_27866_, _29102_, _29104_);
  xor g_59706_(_27866_, _29102_, _29105_);
  xor g_59707_(_27867_, _29102_, _29106_);
  and g_59708_(_27880_, _29105_, _29107_);
  or g_59709_(_27879_, _29106_, _29108_);
  xor g_59710_(_27879_, _29105_, _29109_);
  not g_59711_(_29109_, _29110_);
  xor g_59712_(_28832_, _29110_, _29111_);
  or g_59713_(_27887_, _29111_, _29112_);
  xor g_59714_(_27887_, _29111_, _29113_);
  and g_59715_(_27897_, _29113_, _29115_);
  xor g_59716_(_27896_, _29113_, _29116_);
  or g_59717_(_27890_, _29116_, _29117_);
  xor g_59718_(_27891_, _29116_, _29118_);
  or g_59719_(_26643_, _27892_, _29119_);
  and g_59720_(_29118_, _29119_, _29120_);
  and g_59721_(_28831_, _29120_, _29121_);
  or g_59722_(_29118_, _29119_, _29122_);
  or g_59723_(_28831_, _29116_, _29123_);
  not g_59724_(_29123_, _29124_);
  and g_59725_(_29122_, _29123_, _29126_);
  not g_59726_(_29126_, _29127_);
  or g_59727_(_29121_, _29127_, _29128_);
  not g_59728_(_29128_, _29129_);
  or g_59729_(_27900_, _29128_, _29130_);
  xor g_59730_(_27900_, _29129_, _29131_);
  or g_59731_(_27903_, _29131_, _29132_);
  xor g_59732_(_27904_, _29131_, _29133_);
  or g_59733_(_27910_, _29133_, _29134_);
  xor g_59734_(_27911_, _29133_, _29135_);
  or g_59735_(_27907_, _29135_, _29137_);
  xor g_59736_(_27908_, _29135_, _29138_);
  not g_59737_(_29138_, _29139_);
  or g_59738_(_26662_, _27919_, _29140_);
  and g_59739_(_27917_, _29140_, _29141_);
  xor g_59740_(_29139_, _29141_, _29142_);
  or g_59741_(_28830_, _29142_, _29143_);
  not g_59742_(_29143_, _29144_);
  xor g_59743_(_28830_, _29142_, _29145_);
  not g_59744_(_29145_, _29146_);
  or g_59745_(_26669_, _27922_, _29148_);
  not g_59746_(_29148_, _29149_);
  and g_59747_(_29145_, _29149_, _29150_);
  or g_59748_(_29146_, _29148_, _29151_);
  xor g_59749_(_29145_, _29149_, _29152_);
  and g_59750_(_28829_, _29152_, _29153_);
  xor g_59751_(_28827_, _29152_, _29154_);
  and g_59752_(_27924_, _27929_, _29155_);
  xor g_59753_(_29154_, _29155_, _29156_);
  and g_59754_(_27928_, _29156_, _29157_);
  not g_59755_(_29157_, _29159_);
  xor g_59756_(_27928_, _29156_, _29160_);
  not g_59757_(_29160_, _29161_);
  or g_59758_(_27932_, _29161_, _29162_);
  xor g_59759_(_27932_, _29160_, _29163_);
  or g_59760_(_28825_, _29163_, _29164_);
  xor g_59761_(_28826_, _29163_, _29165_);
  or g_59762_(_28823_, _29165_, _29166_);
  xor g_59763_(_28824_, _29165_, _29167_);
  xor g_59764_(_27942_, _29167_, _29168_);
  xor g_59765_(_27941_, _29167_, _29170_);
  or g_59766_(_27951_, _29168_, _29171_);
  or g_59767_(_27946_, _29168_, _29172_);
  and g_59768_(_29171_, _29172_, _29173_);
  or g_59769_(_27945_, _29170_, _29174_);
  or g_59770_(_27950_, _29174_, _29175_);
  and g_59771_(_29173_, _29175_, _29176_);
  not g_59772_(_29176_, _29177_);
  or g_59773_(_28821_, _29177_, _29178_);
  xor g_59774_(_28822_, _29176_, _29179_);
  xor g_59775_(_28821_, _29176_, _29181_);
  or g_59776_(_28820_, _29181_, _29182_);
  xor g_59777_(_28820_, _29179_, _29183_);
  or g_59778_(_28818_, _29183_, _29184_);
  xor g_59779_(_28818_, _29183_, _29185_);
  xor g_59780_(_28819_, _29183_, _29186_);
  or g_59781_(_28816_, _29186_, _29187_);
  xor g_59782_(_28816_, _29185_, _29188_);
  not g_59783_(_29188_, _29189_);
  xor g_59784_(_27962_, _29188_, _29190_);
  xor g_59785_(_27962_, _29189_, _29192_);
  or g_59786_(_27965_, _29192_, _29193_);
  xor g_59787_(_27965_, _29190_, _29194_);
  or g_59788_(_26726_, _27964_, _29195_);
  and g_59789_(_29194_, _29195_, _29196_);
  or g_59790_(_29194_, _29195_, _29197_);
  not g_59791_(_29197_, _29198_);
  xor g_59792_(_29194_, _29195_, _29199_);
  or g_59793_(_29196_, _29198_, _29200_);
  or g_59794_(_28815_, _29200_, _29201_);
  not g_59795_(_29201_, _29203_);
  xor g_59796_(_28815_, _29199_, _29204_);
  not g_59797_(_29204_, _29205_);
  or g_59798_(_28814_, _29204_, _29206_);
  not g_59799_(_29206_, _29207_);
  xor g_59800_(_28814_, _29205_, _29208_);
  or g_59801_(_26733_, _27969_, _29209_);
  not g_59802_(_29209_, _29210_);
  or g_59803_(_29208_, _29209_, _29211_);
  xor g_59804_(_29208_, _29210_, _29212_);
  not g_59805_(_29212_, _29214_);
  and g_59806_(_27972_, _27974_, _29215_);
  xor g_59807_(_29214_, _29215_, _29216_);
  or g_59808_(_28813_, _29216_, _29217_);
  not g_59809_(_29217_, _29218_);
  xor g_59810_(_28813_, _29216_, _29219_);
  not g_59811_(_29219_, _29220_);
  or g_59812_(_28812_, _29220_, _29221_);
  not g_59813_(_29221_, _29222_);
  xor g_59814_(_28812_, _29219_, _29223_);
  or g_59815_(_27984_, _29223_, _29225_);
  not g_59816_(_29225_, _29226_);
  xor g_59817_(_27983_, _29223_, _29227_);
  or g_59818_(_27980_, _29227_, _29228_);
  not g_59819_(_29228_, _29229_);
  xor g_59820_(_27979_, _29227_, _29230_);
  not g_59821_(_29230_, _29231_);
  and g_59822_(_27986_, _27988_, _29232_);
  xor g_59823_(_29231_, _29232_, _29233_);
  not g_59824_(_29233_, _29234_);
  or g_59825_(_27989_, _29233_, _29236_);
  xor g_59826_(_27989_, _29234_, _29237_);
  not g_59827_(_29237_, _29238_);
  and g_59828_(_27995_, _27998_, _29239_);
  xor g_59829_(_29238_, _29239_, _29240_);
  or g_59830_(_28002_, _29240_, _29241_);
  xor g_59831_(_28002_, _29240_, _29242_);
  xor g_59832_(_28003_, _29240_, _29243_);
  or g_59833_(_28811_, _29243_, _29244_);
  xor g_59834_(_28811_, _29242_, _29245_);
  or g_59835_(_28809_, _29245_, _29247_);
  not g_59836_(_29247_, _29248_);
  xor g_59837_(_28810_, _29245_, _29249_);
  or g_59838_(_28014_, _29249_, _29250_);
  not g_59839_(_29250_, _29251_);
  xor g_59840_(_28013_, _29249_, _29252_);
  not g_59841_(_29252_, _29253_);
  and g_59842_(_28011_, _29253_, _29254_);
  or g_59843_(_28012_, _29252_, _29255_);
  xor g_59844_(_28012_, _29252_, _29256_);
  xor g_59845_(_28011_, _29252_, _29258_);
  or g_59846_(_28808_, _29258_, _29259_);
  xor g_59847_(_28808_, _29256_, _29260_);
  or g_59848_(_28805_, _29260_, _29261_);
  xor g_59849_(_28807_, _29260_, _29262_);
  and g_59850_(_28018_, _28021_, _29263_);
  not g_59851_(_29263_, _29264_);
  xor g_59852_(_29262_, _29264_, _29265_);
  or g_59853_(_28028_, _29265_, _29266_);
  xor g_59854_(_28029_, _29265_, _29267_);
  or g_59855_(_28024_, _29267_, _29269_);
  xor g_59856_(_28025_, _29267_, _29270_);
  and g_59857_(_28034_, _28040_, _29271_);
  xor g_59858_(_29270_, _29271_, _29272_);
  not g_59859_(_29272_, _29273_);
  xor g_59860_(_28038_, _29272_, _29274_);
  xor g_59861_(_28804_, _29274_, _29275_);
  and g_59862_(_28054_, _29275_, _29276_);
  xor g_59863_(_28053_, _29275_, _29277_);
  not g_59864_(_29277_, _29278_);
  or g_59865_(_28055_, _29277_, _29280_);
  xor g_59866_(_28055_, _29278_, _29281_);
  not g_59867_(_29281_, _29282_);
  and g_59868_(_28060_, _28062_, _29283_);
  xor g_59869_(_29282_, _29283_, _29284_);
  not g_59870_(_29284_, _29285_);
  or g_59871_(_28066_, _29284_, _29286_);
  xor g_59872_(_28066_, _29285_, _29287_);
  and g_59873_(_28067_, _28074_, _29288_);
  not g_59874_(_29288_, _29289_);
  xor g_59875_(_29287_, _29289_, _29291_);
  or g_59876_(_28076_, _29291_, _29292_);
  not g_59877_(_29292_, _29293_);
  and g_59878_(_28076_, _29291_, _29294_);
  xor g_59879_(_28076_, _29291_, _29295_);
  or g_59880_(_29293_, _29294_, _29296_);
  or g_59881_(_28084_, _29296_, _29297_);
  xor g_59882_(_28084_, _29295_, _29298_);
  or g_59883_(_28087_, _29298_, _29299_);
  xor g_59884_(_28086_, _29298_, _29300_);
  or g_59885_(_26858_, _28085_, _29302_);
  or g_59886_(_29300_, _29302_, _29303_);
  xor g_59887_(_29300_, _29302_, _29304_);
  not g_59888_(_29304_, _29305_);
  and g_59889_(_28803_, _29304_, _29306_);
  or g_59890_(_28802_, _29305_, _29307_);
  xor g_59891_(_28802_, _29304_, _29308_);
  or g_59892_(_28800_, _29308_, _29309_);
  xor g_59893_(_28801_, _29308_, _29310_);
  not g_59894_(_29310_, _29311_);
  or g_59895_(_28799_, _29310_, _29313_);
  xor g_59896_(_28799_, _29310_, _29314_);
  xor g_59897_(_28799_, _29311_, _29315_);
  or g_59898_(_28096_, _29315_, _29316_);
  xor g_59899_(_28096_, _29314_, _29317_);
  or g_59900_(_28100_, _29317_, _29318_);
  not g_59901_(_29318_, _29319_);
  xor g_59902_(_28099_, _29317_, _29320_);
  or g_59903_(_26878_, _28098_, _29321_);
  not g_59904_(_29321_, _29322_);
  or g_59905_(_29320_, _29321_, _29324_);
  xor g_59906_(_29320_, _29322_, _29325_);
  or g_59907_(_26880_, _28101_, _29326_);
  not g_59908_(_29326_, _29327_);
  or g_59909_(_29325_, _29326_, _29328_);
  xor g_59910_(_29325_, _29326_, _29329_);
  xor g_59911_(_29325_, _29327_, _29330_);
  or g_59912_(_28107_, _29330_, _29331_);
  xor g_59913_(_28107_, _29329_, _29332_);
  not g_59914_(_29332_, _29333_);
  or g_59915_(_26886_, _28106_, _29335_);
  or g_59916_(_29332_, _29335_, _29336_);
  xor g_59917_(_29332_, _29335_, _29337_);
  xor g_59918_(_29333_, _29335_, _29338_);
  or g_59919_(_26889_, _28108_, _29339_);
  or g_59920_(_29338_, _29339_, _29340_);
  xor g_59921_(_29337_, _29339_, _29341_);
  or g_59922_(_28117_, _29341_, _29342_);
  xor g_59923_(_28118_, _29341_, _29343_);
  not g_59924_(_29343_, _29344_);
  or g_59925_(_26897_, _28120_, _29346_);
  and g_59926_(_28112_, _29346_, _29347_);
  xor g_59927_(_29344_, _29347_, _29348_);
  or g_59928_(_28798_, _29348_, _29349_);
  xor g_59929_(_28798_, _29348_, _29350_);
  not g_59930_(_29350_, _29351_);
  and g_59931_(_28126_, _29350_, _29352_);
  or g_59932_(_28124_, _29351_, _29353_);
  xor g_59933_(_28124_, _29350_, _29354_);
  or g_59934_(_28797_, _29354_, _29355_);
  xor g_59935_(_28797_, _29354_, _29357_);
  not g_59936_(_29357_, _29358_);
  or g_59937_(_28796_, _29358_, _29359_);
  not g_59938_(_29359_, _29360_);
  xor g_59939_(_28796_, _29357_, _29361_);
  not g_59940_(_29361_, _29362_);
  or g_59941_(_28132_, _29361_, _29363_);
  not g_59942_(_29363_, _29364_);
  and g_59943_(_28137_, _29362_, _29365_);
  not g_59944_(_29365_, _29366_);
  xor g_59945_(_28137_, _29361_, _29368_);
  and g_59946_(_28132_, _29368_, _29369_);
  or g_59947_(_29364_, _29369_, _29370_);
  or g_59948_(_28140_, _29370_, _29371_);
  not g_59949_(_29371_, _29372_);
  xor g_59950_(_28140_, _29370_, _29373_);
  not g_59951_(_29373_, _29374_);
  or g_59952_(_28148_, _29374_, _29375_);
  not g_59953_(_29375_, _29376_);
  xor g_59954_(_28148_, _29373_, _29377_);
  or g_59955_(_28145_, _29377_, _29379_);
  not g_59956_(_29379_, _29380_);
  xor g_59957_(_28144_, _29377_, _29381_);
  or g_59958_(_28154_, _29374_, _29382_);
  not g_59959_(_29382_, _29383_);
  xor g_59960_(_28155_, _29381_, _29384_);
  and g_59961_(_28160_, _28166_, _29385_);
  xor g_59962_(_29384_, _29385_, _29386_);
  not g_59963_(_29386_, _29387_);
  and g_59964_(_28165_, _29386_, _29388_);
  or g_59965_(_28164_, _29387_, _29390_);
  xor g_59966_(_28164_, _29386_, _29391_);
  or g_59967_(_28168_, _29391_, _29392_);
  not g_59968_(_29392_, _29393_);
  and g_59969_(_28168_, _29391_, _29394_);
  or g_59970_(_29393_, _29394_, _29395_);
  and g_59971_(_28794_, _29395_, _29396_);
  or g_59972_(_28794_, _29395_, _29397_);
  not g_59973_(_29397_, _29398_);
  xor g_59974_(_28794_, _29395_, _29399_);
  or g_59975_(_29396_, _29398_, _29401_);
  or g_59976_(_26945_, _28170_, _29402_);
  or g_59977_(_29401_, _29402_, _29403_);
  not g_59978_(_29403_, _29404_);
  xor g_59979_(_29399_, _29402_, _29405_);
  or g_59980_(_28175_, _29405_, _29406_);
  xor g_59981_(_28176_, _29405_, _29407_);
  xor g_59982_(_28186_, _29407_, _29408_);
  or g_59983_(_28793_, _29408_, _29409_);
  not g_59984_(_29409_, _29410_);
  xor g_59985_(_28793_, _29408_, _29412_);
  not g_59986_(_29412_, _29413_);
  or g_59987_(_28792_, _29413_, _29414_);
  xor g_59988_(_28792_, _29412_, _29415_);
  not g_59989_(_29415_, _29416_);
  or g_59990_(_28791_, _29415_, _29417_);
  xor g_59991_(_28791_, _29416_, _29418_);
  and g_59992_(_28790_, _29418_, _29419_);
  or g_59993_(_28790_, _29418_, _29420_);
  not g_59994_(_29420_, _29421_);
  xor g_59995_(_28790_, _29418_, _29423_);
  or g_59996_(_29419_, _29421_, _29424_);
  or g_59997_(_28198_, _29424_, _29425_);
  xor g_59998_(_28198_, _29423_, _29426_);
  not g_59999_(_29426_, _29427_);
  and g_60000_(_28204_, _28209_, _29428_);
  xor g_60001_(_29427_, _29428_, _29429_);
  xor g_60002_(_29426_, _29428_, _29430_);
  or g_60003_(_28208_, _29429_, _29431_);
  not g_60004_(_29431_, _29432_);
  xor g_60005_(_28208_, _29430_, _29434_);
  not g_60006_(_29434_, _29435_);
  and g_60007_(_28212_, _28215_, _29436_);
  xor g_60008_(_29434_, _29436_, _29437_);
  xor g_60009_(_29435_, _29436_, _29438_);
  or g_60010_(_28789_, _29438_, _29439_);
  xor g_60011_(_28789_, _29438_, _29440_);
  xor g_60012_(_28789_, _29437_, _29441_);
  and g_60013_(_28787_, _29440_, _29442_);
  or g_60014_(_28788_, _29441_, _29443_);
  xor g_60015_(_28787_, _29441_, _29445_);
  not g_60016_(_29445_, _29446_);
  and g_60017_(_28222_, _29446_, _29447_);
  not g_60018_(_29447_, _29448_);
  xor g_60019_(_28221_, _29445_, _29449_);
  xor g_60020_(_28222_, _29445_, _29450_);
  or g_60021_(_28223_, _29450_, _29451_);
  xor g_60022_(_28223_, _29449_, _29452_);
  not g_60023_(_29452_, _29453_);
  or g_60024_(_28227_, _29452_, _29454_);
  xor g_60025_(_28227_, _29453_, _29456_);
  and g_60026_(_28232_, _29456_, _29457_);
  or g_60027_(_28232_, _29456_, _29458_);
  not g_60028_(_29458_, _29459_);
  xor g_60029_(_28232_, _29456_, _29460_);
  or g_60030_(_29457_, _29459_, _29461_);
  or g_60031_(_28230_, _29461_, _29462_);
  not g_60032_(_29462_, _29463_);
  xor g_60033_(_28230_, _29460_, _29464_);
  not g_60034_(_29464_, _29465_);
  and g_60035_(_28234_, _28238_, _29467_);
  xor g_60036_(_29465_, _29467_, _29468_);
  xor g_60037_(_28786_, _29468_, _29469_);
  or g_60038_(_28250_, _29469_, _29470_);
  not g_60039_(_29470_, _29471_);
  xor g_60040_(_28251_, _29469_, _29472_);
  not g_60041_(_29472_, _29473_);
  or g_60042_(_28252_, _29472_, _29474_);
  xor g_60043_(_28252_, _29472_, _29475_);
  xor g_60044_(_28252_, _29473_, _29476_);
  or g_60045_(_28258_, _29476_, _29478_);
  xor g_60046_(_28258_, _29475_, _29479_);
  or g_60047_(_28263_, _29479_, _29480_);
  xor g_60048_(_28264_, _29479_, _29481_);
  or g_60049_(_28262_, _29481_, _29482_);
  xor g_60050_(_28261_, _29481_, _29483_);
  not g_60051_(_29483_, _29484_);
  and g_60052_(_28275_, _29484_, _29485_);
  not g_60053_(_29485_, _29486_);
  xor g_60054_(_28275_, _29484_, _29487_);
  xor g_60055_(_28275_, _29483_, _29489_);
  or g_60056_(_27046_, _28278_, _29490_);
  and g_60057_(_28272_, _29490_, _29491_);
  xor g_60058_(_29487_, _29491_, _29492_);
  or g_60059_(_28783_, _29492_, _29493_);
  xor g_60060_(_28783_, _29492_, _29494_);
  not g_60061_(_29494_, _29495_);
  and g_60062_(_28284_, _28287_, _29496_);
  xor g_60063_(_29494_, _29496_, _29497_);
  or g_60064_(_28291_, _29497_, _29498_);
  xor g_60065_(_28291_, _29497_, _29500_);
  not g_60066_(_29500_, _29501_);
  or g_60067_(_28293_, _29501_, _29502_);
  xor g_60068_(_28293_, _29500_, _29503_);
  not g_60069_(_29503_, _29504_);
  or g_60070_(_28302_, _29503_, _29505_);
  xor g_60071_(_28302_, _29504_, _29506_);
  or g_60072_(_28303_, _29506_, _29507_);
  not g_60073_(_29507_, _29508_);
  xor g_60074_(_28304_, _29506_, _29509_);
  not g_60075_(_29509_, _29511_);
  and g_60076_(_28308_, _28314_, _29512_);
  xor g_60077_(_29511_, _29512_, _29513_);
  or g_60078_(_28782_, _29513_, _29514_);
  xor g_60079_(_28782_, _29513_, _29515_);
  not g_60080_(_29515_, _29516_);
  or g_60081_(_28320_, _29516_, _29517_);
  not g_60082_(_29517_, _29518_);
  xor g_60083_(_28320_, _29515_, _29519_);
  or g_60084_(_28325_, _29519_, _29520_);
  xor g_60085_(_28325_, _29519_, _29522_);
  not g_60086_(_29522_, _29523_);
  or g_60087_(_28329_, _29523_, _29524_);
  xor g_60088_(_28329_, _29522_, _29525_);
  or g_60089_(_28335_, _28338_, _29526_);
  xor g_60090_(_29525_, _29526_, _29527_);
  xor g_60091_(_28781_, _29527_, _29528_);
  xor g_60092_(_28780_, _29527_, _29529_);
  or g_60093_(_28779_, _29528_, _29530_);
  xor g_60094_(_28779_, _29529_, _29531_);
  or g_60095_(_27112_, _28347_, _29533_);
  or g_60096_(_29531_, _29533_, _29534_);
  xor g_60097_(_29531_, _29533_, _29535_);
  xor g_60098_(_28351_, _29535_, _29536_);
  not g_60099_(_29536_, _29537_);
  or g_60100_(_28778_, _29537_, _29538_);
  not g_60101_(_29538_, _29539_);
  xor g_60102_(_28778_, _29536_, _29540_);
  or g_60103_(_27126_, _28352_, _29541_);
  not g_60104_(_29541_, _29542_);
  or g_60105_(_29540_, _29541_, _29544_);
  xor g_60106_(_29540_, _29542_, _29545_);
  or g_60107_(_28360_, _29545_, _29546_);
  not g_60108_(_29546_, _29547_);
  xor g_60109_(_28360_, _29545_, _29548_);
  not g_60110_(_29548_, _29549_);
  and g_60111_(_28364_, _29548_, _29550_);
  not g_60112_(_29550_, _29551_);
  and g_60113_(_28359_, _29548_, _29552_);
  or g_60114_(_28358_, _29549_, _29553_);
  xor g_60115_(_28358_, _29548_, _29555_);
  and g_60116_(_28363_, _29555_, _29556_);
  or g_60117_(_29550_, _29556_, _29557_);
  not g_60118_(_29557_, _29558_);
  and g_60119_(_28371_, _28375_, _29559_);
  xor g_60120_(_29558_, _29559_, _29560_);
  xor g_60121_(_29557_, _29559_, _29561_);
  and g_60122_(_28379_, _29560_, _29562_);
  or g_60123_(_28380_, _29561_, _29563_);
  and g_60124_(_28776_, _29562_, _29564_);
  or g_60125_(_28777_, _29563_, _29566_);
  or g_60126_(_28776_, _29560_, _29567_);
  or g_60127_(_28379_, _29560_, _29568_);
  not g_60128_(_29568_, _29569_);
  and g_60129_(_29567_, _29568_, _29570_);
  not g_60130_(_29570_, _29571_);
  and g_60131_(_29566_, _29570_, _29572_);
  or g_60132_(_29564_, _29571_, _29573_);
  or g_60133_(_28775_, _29573_, _29574_);
  xor g_60134_(_28775_, _29572_, _29575_);
  or g_60135_(_28385_, _29575_, _29577_);
  xor g_60136_(_28386_, _29575_, _29578_);
  or g_60137_(_28390_, _29578_, _29579_);
  xor g_60138_(_28391_, _29578_, _29580_);
  not g_60139_(_29580_, _29581_);
  and g_60140_(_28395_, _29581_, _29582_);
  or g_60141_(_28394_, _29580_, _29583_);
  xor g_60142_(_28395_, _29580_, _29584_);
  not g_60143_(_29584_, _29585_);
  and g_60144_(_28398_, _28402_, _29586_);
  xor g_60145_(_29584_, _29586_, _29588_);
  xor g_60146_(_29585_, _29586_, _29589_);
  or g_60147_(_27176_, _28401_, _29590_);
  not g_60148_(_29590_, _29591_);
  or g_60149_(_27179_, _28403_, _29592_);
  not g_60150_(_29592_, _29593_);
  and g_60151_(_29590_, _29592_, _29594_);
  xor g_60152_(_29588_, _29594_, _29595_);
  xor g_60153_(_29589_, _29594_, _29596_);
  and g_60154_(_28774_, _29596_, _29597_);
  or g_60155_(_28772_, _29595_, _29599_);
  xor g_60156_(_28772_, _29595_, _29600_);
  not g_60157_(_29600_, _29601_);
  or g_60158_(_27186_, _28406_, _29602_);
  or g_60159_(_29601_, _29602_, _29603_);
  xor g_60160_(_29601_, _29602_, _29604_);
  xor g_60161_(_29600_, _29602_, _29605_);
  and g_60162_(_28409_, _28417_, _29606_);
  xor g_60163_(_29604_, _29606_, _29607_);
  or g_60164_(_28414_, _29607_, _29608_);
  xor g_60165_(_28413_, _29607_, _29610_);
  not g_60166_(_29610_, _29611_);
  or g_60167_(_28421_, _29610_, _29612_);
  xor g_60168_(_28421_, _29611_, _29613_);
  not g_60169_(_29613_, _29614_);
  xor g_60170_(_28427_, _29614_, _29615_);
  or g_60171_(_28431_, _29615_, _29616_);
  xor g_60172_(_28431_, _29615_, _29617_);
  xor g_60173_(_28430_, _29615_, _29618_);
  or g_60174_(_28437_, _29618_, _29619_);
  xor g_60175_(_28437_, _29617_, _29621_);
  not g_60176_(_29621_, _29622_);
  or g_60177_(_28438_, _29621_, _29623_);
  xor g_60178_(_28438_, _29622_, _29624_);
  not g_60179_(_29624_, _29625_);
  or g_60180_(_28439_, _29624_, _29626_);
  xor g_60181_(_28439_, _29625_, _29627_);
  not g_60182_(_29627_, _29628_);
  or g_60183_(_28771_, _29627_, _29629_);
  xor g_60184_(_28771_, _29627_, _29630_);
  xor g_60185_(_28771_, _29628_, _29632_);
  or g_60186_(_28770_, _29632_, _29633_);
  xor g_60187_(_28770_, _29630_, _29634_);
  and g_60188_(_28446_, _28450_, _29635_);
  xor g_60189_(_29634_, _29635_, _29636_);
  not g_60190_(_29636_, _29637_);
  or g_60191_(_28449_, _29637_, _29638_);
  xor g_60192_(_28449_, _29636_, _29639_);
  not g_60193_(_29639_, _29640_);
  or g_60194_(_28454_, _29639_, _29641_);
  xor g_60195_(_28454_, _29640_, _29643_);
  or g_60196_(_28458_, _29643_, _29644_);
  xor g_60197_(_28459_, _29643_, _29645_);
  not g_60198_(_29645_, _29646_);
  or g_60199_(_27245_, _28464_, _29647_);
  and g_60200_(_28462_, _29647_, _29648_);
  xor g_60201_(_29645_, _29648_, _29649_);
  xor g_60202_(_29646_, _29648_, _29650_);
  or g_60203_(_28769_, _29650_, _29651_);
  xor g_60204_(_28769_, _29649_, _29652_);
  or g_60205_(_28471_, _29652_, _29654_);
  xor g_60206_(_28470_, _29652_, _29655_);
  or g_60207_(_28472_, _29655_, _29656_);
  xor g_60208_(_28473_, _29655_, _29657_);
  not g_60209_(_29657_, _29658_);
  or g_60210_(_28483_, _29657_, _29659_);
  xor g_60211_(_28483_, _29657_, _29660_);
  xor g_60212_(_28483_, _29658_, _29661_);
  or g_60213_(_28484_, _29661_, _29662_);
  xor g_60214_(_28484_, _29660_, _29663_);
  or g_60215_(_28480_, _29663_, _29665_);
  xor g_60216_(_28481_, _29663_, _29666_);
  or g_60217_(_28486_, _29666_, _29667_);
  xor g_60218_(_28487_, _29666_, _29668_);
  or g_60219_(_27271_, _28482_, _29669_);
  not g_60220_(_29669_, _29670_);
  or g_60221_(_29668_, _29669_, _29671_);
  xor g_60222_(_29668_, _29669_, _29672_);
  xor g_60223_(_29668_, _29670_, _29673_);
  or g_60224_(_27274_, _28489_, _29674_);
  or g_60225_(_29673_, _29674_, _29676_);
  xor g_60226_(_29672_, _29674_, _29677_);
  not g_60227_(_29677_, _29678_);
  or g_60228_(_28768_, _29677_, _29679_);
  xor g_60229_(_28768_, _29677_, _29680_);
  xor g_60230_(_28768_, _29678_, _29681_);
  or g_60231_(_27280_, _28492_, _29682_);
  and g_60232_(_28496_, _29682_, _29683_);
  xor g_60233_(_29681_, _29683_, _29684_);
  xor g_60234_(_29680_, _29683_, _29685_);
  or g_60235_(_28502_, _29685_, _29687_);
  not g_60236_(_29687_, _29688_);
  xor g_60237_(_28503_, _29684_, _29689_);
  xor g_60238_(_28502_, _29684_, _29690_);
  and g_60239_(_27291_, _28497_, _29691_);
  not g_60240_(_29691_, _29692_);
  and g_60241_(_29689_, _29691_, _29693_);
  or g_60242_(_29690_, _29692_, _29694_);
  xor g_60243_(_29690_, _29691_, _29695_);
  or g_60244_(_28766_, _29695_, _29696_);
  xor g_60245_(_28767_, _29695_, _29698_);
  not g_60246_(_29698_, _29699_);
  and g_60247_(_28509_, _28515_, _29700_);
  xor g_60248_(_29699_, _29700_, _29701_);
  or g_60249_(_28514_, _29701_, _29702_);
  xor g_60250_(_28513_, _29701_, _29703_);
  or g_60251_(_28524_, _29703_, _29704_);
  xor g_60252_(_28524_, _29703_, _29705_);
  xor g_60253_(_28525_, _29703_, _29706_);
  or g_60254_(_28531_, _29706_, _29707_);
  not g_60255_(_29707_, _29709_);
  or g_60256_(_28535_, _29706_, _29710_);
  xor g_60257_(_28535_, _29706_, _29711_);
  xor g_60258_(_28535_, _29705_, _29712_);
  and g_60259_(_28531_, _29712_, _29713_);
  or g_60260_(_28530_, _29711_, _29714_);
  and g_60261_(_29707_, _29714_, _29715_);
  or g_60262_(_29709_, _29713_, _29716_);
  or g_60263_(_28538_, _29716_, _29717_);
  xor g_60264_(_28538_, _29715_, _29718_);
  or g_60265_(_27319_, _28536_, _29720_);
  not g_60266_(_29720_, _29721_);
  or g_60267_(_29718_, _29720_, _29722_);
  not g_60268_(_29722_, _29723_);
  xor g_60269_(_29718_, _29720_, _29724_);
  xor g_60270_(_29718_, _29721_, _29725_);
  or g_60271_(_28765_, _29725_, _29726_);
  xor g_60272_(_28765_, _29724_, _29727_);
  or g_60273_(_28764_, _29727_, _29728_);
  not g_60274_(_29728_, _29729_);
  xor g_60275_(_28764_, _29727_, _29731_);
  xor g_60276_(_28763_, _29727_, _29732_);
  or g_60277_(_28761_, _29732_, _29733_);
  not g_60278_(_29733_, _29734_);
  xor g_60279_(_28761_, _29731_, _29735_);
  not g_60280_(_29735_, _29736_);
  and g_60281_(_28547_, _28550_, _29737_);
  or g_60282_(_29735_, _29737_, _29738_);
  xor g_60283_(_29735_, _29737_, _29739_);
  xor g_60284_(_29736_, _29737_, _29740_);
  or g_60285_(_28760_, _29740_, _29742_);
  xor g_60286_(_28760_, _29739_, _29743_);
  or g_60287_(_28759_, _29743_, _29744_);
  or g_60288_(_27343_, _28551_, _29745_);
  or g_60289_(_29743_, _29745_, _29746_);
  xor g_60290_(_29743_, _29745_, _29747_);
  or g_60291_(_28758_, _29747_, _29748_);
  and g_60292_(_29744_, _29748_, _29749_);
  and g_60293_(_28757_, _29749_, _29750_);
  xor g_60294_(_28757_, _29749_, _29751_);
  xor g_60295_(_28756_, _29749_, _29753_);
  or g_60296_(_27353_, _28558_, _29754_);
  or g_60297_(_29753_, _29754_, _29755_);
  xor g_60298_(_29753_, _29754_, _29756_);
  xor g_60299_(_29751_, _29754_, _29757_);
  or g_60300_(_28755_, _29757_, _29758_);
  xor g_60301_(_28755_, _29756_, _29759_);
  not g_60302_(_29759_, _29760_);
  or g_60303_(_28563_, _29759_, _29761_);
  xor g_60304_(_28563_, _29760_, _29762_);
  or g_60305_(_27364_, _28564_, _29764_);
  and g_60306_(_28561_, _29764_, _29765_);
  xor g_60307_(_29762_, _29765_, _29766_);
  not g_60308_(_29766_, _29767_);
  and g_60309_(_28754_, _29766_, _29768_);
  or g_60310_(_28753_, _29767_, _29769_);
  xor g_60311_(_28754_, _29766_, _29770_);
  xor g_60312_(_28753_, _29766_, _29771_);
  or g_60313_(_28568_, _29771_, _29772_);
  not g_60314_(_29772_, _29773_);
  xor g_60315_(_28568_, _29770_, _29775_);
  or g_60316_(_28571_, _29775_, _29776_);
  xor g_60317_(_28572_, _29775_, _29777_);
  or g_60318_(_27375_, _28569_, _29778_);
  or g_60319_(_29777_, _29778_, _29779_);
  xor g_60320_(_29777_, _29778_, _29780_);
  not g_60321_(_29780_, _29781_);
  or g_60322_(_28752_, _29781_, _29782_);
  xor g_60323_(_28752_, _29780_, _29783_);
  not g_60324_(_29783_, _29784_);
  or g_60325_(_28581_, _29783_, _29786_);
  xor g_60326_(_28581_, _29783_, _29787_);
  xor g_60327_(_28581_, _29784_, _29788_);
  or g_60328_(_28579_, _29788_, _29789_);
  not g_60329_(_29789_, _29790_);
  xor g_60330_(_28579_, _29787_, _29791_);
  and g_60331_(_28584_, _29791_, _29792_);
  and g_60332_(_28588_, _29792_, _29793_);
  or g_60333_(_28588_, _29791_, _29794_);
  or g_60334_(_28584_, _29788_, _29795_);
  not g_60335_(_29795_, _29797_);
  and g_60336_(_29794_, _29795_, _29798_);
  not g_60337_(_29798_, _29799_);
  or g_60338_(_29793_, _29799_, _29800_);
  or g_60339_(_28589_, _29800_, _29801_);
  xor g_60340_(_28589_, _29800_, _29802_);
  xor g_60341_(_28590_, _29800_, _29803_);
  and g_60342_(_28594_, _28600_, _29804_);
  xor g_60343_(_29802_, _29804_, _29805_);
  xor g_60344_(_29803_, _29804_, _29806_);
  or g_60345_(_28601_, _29805_, _29808_);
  xor g_60346_(_28601_, _29806_, _29809_);
  not g_60347_(_29809_, _29810_);
  or g_60348_(_28750_, _29809_, _29811_);
  xor g_60349_(_28750_, _29810_, _29812_);
  not g_60350_(_29812_, _29813_);
  or g_60351_(_28749_, _29812_, _29814_);
  xor g_60352_(_28749_, _29813_, _29815_);
  or g_60353_(_27412_, _28605_, _29816_);
  or g_60354_(_29815_, _29816_, _29817_);
  xor g_60355_(_29815_, _29816_, _29819_);
  not g_60356_(_29819_, _29820_);
  and g_60357_(_28748_, _29819_, _29821_);
  or g_60358_(_28747_, _29820_, _29822_);
  xor g_60359_(_28747_, _29819_, _29823_);
  not g_60360_(_29823_, _29824_);
  or g_60361_(_28610_, _29823_, _29825_);
  xor g_60362_(_28610_, _29823_, _29826_);
  xor g_60363_(_28610_, _29824_, _29827_);
  or g_60364_(_27420_, _28607_, _29828_);
  or g_60365_(_29827_, _29828_, _29830_);
  xor g_60366_(_29826_, _29828_, _29831_);
  and g_60367_(_27425_, _28611_, _29832_);
  or g_60368_(_27424_, _28612_, _29833_);
  or g_60369_(_29831_, _29833_, _29834_);
  not g_60370_(_29834_, _29835_);
  xor g_60371_(_29831_, _29832_, _29836_);
  or g_60372_(_28617_, _29836_, _29837_);
  xor g_60373_(_28618_, _29836_, _29838_);
  not g_60374_(_29838_, _29839_);
  or g_60375_(_28619_, _29838_, _29841_);
  xor g_60376_(_28619_, _29838_, _29842_);
  xor g_60377_(_28619_, _29839_, _29843_);
  or g_60378_(_28623_, _29843_, _29844_);
  xor g_60379_(_28623_, _29842_, _29845_);
  or g_60380_(_28628_, _29845_, _29846_);
  xor g_60381_(_28629_, _29845_, _29847_);
  or g_60382_(_27441_, _28625_, _29848_);
  or g_60383_(_29847_, _29848_, _29849_);
  xor g_60384_(_29847_, _29848_, _29850_);
  not g_60385_(_29850_, _29852_);
  and g_60386_(_28746_, _29850_, _29853_);
  or g_60387_(_28745_, _29852_, _29854_);
  xor g_60388_(_28745_, _29850_, _29855_);
  or g_60389_(_28641_, _29855_, _29856_);
  xor g_60390_(_28641_, _29855_, _29857_);
  not g_60391_(_29857_, _29858_);
  or g_60392_(_28643_, _29858_, _29859_);
  xor g_60393_(_28643_, _29857_, _29860_);
  not g_60394_(_29860_, _29861_);
  or g_60395_(_28639_, _29860_, _29863_);
  xor g_60396_(_28639_, _29861_, _29864_);
  or g_60397_(_28645_, _29864_, _29865_);
  xor g_60398_(_28646_, _29864_, _29866_);
  and g_60399_(_28649_, _28652_, _29867_);
  or g_60400_(_29866_, _29867_, _29868_);
  not g_60401_(_29868_, _29869_);
  and g_60402_(_29866_, _29867_, _29870_);
  or g_60403_(_29869_, _29870_, _29871_);
  or g_60404_(_28656_, _29871_, _29872_);
  xor g_60405_(_28657_, _29871_, _29874_);
  or g_60406_(_28662_, _29874_, _29875_);
  xor g_60407_(_28663_, _29874_, _29876_);
  or g_60408_(_28668_, _29876_, _29877_);
  not g_60409_(_29877_, _29878_);
  or g_60410_(_28659_, _29876_, _29879_);
  xor g_60411_(_28660_, _29876_, _29880_);
  or g_60412_(_28671_, _29880_, _29881_);
  xor g_60413_(_28672_, _29880_, _29882_);
  and g_60414_(_28668_, _29882_, _29883_);
  or g_60415_(_29878_, _29883_, _29885_);
  not g_60416_(_29885_, _29886_);
  or g_60417_(_28678_, _29885_, _29887_);
  xor g_60418_(_28678_, _29885_, _29888_);
  xor g_60419_(_28678_, _29886_, _29889_);
  xor g_60420_(_28688_, _29889_, _29890_);
  not g_60421_(_29890_, _29891_);
  xor g_60422_(_28744_, _29891_, _29892_);
  or g_60423_(_28699_, _29892_, _29893_);
  not g_60424_(_29893_, _29894_);
  xor g_60425_(_28699_, _29892_, _29896_);
  xor g_60426_(_28700_, _29892_, _29897_);
  or g_60427_(_28743_, _29897_, _29898_);
  xor g_60428_(_28743_, _29896_, _29899_);
  not g_60429_(_29899_, _29900_);
  or g_60430_(_28742_, _29899_, _29901_);
  xor g_60431_(_28742_, _29900_, _29902_);
  not g_60432_(_29902_, _29903_);
  or g_60433_(_28741_, _29902_, _29904_);
  xor g_60434_(_28741_, _29902_, _29905_);
  xor g_60435_(_28741_, _29903_, _29907_);
  or g_60436_(_28739_, _29907_, _29908_);
  xor g_60437_(_28739_, _29905_, _29909_);
  or g_60438_(_28738_, _29909_, _29910_);
  xor g_60439_(_28738_, _29909_, _29911_);
  not g_60440_(_29911_, _29912_);
  or g_60441_(_27522_, _28704_, _29913_);
  or g_60442_(_29912_, _29913_, _29914_);
  xor g_60443_(_29911_, _29913_, _29915_);
  or g_60444_(_28709_, _29915_, _29916_);
  xor g_60445_(_28707_, _29915_, _29918_);
  or g_60446_(_27529_, _28710_, _29919_);
  or g_60447_(_29918_, _29919_, _29920_);
  xor g_60448_(_29918_, _29919_, _29921_);
  not g_60449_(_29921_, _29922_);
  or g_60450_(_28737_, _29922_, _29923_);
  xor g_60451_(_28737_, _29921_, _29924_);
  and g_60452_(_28736_, _29924_, _29925_);
  or g_60453_(_28736_, _29924_, _29926_);
  not g_60454_(_29926_, _29927_);
  or g_60455_(_29925_, _29927_, _29929_);
  not g_60456_(_29929_, _29930_);
  or g_60457_(_28735_, _29929_, _29931_);
  xor g_60458_(_28735_, _29929_, _29932_);
  xor g_60459_(_28735_, _29930_, _29933_);
  or g_60460_(_28716_, _29933_, _29934_);
  xor g_60461_(_28716_, _29932_, _29935_);
  or g_60462_(_28721_, _29935_, _29936_);
  not g_60463_(_29936_, _29937_);
  xor g_60464_(_28722_, _29935_, _29938_);
  not g_60465_(_29938_, _29940_);
  and g_60466_(_28727_, _28732_, _29941_);
  xor g_60467_(_29940_, _29941_, _29942_);
  or g_60468_(_28734_, _29942_, _29943_);
  xor g_60469_(_28734_, _29942_, out[642]);
  or g_60470_(_28727_, _29938_, _29944_);
  not g_60471_(_29944_, _29945_);
  and g_60472_(_29908_, _29910_, _29946_);
  and g_60473_(_29901_, _29904_, _29947_);
  or g_60474_(_28701_, _29890_, _29948_);
  or g_60475_(_28691_, _29890_, _29950_);
  not g_60476_(_29950_, _29951_);
  and g_60477_(_28681_, _29888_, _29952_);
  or g_60478_(_28682_, _29889_, _29953_);
  and g_60479_(_28687_, _29888_, _29954_);
  or g_60480_(_28685_, _29889_, _29955_);
  or g_60481_(_28600_, _29803_, _29956_);
  not g_60482_(_29956_, _29957_);
  or g_60483_(_29759_, _29764_, _29958_);
  and g_60484_(_29742_, _29746_, _29959_);
  and g_60485_(_29722_, _29726_, _29961_);
  or g_60486_(_28515_, _29698_, _29962_);
  not g_60487_(_29962_, _29963_);
  or g_60488_(_28509_, _29698_, _29964_);
  and g_60489_(_29696_, _29964_, _29965_);
  or g_60490_(_28496_, _29681_, _29966_);
  not g_60491_(_29966_, _29967_);
  or g_60492_(_29681_, _29682_, _29968_);
  not g_60493_(_29968_, _29969_);
  or g_60494_(_29645_, _29647_, _29970_);
  or g_60495_(_28462_, _29645_, _29972_);
  and g_60496_(_29641_, _29644_, _29973_);
  not g_60497_(_29973_, _29974_);
  or g_60498_(_28425_, _29610_, _29975_);
  not g_60499_(_29975_, _29976_);
  or g_60500_(_28426_, _29613_, _29977_);
  and g_60501_(_28418_, _29604_, _29978_);
  not g_60502_(_29978_, _29979_);
  and g_60503_(_29588_, _29591_, _29980_);
  or g_60504_(_29589_, _29590_, _29981_);
  or g_60505_(_28402_, _29584_, _29983_);
  not g_60506_(_29983_, _29984_);
  or g_60507_(_28398_, _29584_, _29985_);
  not g_60508_(_29985_, _29986_);
  or g_60509_(_28372_, _29557_, _29987_);
  or g_60510_(_27148_, _29987_, _29988_);
  or g_60511_(_28370_, _29557_, _29989_);
  not g_60512_(_29989_, _29990_);
  or g_60513_(_28350_, _29531_, _29991_);
  or g_60514_(_27119_, _29991_, _29992_);
  or g_60515_(_27116_, _29991_, _29994_);
  or g_60516_(_28337_, _29525_, _29995_);
  or g_60517_(_28333_, _29525_, _29996_);
  not g_60518_(_29996_, _29997_);
  or g_60519_(_28314_, _29509_, _29998_);
  not g_60520_(_29998_, _29999_);
  or g_60521_(_27075_, _28305_, _30000_);
  or g_60522_(_29509_, _30000_, _30001_);
  or g_60523_(_27069_, _28305_, _30002_);
  or g_60524_(_29509_, _30002_, _30003_);
  and g_60525_(_29507_, _30003_, _30005_);
  and g_60526_(_29502_, _29505_, _30006_);
  or g_60527_(_29489_, _29490_, _30007_);
  or g_60528_(_28272_, _29489_, _30008_);
  and g_60529_(_29480_, _29482_, _30009_);
  or g_60530_(_28242_, _29468_, _30010_);
  or g_60531_(_28238_, _29464_, _30011_);
  or g_60532_(_28234_, _29464_, _30012_);
  or g_60533_(_28215_, _29434_, _30013_);
  or g_60534_(_28212_, _29434_, _30014_);
  not g_60535_(_30014_, _30016_);
  or g_60536_(_28203_, _29426_, _30017_);
  and g_60537_(_29425_, _30017_, _30018_);
  or g_60538_(_28178_, _29405_, _30019_);
  or g_60539_(_28156_, _29381_, _30020_);
  or g_60540_(_26930_, _30020_, _30021_);
  not g_60541_(_30021_, _30022_);
  or g_60542_(_29343_, _29346_, _30023_);
  not g_60543_(_30023_, _30024_);
  or g_60544_(_28112_, _29343_, _30025_);
  not g_60545_(_30025_, _30027_);
  or g_60546_(_28074_, _29287_, _30028_);
  or g_60547_(_28062_, _29281_, _30029_);
  or g_60548_(_28047_, _29274_, _30030_);
  or g_60549_(_26821_, _30030_, _30031_);
  or g_60550_(_28045_, _29274_, _30032_);
  or g_60551_(_28040_, _29270_, _30033_);
  or g_60552_(_26810_, _29267_, _30034_);
  or g_60553_(_28032_, _30034_, _30035_);
  not g_60554_(_30035_, _30036_);
  or g_60555_(_28021_, _29262_, _30038_);
  or g_60556_(_28018_, _29262_, _30039_);
  not g_60557_(_30039_, _30040_);
  or g_60558_(_27998_, _29237_, _30041_);
  or g_60559_(_27988_, _29230_, _30042_);
  or g_60560_(_27986_, _29230_, _30043_);
  not g_60561_(_30043_, _30044_);
  or g_60562_(_27974_, _29212_, _30045_);
  not g_60563_(_30045_, _30046_);
  or g_60564_(_27972_, _29212_, _30047_);
  or g_60565_(_27937_, _29167_, _30049_);
  or g_60566_(_26695_, _30049_, _30050_);
  not g_60567_(_30050_, _30051_);
  or g_60568_(_27929_, _29154_, _30052_);
  not g_60569_(_30052_, _30053_);
  or g_60570_(_27924_, _29154_, _30054_);
  or g_60571_(_29150_, _29153_, _30055_);
  or g_60572_(_27917_, _29133_, _30056_);
  and g_60573_(_29117_, _29122_, _30057_);
  or g_60574_(_27881_, _29106_, _30058_);
  or g_60575_(_27876_, _29100_, _30060_);
  or g_60576_(_27857_, _29093_, _30061_);
  or g_60577_(_27852_, _29093_, _30062_);
  not g_60578_(_30062_, _30063_);
  or g_60579_(_28834_, _29088_, _30064_);
  or g_60580_(_28835_, _29088_, _30065_);
  or g_60581_(_27847_, _29085_, _30066_);
  or g_60582_(_27836_, _29085_, _30067_);
  and g_60583_(_29084_, _30067_, _30068_);
  or g_60584_(_27829_, _29076_, _30069_);
  and g_60585_(_29075_, _30069_, _30071_);
  or g_60586_(_27818_, _29066_, _30072_);
  or g_60587_(_27814_, _29064_, _30073_);
  or g_60588_(_27810_, _29064_, _30074_);
  or g_60589_(_27808_, _29064_, _30075_);
  or g_60590_(_27796_, _29043_, _30076_);
  and g_60591_(_29042_, _30076_, _30077_);
  not g_60592_(_30077_, _30078_);
  and g_60593_(_29029_, _29032_, _30079_);
  or g_60594_(_27772_, _29027_, _30080_);
  or g_60595_(_27769_, _29024_, _30082_);
  or g_60596_(_27763_, _29024_, _30083_);
  or g_60597_(_26508_, _30083_, _30084_);
  or g_60598_(_27750_, _29012_, _30085_);
  or g_60599_(_27738_, _29001_, _30086_);
  not g_60600_(_30086_, _30087_);
  and g_60601_(_27732_, _28999_, _30088_);
  or g_60602_(_29000_, _30088_, _30089_);
  or g_60603_(_27700_, _28976_, _30090_);
  or g_60604_(_27648_, _28920_, _30091_);
  or g_60605_(_27639_, _28907_, _30093_);
  or g_60606_(_26383_, _30093_, _30094_);
  not g_60607_(_30094_, _30095_);
  or g_60608_(_26380_, _30093_, _30096_);
  and g_60609_(_28906_, _28911_, _30097_);
  and g_60610_(_28899_, _28902_, _30098_);
  and g_60611_(_28860_, _28878_, _30099_);
  and g_60612_(_28871_, _30099_, _30100_);
  and g_60613_(_28882_, _30100_, _30101_);
  and g_60614_(_28868_, _28875_, _30102_);
  and g_60615_(_28864_, _30102_, _30104_);
  and g_60616_(_30101_, _30104_, _30105_);
  and g_60617_(_28887_, _30105_, _30106_);
  not g_60618_(_30106_, _30107_);
  or g_60619_(_28890_, _30105_, _30108_);
  or g_60620_(_28891_, _30107_, _30109_);
  not g_60621_(_30109_, _30110_);
  and g_60622_(_30108_, _30109_, _30111_);
  not g_60623_(_30111_, _30112_);
  and g_60624_(_28895_, _28897_, _30113_);
  or g_60625_(_30110_, _30113_, _30115_);
  xor g_60626_(_30112_, _30113_, _30116_);
  xor g_60627_(_30111_, _30113_, _30117_);
  or g_60628_(_30098_, _30117_, _30118_);
  xor g_60629_(_30098_, _30117_, _30119_);
  xor g_60630_(_30098_, _30116_, _30120_);
  or g_60631_(_30097_, _30120_, _30121_);
  xor g_60632_(_30097_, _30119_, _30122_);
  not g_60633_(_30122_, _30123_);
  or g_60634_(_28915_, _30122_, _30124_);
  xor g_60635_(_28915_, _30123_, _30126_);
  not g_60636_(_30126_, _30127_);
  or g_60637_(_30096_, _30126_, _30128_);
  xor g_60638_(_30096_, _30127_, _30129_);
  or g_60639_(_30094_, _30129_, _30130_);
  and g_60640_(_30094_, _30129_, _30131_);
  xor g_60641_(_30095_, _30129_, _30132_);
  or g_60642_(_27645_, _28917_, _30133_);
  or g_60643_(_28920_, _28921_, _30134_);
  and g_60644_(_30133_, _30134_, _30135_);
  xor g_60645_(_30132_, _30135_, _30137_);
  not g_60646_(_30137_, _30138_);
  or g_60647_(_30091_, _30138_, _30139_);
  and g_60648_(_30091_, _30138_, _30140_);
  xor g_60649_(_30091_, _30137_, _30141_);
  xor g_60650_(_28926_, _30141_, _30142_);
  or g_60651_(_28929_, _30142_, _30143_);
  xor g_60652_(_28929_, _30142_, _30144_);
  xor g_60653_(_28930_, _30142_, _30145_);
  or g_60654_(_28942_, _30145_, _30146_);
  xor g_60655_(_28942_, _30144_, _30148_);
  or g_60656_(_28943_, _30148_, _30149_);
  xor g_60657_(_28944_, _30148_, _30150_);
  or g_60658_(_27664_, _28934_, _30151_);
  or g_60659_(_30150_, _30151_, _30152_);
  xor g_60660_(_30150_, _30151_, _30153_);
  not g_60661_(_30153_, _30154_);
  or g_60662_(_27668_, _28934_, _30155_);
  and g_60663_(_28939_, _30155_, _30156_);
  xor g_60664_(_30153_, _30156_, _30157_);
  or g_60665_(_28946_, _30157_, _30159_);
  and g_60666_(_28946_, _30157_, _30160_);
  xor g_60667_(_28945_, _30157_, _30161_);
  not g_60668_(_30161_, _30162_);
  and g_60669_(_28950_, _28952_, _30163_);
  xor g_60670_(_30162_, _30163_, _30164_);
  xor g_60671_(_30161_, _30163_, _30165_);
  or g_60672_(_28958_, _30164_, _30166_);
  not g_60673_(_30166_, _30167_);
  and g_60674_(_28954_, _30164_, _30168_);
  or g_60675_(_28955_, _30165_, _30170_);
  and g_60676_(_28958_, _30168_, _30171_);
  or g_60677_(_28959_, _30170_, _30172_);
  or g_60678_(_28954_, _30164_, _30173_);
  not g_60679_(_30173_, _30174_);
  and g_60680_(_30172_, _30173_, _30175_);
  or g_60681_(_30171_, _30174_, _30176_);
  and g_60682_(_30166_, _30175_, _30177_);
  or g_60683_(_30167_, _30176_, _30178_);
  xor g_60684_(_28962_, _30177_, _30179_);
  not g_60685_(_30179_, _30181_);
  and g_60686_(_28965_, _28968_, _30182_);
  xor g_60687_(_30181_, _30182_, _30183_);
  or g_60688_(_28975_, _30183_, _30184_);
  xor g_60689_(_28974_, _30183_, _30185_);
  or g_60690_(_28976_, _28978_, _30186_);
  or g_60691_(_30185_, _30186_, _30187_);
  xor g_60692_(_30185_, _30186_, _30188_);
  not g_60693_(_30188_, _30189_);
  or g_60694_(_30090_, _30189_, _30190_);
  xor g_60695_(_30090_, _30188_, _30192_);
  xor g_60696_(_28986_, _30192_, _30193_);
  and g_60697_(_28990_, _30193_, _30194_);
  or g_60698_(_28989_, _30193_, _30195_);
  or g_60699_(_28988_, _30193_, _30196_);
  and g_60700_(_30195_, _30196_, _30197_);
  not g_60701_(_30197_, _30198_);
  or g_60702_(_30194_, _30198_, _30199_);
  not g_60703_(_30199_, _30200_);
  or g_60704_(_28997_, _30199_, _30201_);
  not g_60705_(_30201_, _30203_);
  xor g_60706_(_28997_, _30200_, _30204_);
  not g_60707_(_30204_, _30205_);
  or g_60708_(_30089_, _30204_, _30206_);
  xor g_60709_(_30089_, _30205_, _30207_);
  or g_60710_(_30086_, _30207_, _30208_);
  xor g_60711_(_30086_, _30207_, _30209_);
  xor g_60712_(_30087_, _30207_, _30210_);
  or g_60713_(_29005_, _30209_, _30211_);
  not g_60714_(_30211_, _30212_);
  and g_60715_(_29008_, _30212_, _30214_);
  or g_60716_(_29008_, _30210_, _30215_);
  not g_60717_(_30215_, _30216_);
  and g_60718_(_29005_, _30209_, _30217_);
  not g_60719_(_30217_, _30218_);
  or g_60720_(_30216_, _30217_, _30219_);
  or g_60721_(_30214_, _30219_, _30220_);
  not g_60722_(_30220_, _30221_);
  or g_60723_(_27748_, _29012_, _30222_);
  and g_60724_(_29011_, _30222_, _30223_);
  xor g_60725_(_30221_, _30223_, _30225_);
  or g_60726_(_30085_, _30225_, _30226_);
  xor g_60727_(_30085_, _30225_, _30227_);
  not g_60728_(_30227_, _30228_);
  or g_60729_(_29017_, _30228_, _30229_);
  not g_60730_(_30229_, _30230_);
  xor g_60731_(_29017_, _30227_, _30231_);
  or g_60732_(_29021_, _30231_, _30232_);
  xor g_60733_(_29020_, _30231_, _30233_);
  not g_60734_(_30233_, _30234_);
  or g_60735_(_29023_, _30233_, _30236_);
  xor g_60736_(_29023_, _30234_, _30237_);
  not g_60737_(_30237_, _30238_);
  or g_60738_(_30084_, _30237_, _30239_);
  xor g_60739_(_30084_, _30238_, _30240_);
  or g_60740_(_26512_, _30083_, _30241_);
  not g_60741_(_30241_, _30242_);
  or g_60742_(_30240_, _30241_, _30243_);
  xor g_60743_(_30240_, _30242_, _30244_);
  or g_60744_(_30082_, _30244_, _30245_);
  not g_60745_(_30245_, _30247_);
  and g_60746_(_30082_, _30244_, _30248_);
  xor g_60747_(_30082_, _30244_, _30249_);
  or g_60748_(_30247_, _30248_, _30250_);
  or g_60749_(_30080_, _30250_, _30251_);
  xor g_60750_(_30080_, _30249_, _30252_);
  not g_60751_(_30252_, _30253_);
  xor g_60752_(_30079_, _30253_, _30254_);
  not g_60753_(_30254_, _30255_);
  and g_60754_(_29035_, _29038_, _30256_);
  xor g_60755_(_30255_, _30256_, _30258_);
  xor g_60756_(_30078_, _30258_, _30259_);
  or g_60757_(_29049_, _30259_, _30260_);
  or g_60758_(_29043_, _29044_, _30261_);
  or g_60759_(_30259_, _30261_, _30262_);
  and g_60760_(_29054_, _29057_, _30263_);
  not g_60761_(_30263_, _30264_);
  xor g_60762_(_30259_, _30264_, _30265_);
  or g_60763_(_29058_, _30265_, _30266_);
  xor g_60764_(_29058_, _30265_, _30267_);
  not g_60765_(_30267_, _30269_);
  or g_60766_(_29063_, _30269_, _30270_);
  not g_60767_(_30270_, _30271_);
  xor g_60768_(_29063_, _30267_, _30272_);
  not g_60769_(_30272_, _30273_);
  or g_60770_(_30075_, _30272_, _30274_);
  not g_60771_(_30274_, _30275_);
  xor g_60772_(_30075_, _30273_, _30276_);
  not g_60773_(_30276_, _30277_);
  or g_60774_(_30074_, _30276_, _30278_);
  xor g_60775_(_30074_, _30276_, _30280_);
  xor g_60776_(_30074_, _30277_, _30281_);
  or g_60777_(_30073_, _30281_, _30282_);
  xor g_60778_(_30073_, _30280_, _30283_);
  not g_60779_(_30283_, _30284_);
  or g_60780_(_30072_, _30283_, _30285_);
  xor g_60781_(_30072_, _30283_, _30286_);
  xor g_60782_(_30072_, _30284_, _30287_);
  xor g_60783_(_29072_, _30286_, _30288_);
  not g_60784_(_30288_, _30289_);
  or g_60785_(_30071_, _30288_, _30291_);
  xor g_60786_(_30071_, _30288_, _30292_);
  xor g_60787_(_30071_, _30289_, _30293_);
  and g_60788_(_29082_, _30292_, _30294_);
  or g_60789_(_29080_, _30293_, _30295_);
  or g_60790_(_27831_, _29076_, _30296_);
  or g_60791_(_30293_, _30296_, _30297_);
  xor g_60792_(_30292_, _30296_, _30298_);
  and g_60793_(_29080_, _30298_, _30299_);
  or g_60794_(_30294_, _30299_, _30300_);
  not g_60795_(_30300_, _30302_);
  xor g_60796_(_30068_, _30302_, _30303_);
  or g_60797_(_30066_, _30303_, _30304_);
  xor g_60798_(_30066_, _30303_, _30305_);
  not g_60799_(_30305_, _30306_);
  or g_60800_(_30065_, _30306_, _30307_);
  not g_60801_(_30307_, _30308_);
  xor g_60802_(_30065_, _30305_, _30309_);
  not g_60803_(_30309_, _30310_);
  or g_60804_(_30064_, _30309_, _30311_);
  xor g_60805_(_30064_, _30310_, _30313_);
  or g_60806_(_29091_, _30313_, _30314_);
  not g_60807_(_30314_, _30315_);
  xor g_60808_(_29091_, _30313_, _30316_);
  and g_60809_(_30063_, _30316_, _30317_);
  xor g_60810_(_30062_, _30316_, _30318_);
  not g_60811_(_30318_, _30319_);
  or g_60812_(_30061_, _30318_, _30320_);
  xor g_60813_(_30061_, _30319_, _30321_);
  and g_60814_(_29097_, _29099_, _30322_);
  and g_60815_(_30321_, _30322_, _30324_);
  or g_60816_(_29099_, _30321_, _30325_);
  or g_60817_(_29097_, _30318_, _30326_);
  and g_60818_(_30325_, _30326_, _30327_);
  not g_60819_(_30327_, _30328_);
  or g_60820_(_30324_, _30328_, _30329_);
  not g_60821_(_30329_, _30330_);
  and g_60822_(_29101_, _29104_, _30331_);
  or g_60823_(_30329_, _30331_, _30332_);
  not g_60824_(_30332_, _30333_);
  xor g_60825_(_30330_, _30331_, _30335_);
  not g_60826_(_30335_, _30336_);
  or g_60827_(_30060_, _30335_, _30337_);
  xor g_60828_(_30060_, _30335_, _30338_);
  xor g_60829_(_30060_, _30336_, _30339_);
  or g_60830_(_30058_, _30339_, _30340_);
  xor g_60831_(_30058_, _30338_, _30341_);
  or g_60832_(_29108_, _30341_, _30342_);
  xor g_60833_(_29107_, _30341_, _30343_);
  not g_60834_(_30343_, _30344_);
  or g_60835_(_29112_, _30343_, _30346_);
  not g_60836_(_30346_, _30347_);
  and g_60837_(_29115_, _30344_, _30348_);
  xor g_60838_(_29115_, _30343_, _30349_);
  and g_60839_(_29112_, _30349_, _30350_);
  or g_60840_(_30347_, _30350_, _30351_);
  not g_60841_(_30351_, _30352_);
  xor g_60842_(_30057_, _30352_, _30353_);
  or g_60843_(_29123_, _30353_, _30354_);
  not g_60844_(_30354_, _30355_);
  xor g_60845_(_29124_, _30353_, _30357_);
  and g_60846_(_29130_, _29132_, _30358_);
  not g_60847_(_30358_, _30359_);
  xor g_60848_(_30357_, _30359_, _30360_);
  or g_60849_(_29134_, _30360_, _30361_);
  xor g_60850_(_29134_, _30360_, _30362_);
  not g_60851_(_30362_, _30363_);
  or g_60852_(_29137_, _30363_, _30364_);
  not g_60853_(_30364_, _30365_);
  xor g_60854_(_29137_, _30362_, _30366_);
  not g_60855_(_30366_, _30368_);
  or g_60856_(_30056_, _30366_, _30369_);
  xor g_60857_(_30056_, _30366_, _30370_);
  xor g_60858_(_30056_, _30368_, _30371_);
  or g_60859_(_29138_, _29140_, _30372_);
  and g_60860_(_29143_, _30372_, _30373_);
  xor g_60861_(_30371_, _30373_, _30374_);
  not g_60862_(_30374_, _30375_);
  and g_60863_(_30055_, _30374_, _30376_);
  xor g_60864_(_30055_, _30374_, _30377_);
  xor g_60865_(_30055_, _30375_, _30379_);
  or g_60866_(_30054_, _30379_, _30380_);
  not g_60867_(_30380_, _30381_);
  xor g_60868_(_30054_, _30377_, _30382_);
  or g_60869_(_30052_, _30382_, _30383_);
  not g_60870_(_30383_, _30384_);
  xor g_60871_(_30053_, _30382_, _30385_);
  or g_60872_(_29162_, _30385_, _30386_);
  not g_60873_(_30386_, _30387_);
  or g_60874_(_29159_, _30385_, _30388_);
  xor g_60875_(_29157_, _30385_, _30390_);
  not g_60876_(_30390_, _30391_);
  or g_60877_(_29164_, _30390_, _30392_);
  xor g_60878_(_29164_, _30391_, _30393_);
  and g_60879_(_29162_, _30393_, _30394_);
  or g_60880_(_30387_, _30394_, _30395_);
  or g_60881_(_26692_, _30049_, _30396_);
  and g_60882_(_29166_, _30396_, _30397_);
  xor g_60883_(_30395_, _30397_, _30398_);
  and g_60884_(_30051_, _30398_, _30399_);
  not g_60885_(_30399_, _30401_);
  xor g_60886_(_30050_, _30398_, _30402_);
  not g_60887_(_30402_, _30403_);
  xor g_60888_(_29173_, _30403_, _30404_);
  xor g_60889_(_29173_, _30402_, _30405_);
  or g_60890_(_29178_, _30404_, _30406_);
  xor g_60891_(_29178_, _30405_, _30407_);
  not g_60892_(_30407_, _30408_);
  and g_60893_(_29182_, _29184_, _30409_);
  xor g_60894_(_30407_, _30409_, _30410_);
  xor g_60895_(_30408_, _30409_, _30412_);
  or g_60896_(_29187_, _30412_, _30413_);
  xor g_60897_(_29187_, _30412_, _30414_);
  xor g_60898_(_29187_, _30410_, _30415_);
  or g_60899_(_29193_, _30415_, _30416_);
  not g_60900_(_30416_, _30417_);
  or g_60901_(_27959_, _29188_, _30418_);
  or g_60902_(_27958_, _29188_, _30419_);
  not g_60903_(_30419_, _30420_);
  and g_60904_(_30414_, _30420_, _30421_);
  or g_60905_(_30415_, _30419_, _30423_);
  xor g_60906_(_30415_, _30419_, _30424_);
  xor g_60907_(_30415_, _30420_, _30425_);
  or g_60908_(_30418_, _30425_, _30426_);
  xor g_60909_(_30418_, _30424_, _30427_);
  and g_60910_(_29193_, _30427_, _30428_);
  or g_60911_(_30417_, _30428_, _30429_);
  or g_60912_(_29197_, _30429_, _30430_);
  xor g_60913_(_29198_, _30429_, _30431_);
  or g_60914_(_29201_, _30431_, _30432_);
  xor g_60915_(_29203_, _30431_, _30434_);
  or g_60916_(_29206_, _30434_, _30435_);
  xor g_60917_(_29207_, _30434_, _30436_);
  or g_60918_(_29211_, _30436_, _30437_);
  xor g_60919_(_29211_, _30436_, _30438_);
  not g_60920_(_30438_, _30439_);
  or g_60921_(_30047_, _30439_, _30440_);
  xor g_60922_(_30047_, _30438_, _30441_);
  or g_60923_(_30045_, _30441_, _30442_);
  xor g_60924_(_30046_, _30441_, _30443_);
  or g_60925_(_29217_, _30443_, _30445_);
  xor g_60926_(_29218_, _30443_, _30446_);
  or g_60927_(_29221_, _30446_, _30447_);
  xor g_60928_(_29222_, _30446_, _30448_);
  or g_60929_(_29225_, _30448_, _30449_);
  xor g_60930_(_29225_, _30448_, _30450_);
  xor g_60931_(_29226_, _30448_, _30451_);
  and g_60932_(_29228_, _30451_, _30452_);
  or g_60933_(_29229_, _30450_, _30453_);
  and g_60934_(_30043_, _30452_, _30454_);
  or g_60935_(_30044_, _30453_, _30456_);
  or g_60936_(_29228_, _30451_, _30457_);
  not g_60937_(_30457_, _30458_);
  or g_60938_(_30043_, _30451_, _30459_);
  not g_60939_(_30459_, _30460_);
  and g_60940_(_30457_, _30459_, _30461_);
  not g_60941_(_30461_, _30462_);
  and g_60942_(_30456_, _30461_, _30463_);
  or g_60943_(_30454_, _30462_, _30464_);
  or g_60944_(_30042_, _30464_, _30465_);
  xor g_60945_(_30042_, _30463_, _30467_);
  not g_60946_(_30467_, _30468_);
  or g_60947_(_27995_, _29237_, _30469_);
  and g_60948_(_29236_, _30469_, _30470_);
  xor g_60949_(_30468_, _30470_, _30471_);
  xor g_60950_(_30467_, _30470_, _30472_);
  or g_60951_(_30041_, _30471_, _30473_);
  xor g_60952_(_30041_, _30472_, _30474_);
  not g_60953_(_30474_, _30475_);
  and g_60954_(_29241_, _29244_, _30476_);
  xor g_60955_(_30475_, _30476_, _30478_);
  xor g_60956_(_30474_, _30476_, _30479_);
  and g_60957_(_29248_, _30479_, _30480_);
  or g_60958_(_29247_, _30478_, _30481_);
  xor g_60959_(_29247_, _30478_, _30482_);
  xor g_60960_(_29248_, _30478_, _30483_);
  and g_60961_(_29251_, _30482_, _30484_);
  or g_60962_(_29250_, _30483_, _30485_);
  xor g_60963_(_29250_, _30482_, _30486_);
  or g_60964_(_29255_, _30486_, _30487_);
  xor g_60965_(_29254_, _30486_, _30489_);
  not g_60966_(_30489_, _30490_);
  or g_60967_(_29259_, _30489_, _30491_);
  xor g_60968_(_29259_, _30489_, _30492_);
  xor g_60969_(_29259_, _30490_, _30493_);
  or g_60970_(_29261_, _30493_, _30494_);
  xor g_60971_(_29261_, _30492_, _30495_);
  or g_60972_(_30039_, _30495_, _30496_);
  not g_60973_(_30496_, _30497_);
  xor g_60974_(_30039_, _30495_, _30498_);
  xor g_60975_(_30040_, _30495_, _30500_);
  or g_60976_(_30038_, _30500_, _30501_);
  not g_60977_(_30501_, _30502_);
  xor g_60978_(_30038_, _30498_, _30503_);
  and g_60979_(_29266_, _29269_, _30504_);
  xor g_60980_(_30503_, _30504_, _30505_);
  not g_60981_(_30505_, _30506_);
  or g_60982_(_30035_, _30506_, _30507_);
  xor g_60983_(_30036_, _30505_, _30508_);
  xor g_60984_(_30035_, _30505_, _30509_);
  or g_60985_(_30033_, _30509_, _30511_);
  xor g_60986_(_30033_, _30508_, _30512_);
  or g_60987_(_28038_, _29270_, _30513_);
  not g_60988_(_30513_, _30514_);
  or g_60989_(_30512_, _30513_, _30515_);
  not g_60990_(_30515_, _30516_);
  xor g_60991_(_30512_, _30513_, _30517_);
  xor g_60992_(_30512_, _30514_, _30518_);
  and g_60993_(_30032_, _30518_, _30519_);
  and g_60994_(_28046_, _29272_, _30520_);
  or g_60995_(_28045_, _29273_, _30522_);
  and g_60996_(_30517_, _30520_, _30523_);
  or g_60997_(_30518_, _30522_, _30524_);
  or g_60998_(_30519_, _30523_, _30525_);
  not g_60999_(_30525_, _30526_);
  or g_61000_(_30031_, _30525_, _30527_);
  not g_61001_(_30527_, _30528_);
  xor g_61002_(_30031_, _30526_, _30529_);
  not g_61003_(_30529_, _30530_);
  or g_61004_(_26823_, _30030_, _30531_);
  not g_61005_(_30531_, _30533_);
  or g_61006_(_29276_, _30533_, _30534_);
  xor g_61007_(_30529_, _30534_, _30535_);
  not g_61008_(_30535_, _30536_);
  or g_61009_(_28060_, _29281_, _30537_);
  and g_61010_(_29280_, _30537_, _30538_);
  or g_61011_(_30535_, _30538_, _30539_);
  not g_61012_(_30539_, _30540_);
  xor g_61013_(_30536_, _30538_, _30541_);
  or g_61014_(_30029_, _30541_, _30542_);
  not g_61015_(_30542_, _30544_);
  and g_61016_(_30029_, _30541_, _30545_);
  xor g_61017_(_30029_, _30541_, _30546_);
  or g_61018_(_30544_, _30545_, _30547_);
  or g_61019_(_28067_, _29287_, _30548_);
  and g_61020_(_29286_, _30548_, _30549_);
  xor g_61021_(_30546_, _30549_, _30550_);
  or g_61022_(_30028_, _30550_, _30551_);
  not g_61023_(_30551_, _30552_);
  xor g_61024_(_30028_, _30550_, _30553_);
  not g_61025_(_30553_, _30555_);
  and g_61026_(_29293_, _30553_, _30556_);
  or g_61027_(_29292_, _30555_, _30557_);
  xor g_61028_(_29292_, _30553_, _30558_);
  or g_61029_(_29299_, _30558_, _30559_);
  not g_61030_(_30559_, _30560_);
  and g_61031_(_29297_, _30558_, _30561_);
  and g_61032_(_29299_, _30561_, _30562_);
  or g_61033_(_29297_, _30558_, _30563_);
  not g_61034_(_30563_, _30564_);
  or g_61035_(_30562_, _30564_, _30566_);
  or g_61036_(_30560_, _30566_, _30567_);
  not g_61037_(_30567_, _30568_);
  or g_61038_(_29303_, _30567_, _30569_);
  not g_61039_(_30569_, _30570_);
  xor g_61040_(_29303_, _30568_, _30571_);
  or g_61041_(_29307_, _30571_, _30572_);
  xor g_61042_(_29306_, _30571_, _30573_);
  and g_61043_(_29309_, _29313_, _30574_);
  not g_61044_(_30574_, _30575_);
  xor g_61045_(_30573_, _30575_, _30577_);
  not g_61046_(_30577_, _30578_);
  and g_61047_(_29316_, _29318_, _30579_);
  not g_61048_(_30579_, _30580_);
  xor g_61049_(_30577_, _30580_, _30581_);
  or g_61050_(_29324_, _30581_, _30582_);
  not g_61051_(_30582_, _30583_);
  and g_61052_(_29324_, _30581_, _30584_);
  xor g_61053_(_29324_, _30581_, _30585_);
  or g_61054_(_30583_, _30584_, _30586_);
  and g_61055_(_29328_, _29331_, _30588_);
  xor g_61056_(_30585_, _30588_, _30589_);
  not g_61057_(_30589_, _30590_);
  or g_61058_(_29336_, _30589_, _30591_);
  xor g_61059_(_29336_, _30589_, _30592_);
  xor g_61060_(_29336_, _30590_, _30593_);
  and g_61061_(_29340_, _29342_, _30594_);
  xor g_61062_(_30592_, _30594_, _30595_);
  or g_61063_(_30025_, _30595_, _30596_);
  xor g_61064_(_30027_, _30595_, _30597_);
  or g_61065_(_30023_, _30597_, _30599_);
  xor g_61066_(_30024_, _30597_, _30600_);
  not g_61067_(_30600_, _30601_);
  and g_61068_(_29349_, _29353_, _30602_);
  and g_61069_(_30600_, _30602_, _30603_);
  and g_61070_(_29352_, _30601_, _30604_);
  not g_61071_(_30604_, _30605_);
  or g_61072_(_29349_, _30600_, _30606_);
  not g_61073_(_30606_, _30607_);
  or g_61074_(_30604_, _30607_, _30608_);
  or g_61075_(_30603_, _30608_, _30610_);
  or g_61076_(_29355_, _30610_, _30611_);
  xor g_61077_(_29355_, _30610_, _30612_);
  not g_61078_(_30612_, _30613_);
  and g_61079_(_29360_, _30612_, _30614_);
  or g_61080_(_29359_, _30613_, _30615_);
  and g_61081_(_29364_, _30612_, _30616_);
  or g_61082_(_29363_, _30613_, _30617_);
  xor g_61083_(_29363_, _30612_, _30618_);
  and g_61084_(_29359_, _30618_, _30619_);
  or g_61085_(_30614_, _30619_, _30621_);
  not g_61086_(_30621_, _30622_);
  and g_61087_(_29365_, _30622_, _30623_);
  or g_61088_(_29366_, _30621_, _30624_);
  xor g_61089_(_29365_, _30621_, _30625_);
  or g_61090_(_29371_, _30625_, _30626_);
  xor g_61091_(_29371_, _30625_, _30627_);
  xor g_61092_(_29372_, _30625_, _30628_);
  and g_61093_(_29380_, _30627_, _30629_);
  or g_61094_(_29379_, _30628_, _30630_);
  and g_61095_(_29376_, _30627_, _30632_);
  or g_61096_(_29375_, _30628_, _30633_);
  or g_61097_(_30629_, _30632_, _30634_);
  and g_61098_(_29375_, _30628_, _30635_);
  and g_61099_(_29379_, _30635_, _30636_);
  or g_61100_(_30634_, _30636_, _30637_);
  or g_61101_(_29382_, _30637_, _30638_);
  xor g_61102_(_29383_, _30637_, _30639_);
  or g_61103_(_30021_, _30639_, _30640_);
  xor g_61104_(_30022_, _30639_, _30641_);
  or g_61105_(_26933_, _30020_, _30643_);
  or g_61106_(_28166_, _29384_, _30644_);
  and g_61107_(_30643_, _30644_, _30645_);
  xor g_61108_(_30641_, _30645_, _30646_);
  not g_61109_(_30646_, _30647_);
  and g_61110_(_29388_, _30646_, _30648_);
  or g_61111_(_29390_, _30647_, _30649_);
  xor g_61112_(_29388_, _30646_, _30650_);
  xor g_61113_(_29390_, _30646_, _30651_);
  and g_61114_(_29392_, _29397_, _30652_);
  xor g_61115_(_30651_, _30652_, _30654_);
  not g_61116_(_30654_, _30655_);
  and g_61117_(_29404_, _30654_, _30656_);
  or g_61118_(_29403_, _30655_, _30657_);
  xor g_61119_(_29403_, _30654_, _30658_);
  not g_61120_(_30658_, _30659_);
  or g_61121_(_28184_, _29407_, _30660_);
  and g_61122_(_29406_, _30660_, _30661_);
  xor g_61123_(_30659_, _30661_, _30662_);
  or g_61124_(_30019_, _30662_, _30663_);
  not g_61125_(_30663_, _30665_);
  xor g_61126_(_30019_, _30662_, _30666_);
  not g_61127_(_30666_, _30667_);
  and g_61128_(_29409_, _29414_, _30668_);
  xor g_61129_(_30666_, _30668_, _30669_);
  not g_61130_(_30669_, _30670_);
  and g_61131_(_29417_, _29420_, _30671_);
  xor g_61132_(_30670_, _30671_, _30672_);
  not g_61133_(_30672_, _30673_);
  xor g_61134_(_30018_, _30673_, _30674_);
  not g_61135_(_30674_, _30676_);
  or g_61136_(_28209_, _29426_, _30677_);
  or g_61137_(_28199_, _29424_, _30678_);
  or g_61138_(_26973_, _30678_, _30679_);
  and g_61139_(_30677_, _30679_, _30680_);
  xor g_61140_(_30676_, _30680_, _30681_);
  xor g_61141_(_30674_, _30680_, _30682_);
  or g_61142_(_30014_, _30681_, _30683_);
  not g_61143_(_30683_, _30684_);
  and g_61144_(_29431_, _30681_, _30685_);
  or g_61145_(_29432_, _30682_, _30687_);
  and g_61146_(_30014_, _30685_, _30688_);
  or g_61147_(_30016_, _30687_, _30689_);
  or g_61148_(_29431_, _30681_, _30690_);
  not g_61149_(_30690_, _30691_);
  and g_61150_(_30689_, _30690_, _30692_);
  or g_61151_(_30688_, _30691_, _30693_);
  and g_61152_(_30683_, _30692_, _30694_);
  or g_61153_(_30684_, _30693_, _30695_);
  or g_61154_(_30013_, _30695_, _30696_);
  not g_61155_(_30696_, _30698_);
  xor g_61156_(_30013_, _30694_, _30699_);
  not g_61157_(_30699_, _30700_);
  or g_61158_(_29439_, _30699_, _30701_);
  xor g_61159_(_29439_, _30699_, _30702_);
  xor g_61160_(_29439_, _30700_, _30703_);
  and g_61161_(_29442_, _30702_, _30704_);
  or g_61162_(_29443_, _30703_, _30705_);
  xor g_61163_(_29443_, _30702_, _30706_);
  not g_61164_(_30706_, _30707_);
  and g_61165_(_29447_, _30707_, _30709_);
  or g_61166_(_29448_, _30706_, _30710_);
  xor g_61167_(_29447_, _30706_, _30711_);
  and g_61168_(_29451_, _29454_, _30712_);
  xor g_61169_(_30711_, _30712_, _30713_);
  not g_61170_(_30713_, _30714_);
  and g_61171_(_29458_, _29462_, _30715_);
  xor g_61172_(_30713_, _30715_, _30716_);
  or g_61173_(_30012_, _30716_, _30717_);
  not g_61174_(_30717_, _30718_);
  xor g_61175_(_30012_, _30716_, _30720_);
  not g_61176_(_30720_, _30721_);
  or g_61177_(_30011_, _30721_, _30722_);
  xor g_61178_(_30011_, _30720_, _30723_);
  not g_61179_(_30723_, _30724_);
  or g_61180_(_30010_, _30723_, _30725_);
  xor g_61181_(_30010_, _30724_, _30726_);
  or g_61182_(_28243_, _29468_, _30727_);
  or g_61183_(_28247_, _29468_, _30728_);
  and g_61184_(_30727_, _30728_, _30729_);
  xor g_61185_(_30726_, _30729_, _30731_);
  and g_61186_(_29471_, _30731_, _30732_);
  not g_61187_(_30732_, _30733_);
  xor g_61188_(_29470_, _30731_, _30734_);
  not g_61189_(_30734_, _30735_);
  and g_61190_(_29474_, _29478_, _30736_);
  xor g_61191_(_30735_, _30736_, _30737_);
  not g_61192_(_30737_, _30738_);
  xor g_61193_(_30009_, _30738_, _30739_);
  or g_61194_(_29486_, _30739_, _30740_);
  xor g_61195_(_29485_, _30739_, _30742_);
  not g_61196_(_30742_, _30743_);
  or g_61197_(_30008_, _30742_, _30744_);
  xor g_61198_(_30008_, _30742_, _30745_);
  xor g_61199_(_30008_, _30743_, _30746_);
  or g_61200_(_30007_, _30746_, _30747_);
  xor g_61201_(_30007_, _30745_, _30748_);
  or g_61202_(_28284_, _29495_, _30749_);
  and g_61203_(_29493_, _30749_, _30750_);
  xor g_61204_(_30748_, _30750_, _30751_);
  not g_61205_(_30751_, _30753_);
  or g_61206_(_28287_, _29495_, _30754_);
  not g_61207_(_30754_, _30755_);
  and g_61208_(_29498_, _30754_, _30756_);
  xor g_61209_(_30751_, _30756_, _30757_);
  xor g_61210_(_30006_, _30757_, _30758_);
  not g_61211_(_30758_, _30759_);
  xor g_61212_(_30005_, _30758_, _30760_);
  or g_61213_(_30001_, _30760_, _30761_);
  not g_61214_(_30761_, _30762_);
  xor g_61215_(_30001_, _30760_, _30764_);
  and g_61216_(_29999_, _30764_, _30765_);
  not g_61217_(_30765_, _30766_);
  xor g_61218_(_29999_, _30764_, _30767_);
  xor g_61219_(_29998_, _30764_, _30768_);
  xor g_61220_(_29514_, _30767_, _30769_);
  or g_61221_(_29517_, _30769_, _30770_);
  not g_61222_(_30770_, _30771_);
  xor g_61223_(_29518_, _30769_, _30772_);
  or g_61224_(_29524_, _30772_, _30773_);
  or g_61225_(_29520_, _30772_, _30775_);
  and g_61226_(_30773_, _30775_, _30776_);
  not g_61227_(_30776_, _30777_);
  and g_61228_(_29520_, _30772_, _30778_);
  and g_61229_(_29524_, _30778_, _30779_);
  not g_61230_(_30779_, _30780_);
  and g_61231_(_30776_, _30780_, _30781_);
  or g_61232_(_30777_, _30779_, _30782_);
  and g_61233_(_29996_, _30782_, _30783_);
  or g_61234_(_29997_, _30781_, _30784_);
  or g_61235_(_28333_, _29519_, _30786_);
  or g_61236_(_30782_, _30786_, _30787_);
  not g_61237_(_30787_, _30788_);
  and g_61238_(_30784_, _30787_, _30789_);
  or g_61239_(_30783_, _30788_, _30790_);
  or g_61240_(_28339_, _29525_, _30791_);
  or g_61241_(_30790_, _30791_, _30792_);
  xor g_61242_(_30789_, _30791_, _30793_);
  not g_61243_(_30793_, _30794_);
  or g_61244_(_29995_, _30793_, _30795_);
  xor g_61245_(_29995_, _30794_, _30797_);
  or g_61246_(_28344_, _29527_, _30798_);
  and g_61247_(_29530_, _30798_, _30799_);
  xor g_61248_(_30797_, _30799_, _30800_);
  not g_61249_(_30800_, _30801_);
  or g_61250_(_29534_, _30801_, _30802_);
  xor g_61251_(_29534_, _30800_, _30803_);
  not g_61252_(_30803_, _30804_);
  or g_61253_(_29994_, _30803_, _30805_);
  xor g_61254_(_29994_, _30803_, _30806_);
  xor g_61255_(_29994_, _30804_, _30808_);
  or g_61256_(_29992_, _30808_, _30809_);
  xor g_61257_(_29992_, _30806_, _30810_);
  or g_61258_(_29538_, _30810_, _30811_);
  not g_61259_(_30811_, _30812_);
  xor g_61260_(_29538_, _30810_, _30813_);
  xor g_61261_(_29539_, _30810_, _30814_);
  and g_61262_(_29544_, _30814_, _30815_);
  and g_61263_(_29536_, _29542_, _30816_);
  or g_61264_(_29537_, _29541_, _30817_);
  and g_61265_(_30813_, _30816_, _30819_);
  or g_61266_(_30814_, _30817_, _30820_);
  or g_61267_(_30815_, _30819_, _30821_);
  or g_61268_(_29546_, _30821_, _30822_);
  xor g_61269_(_29547_, _30821_, _30823_);
  or g_61270_(_29553_, _30823_, _30824_);
  xor g_61271_(_29552_, _30823_, _30825_);
  or g_61272_(_29551_, _30825_, _30826_);
  not g_61273_(_30826_, _30827_);
  xor g_61274_(_29550_, _30825_, _30828_);
  or g_61275_(_29989_, _30828_, _30830_);
  not g_61276_(_30830_, _30831_);
  xor g_61277_(_29990_, _30828_, _30832_);
  or g_61278_(_28369_, _29557_, _30833_);
  or g_61279_(_27144_, _29987_, _30834_);
  and g_61280_(_30833_, _30834_, _30835_);
  xor g_61281_(_30832_, _30835_, _30836_);
  not g_61282_(_30836_, _30837_);
  or g_61283_(_29988_, _30837_, _30838_);
  xor g_61284_(_29988_, _30836_, _30839_);
  or g_61285_(_29568_, _30839_, _30841_);
  xor g_61286_(_29569_, _30839_, _30842_);
  not g_61287_(_30842_, _30843_);
  or g_61288_(_29567_, _30842_, _30844_);
  xor g_61289_(_29567_, _30842_, _30845_);
  xor g_61290_(_29567_, _30843_, _30846_);
  or g_61291_(_29574_, _30846_, _30847_);
  xor g_61292_(_29574_, _30845_, _30848_);
  not g_61293_(_30848_, _30849_);
  or g_61294_(_29577_, _30848_, _30850_);
  xor g_61295_(_29577_, _30848_, _30852_);
  xor g_61296_(_29577_, _30849_, _30853_);
  and g_61297_(_29579_, _29583_, _30854_);
  xor g_61298_(_30852_, _30854_, _30855_);
  xor g_61299_(_30853_, _30854_, _30856_);
  and g_61300_(_29986_, _30856_, _30857_);
  not g_61301_(_30857_, _30858_);
  xor g_61302_(_29985_, _30855_, _30859_);
  xor g_61303_(_29986_, _30855_, _30860_);
  and g_61304_(_29984_, _30859_, _30861_);
  or g_61305_(_29983_, _30860_, _30863_);
  xor g_61306_(_29983_, _30859_, _30864_);
  or g_61307_(_29981_, _30864_, _30865_);
  xor g_61308_(_29981_, _30864_, _30866_);
  xor g_61309_(_29980_, _30864_, _30867_);
  and g_61310_(_29588_, _29593_, _30868_);
  or g_61311_(_29589_, _29592_, _30869_);
  and g_61312_(_29599_, _30869_, _30870_);
  or g_61313_(_29597_, _30868_, _30871_);
  and g_61314_(_30867_, _30870_, _30872_);
  or g_61315_(_30866_, _30871_, _30874_);
  and g_61316_(_29597_, _30866_, _30875_);
  or g_61317_(_29599_, _30867_, _30876_);
  and g_61318_(_30866_, _30868_, _30877_);
  or g_61319_(_30867_, _30869_, _30878_);
  and g_61320_(_30876_, _30878_, _30879_);
  or g_61321_(_30875_, _30877_, _30880_);
  and g_61322_(_30874_, _30879_, _30881_);
  or g_61323_(_30872_, _30880_, _30882_);
  or g_61324_(_28409_, _29605_, _30883_);
  and g_61325_(_29603_, _30883_, _30885_);
  xor g_61326_(_30881_, _30885_, _30886_);
  or g_61327_(_29979_, _30886_, _30887_);
  xor g_61328_(_29978_, _30886_, _30888_);
  not g_61329_(_30888_, _30889_);
  and g_61330_(_29608_, _29612_, _30890_);
  xor g_61331_(_30889_, _30890_, _30891_);
  or g_61332_(_29977_, _30891_, _30892_);
  xor g_61333_(_29977_, _30891_, _30893_);
  not g_61334_(_30893_, _30894_);
  and g_61335_(_29976_, _30893_, _30896_);
  or g_61336_(_29975_, _30894_, _30897_);
  xor g_61337_(_29976_, _30893_, _30898_);
  xor g_61338_(_29975_, _30893_, _30899_);
  or g_61339_(_29616_, _30899_, _30900_);
  xor g_61340_(_29616_, _30898_, _30901_);
  not g_61341_(_30901_, _30902_);
  or g_61342_(_29619_, _30901_, _30903_);
  not g_61343_(_30903_, _30904_);
  xor g_61344_(_29619_, _30901_, _30905_);
  xor g_61345_(_29619_, _30902_, _30907_);
  or g_61346_(_29623_, _30907_, _30908_);
  not g_61347_(_30908_, _30909_);
  xor g_61348_(_29623_, _30905_, _30910_);
  not g_61349_(_30910_, _30911_);
  or g_61350_(_29626_, _30910_, _30912_);
  xor g_61351_(_29626_, _30911_, _30913_);
  not g_61352_(_30913_, _30914_);
  or g_61353_(_29629_, _30913_, _30915_);
  xor g_61354_(_29629_, _30914_, _30916_);
  not g_61355_(_30916_, _30918_);
  or g_61356_(_28446_, _29634_, _30919_);
  and g_61357_(_29633_, _30919_, _30920_);
  xor g_61358_(_30916_, _30920_, _30921_);
  xor g_61359_(_30918_, _30920_, _30922_);
  or g_61360_(_28450_, _29634_, _30923_);
  not g_61361_(_30923_, _30924_);
  and g_61362_(_29638_, _30923_, _30925_);
  xor g_61363_(_30921_, _30925_, _30926_);
  xor g_61364_(_29973_, _30926_, _30927_);
  xor g_61365_(_29974_, _30926_, _30929_);
  or g_61366_(_29972_, _30929_, _30930_);
  xor g_61367_(_29972_, _30927_, _30931_);
  not g_61368_(_30931_, _30932_);
  or g_61369_(_29970_, _30931_, _30933_);
  xor g_61370_(_29970_, _30932_, _30934_);
  not g_61371_(_30934_, _30935_);
  and g_61372_(_29651_, _29654_, _30936_);
  xor g_61373_(_30935_, _30936_, _30937_);
  not g_61374_(_30937_, _30938_);
  and g_61375_(_29656_, _29659_, _30940_);
  xor g_61376_(_30938_, _30940_, _30941_);
  not g_61377_(_30941_, _30942_);
  and g_61378_(_29662_, _29665_, _30943_);
  xor g_61379_(_30941_, _30943_, _30944_);
  xor g_61380_(_30942_, _30943_, _30945_);
  or g_61381_(_29671_, _30945_, _30946_);
  not g_61382_(_30946_, _30947_);
  or g_61383_(_29667_, _30945_, _30948_);
  xor g_61384_(_29667_, _30944_, _30949_);
  and g_61385_(_29671_, _30949_, _30951_);
  or g_61386_(_30947_, _30951_, _30952_);
  and g_61387_(_29676_, _29679_, _30953_);
  xor g_61388_(_30952_, _30953_, _30954_);
  and g_61389_(_29969_, _30954_, _30955_);
  not g_61390_(_30955_, _30956_);
  xor g_61391_(_29968_, _30954_, _30957_);
  or g_61392_(_29966_, _30957_, _30958_);
  not g_61393_(_30958_, _30959_);
  xor g_61394_(_29967_, _30957_, _30960_);
  not g_61395_(_30960_, _30962_);
  and g_61396_(_29687_, _29694_, _30963_);
  or g_61397_(_29688_, _29693_, _30964_);
  and g_61398_(_30960_, _30963_, _30965_);
  or g_61399_(_30962_, _30964_, _30966_);
  or g_61400_(_29694_, _30960_, _30967_);
  not g_61401_(_30967_, _30968_);
  or g_61402_(_29687_, _30960_, _30969_);
  not g_61403_(_30969_, _30970_);
  and g_61404_(_30967_, _30969_, _30971_);
  not g_61405_(_30971_, _30973_);
  and g_61406_(_30966_, _30971_, _30974_);
  or g_61407_(_30965_, _30973_, _30975_);
  xor g_61408_(_29965_, _30974_, _30976_);
  or g_61409_(_29962_, _30976_, _30977_);
  xor g_61410_(_29963_, _30976_, _30978_);
  or g_61411_(_29704_, _30978_, _30979_);
  not g_61412_(_30979_, _30980_);
  and g_61413_(_29702_, _30978_, _30981_);
  and g_61414_(_29704_, _30981_, _30982_);
  or g_61415_(_29702_, _30978_, _30984_);
  not g_61416_(_30984_, _30985_);
  or g_61417_(_30982_, _30985_, _30986_);
  or g_61418_(_30980_, _30986_, _30987_);
  or g_61419_(_29707_, _30987_, _30988_);
  xor g_61420_(_29709_, _30987_, _30989_);
  not g_61421_(_30989_, _30990_);
  and g_61422_(_29710_, _29717_, _30991_);
  xor g_61423_(_30989_, _30991_, _30992_);
  xor g_61424_(_30990_, _30991_, _30993_);
  xor g_61425_(_29961_, _30992_, _30995_);
  or g_61426_(_29728_, _30995_, _30996_);
  xor g_61427_(_29728_, _30995_, _30997_);
  xor g_61428_(_29729_, _30995_, _30998_);
  and g_61429_(_29734_, _30997_, _30999_);
  or g_61430_(_29733_, _30998_, _31000_);
  xor g_61431_(_29734_, _30997_, _31001_);
  xor g_61432_(_29738_, _31001_, _31002_);
  not g_61433_(_31002_, _31003_);
  xor g_61434_(_29959_, _31003_, _31004_);
  not g_61435_(_31004_, _31006_);
  and g_61436_(_29750_, _31006_, _31007_);
  or g_61437_(_29744_, _31004_, _31008_);
  not g_61438_(_31008_, _31009_);
  xor g_61439_(_29744_, _31004_, _31010_);
  xor g_61440_(_29744_, _31006_, _31011_);
  or g_61441_(_29750_, _31010_, _31012_);
  not g_61442_(_31012_, _31013_);
  or g_61443_(_31007_, _31013_, _31014_);
  and g_61444_(_29755_, _29758_, _31015_);
  xor g_61445_(_31014_, _31015_, _31017_);
  not g_61446_(_31017_, _31018_);
  or g_61447_(_29761_, _31018_, _31019_);
  xor g_61448_(_29761_, _31017_, _31020_);
  or g_61449_(_28561_, _29759_, _31021_);
  not g_61450_(_31021_, _31022_);
  or g_61451_(_31020_, _31021_, _31023_);
  not g_61452_(_31023_, _31024_);
  xor g_61453_(_31020_, _31021_, _31025_);
  xor g_61454_(_31020_, _31022_, _31026_);
  or g_61455_(_29958_, _31026_, _31028_);
  xor g_61456_(_29958_, _31025_, _31029_);
  or g_61457_(_29769_, _31029_, _31030_);
  not g_61458_(_31030_, _31031_);
  xor g_61459_(_29769_, _31029_, _31032_);
  xor g_61460_(_29768_, _31029_, _31033_);
  and g_61461_(_29772_, _29776_, _31034_);
  xor g_61462_(_31032_, _31034_, _31035_);
  or g_61463_(_29782_, _31035_, _31036_);
  not g_61464_(_31036_, _31037_);
  and g_61465_(_29779_, _31035_, _31039_);
  and g_61466_(_29782_, _31039_, _31040_);
  or g_61467_(_29779_, _31035_, _31041_);
  not g_61468_(_31041_, _31042_);
  or g_61469_(_31040_, _31042_, _31043_);
  or g_61470_(_31037_, _31043_, _31044_);
  not g_61471_(_31044_, _31045_);
  or g_61472_(_29786_, _31044_, _31046_);
  xor g_61473_(_29786_, _31044_, _31047_);
  xor g_61474_(_29786_, _31045_, _31048_);
  and g_61475_(_29789_, _29795_, _31050_);
  and g_61476_(_31048_, _31050_, _31051_);
  and g_61477_(_29797_, _31047_, _31052_);
  or g_61478_(_29795_, _31048_, _31053_);
  and g_61479_(_29790_, _31047_, _31054_);
  or g_61480_(_29789_, _31048_, _31055_);
  or g_61481_(_31052_, _31054_, _31056_);
  or g_61482_(_31051_, _31056_, _31057_);
  or g_61483_(_29794_, _31057_, _31058_);
  xor g_61484_(_29794_, _31057_, _31059_);
  not g_61485_(_31059_, _31061_);
  or g_61486_(_29801_, _31061_, _31062_);
  not g_61487_(_31062_, _31063_);
  xor g_61488_(_29801_, _31059_, _31064_);
  not g_61489_(_31064_, _31065_);
  and g_61490_(_29957_, _31065_, _31066_);
  not g_61491_(_31066_, _31067_);
  and g_61492_(_28595_, _29802_, _31068_);
  or g_61493_(_28594_, _29803_, _31069_);
  and g_61494_(_31064_, _31069_, _31070_);
  and g_61495_(_29956_, _31070_, _31072_);
  and g_61496_(_31059_, _31068_, _31073_);
  not g_61497_(_31073_, _31074_);
  or g_61498_(_31072_, _31073_, _31075_);
  or g_61499_(_31066_, _31075_, _31076_);
  not g_61500_(_31076_, _31077_);
  and g_61501_(_29808_, _29811_, _31078_);
  xor g_61502_(_31077_, _31078_, _31079_);
  xor g_61503_(_31076_, _31078_, _31080_);
  and g_61504_(_29814_, _31079_, _31081_);
  or g_61505_(_28749_, _29809_, _31083_);
  not g_61506_(_31083_, _31084_);
  and g_61507_(_31080_, _31084_, _31085_);
  or g_61508_(_31079_, _31083_, _31086_);
  or g_61509_(_31081_, _31085_, _31087_);
  not g_61510_(_31087_, _31088_);
  or g_61511_(_29817_, _31087_, _31089_);
  xor g_61512_(_29817_, _31088_, _31090_);
  or g_61513_(_29822_, _31090_, _31091_);
  not g_61514_(_31091_, _31092_);
  xor g_61515_(_29821_, _31090_, _31094_);
  not g_61516_(_31094_, _31095_);
  and g_61517_(_29825_, _29830_, _31096_);
  xor g_61518_(_31095_, _31096_, _31097_);
  xor g_61519_(_31094_, _31096_, _31098_);
  and g_61520_(_29835_, _31098_, _31099_);
  or g_61521_(_29834_, _31097_, _31100_);
  xor g_61522_(_29834_, _31098_, _31101_);
  not g_61523_(_31101_, _31102_);
  and g_61524_(_29837_, _29841_, _31103_);
  xor g_61525_(_31102_, _31103_, _31105_);
  xor g_61526_(_31101_, _31103_, _31106_);
  or g_61527_(_29844_, _31105_, _31107_);
  xor g_61528_(_29844_, _31106_, _31108_);
  or g_61529_(_29846_, _31108_, _31109_);
  not g_61530_(_31109_, _31110_);
  and g_61531_(_29846_, _31108_, _31111_);
  xor g_61532_(_29846_, _31108_, _31112_);
  or g_61533_(_31110_, _31111_, _31113_);
  or g_61534_(_29849_, _31113_, _31114_);
  xor g_61535_(_29849_, _31112_, _31116_);
  or g_61536_(_29854_, _31116_, _31117_);
  not g_61537_(_31117_, _31118_);
  xor g_61538_(_29853_, _31116_, _31119_);
  not g_61539_(_31119_, _31120_);
  or g_61540_(_29856_, _31119_, _31121_);
  xor g_61541_(_29856_, _31120_, _31122_);
  not g_61542_(_31122_, _31123_);
  or g_61543_(_29859_, _31122_, _31124_);
  xor g_61544_(_29859_, _31123_, _31125_);
  not g_61545_(_31125_, _31127_);
  and g_61546_(_29863_, _29865_, _31128_);
  xor g_61547_(_31127_, _31128_, _31129_);
  xor g_61548_(_29869_, _31129_, _31130_);
  or g_61549_(_29875_, _31130_, _31131_);
  not g_61550_(_31131_, _31132_);
  and g_61551_(_29872_, _31130_, _31133_);
  and g_61552_(_29875_, _31133_, _31134_);
  or g_61553_(_29872_, _31130_, _31135_);
  not g_61554_(_31135_, _31136_);
  or g_61555_(_31134_, _31136_, _31138_);
  or g_61556_(_31132_, _31138_, _31139_);
  not g_61557_(_31139_, _31140_);
  and g_61558_(_29879_, _29881_, _31141_);
  xor g_61559_(_31140_, _31141_, _31142_);
  or g_61560_(_29877_, _31142_, _31143_);
  xor g_61561_(_29878_, _31142_, _31144_);
  not g_61562_(_31144_, _31145_);
  or g_61563_(_29887_, _31144_, _31146_);
  xor g_61564_(_29887_, _31145_, _31147_);
  or g_61565_(_29955_, _31147_, _31149_);
  xor g_61566_(_29954_, _31147_, _31150_);
  or g_61567_(_29953_, _31150_, _31151_);
  xor g_61568_(_29952_, _31150_, _31152_);
  or g_61569_(_28692_, _29890_, _31153_);
  not g_61570_(_31153_, _31154_);
  or g_61571_(_31152_, _31153_, _31155_);
  xor g_61572_(_31152_, _31154_, _31156_);
  or g_61573_(_29950_, _31156_, _31157_);
  xor g_61574_(_29951_, _31156_, _31158_);
  or g_61575_(_29948_, _31158_, _31160_);
  xor g_61576_(_29948_, _31158_, _31161_);
  not g_61577_(_31161_, _31162_);
  and g_61578_(_29893_, _29898_, _31163_);
  xor g_61579_(_31161_, _31163_, _31164_);
  not g_61580_(_31164_, _31165_);
  xor g_61581_(_29947_, _31165_, _31166_);
  not g_61582_(_31166_, _31167_);
  xor g_61583_(_29946_, _31167_, _31168_);
  and g_61584_(_29914_, _31168_, _31169_);
  and g_61585_(_29916_, _31169_, _31171_);
  not g_61586_(_31171_, _31172_);
  or g_61587_(_29916_, _31168_, _31173_);
  or g_61588_(_29914_, _31168_, _31174_);
  and g_61589_(_31173_, _31174_, _31175_);
  not g_61590_(_31175_, _31176_);
  and g_61591_(_31172_, _31175_, _31177_);
  or g_61592_(_31171_, _31176_, _31178_);
  or g_61593_(_29920_, _31178_, _31179_);
  xor g_61594_(_29920_, _31177_, _31180_);
  not g_61595_(_31180_, _31182_);
  or g_61596_(_29923_, _31180_, _31183_);
  xor g_61597_(_29923_, _31182_, _31184_);
  or g_61598_(_29926_, _31184_, _31185_);
  not g_61599_(_31185_, _31186_);
  xor g_61600_(_29926_, _31184_, _31187_);
  xor g_61601_(_29927_, _31184_, _31188_);
  and g_61602_(_29931_, _29934_, _31189_);
  xor g_61603_(_31187_, _31189_, _31190_);
  not g_61604_(_31190_, _31191_);
  and g_61605_(_29937_, _31191_, _31193_);
  or g_61606_(_29936_, _31190_, _31194_);
  xor g_61607_(_29936_, _31190_, _31195_);
  not g_61608_(_31195_, _31196_);
  and g_61609_(_29945_, _31195_, _31197_);
  or g_61610_(_29944_, _31196_, _31198_);
  xor g_61611_(_29944_, _31195_, _31199_);
  or g_61612_(_28732_, _29938_, _31200_);
  and g_61613_(_29943_, _31200_, _31201_);
  xor g_61614_(_31199_, _31201_, out[643]);
  or g_61615_(_29943_, _31199_, _31203_);
  or g_61616_(_31199_, _31200_, _31204_);
  not g_61617_(_31204_, _31205_);
  or g_61618_(_29934_, _31188_, _31206_);
  or g_61619_(_29910_, _31166_, _31207_);
  or g_61620_(_29908_, _31166_, _31208_);
  or g_61621_(_29904_, _31164_, _31209_);
  not g_61622_(_31209_, _31210_);
  or g_61623_(_29901_, _31164_, _31211_);
  or g_61624_(_29898_, _31162_, _31212_);
  not g_61625_(_31212_, _31214_);
  or g_61626_(_29881_, _31139_, _31215_);
  or g_61627_(_29866_, _31129_, _31216_);
  or g_61628_(_28652_, _31216_, _31217_);
  or g_61629_(_28649_, _31216_, _31218_);
  or g_61630_(_29865_, _31125_, _31219_);
  or g_61631_(_29841_, _31101_, _31220_);
  or g_61632_(_29830_, _31094_, _31221_);
  or g_61633_(_29825_, _31094_, _31222_);
  or g_61634_(_29811_, _31076_, _31223_);
  or g_61635_(_29808_, _31076_, _31225_);
  or g_61636_(_29758_, _31014_, _31226_);
  or g_61637_(_29755_, _31011_, _31227_);
  or g_61638_(_29742_, _31002_, _31228_);
  not g_61639_(_31228_, _31229_);
  or g_61640_(_29735_, _30998_, _31230_);
  or g_61641_(_28550_, _31230_, _31231_);
  not g_61642_(_31231_, _31232_);
  or g_61643_(_28547_, _31230_, _31233_);
  not g_61644_(_31233_, _31234_);
  or g_61645_(_29726_, _30993_, _31236_);
  not g_61646_(_31236_, _31237_);
  and g_61647_(_29723_, _30992_, _31238_);
  or g_61648_(_29722_, _30993_, _31239_);
  or g_61649_(_29717_, _30989_, _31240_);
  or g_61650_(_29710_, _30989_, _31241_);
  or g_61651_(_29964_, _30975_, _31242_);
  or g_61652_(_29679_, _30952_, _31243_);
  or g_61653_(_29662_, _30941_, _31244_);
  or g_61654_(_29659_, _30937_, _31245_);
  or g_61655_(_29656_, _30937_, _31247_);
  or g_61656_(_29654_, _30934_, _31248_);
  or g_61657_(_29651_, _30934_, _31249_);
  or g_61658_(_29644_, _30926_, _31250_);
  and g_61659_(_30921_, _30924_, _31251_);
  or g_61660_(_30922_, _30923_, _31252_);
  or g_61661_(_30916_, _30919_, _31253_);
  not g_61662_(_31253_, _31254_);
  or g_61663_(_29633_, _30916_, _31255_);
  or g_61664_(_29612_, _30888_, _31256_);
  or g_61665_(_29608_, _30888_, _31258_);
  or g_61666_(_30882_, _30883_, _31259_);
  or g_61667_(_29603_, _30882_, _31260_);
  and g_61668_(_30865_, _30878_, _31261_);
  and g_61669_(_29582_, _30852_, _31262_);
  or g_61670_(_29583_, _30853_, _31263_);
  or g_61671_(_29579_, _30853_, _31264_);
  and g_61672_(_30847_, _30850_, _31265_);
  or g_61673_(_30832_, _30834_, _31266_);
  or g_61674_(_29530_, _30797_, _31267_);
  not g_61675_(_31267_, _31269_);
  or g_61676_(_30797_, _30798_, _31270_);
  not g_61677_(_31270_, _31271_);
  or g_61678_(_28317_, _29513_, _31272_);
  or g_61679_(_30768_, _31272_, _31273_);
  or g_61680_(_28313_, _29513_, _31274_);
  or g_61681_(_30768_, _31274_, _31275_);
  not g_61682_(_31275_, _31276_);
  or g_61683_(_30003_, _30759_, _31277_);
  not g_61684_(_31277_, _31278_);
  and g_61685_(_29508_, _30758_, _31280_);
  or g_61686_(_29507_, _30759_, _31281_);
  or g_61687_(_29505_, _30757_, _31282_);
  not g_61688_(_31282_, _31283_);
  or g_61689_(_29502_, _30757_, _31284_);
  not g_61690_(_31284_, _31285_);
  or g_61691_(_29498_, _30753_, _31286_);
  not g_61692_(_31286_, _31287_);
  and g_61693_(_30751_, _30755_, _31288_);
  not g_61694_(_31288_, _31289_);
  or g_61695_(_30748_, _30749_, _31291_);
  not g_61696_(_31291_, _31292_);
  or g_61697_(_29482_, _30737_, _31293_);
  not g_61698_(_31293_, _31294_);
  or g_61699_(_29480_, _30737_, _31295_);
  not g_61700_(_31295_, _31296_);
  or g_61701_(_29478_, _30734_, _31297_);
  not g_61702_(_31297_, _31298_);
  or g_61703_(_30726_, _30728_, _31299_);
  not g_61704_(_31299_, _31300_);
  or g_61705_(_30726_, _30727_, _31302_);
  not g_61706_(_31302_, _31303_);
  and g_61707_(_29463_, _30713_, _31304_);
  or g_61708_(_29462_, _30714_, _31305_);
  or g_61709_(_29454_, _30711_, _31306_);
  not g_61710_(_31306_, _31307_);
  or g_61711_(_29451_, _30711_, _31308_);
  not g_61712_(_31308_, _31309_);
  or g_61713_(_30674_, _30677_, _31310_);
  not g_61714_(_31310_, _31311_);
  or g_61715_(_30674_, _30679_, _31313_);
  or g_61716_(_30017_, _30672_, _31314_);
  or g_61717_(_29425_, _30672_, _31315_);
  not g_61718_(_31315_, _31316_);
  and g_61719_(_29421_, _30670_, _31317_);
  not g_61720_(_31317_, _31318_);
  or g_61721_(_29417_, _30669_, _31319_);
  not g_61722_(_31319_, _31320_);
  or g_61723_(_29414_, _30667_, _31321_);
  not g_61724_(_31321_, _31322_);
  or g_61725_(_30658_, _30660_, _31324_);
  or g_61726_(_29406_, _30658_, _31325_);
  or g_61727_(_30641_, _30644_, _31326_);
  or g_61728_(_30641_, _30643_, _31327_);
  not g_61729_(_31327_, _31328_);
  and g_61730_(_30638_, _30640_, _31329_);
  or g_61731_(_29342_, _30593_, _31330_);
  not g_61732_(_31330_, _31331_);
  or g_61733_(_29331_, _30586_, _31332_);
  not g_61734_(_31332_, _31333_);
  or g_61735_(_29328_, _30581_, _31335_);
  or g_61736_(_29309_, _30573_, _31336_);
  or g_61737_(_30547_, _30548_, _31337_);
  or g_61738_(_29286_, _30547_, _31338_);
  and g_61739_(_29276_, _30530_, _31339_);
  not g_61740_(_31339_, _31340_);
  or g_61741_(_29266_, _30503_, _31341_);
  not g_61742_(_31341_, _31342_);
  or g_61743_(_29244_, _30474_, _31343_);
  not g_61744_(_31343_, _31344_);
  or g_61745_(_30467_, _30469_, _31346_);
  and g_61746_(_30437_, _30440_, _31347_);
  and g_61747_(_30432_, _30435_, _31348_);
  not g_61748_(_31348_, _31349_);
  and g_61749_(_30416_, _30430_, _31350_);
  or g_61750_(_29184_, _30407_, _31351_);
  not g_61751_(_31351_, _31352_);
  or g_61752_(_29171_, _30402_, _31353_);
  or g_61753_(_29172_, _30402_, _31354_);
  or g_61754_(_30395_, _30396_, _31355_);
  and g_61755_(_29144_, _30370_, _31357_);
  not g_61756_(_31357_, _31358_);
  or g_61757_(_30371_, _30372_, _31359_);
  not g_61758_(_31359_, _31360_);
  or g_61759_(_29132_, _30357_, _31361_);
  or g_61760_(_29130_, _30357_, _31362_);
  or g_61761_(_29122_, _30351_, _31363_);
  or g_61762_(_29117_, _30351_, _31364_);
  and g_61763_(_30342_, _30346_, _31365_);
  and g_61764_(_30337_, _30340_, _31366_);
  not g_61765_(_31366_, _31368_);
  or g_61766_(_30067_, _30300_, _31369_);
  or g_61767_(_29068_, _30287_, _31370_);
  or g_61768_(_27823_, _31370_, _31371_);
  or g_61769_(_27821_, _31370_, _31372_);
  or g_61770_(_29042_, _30258_, _31373_);
  not g_61771_(_31373_, _31374_);
  and g_61772_(_29039_, _30255_, _31375_);
  not g_61773_(_31375_, _31376_);
  or g_61774_(_29035_, _30254_, _31377_);
  or g_61775_(_29032_, _30252_, _31379_);
  or g_61776_(_29029_, _30252_, _31380_);
  or g_61777_(_30220_, _30222_, _31381_);
  or g_61778_(_29011_, _30220_, _31382_);
  and g_61779_(_30206_, _30208_, _31383_);
  or g_61780_(_27706_, _28981_, _31384_);
  or g_61781_(_30192_, _31384_, _31385_);
  or g_61782_(_28985_, _30192_, _31386_);
  or g_61783_(_28968_, _30179_, _31387_);
  and g_61784_(_30184_, _31387_, _31388_);
  and g_61785_(_28940_, _30153_, _31390_);
  or g_61786_(_28939_, _30154_, _31391_);
  or g_61787_(_30150_, _30155_, _31392_);
  or g_61788_(_28925_, _30140_, _31393_);
  and g_61789_(_30139_, _31393_, _31394_);
  or g_61790_(_30131_, _30133_, _31395_);
  and g_61791_(_30108_, _30118_, _31396_);
  and g_61792_(_30115_, _31396_, _31397_);
  and g_61793_(_30121_, _30124_, _31398_);
  and g_61794_(_31397_, _31398_, _31399_);
  and g_61795_(_30128_, _31399_, _31401_);
  and g_61796_(_30130_, _31401_, _31402_);
  and g_61797_(_31395_, _31402_, _31403_);
  or g_61798_(_30132_, _30134_, _31404_);
  and g_61799_(_31403_, _31404_, _31405_);
  and g_61800_(_31394_, _31405_, _31406_);
  and g_61801_(_30143_, _31406_, _31407_);
  and g_61802_(_30146_, _31407_, _31408_);
  and g_61803_(_30149_, _30152_, _31409_);
  or g_61804_(_31408_, _31409_, _31410_);
  xor g_61805_(_31408_, _31409_, _31412_);
  not g_61806_(_31412_, _31413_);
  or g_61807_(_31392_, _31413_, _31414_);
  xor g_61808_(_31392_, _31412_, _31415_);
  or g_61809_(_31391_, _31415_, _31416_);
  xor g_61810_(_31390_, _31415_, _31417_);
  and g_61811_(_28950_, _30159_, _31418_);
  or g_61812_(_30160_, _31418_, _31419_);
  not g_61813_(_31419_, _31420_);
  and g_61814_(_31417_, _31419_, _31421_);
  or g_61815_(_31417_, _31419_, _31423_);
  xor g_61816_(_31417_, _31420_, _31424_);
  not g_61817_(_31424_, _31425_);
  or g_61818_(_28952_, _30161_, _31426_);
  and g_61819_(_30173_, _31426_, _31427_);
  xor g_61820_(_31425_, _31427_, _31428_);
  or g_61821_(_30166_, _31428_, _31429_);
  xor g_61822_(_30167_, _31428_, _31430_);
  not g_61823_(_31430_, _31431_);
  and g_61824_(_28962_, _28965_, _31432_);
  or g_61825_(_30178_, _31432_, _31434_);
  or g_61826_(_31430_, _31434_, _31435_);
  xor g_61827_(_31430_, _31434_, _31436_);
  xor g_61828_(_31431_, _31434_, _31437_);
  or g_61829_(_31388_, _31437_, _31438_);
  xor g_61830_(_31388_, _31436_, _31439_);
  not g_61831_(_31439_, _31440_);
  or g_61832_(_30187_, _31439_, _31441_);
  xor g_61833_(_30187_, _31440_, _31442_);
  or g_61834_(_30190_, _31442_, _31443_);
  xor g_61835_(_30190_, _31442_, _31445_);
  not g_61836_(_31445_, _31446_);
  or g_61837_(_31386_, _31446_, _31447_);
  xor g_61838_(_31386_, _31446_, _31448_);
  xor g_61839_(_31386_, _31445_, _31449_);
  or g_61840_(_31385_, _31449_, _31450_);
  xor g_61841_(_31385_, _31448_, _31451_);
  not g_61842_(_31451_, _31452_);
  or g_61843_(_30195_, _31451_, _31453_);
  xor g_61844_(_30195_, _31451_, _31454_);
  xor g_61845_(_30195_, _31452_, _31456_);
  or g_61846_(_30196_, _31456_, _31457_);
  xor g_61847_(_30196_, _31454_, _31458_);
  or g_61848_(_30203_, _31458_, _31459_);
  or g_61849_(_30201_, _31454_, _31460_);
  and g_61850_(_31459_, _31460_, _31461_);
  xor g_61851_(_31383_, _31461_, _31462_);
  or g_61852_(_30217_, _31462_, _31463_);
  and g_61853_(_30217_, _31462_, _31464_);
  xor g_61854_(_30218_, _31462_, _31465_);
  xor g_61855_(_30216_, _31465_, _31467_);
  and g_61856_(_31382_, _31467_, _31468_);
  and g_61857_(_31381_, _31468_, _31469_);
  or g_61858_(_31382_, _31465_, _31470_);
  and g_61859_(_31381_, _31470_, _31471_);
  or g_61860_(_31468_, _31471_, _31472_);
  not g_61861_(_31472_, _31473_);
  or g_61862_(_31469_, _31473_, _31474_);
  not g_61863_(_31474_, _31475_);
  or g_61864_(_30226_, _31474_, _31476_);
  and g_61865_(_30226_, _31474_, _31478_);
  xor g_61866_(_30226_, _31474_, _31479_);
  xor g_61867_(_30226_, _31475_, _31480_);
  or g_61868_(_30232_, _31480_, _31481_);
  not g_61869_(_31481_, _31482_);
  or g_61870_(_30230_, _31480_, _31483_);
  or g_61871_(_30229_, _31479_, _31484_);
  and g_61872_(_30232_, _31484_, _31485_);
  and g_61873_(_31483_, _31485_, _31486_);
  or g_61874_(_31482_, _31486_, _31487_);
  not g_61875_(_31487_, _31489_);
  and g_61876_(_30236_, _30239_, _31490_);
  xor g_61877_(_31487_, _31490_, _31491_);
  xor g_61878_(_31489_, _31490_, _31492_);
  or g_61879_(_30243_, _31492_, _31493_);
  xor g_61880_(_30243_, _31491_, _31494_);
  or g_61881_(_30245_, _31494_, _31495_);
  not g_61882_(_31495_, _31496_);
  xor g_61883_(_30247_, _31494_, _31497_);
  not g_61884_(_31497_, _31498_);
  or g_61885_(_30251_, _31497_, _31500_);
  xor g_61886_(_30251_, _31497_, _31501_);
  xor g_61887_(_30251_, _31498_, _31502_);
  or g_61888_(_31380_, _31502_, _31503_);
  xor g_61889_(_31380_, _31501_, _31504_);
  or g_61890_(_31379_, _31504_, _31505_);
  not g_61891_(_31505_, _31506_);
  xor g_61892_(_31379_, _31504_, _31507_);
  not g_61893_(_31507_, _31508_);
  or g_61894_(_31377_, _31508_, _31509_);
  not g_61895_(_31509_, _31511_);
  xor g_61896_(_31377_, _31507_, _31512_);
  not g_61897_(_31512_, _31513_);
  and g_61898_(_31375_, _31513_, _31514_);
  or g_61899_(_31376_, _31512_, _31515_);
  xor g_61900_(_31375_, _31512_, _31516_);
  or g_61901_(_31373_, _31516_, _31517_);
  and g_61902_(_31373_, _31516_, _31518_);
  xor g_61903_(_31374_, _31516_, _31519_);
  or g_61904_(_30076_, _30258_, _31520_);
  and g_61905_(_30262_, _31520_, _31522_);
  xor g_61906_(_31519_, _31522_, _31523_);
  not g_61907_(_31523_, _31524_);
  or g_61908_(_30260_, _31524_, _31525_);
  xor g_61909_(_30260_, _31523_, _31526_);
  not g_61910_(_31526_, _31527_);
  and g_61911_(_30271_, _31527_, _31528_);
  not g_61912_(_31528_, _31529_);
  or g_61913_(_30266_, _31526_, _31530_);
  xor g_61914_(_30266_, _31526_, _31531_);
  not g_61915_(_31531_, _31533_);
  and g_61916_(_30275_, _31531_, _31534_);
  or g_61917_(_30274_, _31533_, _31535_);
  xor g_61918_(_30274_, _31531_, _31536_);
  and g_61919_(_30270_, _31536_, _31537_);
  or g_61920_(_31528_, _31537_, _31538_);
  and g_61921_(_30278_, _30282_, _31539_);
  or g_61922_(_31538_, _31539_, _31540_);
  not g_61923_(_31540_, _31541_);
  and g_61924_(_31538_, _31539_, _31542_);
  xor g_61925_(_31538_, _31539_, _31544_);
  or g_61926_(_31541_, _31542_, _31545_);
  or g_61927_(_30285_, _31545_, _31546_);
  not g_61928_(_31546_, _31547_);
  xor g_61929_(_30285_, _31544_, _31548_);
  not g_61930_(_31548_, _31549_);
  or g_61931_(_31372_, _31548_, _31550_);
  xor g_61932_(_31372_, _31549_, _31551_);
  or g_61933_(_31371_, _31551_, _31552_);
  xor g_61934_(_31371_, _31551_, _31553_);
  xor g_61935_(_30291_, _31553_, _31555_);
  or g_61936_(_30297_, _31555_, _31556_);
  and g_61937_(_30297_, _31555_, _31557_);
  xor g_61938_(_30297_, _31555_, _31558_);
  and g_61939_(_30294_, _31558_, _31559_);
  xor g_61940_(_30295_, _31558_, _31560_);
  or g_61941_(_29084_, _30300_, _31561_);
  not g_61942_(_31561_, _31562_);
  or g_61943_(_31560_, _31561_, _31563_);
  not g_61944_(_31563_, _31564_);
  xor g_61945_(_31560_, _31562_, _31566_);
  not g_61946_(_31566_, _31567_);
  or g_61947_(_31369_, _31566_, _31568_);
  xor g_61948_(_31369_, _31567_, _31569_);
  not g_61949_(_31569_, _31570_);
  or g_61950_(_30304_, _31569_, _31571_);
  xor g_61951_(_30304_, _31570_, _31572_);
  or g_61952_(_30307_, _31572_, _31573_);
  not g_61953_(_31573_, _31574_);
  xor g_61954_(_30308_, _31572_, _31575_);
  not g_61955_(_31575_, _31577_);
  and g_61956_(_30311_, _31575_, _31578_);
  and g_61957_(_30314_, _31578_, _31579_);
  or g_61958_(_30311_, _31575_, _31580_);
  and g_61959_(_30315_, _31577_, _31581_);
  or g_61960_(_30314_, _31575_, _31582_);
  and g_61961_(_31580_, _31582_, _31583_);
  not g_61962_(_31583_, _31584_);
  or g_61963_(_31579_, _31584_, _31585_);
  not g_61964_(_31585_, _31586_);
  and g_61965_(_30317_, _31586_, _31588_);
  xor g_61966_(_30317_, _31586_, _31589_);
  xor g_61967_(_30317_, _31585_, _31590_);
  or g_61968_(_30320_, _31590_, _31591_);
  not g_61969_(_31591_, _31592_);
  xor g_61970_(_30320_, _31589_, _31593_);
  not g_61971_(_31593_, _31594_);
  or g_61972_(_30326_, _31593_, _31595_);
  xor g_61973_(_30326_, _31594_, _31596_);
  not g_61974_(_31596_, _31597_);
  or g_61975_(_30325_, _31596_, _31599_);
  xor g_61976_(_30325_, _31597_, _31600_);
  xor g_61977_(_30333_, _31600_, _31601_);
  xor g_61978_(_31368_, _31601_, _31602_);
  not g_61979_(_31602_, _31603_);
  xor g_61980_(_31365_, _31602_, _31604_);
  and g_61981_(_30348_, _31604_, _31605_);
  not g_61982_(_31605_, _31606_);
  xor g_61983_(_30348_, _31604_, _31607_);
  not g_61984_(_31607_, _31608_);
  or g_61985_(_31364_, _31608_, _31610_);
  not g_61986_(_31610_, _31611_);
  xor g_61987_(_31364_, _31607_, _31612_);
  not g_61988_(_31612_, _31613_);
  or g_61989_(_31363_, _31612_, _31614_);
  xor g_61990_(_31363_, _31612_, _31615_);
  xor g_61991_(_31363_, _31613_, _31616_);
  and g_61992_(_30355_, _31615_, _31617_);
  or g_61993_(_30354_, _31616_, _31618_);
  xor g_61994_(_30354_, _31615_, _31619_);
  not g_61995_(_31619_, _31621_);
  or g_61996_(_31362_, _31619_, _31622_);
  xor g_61997_(_31362_, _31621_, _31623_);
  not g_61998_(_31623_, _31624_);
  or g_61999_(_31361_, _31623_, _31625_);
  xor g_62000_(_31361_, _31623_, _31626_);
  xor g_62001_(_31361_, _31624_, _31627_);
  or g_62002_(_30364_, _31627_, _31628_);
  or g_62003_(_30361_, _31627_, _31629_);
  xor g_62004_(_30361_, _31626_, _31630_);
  or g_62005_(_30369_, _31630_, _31632_);
  xor g_62006_(_30369_, _31630_, _31633_);
  or g_62007_(_30365_, _31633_, _31634_);
  and g_62008_(_31628_, _31634_, _31635_);
  not g_62009_(_31635_, _31636_);
  and g_62010_(_31360_, _31635_, _31637_);
  or g_62011_(_31359_, _31636_, _31638_);
  xor g_62012_(_31359_, _31635_, _31639_);
  not g_62013_(_31639_, _31640_);
  and g_62014_(_31357_, _31640_, _31641_);
  or g_62015_(_31358_, _31639_, _31643_);
  xor g_62016_(_31357_, _31639_, _31644_);
  xor g_62017_(_30376_, _31644_, _31645_);
  or g_62018_(_30380_, _31645_, _31646_);
  not g_62019_(_31646_, _31647_);
  xor g_62020_(_30381_, _31645_, _31648_);
  not g_62021_(_31648_, _31649_);
  and g_62022_(_30383_, _30388_, _31650_);
  xor g_62023_(_31648_, _31650_, _31651_);
  not g_62024_(_31651_, _31652_);
  or g_62025_(_30386_, _31652_, _31654_);
  xor g_62026_(_30386_, _31651_, _31655_);
  not g_62027_(_31655_, _31656_);
  or g_62028_(_29166_, _30395_, _31657_);
  and g_62029_(_30392_, _31657_, _31658_);
  xor g_62030_(_31656_, _31658_, _31659_);
  not g_62031_(_31659_, _31660_);
  or g_62032_(_31355_, _31659_, _31661_);
  xor g_62033_(_31355_, _31660_, _31662_);
  or g_62034_(_30401_, _31662_, _31663_);
  not g_62035_(_31663_, _31665_);
  xor g_62036_(_30399_, _31662_, _31666_);
  not g_62037_(_31666_, _31667_);
  or g_62038_(_31354_, _31666_, _31668_);
  xor g_62039_(_31354_, _31666_, _31669_);
  xor g_62040_(_31354_, _31667_, _31670_);
  or g_62041_(_31353_, _31670_, _31671_);
  xor g_62042_(_31353_, _31669_, _31672_);
  or g_62043_(_29182_, _30407_, _31673_);
  and g_62044_(_30406_, _31673_, _31674_);
  xor g_62045_(_31672_, _31674_, _31676_);
  and g_62046_(_31352_, _31676_, _31677_);
  not g_62047_(_31677_, _31678_);
  xor g_62048_(_31352_, _31676_, _31679_);
  not g_62049_(_31679_, _31680_);
  or g_62050_(_30413_, _31680_, _31681_);
  not g_62051_(_31681_, _31682_);
  xor g_62052_(_30413_, _31679_, _31683_);
  not g_62053_(_31683_, _31684_);
  or g_62054_(_30423_, _31683_, _31685_);
  not g_62055_(_31685_, _31687_);
  or g_62056_(_30426_, _31683_, _31688_);
  xor g_62057_(_30426_, _31683_, _31689_);
  xor g_62058_(_30426_, _31684_, _31690_);
  and g_62059_(_30423_, _31690_, _31691_);
  or g_62060_(_30421_, _31689_, _31692_);
  and g_62061_(_31685_, _31692_, _31693_);
  or g_62062_(_31687_, _31691_, _31694_);
  xor g_62063_(_31350_, _31693_, _31695_);
  xor g_62064_(_31348_, _31695_, _31696_);
  xor g_62065_(_31349_, _31695_, _31698_);
  xor g_62066_(_31347_, _31696_, _31699_);
  or g_62067_(_30445_, _31699_, _31700_);
  not g_62068_(_31700_, _31701_);
  or g_62069_(_30442_, _31699_, _31702_);
  xor g_62070_(_30442_, _31699_, _31703_);
  not g_62071_(_31703_, _31704_);
  or g_62072_(_30447_, _31704_, _31705_);
  not g_62073_(_31705_, _31706_);
  xor g_62074_(_30447_, _31703_, _31707_);
  and g_62075_(_30445_, _31707_, _31709_);
  or g_62076_(_31701_, _31709_, _31710_);
  and g_62077_(_30449_, _30457_, _31711_);
  or g_62078_(_31710_, _31711_, _31712_);
  xor g_62079_(_31710_, _31711_, _31713_);
  and g_62080_(_30460_, _31713_, _31714_);
  xor g_62081_(_30459_, _31713_, _31715_);
  not g_62082_(_31715_, _31716_);
  or g_62083_(_29236_, _30467_, _31717_);
  and g_62084_(_30465_, _31717_, _31718_);
  xor g_62085_(_31716_, _31718_, _31720_);
  or g_62086_(_31346_, _31720_, _31721_);
  xor g_62087_(_31346_, _31720_, _31722_);
  not g_62088_(_31722_, _31723_);
  or g_62089_(_29241_, _30474_, _31724_);
  not g_62090_(_31724_, _31725_);
  and g_62091_(_30473_, _31724_, _31726_);
  xor g_62092_(_31722_, _31726_, _31727_);
  or g_62093_(_31343_, _31727_, _31728_);
  xor g_62094_(_31343_, _31727_, _31729_);
  xor g_62095_(_31344_, _31727_, _31731_);
  and g_62096_(_30481_, _30485_, _31732_);
  or g_62097_(_30480_, _30484_, _31733_);
  and g_62098_(_31731_, _31732_, _31734_);
  or g_62099_(_31729_, _31733_, _31735_);
  and g_62100_(_30484_, _31729_, _31736_);
  or g_62101_(_30485_, _31731_, _31737_);
  and g_62102_(_30480_, _31729_, _31738_);
  or g_62103_(_30481_, _31731_, _31739_);
  and g_62104_(_31737_, _31739_, _31740_);
  or g_62105_(_31736_, _31738_, _31742_);
  and g_62106_(_31735_, _31740_, _31743_);
  or g_62107_(_31734_, _31742_, _31744_);
  or g_62108_(_30487_, _31744_, _31745_);
  not g_62109_(_31745_, _31746_);
  or g_62110_(_30491_, _31744_, _31747_);
  not g_62111_(_31747_, _31748_);
  xor g_62112_(_30491_, _31743_, _31749_);
  and g_62113_(_30487_, _31749_, _31750_);
  or g_62114_(_31746_, _31750_, _31751_);
  not g_62115_(_31751_, _31753_);
  and g_62116_(_30494_, _30496_, _31754_);
  not g_62117_(_31754_, _31755_);
  xor g_62118_(_31751_, _31755_, _31756_);
  xor g_62119_(_31751_, _31754_, _31757_);
  or g_62120_(_31341_, _31756_, _31758_);
  not g_62121_(_31758_, _31759_);
  or g_62122_(_30501_, _31756_, _31760_);
  not g_62123_(_31760_, _31761_);
  and g_62124_(_31758_, _31760_, _31762_);
  not g_62125_(_31762_, _31764_);
  and g_62126_(_30501_, _31756_, _31765_);
  or g_62127_(_30502_, _31757_, _31766_);
  and g_62128_(_31341_, _31765_, _31767_);
  or g_62129_(_31342_, _31766_, _31768_);
  and g_62130_(_31762_, _31768_, _31769_);
  or g_62131_(_31764_, _31767_, _31770_);
  or g_62132_(_29269_, _30503_, _31771_);
  or g_62133_(_31770_, _31771_, _31772_);
  xor g_62134_(_31769_, _31771_, _31773_);
  or g_62135_(_30511_, _31773_, _31775_);
  not g_62136_(_31775_, _31776_);
  and g_62137_(_30507_, _31773_, _31777_);
  and g_62138_(_30511_, _31777_, _31778_);
  or g_62139_(_30507_, _31770_, _31779_);
  not g_62140_(_31779_, _31780_);
  or g_62141_(_31778_, _31780_, _31781_);
  or g_62142_(_31776_, _31781_, _31782_);
  or g_62143_(_30515_, _31782_, _31783_);
  xor g_62144_(_30516_, _31782_, _31784_);
  or g_62145_(_30524_, _31784_, _31786_);
  not g_62146_(_31786_, _31787_);
  or g_62147_(_30527_, _31784_, _31788_);
  xor g_62148_(_30528_, _31784_, _31789_);
  and g_62149_(_30524_, _31789_, _31790_);
  or g_62150_(_31787_, _31790_, _31791_);
  or g_62151_(_30529_, _30531_, _31792_);
  not g_62152_(_31792_, _31793_);
  or g_62153_(_31791_, _31792_, _31794_);
  not g_62154_(_31794_, _31795_);
  xor g_62155_(_31791_, _31793_, _31797_);
  not g_62156_(_31797_, _31798_);
  and g_62157_(_31339_, _31798_, _31799_);
  or g_62158_(_31340_, _31797_, _31800_);
  xor g_62159_(_31339_, _31797_, _31801_);
  xor g_62160_(_30540_, _31801_, _31802_);
  or g_62161_(_30542_, _31802_, _31803_);
  xor g_62162_(_30544_, _31802_, _31804_);
  not g_62163_(_31804_, _31805_);
  or g_62164_(_31338_, _31804_, _31806_);
  xor g_62165_(_31338_, _31804_, _31808_);
  xor g_62166_(_31338_, _31805_, _31809_);
  or g_62167_(_31337_, _31809_, _31810_);
  xor g_62168_(_31337_, _31808_, _31811_);
  or g_62169_(_30552_, _30556_, _31812_);
  xor g_62170_(_31811_, _31812_, _31813_);
  or g_62171_(_30563_, _31813_, _31814_);
  xor g_62172_(_30564_, _31813_, _31815_);
  or g_62173_(_30559_, _31815_, _31816_);
  xor g_62174_(_30560_, _31815_, _31817_);
  or g_62175_(_30569_, _31817_, _31819_);
  xor g_62176_(_30570_, _31817_, _31820_);
  or g_62177_(_31336_, _31820_, _31821_);
  not g_62178_(_31821_, _31822_);
  and g_62179_(_30572_, _31820_, _31823_);
  and g_62180_(_31336_, _31823_, _31824_);
  or g_62181_(_30572_, _31820_, _31825_);
  not g_62182_(_31825_, _31826_);
  or g_62183_(_31824_, _31826_, _31827_);
  or g_62184_(_31822_, _31827_, _31828_);
  not g_62185_(_31828_, _31830_);
  or g_62186_(_29313_, _30573_, _31831_);
  or g_62187_(_29316_, _30577_, _31832_);
  and g_62188_(_31831_, _31832_, _31833_);
  xor g_62189_(_31828_, _31833_, _31834_);
  xor g_62190_(_31830_, _31833_, _31835_);
  or g_62191_(_30582_, _31835_, _31836_);
  and g_62192_(_29319_, _30578_, _31837_);
  not g_62193_(_31837_, _31838_);
  or g_62194_(_31834_, _31837_, _31839_);
  or g_62195_(_30583_, _31839_, _31841_);
  or g_62196_(_31835_, _31838_, _31842_);
  and g_62197_(_31841_, _31842_, _31843_);
  and g_62198_(_31836_, _31843_, _31844_);
  not g_62199_(_31844_, _31845_);
  or g_62200_(_31335_, _31845_, _31846_);
  xor g_62201_(_31335_, _31844_, _31847_);
  or g_62202_(_31332_, _31847_, _31848_);
  xor g_62203_(_31333_, _31847_, _31849_);
  or g_62204_(_29340_, _30593_, _31850_);
  and g_62205_(_30591_, _31850_, _31852_);
  xor g_62206_(_31849_, _31852_, _31853_);
  and g_62207_(_31331_, _31853_, _31854_);
  xor g_62208_(_31330_, _31853_, _31855_);
  and g_62209_(_30596_, _30599_, _31856_);
  xor g_62210_(_31855_, _31856_, _31857_);
  not g_62211_(_31857_, _31858_);
  or g_62212_(_30606_, _31858_, _31859_);
  xor g_62213_(_30606_, _31857_, _31860_);
  or g_62214_(_30605_, _31860_, _31861_);
  xor g_62215_(_30604_, _31860_, _31863_);
  and g_62216_(_30611_, _30615_, _31864_);
  not g_62217_(_31864_, _31865_);
  xor g_62218_(_31863_, _31864_, _31866_);
  xor g_62219_(_31863_, _31865_, _31867_);
  or g_62220_(_30616_, _31866_, _31868_);
  or g_62221_(_30623_, _31868_, _31869_);
  or g_62222_(_30624_, _31867_, _31870_);
  or g_62223_(_30617_, _31867_, _31871_);
  not g_62224_(_31871_, _31872_);
  and g_62225_(_31870_, _31871_, _31874_);
  and g_62226_(_31869_, _31874_, _31875_);
  not g_62227_(_31875_, _31876_);
  or g_62228_(_30626_, _31876_, _31877_);
  xor g_62229_(_30626_, _31875_, _31878_);
  xor g_62230_(_30634_, _31878_, _31879_);
  xor g_62231_(_31329_, _31879_, _31880_);
  not g_62232_(_31880_, _31881_);
  or g_62233_(_31327_, _31881_, _31882_);
  xor g_62234_(_31328_, _31880_, _31883_);
  not g_62235_(_31883_, _31885_);
  or g_62236_(_31326_, _31885_, _31886_);
  xor g_62237_(_31326_, _31883_, _31887_);
  and g_62238_(_29393_, _30650_, _31888_);
  or g_62239_(_29392_, _30651_, _31889_);
  and g_62240_(_30649_, _31889_, _31890_);
  or g_62241_(_30648_, _31888_, _31891_);
  or g_62242_(_31887_, _31890_, _31892_);
  xor g_62243_(_31887_, _31890_, _31893_);
  xor g_62244_(_31887_, _31891_, _31894_);
  and g_62245_(_30656_, _31893_, _31896_);
  not g_62246_(_31896_, _31897_);
  and g_62247_(_29398_, _30650_, _31898_);
  or g_62248_(_29397_, _30651_, _31899_);
  and g_62249_(_31893_, _31898_, _31900_);
  not g_62250_(_31900_, _31901_);
  and g_62251_(_31897_, _31901_, _31902_);
  or g_62252_(_31896_, _31900_, _31903_);
  and g_62253_(_31894_, _31899_, _31904_);
  and g_62254_(_30657_, _31904_, _31905_);
  or g_62255_(_31903_, _31905_, _31907_);
  or g_62256_(_31325_, _31907_, _31908_);
  xor g_62257_(_31325_, _31907_, _31909_);
  not g_62258_(_31909_, _31910_);
  or g_62259_(_31324_, _31910_, _31911_);
  xor g_62260_(_31324_, _31909_, _31912_);
  or g_62261_(_30663_, _31912_, _31913_);
  xor g_62262_(_30665_, _31912_, _31914_);
  and g_62263_(_29410_, _30666_, _31915_);
  not g_62264_(_31915_, _31916_);
  or g_62265_(_31914_, _31916_, _31918_);
  xor g_62266_(_31914_, _31915_, _31919_);
  or g_62267_(_31321_, _31919_, _31920_);
  not g_62268_(_31920_, _31921_);
  xor g_62269_(_31322_, _31919_, _31922_);
  or g_62270_(_31319_, _31922_, _31923_);
  xor g_62271_(_31320_, _31922_, _31924_);
  or g_62272_(_31318_, _31924_, _31925_);
  not g_62273_(_31925_, _31926_);
  xor g_62274_(_31317_, _31924_, _31927_);
  or g_62275_(_31315_, _31927_, _31929_);
  xor g_62276_(_31316_, _31927_, _31930_);
  and g_62277_(_31314_, _31930_, _31931_);
  or g_62278_(_31314_, _31930_, _31932_);
  not g_62279_(_31932_, _31933_);
  xor g_62280_(_31314_, _31930_, _31934_);
  or g_62281_(_31931_, _31933_, _31935_);
  or g_62282_(_31313_, _31935_, _31936_);
  xor g_62283_(_31313_, _31934_, _31937_);
  or g_62284_(_31310_, _31937_, _31938_);
  xor g_62285_(_31311_, _31937_, _31940_);
  or g_62286_(_30690_, _31940_, _31941_);
  xor g_62287_(_30691_, _31940_, _31942_);
  or g_62288_(_30696_, _31942_, _31943_);
  not g_62289_(_31943_, _31944_);
  or g_62290_(_30683_, _31942_, _31945_);
  xor g_62291_(_30683_, _31942_, _31946_);
  xor g_62292_(_30684_, _31942_, _31947_);
  and g_62293_(_30696_, _31947_, _31948_);
  or g_62294_(_30698_, _31946_, _31949_);
  and g_62295_(_31943_, _31949_, _31951_);
  or g_62296_(_31944_, _31948_, _31952_);
  and g_62297_(_30701_, _30705_, _31953_);
  xor g_62298_(_31952_, _31953_, _31954_);
  xor g_62299_(_31951_, _31953_, _31955_);
  and g_62300_(_30710_, _31955_, _31956_);
  and g_62301_(_31308_, _31956_, _31957_);
  and g_62302_(_31309_, _31954_, _31958_);
  or g_62303_(_31308_, _31955_, _31959_);
  and g_62304_(_30709_, _31954_, _31960_);
  or g_62305_(_30710_, _31955_, _31962_);
  or g_62306_(_31958_, _31960_, _31963_);
  or g_62307_(_31957_, _31963_, _31964_);
  or g_62308_(_31306_, _31964_, _31965_);
  xor g_62309_(_31306_, _31964_, _31966_);
  xor g_62310_(_31307_, _31964_, _31967_);
  and g_62311_(_29459_, _30713_, _31968_);
  or g_62312_(_29458_, _30714_, _31969_);
  and g_62313_(_31967_, _31969_, _31970_);
  and g_62314_(_31305_, _31970_, _31971_);
  and g_62315_(_31966_, _31968_, _31973_);
  and g_62316_(_31304_, _31966_, _31974_);
  or g_62317_(_31973_, _31974_, _31975_);
  or g_62318_(_31971_, _31975_, _31976_);
  or g_62319_(_30717_, _31976_, _31977_);
  xor g_62320_(_30718_, _31976_, _31978_);
  not g_62321_(_31978_, _31979_);
  or g_62322_(_30722_, _31978_, _31980_);
  xor g_62323_(_30722_, _31978_, _31981_);
  xor g_62324_(_30722_, _31979_, _31982_);
  or g_62325_(_30725_, _31982_, _31984_);
  xor g_62326_(_30725_, _31981_, _31985_);
  or g_62327_(_31302_, _31985_, _31986_);
  not g_62328_(_31986_, _31987_);
  xor g_62329_(_31303_, _31985_, _31988_);
  or g_62330_(_31299_, _31988_, _31989_);
  not g_62331_(_31989_, _31990_);
  xor g_62332_(_31299_, _31988_, _31991_);
  xor g_62333_(_31300_, _31988_, _31992_);
  or g_62334_(_29474_, _30734_, _31993_);
  and g_62335_(_30733_, _31993_, _31995_);
  xor g_62336_(_31991_, _31995_, _31996_);
  or g_62337_(_31297_, _31996_, _31997_);
  not g_62338_(_31997_, _31998_);
  xor g_62339_(_31298_, _31996_, _31999_);
  or g_62340_(_31295_, _31999_, _32000_);
  xor g_62341_(_31296_, _31999_, _32001_);
  or g_62342_(_31293_, _32001_, _32002_);
  not g_62343_(_32002_, _32003_);
  xor g_62344_(_31294_, _32001_, _32004_);
  and g_62345_(_30740_, _30744_, _32006_);
  not g_62346_(_32006_, _32007_);
  xor g_62347_(_32004_, _32007_, _32008_);
  or g_62348_(_29493_, _30748_, _32009_);
  and g_62349_(_30747_, _32009_, _32010_);
  not g_62350_(_32010_, _32011_);
  xor g_62351_(_32008_, _32011_, _32012_);
  or g_62352_(_31291_, _32012_, _32013_);
  xor g_62353_(_31292_, _32012_, _32014_);
  or g_62354_(_31289_, _32014_, _32015_);
  not g_62355_(_32015_, _32017_);
  xor g_62356_(_31289_, _32014_, _32018_);
  and g_62357_(_31287_, _32018_, _32019_);
  not g_62358_(_32019_, _32020_);
  xor g_62359_(_31286_, _32018_, _32021_);
  or g_62360_(_31284_, _32021_, _32022_);
  xor g_62361_(_31285_, _32021_, _32023_);
  or g_62362_(_31282_, _32023_, _32024_);
  xor g_62363_(_31283_, _32023_, _32025_);
  or g_62364_(_31281_, _32025_, _32026_);
  xor g_62365_(_31280_, _32025_, _32028_);
  or g_62366_(_31277_, _32028_, _32029_);
  not g_62367_(_32029_, _32030_);
  xor g_62368_(_31278_, _32028_, _32031_);
  or g_62369_(_30761_, _32031_, _32032_);
  not g_62370_(_32032_, _32033_);
  xor g_62371_(_30761_, _32031_, _32034_);
  xor g_62372_(_30762_, _32031_, _32035_);
  or g_62373_(_30765_, _32034_, _32036_);
  or g_62374_(_31276_, _32036_, _32037_);
  or g_62375_(_30766_, _32035_, _32039_);
  not g_62376_(_32039_, _32040_);
  or g_62377_(_31275_, _32035_, _32041_);
  and g_62378_(_32039_, _32041_, _32042_);
  and g_62379_(_32037_, _32042_, _32043_);
  not g_62380_(_32043_, _32044_);
  or g_62381_(_31273_, _32044_, _32045_);
  xor g_62382_(_31273_, _32043_, _32046_);
  or g_62383_(_30770_, _32046_, _32047_);
  xor g_62384_(_30771_, _32046_, _32048_);
  xor g_62385_(_30777_, _32048_, _32050_);
  or g_62386_(_30787_, _32050_, _32051_);
  not g_62387_(_32051_, _32052_);
  xor g_62388_(_30788_, _32050_, _32053_);
  and g_62389_(_30792_, _30795_, _32054_);
  not g_62390_(_32054_, _32055_);
  xor g_62391_(_32053_, _32055_, _32056_);
  or g_62392_(_31270_, _32056_, _32057_);
  xor g_62393_(_31271_, _32056_, _32058_);
  or g_62394_(_31267_, _32058_, _32059_);
  not g_62395_(_32059_, _32061_);
  xor g_62396_(_31269_, _32058_, _32062_);
  and g_62397_(_30802_, _30805_, _32063_);
  and g_62398_(_32062_, _32063_, _32064_);
  not g_62399_(_32064_, _32065_);
  or g_62400_(_30805_, _32062_, _32066_);
  not g_62401_(_32066_, _32067_);
  or g_62402_(_30802_, _32062_, _32068_);
  not g_62403_(_32068_, _32069_);
  and g_62404_(_32066_, _32068_, _32070_);
  not g_62405_(_32070_, _32072_);
  and g_62406_(_32065_, _32070_, _32073_);
  or g_62407_(_32064_, _32072_, _32074_);
  and g_62408_(_30809_, _30811_, _32075_);
  or g_62409_(_32074_, _32075_, _32076_);
  xor g_62410_(_32073_, _32075_, _32077_);
  not g_62411_(_32077_, _32078_);
  and g_62412_(_30820_, _30822_, _32079_);
  xor g_62413_(_32078_, _32079_, _32080_);
  or g_62414_(_30824_, _32080_, _32081_);
  not g_62415_(_32081_, _32083_);
  xor g_62416_(_30824_, _32080_, _32084_);
  not g_62417_(_32084_, _32085_);
  and g_62418_(_30827_, _32084_, _32086_);
  or g_62419_(_30826_, _32085_, _32087_);
  xor g_62420_(_30826_, _32084_, _32088_);
  or g_62421_(_30830_, _32088_, _32089_);
  xor g_62422_(_30831_, _32088_, _32090_);
  or g_62423_(_30832_, _30833_, _32091_);
  or g_62424_(_32090_, _32091_, _32092_);
  not g_62425_(_32092_, _32094_);
  and g_62426_(_32090_, _32091_, _32095_);
  xor g_62427_(_32090_, _32091_, _32096_);
  or g_62428_(_32094_, _32095_, _32097_);
  or g_62429_(_31266_, _32097_, _32098_);
  xor g_62430_(_31266_, _32096_, _32099_);
  not g_62431_(_32099_, _32100_);
  or g_62432_(_30838_, _32099_, _32101_);
  xor g_62433_(_30838_, _32100_, _32102_);
  and g_62434_(_30841_, _30844_, _32103_);
  not g_62435_(_32103_, _32105_);
  xor g_62436_(_32102_, _32105_, _32106_);
  xor g_62437_(_31265_, _32106_, _32107_);
  not g_62438_(_32107_, _32108_);
  or g_62439_(_31264_, _32108_, _32109_);
  xor g_62440_(_31264_, _32107_, _32110_);
  or g_62441_(_31263_, _32110_, _32111_);
  xor g_62442_(_31262_, _32110_, _32112_);
  or g_62443_(_30857_, _30861_, _32113_);
  xor g_62444_(_32112_, _32113_, _32114_);
  xor g_62445_(_31261_, _32114_, _32116_);
  and g_62446_(_30875_, _32116_, _32117_);
  xor g_62447_(_30876_, _32116_, _32118_);
  or g_62448_(_31260_, _32118_, _32119_);
  not g_62449_(_32119_, _32120_);
  xor g_62450_(_31260_, _32118_, _32121_);
  not g_62451_(_32121_, _32122_);
  or g_62452_(_31259_, _32122_, _32123_);
  xor g_62453_(_31259_, _32121_, _32124_);
  or g_62454_(_30887_, _32124_, _32125_);
  not g_62455_(_32125_, _32127_);
  and g_62456_(_30887_, _32124_, _32128_);
  xor g_62457_(_30887_, _32124_, _32129_);
  or g_62458_(_32127_, _32128_, _32130_);
  or g_62459_(_31258_, _32130_, _32131_);
  xor g_62460_(_31258_, _32129_, _32132_);
  not g_62461_(_32132_, _32133_);
  or g_62462_(_31256_, _32132_, _32134_);
  xor g_62463_(_31256_, _32132_, _32135_);
  xor g_62464_(_31256_, _32133_, _32136_);
  or g_62465_(_30892_, _32136_, _32138_);
  xor g_62466_(_30892_, _32135_, _32139_);
  or g_62467_(_30897_, _32139_, _32140_);
  xor g_62468_(_30897_, _32139_, _32141_);
  xor g_62469_(_30896_, _32139_, _32142_);
  and g_62470_(_30900_, _30903_, _32143_);
  xor g_62471_(_32141_, _32143_, _32144_);
  not g_62472_(_32144_, _32145_);
  and g_62473_(_30909_, _32145_, _32146_);
  xor g_62474_(_30908_, _32144_, _32147_);
  xor g_62475_(_30909_, _32144_, _32149_);
  and g_62476_(_30912_, _30915_, _32150_);
  xor g_62477_(_32147_, _32150_, _32151_);
  or g_62478_(_31255_, _32151_, _32152_);
  not g_62479_(_32152_, _32153_);
  xor g_62480_(_31255_, _32151_, _32154_);
  and g_62481_(_31254_, _32154_, _32155_);
  not g_62482_(_32155_, _32156_);
  xor g_62483_(_31253_, _32154_, _32157_);
  or g_62484_(_31252_, _32157_, _32158_);
  xor g_62485_(_31251_, _32157_, _32160_);
  not g_62486_(_32160_, _32161_);
  or g_62487_(_29638_, _30922_, _32162_);
  or g_62488_(_29641_, _30926_, _32163_);
  and g_62489_(_32162_, _32163_, _32164_);
  xor g_62490_(_32161_, _32164_, _32165_);
  xor g_62491_(_32160_, _32164_, _32166_);
  or g_62492_(_31250_, _32165_, _32167_);
  xor g_62493_(_31250_, _32166_, _32168_);
  not g_62494_(_32168_, _32169_);
  and g_62495_(_30930_, _30933_, _32171_);
  xor g_62496_(_32169_, _32171_, _32172_);
  or g_62497_(_31249_, _32172_, _32173_);
  not g_62498_(_32173_, _32174_);
  xor g_62499_(_31249_, _32172_, _32175_);
  not g_62500_(_32175_, _32176_);
  or g_62501_(_31248_, _32176_, _32177_);
  xor g_62502_(_31248_, _32175_, _32178_);
  or g_62503_(_31247_, _32178_, _32179_);
  not g_62504_(_32179_, _32180_);
  and g_62505_(_31247_, _32178_, _32182_);
  xor g_62506_(_31247_, _32178_, _32183_);
  or g_62507_(_32180_, _32182_, _32184_);
  or g_62508_(_31245_, _32184_, _32185_);
  xor g_62509_(_31245_, _32183_, _32186_);
  not g_62510_(_32186_, _32187_);
  or g_62511_(_31244_, _32186_, _32188_);
  xor g_62512_(_31244_, _32187_, _32189_);
  not g_62513_(_32189_, _32190_);
  or g_62514_(_29665_, _30941_, _32191_);
  and g_62515_(_30948_, _32191_, _32193_);
  and g_62516_(_30946_, _32193_, _32194_);
  xor g_62517_(_32189_, _32194_, _32195_);
  xor g_62518_(_32190_, _32194_, _32196_);
  or g_62519_(_29676_, _30949_, _32197_);
  or g_62520_(_32196_, _32197_, _32198_);
  xor g_62521_(_32195_, _32197_, _32199_);
  not g_62522_(_32199_, _32200_);
  or g_62523_(_31243_, _32199_, _32201_);
  xor g_62524_(_31243_, _32200_, _32202_);
  or g_62525_(_30956_, _32202_, _32204_);
  not g_62526_(_32204_, _32205_);
  xor g_62527_(_30956_, _32202_, _32206_);
  not g_62528_(_32206_, _32207_);
  and g_62529_(_30959_, _32206_, _32208_);
  or g_62530_(_30958_, _32207_, _32209_);
  xor g_62531_(_30958_, _32206_, _32210_);
  or g_62532_(_30969_, _32210_, _32211_);
  xor g_62533_(_30970_, _32210_, _32212_);
  or g_62534_(_30967_, _32212_, _32213_);
  xor g_62535_(_30968_, _32212_, _32215_);
  or g_62536_(_29696_, _30975_, _32216_);
  or g_62537_(_32215_, _32216_, _32217_);
  not g_62538_(_32217_, _32218_);
  and g_62539_(_32215_, _32216_, _32219_);
  xor g_62540_(_32215_, _32216_, _32220_);
  or g_62541_(_32218_, _32219_, _32221_);
  or g_62542_(_31242_, _32221_, _32222_);
  xor g_62543_(_31242_, _32220_, _32223_);
  not g_62544_(_32223_, _32224_);
  and g_62545_(_30977_, _30984_, _32226_);
  xor g_62546_(_32224_, _32226_, _32227_);
  not g_62547_(_32227_, _32228_);
  and g_62548_(_30979_, _30988_, _32229_);
  xor g_62549_(_32228_, _32229_, _32230_);
  or g_62550_(_31241_, _32230_, _32231_);
  not g_62551_(_32231_, _32232_);
  xor g_62552_(_31241_, _32230_, _32233_);
  not g_62553_(_32233_, _32234_);
  or g_62554_(_31240_, _32234_, _32235_);
  not g_62555_(_32235_, _32237_);
  xor g_62556_(_31240_, _32233_, _32238_);
  or g_62557_(_31239_, _32238_, _32239_);
  not g_62558_(_32239_, _32240_);
  xor g_62559_(_31238_, _32238_, _32241_);
  or g_62560_(_31236_, _32241_, _32242_);
  xor g_62561_(_31237_, _32241_, _32243_);
  not g_62562_(_32243_, _32244_);
  and g_62563_(_30996_, _32243_, _32245_);
  and g_62564_(_31000_, _32245_, _32246_);
  not g_62565_(_32246_, _32248_);
  and g_62566_(_30999_, _32244_, _32249_);
  or g_62567_(_31000_, _32243_, _32250_);
  or g_62568_(_30996_, _32243_, _32251_);
  not g_62569_(_32251_, _32252_);
  and g_62570_(_32250_, _32251_, _32253_);
  or g_62571_(_32249_, _32252_, _32254_);
  and g_62572_(_32248_, _32253_, _32255_);
  or g_62573_(_32246_, _32254_, _32256_);
  and g_62574_(_31234_, _32255_, _32257_);
  or g_62575_(_31233_, _32256_, _32259_);
  xor g_62576_(_31234_, _32255_, _32260_);
  xor g_62577_(_31233_, _32255_, _32261_);
  and g_62578_(_31232_, _32260_, _32262_);
  or g_62579_(_31231_, _32261_, _32263_);
  xor g_62580_(_31231_, _32260_, _32264_);
  or g_62581_(_31228_, _32264_, _32265_);
  xor g_62582_(_31228_, _32264_, _32266_);
  xor g_62583_(_31229_, _32264_, _32267_);
  or g_62584_(_29746_, _31002_, _32268_);
  or g_62585_(_32267_, _32268_, _32270_);
  xor g_62586_(_32266_, _32268_, _32271_);
  not g_62587_(_32271_, _32272_);
  or g_62588_(_31007_, _31009_, _32273_);
  not g_62589_(_32273_, _32274_);
  and g_62590_(_32272_, _32273_, _32275_);
  or g_62591_(_32271_, _32274_, _32276_);
  xor g_62592_(_32271_, _32273_, _32277_);
  or g_62593_(_31227_, _32277_, _32278_);
  not g_62594_(_32278_, _32279_);
  xor g_62595_(_31227_, _32277_, _32281_);
  not g_62596_(_32281_, _32282_);
  or g_62597_(_31226_, _32282_, _32283_);
  xor g_62598_(_31226_, _32281_, _32284_);
  not g_62599_(_32284_, _32285_);
  or g_62600_(_31019_, _32284_, _32286_);
  xor g_62601_(_31019_, _32285_, _32287_);
  or g_62602_(_31023_, _32287_, _32288_);
  xor g_62603_(_31023_, _32287_, _32289_);
  xor g_62604_(_31024_, _32287_, _32290_);
  or g_62605_(_31028_, _32290_, _32292_);
  xor g_62606_(_31028_, _32290_, _32293_);
  xor g_62607_(_31028_, _32289_, _32294_);
  and g_62608_(_29773_, _31032_, _32295_);
  or g_62609_(_29772_, _31033_, _32296_);
  and g_62610_(_32293_, _32295_, _32297_);
  or g_62611_(_32294_, _32296_, _32298_);
  and g_62612_(_31031_, _32293_, _32299_);
  or g_62613_(_31030_, _32294_, _32300_);
  and g_62614_(_32298_, _32300_, _32301_);
  or g_62615_(_32297_, _32299_, _32303_);
  and g_62616_(_31030_, _32294_, _32304_);
  and g_62617_(_32296_, _32304_, _32305_);
  or g_62618_(_32303_, _32305_, _32306_);
  or g_62619_(_31041_, _32306_, _32307_);
  not g_62620_(_32307_, _32308_);
  or g_62621_(_29776_, _31033_, _32309_);
  not g_62622_(_32309_, _32310_);
  or g_62623_(_32306_, _32309_, _32311_);
  xor g_62624_(_32306_, _32309_, _32312_);
  xor g_62625_(_32306_, _32310_, _32314_);
  and g_62626_(_31041_, _32314_, _32315_);
  or g_62627_(_31042_, _32312_, _32316_);
  and g_62628_(_32307_, _32316_, _32317_);
  or g_62629_(_32308_, _32315_, _32318_);
  and g_62630_(_31037_, _32317_, _32319_);
  or g_62631_(_31036_, _32318_, _32320_);
  xor g_62632_(_31037_, _32317_, _32321_);
  xor g_62633_(_31036_, _32317_, _32322_);
  and g_62634_(_31054_, _32321_, _32323_);
  or g_62635_(_31055_, _32322_, _32325_);
  or g_62636_(_31046_, _32318_, _32326_);
  not g_62637_(_32326_, _32327_);
  or g_62638_(_32323_, _32327_, _32328_);
  and g_62639_(_31046_, _32322_, _32329_);
  and g_62640_(_31055_, _32329_, _32330_);
  or g_62641_(_32328_, _32330_, _32331_);
  or g_62642_(_31053_, _32331_, _32332_);
  xor g_62643_(_31053_, _32331_, _32333_);
  xor g_62644_(_31052_, _32331_, _32334_);
  and g_62645_(_31063_, _32333_, _32336_);
  or g_62646_(_31062_, _32334_, _32337_);
  or g_62647_(_31058_, _32334_, _32338_);
  not g_62648_(_32338_, _32339_);
  xor g_62649_(_31058_, _32333_, _32340_);
  or g_62650_(_31074_, _32340_, _32341_);
  not g_62651_(_32341_, _32342_);
  xor g_62652_(_31073_, _32340_, _32343_);
  and g_62653_(_31062_, _32343_, _32344_);
  or g_62654_(_32336_, _32344_, _32345_);
  or g_62655_(_31067_, _32345_, _32347_);
  not g_62656_(_32347_, _32348_);
  xor g_62657_(_31066_, _32345_, _32349_);
  not g_62658_(_32349_, _32350_);
  or g_62659_(_31225_, _32349_, _32351_);
  xor g_62660_(_31225_, _32350_, _32352_);
  not g_62661_(_32352_, _32353_);
  or g_62662_(_31223_, _32352_, _32354_);
  xor g_62663_(_31223_, _32352_, _32355_);
  xor g_62664_(_31223_, _32353_, _32356_);
  and g_62665_(_31086_, _31089_, _32358_);
  xor g_62666_(_32356_, _32358_, _32359_);
  not g_62667_(_32359_, _32360_);
  and g_62668_(_31092_, _32359_, _32361_);
  or g_62669_(_31091_, _32360_, _32362_);
  xor g_62670_(_31091_, _32359_, _32363_);
  not g_62671_(_32363_, _32364_);
  or g_62672_(_31222_, _32363_, _32365_);
  xor g_62673_(_31222_, _32363_, _32366_);
  xor g_62674_(_31222_, _32364_, _32367_);
  or g_62675_(_31221_, _32367_, _32369_);
  not g_62676_(_32369_, _32370_);
  xor g_62677_(_31221_, _32366_, _32371_);
  or g_62678_(_31100_, _32371_, _32372_);
  xor g_62679_(_31099_, _32371_, _32373_);
  or g_62680_(_31220_, _32373_, _32374_);
  not g_62681_(_32374_, _32375_);
  or g_62682_(_29837_, _31101_, _32376_);
  or g_62683_(_32371_, _32376_, _32377_);
  not g_62684_(_32377_, _32378_);
  and g_62685_(_32373_, _32376_, _32380_);
  or g_62686_(_32378_, _32380_, _32381_);
  and g_62687_(_31220_, _32381_, _32382_);
  or g_62688_(_32375_, _32382_, _32383_);
  not g_62689_(_32383_, _32384_);
  and g_62690_(_31107_, _31109_, _32385_);
  xor g_62691_(_32384_, _32385_, _32386_);
  or g_62692_(_31114_, _32386_, _32387_);
  xor g_62693_(_31114_, _32386_, _32388_);
  not g_62694_(_32388_, _32389_);
  and g_62695_(_31117_, _31121_, _32391_);
  xor g_62696_(_32388_, _32391_, _32392_);
  or g_62697_(_29863_, _31122_, _32393_);
  and g_62698_(_31124_, _32393_, _32394_);
  xor g_62699_(_32392_, _32394_, _32395_);
  not g_62700_(_32395_, _32396_);
  or g_62701_(_31219_, _32396_, _32397_);
  xor g_62702_(_31219_, _32395_, _32398_);
  not g_62703_(_32398_, _32399_);
  or g_62704_(_31218_, _32398_, _32400_);
  xor g_62705_(_31218_, _32399_, _32402_);
  not g_62706_(_32402_, _32403_);
  or g_62707_(_31217_, _32402_, _32404_);
  xor g_62708_(_31217_, _32403_, _32405_);
  or g_62709_(_31135_, _32405_, _32406_);
  not g_62710_(_32406_, _32407_);
  xor g_62711_(_31136_, _32405_, _32408_);
  not g_62712_(_32408_, _32409_);
  or g_62713_(_29879_, _31139_, _32410_);
  and g_62714_(_31131_, _32410_, _32411_);
  xor g_62715_(_32409_, _32411_, _32413_);
  or g_62716_(_31215_, _32413_, _32414_);
  not g_62717_(_32414_, _32415_);
  xor g_62718_(_31215_, _32413_, _32416_);
  not g_62719_(_32416_, _32417_);
  and g_62720_(_31143_, _31146_, _32418_);
  xor g_62721_(_32416_, _32418_, _32419_);
  and g_62722_(_31149_, _32419_, _32420_);
  or g_62723_(_31149_, _32419_, _32421_);
  not g_62724_(_32421_, _32422_);
  or g_62725_(_32420_, _32422_, _32424_);
  not g_62726_(_32424_, _32425_);
  and g_62727_(_31151_, _31155_, _32426_);
  or g_62728_(_32424_, _32426_, _32427_);
  xor g_62729_(_32424_, _32426_, _32428_);
  xor g_62730_(_32425_, _32426_, _32429_);
  or g_62731_(_31157_, _32429_, _32430_);
  xor g_62732_(_31157_, _32428_, _32431_);
  not g_62733_(_32431_, _32432_);
  or g_62734_(_31160_, _32431_, _32433_);
  xor g_62735_(_31160_, _32432_, _32435_);
  and g_62736_(_29894_, _31161_, _32436_);
  not g_62737_(_32436_, _32437_);
  or g_62738_(_32435_, _32437_, _32438_);
  xor g_62739_(_32435_, _32436_, _32439_);
  or g_62740_(_31212_, _32439_, _32440_);
  xor g_62741_(_31212_, _32439_, _32441_);
  xor g_62742_(_31214_, _32439_, _32442_);
  or g_62743_(_31211_, _32442_, _32443_);
  not g_62744_(_32443_, _32444_);
  xor g_62745_(_31211_, _32441_, _32446_);
  or g_62746_(_31209_, _32446_, _32447_);
  xor g_62747_(_31210_, _32446_, _32448_);
  not g_62748_(_32448_, _32449_);
  or g_62749_(_31208_, _32448_, _32450_);
  xor g_62750_(_31208_, _32449_, _32451_);
  not g_62751_(_32451_, _32452_);
  or g_62752_(_31207_, _32451_, _32453_);
  xor g_62753_(_31207_, _32451_, _32454_);
  xor g_62754_(_31207_, _32452_, _32455_);
  or g_62755_(_31174_, _32455_, _32457_);
  xor g_62756_(_31174_, _32454_, _32458_);
  or g_62757_(_31173_, _32458_, _32459_);
  not g_62758_(_32459_, _32460_);
  and g_62759_(_31173_, _32458_, _32461_);
  or g_62760_(_32460_, _32461_, _32462_);
  and g_62761_(_31179_, _31183_, _32463_);
  or g_62762_(_32462_, _32463_, _32464_);
  xor g_62763_(_32462_, _32463_, _32465_);
  not g_62764_(_32465_, _32466_);
  or g_62765_(_29931_, _31188_, _32468_);
  and g_62766_(_31185_, _32468_, _32469_);
  xor g_62767_(_32465_, _32469_, _32470_);
  xor g_62768_(_32466_, _32469_, _32471_);
  or g_62769_(_31206_, _32470_, _32472_);
  xor g_62770_(_31206_, _32470_, _32473_);
  xor g_62771_(_31206_, _32471_, _32474_);
  and g_62772_(_31197_, _32473_, _32475_);
  or g_62773_(_31198_, _32474_, _32476_);
  and g_62774_(_31193_, _32473_, _32477_);
  or g_62775_(_31194_, _32474_, _32479_);
  or g_62776_(_32475_, _32477_, _32480_);
  and g_62777_(_31194_, _32474_, _32481_);
  and g_62778_(_31198_, _32481_, _32482_);
  or g_62779_(_32480_, _32482_, _32483_);
  or g_62780_(_31204_, _32483_, _32484_);
  xor g_62781_(_31205_, _32483_, _32485_);
  or g_62782_(_31203_, _32485_, _32486_);
  xor g_62783_(_31203_, _32485_, out[644]);
  or g_62784_(_32466_, _32468_, _32487_);
  not g_62785_(_32487_, _32489_);
  and g_62786_(_31186_, _32465_, _32490_);
  and g_62787_(_32430_, _32433_, _32491_);
  or g_62788_(_32408_, _32410_, _32492_);
  not g_62789_(_32492_, _32493_);
  or g_62790_(_32392_, _32393_, _32494_);
  or g_62791_(_31124_, _32392_, _32495_);
  not g_62792_(_32495_, _32496_);
  or g_62793_(_31121_, _32389_, _32497_);
  and g_62794_(_31118_, _32388_, _32498_);
  or g_62795_(_31117_, _32389_, _32500_);
  and g_62796_(_31110_, _32384_, _32501_);
  or g_62797_(_31089_, _32356_, _32502_);
  not g_62798_(_32502_, _32503_);
  and g_62799_(_32332_, _32338_, _32504_);
  and g_62800_(_32265_, _32270_, _32505_);
  or g_62801_(_30988_, _32227_, _32506_);
  not g_62802_(_32506_, _32507_);
  or g_62803_(_30979_, _32227_, _32508_);
  not g_62804_(_32508_, _32509_);
  or g_62805_(_30984_, _32223_, _32511_);
  or g_62806_(_30977_, _32223_, _32512_);
  not g_62807_(_32512_, _32513_);
  and g_62808_(_30947_, _32190_, _32514_);
  or g_62809_(_30948_, _32189_, _32515_);
  not g_62810_(_32515_, _32516_);
  or g_62811_(_30933_, _32168_, _32517_);
  or g_62812_(_30930_, _32168_, _32518_);
  or g_62813_(_32160_, _32163_, _32519_);
  not g_62814_(_32519_, _32520_);
  or g_62815_(_32160_, _32162_, _32522_);
  not g_62816_(_32522_, _32523_);
  or g_62817_(_30915_, _32149_, _32524_);
  not g_62818_(_32524_, _32525_);
  or g_62819_(_30912_, _32144_, _32526_);
  not g_62820_(_32526_, _32527_);
  or g_62821_(_30900_, _32142_, _32528_);
  and g_62822_(_32140_, _32528_, _32529_);
  or g_62823_(_30878_, _32114_, _32530_);
  or g_62824_(_30865_, _32114_, _32531_);
  not g_62825_(_32531_, _32533_);
  or g_62826_(_30863_, _32112_, _32534_);
  or g_62827_(_30858_, _32112_, _32535_);
  not g_62828_(_32535_, _32536_);
  or g_62829_(_30850_, _32106_, _32537_);
  or g_62830_(_30847_, _32106_, _32538_);
  not g_62831_(_32538_, _32539_);
  or g_62832_(_30844_, _32102_, _32540_);
  or g_62833_(_30841_, _32102_, _32541_);
  or g_62834_(_30822_, _32077_, _32542_);
  not g_62835_(_32542_, _32544_);
  or g_62836_(_30795_, _32053_, _32545_);
  or g_62837_(_30773_, _32048_, _32546_);
  or g_62838_(_30775_, _32048_, _32547_);
  or g_62839_(_32008_, _32009_, _32548_);
  not g_62840_(_32548_, _32549_);
  or g_62841_(_30747_, _32008_, _32550_);
  or g_62842_(_30744_, _32004_, _32551_);
  or g_62843_(_31992_, _31993_, _32552_);
  not g_62844_(_32552_, _32553_);
  and g_62845_(_30732_, _31991_, _32555_);
  or g_62846_(_30733_, _31992_, _32556_);
  and g_62847_(_31984_, _31986_, _32557_);
  and g_62848_(_30704_, _31951_, _32558_);
  or g_62849_(_30705_, _31952_, _32559_);
  or g_62850_(_30638_, _31879_, _32560_);
  not g_62851_(_32560_, _32561_);
  or g_62852_(_30630_, _31878_, _32562_);
  not g_62853_(_32562_, _32563_);
  or g_62854_(_30615_, _31863_, _32564_);
  or g_62855_(_30611_, _31863_, _32566_);
  or g_62856_(_30599_, _31855_, _32567_);
  not g_62857_(_32567_, _32568_);
  or g_62858_(_30596_, _31855_, _32569_);
  not g_62859_(_32569_, _32570_);
  or g_62860_(_31849_, _31850_, _32571_);
  not g_62861_(_32571_, _32572_);
  or g_62862_(_30591_, _31849_, _32573_);
  or g_62863_(_31828_, _31832_, _32574_);
  not g_62864_(_32574_, _32575_);
  or g_62865_(_31828_, _31831_, _32577_);
  not g_62866_(_32577_, _32578_);
  or g_62867_(_30557_, _31811_, _32579_);
  not g_62868_(_32579_, _32580_);
  or g_62869_(_30551_, _31811_, _32581_);
  not g_62870_(_32581_, _32582_);
  and g_62871_(_31806_, _31810_, _32583_);
  not g_62872_(_32583_, _32584_);
  or g_62873_(_29280_, _30535_, _32585_);
  or g_62874_(_31801_, _32585_, _32586_);
  not g_62875_(_32586_, _32588_);
  and g_62876_(_30497_, _31753_, _32589_);
  not g_62877_(_32589_, _32590_);
  or g_62878_(_30494_, _31751_, _32591_);
  and g_62879_(_31722_, _31725_, _32592_);
  or g_62880_(_31715_, _31717_, _32593_);
  or g_62881_(_30465_, _31715_, _32594_);
  and g_62882_(_31700_, _31705_, _32595_);
  or g_62883_(_30440_, _31698_, _32596_);
  and g_62884_(_31702_, _32596_, _32597_);
  or g_62885_(_31672_, _31673_, _32599_);
  or g_62886_(_30406_, _31672_, _32600_);
  or g_62887_(_31655_, _31657_, _32601_);
  not g_62888_(_32601_, _32602_);
  or g_62889_(_30392_, _31655_, _32603_);
  not g_62890_(_32603_, _32604_);
  and g_62891_(_30384_, _31649_, _32605_);
  not g_62892_(_32605_, _32606_);
  and g_62893_(_30374_, _31635_, _32607_);
  not g_62894_(_32607_, _32608_);
  and g_62895_(_29153_, _32607_, _32610_);
  not g_62896_(_32610_, _32611_);
  or g_62897_(_29151_, _32608_, _32612_);
  and g_62898_(_31638_, _31643_, _32613_);
  or g_62899_(_31637_, _31641_, _32614_);
  and g_62900_(_31628_, _31632_, _32615_);
  and g_62901_(_30347_, _31603_, _32616_);
  not g_62902_(_32616_, _32617_);
  or g_62903_(_30340_, _31601_, _32618_);
  not g_62904_(_32618_, _32619_);
  or g_62905_(_30337_, _31601_, _32621_);
  not g_62906_(_32621_, _32622_);
  or g_62907_(_30329_, _31593_, _32623_);
  or g_62908_(_29104_, _32623_, _32624_);
  or g_62909_(_29101_, _30329_, _32625_);
  or g_62910_(_31600_, _32625_, _32626_);
  and g_62911_(_31568_, _31571_, _32627_);
  or g_62912_(_30288_, _31548_, _32628_);
  or g_62913_(_30069_, _32628_, _32629_);
  or g_62914_(_29075_, _32628_, _32630_);
  not g_62915_(_32630_, _32632_);
  and g_62916_(_31529_, _31530_, _32633_);
  or g_62917_(_30239_, _31487_, _32634_);
  not g_62918_(_32634_, _32635_);
  and g_62919_(_30229_, _31476_, _32636_);
  or g_62920_(_31478_, _32636_, _32637_);
  and g_62921_(_30216_, _31463_, _32638_);
  or g_62922_(_31464_, _32638_, _32639_);
  or g_62923_(_30208_, _31461_, _32640_);
  or g_62924_(_27716_, _30193_, _32641_);
  or g_62925_(_28995_, _32641_, _32643_);
  or g_62926_(_31458_, _32643_, _32644_);
  or g_62927_(_30173_, _31424_, _32645_);
  or g_62928_(_31421_, _31426_, _32646_);
  and g_62929_(_31410_, _31414_, _32647_);
  and g_62930_(_31416_, _32647_, _32648_);
  and g_62931_(_31423_, _32648_, _32649_);
  and g_62932_(_32646_, _32649_, _32650_);
  and g_62933_(_32645_, _32650_, _32651_);
  and g_62934_(_31429_, _32651_, _32652_);
  and g_62935_(_31435_, _32652_, _32654_);
  and g_62936_(_31438_, _32654_, _32655_);
  and g_62937_(_31441_, _32655_, _32656_);
  and g_62938_(_31443_, _32656_, _32657_);
  and g_62939_(_31447_, _32657_, _32658_);
  and g_62940_(_31450_, _32658_, _32659_);
  and g_62941_(_31453_, _32659_, _32660_);
  or g_62942_(_32644_, _32660_, _32661_);
  and g_62943_(_31458_, _32643_, _32662_);
  or g_62944_(_27720_, _28995_, _32663_);
  or g_62945_(_30199_, _32663_, _32665_);
  and g_62946_(_30206_, _32665_, _32666_);
  or g_62947_(_32662_, _32666_, _32667_);
  and g_62948_(_31457_, _32660_, _32668_);
  and g_62949_(_32644_, _32668_, _32669_);
  and g_62950_(_32667_, _32669_, _32670_);
  not g_62951_(_32670_, _32671_);
  and g_62952_(_32661_, _32671_, _32672_);
  xor g_62953_(_32640_, _32672_, _32673_);
  xor g_62954_(_31472_, _32673_, _32674_);
  xor g_62955_(_32639_, _32674_, _32676_);
  xor g_62956_(_32637_, _32676_, _32677_);
  or g_62957_(_30236_, _31486_, _32678_);
  and g_62958_(_31481_, _32678_, _32679_);
  xor g_62959_(_32677_, _32679_, _32680_);
  not g_62960_(_32680_, _32681_);
  and g_62961_(_32635_, _32680_, _32682_);
  or g_62962_(_32634_, _32681_, _32683_);
  xor g_62963_(_32634_, _32680_, _32684_);
  not g_62964_(_32684_, _32685_);
  or g_62965_(_31493_, _32684_, _32687_);
  xor g_62966_(_31493_, _32684_, _32688_);
  xor g_62967_(_31493_, _32685_, _32689_);
  and g_62968_(_31496_, _32688_, _32690_);
  or g_62969_(_31495_, _32689_, _32691_);
  xor g_62970_(_31495_, _32688_, _32692_);
  and g_62971_(_31500_, _32692_, _32693_);
  not g_62972_(_32693_, _32694_);
  or g_62973_(_31500_, _32689_, _32695_);
  and g_62974_(_32694_, _32695_, _32696_);
  xor g_62975_(_31503_, _32696_, _32698_);
  or g_62976_(_31509_, _32698_, _32699_);
  not g_62977_(_32699_, _32700_);
  or g_62978_(_31505_, _32698_, _32701_);
  xor g_62979_(_31505_, _32698_, _32702_);
  xor g_62980_(_31506_, _32698_, _32703_);
  and g_62981_(_31509_, _32703_, _32704_);
  or g_62982_(_31511_, _32702_, _32705_);
  or g_62983_(_32700_, _32704_, _32706_);
  and g_62984_(_31515_, _32706_, _32707_);
  and g_62985_(_31514_, _32705_, _32709_);
  or g_62986_(_31515_, _32704_, _32710_);
  and g_62987_(_32699_, _32709_, _32711_);
  or g_62988_(_32707_, _32711_, _32712_);
  or g_62989_(_31518_, _31520_, _32713_);
  and g_62990_(_31517_, _32713_, _32714_);
  not g_62991_(_32714_, _32715_);
  or g_62992_(_32712_, _32714_, _32716_);
  not g_62993_(_32716_, _32717_);
  and g_62994_(_32712_, _32714_, _32718_);
  xor g_62995_(_32712_, _32715_, _32720_);
  or g_62996_(_30262_, _31519_, _32721_);
  and g_62997_(_31525_, _32721_, _32722_);
  and g_62998_(_32720_, _32722_, _32723_);
  not g_62999_(_32723_, _32724_);
  or g_63000_(_32718_, _32722_, _32725_);
  or g_63001_(_32717_, _32725_, _32726_);
  and g_63002_(_32724_, _32726_, _32727_);
  not g_63003_(_32727_, _32728_);
  or g_63004_(_32633_, _32728_, _32729_);
  xor g_63005_(_32633_, _32728_, _32731_);
  xor g_63006_(_32633_, _32727_, _32732_);
  or g_63007_(_31535_, _32732_, _32733_);
  and g_63008_(_31535_, _32732_, _32734_);
  or g_63009_(_31534_, _32731_, _32735_);
  xor g_63010_(_31534_, _32732_, _32736_);
  and g_63011_(_31540_, _32736_, _32737_);
  and g_63012_(_31541_, _32735_, _32738_);
  or g_63013_(_31540_, _32734_, _32739_);
  and g_63014_(_32733_, _32738_, _32740_);
  or g_63015_(_32737_, _32740_, _32742_);
  and g_63016_(_31546_, _32742_, _32743_);
  or g_63017_(_31546_, _32742_, _32744_);
  xor g_63018_(_31546_, _32742_, _32745_);
  xor g_63019_(_31547_, _32742_, _32746_);
  xor g_63020_(_31550_, _32745_, _32747_);
  and g_63021_(_31552_, _32747_, _32748_);
  or g_63022_(_31552_, _32746_, _32749_);
  not g_63023_(_32749_, _32750_);
  or g_63024_(_32748_, _32750_, _32751_);
  xor g_63025_(_32632_, _32751_, _32753_);
  and g_63026_(_32629_, _32753_, _32754_);
  or g_63027_(_32629_, _32753_, _32755_);
  xor g_63028_(_32629_, _32753_, _32756_);
  and g_63029_(_30295_, _31556_, _32757_);
  or g_63030_(_31557_, _32757_, _32758_);
  xor g_63031_(_32756_, _32758_, _32759_);
  or g_63032_(_31563_, _32759_, _32760_);
  xor g_63033_(_31563_, _32759_, _32761_);
  xor g_63034_(_31564_, _32759_, _32762_);
  or g_63035_(_32627_, _32762_, _32764_);
  xor g_63036_(_32627_, _32761_, _32765_);
  and g_63037_(_31573_, _32765_, _32766_);
  or g_63038_(_31573_, _32765_, _32767_);
  xor g_63039_(_31574_, _32765_, _32768_);
  xor g_63040_(_31580_, _32768_, _32769_);
  or g_63041_(_31581_, _32769_, _32770_);
  and g_63042_(_31581_, _32769_, _32771_);
  or g_63043_(_31588_, _32771_, _32772_);
  not g_63044_(_32772_, _32773_);
  and g_63045_(_32770_, _32773_, _32775_);
  not g_63046_(_32775_, _32776_);
  xor g_63047_(_31582_, _32769_, _32777_);
  and g_63048_(_31588_, _32777_, _32778_);
  not g_63049_(_32778_, _32779_);
  and g_63050_(_31591_, _32779_, _32780_);
  or g_63051_(_31592_, _32778_, _32781_);
  and g_63052_(_32776_, _32780_, _32782_);
  or g_63053_(_32775_, _32781_, _32783_);
  or g_63054_(_31591_, _32777_, _32784_);
  and g_63055_(_32783_, _32784_, _32786_);
  xor g_63056_(_31595_, _32786_, _32787_);
  or g_63057_(_31599_, _32787_, _32788_);
  and g_63058_(_31599_, _32787_, _32789_);
  xor g_63059_(_31599_, _32787_, _32790_);
  xor g_63060_(_32626_, _32790_, _32791_);
  or g_63061_(_32624_, _32791_, _32792_);
  and g_63062_(_32624_, _32791_, _32793_);
  xor g_63063_(_32624_, _32791_, _32794_);
  xor g_63064_(_32622_, _32794_, _32795_);
  xor g_63065_(_32621_, _32794_, _32797_);
  and g_63066_(_32619_, _32795_, _32798_);
  or g_63067_(_32618_, _32797_, _32799_);
  and g_63068_(_32618_, _32797_, _32800_);
  not g_63069_(_32800_, _32801_);
  and g_63070_(_32799_, _32801_, _32802_);
  and g_63071_(_32616_, _32802_, _32803_);
  not g_63072_(_32803_, _32804_);
  or g_63073_(_30342_, _31602_, _32805_);
  not g_63074_(_32805_, _32806_);
  or g_63075_(_32802_, _32805_, _32808_);
  not g_63076_(_32808_, _32809_);
  and g_63077_(_32799_, _32805_, _32810_);
  or g_63078_(_32798_, _32806_, _32811_);
  and g_63079_(_32801_, _32810_, _32812_);
  or g_63080_(_32800_, _32811_, _32813_);
  and g_63081_(_32617_, _32813_, _32814_);
  or g_63082_(_32616_, _32812_, _32815_);
  and g_63083_(_32808_, _32814_, _32816_);
  or g_63084_(_32809_, _32815_, _32817_);
  and g_63085_(_32804_, _32817_, _32819_);
  or g_63086_(_32803_, _32816_, _32820_);
  or g_63087_(_31610_, _32820_, _32821_);
  and g_63088_(_31606_, _32819_, _32822_);
  not g_63089_(_32822_, _32823_);
  and g_63090_(_31605_, _32820_, _32824_);
  or g_63091_(_31606_, _32819_, _32825_);
  and g_63092_(_31610_, _32825_, _32826_);
  or g_63093_(_31611_, _32824_, _32827_);
  and g_63094_(_32823_, _32826_, _32828_);
  or g_63095_(_32822_, _32827_, _32830_);
  and g_63096_(_32821_, _32830_, _32831_);
  and g_63097_(_31614_, _31618_, _32832_);
  xor g_63098_(_32831_, _32832_, _32833_);
  or g_63099_(_31622_, _32833_, _32834_);
  not g_63100_(_32834_, _32835_);
  and g_63101_(_31622_, _32833_, _32836_);
  xor g_63102_(_31622_, _32833_, _32837_);
  or g_63103_(_32835_, _32836_, _32838_);
  and g_63104_(_31625_, _31629_, _32839_);
  not g_63105_(_32839_, _32841_);
  and g_63106_(_32838_, _32839_, _32842_);
  or g_63107_(_32837_, _32841_, _32843_);
  or g_63108_(_32836_, _32839_, _32844_);
  not g_63109_(_32844_, _32845_);
  and g_63110_(_32834_, _32845_, _32846_);
  or g_63111_(_32835_, _32844_, _32847_);
  and g_63112_(_32843_, _32847_, _32848_);
  or g_63113_(_32842_, _32846_, _32849_);
  or g_63114_(_32615_, _32849_, _32850_);
  and g_63115_(_32615_, _32849_, _32852_);
  xor g_63116_(_32615_, _32848_, _32853_);
  xor g_63117_(_32614_, _32853_, _32854_);
  or g_63118_(_32612_, _32854_, _32855_);
  and g_63119_(_32612_, _32854_, _32856_);
  xor g_63120_(_32612_, _32854_, _32857_);
  xor g_63121_(_32610_, _32857_, _32858_);
  and g_63122_(_32605_, _32858_, _32859_);
  not g_63123_(_32859_, _32860_);
  and g_63124_(_31647_, _32858_, _32861_);
  xor g_63125_(_31647_, _32858_, _32863_);
  xor g_63126_(_31646_, _32858_, _32864_);
  and g_63127_(_32606_, _32864_, _32865_);
  or g_63128_(_32605_, _32863_, _32866_);
  and g_63129_(_32860_, _32866_, _32867_);
  or g_63130_(_32859_, _32865_, _32868_);
  or g_63131_(_31654_, _32868_, _32869_);
  not g_63132_(_32869_, _32870_);
  or g_63133_(_30388_, _31648_, _32871_);
  not g_63134_(_32871_, _32872_);
  or g_63135_(_32867_, _32871_, _32874_);
  and g_63136_(_32860_, _32871_, _32875_);
  or g_63137_(_32859_, _32872_, _32876_);
  or g_63138_(_32865_, _32876_, _32877_);
  and g_63139_(_31654_, _32877_, _32878_);
  and g_63140_(_32874_, _32878_, _32879_);
  or g_63141_(_32870_, _32879_, _32880_);
  xor g_63142_(_32604_, _32880_, _32881_);
  or g_63143_(_32601_, _32881_, _32882_);
  xor g_63144_(_32602_, _32881_, _32883_);
  not g_63145_(_32883_, _32885_);
  or g_63146_(_31663_, _32883_, _32886_);
  or g_63147_(_31661_, _32883_, _32887_);
  xor g_63148_(_31661_, _32883_, _32888_);
  xor g_63149_(_31661_, _32885_, _32889_);
  and g_63150_(_31663_, _32889_, _32890_);
  or g_63151_(_31665_, _32888_, _32891_);
  and g_63152_(_32886_, _32891_, _32892_);
  xor g_63153_(_31668_, _32892_, _32893_);
  or g_63154_(_31671_, _32893_, _32894_);
  and g_63155_(_31671_, _32893_, _32896_);
  xor g_63156_(_31671_, _32893_, _32897_);
  xor g_63157_(_32600_, _32897_, _32898_);
  or g_63158_(_32599_, _32898_, _32899_);
  not g_63159_(_32899_, _32900_);
  xor g_63160_(_32599_, _32898_, _32901_);
  and g_63161_(_31677_, _32901_, _32902_);
  xor g_63162_(_31677_, _32901_, _32903_);
  xor g_63163_(_31678_, _32901_, _32904_);
  and g_63164_(_31681_, _31685_, _32905_);
  not g_63165_(_32905_, _32907_);
  and g_63166_(_32904_, _32905_, _32908_);
  or g_63167_(_32903_, _32907_, _32909_);
  and g_63168_(_31682_, _32903_, _32910_);
  or g_63169_(_31681_, _32904_, _32911_);
  and g_63170_(_31687_, _32903_, _32912_);
  or g_63171_(_31685_, _32904_, _32913_);
  and g_63172_(_32911_, _32913_, _32914_);
  or g_63173_(_32910_, _32912_, _32915_);
  and g_63174_(_32909_, _32914_, _32916_);
  or g_63175_(_32908_, _32915_, _32918_);
  or g_63176_(_30416_, _31694_, _32919_);
  not g_63177_(_32919_, _32920_);
  and g_63178_(_31688_, _32919_, _32921_);
  xor g_63179_(_32916_, _32921_, _32922_);
  or g_63180_(_30432_, _31695_, _32923_);
  or g_63181_(_30430_, _31694_, _32924_);
  and g_63182_(_32923_, _32924_, _32925_);
  not g_63183_(_32925_, _32926_);
  xor g_63184_(_32922_, _32926_, _32927_);
  not g_63185_(_32927_, _32929_);
  or g_63186_(_30437_, _31698_, _32930_);
  or g_63187_(_30435_, _31695_, _32931_);
  and g_63188_(_32930_, _32931_, _32932_);
  xor g_63189_(_32929_, _32932_, _32933_);
  xor g_63190_(_32597_, _32933_, _32934_);
  not g_63191_(_32934_, _32935_);
  xor g_63192_(_32595_, _32934_, _32936_);
  xor g_63193_(_31712_, _32936_, _32937_);
  and g_63194_(_31714_, _32937_, _32938_);
  xor g_63195_(_31714_, _32937_, _32940_);
  not g_63196_(_32940_, _32941_);
  or g_63197_(_32594_, _32941_, _32942_);
  xor g_63198_(_32594_, _32940_, _32943_);
  not g_63199_(_32943_, _32944_);
  or g_63200_(_32593_, _32943_, _32945_);
  xor g_63201_(_32593_, _32944_, _32946_);
  not g_63202_(_32946_, _32947_);
  or g_63203_(_30473_, _31723_, _32948_);
  not g_63204_(_32948_, _32949_);
  and g_63205_(_31721_, _32948_, _32951_);
  xor g_63206_(_32946_, _32951_, _32952_);
  and g_63207_(_32592_, _32952_, _32953_);
  xor g_63208_(_32592_, _32952_, _32954_);
  not g_63209_(_32954_, _32955_);
  or g_63210_(_31728_, _32955_, _32956_);
  not g_63211_(_32956_, _32957_);
  xor g_63212_(_31728_, _32954_, _32958_);
  not g_63213_(_32958_, _32959_);
  and g_63214_(_31738_, _32959_, _32960_);
  or g_63215_(_31739_, _32958_, _32962_);
  xor g_63216_(_31738_, _32958_, _32963_);
  not g_63217_(_32963_, _32964_);
  and g_63218_(_31737_, _31745_, _32965_);
  xor g_63219_(_32963_, _32965_, _32966_);
  and g_63220_(_31748_, _32966_, _32967_);
  xor g_63221_(_31748_, _32966_, _32968_);
  not g_63222_(_32968_, _32969_);
  or g_63223_(_32591_, _32969_, _32970_);
  not g_63224_(_32970_, _32971_);
  xor g_63225_(_32591_, _32968_, _32973_);
  xor g_63226_(_32590_, _32973_, _32974_);
  not g_63227_(_32974_, _32975_);
  xor g_63228_(_31762_, _32974_, _32976_);
  and g_63229_(_31772_, _32976_, _32977_);
  and g_63230_(_31779_, _32977_, _32978_);
  or g_63231_(_31779_, _32976_, _32979_);
  not g_63232_(_32979_, _32980_);
  or g_63233_(_31772_, _32976_, _32981_);
  and g_63234_(_32979_, _32981_, _32982_);
  not g_63235_(_32982_, _32984_);
  or g_63236_(_32978_, _32984_, _32985_);
  or g_63237_(_31775_, _32985_, _32986_);
  xor g_63238_(_31776_, _32985_, _32987_);
  and g_63239_(_31783_, _31786_, _32988_);
  not g_63240_(_32988_, _32989_);
  xor g_63241_(_32987_, _32989_, _32990_);
  or g_63242_(_31788_, _32990_, _32991_);
  not g_63243_(_32991_, _32992_);
  xor g_63244_(_31788_, _32990_, _32993_);
  not g_63245_(_32993_, _32995_);
  and g_63246_(_31795_, _32993_, _32996_);
  or g_63247_(_31794_, _32995_, _32997_);
  xor g_63248_(_31794_, _32993_, _32998_);
  or g_63249_(_31800_, _32998_, _32999_);
  not g_63250_(_32999_, _33000_);
  xor g_63251_(_31799_, _32998_, _33001_);
  and g_63252_(_32586_, _33001_, _33002_);
  or g_63253_(_32586_, _33001_, _33003_);
  xor g_63254_(_32588_, _33001_, _33004_);
  or g_63255_(_30535_, _30537_, _33006_);
  or g_63256_(_31801_, _33006_, _33007_);
  and g_63257_(_31803_, _33007_, _33008_);
  not g_63258_(_33008_, _33009_);
  xor g_63259_(_33004_, _33009_, _33010_);
  xor g_63260_(_32584_, _33010_, _33011_);
  or g_63261_(_32581_, _33011_, _33012_);
  not g_63262_(_33012_, _33013_);
  xor g_63263_(_32582_, _33011_, _33014_);
  or g_63264_(_32579_, _33014_, _33015_);
  and g_63265_(_32579_, _33014_, _33017_);
  xor g_63266_(_32580_, _33014_, _33018_);
  not g_63267_(_33018_, _33019_);
  or g_63268_(_31814_, _33018_, _33020_);
  xor g_63269_(_31814_, _33019_, _33021_);
  and g_63270_(_31816_, _33021_, _33022_);
  or g_63271_(_31816_, _33018_, _33023_);
  not g_63272_(_33023_, _33024_);
  or g_63273_(_33022_, _33024_, _33025_);
  and g_63274_(_31819_, _31825_, _33026_);
  not g_63275_(_33026_, _33028_);
  xor g_63276_(_33025_, _33028_, _33029_);
  or g_63277_(_31821_, _33029_, _33030_);
  xor g_63278_(_31821_, _33029_, _33031_);
  and g_63279_(_32578_, _33031_, _33032_);
  xor g_63280_(_32577_, _33031_, _33033_);
  not g_63281_(_33033_, _33034_);
  and g_63282_(_32575_, _33034_, _33035_);
  not g_63283_(_33035_, _33036_);
  and g_63284_(_32574_, _33033_, _33037_);
  xor g_63285_(_32575_, _33033_, _33039_);
  not g_63286_(_33039_, _33040_);
  or g_63287_(_31842_, _33039_, _33041_);
  not g_63288_(_33041_, _33042_);
  xor g_63289_(_31842_, _33040_, _33043_);
  not g_63290_(_33043_, _33044_);
  and g_63291_(_31836_, _31846_, _33045_);
  or g_63292_(_33043_, _33045_, _33046_);
  xor g_63293_(_33043_, _33045_, _33047_);
  xor g_63294_(_33044_, _33045_, _33048_);
  or g_63295_(_31848_, _33048_, _33050_);
  xor g_63296_(_31848_, _33047_, _33051_);
  or g_63297_(_32573_, _33051_, _33052_);
  xor g_63298_(_32573_, _33051_, _33053_);
  and g_63299_(_32572_, _33053_, _33054_);
  xor g_63300_(_32571_, _33053_, _33055_);
  not g_63301_(_33055_, _33056_);
  and g_63302_(_31854_, _33056_, _33057_);
  xor g_63303_(_31854_, _33055_, _33058_);
  not g_63304_(_33058_, _33059_);
  and g_63305_(_32570_, _33059_, _33061_);
  xor g_63306_(_32569_, _33058_, _33062_);
  and g_63307_(_32568_, _33062_, _33063_);
  xor g_63308_(_32567_, _33062_, _33064_);
  or g_63309_(_31859_, _33064_, _33065_);
  not g_63310_(_33065_, _33066_);
  xor g_63311_(_31859_, _33064_, _33067_);
  not g_63312_(_33067_, _33068_);
  or g_63313_(_31861_, _33068_, _33069_);
  not g_63314_(_33069_, _33070_);
  xor g_63315_(_31861_, _33067_, _33072_);
  not g_63316_(_33072_, _33073_);
  or g_63317_(_32566_, _33072_, _33074_);
  xor g_63318_(_32566_, _33072_, _33075_);
  xor g_63319_(_32566_, _33073_, _33076_);
  or g_63320_(_32564_, _33076_, _33077_);
  xor g_63321_(_32564_, _33075_, _33078_);
  or g_63322_(_31871_, _33078_, _33079_);
  xor g_63323_(_31872_, _33078_, _33080_);
  not g_63324_(_33080_, _33081_);
  and g_63325_(_31870_, _33080_, _33083_);
  or g_63326_(_31870_, _33080_, _33084_);
  xor g_63327_(_31870_, _33080_, _33085_);
  xor g_63328_(_31870_, _33081_, _33086_);
  or g_63329_(_30633_, _31878_, _33087_);
  and g_63330_(_31877_, _33087_, _33088_);
  xor g_63331_(_33085_, _33088_, _33089_);
  or g_63332_(_32562_, _33089_, _33090_);
  and g_63333_(_32562_, _33089_, _33091_);
  xor g_63334_(_32563_, _33089_, _33092_);
  or g_63335_(_32560_, _33092_, _33094_);
  xor g_63336_(_32561_, _33092_, _33095_);
  or g_63337_(_30640_, _31879_, _33096_);
  and g_63338_(_31882_, _33096_, _33097_);
  or g_63339_(_33095_, _33097_, _33098_);
  xor g_63340_(_33095_, _33097_, _33099_);
  not g_63341_(_33099_, _33100_);
  or g_63342_(_31886_, _33100_, _33101_);
  xor g_63343_(_31886_, _33099_, _33102_);
  xor g_63344_(_31892_, _33102_, _33103_);
  not g_63345_(_33103_, _33105_);
  xor g_63346_(_31902_, _33103_, _33106_);
  or g_63347_(_31908_, _33106_, _33107_);
  not g_63348_(_33107_, _33108_);
  xor g_63349_(_31908_, _33106_, _33109_);
  not g_63350_(_33109_, _33110_);
  or g_63351_(_31911_, _33110_, _33111_);
  xor g_63352_(_31911_, _33109_, _33112_);
  not g_63353_(_33112_, _33113_);
  and g_63354_(_31913_, _31918_, _33114_);
  xor g_63355_(_33113_, _33114_, _33116_);
  or g_63356_(_31920_, _33116_, _33117_);
  xor g_63357_(_31921_, _33116_, _33118_);
  or g_63358_(_31923_, _33118_, _33119_);
  not g_63359_(_33119_, _33120_);
  and g_63360_(_31923_, _33118_, _33121_);
  xor g_63361_(_31923_, _33118_, _33122_);
  or g_63362_(_33120_, _33121_, _33123_);
  and g_63363_(_31926_, _33122_, _33124_);
  or g_63364_(_31925_, _33123_, _33125_);
  or g_63365_(_31929_, _33123_, _33127_);
  xor g_63366_(_31929_, _33122_, _33128_);
  and g_63367_(_31925_, _33128_, _33129_);
  or g_63368_(_33124_, _33129_, _33130_);
  or g_63369_(_31932_, _33130_, _33131_);
  xor g_63370_(_31933_, _33130_, _33132_);
  and g_63371_(_31936_, _31938_, _33133_);
  xor g_63372_(_33132_, _33133_, _33134_);
  not g_63373_(_33134_, _33135_);
  or g_63374_(_31941_, _33135_, _33136_);
  xor g_63375_(_31941_, _33134_, _33138_);
  not g_63376_(_33138_, _33139_);
  or g_63377_(_31945_, _33138_, _33140_);
  not g_63378_(_33140_, _33141_);
  xor g_63379_(_31945_, _33139_, _33142_);
  or g_63380_(_31943_, _33142_, _33143_);
  not g_63381_(_33143_, _33144_);
  or g_63382_(_30701_, _31947_, _33145_);
  not g_63383_(_33145_, _33146_);
  and g_63384_(_33139_, _33146_, _33147_);
  and g_63385_(_33142_, _33145_, _33149_);
  or g_63386_(_33147_, _33149_, _33150_);
  and g_63387_(_31943_, _33150_, _33151_);
  or g_63388_(_33144_, _33151_, _33152_);
  or g_63389_(_32559_, _33152_, _33153_);
  not g_63390_(_33153_, _33154_);
  xor g_63391_(_32559_, _33152_, _33155_);
  xor g_63392_(_32558_, _33152_, _33156_);
  and g_63393_(_31960_, _33155_, _33157_);
  or g_63394_(_31962_, _33156_, _33158_);
  xor g_63395_(_31960_, _33156_, _33160_);
  or g_63396_(_31959_, _33160_, _33161_);
  xor g_63397_(_31959_, _33160_, _33162_);
  xor g_63398_(_31958_, _33160_, _33163_);
  or g_63399_(_31965_, _33163_, _33164_);
  xor g_63400_(_31965_, _33162_, _33165_);
  not g_63401_(_33165_, _33166_);
  and g_63402_(_31973_, _33166_, _33167_);
  not g_63403_(_33167_, _33168_);
  xor g_63404_(_31973_, _33165_, _33169_);
  not g_63405_(_33169_, _33171_);
  and g_63406_(_31974_, _33171_, _33172_);
  xor g_63407_(_31974_, _33169_, _33173_);
  and g_63408_(_31977_, _31980_, _33174_);
  not g_63409_(_33174_, _33175_);
  xor g_63410_(_33173_, _33175_, _33176_);
  xor g_63411_(_33173_, _33174_, _33177_);
  xor g_63412_(_32557_, _33176_, _33178_);
  xor g_63413_(_32557_, _33177_, _33179_);
  and g_63414_(_32555_, _33178_, _33180_);
  or g_63415_(_32556_, _33179_, _33182_);
  and g_63416_(_31990_, _33178_, _33183_);
  not g_63417_(_33183_, _33184_);
  and g_63418_(_33182_, _33184_, _33185_);
  or g_63419_(_33180_, _33183_, _33186_);
  and g_63420_(_31989_, _33179_, _33187_);
  and g_63421_(_32556_, _33187_, _33188_);
  or g_63422_(_33186_, _33188_, _33189_);
  or g_63423_(_32552_, _33189_, _33190_);
  xor g_63424_(_32553_, _33189_, _33191_);
  or g_63425_(_31997_, _33191_, _33193_);
  xor g_63426_(_31998_, _33191_, _33194_);
  or g_63427_(_32000_, _33194_, _33195_);
  xor g_63428_(_32000_, _33194_, _33196_);
  not g_63429_(_33196_, _33197_);
  or g_63430_(_30740_, _32004_, _33198_);
  not g_63431_(_33198_, _33199_);
  and g_63432_(_32002_, _33198_, _33200_);
  xor g_63433_(_33196_, _33200_, _33201_);
  or g_63434_(_32551_, _33201_, _33202_);
  xor g_63435_(_32551_, _33201_, _33204_);
  not g_63436_(_33204_, _33205_);
  or g_63437_(_32550_, _33205_, _33206_);
  xor g_63438_(_32550_, _33204_, _33207_);
  and g_63439_(_32548_, _33207_, _33208_);
  or g_63440_(_32548_, _33207_, _33209_);
  xor g_63441_(_32549_, _33207_, _33210_);
  not g_63442_(_33210_, _33211_);
  and g_63443_(_32013_, _32015_, _33212_);
  xor g_63444_(_33210_, _33212_, _33213_);
  and g_63445_(_32019_, _33213_, _33215_);
  xor g_63446_(_32019_, _33213_, _33216_);
  xor g_63447_(_32020_, _33213_, _33217_);
  or g_63448_(_32022_, _33217_, _33218_);
  not g_63449_(_33218_, _33219_);
  xor g_63450_(_32022_, _33216_, _33220_);
  or g_63451_(_32024_, _33220_, _33221_);
  xor g_63452_(_32024_, _33220_, _33222_);
  not g_63453_(_33222_, _33223_);
  or g_63454_(_32026_, _33223_, _33224_);
  not g_63455_(_33224_, _33226_);
  xor g_63456_(_32026_, _33222_, _33227_);
  or g_63457_(_32029_, _33227_, _33228_);
  xor g_63458_(_32029_, _33227_, _33229_);
  xor g_63459_(_32030_, _33227_, _33230_);
  and g_63460_(_32032_, _33230_, _33231_);
  or g_63461_(_32033_, _33229_, _33232_);
  and g_63462_(_32039_, _33231_, _33233_);
  or g_63463_(_32040_, _33232_, _33234_);
  or g_63464_(_32039_, _33230_, _33235_);
  not g_63465_(_33235_, _33237_);
  or g_63466_(_32032_, _33230_, _33238_);
  not g_63467_(_33238_, _33239_);
  and g_63468_(_33235_, _33238_, _33240_);
  not g_63469_(_33240_, _33241_);
  and g_63470_(_33234_, _33240_, _33242_);
  or g_63471_(_33233_, _33241_, _33243_);
  or g_63472_(_32041_, _33243_, _33244_);
  xor g_63473_(_32041_, _33242_, _33245_);
  not g_63474_(_33245_, _33246_);
  and g_63475_(_32045_, _32047_, _33248_);
  xor g_63476_(_33245_, _33248_, _33249_);
  xor g_63477_(_33246_, _33248_, _33250_);
  or g_63478_(_32547_, _33250_, _33251_);
  xor g_63479_(_32547_, _33249_, _33252_);
  or g_63480_(_32546_, _33252_, _33253_);
  not g_63481_(_33253_, _33254_);
  xor g_63482_(_32546_, _33252_, _33255_);
  not g_63483_(_33255_, _33256_);
  or g_63484_(_30792_, _32050_, _33257_);
  and g_63485_(_32051_, _33257_, _33259_);
  xor g_63486_(_33255_, _33259_, _33260_);
  not g_63487_(_33260_, _33261_);
  or g_63488_(_32545_, _33260_, _33262_);
  xor g_63489_(_32545_, _33260_, _33263_);
  xor g_63490_(_32545_, _33261_, _33264_);
  or g_63491_(_32057_, _33264_, _33265_);
  xor g_63492_(_32057_, _33263_, _33266_);
  or g_63493_(_32059_, _33266_, _33267_);
  xor g_63494_(_32061_, _33266_, _33268_);
  not g_63495_(_33268_, _33270_);
  and g_63496_(_32069_, _33270_, _33271_);
  not g_63497_(_33271_, _33272_);
  xor g_63498_(_32068_, _33268_, _33273_);
  and g_63499_(_32067_, _33273_, _33274_);
  not g_63500_(_33274_, _33275_);
  xor g_63501_(_32067_, _33273_, _33276_);
  or g_63502_(_30820_, _32077_, _33277_);
  not g_63503_(_33277_, _33278_);
  and g_63504_(_32076_, _33277_, _33279_);
  xor g_63505_(_33276_, _33279_, _33281_);
  or g_63506_(_32542_, _33281_, _33282_);
  xor g_63507_(_32542_, _33281_, _33283_);
  xor g_63508_(_32544_, _33281_, _33284_);
  and g_63509_(_32081_, _33284_, _33285_);
  and g_63510_(_32087_, _33285_, _33286_);
  and g_63511_(_32083_, _33283_, _33287_);
  not g_63512_(_33287_, _33288_);
  and g_63513_(_32086_, _33283_, _33289_);
  or g_63514_(_32087_, _33284_, _33290_);
  or g_63515_(_33287_, _33289_, _33292_);
  or g_63516_(_33286_, _33292_, _33293_);
  not g_63517_(_33293_, _33294_);
  or g_63518_(_32092_, _33293_, _33295_);
  not g_63519_(_33295_, _33296_);
  or g_63520_(_32089_, _33293_, _33297_);
  xor g_63521_(_32089_, _33293_, _33298_);
  xor g_63522_(_32089_, _33294_, _33299_);
  and g_63523_(_32092_, _33299_, _33300_);
  or g_63524_(_32094_, _33298_, _33301_);
  and g_63525_(_33295_, _33301_, _33303_);
  or g_63526_(_33296_, _33300_, _33304_);
  and g_63527_(_32098_, _32101_, _33305_);
  xor g_63528_(_33303_, _33305_, _33306_);
  or g_63529_(_32541_, _33306_, _33307_);
  xor g_63530_(_32541_, _33306_, _33308_);
  not g_63531_(_33308_, _33309_);
  or g_63532_(_32540_, _33309_, _33310_);
  not g_63533_(_33310_, _33311_);
  xor g_63534_(_32540_, _33308_, _33312_);
  or g_63535_(_32538_, _33312_, _33314_);
  xor g_63536_(_32539_, _33312_, _33315_);
  not g_63537_(_33315_, _33316_);
  or g_63538_(_32537_, _33315_, _33317_);
  xor g_63539_(_32537_, _33315_, _33318_);
  xor g_63540_(_32537_, _33316_, _33319_);
  and g_63541_(_32109_, _32111_, _33320_);
  xor g_63542_(_33318_, _33320_, _33321_);
  xor g_63543_(_33319_, _33320_, _33322_);
  and g_63544_(_32536_, _33322_, _33323_);
  xor g_63545_(_32535_, _33321_, _33325_);
  not g_63546_(_33325_, _33326_);
  or g_63547_(_32534_, _33326_, _33327_);
  xor g_63548_(_32534_, _33325_, _33328_);
  or g_63549_(_32531_, _33328_, _33329_);
  xor g_63550_(_32533_, _33328_, _33330_);
  or g_63551_(_32530_, _33330_, _33331_);
  xor g_63552_(_32530_, _33330_, _33332_);
  or g_63553_(_32117_, _33332_, _33333_);
  not g_63554_(_33333_, _33334_);
  and g_63555_(_32117_, _33332_, _33336_);
  not g_63556_(_33336_, _33337_);
  xor g_63557_(_32117_, _33332_, _33338_);
  or g_63558_(_33334_, _33336_, _33339_);
  and g_63559_(_32119_, _32123_, _33340_);
  xor g_63560_(_33338_, _33340_, _33341_);
  or g_63561_(_32125_, _33341_, _33342_);
  xor g_63562_(_32127_, _33341_, _33343_);
  not g_63563_(_33343_, _33344_);
  and g_63564_(_32131_, _33343_, _33345_);
  or g_63565_(_32131_, _33343_, _33347_);
  xor g_63566_(_32131_, _33343_, _33348_);
  xor g_63567_(_32131_, _33344_, _33349_);
  and g_63568_(_32134_, _32138_, _33350_);
  xor g_63569_(_33348_, _33350_, _33351_);
  xor g_63570_(_32529_, _33351_, _33352_);
  not g_63571_(_33352_, _33353_);
  and g_63572_(_32146_, _33352_, _33354_);
  not g_63573_(_33354_, _33355_);
  and g_63574_(_30904_, _32141_, _33356_);
  not g_63575_(_33356_, _33358_);
  or g_63576_(_33352_, _33356_, _33359_);
  or g_63577_(_32146_, _33359_, _33360_);
  or g_63578_(_33353_, _33358_, _33361_);
  and g_63579_(_33360_, _33361_, _33362_);
  and g_63580_(_33355_, _33362_, _33363_);
  and g_63581_(_32527_, _33363_, _33364_);
  xor g_63582_(_32526_, _33363_, _33365_);
  or g_63583_(_32524_, _33365_, _33366_);
  not g_63584_(_33366_, _33367_);
  xor g_63585_(_32524_, _33365_, _33369_);
  xor g_63586_(_32525_, _33365_, _33370_);
  and g_63587_(_32155_, _33369_, _33371_);
  and g_63588_(_32152_, _33370_, _33372_);
  and g_63589_(_32156_, _33372_, _33373_);
  and g_63590_(_32153_, _33369_, _33374_);
  or g_63591_(_33373_, _33374_, _33375_);
  or g_63592_(_33371_, _33375_, _33376_);
  not g_63593_(_33376_, _33377_);
  and g_63594_(_32523_, _33377_, _33378_);
  and g_63595_(_32158_, _33376_, _33380_);
  and g_63596_(_32522_, _33380_, _33381_);
  or g_63597_(_32158_, _33376_, _33382_);
  not g_63598_(_33382_, _33383_);
  or g_63599_(_33381_, _33383_, _33384_);
  or g_63600_(_33378_, _33384_, _33385_);
  or g_63601_(_32519_, _33385_, _33386_);
  not g_63602_(_33386_, _33387_);
  xor g_63603_(_32520_, _33385_, _33388_);
  or g_63604_(_32518_, _33388_, _33389_);
  not g_63605_(_33389_, _33391_);
  and g_63606_(_32167_, _33388_, _33392_);
  and g_63607_(_32518_, _33392_, _33393_);
  or g_63608_(_32167_, _33388_, _33394_);
  not g_63609_(_33394_, _33395_);
  or g_63610_(_33393_, _33395_, _33396_);
  or g_63611_(_33391_, _33396_, _33397_);
  not g_63612_(_33397_, _33398_);
  or g_63613_(_32517_, _33397_, _33399_);
  xor g_63614_(_32517_, _33397_, _33400_);
  xor g_63615_(_32517_, _33398_, _33402_);
  and g_63616_(_32173_, _32177_, _33403_);
  xor g_63617_(_33400_, _33403_, _33404_);
  or g_63618_(_32179_, _33404_, _33405_);
  xor g_63619_(_32180_, _33404_, _33406_);
  and g_63620_(_32185_, _33406_, _33407_);
  or g_63621_(_32185_, _33404_, _33408_);
  not g_63622_(_33408_, _33409_);
  or g_63623_(_33407_, _33409_, _33410_);
  or g_63624_(_32189_, _32191_, _33411_);
  and g_63625_(_32188_, _33411_, _33413_);
  not g_63626_(_33413_, _33414_);
  xor g_63627_(_33410_, _33414_, _33415_);
  or g_63628_(_32515_, _33415_, _33416_);
  xor g_63629_(_32516_, _33415_, _33417_);
  not g_63630_(_33417_, _33418_);
  and g_63631_(_32514_, _33418_, _33419_);
  xor g_63632_(_32514_, _33417_, _33420_);
  and g_63633_(_32198_, _32201_, _33421_);
  not g_63634_(_33421_, _33422_);
  xor g_63635_(_33420_, _33421_, _33424_);
  xor g_63636_(_33420_, _33422_, _33425_);
  and g_63637_(_32204_, _33425_, _33426_);
  and g_63638_(_32209_, _33426_, _33427_);
  and g_63639_(_32208_, _33424_, _33428_);
  or g_63640_(_32209_, _33425_, _33429_);
  and g_63641_(_32205_, _33424_, _33430_);
  or g_63642_(_32204_, _33425_, _33431_);
  or g_63643_(_33428_, _33430_, _33432_);
  or g_63644_(_33427_, _33432_, _33433_);
  and g_63645_(_32211_, _33433_, _33435_);
  or g_63646_(_32211_, _33433_, _33436_);
  xor g_63647_(_32211_, _33433_, _33437_);
  and g_63648_(_32213_, _32217_, _33438_);
  xor g_63649_(_33437_, _33438_, _33439_);
  or g_63650_(_32222_, _33439_, _33440_);
  not g_63651_(_33440_, _33441_);
  xor g_63652_(_32222_, _33439_, _33442_);
  and g_63653_(_32513_, _33442_, _33443_);
  xor g_63654_(_32512_, _33442_, _33444_);
  or g_63655_(_32511_, _33444_, _33446_);
  not g_63656_(_33446_, _33447_);
  xor g_63657_(_32511_, _33444_, _33448_);
  not g_63658_(_33448_, _33449_);
  and g_63659_(_32509_, _33448_, _33450_);
  or g_63660_(_32508_, _33449_, _33451_);
  and g_63661_(_32508_, _33449_, _33452_);
  xor g_63662_(_32509_, _33448_, _33453_);
  xor g_63663_(_32508_, _33448_, _33454_);
  or g_63664_(_32506_, _33454_, _33455_);
  not g_63665_(_33455_, _33457_);
  and g_63666_(_32232_, _33453_, _33458_);
  xor g_63667_(_32231_, _33454_, _33459_);
  xor g_63668_(_32231_, _33453_, _33460_);
  and g_63669_(_32506_, _33460_, _33461_);
  or g_63670_(_32507_, _33459_, _33462_);
  and g_63671_(_33455_, _33462_, _33463_);
  or g_63672_(_33457_, _33461_, _33464_);
  and g_63673_(_32235_, _32239_, _33465_);
  and g_63674_(_33464_, _33465_, _33466_);
  and g_63675_(_32237_, _33463_, _33468_);
  or g_63676_(_32235_, _33464_, _33469_);
  and g_63677_(_32240_, _33463_, _33470_);
  or g_63678_(_32239_, _33464_, _33471_);
  or g_63679_(_33468_, _33470_, _33472_);
  or g_63680_(_33466_, _33472_, _33473_);
  and g_63681_(_32242_, _32251_, _33474_);
  not g_63682_(_33474_, _33475_);
  xor g_63683_(_33473_, _33475_, _33476_);
  or g_63684_(_32250_, _33476_, _33477_);
  xor g_63685_(_32250_, _33476_, _33479_);
  xor g_63686_(_32249_, _33476_, _33480_);
  or g_63687_(_32263_, _33480_, _33481_);
  not g_63688_(_33481_, _33482_);
  and g_63689_(_32259_, _33480_, _33483_);
  or g_63690_(_32257_, _33479_, _33484_);
  and g_63691_(_32263_, _33483_, _33485_);
  or g_63692_(_32262_, _33484_, _33486_);
  and g_63693_(_32257_, _33479_, _33487_);
  not g_63694_(_33487_, _33488_);
  and g_63695_(_33486_, _33488_, _33490_);
  or g_63696_(_33485_, _33487_, _33491_);
  and g_63697_(_33481_, _33490_, _33492_);
  or g_63698_(_33482_, _33491_, _33493_);
  xor g_63699_(_32505_, _33493_, _33494_);
  xor g_63700_(_32505_, _33492_, _33495_);
  and g_63701_(_31007_, _32272_, _33496_);
  and g_63702_(_33494_, _33496_, _33497_);
  not g_63703_(_33497_, _33498_);
  or g_63704_(_31008_, _32271_, _33499_);
  not g_63705_(_33499_, _33501_);
  and g_63706_(_33494_, _33501_, _33502_);
  not g_63707_(_33502_, _33503_);
  and g_63708_(_32276_, _33495_, _33504_);
  or g_63709_(_32275_, _33494_, _33505_);
  and g_63710_(_33503_, _33505_, _33506_);
  or g_63711_(_33502_, _33504_, _33507_);
  and g_63712_(_33498_, _33506_, _33508_);
  or g_63713_(_33497_, _33507_, _33509_);
  and g_63714_(_32278_, _33509_, _33510_);
  and g_63715_(_32279_, _33508_, _33512_);
  or g_63716_(_32278_, _33509_, _33513_);
  xor g_63717_(_32279_, _33509_, _33514_);
  not g_63718_(_33514_, _33515_);
  and g_63719_(_32283_, _32286_, _33516_);
  xor g_63720_(_33515_, _33516_, _33517_);
  xor g_63721_(_33514_, _33516_, _33518_);
  or g_63722_(_32288_, _33517_, _33519_);
  xor g_63723_(_32288_, _33518_, _33520_);
  not g_63724_(_33520_, _33521_);
  or g_63725_(_32292_, _33520_, _33523_);
  not g_63726_(_33523_, _33524_);
  xor g_63727_(_32292_, _33520_, _33525_);
  and g_63728_(_32301_, _33525_, _33526_);
  not g_63729_(_33526_, _33527_);
  or g_63730_(_32301_, _33521_, _33528_);
  and g_63731_(_33527_, _33528_, _33529_);
  or g_63732_(_32311_, _33529_, _33530_);
  xor g_63733_(_32311_, _33529_, _33531_);
  and g_63734_(_32319_, _33531_, _33532_);
  and g_63735_(_32308_, _33531_, _33534_);
  not g_63736_(_33534_, _33535_);
  xor g_63737_(_32307_, _33531_, _33536_);
  and g_63738_(_32320_, _33536_, _33537_);
  or g_63739_(_33532_, _33537_, _33538_);
  xor g_63740_(_32328_, _33538_, _33539_);
  not g_63741_(_33539_, _33540_);
  xor g_63742_(_32504_, _33539_, _33541_);
  and g_63743_(_32336_, _33541_, _33542_);
  xor g_63744_(_32336_, _33541_, _33543_);
  xor g_63745_(_32337_, _33541_, _33545_);
  and g_63746_(_32342_, _33543_, _33546_);
  or g_63747_(_32341_, _33545_, _33547_);
  xor g_63748_(_32342_, _33543_, _33548_);
  xor g_63749_(_32341_, _33543_, _33549_);
  and g_63750_(_32347_, _32351_, _33550_);
  xor g_63751_(_33548_, _33550_, _33551_);
  not g_63752_(_33551_, _33552_);
  and g_63753_(_31085_, _32355_, _33553_);
  or g_63754_(_31086_, _32356_, _33554_);
  and g_63755_(_32354_, _33554_, _33556_);
  xor g_63756_(_33552_, _33556_, _33557_);
  or g_63757_(_32502_, _33557_, _33558_);
  xor g_63758_(_32502_, _33557_, _33559_);
  xor g_63759_(_32503_, _33557_, _33560_);
  and g_63760_(_32361_, _33559_, _33561_);
  or g_63761_(_32362_, _33560_, _33562_);
  xor g_63762_(_32362_, _33559_, _33563_);
  or g_63763_(_32365_, _33563_, _33564_);
  xor g_63764_(_32365_, _33563_, _33565_);
  not g_63765_(_33565_, _33567_);
  and g_63766_(_32370_, _33565_, _33568_);
  or g_63767_(_32369_, _33567_, _33569_);
  xor g_63768_(_32369_, _33565_, _33570_);
  and g_63769_(_32372_, _33570_, _33571_);
  and g_63770_(_32377_, _33571_, _33572_);
  or g_63771_(_32372_, _33570_, _33573_);
  not g_63772_(_33573_, _33574_);
  or g_63773_(_32377_, _33570_, _33575_);
  and g_63774_(_33573_, _33575_, _33576_);
  not g_63775_(_33576_, _33578_);
  or g_63776_(_33572_, _33578_, _33579_);
  not g_63777_(_33579_, _33580_);
  or g_63778_(_31107_, _32383_, _33581_);
  not g_63779_(_33581_, _33582_);
  and g_63780_(_32374_, _33581_, _33583_);
  xor g_63781_(_33579_, _33583_, _33584_);
  not g_63782_(_33584_, _33585_);
  and g_63783_(_32501_, _33584_, _33586_);
  not g_63784_(_33586_, _33587_);
  xor g_63785_(_32501_, _33584_, _33589_);
  xor g_63786_(_32501_, _33585_, _33590_);
  or g_63787_(_32387_, _33590_, _33591_);
  xor g_63788_(_32387_, _33589_, _33592_);
  or g_63789_(_32500_, _33592_, _33593_);
  xor g_63790_(_32498_, _33592_, _33594_);
  or g_63791_(_32497_, _33594_, _33595_);
  not g_63792_(_33595_, _33596_);
  xor g_63793_(_32497_, _33594_, _33597_);
  and g_63794_(_32496_, _33597_, _33598_);
  xor g_63795_(_32496_, _33597_, _33600_);
  xor g_63796_(_32495_, _33597_, _33601_);
  or g_63797_(_32494_, _33601_, _33602_);
  xor g_63798_(_32494_, _33600_, _33603_);
  not g_63799_(_33603_, _33604_);
  or g_63800_(_32397_, _33603_, _33605_);
  xor g_63801_(_32397_, _33604_, _33606_);
  not g_63802_(_33606_, _33607_);
  and g_63803_(_32400_, _32404_, _33608_);
  or g_63804_(_33606_, _33608_, _33609_);
  xor g_63805_(_33606_, _33608_, _33611_);
  xor g_63806_(_33607_, _33608_, _33612_);
  or g_63807_(_31131_, _32408_, _33613_);
  and g_63808_(_32406_, _33613_, _33614_);
  xor g_63809_(_33611_, _33614_, _33615_);
  not g_63810_(_33615_, _33616_);
  and g_63811_(_32493_, _33616_, _33617_);
  xor g_63812_(_32492_, _33615_, _33618_);
  and g_63813_(_32415_, _33618_, _33619_);
  xor g_63814_(_32414_, _33618_, _33620_);
  not g_63815_(_33620_, _33622_);
  or g_63816_(_31143_, _32413_, _33623_);
  not g_63817_(_33623_, _33624_);
  and g_63818_(_33622_, _33624_, _33625_);
  xor g_63819_(_33620_, _33623_, _33626_);
  or g_63820_(_31146_, _32417_, _33627_);
  not g_63821_(_33627_, _33628_);
  and g_63822_(_32421_, _33627_, _33629_);
  xor g_63823_(_33626_, _33629_, _33630_);
  not g_63824_(_33630_, _33631_);
  xor g_63825_(_32427_, _33631_, _33633_);
  not g_63826_(_33633_, _33634_);
  xor g_63827_(_32491_, _33633_, _33635_);
  xor g_63828_(_32491_, _33634_, _33636_);
  or g_63829_(_32438_, _33636_, _33637_);
  not g_63830_(_33637_, _33638_);
  xor g_63831_(_32438_, _33635_, _33639_);
  not g_63832_(_33639_, _33640_);
  or g_63833_(_32440_, _33639_, _33641_);
  xor g_63834_(_32440_, _33639_, _33642_);
  xor g_63835_(_32440_, _33640_, _33644_);
  and g_63836_(_32444_, _33642_, _33645_);
  or g_63837_(_32443_, _33644_, _33646_);
  xor g_63838_(_32444_, _33642_, _33647_);
  xor g_63839_(_32443_, _33642_, _33648_);
  or g_63840_(_32447_, _33648_, _33649_);
  not g_63841_(_33649_, _33650_);
  xor g_63842_(_32447_, _33647_, _33651_);
  and g_63843_(_32450_, _33651_, _33652_);
  or g_63844_(_32450_, _33651_, _33653_);
  not g_63845_(_33653_, _33655_);
  or g_63846_(_33652_, _33655_, _33656_);
  not g_63847_(_33656_, _33657_);
  and g_63848_(_32453_, _32457_, _33658_);
  xor g_63849_(_33657_, _33658_, _33659_);
  xor g_63850_(_33656_, _33658_, _33660_);
  and g_63851_(_32460_, _33660_, _33661_);
  not g_63852_(_33661_, _33662_);
  xor g_63853_(_32459_, _33659_, _33663_);
  xor g_63854_(_32464_, _33663_, _33664_);
  not g_63855_(_33664_, _33666_);
  and g_63856_(_32490_, _33666_, _33667_);
  xor g_63857_(_32490_, _33664_, _33668_);
  not g_63858_(_33668_, _33669_);
  and g_63859_(_32489_, _33669_, _33670_);
  xor g_63860_(_32489_, _33668_, _33671_);
  not g_63861_(_33671_, _33672_);
  or g_63862_(_32472_, _33671_, _33673_);
  and g_63863_(_32472_, _33671_, _33674_);
  xor g_63864_(_32472_, _33672_, _33675_);
  not g_63865_(_33675_, _33677_);
  xor g_63866_(_32480_, _33675_, _33678_);
  xor g_63867_(_32480_, _33677_, _33679_);
  or g_63868_(_32484_, _33678_, _33680_);
  xor g_63869_(_32484_, _33679_, _33681_);
  or g_63870_(_32486_, _33681_, _33682_);
  xor g_63871_(_32486_, _33681_, out[645]);
  and g_63872_(_32475_, _33677_, _33683_);
  or g_63873_(_32476_, _33675_, _33684_);
  or g_63874_(_32462_, _33659_, _33685_);
  or g_63875_(_31183_, _33685_, _33687_);
  not g_63876_(_33687_, _33688_);
  or g_63877_(_31179_, _33685_, _33689_);
  or g_63878_(_32457_, _33656_, _33690_);
  not g_63879_(_33690_, _33691_);
  or g_63880_(_32453_, _33656_, _33692_);
  or g_63881_(_32433_, _33633_, _33693_);
  or g_63882_(_32430_, _33630_, _33694_);
  not g_63883_(_33694_, _33695_);
  or g_63884_(_31155_, _32424_, _33696_);
  or g_63885_(_33630_, _33696_, _33698_);
  not g_63886_(_33698_, _33699_);
  or g_63887_(_31151_, _32424_, _33700_);
  not g_63888_(_33700_, _33701_);
  and g_63889_(_33631_, _33701_, _33702_);
  not g_63890_(_33702_, _33703_);
  and g_63891_(_32422_, _33626_, _33704_);
  and g_63892_(_33626_, _33628_, _33705_);
  or g_63893_(_33612_, _33613_, _33706_);
  and g_63894_(_32407_, _33611_, _33707_);
  or g_63895_(_32406_, _33612_, _33709_);
  and g_63896_(_33591_, _33593_, _33710_);
  not g_63897_(_33710_, _33711_);
  and g_63898_(_33580_, _33582_, _33712_);
  and g_63899_(_33552_, _33553_, _33713_);
  or g_63900_(_33551_, _33554_, _33714_);
  or g_63901_(_32351_, _33549_, _33715_);
  not g_63902_(_33715_, _33716_);
  and g_63903_(_32348_, _33548_, _33717_);
  or g_63904_(_32347_, _33549_, _33718_);
  and g_63905_(_32339_, _33540_, _33720_);
  or g_63906_(_32332_, _33539_, _33721_);
  or g_63907_(_32325_, _33538_, _33722_);
  not g_63908_(_33722_, _33723_);
  or g_63909_(_32326_, _33538_, _33724_);
  not g_63910_(_33724_, _33725_);
  or g_63911_(_32298_, _33520_, _33726_);
  or g_63912_(_32300_, _33520_, _33727_);
  not g_63913_(_33727_, _33728_);
  or g_63914_(_32286_, _33514_, _33729_);
  not g_63915_(_33729_, _33731_);
  or g_63916_(_32270_, _33493_, _33732_);
  and g_63917_(_33503_, _33732_, _33733_);
  not g_63918_(_33733_, _33734_);
  or g_63919_(_32251_, _33473_, _33735_);
  or g_63920_(_32242_, _33473_, _33736_);
  and g_63921_(_32506_, _33451_, _33737_);
  or g_63922_(_33452_, _33737_, _33738_);
  or g_63923_(_32201_, _33420_, _33739_);
  or g_63924_(_33410_, _33411_, _33740_);
  not g_63925_(_33740_, _33742_);
  or g_63926_(_32188_, _33407_, _33743_);
  and g_63927_(_33408_, _33743_, _33744_);
  not g_63928_(_33744_, _33745_);
  or g_63929_(_32177_, _33402_, _33746_);
  and g_63930_(_32174_, _33400_, _33747_);
  or g_63931_(_32173_, _33402_, _33748_);
  or g_63932_(_32528_, _33351_, _33749_);
  not g_63933_(_33749_, _33750_);
  or g_63934_(_32123_, _33339_, _33751_);
  or g_63935_(_32111_, _33319_, _33753_);
  or g_63936_(_32109_, _33312_, _33754_);
  or g_63937_(_32101_, _33304_, _33755_);
  and g_63938_(_33276_, _33278_, _33756_);
  not g_63939_(_33756_, _33757_);
  and g_63940_(_30812_, _32073_, _33758_);
  and g_63941_(_33276_, _33758_, _33759_);
  or g_63942_(_30809_, _32074_, _33760_);
  not g_63943_(_33760_, _33761_);
  and g_63944_(_33273_, _33761_, _33762_);
  and g_63945_(_33262_, _33265_, _33764_);
  or g_63946_(_33256_, _33257_, _33765_);
  not g_63947_(_33765_, _33766_);
  and g_63948_(_32052_, _33255_, _33767_);
  or g_63949_(_32047_, _33245_, _33768_);
  not g_63950_(_33768_, _33769_);
  or g_63951_(_32045_, _33243_, _33770_);
  and g_63952_(_32017_, _33211_, _33771_);
  not g_63953_(_33771_, _33772_);
  and g_63954_(_32003_, _33196_, _33773_);
  not g_63955_(_33773_, _33775_);
  and g_63956_(_33193_, _33195_, _33776_);
  and g_63957_(_31987_, _33177_, _33777_);
  not g_63958_(_33777_, _33778_);
  or g_63959_(_31984_, _33176_, _33779_);
  or g_63960_(_31980_, _33173_, _33780_);
  or g_63961_(_31977_, _33173_, _33781_);
  or g_63962_(_31938_, _33132_, _33782_);
  not g_63963_(_33782_, _33783_);
  or g_63964_(_31936_, _33132_, _33784_);
  not g_63965_(_33784_, _33786_);
  or g_63966_(_31913_, _33112_, _33787_);
  or g_63967_(_31897_, _33105_, _33788_);
  or g_63968_(_31901_, _33105_, _33789_);
  or g_63969_(_31887_, _31889_, _33790_);
  or g_63970_(_33102_, _33790_, _33791_);
  not g_63971_(_33791_, _33792_);
  or g_63972_(_30649_, _31887_, _33793_);
  or g_63973_(_33102_, _33793_, _33794_);
  or g_63974_(_33086_, _33087_, _33795_);
  and g_63975_(_33077_, _33079_, _33797_);
  not g_63976_(_33797_, _33798_);
  and g_63977_(_33050_, _33052_, _33799_);
  or g_63978_(_31825_, _33025_, _33800_);
  or g_63979_(_31810_, _33010_, _33801_);
  or g_63980_(_31806_, _33010_, _33802_);
  or g_63981_(_31803_, _33004_, _33803_);
  and g_63982_(_33802_, _33803_, _33804_);
  and g_63983_(_33003_, _33007_, _33805_);
  or g_63984_(_33002_, _33805_, _33806_);
  not g_63985_(_33806_, _33808_);
  and g_63986_(_32997_, _32999_, _33809_);
  or g_63987_(_32996_, _33000_, _33810_);
  or g_63988_(_31786_, _32987_, _33811_);
  or g_63989_(_31783_, _32987_, _33812_);
  and g_63990_(_31759_, _32974_, _33813_);
  or g_63991_(_31758_, _32975_, _33814_);
  and g_63992_(_31761_, _32974_, _33815_);
  and g_63993_(_32589_, _32968_, _33816_);
  or g_63994_(_31737_, _32963_, _33817_);
  and g_63995_(_32947_, _32949_, _33819_);
  or g_63996_(_31710_, _32936_, _33820_);
  not g_63997_(_33820_, _33821_);
  or g_63998_(_30449_, _33820_, _33822_);
  not g_63999_(_33822_, _33823_);
  and g_64000_(_31706_, _32934_, _33824_);
  not g_64001_(_33824_, _33825_);
  or g_64002_(_31700_, _32935_, _33826_);
  or g_64003_(_31702_, _32933_, _33827_);
  or g_64004_(_32596_, _32933_, _33828_);
  or g_64005_(_32927_, _32930_, _33830_);
  or g_64006_(_32922_, _32924_, _33831_);
  and g_64007_(_32916_, _32920_, _33832_);
  not g_64008_(_33832_, _33833_);
  and g_64009_(_33831_, _33833_, _33834_);
  or g_64010_(_32900_, _32902_, _33835_);
  or g_64011_(_32600_, _32896_, _33836_);
  and g_64012_(_32894_, _33836_, _33837_);
  and g_64013_(_31668_, _32886_, _33838_);
  or g_64014_(_32890_, _33838_, _33839_);
  and g_64015_(_32882_, _32887_, _33841_);
  or g_64016_(_32603_, _32879_, _33842_);
  and g_64017_(_32869_, _33842_, _33843_);
  or g_64018_(_32865_, _32875_, _33844_);
  and g_64019_(_32611_, _32855_, _33845_);
  or g_64020_(_32856_, _33845_, _33846_);
  and g_64021_(_31617_, _32831_, _33847_);
  and g_64022_(_31614_, _32821_, _33848_);
  or g_64023_(_32828_, _33848_, _33849_);
  or g_64024_(_32621_, _32793_, _33850_);
  and g_64025_(_32792_, _33850_, _33852_);
  or g_64026_(_32626_, _32789_, _33853_);
  and g_64027_(_32788_, _33853_, _33854_);
  and g_64028_(_31595_, _32784_, _33855_);
  or g_64029_(_32782_, _33855_, _33856_);
  and g_64030_(_32770_, _32772_, _33857_);
  or g_64031_(_31580_, _32766_, _33858_);
  and g_64032_(_32767_, _33858_, _33859_);
  and g_64033_(_32760_, _32764_, _33860_);
  and g_64034_(_31559_, _32756_, _33861_);
  or g_64035_(_31556_, _32754_, _33863_);
  and g_64036_(_32755_, _33863_, _33864_);
  and g_64037_(_31550_, _32744_, _33865_);
  or g_64038_(_32743_, _33865_, _33866_);
  and g_64039_(_32699_, _32710_, _33867_);
  or g_64040_(_31503_, _32693_, _33868_);
  and g_64041_(_32695_, _33868_, _33869_);
  and g_64042_(_32687_, _32691_, _33870_);
  or g_64043_(_32682_, _33870_, _33871_);
  or g_64044_(_32683_, _32690_, _33872_);
  and g_64045_(_33871_, _33872_, _33874_);
  xor g_64046_(_33869_, _33874_, _33875_);
  xor g_64047_(_32701_, _33875_, _33876_);
  xor g_64048_(_33867_, _33876_, _33877_);
  and g_64049_(_32716_, _32725_, _33878_);
  xor g_64050_(_33877_, _33878_, _33879_);
  and g_64051_(_32729_, _33879_, _33880_);
  and g_64052_(_31530_, _33879_, _33881_);
  not g_64053_(_33881_, _33882_);
  and g_64054_(_31528_, _32727_, _33883_);
  and g_64055_(_33882_, _33883_, _33885_);
  or g_64056_(_33880_, _33885_, _33886_);
  and g_64057_(_32733_, _32739_, _33887_);
  xor g_64058_(_33886_, _33887_, _33888_);
  xor g_64059_(_33866_, _33888_, _33889_);
  and g_64060_(_32630_, _32749_, _33890_);
  or g_64061_(_32748_, _33890_, _33891_);
  xor g_64062_(_33889_, _33891_, _33892_);
  xor g_64063_(_33864_, _33892_, _33893_);
  xor g_64064_(_33861_, _33893_, _33894_);
  xor g_64065_(_33860_, _33894_, _33896_);
  xor g_64066_(_33859_, _33896_, _33897_);
  xor g_64067_(_33857_, _33897_, _33898_);
  xor g_64068_(_33856_, _33898_, _33899_);
  xor g_64069_(_33854_, _33899_, _33900_);
  xor g_64070_(_33852_, _33900_, _33901_);
  or g_64071_(_31606_, _32816_, _33902_);
  and g_64072_(_32804_, _33902_, _33903_);
  and g_64073_(_32801_, _32811_, _33904_);
  xor g_64074_(_33903_, _33904_, _33905_);
  xor g_64075_(_33901_, _33905_, _33907_);
  xor g_64076_(_33849_, _33907_, _33908_);
  xor g_64077_(_33847_, _33908_, _33909_);
  and g_64078_(_32834_, _32844_, _33910_);
  xor g_64079_(_33909_, _33910_, _33911_);
  or g_64080_(_32613_, _32852_, _33912_);
  and g_64081_(_32850_, _33912_, _33913_);
  xor g_64082_(_33911_, _33913_, _33914_);
  xor g_64083_(_33846_, _33914_, _33915_);
  xor g_64084_(_32861_, _33915_, _33916_);
  xor g_64085_(_33844_, _33916_, _33918_);
  xor g_64086_(_33843_, _33918_, _33919_);
  xor g_64087_(_33841_, _33919_, _33920_);
  xor g_64088_(_33839_, _33920_, _33921_);
  xor g_64089_(_33837_, _33921_, _33922_);
  and g_64090_(_33835_, _33922_, _33923_);
  xor g_64091_(_33835_, _33922_, _33924_);
  not g_64092_(_33924_, _33925_);
  or g_64093_(_32911_, _33925_, _33926_);
  xor g_64094_(_32910_, _33924_, _33927_);
  xor g_64095_(_32911_, _33924_, _33929_);
  or g_64096_(_31688_, _32918_, _33930_);
  and g_64097_(_32913_, _33930_, _33931_);
  or g_64098_(_33929_, _33931_, _33932_);
  xor g_64099_(_33927_, _33931_, _33933_);
  and g_64100_(_33834_, _33933_, _33934_);
  or g_64101_(_33834_, _33933_, _33935_);
  xor g_64102_(_33834_, _33933_, _33936_);
  or g_64103_(_32922_, _32923_, _33937_);
  or g_64104_(_32927_, _32931_, _33938_);
  and g_64105_(_33937_, _33938_, _33940_);
  xor g_64106_(_33936_, _33940_, _33941_);
  or g_64107_(_33830_, _33941_, _33942_);
  and g_64108_(_33830_, _33941_, _33943_);
  xor g_64109_(_33830_, _33941_, _33944_);
  xor g_64110_(_33828_, _33944_, _33945_);
  or g_64111_(_33827_, _33945_, _33946_);
  xor g_64112_(_33827_, _33945_, _33947_);
  not g_64113_(_33947_, _33948_);
  or g_64114_(_33826_, _33948_, _33949_);
  xor g_64115_(_33826_, _33947_, _33951_);
  or g_64116_(_33825_, _33951_, _33952_);
  xor g_64117_(_33825_, _33951_, _33953_);
  and g_64118_(_33823_, _33953_, _33954_);
  or g_64119_(_33823_, _33953_, _33955_);
  xor g_64120_(_33822_, _33953_, _33956_);
  not g_64121_(_33956_, _33957_);
  and g_64122_(_30458_, _33821_, _33958_);
  or g_64123_(_32938_, _33958_, _33959_);
  xor g_64124_(_33956_, _33959_, _33960_);
  and g_64125_(_32942_, _33960_, _33962_);
  or g_64126_(_32942_, _33960_, _33963_);
  xor g_64127_(_32942_, _33960_, _33964_);
  not g_64128_(_33964_, _33965_);
  or g_64129_(_31721_, _32946_, _33966_);
  and g_64130_(_32945_, _33966_, _33967_);
  xor g_64131_(_33964_, _33967_, _33968_);
  not g_64132_(_33968_, _33969_);
  and g_64133_(_33819_, _33969_, _33970_);
  xor g_64134_(_33819_, _33969_, _33971_);
  xor g_64135_(_33819_, _33968_, _33973_);
  and g_64136_(_32957_, _33971_, _33974_);
  or g_64137_(_32956_, _33973_, _33975_);
  and g_64138_(_32953_, _33971_, _33976_);
  xor g_64139_(_32953_, _33973_, _33977_);
  and g_64140_(_32956_, _33977_, _33978_);
  or g_64141_(_33974_, _33978_, _33979_);
  xor g_64142_(_32960_, _33979_, _33980_);
  or g_64143_(_33817_, _33980_, _33981_);
  and g_64144_(_33817_, _33980_, _33982_);
  xor g_64145_(_33817_, _33980_, _33984_);
  and g_64146_(_32967_, _33984_, _33985_);
  and g_64147_(_31746_, _32964_, _33986_);
  or g_64148_(_31745_, _32963_, _33987_);
  xor g_64149_(_33984_, _33986_, _33988_);
  or g_64150_(_32967_, _33988_, _33989_);
  not g_64151_(_33989_, _33990_);
  or g_64152_(_33985_, _33990_, _33991_);
  xor g_64153_(_32970_, _33991_, _33992_);
  and g_64154_(_33816_, _33992_, _33993_);
  or g_64155_(_33816_, _33992_, _33995_);
  xor g_64156_(_33816_, _33992_, _33996_);
  xor g_64157_(_33815_, _33996_, _33997_);
  and g_64158_(_33813_, _33997_, _33998_);
  xor g_64159_(_33813_, _33997_, _33999_);
  xor g_64160_(_33814_, _33997_, _34000_);
  or g_64161_(_32981_, _34000_, _34001_);
  xor g_64162_(_32981_, _33999_, _34002_);
  or g_64163_(_32979_, _34002_, _34003_);
  xor g_64164_(_32980_, _34002_, _34004_);
  or g_64165_(_32986_, _34004_, _34006_);
  and g_64166_(_32986_, _34004_, _34007_);
  xor g_64167_(_32986_, _34004_, _34008_);
  xor g_64168_(_33812_, _34008_, _34009_);
  xor g_64169_(_33811_, _34009_, _34010_);
  xor g_64170_(_32991_, _34010_, _34011_);
  xor g_64171_(_32992_, _34010_, _34012_);
  and g_64172_(_33809_, _34011_, _34013_);
  or g_64173_(_33810_, _34012_, _34014_);
  and g_64174_(_33810_, _34012_, _34015_);
  or g_64175_(_33809_, _34011_, _34017_);
  or g_64176_(_33808_, _34015_, _34018_);
  and g_64177_(_34014_, _34018_, _34019_);
  or g_64178_(_34013_, _34018_, _34020_);
  and g_64179_(_33806_, _34020_, _34021_);
  and g_64180_(_34017_, _34019_, _34022_);
  or g_64181_(_34021_, _34022_, _34023_);
  or g_64182_(_33804_, _34023_, _34024_);
  xor g_64183_(_33804_, _34023_, _34025_);
  not g_64184_(_34025_, _34026_);
  or g_64185_(_33801_, _34026_, _34028_);
  xor g_64186_(_33801_, _34025_, _34029_);
  or g_64187_(_33012_, _34029_, _34030_);
  and g_64188_(_33012_, _34029_, _34031_);
  xor g_64189_(_33013_, _34029_, _34032_);
  or g_64190_(_31814_, _33017_, _34033_);
  and g_64191_(_33015_, _34033_, _34034_);
  not g_64192_(_34034_, _34035_);
  xor g_64193_(_34032_, _34035_, _34036_);
  and g_64194_(_31819_, _33023_, _34037_);
  or g_64195_(_33022_, _34037_, _34039_);
  not g_64196_(_34039_, _34040_);
  or g_64197_(_34036_, _34039_, _34041_);
  xor g_64198_(_34036_, _34039_, _34042_);
  xor g_64199_(_34036_, _34040_, _34043_);
  or g_64200_(_33800_, _34043_, _34044_);
  xor g_64201_(_33800_, _34042_, _34045_);
  or g_64202_(_33030_, _34045_, _34046_);
  xor g_64203_(_33030_, _34045_, _34047_);
  or g_64204_(_33032_, _34047_, _34048_);
  and g_64205_(_33032_, _34047_, _34050_);
  xor g_64206_(_33032_, _34047_, _34051_);
  or g_64207_(_31842_, _33037_, _34052_);
  and g_64208_(_33036_, _34052_, _34053_);
  not g_64209_(_34053_, _34054_);
  xor g_64210_(_34051_, _34054_, _34055_);
  not g_64211_(_34055_, _34056_);
  or g_64212_(_33046_, _34056_, _34057_);
  xor g_64213_(_33046_, _34055_, _34058_);
  or g_64214_(_33799_, _34058_, _34059_);
  xor g_64215_(_33799_, _34058_, _34061_);
  and g_64216_(_33057_, _34061_, _34062_);
  not g_64217_(_34062_, _34063_);
  and g_64218_(_33054_, _34061_, _34064_);
  xor g_64219_(_33054_, _34061_, _34065_);
  or g_64220_(_33057_, _34065_, _34066_);
  and g_64221_(_34063_, _34066_, _34067_);
  and g_64222_(_33063_, _34067_, _34068_);
  not g_64223_(_34068_, _34069_);
  xor g_64224_(_33061_, _34067_, _34070_);
  or g_64225_(_33063_, _34070_, _34072_);
  and g_64226_(_34069_, _34072_, _34073_);
  not g_64227_(_34073_, _34074_);
  xor g_64228_(_33065_, _34073_, _34075_);
  and g_64229_(_33069_, _34075_, _34076_);
  and g_64230_(_33070_, _34073_, _34077_);
  or g_64231_(_33069_, _34074_, _34078_);
  or g_64232_(_34076_, _34077_, _34079_);
  xor g_64233_(_33074_, _34079_, _34080_);
  and g_64234_(_33798_, _34080_, _34081_);
  xor g_64235_(_33798_, _34080_, _34083_);
  and g_64236_(_31877_, _33084_, _34084_);
  or g_64237_(_33083_, _34084_, _34085_);
  not g_64238_(_34085_, _34086_);
  and g_64239_(_34083_, _34086_, _34087_);
  xor g_64240_(_34083_, _34086_, _34088_);
  xor g_64241_(_34083_, _34085_, _34089_);
  or g_64242_(_33795_, _34089_, _34090_);
  and g_64243_(_33795_, _34089_, _34091_);
  xor g_64244_(_33795_, _34088_, _34092_);
  not g_64245_(_34092_, _34094_);
  or g_64246_(_32560_, _33091_, _34095_);
  and g_64247_(_33090_, _34095_, _34096_);
  xor g_64248_(_34092_, _34096_, _34097_);
  xor g_64249_(_34094_, _34096_, _34098_);
  or g_64250_(_33098_, _34098_, _34099_);
  xor g_64251_(_33098_, _34097_, _34100_);
  xor g_64252_(_33101_, _34100_, _34101_);
  xor g_64253_(_33794_, _34101_, _34102_);
  or g_64254_(_33791_, _34102_, _34103_);
  xor g_64255_(_33792_, _34102_, _34105_);
  or g_64256_(_33789_, _34105_, _34106_);
  xor g_64257_(_33789_, _34105_, _34107_);
  not g_64258_(_34107_, _34108_);
  or g_64259_(_33788_, _34108_, _34109_);
  xor g_64260_(_33788_, _34108_, _34110_);
  xor g_64261_(_33788_, _34107_, _34111_);
  and g_64262_(_33108_, _34110_, _34112_);
  xor g_64263_(_33107_, _34110_, _34113_);
  and g_64264_(_33111_, _34113_, _34114_);
  or g_64265_(_33111_, _34111_, _34116_);
  not g_64266_(_34116_, _34117_);
  or g_64267_(_34114_, _34117_, _34118_);
  not g_64268_(_34118_, _34119_);
  xor g_64269_(_33787_, _34119_, _34120_);
  xor g_64270_(_33787_, _34118_, _34121_);
  or g_64271_(_31918_, _33112_, _34122_);
  and g_64272_(_33117_, _34122_, _34123_);
  xor g_64273_(_34121_, _34123_, _34124_);
  or g_64274_(_33119_, _34124_, _34125_);
  xor g_64275_(_33120_, _34124_, _34127_);
  not g_64276_(_34127_, _34128_);
  and g_64277_(_33125_, _33127_, _34129_);
  or g_64278_(_34127_, _34129_, _34130_);
  xor g_64279_(_34127_, _34129_, _34131_);
  xor g_64280_(_34128_, _34129_, _34132_);
  or g_64281_(_33131_, _34132_, _34133_);
  xor g_64282_(_33131_, _34131_, _34134_);
  and g_64283_(_33784_, _34134_, _34135_);
  and g_64284_(_33786_, _34131_, _34136_);
  or g_64285_(_33784_, _34132_, _34138_);
  or g_64286_(_34135_, _34136_, _34139_);
  xor g_64287_(_33783_, _34139_, _34140_);
  not g_64288_(_34140_, _34141_);
  or g_64289_(_33136_, _34140_, _34142_);
  xor g_64290_(_33136_, _34141_, _34143_);
  or g_64291_(_33141_, _34143_, _34144_);
  or g_64292_(_33140_, _34141_, _34145_);
  and g_64293_(_34144_, _34145_, _34146_);
  xor g_64294_(_33143_, _34146_, _34147_);
  and g_64295_(_33147_, _34147_, _34149_);
  xor g_64296_(_33147_, _34147_, _34150_);
  and g_64297_(_33154_, _34150_, _34151_);
  xor g_64298_(_33154_, _34150_, _34152_);
  and g_64299_(_33157_, _34152_, _34153_);
  xor g_64300_(_33158_, _34152_, _34154_);
  and g_64301_(_33161_, _33164_, _34155_);
  or g_64302_(_34154_, _34155_, _34156_);
  xor g_64303_(_34154_, _34155_, _34157_);
  and g_64304_(_33167_, _34157_, _34158_);
  xor g_64305_(_33168_, _34157_, _34160_);
  not g_64306_(_34160_, _34161_);
  and g_64307_(_33172_, _34161_, _34162_);
  xor g_64308_(_33172_, _34160_, _34163_);
  or g_64309_(_33781_, _34163_, _34164_);
  xor g_64310_(_33781_, _34163_, _34165_);
  not g_64311_(_34165_, _34166_);
  or g_64312_(_33780_, _34166_, _34167_);
  xor g_64313_(_33780_, _34165_, _34168_);
  or g_64314_(_33779_, _34168_, _34169_);
  xor g_64315_(_33779_, _34168_, _34171_);
  or g_64316_(_33777_, _34171_, _34172_);
  and g_64317_(_33777_, _34171_, _34173_);
  xor g_64318_(_33778_, _34171_, _34174_);
  and g_64319_(_33185_, _33190_, _34175_);
  not g_64320_(_34175_, _34176_);
  xor g_64321_(_34174_, _34176_, _34177_);
  or g_64322_(_33776_, _34177_, _34178_);
  xor g_64323_(_33776_, _34177_, _34179_);
  or g_64324_(_33773_, _34179_, _34180_);
  and g_64325_(_33773_, _34179_, _34182_);
  xor g_64326_(_33775_, _34179_, _34183_);
  and g_64327_(_33196_, _33199_, _34184_);
  or g_64328_(_33197_, _33198_, _34185_);
  and g_64329_(_33202_, _34185_, _34186_);
  xor g_64330_(_34183_, _34186_, _34187_);
  not g_64331_(_34187_, _34188_);
  or g_64332_(_33206_, _34188_, _34189_);
  xor g_64333_(_33206_, _34187_, _34190_);
  and g_64334_(_32013_, _33209_, _34191_);
  or g_64335_(_33208_, _34191_, _34193_);
  or g_64336_(_34190_, _34193_, _34194_);
  xor g_64337_(_34190_, _34193_, _34195_);
  and g_64338_(_33771_, _34195_, _34196_);
  or g_64339_(_33771_, _34195_, _34197_);
  xor g_64340_(_33771_, _34195_, _34198_);
  xor g_64341_(_33772_, _34195_, _34199_);
  xor g_64342_(_33215_, _34199_, _34200_);
  or g_64343_(_33219_, _34200_, _34201_);
  or g_64344_(_33218_, _34198_, _34202_);
  and g_64345_(_34201_, _34202_, _34204_);
  not g_64346_(_34204_, _34205_);
  or g_64347_(_33224_, _34204_, _34206_);
  xor g_64348_(_33221_, _34205_, _34207_);
  xor g_64349_(_33221_, _34204_, _34208_);
  and g_64350_(_33224_, _34207_, _34209_);
  or g_64351_(_33226_, _34208_, _34210_);
  and g_64352_(_34206_, _34210_, _34211_);
  not g_64353_(_34211_, _34212_);
  and g_64354_(_33239_, _34211_, _34213_);
  or g_64355_(_33238_, _34212_, _34215_);
  xor g_64356_(_33228_, _34211_, _34216_);
  and g_64357_(_33238_, _34216_, _34217_);
  or g_64358_(_34213_, _34217_, _34218_);
  xor g_64359_(_33237_, _34218_, _34219_);
  or g_64360_(_33244_, _34219_, _34220_);
  and g_64361_(_33244_, _34219_, _34221_);
  xor g_64362_(_33244_, _34219_, _34222_);
  xor g_64363_(_33770_, _34222_, _34223_);
  or g_64364_(_33768_, _34223_, _34224_);
  xor g_64365_(_33769_, _34223_, _34226_);
  and g_64366_(_33251_, _34226_, _34227_);
  or g_64367_(_33251_, _34226_, _34228_);
  xor g_64368_(_33251_, _34226_, _34229_);
  xor g_64369_(_33254_, _34229_, _34230_);
  or g_64370_(_33767_, _34230_, _34231_);
  and g_64371_(_33767_, _34229_, _34232_);
  not g_64372_(_34232_, _34233_);
  and g_64373_(_34231_, _34233_, _34234_);
  xor g_64374_(_33765_, _34234_, _34235_);
  not g_64375_(_34235_, _34237_);
  or g_64376_(_33764_, _34235_, _34238_);
  xor g_64377_(_33764_, _34235_, _34239_);
  xor g_64378_(_33764_, _34237_, _34240_);
  or g_64379_(_33267_, _34240_, _34241_);
  xor g_64380_(_33267_, _34240_, _34242_);
  xor g_64381_(_33267_, _34239_, _34243_);
  and g_64382_(_33272_, _34243_, _34244_);
  or g_64383_(_33271_, _34242_, _34245_);
  and g_64384_(_33271_, _34239_, _34246_);
  not g_64385_(_34246_, _34248_);
  and g_64386_(_34245_, _34248_, _34249_);
  or g_64387_(_34244_, _34246_, _34250_);
  and g_64388_(_33762_, _34249_, _34251_);
  not g_64389_(_34251_, _34252_);
  and g_64390_(_33275_, _34249_, _34253_);
  and g_64391_(_33274_, _34250_, _34254_);
  or g_64392_(_33762_, _34254_, _34255_);
  or g_64393_(_34253_, _34255_, _34256_);
  and g_64394_(_34252_, _34256_, _34257_);
  xor g_64395_(_33759_, _34257_, _34259_);
  and g_64396_(_33756_, _34259_, _34260_);
  xor g_64397_(_33757_, _34259_, _34261_);
  and g_64398_(_33282_, _34261_, _34262_);
  or g_64399_(_33282_, _34261_, _34263_);
  xor g_64400_(_33282_, _34261_, _34264_);
  xor g_64401_(_33288_, _34264_, _34265_);
  or g_64402_(_33290_, _34265_, _34266_);
  and g_64403_(_33290_, _34265_, _34267_);
  xor g_64404_(_33290_, _34265_, _34268_);
  xor g_64405_(_33297_, _34268_, _34270_);
  and g_64406_(_32098_, _33295_, _34271_);
  or g_64407_(_33300_, _34271_, _34272_);
  not g_64408_(_34272_, _34273_);
  or g_64409_(_34270_, _34272_, _34274_);
  and g_64410_(_34270_, _34272_, _34275_);
  xor g_64411_(_34270_, _34272_, _34276_);
  xor g_64412_(_34270_, _34273_, _34277_);
  xor g_64413_(_33755_, _34277_, _34278_);
  xor g_64414_(_33755_, _34276_, _34279_);
  or g_64415_(_33307_, _34279_, _34281_);
  xor g_64416_(_33307_, _34278_, _34282_);
  or g_64417_(_33310_, _34282_, _34283_);
  xor g_64418_(_33311_, _34282_, _34284_);
  and g_64419_(_33314_, _33317_, _34285_);
  not g_64420_(_34285_, _34286_);
  or g_64421_(_34284_, _34285_, _34287_);
  xor g_64422_(_34284_, _34286_, _34288_);
  not g_64423_(_34288_, _34289_);
  or g_64424_(_33754_, _34288_, _34290_);
  xor g_64425_(_33754_, _34288_, _34292_);
  xor g_64426_(_33754_, _34289_, _34293_);
  or g_64427_(_33753_, _34293_, _34294_);
  xor g_64428_(_33753_, _34293_, _34295_);
  xor g_64429_(_33753_, _34292_, _34296_);
  and g_64430_(_33323_, _34295_, _34297_);
  xor g_64431_(_33323_, _34296_, _34298_);
  or g_64432_(_33327_, _34298_, _34299_);
  and g_64433_(_33327_, _34298_, _34300_);
  xor g_64434_(_33327_, _34298_, _34301_);
  xor g_64435_(_33329_, _34301_, _34303_);
  or g_64436_(_33331_, _34303_, _34304_);
  xor g_64437_(_33331_, _34303_, _34305_);
  and g_64438_(_32120_, _33333_, _34306_);
  or g_64439_(_32119_, _33334_, _34307_);
  and g_64440_(_33337_, _34307_, _34308_);
  or g_64441_(_33336_, _34306_, _34309_);
  and g_64442_(_34305_, _34309_, _34310_);
  xor g_64443_(_34305_, _34308_, _34311_);
  or g_64444_(_33751_, _34311_, _34312_);
  and g_64445_(_33751_, _34311_, _34314_);
  xor g_64446_(_33751_, _34311_, _34315_);
  xor g_64447_(_33342_, _34315_, _34316_);
  and g_64448_(_32134_, _33347_, _34317_);
  or g_64449_(_33345_, _34317_, _34318_);
  not g_64450_(_34318_, _34319_);
  or g_64451_(_34316_, _34318_, _34320_);
  xor g_64452_(_34316_, _34319_, _34321_);
  or g_64453_(_32140_, _33351_, _34322_);
  or g_64454_(_32138_, _33349_, _34323_);
  and g_64455_(_34322_, _34323_, _34325_);
  not g_64456_(_34325_, _34326_);
  or g_64457_(_34321_, _34325_, _34327_);
  xor g_64458_(_34321_, _34326_, _34328_);
  or g_64459_(_33749_, _34328_, _34329_);
  and g_64460_(_33749_, _34328_, _34330_);
  xor g_64461_(_33750_, _34328_, _34331_);
  xor g_64462_(_33361_, _34331_, _34332_);
  or g_64463_(_33354_, _34332_, _34333_);
  and g_64464_(_33354_, _34332_, _34334_);
  xor g_64465_(_33354_, _34332_, _34336_);
  xor g_64466_(_33364_, _34336_, _34337_);
  and g_64467_(_33374_, _34337_, _34338_);
  and g_64468_(_33367_, _34337_, _34339_);
  xor g_64469_(_33367_, _34337_, _34340_);
  or g_64470_(_33374_, _34340_, _34341_);
  not g_64471_(_34341_, _34342_);
  or g_64472_(_34338_, _34342_, _34343_);
  xor g_64473_(_33371_, _34343_, _34344_);
  or g_64474_(_33382_, _34344_, _34345_);
  xor g_64475_(_33382_, _34344_, _34347_);
  and g_64476_(_33378_, _34347_, _34348_);
  or g_64477_(_33378_, _34347_, _34349_);
  xor g_64478_(_33378_, _34347_, _34350_);
  xor g_64479_(_33386_, _34350_, _34351_);
  and g_64480_(_33394_, _34351_, _34352_);
  or g_64481_(_33394_, _34351_, _34353_);
  xor g_64482_(_33394_, _34351_, _34354_);
  xor g_64483_(_33389_, _34354_, _34355_);
  or g_64484_(_33748_, _34355_, _34356_);
  or g_64485_(_33399_, _34355_, _34358_);
  xor g_64486_(_33399_, _34355_, _34359_);
  or g_64487_(_33747_, _34359_, _34360_);
  and g_64488_(_34356_, _34360_, _34361_);
  not g_64489_(_34361_, _34362_);
  and g_64490_(_33746_, _34362_, _34363_);
  not g_64491_(_34363_, _34364_);
  or g_64492_(_33746_, _34355_, _34365_);
  and g_64493_(_34364_, _34365_, _34366_);
  xor g_64494_(_33405_, _34366_, _34367_);
  or g_64495_(_33744_, _34367_, _34369_);
  xor g_64496_(_33745_, _34367_, _34370_);
  or g_64497_(_33740_, _34370_, _34371_);
  and g_64498_(_33740_, _34370_, _34372_);
  xor g_64499_(_33742_, _34370_, _34373_);
  xor g_64500_(_33416_, _34373_, _34374_);
  and g_64501_(_33419_, _34374_, _34375_);
  xor g_64502_(_33419_, _34374_, _34376_);
  or g_64503_(_32198_, _33417_, _34377_);
  not g_64504_(_34377_, _34378_);
  and g_64505_(_34376_, _34378_, _34380_);
  xor g_64506_(_34376_, _34378_, _34381_);
  xor g_64507_(_34376_, _34377_, _34382_);
  or g_64508_(_33739_, _34382_, _34383_);
  xor g_64509_(_33739_, _34381_, _34384_);
  or g_64510_(_33431_, _34384_, _34385_);
  and g_64511_(_33431_, _34384_, _34386_);
  xor g_64512_(_33430_, _34384_, _34387_);
  xor g_64513_(_33428_, _34387_, _34388_);
  and g_64514_(_32213_, _33436_, _34389_);
  or g_64515_(_33435_, _34389_, _34391_);
  or g_64516_(_34388_, _34391_, _34392_);
  xor g_64517_(_34388_, _34391_, _34393_);
  and g_64518_(_32218_, _33437_, _34394_);
  or g_64519_(_33441_, _34394_, _34395_);
  and g_64520_(_34393_, _34395_, _34396_);
  xor g_64521_(_34393_, _34395_, _34397_);
  and g_64522_(_33443_, _34397_, _34398_);
  xor g_64523_(_33443_, _34397_, _34399_);
  xor g_64524_(_33446_, _34399_, _34400_);
  xor g_64525_(_33738_, _34400_, _34402_);
  or g_64526_(_33458_, _34402_, _34403_);
  not g_64527_(_34403_, _34404_);
  and g_64528_(_33458_, _34402_, _34405_);
  xor g_64529_(_33458_, _34402_, _34406_);
  xor g_64530_(_33469_, _34406_, _34407_);
  or g_64531_(_33471_, _34407_, _34408_);
  and g_64532_(_33471_, _34407_, _34409_);
  xor g_64533_(_33471_, _34407_, _34410_);
  xor g_64534_(_33736_, _34410_, _34411_);
  or g_64535_(_33735_, _34411_, _34413_);
  and g_64536_(_33735_, _34411_, _34414_);
  xor g_64537_(_33735_, _34411_, _34415_);
  not g_64538_(_34415_, _34416_);
  or g_64539_(_33488_, _34416_, _34417_);
  not g_64540_(_34417_, _34418_);
  and g_64541_(_33477_, _34415_, _34419_);
  not g_64542_(_34419_, _34420_);
  or g_64543_(_33477_, _34415_, _34421_);
  and g_64544_(_33488_, _34421_, _34422_);
  and g_64545_(_34420_, _34422_, _34424_);
  or g_64546_(_34418_, _34424_, _34425_);
  or g_64547_(_32265_, _33493_, _34426_);
  and g_64548_(_33481_, _34426_, _34427_);
  xor g_64549_(_34425_, _34427_, _34428_);
  and g_64550_(_33734_, _34428_, _34429_);
  xor g_64551_(_33734_, _34428_, _34430_);
  xor g_64552_(_33733_, _34428_, _34431_);
  and g_64553_(_33497_, _34430_, _34432_);
  or g_64554_(_33498_, _34431_, _34433_);
  and g_64555_(_33498_, _34431_, _34435_);
  or g_64556_(_33497_, _34430_, _34436_);
  and g_64557_(_34433_, _34436_, _34437_);
  or g_64558_(_34432_, _34435_, _34438_);
  or g_64559_(_32283_, _33510_, _34439_);
  not g_64560_(_34439_, _34440_);
  and g_64561_(_33513_, _34439_, _34441_);
  or g_64562_(_33512_, _34440_, _34442_);
  and g_64563_(_34438_, _34441_, _34443_);
  or g_64564_(_34437_, _34442_, _34444_);
  and g_64565_(_34436_, _34442_, _34446_);
  or g_64566_(_34435_, _34441_, _34447_);
  and g_64567_(_34433_, _34446_, _34448_);
  or g_64568_(_34432_, _34447_, _34449_);
  and g_64569_(_34444_, _34449_, _34450_);
  or g_64570_(_34443_, _34448_, _34451_);
  and g_64571_(_33729_, _34451_, _34452_);
  or g_64572_(_33729_, _34451_, _34453_);
  xor g_64573_(_33731_, _34450_, _34454_);
  and g_64574_(_33519_, _33523_, _34455_);
  not g_64575_(_34455_, _34457_);
  xor g_64576_(_34454_, _34457_, _34458_);
  and g_64577_(_33728_, _34458_, _34459_);
  xor g_64578_(_33727_, _34458_, _34460_);
  or g_64579_(_33726_, _34460_, _34461_);
  xor g_64580_(_33726_, _34460_, _34462_);
  not g_64581_(_34462_, _34463_);
  or g_64582_(_33530_, _34463_, _34464_);
  xor g_64583_(_33530_, _34462_, _34465_);
  or g_64584_(_33535_, _34465_, _34466_);
  xor g_64585_(_33535_, _34465_, _34468_);
  or g_64586_(_33532_, _34468_, _34469_);
  and g_64587_(_33532_, _34468_, _34470_);
  xor g_64588_(_33532_, _34468_, _34471_);
  xor g_64589_(_33724_, _34471_, _34472_);
  and g_64590_(_33722_, _34472_, _34473_);
  or g_64591_(_33722_, _34472_, _34474_);
  xor g_64592_(_33723_, _34472_, _34475_);
  xor g_64593_(_33721_, _34475_, _34476_);
  and g_64594_(_33720_, _34476_, _34477_);
  xor g_64595_(_33720_, _34476_, _34479_);
  not g_64596_(_34479_, _34480_);
  and g_64597_(_33542_, _34479_, _34481_);
  xor g_64598_(_33542_, _34479_, _34482_);
  not g_64599_(_34482_, _34483_);
  and g_64600_(_33717_, _34482_, _34484_);
  or g_64601_(_33718_, _34483_, _34485_);
  and g_64602_(_33546_, _34479_, _34486_);
  or g_64603_(_33547_, _34480_, _34487_);
  or g_64604_(_33546_, _34482_, _34488_);
  and g_64605_(_34487_, _34488_, _34490_);
  or g_64606_(_33717_, _34490_, _34491_);
  and g_64607_(_34485_, _34491_, _34492_);
  xor g_64608_(_33715_, _34492_, _34493_);
  or g_64609_(_33714_, _34493_, _34494_);
  not g_64610_(_34494_, _34495_);
  or g_64611_(_32354_, _33551_, _34496_);
  not g_64612_(_34496_, _34497_);
  or g_64613_(_34493_, _34496_, _34498_);
  xor g_64614_(_34493_, _34496_, _34499_);
  xor g_64615_(_34493_, _34497_, _34501_);
  and g_64616_(_33714_, _34501_, _34502_);
  or g_64617_(_33713_, _34499_, _34503_);
  and g_64618_(_34494_, _34503_, _34504_);
  or g_64619_(_34495_, _34502_, _34505_);
  and g_64620_(_33561_, _34504_, _34506_);
  or g_64621_(_33562_, _34505_, _34507_);
  xor g_64622_(_33558_, _34504_, _34508_);
  and g_64623_(_33562_, _34508_, _34509_);
  or g_64624_(_34506_, _34509_, _34510_);
  not g_64625_(_34510_, _34512_);
  and g_64626_(_33568_, _34512_, _34513_);
  or g_64627_(_33569_, _34510_, _34514_);
  xor g_64628_(_33564_, _34510_, _34515_);
  or g_64629_(_33568_, _34515_, _34516_);
  and g_64630_(_34514_, _34516_, _34517_);
  xor g_64631_(_33573_, _34517_, _34518_);
  and g_64632_(_33575_, _34518_, _34519_);
  not g_64633_(_34519_, _34520_);
  or g_64634_(_33575_, _34518_, _34521_);
  xor g_64635_(_33575_, _34518_, _34523_);
  or g_64636_(_32374_, _33579_, _34524_);
  or g_64637_(_34523_, _34524_, _34525_);
  not g_64638_(_34525_, _34526_);
  and g_64639_(_34521_, _34524_, _34527_);
  and g_64640_(_34520_, _34527_, _34528_);
  or g_64641_(_34526_, _34528_, _34529_);
  and g_64642_(_33712_, _34529_, _34530_);
  or g_64643_(_33712_, _34529_, _34531_);
  xor g_64644_(_33712_, _34529_, _34532_);
  xor g_64645_(_33587_, _34532_, _34534_);
  xor g_64646_(_33586_, _34532_, _34535_);
  and g_64647_(_33711_, _34535_, _34536_);
  xor g_64648_(_33710_, _34534_, _34537_);
  xor g_64649_(_33710_, _34535_, _34538_);
  and g_64650_(_33598_, _34538_, _34539_);
  not g_64651_(_34539_, _34540_);
  and g_64652_(_33595_, _34538_, _34541_);
  or g_64653_(_33596_, _34537_, _34542_);
  and g_64654_(_33596_, _34537_, _34543_);
  or g_64655_(_33598_, _34543_, _34545_);
  or g_64656_(_34541_, _34545_, _34546_);
  and g_64657_(_34540_, _34546_, _34547_);
  not g_64658_(_34547_, _34548_);
  and g_64659_(_33602_, _33605_, _34549_);
  or g_64660_(_34547_, _34549_, _34550_);
  xor g_64661_(_34547_, _34549_, _34551_);
  xor g_64662_(_34548_, _34549_, _34552_);
  or g_64663_(_33609_, _34552_, _34553_);
  xor g_64664_(_33609_, _34551_, _34554_);
  and g_64665_(_33709_, _34554_, _34556_);
  or g_64666_(_33709_, _34554_, _34557_);
  xor g_64667_(_33707_, _34554_, _34558_);
  xor g_64668_(_33706_, _34558_, _34559_);
  and g_64669_(_33617_, _34559_, _34560_);
  xor g_64670_(_33617_, _34559_, _34561_);
  or g_64671_(_33619_, _34561_, _34562_);
  and g_64672_(_33619_, _34559_, _34563_);
  not g_64673_(_34563_, _34564_);
  and g_64674_(_34562_, _34564_, _34565_);
  or g_64675_(_33625_, _34565_, _34567_);
  and g_64676_(_33625_, _34561_, _34568_);
  not g_64677_(_34568_, _34569_);
  and g_64678_(_34567_, _34569_, _34570_);
  xor g_64679_(_33705_, _34570_, _34571_);
  or g_64680_(_33704_, _34571_, _34572_);
  and g_64681_(_33704_, _34571_, _34573_);
  xor g_64682_(_33704_, _34571_, _34574_);
  xor g_64683_(_33703_, _34574_, _34575_);
  or g_64684_(_33698_, _34575_, _34576_);
  xor g_64685_(_33699_, _34575_, _34578_);
  or g_64686_(_33694_, _34578_, _34579_);
  xor g_64687_(_33695_, _34578_, _34580_);
  or g_64688_(_33693_, _34580_, _34581_);
  xor g_64689_(_33693_, _34580_, _34582_);
  xor g_64690_(_33637_, _34582_, _34583_);
  xor g_64691_(_33638_, _34582_, _34584_);
  and g_64692_(_33645_, _34584_, _34585_);
  or g_64693_(_33646_, _34583_, _34586_);
  and g_64694_(_33637_, _33641_, _34587_);
  not g_64695_(_34587_, _34589_);
  and g_64696_(_34582_, _34589_, _34590_);
  xor g_64697_(_34582_, _34587_, _34591_);
  and g_64698_(_33646_, _34591_, _34592_);
  not g_64699_(_34592_, _34593_);
  and g_64700_(_34586_, _34593_, _34594_);
  or g_64701_(_34585_, _34592_, _34595_);
  or g_64702_(_33653_, _34595_, _34596_);
  and g_64703_(_33649_, _34594_, _34597_);
  not g_64704_(_34597_, _34598_);
  and g_64705_(_33650_, _34595_, _34600_);
  or g_64706_(_33649_, _34594_, _34601_);
  and g_64707_(_33653_, _34601_, _34602_);
  or g_64708_(_33655_, _34600_, _34603_);
  and g_64709_(_34598_, _34602_, _34604_);
  or g_64710_(_34597_, _34603_, _34605_);
  and g_64711_(_34596_, _34605_, _34606_);
  xor g_64712_(_33692_, _34606_, _34607_);
  or g_64713_(_33690_, _34607_, _34608_);
  xor g_64714_(_33691_, _34607_, _34609_);
  or g_64715_(_33662_, _34609_, _34611_);
  xor g_64716_(_33661_, _34609_, _34612_);
  and g_64717_(_33689_, _34612_, _34613_);
  not g_64718_(_34613_, _34614_);
  or g_64719_(_33689_, _34612_, _34615_);
  not g_64720_(_34615_, _34616_);
  and g_64721_(_34614_, _34615_, _34617_);
  or g_64722_(_34613_, _34616_, _34618_);
  and g_64723_(_33688_, _34618_, _34619_);
  and g_64724_(_33687_, _34615_, _34620_);
  and g_64725_(_34614_, _34620_, _34622_);
  or g_64726_(_33667_, _34622_, _34623_);
  or g_64727_(_34619_, _34623_, _34624_);
  and g_64728_(_33667_, _34617_, _34625_);
  not g_64729_(_34625_, _34626_);
  and g_64730_(_34624_, _34626_, _34627_);
  xor g_64731_(_33670_, _34627_, _34628_);
  and g_64732_(_32479_, _33673_, _34629_);
  or g_64733_(_33674_, _34629_, _34630_);
  not g_64734_(_34630_, _34631_);
  and g_64735_(_34628_, _34631_, _34633_);
  xor g_64736_(_34628_, _34631_, _34634_);
  and g_64737_(_33683_, _34634_, _34635_);
  xor g_64738_(_33684_, _34634_, _34636_);
  and g_64739_(_33680_, _33682_, _34637_);
  or g_64740_(_34636_, _34637_, _34638_);
  xor g_64741_(_34636_, _34637_, out[646]);
  or g_64742_(_34633_, _34635_, _34639_);
  and g_64743_(_33670_, _34624_, _34640_);
  or g_64744_(_34625_, _34640_, _34641_);
  or g_64745_(_34613_, _34620_, _34643_);
  and g_64746_(_34608_, _34611_, _34644_);
  and g_64747_(_33692_, _34596_, _34645_);
  or g_64748_(_34604_, _34645_, _34646_);
  or g_64749_(_33649_, _34591_, _34647_);
  and g_64750_(_34586_, _34647_, _34648_);
  and g_64751_(_34579_, _34581_, _34649_);
  and g_64752_(_33702_, _34572_, _34650_);
  or g_64753_(_34573_, _34650_, _34651_);
  and g_64754_(_33705_, _34567_, _34652_);
  or g_64755_(_34568_, _34652_, _34654_);
  or g_64756_(_34560_, _34563_, _34655_);
  and g_64757_(_34550_, _34553_, _34656_);
  and g_64758_(_34542_, _34545_, _34657_);
  and g_64759_(_33586_, _34531_, _34658_);
  or g_64760_(_34530_, _34658_, _34659_);
  or g_64761_(_34519_, _34527_, _34660_);
  and g_64762_(_33574_, _34516_, _34661_);
  or g_64763_(_34513_, _34661_, _34662_);
  and g_64764_(_33564_, _34507_, _34663_);
  or g_64765_(_34509_, _34663_, _34665_);
  or g_64766_(_33558_, _34502_, _34666_);
  and g_64767_(_34494_, _34666_, _34667_);
  or g_64768_(_33716_, _34484_, _34668_);
  and g_64769_(_34491_, _34668_, _34669_);
  or g_64770_(_34477_, _34481_, _34670_);
  or g_64771_(_34486_, _34670_, _34671_);
  or g_64772_(_33721_, _34473_, _34672_);
  and g_64773_(_34474_, _34672_, _34673_);
  and g_64774_(_33725_, _34469_, _34674_);
  or g_64775_(_34470_, _34674_, _34676_);
  and g_64776_(_34464_, _34466_, _34677_);
  and g_64777_(_33524_, _34454_, _34678_);
  and g_64778_(_33519_, _34453_, _34679_);
  or g_64779_(_34452_, _34679_, _34680_);
  or g_64780_(_34432_, _34446_, _34681_);
  or g_64781_(_34425_, _34426_, _34682_);
  or g_64782_(_33481_, _34424_, _34683_);
  and g_64783_(_34417_, _34683_, _34684_);
  or g_64784_(_33736_, _34409_, _34685_);
  and g_64785_(_34408_, _34685_, _34687_);
  or g_64786_(_33469_, _34404_, _34688_);
  not g_64787_(_34688_, _34689_);
  or g_64788_(_34405_, _34689_, _34690_);
  or g_64789_(_33455_, _34400_, _34691_);
  or g_64790_(_33447_, _33450_, _34692_);
  and g_64791_(_34399_, _34692_, _34693_);
  or g_64792_(_34396_, _34398_, _34694_);
  or g_64793_(_34375_, _34380_, _34695_);
  or g_64794_(_33416_, _34372_, _34696_);
  and g_64795_(_34371_, _34696_, _34698_);
  and g_64796_(_34356_, _34358_, _34699_);
  and g_64797_(_33389_, _34353_, _34700_);
  or g_64798_(_34352_, _34700_, _34701_);
  or g_64799_(_33387_, _34348_, _34702_);
  and g_64800_(_34349_, _34702_, _34703_);
  and g_64801_(_33371_, _34341_, _34704_);
  or g_64802_(_34338_, _34704_, _34705_);
  or g_64803_(_33364_, _34334_, _34706_);
  and g_64804_(_34333_, _34706_, _34707_);
  or g_64805_(_33342_, _34314_, _34709_);
  and g_64806_(_34312_, _34709_, _34710_);
  or g_64807_(_33329_, _34300_, _34711_);
  and g_64808_(_34299_, _34711_, _34712_);
  and g_64809_(_34290_, _34294_, _34713_);
  and g_64810_(_34281_, _34283_, _34714_);
  and g_64811_(_33755_, _34274_, _34715_);
  or g_64812_(_34275_, _34715_, _34716_);
  or g_64813_(_33297_, _34267_, _34717_);
  and g_64814_(_34266_, _34717_, _34718_);
  or g_64815_(_33288_, _34262_, _34720_);
  and g_64816_(_34263_, _34720_, _34721_);
  and g_64817_(_33759_, _34256_, _34722_);
  or g_64818_(_34251_, _34722_, _34723_);
  and g_64819_(_33274_, _34245_, _34724_);
  or g_64820_(_34246_, _34724_, _34725_);
  and g_64821_(_33766_, _34231_, _34726_);
  or g_64822_(_34232_, _34726_, _34727_);
  or g_64823_(_33253_, _34227_, _34728_);
  and g_64824_(_34228_, _34728_, _34729_);
  or g_64825_(_33770_, _34221_, _34731_);
  and g_64826_(_34220_, _34731_, _34732_);
  or g_64827_(_33235_, _34217_, _34733_);
  and g_64828_(_34215_, _34733_, _34734_);
  and g_64829_(_33228_, _34206_, _34735_);
  or g_64830_(_34209_, _34735_, _34736_);
  and g_64831_(_33218_, _33221_, _34737_);
  or g_64832_(_34200_, _34737_, _34738_);
  and g_64833_(_33215_, _34197_, _34739_);
  or g_64834_(_34196_, _34739_, _34740_);
  and g_64835_(_34189_, _34194_, _34742_);
  or g_64836_(_33202_, _34183_, _34743_);
  or g_64837_(_34182_, _34184_, _34744_);
  and g_64838_(_34180_, _34744_, _34745_);
  or g_64839_(_33183_, _34173_, _34746_);
  and g_64840_(_34172_, _34746_, _34747_);
  and g_64841_(_34167_, _34169_, _34748_);
  or g_64842_(_34158_, _34162_, _34749_);
  or g_64843_(_34151_, _34153_, _34750_);
  or g_64844_(_33782_, _34135_, _34751_);
  and g_64845_(_34138_, _34751_, _34753_);
  or g_64846_(_33117_, _34120_, _34754_);
  and g_64847_(_34125_, _34754_, _34755_);
  or g_64848_(_34120_, _34122_, _34756_);
  and g_64849_(_34106_, _34109_, _34757_);
  and g_64850_(_33101_, _33794_, _34758_);
  or g_64851_(_34100_, _34758_, _34759_);
  or g_64852_(_33094_, _34092_, _34760_);
  and g_64853_(_33090_, _34090_, _34761_);
  or g_64854_(_34091_, _34761_, _34762_);
  or g_64855_(_34081_, _34087_, _34764_);
  or g_64856_(_33074_, _34076_, _34765_);
  and g_64857_(_34078_, _34765_, _34766_);
  and g_64858_(_33066_, _34072_, _34767_);
  or g_64859_(_34068_, _34767_, _34768_);
  and g_64860_(_33061_, _34066_, _34769_);
  or g_64861_(_34062_, _34769_, _34770_);
  and g_64862_(_34057_, _34059_, _34771_);
  and g_64863_(_34044_, _34046_, _34772_);
  and g_64864_(_33042_, _34051_, _34773_);
  xor g_64865_(_34772_, _34773_, _34775_);
  and g_64866_(_33035_, _34048_, _34776_);
  or g_64867_(_34050_, _34776_, _34777_);
  and g_64868_(_34024_, _34028_, _34778_);
  and g_64869_(_32991_, _33811_, _34779_);
  or g_64870_(_34009_, _34779_, _34780_);
  and g_64871_(_33815_, _33995_, _34781_);
  or g_64872_(_33993_, _34781_, _34782_);
  and g_64873_(_32971_, _33989_, _34783_);
  or g_64874_(_33985_, _34783_, _34784_);
  and g_64875_(_33981_, _33987_, _34786_);
  or g_64876_(_33982_, _34786_, _34787_);
  and g_64877_(_32962_, _33975_, _34788_);
  or g_64878_(_33978_, _34788_, _34789_);
  or g_64879_(_33970_, _33976_, _34790_);
  or g_64880_(_33965_, _33966_, _34791_);
  and g_64881_(_32938_, _33957_, _34792_);
  and g_64882_(_33955_, _33958_, _34793_);
  or g_64883_(_33954_, _34793_, _34794_);
  and g_64884_(_33949_, _33952_, _34795_);
  or g_64885_(_33828_, _33943_, _34797_);
  and g_64886_(_33942_, _34797_, _34798_);
  or g_64887_(_33934_, _33940_, _34799_);
  and g_64888_(_33935_, _34799_, _34800_);
  and g_64889_(_33926_, _33932_, _34801_);
  or g_64890_(_33923_, _34801_, _34802_);
  and g_64891_(_33923_, _33932_, _34803_);
  not g_64892_(_34803_, _34804_);
  and g_64893_(_34802_, _34804_, _34805_);
  xor g_64894_(_34800_, _34805_, _34806_);
  xor g_64895_(_34798_, _34806_, _34808_);
  xor g_64896_(_33946_, _34808_, _34809_);
  xor g_64897_(_34795_, _34809_, _34810_);
  xor g_64898_(_34794_, _34810_, _34811_);
  xor g_64899_(_34792_, _34811_, _34812_);
  or g_64900_(_32945_, _33962_, _34813_);
  and g_64901_(_33963_, _34813_, _34814_);
  xor g_64902_(_34812_, _34814_, _34815_);
  xor g_64903_(_34791_, _34815_, _34816_);
  xor g_64904_(_34790_, _34816_, _34817_);
  xor g_64905_(_34789_, _34817_, _34819_);
  xor g_64906_(_34787_, _34819_, _34820_);
  xor g_64907_(_34784_, _34820_, _34821_);
  xor g_64908_(_34782_, _34821_, _34822_);
  xor g_64909_(_33998_, _34822_, _34823_);
  xor g_64910_(_34001_, _34823_, _34824_);
  xor g_64911_(_34003_, _34824_, _34825_);
  or g_64912_(_33812_, _34007_, _34826_);
  and g_64913_(_34006_, _34826_, _34827_);
  xor g_64914_(_34825_, _34827_, _34828_);
  xor g_64915_(_34780_, _34828_, _34830_);
  xor g_64916_(_34019_, _34830_, _34831_);
  xor g_64917_(_34778_, _34831_, _34832_);
  or g_64918_(_33015_, _34031_, _34833_);
  and g_64919_(_34030_, _34833_, _34834_);
  xor g_64920_(_34832_, _34834_, _34835_);
  or g_64921_(_33020_, _34032_, _34836_);
  and g_64922_(_34041_, _34836_, _34837_);
  xor g_64923_(_34835_, _34837_, _34838_);
  xor g_64924_(_34777_, _34838_, _34839_);
  xor g_64925_(_34775_, _34839_, _34841_);
  xor g_64926_(_34771_, _34841_, _34842_);
  xor g_64927_(_34064_, _34842_, _34843_);
  xor g_64928_(_34770_, _34843_, _34844_);
  xor g_64929_(_34768_, _34844_, _34845_);
  xor g_64930_(_34766_, _34845_, _34846_);
  xor g_64931_(_34764_, _34846_, _34847_);
  xor g_64932_(_34762_, _34847_, _34848_);
  xor g_64933_(_34760_, _34848_, _34849_);
  xor g_64934_(_34099_, _34849_, _34850_);
  xor g_64935_(_34759_, _34850_, _34852_);
  xor g_64936_(_34103_, _34852_, _34853_);
  xor g_64937_(_34757_, _34853_, _34854_);
  xor g_64938_(_34112_, _34854_, _34855_);
  or g_64939_(_33787_, _34114_, _34856_);
  and g_64940_(_34116_, _34856_, _34857_);
  xor g_64941_(_34855_, _34857_, _34858_);
  xor g_64942_(_34756_, _34858_, _34859_);
  xor g_64943_(_34755_, _34859_, _34860_);
  xor g_64944_(_34130_, _34860_, _34861_);
  xor g_64945_(_34133_, _34861_, _34863_);
  xor g_64946_(_34753_, _34863_, _34864_);
  and g_64947_(_33140_, _33143_, _34865_);
  or g_64948_(_34143_, _34865_, _34866_);
  and g_64949_(_34142_, _34866_, _34867_);
  xor g_64950_(_34864_, _34867_, _34868_);
  xor g_64951_(_34149_, _34868_, _34869_);
  xor g_64952_(_34750_, _34869_, _34870_);
  xor g_64953_(_34156_, _34870_, _34871_);
  xor g_64954_(_34749_, _34871_, _34872_);
  xor g_64955_(_34164_, _34872_, _34874_);
  xor g_64956_(_34748_, _34874_, _34875_);
  xor g_64957_(_34747_, _34875_, _34876_);
  and g_64958_(_33182_, _33190_, _34877_);
  or g_64959_(_34174_, _34877_, _34878_);
  and g_64960_(_34178_, _34878_, _34879_);
  xor g_64961_(_34876_, _34879_, _34880_);
  xor g_64962_(_34745_, _34880_, _34881_);
  xor g_64963_(_34743_, _34881_, _34882_);
  xor g_64964_(_34742_, _34882_, _34883_);
  xor g_64965_(_34740_, _34883_, _34885_);
  xor g_64966_(_34738_, _34885_, _34886_);
  xor g_64967_(_34736_, _34886_, _34887_);
  xor g_64968_(_34734_, _34887_, _34888_);
  xor g_64969_(_34732_, _34888_, _34889_);
  xor g_64970_(_34224_, _34889_, _34890_);
  xor g_64971_(_34729_, _34890_, _34891_);
  xor g_64972_(_34727_, _34891_, _34892_);
  xor g_64973_(_34238_, _34892_, _34893_);
  xor g_64974_(_34241_, _34893_, _34894_);
  xor g_64975_(_34725_, _34894_, _34896_);
  xor g_64976_(_34723_, _34896_, _34897_);
  xor g_64977_(_34260_, _34897_, _34898_);
  xor g_64978_(_34721_, _34898_, _34899_);
  xor g_64979_(_34718_, _34899_, _34900_);
  xor g_64980_(_34716_, _34900_, _34901_);
  xor g_64981_(_34714_, _34901_, _34902_);
  xor g_64982_(_34287_, _34902_, _34903_);
  xor g_64983_(_34713_, _34903_, _34904_);
  xor g_64984_(_34297_, _34904_, _34905_);
  xor g_64985_(_34712_, _34905_, _34907_);
  xor g_64986_(_34304_, _34907_, _34908_);
  xor g_64987_(_34310_, _34908_, _34909_);
  xor g_64988_(_34710_, _34909_, _34910_);
  and g_64989_(_34320_, _34327_, _34911_);
  or g_64990_(_33361_, _34330_, _34912_);
  and g_64991_(_34329_, _34912_, _34913_);
  xor g_64992_(_34911_, _34913_, _34914_);
  xor g_64993_(_34910_, _34914_, _34915_);
  xor g_64994_(_34707_, _34915_, _34916_);
  xor g_64995_(_34339_, _34916_, _34918_);
  xor g_64996_(_34705_, _34918_, _34919_);
  xor g_64997_(_34345_, _34919_, _34920_);
  xor g_64998_(_34703_, _34920_, _34921_);
  xor g_64999_(_34701_, _34921_, _34922_);
  xor g_65000_(_34699_, _34922_, _34923_);
  and g_65001_(_33405_, _34365_, _34924_);
  or g_65002_(_34363_, _34924_, _34925_);
  xor g_65003_(_34369_, _34925_, _34926_);
  xor g_65004_(_34923_, _34926_, _34927_);
  xor g_65005_(_34698_, _34927_, _34929_);
  xor g_65006_(_34695_, _34929_, _34930_);
  xor g_65007_(_34383_, _34930_, _34931_);
  or g_65008_(_33429_, _34386_, _34932_);
  and g_65009_(_34385_, _34932_, _34933_);
  xor g_65010_(_34931_, _34933_, _34934_);
  xor g_65011_(_34392_, _34934_, _34935_);
  xor g_65012_(_34694_, _34935_, _34936_);
  xor g_65013_(_34693_, _34936_, _34937_);
  xor g_65014_(_34691_, _34937_, _34938_);
  xor g_65015_(_34690_, _34938_, _34940_);
  xor g_65016_(_34687_, _34940_, _34941_);
  or g_65017_(_33477_, _34414_, _34942_);
  and g_65018_(_34413_, _34942_, _34943_);
  xor g_65019_(_34941_, _34943_, _34944_);
  xor g_65020_(_34684_, _34944_, _34945_);
  xor g_65021_(_34682_, _34945_, _34946_);
  xor g_65022_(_34429_, _34946_, _34947_);
  xor g_65023_(_34681_, _34947_, _34948_);
  xor g_65024_(_34680_, _34948_, _34949_);
  xor g_65025_(_34678_, _34949_, _34951_);
  xor g_65026_(_34459_, _34951_, _34952_);
  xor g_65027_(_34461_, _34952_, _34953_);
  xor g_65028_(_34677_, _34953_, _34954_);
  xor g_65029_(_34676_, _34954_, _34955_);
  xor g_65030_(_34673_, _34955_, _34956_);
  xor g_65031_(_34671_, _34956_, _34957_);
  xor g_65032_(_34669_, _34957_, _34958_);
  xor g_65033_(_34498_, _34958_, _34959_);
  xor g_65034_(_34667_, _34959_, _34960_);
  xor g_65035_(_34665_, _34960_, _34962_);
  xor g_65036_(_34662_, _34962_, _34963_);
  xor g_65037_(_34660_, _34963_, _34964_);
  xor g_65038_(_34659_, _34964_, _34965_);
  xor g_65039_(_34536_, _34965_, _34966_);
  xor g_65040_(_34657_, _34966_, _34967_);
  xor g_65041_(_34656_, _34967_, _34968_);
  or g_65042_(_33706_, _34556_, _34969_);
  and g_65043_(_34557_, _34969_, _34970_);
  xor g_65044_(_34968_, _34970_, _34971_);
  xor g_65045_(_34655_, _34971_, _34973_);
  xor g_65046_(_34654_, _34973_, _34974_);
  xor g_65047_(_34651_, _34974_, _34975_);
  xor g_65048_(_34576_, _34975_, _34976_);
  xor g_65049_(_34649_, _34976_, _34977_);
  xor g_65050_(_34590_, _34977_, _34978_);
  xor g_65051_(_34648_, _34978_, _34979_);
  xor g_65052_(_34646_, _34979_, _34980_);
  xor g_65053_(_34644_, _34980_, _34981_);
  xor g_65054_(_34643_, _34981_, _34982_);
  xor g_65055_(_34641_, _34982_, _34984_);
  xor g_65056_(_34639_, _34984_, _34985_);
  xor g_65057_(_34638_, _34985_, out[647]);
  buf b_0_(set1[16], out[336]);
  buf b_1_(set1[236], out[556]);
  buf b_2_(set2[96], out[96]);
  buf b_3_(set1[83], out[403]);
  buf b_4_(set1[89], out[409]);
  buf b_5_(set1[32], out[352]);
  buf b_6_(set1[187], out[507]);
  buf b_7_(set1[192], out[512]);
  buf b_8_(set1[149], out[469]);
  buf b_9_(set1[210], out[530]);
  buf b_10_(set1[74], out[394]);
  buf b_11_(set2[8], out[8]);
  buf b_12_(set2[293], out[293]);
  buf b_13_(set2[173], out[173]);
  buf b_14_(set2[2], out[2]);
  buf b_15_(set1[229], out[549]);
  buf b_16_(set1[203], out[523]);
  buf b_17_(set2[84], out[84]);
  buf b_18_(set1[208], out[528]);
  buf b_19_(set2[197], out[197]);
  buf b_20_(set1[268], out[588]);
  buf b_21_(set1[13], out[333]);
  buf b_22_(set1[59], out[379]);
  buf b_23_(set2[125], out[125]);
  buf b_24_(set2[238], out[238]);
  buf b_25_(set1[305], out[625]);
  buf b_26_(set1[297], out[617]);
  buf b_27_(set1[176], out[496]);
  buf b_28_(set1[116], out[436]);
  buf b_29_(set2[62], out[62]);
  buf b_30_(set2[272], out[272]);
  buf b_31_(set1[53], out[373]);
  buf b_32_(set2[1], out[1]);
  buf b_33_(set1[272], out[592]);
  buf b_34_(set2[160], out[160]);
  buf b_35_(set2[203], out[203]);
  buf b_36_(set2[95], out[95]);
  buf b_37_(set1[247], out[567]);
  buf b_38_(set1[121], out[441]);
  buf b_39_(set1[278], out[598]);
  buf b_40_(set2[6], out[6]);
  buf b_41_(set1[61], out[381]);
  buf b_42_(set2[101], out[101]);
  buf b_43_(set2[318], out[318]);
  buf b_44_(set2[130], out[130]);
  buf b_45_(set1[174], out[494]);
  buf b_46_(set1[310], out[630]);
  buf b_47_(set1[46], out[366]);
  buf b_48_(set2[91], out[91]);
  buf b_49_(set2[186], out[186]);
  buf b_50_(set2[260], out[260]);
  buf b_51_(set1[287], out[607]);
  buf b_52_(set1[237], out[557]);
  buf b_53_(set1[10], out[330]);
  buf b_54_(set2[19], out[19]);
  buf b_55_(set2[176], out[176]);
  buf b_56_(set2[75], out[75]);
  buf b_57_(set2[16], out[16]);
  buf b_58_(set2[282], out[282]);
  buf b_59_(set1[25], out[345]);
  buf b_60_(set2[283], out[283]);
  buf b_61_(set1[199], out[519]);
  buf b_62_(set1[180], out[500]);
  buf b_63_(set2[123], out[123]);
  buf b_64_(set1[110], out[430]);
  buf b_65_(set1[201], out[521]);
  buf b_66_(set1[8], out[328]);
  buf b_67_(set1[289], out[609]);
  buf b_68_(set1[154], out[474]);
  buf b_69_(set1[148], out[468]);
  buf b_70_(set1[280], out[600]);
  buf b_71_(set1[298], out[618]);
  buf b_72_(set1[197], out[517]);
  buf b_73_(set2[247], out[247]);
  buf b_74_(set1[266], out[586]);
  buf b_75_(set1[14], out[334]);
  buf b_76_(set1[193], out[513]);
  buf b_77_(set2[134], out[134]);
  buf b_78_(set1[168], out[488]);
  buf b_79_(set2[33], out[33]);
  buf b_80_(set1[233], out[553]);
  buf b_81_(set1[250], out[570]);
  buf b_82_(set2[194], out[194]);
  buf b_83_(set2[26], out[26]);
  buf b_84_(set1[99], out[419]);
  buf b_85_(set2[222], out[222]);
  buf b_86_(set1[196], out[516]);
  buf b_87_(set2[154], out[154]);
  buf b_88_(set2[126], out[126]);
  buf b_89_(set2[199], out[199]);
  buf b_90_(set1[293], out[613]);
  buf b_91_(set1[246], out[566]);
  buf b_92_(set1[317], out[637]);
  buf b_93_(set2[7], out[7]);
  buf b_94_(set1[101], out[421]);
  buf b_95_(set1[173], out[493]);
  buf b_96_(set1[274], out[594]);
  buf b_97_(set2[40], out[40]);
  buf b_98_(set1[43], out[363]);
  buf b_99_(set2[70], out[70]);
  buf b_100_(set1[105], out[425]);
  buf b_101_(set2[202], out[202]);
  buf b_102_(set1[270], out[590]);
  buf b_103_(set2[147], out[147]);
  buf b_104_(set1[33], out[353]);
  buf b_105_(set1[302], out[622]);
  buf b_106_(set2[259], out[259]);
  buf b_107_(set1[189], out[509]);
  buf b_108_(set1[241], out[561]);
  buf b_109_(set2[139], out[139]);
  buf b_110_(set1[67], out[387]);
  buf b_111_(set2[48], out[48]);
  buf b_112_(set2[77], out[77]);
  buf b_113_(set1[273], out[593]);
  buf b_114_(set2[56], out[56]);
  buf b_115_(set1[2], out[322]);
  buf b_116_(set1[151], out[471]);
  buf b_117_(set2[265], out[265]);
  buf b_118_(set2[122], out[122]);
  buf b_119_(set2[28], out[28]);
  buf b_120_(set1[172], out[492]);
  buf b_121_(set1[31], out[351]);
  buf b_122_(set2[217], out[217]);
  buf b_123_(set1[0], out[320]);
  buf b_124_(set2[234], out[234]);
  buf b_125_(set2[220], out[220]);
  buf b_126_(set1[143], out[463]);
  buf b_127_(set1[198], out[518]);
  buf b_128_(set2[97], out[97]);
  buf b_129_(set2[67], out[67]);
  buf b_130_(set1[249], out[569]);
  buf b_131_(set2[214], out[214]);
  buf b_132_(set2[221], out[221]);
  buf b_133_(set1[97], out[417]);
  buf b_134_(set2[142], out[142]);
  buf b_135_(set1[69], out[389]);
  buf b_136_(set1[122], out[442]);
  buf b_137_(set2[10], out[10]);
  buf b_138_(set2[307], out[307]);
  buf b_139_(set1[158], out[478]);
  buf b_140_(set1[87], out[407]);
  buf b_141_(set1[19], out[339]);
  buf b_142_(set2[37], out[37]);
  buf b_143_(set1[29], out[349]);
  buf b_144_(set1[37], out[357]);
  buf b_145_(set1[161], out[481]);
  buf b_146_(set1[66], out[386]);
  buf b_147_(set2[213], out[213]);
  buf b_148_(set1[75], out[395]);
  buf b_149_(set2[49], out[49]);
  buf b_150_(set1[186], out[506]);
  buf b_151_(set1[243], out[563]);
  buf b_152_(set1[256], out[576]);
  buf b_153_(set1[221], out[541]);
  buf b_154_(set2[105], out[105]);
  buf b_155_(set1[160], out[480]);
  buf b_156_(set2[74], out[74]);
  buf b_157_(set2[11], out[11]);
  buf b_158_(set1[79], out[399]);
  buf b_159_(set2[86], out[86]);
  buf b_160_(set1[182], out[502]);
  buf b_161_(set2[58], out[58]);
  buf b_162_(set1[294], out[614]);
  buf b_163_(set1[82], out[402]);
  buf b_164_(set2[157], out[157]);
  buf b_165_(set1[77], out[397]);
  buf b_166_(set1[24], out[344]);
  buf b_167_(set1[52], out[372]);
  buf b_168_(set2[137], out[137]);
  buf b_169_(set2[188], out[188]);
  buf b_170_(set2[291], out[291]);
  buf b_171_(set2[136], out[136]);
  buf b_172_(set1[138], out[458]);
  buf b_173_(set2[79], out[79]);
  buf b_174_(set2[177], out[177]);
  buf b_175_(set2[5], out[5]);
  buf b_176_(set2[195], out[195]);
  buf b_177_(set2[280], out[280]);
  buf b_178_(set2[191], out[191]);
  buf b_179_(set1[164], out[484]);
  buf b_180_(set2[78], out[78]);
  buf b_181_(set1[130], out[450]);
  buf b_182_(set1[42], out[362]);
  buf b_183_(set2[216], out[216]);
  buf b_184_(set2[120], out[120]);
  buf b_185_(set1[240], out[560]);
  buf b_186_(set1[146], out[466]);
  buf b_187_(set1[106], out[426]);
  buf b_188_(set2[35], out[35]);
  buf b_189_(set1[222], out[542]);
  buf b_190_(set2[66], out[66]);
  buf b_191_(set2[218], out[218]);
  buf b_192_(set2[183], out[183]);
  buf b_193_(set2[76], out[76]);
  buf b_194_(set2[290], out[290]);
  buf b_195_(set2[106], out[106]);
  buf b_196_(set1[21], out[341]);
  buf b_197_(set2[179], out[179]);
  buf b_198_(set2[0], out[0]);
  buf b_199_(set1[60], out[380]);
  buf b_200_(set1[184], out[504]);
  buf b_201_(set2[192], out[192]);
  buf b_202_(set1[288], out[608]);
  buf b_203_(set2[207], out[207]);
  buf b_204_(set1[284], out[604]);
  buf b_205_(set2[243], out[243]);
  buf b_206_(set1[141], out[461]);
  buf b_207_(set1[26], out[346]);
  buf b_208_(set1[23], out[343]);
  buf b_209_(set2[145], out[145]);
  buf b_210_(set2[21], out[21]);
  buf b_211_(set1[163], out[483]);
  buf b_212_(set2[9], out[9]);
  buf b_213_(set1[132], out[452]);
  buf b_214_(set2[289], out[289]);
  buf b_215_(set2[187], out[187]);
  buf b_216_(set1[185], out[505]);
  buf b_217_(set2[23], out[23]);
  buf b_218_(set1[114], out[434]);
  buf b_219_(set1[27], out[347]);
  buf b_220_(set2[275], out[275]);
  buf b_221_(set1[118], out[438]);
  buf b_222_(set2[317], out[317]);
  buf b_223_(set2[132], out[132]);
  buf b_224_(set2[273], out[273]);
  buf b_225_(set1[126], out[446]);
  buf b_226_(set1[167], out[487]);
  buf b_227_(set2[248], out[248]);
  buf b_228_(set2[205], out[205]);
  buf b_229_(set2[146], out[146]);
  buf b_230_(set2[242], out[242]);
  buf b_231_(set1[157], out[477]);
  buf b_232_(set2[287], out[287]);
  buf b_233_(set1[142], out[462]);
  buf b_234_(set2[198], out[198]);
  buf b_235_(set2[211], out[211]);
  buf b_236_(set1[4], out[324]);
  buf b_237_(set1[57], out[377]);
  buf b_238_(set1[145], out[465]);
  buf b_239_(set1[311], out[631]);
  buf b_240_(set2[210], out[210]);
  buf b_241_(set1[245], out[565]);
  buf b_242_(set2[72], out[72]);
  buf b_243_(set2[215], out[215]);
  buf b_244_(set2[85], out[85]);
  buf b_245_(set1[314], out[634]);
  buf b_246_(set1[51], out[371]);
  buf b_247_(set1[152], out[472]);
  buf b_248_(set1[307], out[627]);
  buf b_249_(set1[205], out[525]);
  buf b_250_(set1[1], out[321]);
  buf b_251_(set1[251], out[571]);
  buf b_252_(set2[90], out[90]);
  buf b_253_(set2[309], out[309]);
  buf b_254_(set2[231], out[231]);
  buf b_255_(set2[219], out[219]);
  buf b_256_(set1[153], out[473]);
  buf b_257_(set2[174], out[174]);
  buf b_258_(set1[36], out[356]);
  buf b_259_(set1[178], out[498]);
  buf b_260_(set2[261], out[261]);
  buf b_261_(set1[226], out[546]);
  buf b_262_(set2[201], out[201]);
  buf b_263_(set1[188], out[508]);
  buf b_264_(set1[107], out[427]);
  buf b_265_(set2[153], out[153]);
  buf b_266_(set1[104], out[424]);
  buf b_267_(set2[271], out[271]);
  buf b_268_(set1[228], out[548]);
  buf b_269_(set1[85], out[405]);
  buf b_270_(set2[94], out[94]);
  buf b_271_(set1[177], out[497]);
  buf b_272_(set2[31], out[31]);
  buf b_273_(set2[249], out[249]);
  buf b_274_(set2[257], out[257]);
  buf b_275_(set2[232], out[232]);
  buf b_276_(set2[117], out[117]);
  buf b_277_(set2[165], out[165]);
  buf b_278_(set1[296], out[616]);
  buf b_279_(set2[241], out[241]);
  buf b_280_(set1[80], out[400]);
  buf b_281_(set2[20], out[20]);
  buf b_282_(set1[109], out[429]);
  buf b_283_(set1[211], out[531]);
  buf b_284_(set1[252], out[572]);
  buf b_285_(set1[235], out[555]);
  buf b_286_(set2[223], out[223]);
  buf b_287_(set1[119], out[439]);
  buf b_288_(set2[111], out[111]);
  buf b_289_(set2[171], out[171]);
  buf b_290_(set2[29], out[29]);
  buf b_291_(set2[180], out[180]);
  buf b_292_(set1[253], out[573]);
  buf b_293_(set2[38], out[38]);
  buf b_294_(set1[72], out[392]);
  buf b_295_(set1[219], out[539]);
  buf b_296_(set2[69], out[69]);
  buf b_297_(set1[238], out[558]);
  buf b_298_(set2[233], out[233]);
  buf b_299_(set1[18], out[338]);
  buf b_300_(set2[254], out[254]);
  buf b_301_(set1[300], out[620]);
  buf b_302_(set2[12], out[12]);
  buf b_303_(set2[140], out[140]);
  buf b_304_(set2[112], out[112]);
  buf b_305_(set1[98], out[418]);
  buf b_306_(set1[86], out[406]);
  buf b_307_(set2[109], out[109]);
  buf b_308_(set1[166], out[486]);
  buf b_309_(set1[195], out[515]);
  buf b_310_(set2[108], out[108]);
  buf b_311_(set1[303], out[623]);
  buf b_312_(set2[301], out[301]);
  buf b_313_(set2[305], out[305]);
  buf b_314_(set2[288], out[288]);
  buf b_315_(set2[274], out[274]);
  buf b_316_(set2[292], out[292]);
  buf b_317_(set1[102], out[422]);
  buf b_318_(set2[107], out[107]);
  buf b_319_(set2[189], out[189]);
  buf b_320_(set1[136], out[456]);
  buf b_321_(set1[55], out[375]);
  buf b_322_(set2[4], out[4]);
  buf b_323_(set1[123], out[443]);
  buf b_324_(set2[151], out[151]);
  buf b_325_(set2[267], out[267]);
  buf b_326_(set1[214], out[534]);
  buf b_327_(set1[115], out[435]);
  buf b_328_(set1[7], out[327]);
  buf b_329_(set2[299], out[299]);
  buf b_330_(set2[59], out[59]);
  buf b_331_(set1[30], out[350]);
  buf b_332_(set2[286], out[286]);
  buf b_333_(set2[319], out[319]);
  buf b_334_(set1[11], out[331]);
  buf b_335_(set2[68], out[68]);
  buf b_336_(set2[279], out[279]);
  buf b_337_(set1[56], out[376]);
  buf b_338_(set2[181], out[181]);
  buf b_339_(set2[81], out[81]);
  buf b_340_(set2[206], out[206]);
  buf b_341_(set1[34], out[354]);
  buf b_342_(set1[81], out[401]);
  buf b_343_(set2[270], out[270]);
  buf b_344_(set2[295], out[295]);
  buf b_345_(set1[282], out[602]);
  buf b_346_(set1[48], out[368]);
  buf b_347_(set1[234], out[554]);
  buf b_348_(set1[54], out[374]);
  buf b_349_(set1[84], out[404]);
  buf b_350_(set2[22], out[22]);
  buf b_351_(set1[230], out[550]);
  buf b_352_(set1[15], out[335]);
  buf b_353_(set2[196], out[196]);
  buf b_354_(set2[235], out[235]);
  buf b_355_(set1[58], out[378]);
  buf b_356_(set1[262], out[582]);
  buf b_357_(set1[108], out[428]);
  buf b_358_(set1[275], out[595]);
  buf b_359_(set2[30], out[30]);
  buf b_360_(set2[266], out[266]);
  buf b_361_(set1[204], out[524]);
  buf b_362_(set2[298], out[298]);
  buf b_363_(set1[242], out[562]);
  buf b_364_(set2[264], out[264]);
  buf b_365_(set2[3], out[3]);
  buf b_366_(set1[22], out[342]);
  buf b_367_(set1[181], out[501]);
  buf b_368_(set1[73], out[393]);
  buf b_369_(set2[277], out[277]);
  buf b_370_(set1[92], out[412]);
  buf b_371_(set1[50], out[370]);
  buf b_372_(set2[306], out[306]);
  buf b_373_(set2[212], out[212]);
  buf b_374_(set1[68], out[388]);
  buf b_375_(set2[312], out[312]);
  buf b_376_(set1[169], out[489]);
  buf b_377_(set1[183], out[503]);
  buf b_378_(set1[231], out[551]);
  buf b_379_(set1[291], out[611]);
  buf b_380_(set1[227], out[547]);
  buf b_381_(set2[226], out[226]);
  buf b_382_(set2[46], out[46]);
  buf b_383_(set2[100], out[100]);
  buf b_384_(set2[164], out[164]);
  buf b_385_(set2[71], out[71]);
  buf b_386_(set2[315], out[315]);
  buf b_387_(set1[120], out[440]);
  buf b_388_(set1[147], out[467]);
  buf b_389_(set2[115], out[115]);
  buf b_390_(set1[9], out[329]);
  buf b_391_(set2[303], out[303]);
  buf b_392_(set2[159], out[159]);
  buf b_393_(set1[313], out[633]);
  buf b_394_(set2[162], out[162]);
  buf b_395_(set1[304], out[624]);
  buf b_396_(set2[281], out[281]);
  buf b_397_(set1[47], out[367]);
  buf b_398_(set2[73], out[73]);
  buf b_399_(set1[129], out[449]);
  buf b_400_(set2[113], out[113]);
  buf b_401_(set2[65], out[65]);
  buf b_402_(set2[161], out[161]);
  buf b_403_(set1[103], out[423]);
  buf b_404_(set2[155], out[155]);
  buf b_405_(set1[283], out[603]);
  buf b_406_(set1[135], out[455]);
  buf b_407_(set2[163], out[163]);
  buf b_408_(set1[41], out[361]);
  buf b_409_(set2[253], out[253]);
  buf b_410_(set1[315], out[635]);
  buf b_411_(set2[294], out[294]);
  buf b_412_(set1[95], out[415]);
  buf b_413_(set1[260], out[580]);
  buf b_414_(set1[206], out[526]);
  buf b_415_(set1[318], out[638]);
  buf b_416_(set2[184], out[184]);
  buf b_417_(set1[3], out[323]);
  buf b_418_(set2[172], out[172]);
  buf b_419_(set2[64], out[64]);
  buf b_420_(set1[209], out[529]);
  buf b_421_(set1[90], out[410]);
  buf b_422_(set2[103], out[103]);
  buf b_423_(set2[83], out[83]);
  buf b_424_(set2[310], out[310]);
  buf b_425_(set1[281], out[601]);
  buf b_426_(set2[193], out[193]);
  buf b_427_(set1[111], out[431]);
  buf b_428_(set2[239], out[239]);
  buf b_429_(set2[209], out[209]);
  buf b_430_(set1[117], out[437]);
  buf b_431_(set1[261], out[581]);
  buf b_432_(set2[190], out[190]);
  buf b_433_(set2[169], out[169]);
  buf b_434_(set1[78], out[398]);
  buf b_435_(set2[55], out[55]);
  buf b_436_(set2[53], out[53]);
  buf b_437_(set2[240], out[240]);
  buf b_438_(set1[218], out[538]);
  buf b_439_(set2[224], out[224]);
  buf b_440_(set2[44], out[44]);
  buf b_441_(set2[263], out[263]);
  buf b_442_(set2[237], out[237]);
  buf b_443_(set1[213], out[533]);
  buf b_444_(set1[265], out[585]);
  buf b_445_(set1[88], out[408]);
  buf b_446_(set1[76], out[396]);
  buf b_447_(set1[264], out[584]);
  buf b_448_(set2[54], out[54]);
  buf b_449_(set1[215], out[535]);
  buf b_450_(set2[27], out[27]);
  buf b_451_(set2[276], out[276]);
  buf b_452_(set2[278], out[278]);
  buf b_453_(set2[297], out[297]);
  buf b_454_(set2[230], out[230]);
  buf b_455_(set1[12], out[332]);
  buf b_456_(set2[296], out[296]);
  buf b_457_(set1[171], out[491]);
  buf b_458_(set2[143], out[143]);
  buf b_459_(set2[314], out[314]);
  buf b_460_(set1[194], out[514]);
  buf b_461_(set1[128], out[448]);
  buf b_462_(set2[87], out[87]);
  buf b_463_(set2[41], out[41]);
  buf b_464_(set1[306], out[626]);
  buf b_465_(set1[257], out[577]);
  buf b_466_(set1[179], out[499]);
  buf b_467_(set2[128], out[128]);
  buf b_468_(set1[277], out[597]);
  buf b_469_(set1[225], out[545]);
  buf b_470_(set1[159], out[479]);
  buf b_471_(set1[165], out[485]);
  buf b_472_(set2[150], out[150]);
  buf b_473_(set1[62], out[382]);
  buf b_474_(set2[149], out[149]);
  buf b_475_(set2[138], out[138]);
  buf b_476_(set1[39], out[359]);
  buf b_477_(set2[135], out[135]);
  buf b_478_(set1[239], out[559]);
  buf b_479_(set2[127], out[127]);
  buf b_480_(set1[28], out[348]);
  buf b_481_(set2[63], out[63]);
  buf b_482_(set2[13], out[13]);
  buf b_483_(set2[229], out[229]);
  buf b_484_(set2[285], out[285]);
  buf b_485_(set2[47], out[47]);
  buf b_486_(set2[102], out[102]);
  buf b_487_(set2[185], out[185]);
  buf b_488_(set1[212], out[532]);
  buf b_489_(set1[267], out[587]);
  buf b_490_(set1[191], out[511]);
  buf b_491_(set1[125], out[445]);
  buf b_492_(set2[51], out[51]);
  buf b_493_(set2[110], out[110]);
  buf b_494_(set1[96], out[416]);
  buf b_495_(set2[227], out[227]);
  buf b_496_(set2[114], out[114]);
  buf b_497_(set1[309], out[629]);
  buf b_498_(set2[131], out[131]);
  buf b_499_(set1[279], out[599]);
  buf b_500_(set2[178], out[178]);
  buf b_501_(set1[49], out[369]);
  buf b_502_(set1[144], out[464]);
  buf b_503_(set2[98], out[98]);
  buf b_504_(set1[276], out[596]);
  buf b_505_(set2[302], out[302]);
  buf b_506_(set2[15], out[15]);
  buf b_507_(set1[162], out[482]);
  buf b_508_(set1[137], out[457]);
  buf b_509_(set2[208], out[208]);
  buf b_510_(set2[119], out[119]);
  buf b_511_(set2[182], out[182]);
  buf b_512_(set1[127], out[447]);
  buf b_513_(set1[224], out[544]);
  buf b_514_(set2[50], out[50]);
  buf b_515_(set1[170], out[490]);
  buf b_516_(set2[141], out[141]);
  buf b_517_(set1[113], out[433]);
  buf b_518_(set1[316], out[636]);
  buf b_519_(set2[116], out[116]);
  buf b_520_(set2[255], out[255]);
  buf b_521_(set2[118], out[118]);
  buf b_522_(set1[190], out[510]);
  buf b_523_(set1[232], out[552]);
  buf b_524_(set1[295], out[615]);
  buf b_525_(set1[258], out[578]);
  buf b_526_(set2[39], out[39]);
  buf b_527_(set2[80], out[80]);
  buf b_528_(set1[150], out[470]);
  buf b_529_(set1[45], out[365]);
  buf b_530_(set1[286], out[606]);
  buf b_531_(set1[202], out[522]);
  buf b_532_(set1[20], out[340]);
  buf b_533_(set2[89], out[89]);
  buf b_534_(set1[290], out[610]);
  buf b_535_(set1[216], out[536]);
  buf b_536_(set1[17], out[337]);
  buf b_537_(set2[269], out[269]);
  buf b_538_(set2[158], out[158]);
  buf b_539_(set2[313], out[313]);
  buf b_540_(set1[200], out[520]);
  buf b_541_(set1[5], out[325]);
  buf b_542_(set1[93], out[413]);
  buf b_543_(set1[271], out[591]);
  buf b_544_(set2[34], out[34]);
  buf b_545_(set1[131], out[451]);
  buf b_546_(set1[223], out[543]);
  buf b_547_(set2[316], out[316]);
  buf b_548_(set2[93], out[93]);
  buf b_549_(set1[255], out[575]);
  buf b_550_(set2[268], out[268]);
  buf b_551_(set2[236], out[236]);
  buf b_552_(set2[36], out[36]);
  buf b_553_(set2[200], out[200]);
  buf b_554_(set1[263], out[583]);
  buf b_555_(set2[82], out[82]);
  buf b_556_(set2[88], out[88]);
  buf b_557_(set1[63], out[383]);
  buf b_558_(set1[285], out[605]);
  buf b_559_(set1[319], out[639]);
  buf b_560_(set2[170], out[170]);
  buf b_561_(set1[100], out[420]);
  buf b_562_(set1[64], out[384]);
  buf b_563_(set1[44], out[364]);
  buf b_564_(set1[94], out[414]);
  buf b_565_(set2[124], out[124]);
  buf b_566_(set1[156], out[476]);
  buf b_567_(set1[155], out[475]);
  buf b_568_(set2[225], out[225]);
  buf b_569_(set2[152], out[152]);
  buf b_570_(set2[18], out[18]);
  buf b_571_(set1[244], out[564]);
  buf b_572_(set2[244], out[244]);
  buf b_573_(set2[32], out[32]);
  buf b_574_(set1[124], out[444]);
  buf b_575_(set2[92], out[92]);
  buf b_576_(set1[65], out[385]);
  buf b_577_(set1[91], out[411]);
  buf b_578_(set2[52], out[52]);
  buf b_579_(set2[245], out[245]);
  buf b_580_(set2[14], out[14]);
  buf b_581_(set1[40], out[360]);
  buf b_582_(set2[168], out[168]);
  buf b_583_(set1[140], out[460]);
  buf b_584_(set2[99], out[99]);
  buf b_585_(set1[70], out[390]);
  buf b_586_(set1[292], out[612]);
  buf b_587_(set2[60], out[60]);
  buf b_588_(set2[144], out[144]);
  buf b_589_(set1[217], out[537]);
  buf b_590_(set2[252], out[252]);
  buf b_591_(set1[139], out[459]);
  buf b_592_(set1[134], out[454]);
  buf b_593_(set2[121], out[121]);
  buf b_594_(set2[133], out[133]);
  buf b_595_(set1[207], out[527]);
  buf b_596_(set1[308], out[628]);
  buf b_597_(set2[148], out[148]);
  buf b_598_(set1[259], out[579]);
  buf b_599_(set1[301], out[621]);
  buf b_600_(set2[24], out[24]);
  buf b_601_(set2[308], out[308]);
  buf b_602_(set2[258], out[258]);
  buf b_603_(set1[71], out[391]);
  buf b_604_(set2[166], out[166]);
  buf b_605_(set2[262], out[262]);
  buf b_606_(set1[248], out[568]);
  buf b_607_(set2[129], out[129]);
  buf b_608_(set2[61], out[61]);
  buf b_609_(set2[228], out[228]);
  buf b_610_(set2[304], out[304]);
  buf b_611_(set2[167], out[167]);
  buf b_612_(set2[42], out[42]);
  buf b_613_(set2[25], out[25]);
  buf b_614_(set1[220], out[540]);
  buf b_615_(set1[112], out[432]);
  buf b_616_(set2[43], out[43]);
  buf b_617_(set1[254], out[574]);
  buf b_618_(set2[156], out[156]);
  buf b_619_(set2[204], out[204]);
  buf b_620_(set1[133], out[453]);
  buf b_621_(set1[175], out[495]);
  buf b_622_(set1[312], out[632]);
  buf b_623_(set2[45], out[45]);
  buf b_624_(set2[175], out[175]);
  buf b_625_(set2[17], out[17]);
  buf b_626_(set2[104], out[104]);
  buf b_627_(set2[284], out[284]);
  buf b_628_(set1[6], out[326]);
  buf b_629_(set2[311], out[311]);
  buf b_630_(set2[256], out[256]);
  buf b_631_(set1[269], out[589]);
  buf b_632_(set2[246], out[246]);
  buf b_633_(set1[35], out[355]);
  buf b_634_(set2[250], out[250]);
  buf b_635_(set1[299], out[619]);
  buf b_636_(set1[38], out[358]);
  buf b_637_(set2[57], out[57]);
  buf b_638_(set2[300], out[300]);
  buf b_639_(set2[251], out[251]);

endmodule
