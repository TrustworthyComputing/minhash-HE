module min_hash(
  input wire [479:0] set1,
  input wire [479:0] set2,
  output wire [975:0] out
);
  wire [15:0] set1_unflattened[30];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  wire [15:0] set2_unflattened[30];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  wire [15:0] array_index_512818;
  wire [15:0] array_index_512819;
  wire [11:0] add_512826;
  wire [11:0] add_512829;
  wire [15:0] array_index_512834;
  wire [15:0] array_index_512837;
  wire [10:0] add_512841;
  wire [10:0] add_512844;
  wire [11:0] add_512860;
  wire [11:0] sel_512862;
  wire [11:0] add_512865;
  wire [11:0] sel_512867;
  wire [15:0] array_index_512880;
  wire [15:0] array_index_512883;
  wire [10:0] add_512887;
  wire [10:0] add_512889;
  wire [10:0] add_512891;
  wire [11:0] sel_512894;
  wire [10:0] add_512896;
  wire [11:0] sel_512899;
  wire [11:0] add_512916;
  wire [11:0] sel_512918;
  wire [11:0] add_512921;
  wire [11:0] sel_512923;
  wire [15:0] array_index_512942;
  wire [15:0] array_index_512945;
  wire [10:0] add_512949;
  wire [10:0] add_512951;
  wire [10:0] add_512953;
  wire [11:0] sel_512955;
  wire [10:0] add_512957;
  wire [11:0] sel_512959;
  wire [10:0] add_512961;
  wire [11:0] sel_512964;
  wire [10:0] add_512966;
  wire [11:0] sel_512969;
  wire [11:0] add_512990;
  wire [11:0] sel_512992;
  wire [11:0] add_512995;
  wire [11:0] sel_512997;
  wire [15:0] array_index_513022;
  wire [15:0] array_index_513025;
  wire [11:0] add_513029;
  wire [11:0] add_513031;
  wire [10:0] add_513033;
  wire [11:0] sel_513035;
  wire [10:0] add_513037;
  wire [11:0] sel_513039;
  wire [10:0] add_513041;
  wire [11:0] sel_513043;
  wire [10:0] add_513045;
  wire [11:0] sel_513047;
  wire [10:0] add_513049;
  wire [11:0] sel_513052;
  wire [10:0] add_513054;
  wire [11:0] sel_513057;
  wire [11:0] add_513082;
  wire [11:0] sel_513084;
  wire [11:0] add_513087;
  wire [11:0] sel_513089;
  wire [15:0] array_index_513120;
  wire [15:0] array_index_513123;
  wire [7:0] add_513127;
  wire [7:0] add_513130;
  wire [11:0] add_513133;
  wire [11:0] sel_513135;
  wire [11:0] add_513137;
  wire [11:0] sel_513139;
  wire [10:0] add_513141;
  wire [11:0] sel_513143;
  wire [10:0] add_513145;
  wire [11:0] sel_513147;
  wire [10:0] add_513149;
  wire [11:0] sel_513151;
  wire [10:0] add_513153;
  wire [11:0] sel_513155;
  wire [10:0] add_513157;
  wire [11:0] sel_513160;
  wire [10:0] add_513162;
  wire [11:0] sel_513165;
  wire [11:0] add_513194;
  wire [11:0] sel_513196;
  wire [11:0] add_513199;
  wire [11:0] sel_513201;
  wire [15:0] array_index_513238;
  wire [15:0] array_index_513241;
  wire [11:0] add_513245;
  wire [11:0] add_513247;
  wire [7:0] add_513249;
  wire [11:0] sel_513252;
  wire [7:0] add_513254;
  wire [11:0] sel_513257;
  wire [11:0] add_513259;
  wire [11:0] sel_513261;
  wire [11:0] add_513263;
  wire [11:0] sel_513265;
  wire [10:0] add_513267;
  wire [11:0] sel_513269;
  wire [10:0] add_513271;
  wire [11:0] sel_513273;
  wire [10:0] add_513275;
  wire [11:0] sel_513277;
  wire [10:0] add_513279;
  wire [11:0] sel_513281;
  wire [10:0] add_513283;
  wire [11:0] sel_513286;
  wire [10:0] add_513288;
  wire [11:0] sel_513291;
  wire [11:0] add_513324;
  wire [11:0] sel_513326;
  wire [11:0] add_513329;
  wire [11:0] sel_513331;
  wire [15:0] array_index_513374;
  wire [15:0] array_index_513377;
  wire [9:0] add_513381;
  wire [9:0] add_513384;
  wire [11:0] add_513387;
  wire [11:0] sel_513389;
  wire [11:0] add_513391;
  wire [11:0] sel_513393;
  wire [7:0] add_513395;
  wire [11:0] sel_513398;
  wire [7:0] add_513400;
  wire [11:0] sel_513403;
  wire [11:0] add_513405;
  wire [11:0] sel_513407;
  wire [11:0] add_513409;
  wire [11:0] sel_513411;
  wire [10:0] add_513413;
  wire [11:0] sel_513415;
  wire [10:0] add_513417;
  wire [11:0] sel_513419;
  wire [10:0] add_513421;
  wire [11:0] sel_513423;
  wire [10:0] add_513425;
  wire [11:0] sel_513427;
  wire [10:0] add_513429;
  wire [11:0] sel_513432;
  wire [10:0] add_513434;
  wire [11:0] sel_513437;
  wire [11:0] add_513474;
  wire [11:0] sel_513476;
  wire [11:0] add_513479;
  wire [11:0] sel_513481;
  wire [15:0] array_index_513530;
  wire [15:0] array_index_513533;
  wire [11:0] add_513537;
  wire [11:0] add_513539;
  wire [9:0] add_513541;
  wire [11:0] sel_513544;
  wire [9:0] add_513546;
  wire [11:0] sel_513549;
  wire [11:0] add_513551;
  wire [11:0] sel_513553;
  wire [11:0] add_513555;
  wire [11:0] sel_513557;
  wire [7:0] add_513559;
  wire [11:0] sel_513562;
  wire [7:0] add_513564;
  wire [11:0] sel_513567;
  wire [11:0] add_513569;
  wire [11:0] sel_513571;
  wire [11:0] add_513573;
  wire [11:0] sel_513575;
  wire [10:0] add_513577;
  wire [11:0] sel_513579;
  wire [10:0] add_513581;
  wire [11:0] sel_513583;
  wire [10:0] add_513585;
  wire [11:0] sel_513587;
  wire [10:0] add_513589;
  wire [11:0] sel_513591;
  wire [10:0] add_513593;
  wire [11:0] sel_513596;
  wire [10:0] add_513598;
  wire [11:0] sel_513601;
  wire [11:0] add_513642;
  wire [11:0] sel_513644;
  wire [11:0] add_513647;
  wire [11:0] sel_513649;
  wire [15:0] array_index_513702;
  wire [15:0] array_index_513705;
  wire [11:0] add_513709;
  wire [11:0] add_513711;
  wire [11:0] add_513713;
  wire [11:0] sel_513715;
  wire [11:0] add_513717;
  wire [11:0] sel_513719;
  wire [9:0] add_513721;
  wire [11:0] sel_513724;
  wire [9:0] add_513726;
  wire [11:0] sel_513729;
  wire [11:0] add_513731;
  wire [11:0] sel_513733;
  wire [11:0] add_513735;
  wire [11:0] sel_513737;
  wire [7:0] add_513739;
  wire [11:0] sel_513742;
  wire [7:0] add_513744;
  wire [11:0] sel_513747;
  wire [11:0] add_513749;
  wire [11:0] sel_513751;
  wire [11:0] add_513753;
  wire [11:0] sel_513755;
  wire [10:0] add_513757;
  wire [11:0] sel_513759;
  wire [10:0] add_513761;
  wire [11:0] sel_513763;
  wire [10:0] add_513765;
  wire [11:0] sel_513767;
  wire [10:0] add_513769;
  wire [11:0] sel_513771;
  wire [10:0] add_513773;
  wire [11:0] sel_513776;
  wire [10:0] add_513778;
  wire [11:0] sel_513781;
  wire [11:0] add_513826;
  wire [11:0] sel_513828;
  wire [11:0] add_513831;
  wire [11:0] sel_513833;
  wire [15:0] array_index_513890;
  wire [15:0] array_index_513893;
  wire [10:0] add_513897;
  wire [10:0] add_513899;
  wire [11:0] add_513901;
  wire [11:0] sel_513903;
  wire [11:0] add_513905;
  wire [11:0] sel_513907;
  wire [11:0] add_513909;
  wire [11:0] sel_513911;
  wire [11:0] add_513913;
  wire [11:0] sel_513915;
  wire [9:0] add_513917;
  wire [11:0] sel_513920;
  wire [9:0] add_513922;
  wire [11:0] sel_513925;
  wire [11:0] add_513927;
  wire [11:0] sel_513929;
  wire [11:0] add_513931;
  wire [11:0] sel_513933;
  wire [7:0] add_513935;
  wire [11:0] sel_513938;
  wire [7:0] add_513940;
  wire [11:0] sel_513943;
  wire [11:0] add_513945;
  wire [11:0] sel_513947;
  wire [11:0] add_513949;
  wire [11:0] sel_513951;
  wire [10:0] add_513953;
  wire [11:0] sel_513955;
  wire [10:0] add_513957;
  wire [11:0] sel_513959;
  wire [10:0] add_513961;
  wire [11:0] sel_513963;
  wire [10:0] add_513965;
  wire [11:0] sel_513967;
  wire [10:0] add_513969;
  wire [11:0] sel_513972;
  wire [10:0] add_513974;
  wire [11:0] sel_513977;
  wire [11:0] add_514026;
  wire [11:0] sel_514028;
  wire [11:0] add_514031;
  wire [11:0] sel_514033;
  wire [15:0] array_index_514096;
  wire [15:0] array_index_514099;
  wire [11:0] add_514103;
  wire [11:0] add_514105;
  wire [10:0] add_514107;
  wire [11:0] sel_514109;
  wire [10:0] add_514111;
  wire [11:0] sel_514113;
  wire [11:0] add_514115;
  wire [11:0] sel_514117;
  wire [11:0] add_514119;
  wire [11:0] sel_514121;
  wire [11:0] add_514123;
  wire [11:0] sel_514125;
  wire [11:0] add_514127;
  wire [11:0] sel_514129;
  wire [9:0] add_514131;
  wire [11:0] sel_514134;
  wire [9:0] add_514136;
  wire [11:0] sel_514139;
  wire [11:0] add_514141;
  wire [11:0] sel_514143;
  wire [11:0] add_514145;
  wire [11:0] sel_514147;
  wire [7:0] add_514149;
  wire [11:0] sel_514152;
  wire [7:0] add_514154;
  wire [11:0] sel_514157;
  wire [11:0] add_514159;
  wire [11:0] sel_514161;
  wire [11:0] add_514163;
  wire [11:0] sel_514165;
  wire [10:0] add_514167;
  wire [11:0] sel_514169;
  wire [10:0] add_514171;
  wire [11:0] sel_514173;
  wire [10:0] add_514175;
  wire [11:0] sel_514177;
  wire [10:0] add_514179;
  wire [11:0] sel_514181;
  wire [10:0] add_514183;
  wire [11:0] sel_514186;
  wire [10:0] add_514188;
  wire [11:0] sel_514191;
  wire [11:0] add_514244;
  wire [11:0] sel_514246;
  wire [11:0] add_514249;
  wire [11:0] sel_514251;
  wire [15:0] array_index_514318;
  wire [15:0] array_index_514321;
  wire [9:0] add_514325;
  wire [9:0] add_514327;
  wire [11:0] add_514329;
  wire [11:0] sel_514331;
  wire [11:0] add_514333;
  wire [11:0] sel_514335;
  wire [10:0] add_514337;
  wire [11:0] sel_514339;
  wire [10:0] add_514341;
  wire [11:0] sel_514343;
  wire [11:0] add_514345;
  wire [11:0] sel_514347;
  wire [11:0] add_514349;
  wire [11:0] sel_514351;
  wire [11:0] add_514353;
  wire [11:0] sel_514355;
  wire [11:0] add_514357;
  wire [11:0] sel_514359;
  wire [9:0] add_514361;
  wire [11:0] sel_514364;
  wire [9:0] add_514366;
  wire [11:0] sel_514369;
  wire [11:0] add_514371;
  wire [11:0] sel_514373;
  wire [11:0] add_514375;
  wire [11:0] sel_514377;
  wire [7:0] add_514379;
  wire [11:0] sel_514382;
  wire [7:0] add_514384;
  wire [11:0] sel_514387;
  wire [11:0] add_514389;
  wire [11:0] sel_514391;
  wire [11:0] add_514393;
  wire [11:0] sel_514395;
  wire [10:0] add_514397;
  wire [11:0] sel_514399;
  wire [10:0] add_514401;
  wire [11:0] sel_514403;
  wire [10:0] add_514405;
  wire [11:0] sel_514407;
  wire [10:0] add_514409;
  wire [11:0] sel_514411;
  wire [10:0] add_514413;
  wire [11:0] sel_514416;
  wire [10:0] add_514418;
  wire [11:0] sel_514421;
  wire [11:0] add_514478;
  wire [11:0] sel_514480;
  wire [11:0] add_514483;
  wire [11:0] sel_514485;
  wire [15:0] array_index_514558;
  wire [15:0] array_index_514561;
  wire [10:0] add_514565;
  wire [10:0] add_514567;
  wire [9:0] add_514569;
  wire [11:0] sel_514571;
  wire [9:0] add_514573;
  wire [11:0] sel_514575;
  wire [11:0] add_514577;
  wire [11:0] sel_514579;
  wire [11:0] add_514581;
  wire [11:0] sel_514583;
  wire [10:0] add_514585;
  wire [11:0] sel_514587;
  wire [10:0] add_514589;
  wire [11:0] sel_514591;
  wire [11:0] add_514593;
  wire [11:0] sel_514595;
  wire [11:0] add_514597;
  wire [11:0] sel_514599;
  wire [11:0] add_514601;
  wire [11:0] sel_514603;
  wire [11:0] add_514605;
  wire [11:0] sel_514607;
  wire [9:0] add_514609;
  wire [11:0] sel_514612;
  wire [9:0] add_514614;
  wire [11:0] sel_514617;
  wire [11:0] add_514619;
  wire [11:0] sel_514621;
  wire [11:0] add_514623;
  wire [11:0] sel_514625;
  wire [7:0] add_514627;
  wire [11:0] sel_514630;
  wire [7:0] add_514632;
  wire [11:0] sel_514635;
  wire [11:0] add_514637;
  wire [11:0] sel_514639;
  wire [11:0] add_514641;
  wire [11:0] sel_514643;
  wire [10:0] add_514645;
  wire [11:0] sel_514647;
  wire [10:0] add_514649;
  wire [11:0] sel_514651;
  wire [10:0] add_514653;
  wire [11:0] sel_514655;
  wire [10:0] add_514657;
  wire [11:0] sel_514659;
  wire [10:0] add_514661;
  wire [11:0] sel_514664;
  wire [10:0] add_514666;
  wire [11:0] sel_514669;
  wire [11:0] add_514730;
  wire [11:0] sel_514732;
  wire [11:0] add_514735;
  wire [11:0] sel_514737;
  wire [15:0] array_index_514818;
  wire [15:0] array_index_514821;
  wire [8:0] add_514825;
  wire [8:0] add_514828;
  wire [10:0] add_514831;
  wire [11:0] sel_514833;
  wire [10:0] add_514835;
  wire [11:0] sel_514837;
  wire [9:0] add_514839;
  wire [11:0] sel_514841;
  wire [9:0] add_514843;
  wire [11:0] sel_514845;
  wire [11:0] add_514847;
  wire [11:0] sel_514849;
  wire [11:0] add_514851;
  wire [11:0] sel_514853;
  wire [10:0] add_514855;
  wire [11:0] sel_514857;
  wire [10:0] add_514859;
  wire [11:0] sel_514861;
  wire [11:0] add_514863;
  wire [11:0] sel_514865;
  wire [11:0] add_514867;
  wire [11:0] sel_514869;
  wire [11:0] add_514871;
  wire [11:0] sel_514873;
  wire [11:0] add_514875;
  wire [11:0] sel_514877;
  wire [9:0] add_514879;
  wire [11:0] sel_514882;
  wire [9:0] add_514884;
  wire [11:0] sel_514887;
  wire [11:0] add_514889;
  wire [11:0] sel_514891;
  wire [11:0] add_514893;
  wire [11:0] sel_514895;
  wire [7:0] add_514897;
  wire [11:0] sel_514900;
  wire [7:0] add_514902;
  wire [11:0] sel_514905;
  wire [11:0] add_514907;
  wire [11:0] sel_514909;
  wire [11:0] add_514911;
  wire [11:0] sel_514913;
  wire [10:0] add_514915;
  wire [11:0] sel_514917;
  wire [10:0] add_514919;
  wire [11:0] sel_514921;
  wire [10:0] add_514923;
  wire [11:0] sel_514925;
  wire [10:0] add_514927;
  wire [11:0] sel_514929;
  wire [10:0] add_514931;
  wire [11:0] sel_514934;
  wire [10:0] add_514936;
  wire [11:0] sel_514939;
  wire [11:0] add_515004;
  wire [11:0] sel_515006;
  wire [11:0] add_515009;
  wire [11:0] sel_515011;
  wire [15:0] array_index_515098;
  wire [15:0] array_index_515101;
  wire [11:0] add_515105;
  wire [11:0] add_515107;
  wire [8:0] add_515109;
  wire [11:0] sel_515112;
  wire [8:0] add_515114;
  wire [11:0] sel_515117;
  wire [10:0] add_515119;
  wire [11:0] sel_515121;
  wire [10:0] add_515123;
  wire [11:0] sel_515125;
  wire [9:0] add_515127;
  wire [11:0] sel_515129;
  wire [9:0] add_515131;
  wire [11:0] sel_515133;
  wire [11:0] add_515135;
  wire [11:0] sel_515137;
  wire [11:0] add_515139;
  wire [11:0] sel_515141;
  wire [10:0] add_515143;
  wire [11:0] sel_515145;
  wire [10:0] add_515147;
  wire [11:0] sel_515149;
  wire [11:0] add_515151;
  wire [11:0] sel_515153;
  wire [11:0] add_515155;
  wire [11:0] sel_515157;
  wire [11:0] add_515159;
  wire [11:0] sel_515161;
  wire [11:0] add_515163;
  wire [11:0] sel_515165;
  wire [9:0] add_515167;
  wire [11:0] sel_515170;
  wire [9:0] add_515172;
  wire [11:0] sel_515175;
  wire [11:0] add_515177;
  wire [11:0] sel_515179;
  wire [11:0] add_515181;
  wire [11:0] sel_515183;
  wire [7:0] add_515185;
  wire [11:0] sel_515188;
  wire [7:0] add_515190;
  wire [11:0] sel_515193;
  wire [11:0] add_515195;
  wire [11:0] sel_515197;
  wire [11:0] add_515199;
  wire [11:0] sel_515201;
  wire [10:0] add_515203;
  wire [11:0] sel_515205;
  wire [10:0] add_515207;
  wire [11:0] sel_515209;
  wire [10:0] add_515211;
  wire [11:0] sel_515213;
  wire [10:0] add_515215;
  wire [11:0] sel_515217;
  wire [10:0] add_515219;
  wire [11:0] sel_515222;
  wire [10:0] add_515224;
  wire [11:0] sel_515227;
  wire [11:0] add_515298;
  wire [11:0] sel_515300;
  wire [11:0] add_515303;
  wire [11:0] sel_515305;
  wire [8:0] add_515307;
  wire [8:0] add_515309;
  wire [15:0] array_index_515398;
  wire [15:0] array_index_515401;
  wire [11:0] add_515411;
  wire [11:0] sel_515413;
  wire [11:0] add_515415;
  wire [11:0] sel_515417;
  wire [8:0] add_515419;
  wire [11:0] sel_515422;
  wire [8:0] add_515424;
  wire [11:0] sel_515427;
  wire [10:0] add_515429;
  wire [11:0] sel_515431;
  wire [10:0] add_515433;
  wire [11:0] sel_515435;
  wire [9:0] add_515437;
  wire [11:0] sel_515439;
  wire [9:0] add_515441;
  wire [11:0] sel_515443;
  wire [11:0] add_515445;
  wire [11:0] sel_515447;
  wire [11:0] add_515449;
  wire [11:0] sel_515451;
  wire [10:0] add_515453;
  wire [11:0] sel_515455;
  wire [10:0] add_515457;
  wire [11:0] sel_515459;
  wire [11:0] add_515461;
  wire [11:0] sel_515463;
  wire [11:0] add_515465;
  wire [11:0] sel_515467;
  wire [11:0] add_515469;
  wire [11:0] sel_515471;
  wire [11:0] add_515473;
  wire [11:0] sel_515475;
  wire [9:0] add_515477;
  wire [11:0] sel_515480;
  wire [9:0] add_515482;
  wire [11:0] sel_515485;
  wire [11:0] add_515487;
  wire [11:0] sel_515489;
  wire [11:0] add_515491;
  wire [11:0] sel_515493;
  wire [7:0] add_515495;
  wire [11:0] sel_515498;
  wire [7:0] add_515500;
  wire [11:0] sel_515503;
  wire [11:0] add_515505;
  wire [11:0] sel_515507;
  wire [11:0] add_515509;
  wire [11:0] sel_515511;
  wire [10:0] add_515513;
  wire [11:0] sel_515515;
  wire [10:0] add_515517;
  wire [11:0] sel_515519;
  wire [10:0] add_515521;
  wire [11:0] sel_515523;
  wire [10:0] add_515525;
  wire [11:0] sel_515527;
  wire [10:0] add_515529;
  wire [11:0] sel_515532;
  wire [10:0] add_515534;
  wire [11:0] sel_515537;
  wire [11:0] add_515545;
  wire [11:0] add_515547;
  wire [11:0] add_515618;
  wire [11:0] sel_515620;
  wire [11:0] add_515623;
  wire [11:0] sel_515625;
  wire [8:0] add_515633;
  wire [11:0] sel_515635;
  wire [8:0] add_515637;
  wire [11:0] sel_515639;
  wire [15:0] array_index_515726;
  wire [15:0] array_index_515729;
  wire [10:0] add_515733;
  wire [10:0] add_515735;
  wire [11:0] add_515747;
  wire [11:0] sel_515749;
  wire [11:0] add_515751;
  wire [11:0] sel_515753;
  wire [8:0] add_515755;
  wire [11:0] sel_515758;
  wire [8:0] add_515760;
  wire [11:0] sel_515763;
  wire [10:0] add_515765;
  wire [11:0] sel_515767;
  wire [10:0] add_515769;
  wire [11:0] sel_515771;
  wire [9:0] add_515773;
  wire [11:0] sel_515775;
  wire [9:0] add_515777;
  wire [11:0] sel_515779;
  wire [11:0] add_515781;
  wire [11:0] sel_515783;
  wire [11:0] add_515785;
  wire [11:0] sel_515787;
  wire [10:0] add_515789;
  wire [11:0] sel_515791;
  wire [10:0] add_515793;
  wire [11:0] sel_515795;
  wire [11:0] add_515797;
  wire [11:0] sel_515799;
  wire [11:0] add_515801;
  wire [11:0] sel_515803;
  wire [11:0] add_515805;
  wire [11:0] sel_515807;
  wire [11:0] add_515809;
  wire [11:0] sel_515811;
  wire [9:0] add_515813;
  wire [11:0] sel_515816;
  wire [9:0] add_515818;
  wire [11:0] sel_515821;
  wire [11:0] add_515823;
  wire [11:0] sel_515825;
  wire [11:0] add_515827;
  wire [11:0] sel_515829;
  wire [7:0] add_515831;
  wire [11:0] sel_515834;
  wire [7:0] add_515836;
  wire [11:0] sel_515839;
  wire [11:0] add_515841;
  wire [11:0] sel_515843;
  wire [11:0] add_515845;
  wire [11:0] sel_515847;
  wire [10:0] add_515849;
  wire [11:0] sel_515851;
  wire [10:0] add_515853;
  wire [11:0] sel_515855;
  wire [10:0] add_515857;
  wire [11:0] sel_515859;
  wire [10:0] add_515861;
  wire [11:0] sel_515863;
  wire [10:0] add_515865;
  wire [11:0] sel_515868;
  wire [10:0] add_515870;
  wire [11:0] sel_515873;
  wire [11:0] add_515887;
  wire [11:0] sel_515889;
  wire [11:0] add_515891;
  wire [11:0] sel_515893;
  wire [11:0] add_515962;
  wire [11:0] sel_515964;
  wire [11:0] add_515967;
  wire [11:0] sel_515969;
  wire [11:0] add_515971;
  wire [11:0] add_515973;
  wire [8:0] add_515987;
  wire [11:0] sel_515989;
  wire [8:0] add_515991;
  wire [11:0] sel_515993;
  wire [15:0] array_index_516080;
  wire [15:0] array_index_516083;
  wire [10:0] add_516093;
  wire [11:0] sel_516095;
  wire [10:0] add_516097;
  wire [11:0] sel_516099;
  wire [11:0] add_516109;
  wire [11:0] sel_516111;
  wire [11:0] add_516113;
  wire [11:0] sel_516115;
  wire [8:0] add_516117;
  wire [11:0] sel_516120;
  wire [8:0] add_516122;
  wire [11:0] sel_516125;
  wire [10:0] add_516127;
  wire [11:0] sel_516129;
  wire [10:0] add_516131;
  wire [11:0] sel_516133;
  wire [9:0] add_516135;
  wire [11:0] sel_516137;
  wire [9:0] add_516139;
  wire [11:0] sel_516141;
  wire [11:0] add_516143;
  wire [11:0] sel_516145;
  wire [11:0] add_516147;
  wire [11:0] sel_516149;
  wire [10:0] add_516151;
  wire [11:0] sel_516153;
  wire [10:0] add_516155;
  wire [11:0] sel_516157;
  wire [11:0] add_516159;
  wire [11:0] sel_516161;
  wire [11:0] add_516163;
  wire [11:0] sel_516165;
  wire [11:0] add_516167;
  wire [11:0] sel_516169;
  wire [11:0] add_516171;
  wire [11:0] sel_516173;
  wire [9:0] add_516175;
  wire [11:0] sel_516178;
  wire [9:0] add_516180;
  wire [11:0] sel_516183;
  wire [11:0] add_516185;
  wire [11:0] sel_516187;
  wire [11:0] add_516189;
  wire [11:0] sel_516191;
  wire [7:0] add_516193;
  wire [11:0] sel_516196;
  wire [7:0] add_516198;
  wire [11:0] sel_516201;
  wire [11:0] add_516203;
  wire [11:0] sel_516205;
  wire [11:0] add_516207;
  wire [11:0] sel_516209;
  wire [10:0] add_516211;
  wire [11:0] sel_516213;
  wire [10:0] add_516215;
  wire [11:0] sel_516217;
  wire [10:0] add_516219;
  wire [11:0] sel_516221;
  wire [10:0] add_516223;
  wire [11:0] sel_516225;
  wire [10:0] add_516227;
  wire [11:0] sel_516230;
  wire [10:0] add_516232;
  wire [11:0] sel_516235;
  wire [11:0] add_516243;
  wire [11:0] add_516245;
  wire [11:0] add_516257;
  wire [11:0] sel_516259;
  wire [11:0] add_516261;
  wire [11:0] sel_516263;
  wire [11:0] add_516332;
  wire [11:0] sel_516334;
  wire [11:0] add_516337;
  wire [11:0] sel_516339;
  wire [11:0] add_516347;
  wire [11:0] sel_516349;
  wire [11:0] add_516351;
  wire [11:0] sel_516353;
  wire [8:0] add_516365;
  wire [11:0] sel_516367;
  wire [8:0] add_516369;
  wire [11:0] sel_516371;
  wire [15:0] array_index_516458;
  wire [15:0] array_index_516461;
  wire [11:0] add_516465;
  wire [11:0] add_516467;
  wire [10:0] add_516479;
  wire [11:0] sel_516481;
  wire [10:0] add_516483;
  wire [11:0] sel_516485;
  wire [11:0] add_516495;
  wire [11:0] sel_516497;
  wire [11:0] add_516499;
  wire [11:0] sel_516501;
  wire [8:0] add_516503;
  wire [11:0] sel_516506;
  wire [8:0] add_516508;
  wire [11:0] sel_516511;
  wire [10:0] add_516513;
  wire [11:0] sel_516515;
  wire [10:0] add_516517;
  wire [11:0] sel_516519;
  wire [9:0] add_516521;
  wire [11:0] sel_516523;
  wire [9:0] add_516525;
  wire [11:0] sel_516527;
  wire [11:0] add_516529;
  wire [11:0] sel_516531;
  wire [11:0] add_516533;
  wire [11:0] sel_516535;
  wire [10:0] add_516537;
  wire [11:0] sel_516539;
  wire [10:0] add_516541;
  wire [11:0] sel_516543;
  wire [11:0] add_516545;
  wire [11:0] sel_516547;
  wire [11:0] add_516549;
  wire [11:0] sel_516551;
  wire [11:0] add_516553;
  wire [11:0] sel_516555;
  wire [11:0] add_516557;
  wire [11:0] sel_516559;
  wire [9:0] add_516561;
  wire [11:0] sel_516564;
  wire [9:0] add_516566;
  wire [11:0] sel_516569;
  wire [11:0] add_516571;
  wire [11:0] sel_516573;
  wire [11:0] add_516575;
  wire [11:0] sel_516577;
  wire [7:0] add_516579;
  wire [11:0] sel_516582;
  wire [7:0] add_516584;
  wire [11:0] sel_516587;
  wire [11:0] add_516589;
  wire [11:0] sel_516591;
  wire [11:0] add_516593;
  wire [11:0] sel_516595;
  wire [10:0] add_516597;
  wire [11:0] sel_516599;
  wire [10:0] add_516601;
  wire [11:0] sel_516603;
  wire [10:0] add_516605;
  wire [11:0] sel_516607;
  wire [10:0] add_516609;
  wire [11:0] sel_516611;
  wire [10:0] add_516613;
  wire [11:0] sel_516616;
  wire [10:0] add_516618;
  wire [11:0] sel_516621;
  wire [11:0] add_516635;
  wire [11:0] sel_516637;
  wire [11:0] add_516639;
  wire [11:0] sel_516641;
  wire [11:0] add_516651;
  wire [11:0] sel_516653;
  wire [11:0] add_516655;
  wire [11:0] sel_516657;
  wire [11:0] add_516726;
  wire [11:0] sel_516728;
  wire [11:0] add_516731;
  wire [11:0] sel_516733;
  wire [11:0] add_516735;
  wire [11:0] add_516737;
  wire [11:0] add_516749;
  wire [11:0] sel_516751;
  wire [11:0] add_516753;
  wire [11:0] sel_516755;
  wire [8:0] add_516767;
  wire [11:0] sel_516769;
  wire [8:0] add_516771;
  wire [11:0] sel_516773;
  wire [15:0] array_index_516860;
  wire [15:0] array_index_516863;
  wire [11:0] add_516873;
  wire [11:0] sel_516875;
  wire [11:0] add_516877;
  wire [11:0] sel_516879;
  wire [10:0] add_516889;
  wire [11:0] sel_516891;
  wire [10:0] add_516893;
  wire [11:0] sel_516895;
  wire [11:0] add_516905;
  wire [11:0] sel_516907;
  wire [11:0] add_516909;
  wire [11:0] sel_516911;
  wire [8:0] add_516913;
  wire [11:0] sel_516916;
  wire [8:0] add_516918;
  wire [11:0] sel_516921;
  wire [10:0] add_516923;
  wire [11:0] sel_516925;
  wire [10:0] add_516927;
  wire [11:0] sel_516929;
  wire [9:0] add_516931;
  wire [11:0] sel_516933;
  wire [9:0] add_516935;
  wire [11:0] sel_516937;
  wire [11:0] add_516939;
  wire [11:0] sel_516941;
  wire [11:0] add_516943;
  wire [11:0] sel_516945;
  wire [10:0] add_516947;
  wire [11:0] sel_516949;
  wire [10:0] add_516951;
  wire [11:0] sel_516953;
  wire [11:0] add_516955;
  wire [11:0] sel_516957;
  wire [11:0] add_516959;
  wire [11:0] sel_516961;
  wire [11:0] add_516963;
  wire [11:0] sel_516965;
  wire [11:0] add_516967;
  wire [11:0] sel_516969;
  wire [9:0] add_516971;
  wire [11:0] sel_516974;
  wire [9:0] add_516976;
  wire [11:0] sel_516979;
  wire [11:0] add_516981;
  wire [11:0] sel_516983;
  wire [11:0] add_516985;
  wire [11:0] sel_516987;
  wire [7:0] add_516989;
  wire [11:0] sel_516992;
  wire [7:0] add_516994;
  wire [11:0] sel_516997;
  wire [11:0] add_516999;
  wire [11:0] sel_517001;
  wire [11:0] add_517003;
  wire [11:0] sel_517005;
  wire [10:0] add_517007;
  wire [11:0] sel_517009;
  wire [10:0] add_517011;
  wire [11:0] sel_517013;
  wire [10:0] add_517015;
  wire [11:0] sel_517017;
  wire [10:0] add_517019;
  wire [11:0] sel_517021;
  wire [10:0] add_517023;
  wire [11:0] sel_517026;
  wire [10:0] add_517028;
  wire [11:0] sel_517031;
  wire [11:0] add_517039;
  wire [11:0] add_517041;
  wire [11:0] add_517053;
  wire [11:0] sel_517055;
  wire [11:0] add_517057;
  wire [11:0] sel_517059;
  wire [11:0] add_517069;
  wire [11:0] sel_517071;
  wire [11:0] add_517073;
  wire [11:0] sel_517075;
  wire [11:0] add_517144;
  wire [11:0] sel_517146;
  wire [11:0] add_517149;
  wire [11:0] sel_517151;
  wire [11:0] add_517159;
  wire [11:0] sel_517161;
  wire [11:0] add_517163;
  wire [11:0] sel_517165;
  wire [11:0] add_517175;
  wire [11:0] sel_517177;
  wire [11:0] add_517179;
  wire [11:0] sel_517181;
  wire [8:0] add_517193;
  wire [11:0] sel_517195;
  wire [8:0] add_517197;
  wire [11:0] sel_517199;
  wire [15:0] array_index_517286;
  wire [15:0] array_index_517289;
  wire [11:0] add_517293;
  wire [11:0] add_517295;
  wire [11:0] add_517307;
  wire [11:0] sel_517309;
  wire [11:0] add_517311;
  wire [11:0] sel_517313;
  wire [10:0] add_517323;
  wire [11:0] sel_517325;
  wire [10:0] add_517327;
  wire [11:0] sel_517329;
  wire [11:0] add_517339;
  wire [11:0] sel_517341;
  wire [11:0] add_517343;
  wire [11:0] sel_517345;
  wire [8:0] add_517347;
  wire [11:0] sel_517350;
  wire [8:0] add_517352;
  wire [11:0] sel_517355;
  wire [10:0] add_517357;
  wire [11:0] sel_517359;
  wire [10:0] add_517361;
  wire [11:0] sel_517363;
  wire [9:0] add_517365;
  wire [11:0] sel_517367;
  wire [9:0] add_517369;
  wire [11:0] sel_517371;
  wire [11:0] add_517373;
  wire [11:0] sel_517375;
  wire [11:0] add_517377;
  wire [11:0] sel_517379;
  wire [10:0] add_517381;
  wire [11:0] sel_517383;
  wire [10:0] add_517385;
  wire [11:0] sel_517387;
  wire [11:0] add_517389;
  wire [11:0] sel_517391;
  wire [11:0] add_517393;
  wire [11:0] sel_517395;
  wire [11:0] add_517397;
  wire [11:0] sel_517399;
  wire [11:0] add_517401;
  wire [11:0] sel_517403;
  wire [9:0] add_517405;
  wire [11:0] sel_517408;
  wire [9:0] add_517410;
  wire [11:0] sel_517413;
  wire [11:0] add_517415;
  wire [11:0] sel_517417;
  wire [11:0] add_517419;
  wire [11:0] sel_517421;
  wire [7:0] add_517423;
  wire [11:0] sel_517426;
  wire [7:0] add_517428;
  wire [11:0] sel_517431;
  wire [11:0] add_517433;
  wire [11:0] sel_517435;
  wire [11:0] add_517437;
  wire [11:0] sel_517439;
  wire [10:0] add_517441;
  wire [11:0] sel_517443;
  wire [10:0] add_517445;
  wire [11:0] sel_517447;
  wire [10:0] add_517449;
  wire [11:0] sel_517451;
  wire [10:0] add_517453;
  wire [11:0] sel_517455;
  wire [10:0] add_517457;
  wire [11:0] sel_517460;
  wire [10:0] add_517462;
  wire [11:0] sel_517465;
  wire [11:0] add_517479;
  wire [11:0] sel_517481;
  wire [11:0] add_517483;
  wire [11:0] sel_517485;
  wire [11:0] add_517495;
  wire [11:0] sel_517497;
  wire [11:0] add_517499;
  wire [11:0] sel_517501;
  wire [11:0] add_517511;
  wire [11:0] sel_517513;
  wire [11:0] add_517515;
  wire [11:0] sel_517517;
  wire [11:0] add_517586;
  wire [11:0] sel_517588;
  wire [11:0] add_517591;
  wire [11:0] sel_517593;
  wire [11:0] add_517595;
  wire [11:0] add_517597;
  wire [11:0] add_517609;
  wire [11:0] sel_517611;
  wire [11:0] add_517613;
  wire [11:0] sel_517615;
  wire [11:0] add_517625;
  wire [11:0] sel_517627;
  wire [11:0] add_517629;
  wire [11:0] sel_517631;
  wire [8:0] add_517643;
  wire [11:0] sel_517645;
  wire [8:0] add_517647;
  wire [11:0] sel_517649;
  wire [15:0] array_index_517736;
  wire [15:0] array_index_517739;
  wire [11:0] add_517749;
  wire [11:0] sel_517751;
  wire [11:0] add_517753;
  wire [11:0] sel_517755;
  wire [11:0] add_517765;
  wire [11:0] sel_517767;
  wire [11:0] add_517769;
  wire [11:0] sel_517771;
  wire [10:0] add_517781;
  wire [11:0] sel_517783;
  wire [10:0] add_517785;
  wire [11:0] sel_517787;
  wire [11:0] add_517797;
  wire [11:0] sel_517799;
  wire [11:0] add_517801;
  wire [11:0] sel_517803;
  wire [8:0] add_517805;
  wire [11:0] sel_517808;
  wire [8:0] add_517810;
  wire [11:0] sel_517813;
  wire [10:0] add_517815;
  wire [11:0] sel_517817;
  wire [10:0] add_517819;
  wire [11:0] sel_517821;
  wire [9:0] add_517823;
  wire [11:0] sel_517825;
  wire [9:0] add_517827;
  wire [11:0] sel_517829;
  wire [11:0] add_517831;
  wire [11:0] sel_517833;
  wire [11:0] add_517835;
  wire [11:0] sel_517837;
  wire [10:0] add_517839;
  wire [11:0] sel_517841;
  wire [10:0] add_517843;
  wire [11:0] sel_517845;
  wire [11:0] add_517847;
  wire [11:0] sel_517849;
  wire [11:0] add_517851;
  wire [11:0] sel_517853;
  wire [11:0] add_517855;
  wire [11:0] sel_517857;
  wire [11:0] add_517859;
  wire [11:0] sel_517861;
  wire [9:0] add_517863;
  wire [11:0] sel_517866;
  wire [9:0] add_517868;
  wire [11:0] sel_517871;
  wire [11:0] add_517873;
  wire [11:0] sel_517875;
  wire [11:0] add_517877;
  wire [11:0] sel_517879;
  wire [7:0] add_517881;
  wire [11:0] sel_517884;
  wire [7:0] add_517886;
  wire [11:0] sel_517889;
  wire [11:0] add_517891;
  wire [11:0] sel_517893;
  wire [11:0] add_517895;
  wire [11:0] sel_517897;
  wire [10:0] add_517899;
  wire [11:0] sel_517901;
  wire [10:0] add_517903;
  wire [11:0] sel_517905;
  wire [10:0] add_517907;
  wire [11:0] sel_517909;
  wire [10:0] add_517911;
  wire [11:0] sel_517913;
  wire [10:0] add_517915;
  wire [11:0] sel_517918;
  wire [10:0] add_517920;
  wire [11:0] sel_517923;
  wire [10:0] add_517931;
  wire [10:0] add_517933;
  wire [11:0] add_517945;
  wire [11:0] sel_517947;
  wire [11:0] add_517949;
  wire [11:0] sel_517951;
  wire [11:0] add_517961;
  wire [11:0] sel_517963;
  wire [11:0] add_517965;
  wire [11:0] sel_517967;
  wire [11:0] add_517977;
  wire [11:0] sel_517979;
  wire [11:0] add_517981;
  wire [11:0] sel_517983;
  wire [11:0] add_518052;
  wire [11:0] sel_518054;
  wire [11:0] add_518057;
  wire [11:0] sel_518059;
  wire [11:0] add_518067;
  wire [11:0] sel_518069;
  wire [11:0] add_518071;
  wire [11:0] sel_518073;
  wire [11:0] add_518083;
  wire [11:0] sel_518085;
  wire [11:0] add_518087;
  wire [11:0] sel_518089;
  wire [11:0] add_518099;
  wire [11:0] sel_518101;
  wire [11:0] add_518103;
  wire [11:0] sel_518105;
  wire [8:0] add_518117;
  wire [11:0] sel_518119;
  wire [8:0] add_518121;
  wire [11:0] sel_518123;
  wire [15:0] array_index_518210;
  wire [15:0] array_index_518213;
  wire [11:0] add_518217;
  wire [11:0] add_518219;
  wire [11:0] add_518233;
  wire [11:0] sel_518235;
  wire [11:0] add_518237;
  wire [11:0] sel_518239;
  wire [11:0] add_518249;
  wire [11:0] sel_518251;
  wire [11:0] add_518253;
  wire [11:0] sel_518255;
  wire [10:0] add_518265;
  wire [11:0] sel_518267;
  wire [10:0] add_518269;
  wire [11:0] sel_518271;
  wire [11:0] add_518281;
  wire [11:0] sel_518283;
  wire [11:0] add_518285;
  wire [11:0] sel_518287;
  wire [8:0] add_518289;
  wire [11:0] sel_518292;
  wire [8:0] add_518294;
  wire [11:0] sel_518297;
  wire [10:0] add_518299;
  wire [11:0] sel_518301;
  wire [10:0] add_518303;
  wire [11:0] sel_518305;
  wire [9:0] add_518307;
  wire [11:0] sel_518309;
  wire [9:0] add_518311;
  wire [11:0] sel_518313;
  wire [11:0] add_518315;
  wire [11:0] sel_518317;
  wire [11:0] add_518319;
  wire [11:0] sel_518321;
  wire [10:0] add_518323;
  wire [11:0] sel_518325;
  wire [10:0] add_518327;
  wire [11:0] sel_518329;
  wire [11:0] add_518331;
  wire [11:0] sel_518333;
  wire [11:0] add_518335;
  wire [11:0] sel_518337;
  wire [11:0] add_518339;
  wire [11:0] sel_518341;
  wire [11:0] add_518343;
  wire [11:0] sel_518345;
  wire [9:0] add_518347;
  wire [11:0] sel_518350;
  wire [9:0] add_518352;
  wire [11:0] sel_518355;
  wire [11:0] add_518357;
  wire [11:0] sel_518359;
  wire [11:0] add_518361;
  wire [11:0] sel_518363;
  wire [7:0] add_518365;
  wire [11:0] sel_518368;
  wire [7:0] add_518370;
  wire [11:0] sel_518373;
  wire [11:0] add_518375;
  wire [11:0] sel_518377;
  wire [11:0] add_518379;
  wire [11:0] sel_518381;
  wire [10:0] add_518383;
  wire [11:0] sel_518385;
  wire [10:0] add_518387;
  wire [11:0] sel_518389;
  wire [10:0] add_518391;
  wire [11:0] sel_518393;
  wire [10:0] add_518395;
  wire [11:0] sel_518397;
  wire [10:0] add_518399;
  wire [11:0] sel_518402;
  wire [10:0] add_518404;
  wire [11:0] sel_518407;
  wire [10:0] add_518421;
  wire [11:0] sel_518423;
  wire [10:0] add_518425;
  wire [11:0] sel_518427;
  wire [11:0] add_518437;
  wire [11:0] sel_518439;
  wire [11:0] add_518441;
  wire [11:0] sel_518443;
  wire [11:0] add_518453;
  wire [11:0] sel_518455;
  wire [11:0] add_518457;
  wire [11:0] sel_518459;
  wire [11:0] add_518469;
  wire [11:0] sel_518471;
  wire [11:0] add_518473;
  wire [11:0] sel_518475;
  wire [11:0] add_518544;
  wire [11:0] sel_518546;
  wire [11:0] add_518549;
  wire [11:0] sel_518551;
  wire [10:0] add_518553;
  wire [10:0] add_518555;
  wire [11:0] add_518567;
  wire [11:0] sel_518569;
  wire [11:0] add_518571;
  wire [11:0] sel_518573;
  wire [11:0] add_518583;
  wire [11:0] sel_518585;
  wire [11:0] add_518587;
  wire [11:0] sel_518589;
  wire [11:0] add_518599;
  wire [11:0] sel_518601;
  wire [11:0] add_518603;
  wire [11:0] sel_518605;
  wire [8:0] add_518617;
  wire [11:0] sel_518619;
  wire [8:0] add_518621;
  wire [11:0] sel_518623;
  wire [15:0] array_index_518710;
  wire [15:0] array_index_518713;
  wire [11:0] add_518723;
  wire [11:0] sel_518725;
  wire [11:0] add_518727;
  wire [11:0] sel_518729;
  wire [11:0] add_518741;
  wire [11:0] sel_518743;
  wire [11:0] add_518745;
  wire [11:0] sel_518747;
  wire [11:0] add_518757;
  wire [11:0] sel_518759;
  wire [11:0] add_518761;
  wire [11:0] sel_518763;
  wire [10:0] add_518773;
  wire [11:0] sel_518775;
  wire [10:0] add_518777;
  wire [11:0] sel_518779;
  wire [11:0] add_518789;
  wire [11:0] sel_518791;
  wire [11:0] add_518793;
  wire [11:0] sel_518795;
  wire [8:0] add_518797;
  wire [11:0] sel_518800;
  wire [8:0] add_518802;
  wire [11:0] sel_518805;
  wire [10:0] add_518807;
  wire [11:0] sel_518809;
  wire [10:0] add_518811;
  wire [11:0] sel_518813;
  wire [9:0] add_518815;
  wire [11:0] sel_518817;
  wire [9:0] add_518819;
  wire [11:0] sel_518821;
  wire [11:0] add_518823;
  wire [11:0] sel_518825;
  wire [11:0] add_518827;
  wire [11:0] sel_518829;
  wire [10:0] add_518831;
  wire [11:0] sel_518833;
  wire [10:0] add_518835;
  wire [11:0] sel_518837;
  wire [11:0] add_518839;
  wire [11:0] sel_518841;
  wire [11:0] add_518843;
  wire [11:0] sel_518845;
  wire [11:0] add_518847;
  wire [11:0] sel_518849;
  wire [11:0] add_518851;
  wire [11:0] sel_518853;
  wire [9:0] add_518855;
  wire [11:0] sel_518858;
  wire [9:0] add_518860;
  wire [11:0] sel_518863;
  wire [11:0] add_518865;
  wire [11:0] sel_518867;
  wire [11:0] add_518869;
  wire [11:0] sel_518871;
  wire [7:0] add_518873;
  wire [11:0] sel_518876;
  wire [7:0] add_518878;
  wire [11:0] sel_518881;
  wire [11:0] add_518883;
  wire [11:0] sel_518885;
  wire [11:0] add_518887;
  wire [11:0] sel_518889;
  wire [10:0] add_518891;
  wire [11:0] sel_518893;
  wire [10:0] add_518895;
  wire [11:0] sel_518897;
  wire [10:0] add_518899;
  wire [11:0] sel_518901;
  wire [10:0] add_518903;
  wire [11:0] sel_518905;
  wire [10:0] add_518907;
  wire [11:0] sel_518910;
  wire [10:0] add_518912;
  wire [11:0] sel_518915;
  wire [11:0] add_518923;
  wire [11:0] add_518925;
  wire [10:0] add_518939;
  wire [11:0] sel_518941;
  wire [10:0] add_518943;
  wire [11:0] sel_518945;
  wire [11:0] add_518955;
  wire [11:0] sel_518957;
  wire [11:0] add_518959;
  wire [11:0] sel_518961;
  wire [11:0] add_518971;
  wire [11:0] sel_518973;
  wire [11:0] add_518975;
  wire [11:0] sel_518977;
  wire [11:0] add_518987;
  wire [11:0] sel_518989;
  wire [11:0] add_518991;
  wire [11:0] sel_518993;
  wire [11:0] add_519062;
  wire [11:0] sel_519064;
  wire [11:0] add_519067;
  wire [11:0] sel_519069;
  wire [10:0] add_519077;
  wire [11:0] sel_519079;
  wire [10:0] add_519081;
  wire [11:0] sel_519083;
  wire [11:0] add_519093;
  wire [11:0] sel_519095;
  wire [11:0] add_519097;
  wire [11:0] sel_519099;
  wire [11:0] add_519109;
  wire [11:0] sel_519111;
  wire [11:0] add_519113;
  wire [11:0] sel_519115;
  wire [11:0] add_519125;
  wire [11:0] sel_519127;
  wire [11:0] add_519129;
  wire [11:0] sel_519131;
  wire [8:0] add_519143;
  wire [11:0] sel_519145;
  wire [8:0] add_519147;
  wire [11:0] sel_519149;
  wire [15:0] array_index_519236;
  wire [15:0] array_index_519239;
  wire [11:0] add_519243;
  wire [11:0] add_519245;
  wire [11:0] add_519257;
  wire [11:0] sel_519259;
  wire [11:0] add_519261;
  wire [11:0] sel_519263;
  wire [11:0] add_519275;
  wire [11:0] sel_519277;
  wire [11:0] add_519279;
  wire [11:0] sel_519281;
  wire [11:0] add_519291;
  wire [11:0] sel_519293;
  wire [11:0] add_519295;
  wire [11:0] sel_519297;
  wire [10:0] add_519307;
  wire [11:0] sel_519309;
  wire [10:0] add_519311;
  wire [11:0] sel_519313;
  wire [11:0] add_519323;
  wire [11:0] sel_519325;
  wire [11:0] add_519327;
  wire [11:0] sel_519329;
  wire [8:0] add_519331;
  wire [11:0] sel_519334;
  wire [8:0] add_519336;
  wire [11:0] sel_519339;
  wire [10:0] add_519341;
  wire [11:0] sel_519343;
  wire [10:0] add_519345;
  wire [11:0] sel_519347;
  wire [9:0] add_519349;
  wire [11:0] sel_519351;
  wire [9:0] add_519353;
  wire [11:0] sel_519355;
  wire [11:0] add_519357;
  wire [11:0] sel_519359;
  wire [11:0] add_519361;
  wire [11:0] sel_519363;
  wire [10:0] add_519365;
  wire [11:0] sel_519367;
  wire [10:0] add_519369;
  wire [11:0] sel_519371;
  wire [11:0] add_519373;
  wire [11:0] sel_519375;
  wire [11:0] add_519377;
  wire [11:0] sel_519379;
  wire [11:0] add_519381;
  wire [11:0] sel_519383;
  wire [11:0] add_519385;
  wire [11:0] sel_519387;
  wire [9:0] add_519389;
  wire [11:0] sel_519392;
  wire [9:0] add_519394;
  wire [11:0] sel_519397;
  wire [11:0] add_519399;
  wire [11:0] sel_519401;
  wire [11:0] add_519403;
  wire [11:0] sel_519405;
  wire [7:0] add_519407;
  wire [11:0] sel_519410;
  wire [7:0] add_519412;
  wire [11:0] sel_519415;
  wire [11:0] add_519417;
  wire [11:0] sel_519419;
  wire [11:0] add_519421;
  wire [11:0] sel_519423;
  wire [10:0] add_519425;
  wire [11:0] sel_519427;
  wire [10:0] add_519429;
  wire [11:0] sel_519431;
  wire [10:0] add_519433;
  wire [11:0] sel_519435;
  wire [10:0] add_519437;
  wire [11:0] sel_519439;
  wire [10:0] add_519441;
  wire [11:0] sel_519444;
  wire [10:0] add_519446;
  wire [11:0] sel_519449;
  wire [11:0] add_519463;
  wire [11:0] sel_519465;
  wire [11:0] add_519467;
  wire [11:0] sel_519469;
  wire [10:0] add_519481;
  wire [11:0] sel_519483;
  wire [10:0] add_519485;
  wire [11:0] sel_519487;
  wire [11:0] add_519497;
  wire [11:0] sel_519499;
  wire [11:0] add_519501;
  wire [11:0] sel_519503;
  wire [11:0] add_519513;
  wire [11:0] sel_519515;
  wire [11:0] add_519517;
  wire [11:0] sel_519519;
  wire [11:0] add_519529;
  wire [11:0] sel_519531;
  wire [11:0] add_519533;
  wire [11:0] sel_519535;
  wire [11:0] add_519604;
  wire [11:0] sel_519606;
  wire [11:0] add_519609;
  wire [11:0] sel_519611;
  wire [10:0] add_519613;
  wire [10:0] add_519615;
  wire [10:0] add_519627;
  wire [11:0] sel_519629;
  wire [10:0] add_519631;
  wire [11:0] sel_519633;
  wire [11:0] add_519643;
  wire [11:0] sel_519645;
  wire [11:0] add_519647;
  wire [11:0] sel_519649;
  wire [11:0] add_519659;
  wire [11:0] sel_519661;
  wire [11:0] add_519663;
  wire [11:0] sel_519665;
  wire [11:0] add_519675;
  wire [11:0] sel_519677;
  wire [11:0] add_519679;
  wire [11:0] sel_519681;
  wire [8:0] add_519693;
  wire [11:0] sel_519695;
  wire [8:0] add_519697;
  wire [11:0] sel_519699;
  wire [15:0] array_index_519786;
  wire [15:0] array_index_519789;
  wire [11:0] add_519799;
  wire [11:0] sel_519801;
  wire [11:0] add_519803;
  wire [11:0] sel_519805;
  wire [11:0] add_519815;
  wire [11:0] sel_519817;
  wire [11:0] add_519819;
  wire [11:0] sel_519821;
  wire [11:0] add_519833;
  wire [11:0] sel_519835;
  wire [11:0] add_519837;
  wire [11:0] sel_519839;
  wire [11:0] add_519849;
  wire [11:0] sel_519851;
  wire [11:0] add_519853;
  wire [11:0] sel_519855;
  wire [10:0] add_519865;
  wire [11:0] sel_519867;
  wire [10:0] add_519869;
  wire [11:0] sel_519871;
  wire [11:0] add_519881;
  wire [11:0] sel_519883;
  wire [11:0] add_519885;
  wire [11:0] sel_519887;
  wire [8:0] add_519889;
  wire [11:0] sel_519892;
  wire [8:0] add_519894;
  wire [11:0] sel_519897;
  wire [10:0] add_519899;
  wire [11:0] sel_519901;
  wire [10:0] add_519903;
  wire [11:0] sel_519905;
  wire [9:0] add_519907;
  wire [11:0] sel_519909;
  wire [9:0] add_519911;
  wire [11:0] sel_519913;
  wire [11:0] add_519915;
  wire [11:0] sel_519917;
  wire [11:0] add_519919;
  wire [11:0] sel_519921;
  wire [10:0] add_519923;
  wire [11:0] sel_519925;
  wire [10:0] add_519927;
  wire [11:0] sel_519929;
  wire [11:0] add_519931;
  wire [11:0] sel_519933;
  wire [11:0] add_519935;
  wire [11:0] sel_519937;
  wire [11:0] add_519939;
  wire [11:0] sel_519941;
  wire [11:0] add_519943;
  wire [11:0] sel_519945;
  wire [9:0] add_519947;
  wire [11:0] sel_519950;
  wire [9:0] add_519952;
  wire [11:0] sel_519955;
  wire [11:0] add_519957;
  wire [11:0] sel_519959;
  wire [11:0] add_519961;
  wire [11:0] sel_519963;
  wire [7:0] add_519965;
  wire [11:0] sel_519968;
  wire [7:0] add_519970;
  wire [11:0] sel_519973;
  wire [11:0] add_519975;
  wire [11:0] sel_519977;
  wire [11:0] add_519979;
  wire [11:0] sel_519981;
  wire [10:0] add_519983;
  wire [11:0] sel_519985;
  wire [10:0] add_519987;
  wire [11:0] sel_519989;
  wire [10:0] add_519991;
  wire [11:0] sel_519993;
  wire [10:0] add_519995;
  wire [11:0] sel_519997;
  wire [10:0] add_519999;
  wire [11:0] sel_520002;
  wire [10:0] add_520004;
  wire [11:0] sel_520007;
  wire [11:0] add_520015;
  wire [11:0] add_520017;
  wire [11:0] add_520031;
  wire [11:0] sel_520033;
  wire [11:0] add_520035;
  wire [11:0] sel_520037;
  wire [10:0] add_520049;
  wire [11:0] sel_520051;
  wire [10:0] add_520053;
  wire [11:0] sel_520055;
  wire [11:0] add_520065;
  wire [11:0] sel_520067;
  wire [11:0] add_520069;
  wire [11:0] sel_520071;
  wire [11:0] add_520081;
  wire [11:0] sel_520083;
  wire [11:0] add_520085;
  wire [11:0] sel_520087;
  wire [11:0] add_520097;
  wire [11:0] sel_520099;
  wire [11:0] add_520101;
  wire [11:0] sel_520103;
  wire [11:0] add_520172;
  wire [11:0] sel_520174;
  wire [11:0] add_520177;
  wire [11:0] sel_520179;
  wire [10:0] add_520187;
  wire [11:0] sel_520189;
  wire [10:0] add_520191;
  wire [11:0] sel_520193;
  wire [10:0] add_520203;
  wire [11:0] sel_520205;
  wire [10:0] add_520207;
  wire [11:0] sel_520209;
  wire [11:0] add_520219;
  wire [11:0] sel_520221;
  wire [11:0] add_520223;
  wire [11:0] sel_520225;
  wire [11:0] add_520235;
  wire [11:0] sel_520237;
  wire [11:0] add_520239;
  wire [11:0] sel_520241;
  wire [11:0] add_520251;
  wire [11:0] sel_520253;
  wire [11:0] add_520255;
  wire [11:0] sel_520257;
  wire [8:0] add_520269;
  wire [11:0] sel_520271;
  wire [8:0] add_520273;
  wire [11:0] sel_520275;
  wire [15:0] array_index_520362;
  wire [15:0] array_index_520365;
  wire [8:0] add_520369;
  wire [8:0] add_520371;
  wire [11:0] add_520383;
  wire [11:0] sel_520385;
  wire [11:0] add_520387;
  wire [11:0] sel_520389;
  wire [11:0] add_520399;
  wire [11:0] sel_520401;
  wire [11:0] add_520403;
  wire [11:0] sel_520405;
  wire [11:0] add_520417;
  wire [11:0] sel_520419;
  wire [11:0] add_520421;
  wire [11:0] sel_520423;
  wire [11:0] add_520433;
  wire [11:0] sel_520435;
  wire [11:0] add_520437;
  wire [11:0] sel_520439;
  wire [10:0] add_520449;
  wire [11:0] sel_520451;
  wire [10:0] add_520453;
  wire [11:0] sel_520455;
  wire [11:0] add_520465;
  wire [11:0] sel_520467;
  wire [11:0] add_520469;
  wire [11:0] sel_520471;
  wire [8:0] add_520473;
  wire [11:0] sel_520476;
  wire [8:0] add_520478;
  wire [11:0] sel_520481;
  wire [10:0] add_520483;
  wire [11:0] sel_520485;
  wire [10:0] add_520487;
  wire [11:0] sel_520489;
  wire [9:0] add_520491;
  wire [11:0] sel_520493;
  wire [9:0] add_520495;
  wire [11:0] sel_520497;
  wire [11:0] add_520499;
  wire [11:0] sel_520501;
  wire [11:0] add_520503;
  wire [11:0] sel_520505;
  wire [10:0] add_520507;
  wire [11:0] sel_520509;
  wire [10:0] add_520511;
  wire [11:0] sel_520513;
  wire [11:0] add_520515;
  wire [11:0] sel_520517;
  wire [11:0] add_520519;
  wire [11:0] sel_520521;
  wire [11:0] add_520523;
  wire [11:0] sel_520525;
  wire [11:0] add_520527;
  wire [11:0] sel_520529;
  wire [9:0] add_520531;
  wire [11:0] sel_520534;
  wire [9:0] add_520536;
  wire [11:0] sel_520539;
  wire [11:0] add_520541;
  wire [11:0] sel_520543;
  wire [11:0] add_520545;
  wire [11:0] sel_520547;
  wire [7:0] add_520549;
  wire [11:0] sel_520552;
  wire [7:0] add_520554;
  wire [11:0] sel_520557;
  wire [11:0] add_520559;
  wire [11:0] sel_520561;
  wire [11:0] add_520563;
  wire [11:0] sel_520565;
  wire [10:0] add_520567;
  wire [11:0] sel_520569;
  wire [10:0] add_520571;
  wire [11:0] sel_520573;
  wire [10:0] add_520575;
  wire [11:0] sel_520577;
  wire [10:0] add_520579;
  wire [11:0] sel_520581;
  wire [10:0] add_520583;
  wire [11:0] sel_520586;
  wire [10:0] add_520588;
  wire [11:0] sel_520591;
  wire [11:0] add_520605;
  wire [11:0] sel_520607;
  wire [11:0] add_520609;
  wire [11:0] sel_520611;
  wire [11:0] add_520623;
  wire [11:0] sel_520625;
  wire [11:0] add_520627;
  wire [11:0] sel_520629;
  wire [10:0] add_520641;
  wire [11:0] sel_520643;
  wire [10:0] add_520645;
  wire [11:0] sel_520647;
  wire [11:0] add_520657;
  wire [11:0] sel_520659;
  wire [11:0] add_520661;
  wire [11:0] sel_520663;
  wire [11:0] add_520673;
  wire [11:0] sel_520675;
  wire [11:0] add_520677;
  wire [11:0] sel_520679;
  wire [11:0] add_520689;
  wire [11:0] sel_520691;
  wire [11:0] add_520693;
  wire [11:0] sel_520695;
  wire [11:0] add_520764;
  wire [11:0] sel_520766;
  wire [11:0] add_520769;
  wire [11:0] sel_520771;
  wire [11:0] add_520773;
  wire [11:0] add_520775;
  wire [10:0] add_520789;
  wire [11:0] sel_520791;
  wire [10:0] add_520793;
  wire [11:0] sel_520795;
  wire [10:0] add_520805;
  wire [11:0] sel_520807;
  wire [10:0] add_520809;
  wire [11:0] sel_520811;
  wire [11:0] add_520821;
  wire [11:0] sel_520823;
  wire [11:0] add_520825;
  wire [11:0] sel_520827;
  wire [11:0] add_520837;
  wire [11:0] sel_520839;
  wire [11:0] add_520841;
  wire [11:0] sel_520843;
  wire [11:0] add_520853;
  wire [11:0] sel_520855;
  wire [11:0] add_520857;
  wire [11:0] sel_520859;
  wire [8:0] add_520871;
  wire [11:0] sel_520873;
  wire [8:0] add_520875;
  wire [11:0] sel_520877;
  wire [15:0] array_index_520964;
  wire [15:0] array_index_520967;
  wire [8:0] add_520977;
  wire [11:0] sel_520979;
  wire [8:0] add_520981;
  wire [11:0] sel_520983;
  wire [11:0] add_520993;
  wire [11:0] sel_520995;
  wire [11:0] add_520997;
  wire [11:0] sel_520999;
  wire [11:0] add_521009;
  wire [11:0] sel_521011;
  wire [11:0] add_521013;
  wire [11:0] sel_521015;
  wire [11:0] add_521027;
  wire [11:0] sel_521029;
  wire [11:0] add_521031;
  wire [11:0] sel_521033;
  wire [11:0] add_521043;
  wire [11:0] sel_521045;
  wire [11:0] add_521047;
  wire [11:0] sel_521049;
  wire [10:0] add_521059;
  wire [11:0] sel_521061;
  wire [10:0] add_521063;
  wire [11:0] sel_521065;
  wire [11:0] add_521075;
  wire [11:0] sel_521077;
  wire [11:0] add_521079;
  wire [11:0] sel_521081;
  wire [8:0] add_521083;
  wire [11:0] sel_521086;
  wire [8:0] add_521088;
  wire [11:0] sel_521091;
  wire [10:0] add_521093;
  wire [11:0] sel_521095;
  wire [10:0] add_521097;
  wire [11:0] sel_521099;
  wire [9:0] add_521101;
  wire [11:0] sel_521103;
  wire [9:0] add_521105;
  wire [11:0] sel_521107;
  wire [11:0] add_521109;
  wire [11:0] sel_521111;
  wire [11:0] add_521113;
  wire [11:0] sel_521115;
  wire [10:0] add_521117;
  wire [11:0] sel_521119;
  wire [10:0] add_521121;
  wire [11:0] sel_521123;
  wire [11:0] add_521125;
  wire [11:0] sel_521127;
  wire [11:0] add_521129;
  wire [11:0] sel_521131;
  wire [11:0] add_521133;
  wire [11:0] sel_521135;
  wire [11:0] add_521137;
  wire [11:0] sel_521139;
  wire [9:0] add_521141;
  wire [11:0] sel_521144;
  wire [9:0] add_521146;
  wire [11:0] sel_521149;
  wire [11:0] add_521151;
  wire [11:0] sel_521153;
  wire [11:0] add_521155;
  wire [11:0] sel_521157;
  wire [7:0] add_521159;
  wire [11:0] sel_521162;
  wire [7:0] add_521164;
  wire [11:0] sel_521167;
  wire [11:0] add_521169;
  wire [11:0] sel_521171;
  wire [11:0] add_521173;
  wire [11:0] sel_521175;
  wire [10:0] add_521177;
  wire [11:0] sel_521179;
  wire [10:0] add_521181;
  wire [11:0] sel_521183;
  wire [10:0] add_521185;
  wire [11:0] sel_521187;
  wire [10:0] add_521189;
  wire [11:0] sel_521191;
  wire [10:0] add_521193;
  wire [11:0] sel_521196;
  wire [10:0] add_521198;
  wire [11:0] sel_521201;
  wire [8:0] add_521209;
  wire [8:0] add_521211;
  wire [11:0] add_521223;
  wire [11:0] sel_521225;
  wire [11:0] add_521227;
  wire [11:0] sel_521229;
  wire [11:0] add_521241;
  wire [11:0] sel_521243;
  wire [11:0] add_521245;
  wire [11:0] sel_521247;
  wire [10:0] add_521259;
  wire [11:0] sel_521261;
  wire [10:0] add_521263;
  wire [11:0] sel_521265;
  wire [11:0] add_521275;
  wire [11:0] sel_521277;
  wire [11:0] add_521279;
  wire [11:0] sel_521281;
  wire [11:0] add_521291;
  wire [11:0] sel_521293;
  wire [11:0] add_521295;
  wire [11:0] sel_521297;
  wire [11:0] add_521307;
  wire [11:0] sel_521309;
  wire [11:0] add_521311;
  wire [11:0] sel_521313;
  wire [11:0] add_521382;
  wire [11:0] sel_521384;
  wire [11:0] add_521387;
  wire [11:0] sel_521389;
  wire [11:0] add_521397;
  wire [11:0] sel_521399;
  wire [11:0] add_521401;
  wire [11:0] sel_521403;
  wire [10:0] add_521415;
  wire [11:0] sel_521417;
  wire [10:0] add_521419;
  wire [11:0] sel_521421;
  wire [10:0] add_521431;
  wire [11:0] sel_521433;
  wire [10:0] add_521435;
  wire [11:0] sel_521437;
  wire [11:0] add_521447;
  wire [11:0] sel_521449;
  wire [11:0] add_521451;
  wire [11:0] sel_521453;
  wire [11:0] add_521463;
  wire [11:0] sel_521465;
  wire [11:0] add_521467;
  wire [11:0] sel_521469;
  wire [11:0] add_521479;
  wire [11:0] sel_521481;
  wire [11:0] add_521483;
  wire [11:0] sel_521485;
  wire [8:0] add_521497;
  wire [11:0] sel_521499;
  wire [8:0] add_521501;
  wire [11:0] sel_521503;
  wire [15:0] array_index_521590;
  wire [15:0] array_index_521593;
  wire [8:0] add_521597;
  wire [8:0] add_521599;
  wire [8:0] add_521613;
  wire [11:0] sel_521615;
  wire [8:0] add_521617;
  wire [11:0] sel_521619;
  wire [11:0] add_521629;
  wire [11:0] sel_521631;
  wire [11:0] add_521633;
  wire [11:0] sel_521635;
  wire [11:0] add_521645;
  wire [11:0] sel_521647;
  wire [11:0] add_521649;
  wire [11:0] sel_521651;
  wire [11:0] add_521663;
  wire [11:0] sel_521665;
  wire [11:0] add_521667;
  wire [11:0] sel_521669;
  wire [11:0] add_521679;
  wire [11:0] sel_521681;
  wire [11:0] add_521683;
  wire [11:0] sel_521685;
  wire [10:0] add_521695;
  wire [11:0] sel_521697;
  wire [10:0] add_521699;
  wire [11:0] sel_521701;
  wire [11:0] add_521711;
  wire [11:0] sel_521713;
  wire [11:0] add_521715;
  wire [11:0] sel_521717;
  wire [8:0] add_521719;
  wire [11:0] sel_521722;
  wire [8:0] add_521724;
  wire [11:0] sel_521727;
  wire [10:0] add_521729;
  wire [11:0] sel_521731;
  wire [10:0] add_521733;
  wire [11:0] sel_521735;
  wire [9:0] add_521737;
  wire [11:0] sel_521739;
  wire [9:0] add_521741;
  wire [11:0] sel_521743;
  wire [11:0] add_521745;
  wire [11:0] sel_521747;
  wire [11:0] add_521749;
  wire [11:0] sel_521751;
  wire [10:0] add_521753;
  wire [11:0] sel_521755;
  wire [10:0] add_521757;
  wire [11:0] sel_521759;
  wire [11:0] add_521761;
  wire [11:0] sel_521763;
  wire [11:0] add_521765;
  wire [11:0] sel_521767;
  wire [11:0] add_521769;
  wire [11:0] sel_521771;
  wire [11:0] add_521773;
  wire [11:0] sel_521775;
  wire [9:0] add_521777;
  wire [11:0] sel_521780;
  wire [9:0] add_521782;
  wire [11:0] sel_521785;
  wire [11:0] add_521787;
  wire [11:0] sel_521789;
  wire [11:0] add_521791;
  wire [11:0] sel_521793;
  wire [7:0] add_521795;
  wire [11:0] sel_521798;
  wire [7:0] add_521800;
  wire [11:0] sel_521803;
  wire [11:0] add_521805;
  wire [11:0] sel_521807;
  wire [11:0] add_521809;
  wire [11:0] sel_521811;
  wire [10:0] add_521813;
  wire [11:0] sel_521815;
  wire [10:0] add_521817;
  wire [11:0] sel_521819;
  wire [10:0] add_521821;
  wire [11:0] sel_521823;
  wire [10:0] add_521825;
  wire [11:0] sel_521827;
  wire [10:0] add_521829;
  wire [11:0] sel_521832;
  wire [10:0] add_521834;
  wire [11:0] sel_521837;
  wire [8:0] add_521851;
  wire [11:0] sel_521853;
  wire [8:0] add_521855;
  wire [11:0] sel_521857;
  wire [11:0] add_521867;
  wire [11:0] sel_521869;
  wire [11:0] add_521871;
  wire [11:0] sel_521873;
  wire [11:0] add_521885;
  wire [11:0] sel_521887;
  wire [11:0] add_521889;
  wire [11:0] sel_521891;
  wire [10:0] add_521903;
  wire [11:0] sel_521905;
  wire [10:0] add_521907;
  wire [11:0] sel_521909;
  wire [11:0] add_521919;
  wire [11:0] sel_521921;
  wire [11:0] add_521923;
  wire [11:0] sel_521925;
  wire [11:0] add_521935;
  wire [11:0] sel_521937;
  wire [11:0] add_521939;
  wire [11:0] sel_521941;
  wire [11:0] add_521951;
  wire [11:0] sel_521953;
  wire [11:0] add_521955;
  wire [11:0] sel_521957;
  wire [11:0] add_522025;
  wire [11:0] sel_522027;
  wire [11:0] add_522029;
  wire [11:0] sel_522031;
  wire [9:0] add_522033;
  wire [9:0] add_522035;
  wire [11:0] add_522049;
  wire [11:0] sel_522051;
  wire [11:0] add_522053;
  wire [11:0] sel_522055;
  wire [10:0] add_522067;
  wire [11:0] sel_522069;
  wire [10:0] add_522071;
  wire [11:0] sel_522073;
  wire [10:0] add_522083;
  wire [11:0] sel_522085;
  wire [10:0] add_522087;
  wire [11:0] sel_522089;
  wire [11:0] add_522099;
  wire [11:0] sel_522101;
  wire [11:0] add_522103;
  wire [11:0] sel_522105;
  wire [11:0] add_522115;
  wire [11:0] sel_522117;
  wire [11:0] add_522119;
  wire [11:0] sel_522121;
  wire [11:0] add_522131;
  wire [11:0] sel_522133;
  wire [11:0] add_522135;
  wire [11:0] sel_522137;
  wire [8:0] add_522149;
  wire [11:0] sel_522151;
  wire [8:0] add_522153;
  wire [11:0] sel_522155;
  wire [8:0] add_522253;
  wire [11:0] sel_522255;
  wire [8:0] add_522257;
  wire [11:0] sel_522259;
  wire [8:0] add_522271;
  wire [11:0] sel_522273;
  wire [8:0] add_522275;
  wire [11:0] sel_522277;
  wire [11:0] add_522287;
  wire [11:0] sel_522289;
  wire [11:0] add_522291;
  wire [11:0] sel_522293;
  wire [11:0] add_522303;
  wire [11:0] sel_522305;
  wire [11:0] add_522307;
  wire [11:0] sel_522309;
  wire [11:0] add_522321;
  wire [11:0] sel_522323;
  wire [11:0] add_522325;
  wire [11:0] sel_522327;
  wire [11:0] add_522337;
  wire [11:0] sel_522339;
  wire [11:0] add_522341;
  wire [11:0] sel_522343;
  wire [10:0] add_522353;
  wire [11:0] sel_522355;
  wire [10:0] add_522357;
  wire [11:0] sel_522359;
  wire [11:0] add_522369;
  wire [11:0] sel_522371;
  wire [11:0] add_522373;
  wire [11:0] sel_522375;
  wire [8:0] add_522377;
  wire [11:0] sel_522380;
  wire [8:0] add_522382;
  wire [11:0] sel_522385;
  wire [10:0] add_522387;
  wire [11:0] sel_522389;
  wire [10:0] add_522391;
  wire [11:0] sel_522393;
  wire [9:0] add_522395;
  wire [11:0] sel_522397;
  wire [9:0] add_522399;
  wire [11:0] sel_522401;
  wire [11:0] add_522403;
  wire [11:0] sel_522405;
  wire [11:0] add_522407;
  wire [11:0] sel_522409;
  wire [10:0] add_522411;
  wire [11:0] sel_522413;
  wire [10:0] add_522415;
  wire [11:0] sel_522417;
  wire [11:0] add_522419;
  wire [11:0] sel_522421;
  wire [11:0] add_522423;
  wire [11:0] sel_522425;
  wire [11:0] add_522427;
  wire [11:0] sel_522429;
  wire [11:0] add_522431;
  wire [11:0] sel_522433;
  wire [9:0] add_522435;
  wire [11:0] sel_522438;
  wire [9:0] add_522440;
  wire [11:0] sel_522443;
  wire [11:0] add_522445;
  wire [11:0] sel_522447;
  wire [11:0] add_522449;
  wire [11:0] sel_522451;
  wire [7:0] add_522453;
  wire [11:0] sel_522456;
  wire [7:0] add_522458;
  wire [11:0] sel_522461;
  wire [11:0] add_522463;
  wire [11:0] sel_522465;
  wire [11:0] add_522467;
  wire [11:0] sel_522469;
  wire [10:0] add_522471;
  wire [11:0] sel_522473;
  wire [10:0] add_522475;
  wire [11:0] sel_522477;
  wire [10:0] add_522479;
  wire [11:0] sel_522481;
  wire [10:0] add_522483;
  wire [11:0] sel_522485;
  wire [10:0] add_522487;
  wire [11:0] sel_522490;
  wire [10:0] add_522492;
  wire [11:0] sel_522495;
  wire [11:0] add_522499;
  wire [11:0] add_522501;
  wire [8:0] add_522515;
  wire [11:0] sel_522517;
  wire [8:0] add_522519;
  wire [11:0] sel_522521;
  wire [11:0] add_522531;
  wire [11:0] sel_522533;
  wire [11:0] add_522535;
  wire [11:0] sel_522537;
  wire [11:0] add_522549;
  wire [11:0] sel_522551;
  wire [11:0] add_522553;
  wire [11:0] sel_522555;
  wire [10:0] add_522567;
  wire [11:0] sel_522569;
  wire [10:0] add_522571;
  wire [11:0] sel_522573;
  wire [11:0] add_522583;
  wire [11:0] sel_522585;
  wire [11:0] add_522587;
  wire [11:0] sel_522589;
  wire [11:0] add_522599;
  wire [11:0] sel_522601;
  wire [11:0] add_522603;
  wire [11:0] sel_522605;
  wire [11:0] add_522615;
  wire [11:0] sel_522617;
  wire [11:0] add_522619;
  wire [11:0] sel_522621;
  wire [9:0] add_522697;
  wire [11:0] sel_522699;
  wire [9:0] add_522701;
  wire [11:0] sel_522703;
  wire [11:0] add_522715;
  wire [11:0] sel_522717;
  wire [11:0] add_522719;
  wire [11:0] sel_522721;
  wire [10:0] add_522733;
  wire [11:0] sel_522735;
  wire [10:0] add_522737;
  wire [11:0] sel_522739;
  wire [10:0] add_522749;
  wire [11:0] sel_522751;
  wire [10:0] add_522753;
  wire [11:0] sel_522755;
  wire [11:0] add_522765;
  wire [11:0] sel_522767;
  wire [11:0] add_522769;
  wire [11:0] sel_522771;
  wire [11:0] add_522781;
  wire [11:0] sel_522783;
  wire [11:0] add_522785;
  wire [11:0] sel_522787;
  wire [11:0] add_522797;
  wire [11:0] sel_522799;
  wire [11:0] add_522801;
  wire [11:0] sel_522803;
  wire [8:0] add_522815;
  wire [11:0] sel_522817;
  wire [8:0] add_522819;
  wire [11:0] sel_522821;
  wire [10:0] add_522907;
  wire [10:0] add_522909;
  wire [8:0] add_522921;
  wire [11:0] sel_522923;
  wire [8:0] add_522925;
  wire [11:0] sel_522927;
  wire [8:0] add_522939;
  wire [11:0] sel_522941;
  wire [8:0] add_522943;
  wire [11:0] sel_522945;
  wire [11:0] add_522955;
  wire [11:0] sel_522957;
  wire [11:0] add_522959;
  wire [11:0] sel_522961;
  wire [11:0] add_522971;
  wire [11:0] sel_522973;
  wire [11:0] add_522975;
  wire [11:0] sel_522977;
  wire [11:0] add_522989;
  wire [11:0] sel_522991;
  wire [11:0] add_522993;
  wire [11:0] sel_522995;
  wire [11:0] add_523005;
  wire [11:0] sel_523007;
  wire [11:0] add_523009;
  wire [11:0] sel_523011;
  wire [10:0] add_523021;
  wire [11:0] sel_523023;
  wire [10:0] add_523025;
  wire [11:0] sel_523027;
  wire [11:0] add_523037;
  wire [11:0] sel_523039;
  wire [11:0] add_523041;
  wire [11:0] sel_523043;
  wire [8:0] add_523045;
  wire [11:0] sel_523048;
  wire [8:0] add_523050;
  wire [11:0] sel_523053;
  wire [10:0] add_523055;
  wire [11:0] sel_523057;
  wire [10:0] add_523059;
  wire [11:0] sel_523061;
  wire [9:0] add_523063;
  wire [11:0] sel_523065;
  wire [9:0] add_523067;
  wire [11:0] sel_523069;
  wire [11:0] add_523071;
  wire [11:0] sel_523073;
  wire [11:0] add_523075;
  wire [11:0] sel_523077;
  wire [10:0] add_523079;
  wire [11:0] sel_523081;
  wire [10:0] add_523083;
  wire [11:0] sel_523085;
  wire [11:0] add_523087;
  wire [11:0] sel_523089;
  wire [11:0] add_523091;
  wire [11:0] sel_523093;
  wire [11:0] add_523095;
  wire [11:0] sel_523097;
  wire [11:0] add_523099;
  wire [11:0] sel_523101;
  wire [9:0] add_523103;
  wire [11:0] sel_523106;
  wire [9:0] add_523108;
  wire [11:0] sel_523111;
  wire [11:0] add_523113;
  wire [11:0] sel_523115;
  wire [11:0] add_523117;
  wire [11:0] sel_523119;
  wire [7:0] add_523121;
  wire [11:0] sel_523124;
  wire [7:0] add_523126;
  wire [11:0] sel_523129;
  wire [11:0] add_523131;
  wire [11:0] sel_523133;
  wire [11:0] add_523135;
  wire [11:0] sel_523137;
  wire [10:0] add_523139;
  wire [11:0] sel_523141;
  wire [10:0] add_523143;
  wire [11:0] sel_523145;
  wire [10:0] add_523147;
  wire [11:0] sel_523149;
  wire [10:0] add_523151;
  wire [11:0] sel_523153;
  wire [1:0] concat_523156;
  wire [11:0] add_523165;
  wire [11:0] sel_523167;
  wire [11:0] add_523169;
  wire [11:0] sel_523171;
  wire [8:0] add_523183;
  wire [11:0] sel_523185;
  wire [8:0] add_523187;
  wire [11:0] sel_523189;
  wire [11:0] add_523199;
  wire [11:0] sel_523201;
  wire [11:0] add_523203;
  wire [11:0] sel_523205;
  wire [11:0] add_523217;
  wire [11:0] sel_523219;
  wire [11:0] add_523221;
  wire [11:0] sel_523223;
  wire [10:0] add_523235;
  wire [11:0] sel_523237;
  wire [10:0] add_523239;
  wire [11:0] sel_523241;
  wire [11:0] add_523251;
  wire [11:0] sel_523253;
  wire [11:0] add_523255;
  wire [11:0] sel_523257;
  wire [11:0] add_523267;
  wire [11:0] sel_523269;
  wire [11:0] add_523271;
  wire [11:0] sel_523273;
  wire [11:0] add_523283;
  wire [11:0] sel_523285;
  wire [11:0] add_523287;
  wire [11:0] sel_523289;
  wire [1:0] add_523353;
  wire [10:0] add_523355;
  wire [10:0] add_523357;
  wire [9:0] add_523371;
  wire [11:0] sel_523373;
  wire [9:0] add_523375;
  wire [11:0] sel_523377;
  wire [11:0] add_523389;
  wire [11:0] sel_523391;
  wire [11:0] add_523393;
  wire [11:0] sel_523395;
  wire [10:0] add_523407;
  wire [11:0] sel_523409;
  wire [10:0] add_523411;
  wire [11:0] sel_523413;
  wire [10:0] add_523423;
  wire [11:0] sel_523425;
  wire [10:0] add_523427;
  wire [11:0] sel_523429;
  wire [11:0] add_523439;
  wire [11:0] sel_523441;
  wire [11:0] add_523443;
  wire [11:0] sel_523445;
  wire [11:0] add_523455;
  wire [11:0] sel_523457;
  wire [11:0] add_523459;
  wire [11:0] sel_523461;
  wire [11:0] add_523471;
  wire [11:0] sel_523473;
  wire [11:0] add_523475;
  wire [11:0] sel_523477;
  wire [8:0] add_523489;
  wire [11:0] sel_523491;
  wire [8:0] add_523493;
  wire [11:0] sel_523495;
  wire [10:0] add_523581;
  wire [11:0] sel_523583;
  wire [10:0] add_523585;
  wire [11:0] sel_523587;
  wire [8:0] add_523597;
  wire [11:0] sel_523599;
  wire [8:0] add_523601;
  wire [11:0] sel_523603;
  wire [8:0] add_523615;
  wire [11:0] sel_523617;
  wire [8:0] add_523619;
  wire [11:0] sel_523621;
  wire [11:0] add_523631;
  wire [11:0] sel_523633;
  wire [11:0] add_523635;
  wire [11:0] sel_523637;
  wire [11:0] add_523647;
  wire [11:0] sel_523649;
  wire [11:0] add_523651;
  wire [11:0] sel_523653;
  wire [11:0] add_523665;
  wire [11:0] sel_523667;
  wire [11:0] add_523669;
  wire [11:0] sel_523671;
  wire [11:0] add_523681;
  wire [11:0] sel_523683;
  wire [11:0] add_523685;
  wire [11:0] sel_523687;
  wire [10:0] add_523697;
  wire [11:0] sel_523699;
  wire [10:0] add_523701;
  wire [11:0] sel_523703;
  wire [11:0] add_523713;
  wire [11:0] sel_523715;
  wire [11:0] add_523717;
  wire [11:0] sel_523719;
  wire [8:0] add_523721;
  wire [11:0] sel_523724;
  wire [8:0] add_523726;
  wire [11:0] sel_523729;
  wire [10:0] add_523731;
  wire [11:0] sel_523733;
  wire [10:0] add_523735;
  wire [11:0] sel_523737;
  wire [9:0] add_523739;
  wire [11:0] sel_523741;
  wire [9:0] add_523743;
  wire [11:0] sel_523745;
  wire [11:0] add_523747;
  wire [11:0] sel_523749;
  wire [11:0] add_523751;
  wire [11:0] sel_523753;
  wire [10:0] add_523755;
  wire [11:0] sel_523757;
  wire [10:0] add_523759;
  wire [11:0] sel_523761;
  wire [11:0] add_523763;
  wire [11:0] sel_523765;
  wire [11:0] add_523767;
  wire [11:0] sel_523769;
  wire [11:0] add_523771;
  wire [11:0] sel_523773;
  wire [11:0] add_523775;
  wire [11:0] sel_523777;
  wire [9:0] add_523779;
  wire [11:0] sel_523782;
  wire [9:0] add_523784;
  wire [11:0] sel_523787;
  wire [11:0] add_523789;
  wire [11:0] sel_523791;
  wire [11:0] add_523793;
  wire [11:0] sel_523795;
  wire [7:0] add_523797;
  wire [11:0] sel_523800;
  wire [7:0] add_523802;
  wire [11:0] sel_523805;
  wire [11:0] add_523807;
  wire [11:0] sel_523809;
  wire [11:0] add_523811;
  wire [11:0] sel_523813;
  wire [10:0] add_523815;
  wire [11:0] sel_523817;
  wire [10:0] add_523819;
  wire [11:0] sel_523821;
  wire [2:0] concat_523824;
  wire [11:0] add_523827;
  wire [11:0] add_523829;
  wire [11:0] add_523843;
  wire [11:0] sel_523845;
  wire [11:0] add_523847;
  wire [11:0] sel_523849;
  wire [8:0] add_523861;
  wire [11:0] sel_523863;
  wire [8:0] add_523865;
  wire [11:0] sel_523867;
  wire [11:0] add_523877;
  wire [11:0] sel_523879;
  wire [11:0] add_523881;
  wire [11:0] sel_523883;
  wire [11:0] add_523895;
  wire [11:0] sel_523897;
  wire [11:0] add_523899;
  wire [11:0] sel_523901;
  wire [10:0] add_523913;
  wire [11:0] sel_523915;
  wire [10:0] add_523917;
  wire [11:0] sel_523919;
  wire [11:0] add_523929;
  wire [11:0] sel_523931;
  wire [11:0] add_523933;
  wire [11:0] sel_523935;
  wire [11:0] add_523945;
  wire [11:0] sel_523947;
  wire [11:0] add_523949;
  wire [11:0] sel_523951;
  wire [11:0] add_523961;
  wire [11:0] sel_523963;
  wire [11:0] add_523965;
  wire [11:0] sel_523967;
  wire [2:0] add_524027;
  wire [10:0] add_524035;
  wire [11:0] sel_524037;
  wire [10:0] add_524039;
  wire [11:0] sel_524041;
  wire [9:0] add_524053;
  wire [11:0] sel_524055;
  wire [9:0] add_524057;
  wire [11:0] sel_524059;
  wire [11:0] add_524071;
  wire [11:0] sel_524073;
  wire [11:0] add_524075;
  wire [11:0] sel_524077;
  wire [10:0] add_524089;
  wire [11:0] sel_524091;
  wire [10:0] add_524093;
  wire [11:0] sel_524095;
  wire [10:0] add_524105;
  wire [11:0] sel_524107;
  wire [10:0] add_524109;
  wire [11:0] sel_524111;
  wire [11:0] add_524121;
  wire [11:0] sel_524123;
  wire [11:0] add_524125;
  wire [11:0] sel_524127;
  wire [11:0] add_524137;
  wire [11:0] sel_524139;
  wire [11:0] add_524141;
  wire [11:0] sel_524143;
  wire [11:0] add_524153;
  wire [11:0] sel_524155;
  wire [11:0] add_524157;
  wire [11:0] sel_524159;
  wire [8:0] add_524171;
  wire [11:0] sel_524173;
  wire [8:0] add_524175;
  wire [11:0] sel_524177;
  wire [11:0] add_524251;
  wire [11:0] add_524253;
  wire [10:0] add_524265;
  wire [11:0] sel_524267;
  wire [10:0] add_524269;
  wire [11:0] sel_524271;
  wire [8:0] add_524281;
  wire [11:0] sel_524283;
  wire [8:0] add_524285;
  wire [11:0] sel_524287;
  wire [8:0] add_524299;
  wire [11:0] sel_524301;
  wire [8:0] add_524303;
  wire [11:0] sel_524305;
  wire [11:0] add_524315;
  wire [11:0] sel_524317;
  wire [11:0] add_524319;
  wire [11:0] sel_524321;
  wire [11:0] add_524331;
  wire [11:0] sel_524333;
  wire [11:0] add_524335;
  wire [11:0] sel_524337;
  wire [11:0] add_524349;
  wire [11:0] sel_524351;
  wire [11:0] add_524353;
  wire [11:0] sel_524355;
  wire [11:0] add_524365;
  wire [11:0] sel_524367;
  wire [11:0] add_524369;
  wire [11:0] sel_524371;
  wire [10:0] add_524381;
  wire [11:0] sel_524383;
  wire [10:0] add_524385;
  wire [11:0] sel_524387;
  wire [11:0] add_524397;
  wire [11:0] sel_524399;
  wire [11:0] add_524401;
  wire [11:0] sel_524403;
  wire [8:0] add_524405;
  wire [11:0] sel_524408;
  wire [8:0] add_524410;
  wire [11:0] sel_524413;
  wire [10:0] add_524415;
  wire [11:0] sel_524417;
  wire [10:0] add_524419;
  wire [11:0] sel_524421;
  wire [9:0] add_524423;
  wire [11:0] sel_524425;
  wire [9:0] add_524427;
  wire [11:0] sel_524429;
  wire [11:0] add_524431;
  wire [11:0] sel_524433;
  wire [11:0] add_524435;
  wire [11:0] sel_524437;
  wire [10:0] add_524439;
  wire [11:0] sel_524441;
  wire [10:0] add_524443;
  wire [11:0] sel_524445;
  wire [11:0] add_524447;
  wire [11:0] sel_524449;
  wire [11:0] add_524451;
  wire [11:0] sel_524453;
  wire [11:0] add_524455;
  wire [11:0] sel_524457;
  wire [11:0] add_524459;
  wire [11:0] sel_524461;
  wire [9:0] add_524463;
  wire [11:0] sel_524466;
  wire [9:0] add_524468;
  wire [11:0] sel_524471;
  wire [11:0] add_524473;
  wire [11:0] sel_524475;
  wire [11:0] add_524477;
  wire [11:0] sel_524479;
  wire [7:0] add_524481;
  wire [11:0] sel_524484;
  wire [7:0] add_524486;
  wire [11:0] sel_524489;
  wire [11:0] add_524491;
  wire [11:0] sel_524493;
  wire [11:0] add_524495;
  wire [11:0] sel_524497;
  wire [3:0] concat_524500;
  wire [11:0] add_524509;
  wire [11:0] sel_524511;
  wire [11:0] add_524513;
  wire [11:0] sel_524515;
  wire [11:0] add_524527;
  wire [11:0] sel_524529;
  wire [11:0] add_524531;
  wire [11:0] sel_524533;
  wire [8:0] add_524545;
  wire [11:0] sel_524547;
  wire [8:0] add_524549;
  wire [11:0] sel_524551;
  wire [11:0] add_524561;
  wire [11:0] sel_524563;
  wire [11:0] add_524565;
  wire [11:0] sel_524567;
  wire [11:0] add_524579;
  wire [11:0] sel_524581;
  wire [11:0] add_524583;
  wire [11:0] sel_524585;
  wire [10:0] add_524597;
  wire [11:0] sel_524599;
  wire [10:0] add_524601;
  wire [11:0] sel_524603;
  wire [11:0] add_524613;
  wire [11:0] sel_524615;
  wire [11:0] add_524617;
  wire [11:0] sel_524619;
  wire [11:0] add_524629;
  wire [11:0] sel_524631;
  wire [11:0] add_524633;
  wire [11:0] sel_524635;
  wire [11:0] add_524645;
  wire [11:0] sel_524647;
  wire [11:0] add_524649;
  wire [11:0] sel_524651;
  wire [3:0] add_524707;
  wire [10:0] add_524709;
  wire [10:0] add_524711;
  wire [10:0] add_524723;
  wire [11:0] sel_524725;
  wire [10:0] add_524727;
  wire [11:0] sel_524729;
  wire [9:0] add_524741;
  wire [11:0] sel_524743;
  wire [9:0] add_524745;
  wire [11:0] sel_524747;
  wire [11:0] add_524759;
  wire [11:0] sel_524761;
  wire [11:0] add_524763;
  wire [11:0] sel_524765;
  wire [10:0] add_524777;
  wire [11:0] sel_524779;
  wire [10:0] add_524781;
  wire [11:0] sel_524783;
  wire [10:0] add_524793;
  wire [11:0] sel_524795;
  wire [10:0] add_524797;
  wire [11:0] sel_524799;
  wire [11:0] add_524809;
  wire [11:0] sel_524811;
  wire [11:0] add_524813;
  wire [11:0] sel_524815;
  wire [11:0] add_524825;
  wire [11:0] sel_524827;
  wire [11:0] add_524829;
  wire [11:0] sel_524831;
  wire [11:0] add_524841;
  wire [11:0] sel_524843;
  wire [11:0] add_524845;
  wire [11:0] sel_524847;
  wire [8:0] add_524859;
  wire [11:0] sel_524861;
  wire [8:0] add_524863;
  wire [11:0] sel_524865;
  wire [11:0] add_524939;
  wire [11:0] sel_524941;
  wire [11:0] add_524943;
  wire [11:0] sel_524945;
  wire [10:0] add_524955;
  wire [11:0] sel_524957;
  wire [10:0] add_524959;
  wire [11:0] sel_524961;
  wire [8:0] add_524971;
  wire [11:0] sel_524973;
  wire [8:0] add_524975;
  wire [11:0] sel_524977;
  wire [8:0] add_524989;
  wire [11:0] sel_524991;
  wire [8:0] add_524993;
  wire [11:0] sel_524995;
  wire [11:0] add_525005;
  wire [11:0] sel_525007;
  wire [11:0] add_525009;
  wire [11:0] sel_525011;
  wire [11:0] add_525021;
  wire [11:0] sel_525023;
  wire [11:0] add_525025;
  wire [11:0] sel_525027;
  wire [11:0] add_525039;
  wire [11:0] sel_525041;
  wire [11:0] add_525043;
  wire [11:0] sel_525045;
  wire [11:0] add_525055;
  wire [11:0] sel_525057;
  wire [11:0] add_525059;
  wire [11:0] sel_525061;
  wire [10:0] add_525071;
  wire [11:0] sel_525073;
  wire [10:0] add_525075;
  wire [11:0] sel_525077;
  wire [11:0] add_525087;
  wire [11:0] sel_525089;
  wire [11:0] add_525091;
  wire [11:0] sel_525093;
  wire [8:0] add_525095;
  wire [11:0] sel_525098;
  wire [8:0] add_525100;
  wire [11:0] sel_525103;
  wire [10:0] add_525105;
  wire [11:0] sel_525107;
  wire [10:0] add_525109;
  wire [11:0] sel_525111;
  wire [9:0] add_525113;
  wire [11:0] sel_525115;
  wire [9:0] add_525117;
  wire [11:0] sel_525119;
  wire [11:0] add_525121;
  wire [11:0] sel_525123;
  wire [11:0] add_525125;
  wire [11:0] sel_525127;
  wire [10:0] add_525129;
  wire [11:0] sel_525131;
  wire [10:0] add_525133;
  wire [11:0] sel_525135;
  wire [11:0] add_525137;
  wire [11:0] sel_525139;
  wire [11:0] add_525141;
  wire [11:0] sel_525143;
  wire [11:0] add_525145;
  wire [11:0] sel_525147;
  wire [11:0] add_525149;
  wire [11:0] sel_525151;
  wire [9:0] add_525153;
  wire [11:0] sel_525156;
  wire [9:0] add_525158;
  wire [11:0] sel_525161;
  wire [11:0] add_525163;
  wire [11:0] sel_525165;
  wire [11:0] add_525167;
  wire [11:0] sel_525169;
  wire [7:0] add_525171;
  wire [11:0] sel_525174;
  wire [7:0] add_525176;
  wire [11:0] sel_525179;
  wire [4:0] concat_525182;
  wire [11:0] add_525185;
  wire [11:0] add_525187;
  wire [11:0] add_525201;
  wire [11:0] sel_525203;
  wire [11:0] add_525205;
  wire [11:0] sel_525207;
  wire [11:0] add_525219;
  wire [11:0] sel_525221;
  wire [11:0] add_525223;
  wire [11:0] sel_525225;
  wire [8:0] add_525237;
  wire [11:0] sel_525239;
  wire [8:0] add_525241;
  wire [11:0] sel_525243;
  wire [11:0] add_525253;
  wire [11:0] sel_525255;
  wire [11:0] add_525257;
  wire [11:0] sel_525259;
  wire [11:0] add_525271;
  wire [11:0] sel_525273;
  wire [11:0] add_525275;
  wire [11:0] sel_525277;
  wire [10:0] add_525289;
  wire [11:0] sel_525291;
  wire [10:0] add_525293;
  wire [11:0] sel_525295;
  wire [11:0] add_525305;
  wire [11:0] sel_525307;
  wire [11:0] add_525309;
  wire [11:0] sel_525311;
  wire [11:0] add_525321;
  wire [11:0] sel_525323;
  wire [11:0] add_525325;
  wire [11:0] sel_525327;
  wire [11:0] add_525337;
  wire [11:0] sel_525339;
  wire [11:0] add_525341;
  wire [11:0] sel_525343;
  wire [4:0] add_525395;
  wire [10:0] add_525403;
  wire [11:0] sel_525405;
  wire [10:0] add_525407;
  wire [11:0] sel_525409;
  wire [10:0] add_525419;
  wire [11:0] sel_525421;
  wire [10:0] add_525423;
  wire [11:0] sel_525425;
  wire [9:0] add_525437;
  wire [11:0] sel_525439;
  wire [9:0] add_525441;
  wire [11:0] sel_525443;
  wire [11:0] add_525455;
  wire [11:0] sel_525457;
  wire [11:0] add_525459;
  wire [11:0] sel_525461;
  wire [10:0] add_525473;
  wire [11:0] sel_525475;
  wire [10:0] add_525477;
  wire [11:0] sel_525479;
  wire [10:0] add_525489;
  wire [11:0] sel_525491;
  wire [10:0] add_525493;
  wire [11:0] sel_525495;
  wire [11:0] add_525505;
  wire [11:0] sel_525507;
  wire [11:0] add_525509;
  wire [11:0] sel_525511;
  wire [11:0] add_525521;
  wire [11:0] sel_525523;
  wire [11:0] add_525525;
  wire [11:0] sel_525527;
  wire [11:0] add_525537;
  wire [11:0] sel_525539;
  wire [11:0] add_525541;
  wire [11:0] sel_525543;
  wire [8:0] add_525555;
  wire [11:0] sel_525557;
  wire [8:0] add_525559;
  wire [11:0] sel_525561;
  wire [7:0] add_525623;
  wire [7:0] add_525625;
  wire [11:0] add_525637;
  wire [11:0] sel_525639;
  wire [11:0] add_525641;
  wire [11:0] sel_525643;
  wire [10:0] add_525653;
  wire [11:0] sel_525655;
  wire [10:0] add_525657;
  wire [11:0] sel_525659;
  wire [8:0] add_525669;
  wire [11:0] sel_525671;
  wire [8:0] add_525673;
  wire [11:0] sel_525675;
  wire [8:0] add_525687;
  wire [11:0] sel_525689;
  wire [8:0] add_525691;
  wire [11:0] sel_525693;
  wire [11:0] add_525703;
  wire [11:0] sel_525705;
  wire [11:0] add_525707;
  wire [11:0] sel_525709;
  wire [11:0] add_525719;
  wire [11:0] sel_525721;
  wire [11:0] add_525723;
  wire [11:0] sel_525725;
  wire [11:0] add_525737;
  wire [11:0] sel_525739;
  wire [11:0] add_525741;
  wire [11:0] sel_525743;
  wire [11:0] add_525753;
  wire [11:0] sel_525755;
  wire [11:0] add_525757;
  wire [11:0] sel_525759;
  wire [10:0] add_525769;
  wire [11:0] sel_525771;
  wire [10:0] add_525773;
  wire [11:0] sel_525775;
  wire [11:0] add_525785;
  wire [11:0] sel_525787;
  wire [11:0] add_525789;
  wire [11:0] sel_525791;
  wire [8:0] add_525793;
  wire [11:0] sel_525796;
  wire [8:0] add_525798;
  wire [11:0] sel_525801;
  wire [10:0] add_525803;
  wire [11:0] sel_525805;
  wire [10:0] add_525807;
  wire [11:0] sel_525809;
  wire [9:0] add_525811;
  wire [11:0] sel_525813;
  wire [9:0] add_525815;
  wire [11:0] sel_525817;
  wire [11:0] add_525819;
  wire [11:0] sel_525821;
  wire [11:0] add_525823;
  wire [11:0] sel_525825;
  wire [10:0] add_525827;
  wire [11:0] sel_525829;
  wire [10:0] add_525831;
  wire [11:0] sel_525833;
  wire [11:0] add_525835;
  wire [11:0] sel_525837;
  wire [11:0] add_525839;
  wire [11:0] sel_525841;
  wire [11:0] add_525843;
  wire [11:0] sel_525845;
  wire [11:0] add_525847;
  wire [11:0] sel_525849;
  wire [9:0] add_525851;
  wire [11:0] sel_525854;
  wire [9:0] add_525856;
  wire [11:0] sel_525859;
  wire [11:0] add_525861;
  wire [11:0] sel_525863;
  wire [11:0] add_525865;
  wire [11:0] sel_525867;
  wire [5:0] concat_525870;
  wire [11:0] add_525879;
  wire [11:0] sel_525881;
  wire [11:0] add_525883;
  wire [11:0] sel_525885;
  wire [11:0] add_525897;
  wire [11:0] sel_525899;
  wire [11:0] add_525901;
  wire [11:0] sel_525903;
  wire [11:0] add_525915;
  wire [11:0] sel_525917;
  wire [11:0] add_525919;
  wire [11:0] sel_525921;
  wire [8:0] add_525933;
  wire [11:0] sel_525935;
  wire [8:0] add_525937;
  wire [11:0] sel_525939;
  wire [11:0] add_525949;
  wire [11:0] sel_525951;
  wire [11:0] add_525953;
  wire [11:0] sel_525955;
  wire [11:0] add_525967;
  wire [11:0] sel_525969;
  wire [11:0] add_525971;
  wire [11:0] sel_525973;
  wire [10:0] add_525985;
  wire [11:0] sel_525987;
  wire [10:0] add_525989;
  wire [11:0] sel_525991;
  wire [11:0] add_526001;
  wire [11:0] sel_526003;
  wire [11:0] add_526005;
  wire [11:0] sel_526007;
  wire [11:0] add_526017;
  wire [11:0] sel_526019;
  wire [11:0] add_526021;
  wire [11:0] sel_526023;
  wire [11:0] add_526033;
  wire [11:0] sel_526035;
  wire [11:0] add_526037;
  wire [11:0] sel_526039;
  wire [5:0] add_526087;
  wire [11:0] add_526089;
  wire [11:0] add_526091;
  wire [10:0] add_526105;
  wire [11:0] sel_526107;
  wire [10:0] add_526109;
  wire [11:0] sel_526111;
  wire [10:0] add_526121;
  wire [11:0] sel_526123;
  wire [10:0] add_526125;
  wire [11:0] sel_526127;
  wire [9:0] add_526139;
  wire [11:0] sel_526141;
  wire [9:0] add_526143;
  wire [11:0] sel_526145;
  wire [11:0] add_526157;
  wire [11:0] sel_526159;
  wire [11:0] add_526161;
  wire [11:0] sel_526163;
  wire [10:0] add_526175;
  wire [11:0] sel_526177;
  wire [10:0] add_526179;
  wire [11:0] sel_526181;
  wire [10:0] add_526191;
  wire [11:0] sel_526193;
  wire [10:0] add_526195;
  wire [11:0] sel_526197;
  wire [11:0] add_526207;
  wire [11:0] sel_526209;
  wire [11:0] add_526211;
  wire [11:0] sel_526213;
  wire [11:0] add_526223;
  wire [11:0] sel_526225;
  wire [11:0] add_526227;
  wire [11:0] sel_526229;
  wire [11:0] add_526239;
  wire [11:0] sel_526241;
  wire [11:0] add_526243;
  wire [11:0] sel_526245;
  wire [8:0] add_526257;
  wire [11:0] sel_526259;
  wire [8:0] add_526261;
  wire [11:0] sel_526263;
  wire [7:0] add_526325;
  wire [11:0] sel_526327;
  wire [7:0] add_526329;
  wire [11:0] sel_526331;
  wire [11:0] add_526341;
  wire [11:0] sel_526343;
  wire [11:0] add_526345;
  wire [11:0] sel_526347;
  wire [10:0] add_526357;
  wire [11:0] sel_526359;
  wire [10:0] add_526361;
  wire [11:0] sel_526363;
  wire [8:0] add_526373;
  wire [11:0] sel_526375;
  wire [8:0] add_526377;
  wire [11:0] sel_526379;
  wire [8:0] add_526391;
  wire [11:0] sel_526393;
  wire [8:0] add_526395;
  wire [11:0] sel_526397;
  wire [11:0] add_526407;
  wire [11:0] sel_526409;
  wire [11:0] add_526411;
  wire [11:0] sel_526413;
  wire [11:0] add_526423;
  wire [11:0] sel_526425;
  wire [11:0] add_526427;
  wire [11:0] sel_526429;
  wire [11:0] add_526441;
  wire [11:0] sel_526443;
  wire [11:0] add_526445;
  wire [11:0] sel_526447;
  wire [11:0] add_526457;
  wire [11:0] sel_526459;
  wire [11:0] add_526461;
  wire [11:0] sel_526463;
  wire [10:0] add_526473;
  wire [11:0] sel_526475;
  wire [10:0] add_526477;
  wire [11:0] sel_526479;
  wire [11:0] add_526489;
  wire [11:0] sel_526491;
  wire [11:0] add_526493;
  wire [11:0] sel_526495;
  wire [8:0] add_526497;
  wire [11:0] sel_526500;
  wire [8:0] add_526502;
  wire [11:0] sel_526505;
  wire [10:0] add_526507;
  wire [11:0] sel_526509;
  wire [10:0] add_526511;
  wire [11:0] sel_526513;
  wire [9:0] add_526515;
  wire [11:0] sel_526517;
  wire [9:0] add_526519;
  wire [11:0] sel_526521;
  wire [11:0] add_526523;
  wire [11:0] sel_526525;
  wire [11:0] add_526527;
  wire [11:0] sel_526529;
  wire [10:0] add_526531;
  wire [11:0] sel_526533;
  wire [10:0] add_526535;
  wire [11:0] sel_526537;
  wire [11:0] add_526539;
  wire [11:0] sel_526541;
  wire [11:0] add_526543;
  wire [11:0] sel_526545;
  wire [11:0] add_526547;
  wire [11:0] sel_526549;
  wire [11:0] add_526551;
  wire [11:0] sel_526553;
  wire [9:0] add_526555;
  wire [11:0] sel_526558;
  wire [9:0] add_526560;
  wire [11:0] sel_526563;
  wire [6:0] concat_526566;
  wire [10:0] add_526569;
  wire [10:0] add_526571;
  wire [11:0] add_526583;
  wire [11:0] sel_526585;
  wire [11:0] add_526587;
  wire [11:0] sel_526589;
  wire [11:0] add_526601;
  wire [11:0] sel_526603;
  wire [11:0] add_526605;
  wire [11:0] sel_526607;
  wire [11:0] add_526619;
  wire [11:0] sel_526621;
  wire [11:0] add_526623;
  wire [11:0] sel_526625;
  wire [8:0] add_526637;
  wire [11:0] sel_526639;
  wire [8:0] add_526641;
  wire [11:0] sel_526643;
  wire [11:0] add_526653;
  wire [11:0] sel_526655;
  wire [11:0] add_526657;
  wire [11:0] sel_526659;
  wire [11:0] add_526671;
  wire [11:0] sel_526673;
  wire [11:0] add_526675;
  wire [11:0] sel_526677;
  wire [10:0] add_526689;
  wire [11:0] sel_526691;
  wire [10:0] add_526693;
  wire [11:0] sel_526695;
  wire [11:0] add_526705;
  wire [11:0] sel_526707;
  wire [11:0] add_526709;
  wire [11:0] sel_526711;
  wire [11:0] add_526721;
  wire [11:0] sel_526723;
  wire [11:0] add_526725;
  wire [11:0] sel_526727;
  wire [11:0] add_526737;
  wire [11:0] sel_526739;
  wire [11:0] add_526741;
  wire [11:0] sel_526743;
  wire [6:0] add_526787;
  wire [11:0] add_526795;
  wire [11:0] sel_526797;
  wire [11:0] add_526799;
  wire [11:0] sel_526801;
  wire [10:0] add_526813;
  wire [11:0] sel_526815;
  wire [10:0] add_526817;
  wire [11:0] sel_526819;
  wire [10:0] add_526829;
  wire [11:0] sel_526831;
  wire [10:0] add_526833;
  wire [11:0] sel_526835;
  wire [9:0] add_526847;
  wire [11:0] sel_526849;
  wire [9:0] add_526851;
  wire [11:0] sel_526853;
  wire [11:0] add_526865;
  wire [11:0] sel_526867;
  wire [11:0] add_526869;
  wire [11:0] sel_526871;
  wire [10:0] add_526883;
  wire [11:0] sel_526885;
  wire [10:0] add_526887;
  wire [11:0] sel_526889;
  wire [10:0] add_526899;
  wire [11:0] sel_526901;
  wire [10:0] add_526903;
  wire [11:0] sel_526905;
  wire [11:0] add_526915;
  wire [11:0] sel_526917;
  wire [11:0] add_526919;
  wire [11:0] sel_526921;
  wire [11:0] add_526931;
  wire [11:0] sel_526933;
  wire [11:0] add_526935;
  wire [11:0] sel_526937;
  wire [11:0] add_526947;
  wire [11:0] sel_526949;
  wire [11:0] add_526951;
  wire [11:0] sel_526953;
  wire [8:0] add_526965;
  wire [11:0] sel_526967;
  wire [8:0] add_526969;
  wire [11:0] sel_526971;
  wire [9:0] add_527021;
  wire [9:0] add_527023;
  wire [7:0] add_527037;
  wire [11:0] sel_527039;
  wire [7:0] add_527041;
  wire [11:0] sel_527043;
  wire [11:0] add_527053;
  wire [11:0] sel_527055;
  wire [11:0] add_527057;
  wire [11:0] sel_527059;
  wire [10:0] add_527069;
  wire [11:0] sel_527071;
  wire [10:0] add_527073;
  wire [11:0] sel_527075;
  wire [8:0] add_527085;
  wire [11:0] sel_527087;
  wire [8:0] add_527089;
  wire [11:0] sel_527091;
  wire [8:0] add_527103;
  wire [11:0] sel_527105;
  wire [8:0] add_527107;
  wire [11:0] sel_527109;
  wire [11:0] add_527119;
  wire [11:0] sel_527121;
  wire [11:0] add_527123;
  wire [11:0] sel_527125;
  wire [11:0] add_527135;
  wire [11:0] sel_527137;
  wire [11:0] add_527139;
  wire [11:0] sel_527141;
  wire [11:0] add_527153;
  wire [11:0] sel_527155;
  wire [11:0] add_527157;
  wire [11:0] sel_527159;
  wire [11:0] add_527169;
  wire [11:0] sel_527171;
  wire [11:0] add_527173;
  wire [11:0] sel_527175;
  wire [10:0] add_527185;
  wire [11:0] sel_527187;
  wire [10:0] add_527189;
  wire [11:0] sel_527191;
  wire [11:0] add_527201;
  wire [11:0] sel_527203;
  wire [11:0] add_527205;
  wire [11:0] sel_527207;
  wire [8:0] add_527209;
  wire [11:0] sel_527212;
  wire [8:0] add_527214;
  wire [11:0] sel_527217;
  wire [10:0] add_527219;
  wire [11:0] sel_527221;
  wire [10:0] add_527223;
  wire [11:0] sel_527225;
  wire [9:0] add_527227;
  wire [11:0] sel_527229;
  wire [9:0] add_527231;
  wire [11:0] sel_527233;
  wire [11:0] add_527235;
  wire [11:0] sel_527237;
  wire [11:0] add_527239;
  wire [11:0] sel_527241;
  wire [10:0] add_527243;
  wire [11:0] sel_527245;
  wire [10:0] add_527247;
  wire [11:0] sel_527249;
  wire [11:0] add_527251;
  wire [11:0] sel_527253;
  wire [11:0] add_527255;
  wire [11:0] sel_527257;
  wire [11:0] add_527259;
  wire [11:0] sel_527261;
  wire [11:0] add_527263;
  wire [11:0] sel_527265;
  wire [7:0] concat_527268;
  wire [10:0] add_527277;
  wire [11:0] sel_527279;
  wire [10:0] add_527281;
  wire [11:0] sel_527283;
  wire [11:0] add_527293;
  wire [11:0] sel_527295;
  wire [11:0] add_527297;
  wire [11:0] sel_527299;
  wire [11:0] add_527311;
  wire [11:0] sel_527313;
  wire [11:0] add_527315;
  wire [11:0] sel_527317;
  wire [11:0] add_527329;
  wire [11:0] sel_527331;
  wire [11:0] add_527333;
  wire [11:0] sel_527335;
  wire [8:0] add_527347;
  wire [11:0] sel_527349;
  wire [8:0] add_527351;
  wire [11:0] sel_527353;
  wire [11:0] add_527363;
  wire [11:0] sel_527365;
  wire [11:0] add_527367;
  wire [11:0] sel_527369;
  wire [11:0] add_527381;
  wire [11:0] sel_527383;
  wire [11:0] add_527385;
  wire [11:0] sel_527387;
  wire [10:0] add_527399;
  wire [11:0] sel_527401;
  wire [10:0] add_527403;
  wire [11:0] sel_527405;
  wire [11:0] add_527415;
  wire [11:0] sel_527417;
  wire [11:0] add_527419;
  wire [11:0] sel_527421;
  wire [11:0] add_527431;
  wire [11:0] sel_527433;
  wire [11:0] add_527435;
  wire [11:0] sel_527437;
  wire [11:0] add_527447;
  wire [11:0] sel_527449;
  wire [11:0] add_527451;
  wire [11:0] sel_527453;
  wire [7:0] add_527493;
  wire [11:0] add_527495;
  wire [11:0] add_527497;
  wire [11:0] add_527511;
  wire [11:0] sel_527513;
  wire [11:0] add_527515;
  wire [11:0] sel_527517;
  wire [10:0] add_527529;
  wire [11:0] sel_527531;
  wire [10:0] add_527533;
  wire [11:0] sel_527535;
  wire [10:0] add_527545;
  wire [11:0] sel_527547;
  wire [10:0] add_527549;
  wire [11:0] sel_527551;
  wire [9:0] add_527563;
  wire [11:0] sel_527565;
  wire [9:0] add_527567;
  wire [11:0] sel_527569;
  wire [11:0] add_527581;
  wire [11:0] sel_527583;
  wire [11:0] add_527585;
  wire [11:0] sel_527587;
  wire [10:0] add_527599;
  wire [11:0] sel_527601;
  wire [10:0] add_527603;
  wire [11:0] sel_527605;
  wire [10:0] add_527615;
  wire [11:0] sel_527617;
  wire [10:0] add_527619;
  wire [11:0] sel_527621;
  wire [11:0] add_527631;
  wire [11:0] sel_527633;
  wire [11:0] add_527635;
  wire [11:0] sel_527637;
  wire [11:0] add_527647;
  wire [11:0] sel_527649;
  wire [11:0] add_527651;
  wire [11:0] sel_527653;
  wire [11:0] add_527663;
  wire [11:0] sel_527665;
  wire [11:0] add_527667;
  wire [11:0] sel_527669;
  wire [8:0] add_527681;
  wire [11:0] sel_527683;
  wire [8:0] add_527685;
  wire [11:0] sel_527687;
  wire [9:0] add_527735;
  wire [11:0] sel_527737;
  wire [9:0] add_527739;
  wire [11:0] sel_527741;
  wire [7:0] add_527753;
  wire [11:0] sel_527755;
  wire [7:0] add_527757;
  wire [11:0] sel_527759;
  wire [11:0] add_527769;
  wire [11:0] sel_527771;
  wire [11:0] add_527773;
  wire [11:0] sel_527775;
  wire [10:0] add_527785;
  wire [11:0] sel_527787;
  wire [10:0] add_527789;
  wire [11:0] sel_527791;
  wire [8:0] add_527801;
  wire [11:0] sel_527803;
  wire [8:0] add_527805;
  wire [11:0] sel_527807;
  wire [8:0] add_527819;
  wire [11:0] sel_527821;
  wire [8:0] add_527823;
  wire [11:0] sel_527825;
  wire [11:0] add_527835;
  wire [11:0] sel_527837;
  wire [11:0] add_527839;
  wire [11:0] sel_527841;
  wire [11:0] add_527851;
  wire [11:0] sel_527853;
  wire [11:0] add_527855;
  wire [11:0] sel_527857;
  wire [11:0] add_527869;
  wire [11:0] sel_527871;
  wire [11:0] add_527873;
  wire [11:0] sel_527875;
  wire [11:0] add_527885;
  wire [11:0] sel_527887;
  wire [11:0] add_527889;
  wire [11:0] sel_527891;
  wire [10:0] add_527901;
  wire [11:0] sel_527903;
  wire [10:0] add_527905;
  wire [11:0] sel_527907;
  wire [11:0] add_527917;
  wire [11:0] sel_527919;
  wire [11:0] add_527921;
  wire [11:0] sel_527923;
  wire [8:0] add_527925;
  wire [11:0] sel_527928;
  wire [8:0] add_527930;
  wire [11:0] sel_527933;
  wire [10:0] add_527935;
  wire [11:0] sel_527937;
  wire [10:0] add_527939;
  wire [11:0] sel_527941;
  wire [9:0] add_527943;
  wire [11:0] sel_527945;
  wire [9:0] add_527947;
  wire [11:0] sel_527949;
  wire [11:0] add_527951;
  wire [11:0] sel_527953;
  wire [11:0] add_527955;
  wire [11:0] sel_527957;
  wire [10:0] add_527959;
  wire [11:0] sel_527961;
  wire [10:0] add_527963;
  wire [11:0] sel_527965;
  wire [11:0] add_527967;
  wire [11:0] sel_527969;
  wire [11:0] add_527971;
  wire [11:0] sel_527973;
  wire [8:0] concat_527976;
  wire [10:0] add_527989;
  wire [11:0] sel_527991;
  wire [10:0] add_527993;
  wire [11:0] sel_527995;
  wire [11:0] add_528005;
  wire [11:0] sel_528007;
  wire [11:0] add_528009;
  wire [11:0] sel_528011;
  wire [11:0] add_528023;
  wire [11:0] sel_528025;
  wire [11:0] add_528027;
  wire [11:0] sel_528029;
  wire [11:0] add_528041;
  wire [11:0] sel_528043;
  wire [11:0] add_528045;
  wire [11:0] sel_528047;
  wire [8:0] add_528059;
  wire [11:0] sel_528061;
  wire [8:0] add_528063;
  wire [11:0] sel_528065;
  wire [11:0] add_528075;
  wire [11:0] sel_528077;
  wire [11:0] add_528079;
  wire [11:0] sel_528081;
  wire [11:0] add_528093;
  wire [11:0] sel_528095;
  wire [11:0] add_528097;
  wire [11:0] sel_528099;
  wire [10:0] add_528111;
  wire [11:0] sel_528113;
  wire [10:0] add_528115;
  wire [11:0] sel_528117;
  wire [11:0] add_528127;
  wire [11:0] sel_528129;
  wire [11:0] add_528131;
  wire [11:0] sel_528133;
  wire [11:0] add_528143;
  wire [11:0] sel_528145;
  wire [11:0] add_528147;
  wire [11:0] sel_528149;
  wire [11:0] add_528159;
  wire [11:0] sel_528161;
  wire [11:0] add_528163;
  wire [11:0] sel_528165;
  wire [8:0] add_528201;
  wire [11:0] add_528203;
  wire [11:0] sel_528205;
  wire [11:0] add_528207;
  wire [11:0] sel_528209;
  wire [11:0] add_528221;
  wire [11:0] sel_528223;
  wire [11:0] add_528225;
  wire [11:0] sel_528227;
  wire [10:0] add_528239;
  wire [11:0] sel_528241;
  wire [10:0] add_528243;
  wire [11:0] sel_528245;
  wire [10:0] add_528255;
  wire [11:0] sel_528257;
  wire [10:0] add_528259;
  wire [11:0] sel_528261;
  wire [9:0] add_528273;
  wire [11:0] sel_528275;
  wire [9:0] add_528277;
  wire [11:0] sel_528279;
  wire [11:0] add_528291;
  wire [11:0] sel_528293;
  wire [11:0] add_528295;
  wire [11:0] sel_528297;
  wire [10:0] add_528309;
  wire [11:0] sel_528311;
  wire [10:0] add_528313;
  wire [11:0] sel_528315;
  wire [10:0] add_528325;
  wire [11:0] sel_528327;
  wire [10:0] add_528329;
  wire [11:0] sel_528331;
  wire [11:0] add_528341;
  wire [11:0] sel_528343;
  wire [11:0] add_528345;
  wire [11:0] sel_528347;
  wire [11:0] add_528357;
  wire [11:0] sel_528359;
  wire [11:0] add_528361;
  wire [11:0] sel_528363;
  wire [11:0] add_528373;
  wire [11:0] sel_528375;
  wire [11:0] add_528377;
  wire [11:0] sel_528379;
  wire [8:0] add_528391;
  wire [11:0] sel_528393;
  wire [8:0] add_528395;
  wire [11:0] sel_528397;
  wire [9:0] add_528441;
  wire [11:0] sel_528443;
  wire [9:0] add_528445;
  wire [11:0] sel_528447;
  wire [7:0] add_528459;
  wire [11:0] sel_528461;
  wire [7:0] add_528463;
  wire [11:0] sel_528465;
  wire [11:0] add_528475;
  wire [11:0] sel_528477;
  wire [11:0] add_528479;
  wire [11:0] sel_528481;
  wire [10:0] add_528491;
  wire [11:0] sel_528493;
  wire [10:0] add_528495;
  wire [11:0] sel_528497;
  wire [8:0] add_528507;
  wire [11:0] sel_528509;
  wire [8:0] add_528511;
  wire [11:0] sel_528513;
  wire [8:0] add_528525;
  wire [11:0] sel_528527;
  wire [8:0] add_528529;
  wire [11:0] sel_528531;
  wire [11:0] add_528541;
  wire [11:0] sel_528543;
  wire [11:0] add_528545;
  wire [11:0] sel_528547;
  wire [11:0] add_528557;
  wire [11:0] sel_528559;
  wire [11:0] add_528561;
  wire [11:0] sel_528563;
  wire [11:0] add_528575;
  wire [11:0] sel_528577;
  wire [11:0] add_528579;
  wire [11:0] sel_528581;
  wire [11:0] add_528591;
  wire [11:0] sel_528593;
  wire [11:0] add_528595;
  wire [11:0] sel_528597;
  wire [10:0] add_528607;
  wire [11:0] sel_528609;
  wire [10:0] add_528611;
  wire [11:0] sel_528613;
  wire [11:0] add_528623;
  wire [11:0] sel_528625;
  wire [11:0] add_528627;
  wire [11:0] sel_528629;
  wire [8:0] add_528631;
  wire [11:0] sel_528634;
  wire [8:0] add_528636;
  wire [11:0] sel_528639;
  wire [10:0] add_528641;
  wire [11:0] sel_528643;
  wire [10:0] add_528645;
  wire [11:0] sel_528647;
  wire [9:0] add_528649;
  wire [11:0] sel_528651;
  wire [9:0] add_528653;
  wire [11:0] sel_528655;
  wire [11:0] add_528657;
  wire [11:0] sel_528659;
  wire [11:0] add_528661;
  wire [11:0] sel_528663;
  wire [10:0] add_528665;
  wire [11:0] sel_528667;
  wire [10:0] add_528669;
  wire [11:0] sel_528671;
  wire [9:0] concat_528674;
  wire [10:0] add_528685;
  wire [11:0] sel_528687;
  wire [10:0] add_528689;
  wire [11:0] sel_528691;
  wire [11:0] add_528701;
  wire [11:0] sel_528703;
  wire [11:0] add_528705;
  wire [11:0] sel_528707;
  wire [11:0] add_528719;
  wire [11:0] sel_528721;
  wire [11:0] add_528723;
  wire [11:0] sel_528725;
  wire [11:0] add_528737;
  wire [11:0] sel_528739;
  wire [11:0] add_528741;
  wire [11:0] sel_528743;
  wire [8:0] add_528755;
  wire [11:0] sel_528757;
  wire [8:0] add_528759;
  wire [11:0] sel_528761;
  wire [11:0] add_528771;
  wire [11:0] sel_528773;
  wire [11:0] add_528775;
  wire [11:0] sel_528777;
  wire [11:0] add_528789;
  wire [11:0] sel_528791;
  wire [11:0] add_528793;
  wire [11:0] sel_528795;
  wire [10:0] add_528807;
  wire [11:0] sel_528809;
  wire [10:0] add_528811;
  wire [11:0] sel_528813;
  wire [11:0] add_528823;
  wire [11:0] sel_528825;
  wire [11:0] add_528827;
  wire [11:0] sel_528829;
  wire [11:0] add_528839;
  wire [11:0] sel_528841;
  wire [11:0] add_528843;
  wire [11:0] sel_528845;
  wire [11:0] add_528855;
  wire [11:0] sel_528857;
  wire [11:0] add_528859;
  wire [11:0] sel_528861;
  wire [9:0] add_528893;
  wire [11:0] add_528895;
  wire [11:0] sel_528897;
  wire [11:0] add_528899;
  wire [11:0] sel_528901;
  wire [11:0] add_528913;
  wire [11:0] sel_528915;
  wire [11:0] add_528917;
  wire [11:0] sel_528919;
  wire [10:0] add_528931;
  wire [11:0] sel_528933;
  wire [10:0] add_528935;
  wire [11:0] sel_528937;
  wire [10:0] add_528947;
  wire [11:0] sel_528949;
  wire [10:0] add_528951;
  wire [11:0] sel_528953;
  wire [9:0] add_528965;
  wire [11:0] sel_528967;
  wire [9:0] add_528969;
  wire [11:0] sel_528971;
  wire [11:0] add_528983;
  wire [11:0] sel_528985;
  wire [11:0] add_528987;
  wire [11:0] sel_528989;
  wire [10:0] add_529001;
  wire [11:0] sel_529003;
  wire [10:0] add_529005;
  wire [11:0] sel_529007;
  wire [10:0] add_529017;
  wire [11:0] sel_529019;
  wire [10:0] add_529021;
  wire [11:0] sel_529023;
  wire [11:0] add_529033;
  wire [11:0] sel_529035;
  wire [11:0] add_529037;
  wire [11:0] sel_529039;
  wire [11:0] add_529049;
  wire [11:0] sel_529051;
  wire [11:0] add_529053;
  wire [11:0] sel_529055;
  wire [11:0] add_529065;
  wire [11:0] sel_529067;
  wire [11:0] add_529069;
  wire [11:0] sel_529071;
  wire [8:0] add_529083;
  wire [11:0] sel_529085;
  wire [8:0] add_529087;
  wire [11:0] sel_529089;
  wire [9:0] add_529129;
  wire [11:0] sel_529131;
  wire [9:0] add_529133;
  wire [11:0] sel_529135;
  wire [7:0] add_529147;
  wire [11:0] sel_529149;
  wire [7:0] add_529151;
  wire [11:0] sel_529153;
  wire [11:0] add_529163;
  wire [11:0] sel_529165;
  wire [11:0] add_529167;
  wire [11:0] sel_529169;
  wire [10:0] add_529179;
  wire [11:0] sel_529181;
  wire [10:0] add_529183;
  wire [11:0] sel_529185;
  wire [8:0] add_529195;
  wire [11:0] sel_529197;
  wire [8:0] add_529199;
  wire [11:0] sel_529201;
  wire [8:0] add_529213;
  wire [11:0] sel_529215;
  wire [8:0] add_529217;
  wire [11:0] sel_529219;
  wire [11:0] add_529229;
  wire [11:0] sel_529231;
  wire [11:0] add_529233;
  wire [11:0] sel_529235;
  wire [11:0] add_529245;
  wire [11:0] sel_529247;
  wire [11:0] add_529249;
  wire [11:0] sel_529251;
  wire [11:0] add_529263;
  wire [11:0] sel_529265;
  wire [11:0] add_529267;
  wire [11:0] sel_529269;
  wire [11:0] add_529279;
  wire [11:0] sel_529281;
  wire [11:0] add_529283;
  wire [11:0] sel_529285;
  wire [10:0] add_529295;
  wire [11:0] sel_529297;
  wire [10:0] add_529299;
  wire [11:0] sel_529301;
  wire [11:0] add_529311;
  wire [11:0] sel_529313;
  wire [11:0] add_529315;
  wire [11:0] sel_529317;
  wire [8:0] add_529319;
  wire [11:0] sel_529322;
  wire [8:0] add_529324;
  wire [11:0] sel_529327;
  wire [10:0] add_529329;
  wire [11:0] sel_529331;
  wire [10:0] add_529333;
  wire [11:0] sel_529335;
  wire [9:0] add_529337;
  wire [11:0] sel_529339;
  wire [9:0] add_529341;
  wire [11:0] sel_529343;
  wire [11:0] add_529345;
  wire [11:0] sel_529347;
  wire [11:0] add_529349;
  wire [11:0] sel_529351;
  wire [10:0] concat_529354;
  wire [10:0] add_529365;
  wire [11:0] sel_529367;
  wire [10:0] add_529369;
  wire [11:0] sel_529371;
  wire [11:0] add_529381;
  wire [11:0] sel_529383;
  wire [11:0] add_529385;
  wire [11:0] sel_529387;
  wire [11:0] add_529399;
  wire [11:0] sel_529401;
  wire [11:0] add_529403;
  wire [11:0] sel_529405;
  wire [11:0] add_529417;
  wire [11:0] sel_529419;
  wire [11:0] add_529421;
  wire [11:0] sel_529423;
  wire [8:0] add_529435;
  wire [11:0] sel_529437;
  wire [8:0] add_529439;
  wire [11:0] sel_529441;
  wire [11:0] add_529451;
  wire [11:0] sel_529453;
  wire [11:0] add_529455;
  wire [11:0] sel_529457;
  wire [11:0] add_529469;
  wire [11:0] sel_529471;
  wire [11:0] add_529473;
  wire [11:0] sel_529475;
  wire [10:0] add_529487;
  wire [11:0] sel_529489;
  wire [10:0] add_529491;
  wire [11:0] sel_529493;
  wire [11:0] add_529503;
  wire [11:0] sel_529505;
  wire [11:0] add_529507;
  wire [11:0] sel_529509;
  wire [11:0] add_529519;
  wire [11:0] sel_529521;
  wire [11:0] add_529523;
  wire [11:0] sel_529525;
  wire [11:0] add_529535;
  wire [11:0] sel_529537;
  wire [11:0] add_529539;
  wire [11:0] sel_529541;
  wire [10:0] add_529569;
  wire [11:0] add_529571;
  wire [11:0] sel_529573;
  wire [11:0] add_529575;
  wire [11:0] sel_529577;
  wire [11:0] add_529589;
  wire [11:0] sel_529591;
  wire [11:0] add_529593;
  wire [11:0] sel_529595;
  wire [10:0] add_529607;
  wire [11:0] sel_529609;
  wire [10:0] add_529611;
  wire [11:0] sel_529613;
  wire [10:0] add_529623;
  wire [11:0] sel_529625;
  wire [10:0] add_529627;
  wire [11:0] sel_529629;
  wire [9:0] add_529641;
  wire [11:0] sel_529643;
  wire [9:0] add_529645;
  wire [11:0] sel_529647;
  wire [11:0] add_529659;
  wire [11:0] sel_529661;
  wire [11:0] add_529663;
  wire [11:0] sel_529665;
  wire [10:0] add_529677;
  wire [11:0] sel_529679;
  wire [10:0] add_529681;
  wire [11:0] sel_529683;
  wire [10:0] add_529693;
  wire [11:0] sel_529695;
  wire [10:0] add_529697;
  wire [11:0] sel_529699;
  wire [11:0] add_529709;
  wire [11:0] sel_529711;
  wire [11:0] add_529713;
  wire [11:0] sel_529715;
  wire [11:0] add_529725;
  wire [11:0] sel_529727;
  wire [11:0] add_529729;
  wire [11:0] sel_529731;
  wire [11:0] add_529741;
  wire [11:0] sel_529743;
  wire [11:0] add_529745;
  wire [11:0] sel_529747;
  wire [8:0] add_529759;
  wire [11:0] sel_529761;
  wire [8:0] add_529763;
  wire [11:0] sel_529765;
  wire [9:0] add_529799;
  wire [11:0] sel_529801;
  wire [9:0] add_529803;
  wire [11:0] sel_529805;
  wire [7:0] add_529817;
  wire [11:0] sel_529819;
  wire [7:0] add_529821;
  wire [11:0] sel_529823;
  wire [11:0] add_529833;
  wire [11:0] sel_529835;
  wire [11:0] add_529837;
  wire [11:0] sel_529839;
  wire [10:0] add_529849;
  wire [11:0] sel_529851;
  wire [10:0] add_529853;
  wire [11:0] sel_529855;
  wire [8:0] add_529865;
  wire [11:0] sel_529867;
  wire [8:0] add_529869;
  wire [11:0] sel_529871;
  wire [8:0] add_529883;
  wire [11:0] sel_529885;
  wire [8:0] add_529887;
  wire [11:0] sel_529889;
  wire [11:0] add_529899;
  wire [11:0] sel_529901;
  wire [11:0] add_529903;
  wire [11:0] sel_529905;
  wire [11:0] add_529915;
  wire [11:0] sel_529917;
  wire [11:0] add_529919;
  wire [11:0] sel_529921;
  wire [11:0] add_529933;
  wire [11:0] sel_529935;
  wire [11:0] add_529937;
  wire [11:0] sel_529939;
  wire [11:0] add_529949;
  wire [11:0] sel_529951;
  wire [11:0] add_529953;
  wire [11:0] sel_529955;
  wire [10:0] add_529965;
  wire [11:0] sel_529967;
  wire [10:0] add_529969;
  wire [11:0] sel_529971;
  wire [11:0] add_529981;
  wire [11:0] sel_529983;
  wire [11:0] add_529985;
  wire [11:0] sel_529987;
  wire [8:0] add_529989;
  wire [11:0] sel_529992;
  wire [8:0] add_529994;
  wire [11:0] sel_529997;
  wire [10:0] add_529999;
  wire [11:0] sel_530001;
  wire [10:0] add_530003;
  wire [11:0] sel_530005;
  wire [9:0] add_530007;
  wire [11:0] sel_530009;
  wire [9:0] add_530011;
  wire [11:0] sel_530013;
  wire [11:0] concat_530016;
  wire [10:0] add_530027;
  wire [11:0] sel_530029;
  wire [10:0] add_530031;
  wire [11:0] sel_530033;
  wire [11:0] add_530043;
  wire [11:0] sel_530045;
  wire [11:0] add_530047;
  wire [11:0] sel_530049;
  wire [11:0] add_530061;
  wire [11:0] sel_530063;
  wire [11:0] add_530065;
  wire [11:0] sel_530067;
  wire [11:0] add_530079;
  wire [11:0] sel_530081;
  wire [11:0] add_530083;
  wire [11:0] sel_530085;
  wire [8:0] add_530097;
  wire [11:0] sel_530099;
  wire [8:0] add_530101;
  wire [11:0] sel_530103;
  wire [11:0] add_530113;
  wire [11:0] sel_530115;
  wire [11:0] add_530117;
  wire [11:0] sel_530119;
  wire [11:0] add_530131;
  wire [11:0] sel_530133;
  wire [11:0] add_530135;
  wire [11:0] sel_530137;
  wire [10:0] add_530149;
  wire [11:0] sel_530151;
  wire [10:0] add_530153;
  wire [11:0] sel_530155;
  wire [11:0] add_530165;
  wire [11:0] sel_530167;
  wire [11:0] add_530169;
  wire [11:0] sel_530171;
  wire [11:0] add_530181;
  wire [11:0] sel_530183;
  wire [11:0] add_530185;
  wire [11:0] sel_530187;
  wire [11:0] add_530197;
  wire [11:0] sel_530199;
  wire [11:0] add_530201;
  wire [11:0] sel_530203;
  wire [11:0] add_530227;
  wire [11:0] add_530229;
  wire [11:0] sel_530231;
  wire [11:0] add_530233;
  wire [11:0] sel_530235;
  wire [11:0] add_530247;
  wire [11:0] sel_530249;
  wire [11:0] add_530251;
  wire [11:0] sel_530253;
  wire [10:0] add_530265;
  wire [11:0] sel_530267;
  wire [10:0] add_530269;
  wire [11:0] sel_530271;
  wire [10:0] add_530281;
  wire [11:0] sel_530283;
  wire [10:0] add_530285;
  wire [11:0] sel_530287;
  wire [9:0] add_530299;
  wire [11:0] sel_530301;
  wire [9:0] add_530303;
  wire [11:0] sel_530305;
  wire [11:0] add_530317;
  wire [11:0] sel_530319;
  wire [11:0] add_530321;
  wire [11:0] sel_530323;
  wire [10:0] add_530335;
  wire [11:0] sel_530337;
  wire [10:0] add_530339;
  wire [11:0] sel_530341;
  wire [10:0] add_530351;
  wire [11:0] sel_530353;
  wire [10:0] add_530355;
  wire [11:0] sel_530357;
  wire [11:0] add_530367;
  wire [11:0] sel_530369;
  wire [11:0] add_530371;
  wire [11:0] sel_530373;
  wire [11:0] add_530383;
  wire [11:0] sel_530385;
  wire [11:0] add_530387;
  wire [11:0] sel_530389;
  wire [11:0] add_530399;
  wire [11:0] sel_530401;
  wire [11:0] add_530403;
  wire [11:0] sel_530405;
  wire [8:0] add_530417;
  wire [11:0] sel_530419;
  wire [8:0] add_530421;
  wire [11:0] sel_530423;
  wire [9:0] add_530453;
  wire [11:0] sel_530455;
  wire [9:0] add_530457;
  wire [11:0] sel_530459;
  wire [7:0] add_530471;
  wire [11:0] sel_530473;
  wire [7:0] add_530475;
  wire [11:0] sel_530477;
  wire [11:0] add_530487;
  wire [11:0] sel_530489;
  wire [11:0] add_530491;
  wire [11:0] sel_530493;
  wire [10:0] add_530503;
  wire [11:0] sel_530505;
  wire [10:0] add_530507;
  wire [11:0] sel_530509;
  wire [8:0] add_530519;
  wire [11:0] sel_530521;
  wire [8:0] add_530523;
  wire [11:0] sel_530525;
  wire [8:0] add_530537;
  wire [11:0] sel_530539;
  wire [8:0] add_530541;
  wire [11:0] sel_530543;
  wire [11:0] add_530553;
  wire [11:0] sel_530555;
  wire [11:0] add_530557;
  wire [11:0] sel_530559;
  wire [11:0] add_530569;
  wire [11:0] sel_530571;
  wire [11:0] add_530573;
  wire [11:0] sel_530575;
  wire [11:0] add_530587;
  wire [11:0] sel_530589;
  wire [11:0] add_530591;
  wire [11:0] sel_530593;
  wire [11:0] add_530603;
  wire [11:0] sel_530605;
  wire [11:0] add_530607;
  wire [11:0] sel_530609;
  wire [10:0] add_530619;
  wire [11:0] sel_530621;
  wire [10:0] add_530623;
  wire [11:0] sel_530625;
  wire [11:0] add_530635;
  wire [11:0] sel_530637;
  wire [11:0] add_530639;
  wire [11:0] sel_530641;
  wire [8:0] add_530643;
  wire [11:0] sel_530646;
  wire [8:0] add_530648;
  wire [11:0] sel_530651;
  wire [10:0] add_530653;
  wire [11:0] sel_530655;
  wire [10:0] add_530657;
  wire [11:0] sel_530659;
  wire [12:0] concat_530662;
  wire [10:0] add_530673;
  wire [11:0] sel_530675;
  wire [10:0] add_530677;
  wire [11:0] sel_530679;
  wire [11:0] add_530689;
  wire [11:0] sel_530691;
  wire [11:0] add_530693;
  wire [11:0] sel_530695;
  wire [11:0] add_530707;
  wire [11:0] sel_530709;
  wire [11:0] add_530711;
  wire [11:0] sel_530713;
  wire [11:0] add_530725;
  wire [11:0] sel_530727;
  wire [11:0] add_530729;
  wire [11:0] sel_530731;
  wire [8:0] add_530743;
  wire [11:0] sel_530745;
  wire [8:0] add_530747;
  wire [11:0] sel_530749;
  wire [11:0] add_530759;
  wire [11:0] sel_530761;
  wire [11:0] add_530763;
  wire [11:0] sel_530765;
  wire [11:0] add_530777;
  wire [11:0] sel_530779;
  wire [11:0] add_530781;
  wire [11:0] sel_530783;
  wire [10:0] add_530795;
  wire [11:0] sel_530797;
  wire [10:0] add_530799;
  wire [11:0] sel_530801;
  wire [11:0] add_530811;
  wire [11:0] sel_530813;
  wire [11:0] add_530815;
  wire [11:0] sel_530817;
  wire [11:0] add_530827;
  wire [11:0] sel_530829;
  wire [11:0] add_530831;
  wire [11:0] sel_530833;
  wire [11:0] add_530843;
  wire [11:0] sel_530845;
  wire [11:0] add_530847;
  wire [11:0] sel_530849;
  wire [12:0] add_530869;
  wire [11:0] add_530871;
  wire [11:0] sel_530873;
  wire [11:0] add_530875;
  wire [11:0] sel_530877;
  wire [11:0] add_530889;
  wire [11:0] sel_530891;
  wire [11:0] add_530893;
  wire [11:0] sel_530895;
  wire [10:0] add_530907;
  wire [11:0] sel_530909;
  wire [10:0] add_530911;
  wire [11:0] sel_530913;
  wire [10:0] add_530923;
  wire [11:0] sel_530925;
  wire [10:0] add_530927;
  wire [11:0] sel_530929;
  wire [9:0] add_530941;
  wire [11:0] sel_530943;
  wire [9:0] add_530945;
  wire [11:0] sel_530947;
  wire [11:0] add_530959;
  wire [11:0] sel_530961;
  wire [11:0] add_530963;
  wire [11:0] sel_530965;
  wire [10:0] add_530977;
  wire [11:0] sel_530979;
  wire [10:0] add_530981;
  wire [11:0] sel_530983;
  wire [10:0] add_530993;
  wire [11:0] sel_530995;
  wire [10:0] add_530997;
  wire [11:0] sel_530999;
  wire [11:0] add_531009;
  wire [11:0] sel_531011;
  wire [11:0] add_531013;
  wire [11:0] sel_531015;
  wire [11:0] add_531025;
  wire [11:0] sel_531027;
  wire [11:0] add_531029;
  wire [11:0] sel_531031;
  wire [11:0] add_531041;
  wire [11:0] sel_531043;
  wire [11:0] add_531045;
  wire [11:0] sel_531047;
  wire [8:0] add_531059;
  wire [11:0] sel_531061;
  wire [8:0] add_531063;
  wire [11:0] sel_531065;
  wire [9:0] add_531089;
  wire [11:0] sel_531091;
  wire [9:0] add_531093;
  wire [11:0] sel_531095;
  wire [7:0] add_531107;
  wire [11:0] sel_531109;
  wire [7:0] add_531111;
  wire [11:0] sel_531113;
  wire [11:0] add_531123;
  wire [11:0] sel_531125;
  wire [11:0] add_531127;
  wire [11:0] sel_531129;
  wire [10:0] add_531139;
  wire [11:0] sel_531141;
  wire [10:0] add_531143;
  wire [11:0] sel_531145;
  wire [8:0] add_531155;
  wire [11:0] sel_531157;
  wire [8:0] add_531159;
  wire [11:0] sel_531161;
  wire [8:0] add_531173;
  wire [11:0] sel_531175;
  wire [8:0] add_531177;
  wire [11:0] sel_531179;
  wire [11:0] add_531189;
  wire [11:0] sel_531191;
  wire [11:0] add_531193;
  wire [11:0] sel_531195;
  wire [11:0] add_531205;
  wire [11:0] sel_531207;
  wire [11:0] add_531209;
  wire [11:0] sel_531211;
  wire [11:0] add_531223;
  wire [11:0] sel_531225;
  wire [11:0] add_531227;
  wire [11:0] sel_531229;
  wire [11:0] add_531239;
  wire [11:0] sel_531241;
  wire [11:0] add_531243;
  wire [11:0] sel_531245;
  wire [10:0] add_531255;
  wire [11:0] sel_531257;
  wire [10:0] add_531259;
  wire [11:0] sel_531261;
  wire [11:0] add_531271;
  wire [11:0] sel_531273;
  wire [11:0] add_531275;
  wire [11:0] sel_531277;
  wire [8:0] add_531279;
  wire [11:0] sel_531282;
  wire [8:0] add_531284;
  wire [11:0] sel_531287;
  wire [13:0] concat_531290;
  wire [10:0] add_531301;
  wire [11:0] sel_531303;
  wire [10:0] add_531305;
  wire [11:0] sel_531307;
  wire [11:0] add_531317;
  wire [11:0] sel_531319;
  wire [11:0] add_531321;
  wire [11:0] sel_531323;
  wire [11:0] add_531335;
  wire [11:0] sel_531337;
  wire [11:0] add_531339;
  wire [11:0] sel_531341;
  wire [11:0] add_531353;
  wire [11:0] sel_531355;
  wire [11:0] add_531357;
  wire [11:0] sel_531359;
  wire [8:0] add_531371;
  wire [11:0] sel_531373;
  wire [8:0] add_531375;
  wire [11:0] sel_531377;
  wire [11:0] add_531387;
  wire [11:0] sel_531389;
  wire [11:0] add_531391;
  wire [11:0] sel_531393;
  wire [11:0] add_531405;
  wire [11:0] sel_531407;
  wire [11:0] add_531409;
  wire [11:0] sel_531411;
  wire [10:0] add_531423;
  wire [11:0] sel_531425;
  wire [10:0] add_531427;
  wire [11:0] sel_531429;
  wire [11:0] add_531439;
  wire [11:0] sel_531441;
  wire [11:0] add_531443;
  wire [11:0] sel_531445;
  wire [11:0] add_531455;
  wire [11:0] sel_531457;
  wire [11:0] add_531459;
  wire [11:0] sel_531461;
  wire [11:0] add_531471;
  wire [11:0] sel_531473;
  wire [11:0] add_531475;
  wire [11:0] sel_531477;
  wire [13:0] add_531493;
  wire [11:0] add_531495;
  wire [11:0] sel_531497;
  wire [11:0] add_531499;
  wire [11:0] sel_531501;
  wire [11:0] add_531513;
  wire [11:0] sel_531515;
  wire [11:0] add_531517;
  wire [11:0] sel_531519;
  wire [10:0] add_531531;
  wire [11:0] sel_531533;
  wire [10:0] add_531535;
  wire [11:0] sel_531537;
  wire [10:0] add_531547;
  wire [11:0] sel_531549;
  wire [10:0] add_531551;
  wire [11:0] sel_531553;
  wire [9:0] add_531565;
  wire [11:0] sel_531567;
  wire [9:0] add_531569;
  wire [11:0] sel_531571;
  wire [11:0] add_531583;
  wire [11:0] sel_531585;
  wire [11:0] add_531587;
  wire [11:0] sel_531589;
  wire [10:0] add_531601;
  wire [11:0] sel_531603;
  wire [10:0] add_531605;
  wire [11:0] sel_531607;
  wire [10:0] add_531617;
  wire [11:0] sel_531619;
  wire [10:0] add_531621;
  wire [11:0] sel_531623;
  wire [11:0] add_531633;
  wire [11:0] sel_531635;
  wire [11:0] add_531637;
  wire [11:0] sel_531639;
  wire [11:0] add_531649;
  wire [11:0] sel_531651;
  wire [11:0] add_531653;
  wire [11:0] sel_531655;
  wire [11:0] add_531665;
  wire [11:0] sel_531667;
  wire [11:0] add_531669;
  wire [11:0] sel_531671;
  wire [8:0] add_531683;
  wire [11:0] sel_531685;
  wire [8:0] add_531687;
  wire [11:0] sel_531689;
  wire [9:0] add_531705;
  wire [11:0] sel_531707;
  wire [9:0] add_531709;
  wire [11:0] sel_531711;
  wire [7:0] add_531723;
  wire [11:0] sel_531725;
  wire [7:0] add_531727;
  wire [11:0] sel_531729;
  wire [11:0] add_531739;
  wire [11:0] sel_531741;
  wire [11:0] add_531743;
  wire [11:0] sel_531745;
  wire [10:0] add_531755;
  wire [11:0] sel_531757;
  wire [10:0] add_531759;
  wire [11:0] sel_531761;
  wire [8:0] add_531771;
  wire [11:0] sel_531773;
  wire [8:0] add_531775;
  wire [11:0] sel_531777;
  wire [8:0] add_531789;
  wire [11:0] sel_531791;
  wire [8:0] add_531793;
  wire [11:0] sel_531795;
  wire [11:0] add_531805;
  wire [11:0] sel_531807;
  wire [11:0] add_531809;
  wire [11:0] sel_531811;
  wire [11:0] add_531821;
  wire [11:0] sel_531823;
  wire [11:0] add_531825;
  wire [11:0] sel_531827;
  wire [11:0] add_531839;
  wire [11:0] sel_531841;
  wire [11:0] add_531843;
  wire [11:0] sel_531845;
  wire [11:0] add_531855;
  wire [11:0] sel_531857;
  wire [11:0] add_531859;
  wire [11:0] sel_531861;
  wire [10:0] add_531871;
  wire [11:0] sel_531873;
  wire [10:0] add_531875;
  wire [11:0] sel_531877;
  wire [11:0] add_531887;
  wire [11:0] sel_531889;
  wire [11:0] add_531891;
  wire [11:0] sel_531893;
  wire [14:0] concat_531896;
  wire [10:0] add_531907;
  wire [11:0] sel_531909;
  wire [10:0] add_531911;
  wire [11:0] sel_531913;
  wire [11:0] add_531923;
  wire [11:0] sel_531925;
  wire [11:0] add_531927;
  wire [11:0] sel_531929;
  wire [11:0] add_531941;
  wire [11:0] sel_531943;
  wire [11:0] add_531945;
  wire [11:0] sel_531947;
  wire [11:0] add_531959;
  wire [11:0] sel_531961;
  wire [11:0] add_531963;
  wire [11:0] sel_531965;
  wire [8:0] add_531977;
  wire [11:0] sel_531979;
  wire [8:0] add_531981;
  wire [11:0] sel_531983;
  wire [11:0] add_531993;
  wire [11:0] sel_531995;
  wire [11:0] add_531997;
  wire [11:0] sel_531999;
  wire [11:0] add_532011;
  wire [11:0] sel_532013;
  wire [11:0] add_532015;
  wire [11:0] sel_532017;
  wire [10:0] add_532029;
  wire [11:0] sel_532031;
  wire [10:0] add_532033;
  wire [11:0] sel_532035;
  wire [11:0] add_532045;
  wire [11:0] sel_532047;
  wire [11:0] add_532049;
  wire [11:0] sel_532051;
  wire [11:0] add_532061;
  wire [11:0] sel_532063;
  wire [11:0] add_532065;
  wire [11:0] sel_532067;
  wire [11:0] add_532077;
  wire [11:0] sel_532079;
  wire [11:0] add_532081;
  wire [11:0] sel_532083;
  wire [14:0] add_532095;
  wire [11:0] add_532097;
  wire [11:0] sel_532099;
  wire [11:0] add_532101;
  wire [11:0] sel_532103;
  wire [11:0] add_532115;
  wire [11:0] sel_532117;
  wire [11:0] add_532119;
  wire [11:0] sel_532121;
  wire [10:0] add_532133;
  wire [11:0] sel_532135;
  wire [10:0] add_532137;
  wire [11:0] sel_532139;
  wire [10:0] add_532149;
  wire [11:0] sel_532151;
  wire [10:0] add_532153;
  wire [11:0] sel_532155;
  wire [9:0] add_532167;
  wire [11:0] sel_532169;
  wire [9:0] add_532171;
  wire [11:0] sel_532173;
  wire [11:0] add_532185;
  wire [11:0] sel_532187;
  wire [11:0] add_532189;
  wire [11:0] sel_532191;
  wire [10:0] add_532203;
  wire [11:0] sel_532205;
  wire [10:0] add_532207;
  wire [11:0] sel_532209;
  wire [10:0] add_532219;
  wire [11:0] sel_532221;
  wire [10:0] add_532223;
  wire [11:0] sel_532225;
  wire [11:0] add_532235;
  wire [11:0] sel_532237;
  wire [11:0] add_532239;
  wire [11:0] sel_532241;
  wire [11:0] add_532251;
  wire [11:0] sel_532253;
  wire [11:0] add_532255;
  wire [11:0] sel_532257;
  wire [11:0] add_532267;
  wire [11:0] sel_532269;
  wire [11:0] add_532271;
  wire [11:0] sel_532273;
  wire [8:0] add_532285;
  wire [11:0] sel_532287;
  wire [8:0] add_532289;
  wire [11:0] sel_532291;
  wire [9:0] add_532301;
  wire [11:0] sel_532303;
  wire [9:0] add_532305;
  wire [11:0] sel_532307;
  wire [7:0] add_532319;
  wire [11:0] sel_532321;
  wire [7:0] add_532323;
  wire [11:0] sel_532325;
  wire [11:0] add_532335;
  wire [11:0] sel_532337;
  wire [11:0] add_532339;
  wire [11:0] sel_532341;
  wire [10:0] add_532351;
  wire [11:0] sel_532353;
  wire [10:0] add_532355;
  wire [11:0] sel_532357;
  wire [8:0] add_532367;
  wire [11:0] sel_532369;
  wire [8:0] add_532371;
  wire [11:0] sel_532373;
  wire [8:0] add_532385;
  wire [11:0] sel_532387;
  wire [8:0] add_532389;
  wire [11:0] sel_532391;
  wire [11:0] add_532401;
  wire [11:0] sel_532403;
  wire [11:0] add_532405;
  wire [11:0] sel_532407;
  wire [11:0] add_532417;
  wire [11:0] sel_532419;
  wire [11:0] add_532421;
  wire [11:0] sel_532423;
  wire [11:0] add_532435;
  wire [11:0] sel_532437;
  wire [11:0] add_532439;
  wire [11:0] sel_532441;
  wire [11:0] add_532451;
  wire [11:0] sel_532453;
  wire [11:0] add_532455;
  wire [11:0] sel_532457;
  wire [10:0] add_532467;
  wire [11:0] sel_532469;
  wire [10:0] add_532471;
  wire [11:0] sel_532473;
  wire [15:0] concat_532484;
  wire [10:0] add_532495;
  wire [11:0] sel_532497;
  wire [10:0] add_532499;
  wire [11:0] sel_532501;
  wire [11:0] add_532511;
  wire [11:0] sel_532513;
  wire [11:0] add_532515;
  wire [11:0] sel_532517;
  wire [11:0] add_532529;
  wire [11:0] sel_532531;
  wire [11:0] add_532533;
  wire [11:0] sel_532535;
  wire [11:0] add_532547;
  wire [11:0] sel_532549;
  wire [11:0] add_532551;
  wire [11:0] sel_532553;
  wire [8:0] add_532565;
  wire [11:0] sel_532567;
  wire [8:0] add_532569;
  wire [11:0] sel_532571;
  wire [11:0] add_532581;
  wire [11:0] sel_532583;
  wire [11:0] add_532585;
  wire [11:0] sel_532587;
  wire [11:0] add_532599;
  wire [11:0] sel_532601;
  wire [11:0] add_532603;
  wire [11:0] sel_532605;
  wire [10:0] add_532617;
  wire [11:0] sel_532619;
  wire [10:0] add_532621;
  wire [11:0] sel_532623;
  wire [11:0] add_532633;
  wire [11:0] sel_532635;
  wire [11:0] add_532637;
  wire [11:0] sel_532639;
  wire [11:0] add_532649;
  wire [11:0] sel_532651;
  wire [11:0] add_532653;
  wire [11:0] sel_532655;
  wire [11:0] add_532665;
  wire [11:0] sel_532667;
  wire [11:0] add_532669;
  wire [11:0] sel_532671;
  wire [15:0] add_532677;
  wire [11:0] add_532679;
  wire [11:0] sel_532681;
  wire [11:0] add_532683;
  wire [11:0] sel_532685;
  wire [11:0] add_532697;
  wire [11:0] sel_532699;
  wire [11:0] add_532701;
  wire [11:0] sel_532703;
  wire [10:0] add_532715;
  wire [11:0] sel_532717;
  wire [10:0] add_532719;
  wire [11:0] sel_532721;
  wire [10:0] add_532731;
  wire [11:0] sel_532733;
  wire [10:0] add_532735;
  wire [11:0] sel_532737;
  wire [9:0] add_532749;
  wire [11:0] sel_532751;
  wire [9:0] add_532753;
  wire [11:0] sel_532755;
  wire [11:0] add_532767;
  wire [11:0] sel_532769;
  wire [11:0] add_532771;
  wire [11:0] sel_532773;
  wire [10:0] add_532785;
  wire [11:0] sel_532787;
  wire [10:0] add_532789;
  wire [11:0] sel_532791;
  wire [10:0] add_532801;
  wire [11:0] sel_532803;
  wire [10:0] add_532805;
  wire [11:0] sel_532807;
  wire [11:0] add_532817;
  wire [11:0] sel_532819;
  wire [11:0] add_532821;
  wire [11:0] sel_532823;
  wire [11:0] add_532833;
  wire [11:0] sel_532835;
  wire [11:0] add_532837;
  wire [11:0] sel_532839;
  wire [11:0] add_532849;
  wire [11:0] sel_532851;
  wire [11:0] add_532853;
  wire [11:0] sel_532855;
  wire [15:0] sel_532868;
  wire [9:0] add_532875;
  wire [11:0] sel_532877;
  wire [9:0] add_532879;
  wire [11:0] sel_532881;
  wire [7:0] add_532893;
  wire [11:0] sel_532895;
  wire [7:0] add_532897;
  wire [11:0] sel_532899;
  wire [11:0] add_532909;
  wire [11:0] sel_532911;
  wire [11:0] add_532913;
  wire [11:0] sel_532915;
  wire [10:0] add_532925;
  wire [11:0] sel_532927;
  wire [10:0] add_532929;
  wire [11:0] sel_532931;
  wire [8:0] add_532941;
  wire [11:0] sel_532943;
  wire [8:0] add_532945;
  wire [11:0] sel_532947;
  wire [8:0] add_532959;
  wire [11:0] sel_532961;
  wire [8:0] add_532963;
  wire [11:0] sel_532965;
  wire [11:0] add_532975;
  wire [11:0] sel_532977;
  wire [11:0] add_532979;
  wire [11:0] sel_532981;
  wire [11:0] add_532991;
  wire [11:0] sel_532993;
  wire [11:0] add_532995;
  wire [11:0] sel_532997;
  wire [11:0] add_533009;
  wire [11:0] sel_533011;
  wire [11:0] add_533013;
  wire [11:0] sel_533015;
  wire [11:0] add_533025;
  wire [11:0] sel_533027;
  wire [11:0] add_533029;
  wire [11:0] sel_533031;
  wire [10:0] add_533041;
  wire [11:0] sel_533043;
  wire [10:0] add_533045;
  wire [11:0] sel_533047;
  wire [15:0] add_533051;
  wire [10:0] add_533061;
  wire [11:0] sel_533063;
  wire [10:0] add_533065;
  wire [11:0] sel_533067;
  wire [11:0] add_533077;
  wire [11:0] sel_533079;
  wire [11:0] add_533081;
  wire [11:0] sel_533083;
  wire [11:0] add_533095;
  wire [11:0] sel_533097;
  wire [11:0] add_533099;
  wire [11:0] sel_533101;
  wire [11:0] add_533113;
  wire [11:0] sel_533115;
  wire [11:0] add_533117;
  wire [11:0] sel_533119;
  wire [8:0] add_533131;
  wire [11:0] sel_533133;
  wire [8:0] add_533135;
  wire [11:0] sel_533137;
  wire [11:0] add_533147;
  wire [11:0] sel_533149;
  wire [11:0] add_533151;
  wire [11:0] sel_533153;
  wire [11:0] add_533165;
  wire [11:0] sel_533167;
  wire [11:0] add_533169;
  wire [11:0] sel_533171;
  wire [10:0] add_533183;
  wire [11:0] sel_533185;
  wire [10:0] add_533187;
  wire [11:0] sel_533189;
  wire [11:0] add_533199;
  wire [11:0] sel_533201;
  wire [11:0] add_533203;
  wire [11:0] sel_533205;
  wire [11:0] add_533215;
  wire [11:0] sel_533217;
  wire [11:0] add_533219;
  wire [11:0] sel_533221;
  wire [15:0] sel_533232;
  wire [11:0] add_533235;
  wire [11:0] sel_533237;
  wire [11:0] add_533239;
  wire [11:0] sel_533241;
  wire [11:0] add_533253;
  wire [11:0] sel_533255;
  wire [11:0] add_533257;
  wire [11:0] sel_533259;
  wire [10:0] add_533271;
  wire [11:0] sel_533273;
  wire [10:0] add_533275;
  wire [11:0] sel_533277;
  wire [10:0] add_533287;
  wire [11:0] sel_533289;
  wire [10:0] add_533291;
  wire [11:0] sel_533293;
  wire [9:0] add_533305;
  wire [11:0] sel_533307;
  wire [9:0] add_533309;
  wire [11:0] sel_533311;
  wire [11:0] add_533323;
  wire [11:0] sel_533325;
  wire [11:0] add_533327;
  wire [11:0] sel_533329;
  wire [10:0] add_533341;
  wire [11:0] sel_533343;
  wire [10:0] add_533345;
  wire [11:0] sel_533347;
  wire [10:0] add_533357;
  wire [11:0] sel_533359;
  wire [10:0] add_533361;
  wire [11:0] sel_533363;
  wire [11:0] add_533373;
  wire [11:0] sel_533375;
  wire [11:0] add_533377;
  wire [11:0] sel_533379;
  wire [11:0] add_533389;
  wire [11:0] sel_533391;
  wire [11:0] add_533393;
  wire [11:0] sel_533395;
  wire [11:0] add_533405;
  wire [11:0] sel_533407;
  wire [11:0] add_533409;
  wire [11:0] sel_533411;
  wire [15:0] add_533417;
  wire [9:0] add_533423;
  wire [11:0] sel_533425;
  wire [9:0] add_533427;
  wire [11:0] sel_533429;
  wire [7:0] add_533441;
  wire [11:0] sel_533443;
  wire [7:0] add_533445;
  wire [11:0] sel_533447;
  wire [11:0] add_533457;
  wire [11:0] sel_533459;
  wire [11:0] add_533461;
  wire [11:0] sel_533463;
  wire [10:0] add_533473;
  wire [11:0] sel_533475;
  wire [10:0] add_533477;
  wire [11:0] sel_533479;
  wire [8:0] add_533489;
  wire [11:0] sel_533491;
  wire [8:0] add_533493;
  wire [11:0] sel_533495;
  wire [8:0] add_533507;
  wire [11:0] sel_533509;
  wire [8:0] add_533511;
  wire [11:0] sel_533513;
  wire [11:0] add_533523;
  wire [11:0] sel_533525;
  wire [11:0] add_533527;
  wire [11:0] sel_533529;
  wire [11:0] add_533539;
  wire [11:0] sel_533541;
  wire [11:0] add_533543;
  wire [11:0] sel_533545;
  wire [11:0] add_533557;
  wire [11:0] sel_533559;
  wire [11:0] add_533561;
  wire [11:0] sel_533563;
  wire [11:0] add_533573;
  wire [11:0] sel_533575;
  wire [11:0] add_533577;
  wire [11:0] sel_533579;
  wire [15:0] sel_533590;
  wire [10:0] add_533601;
  wire [11:0] sel_533603;
  wire [10:0] add_533605;
  wire [11:0] sel_533607;
  wire [11:0] add_533617;
  wire [11:0] sel_533619;
  wire [11:0] add_533621;
  wire [11:0] sel_533623;
  wire [11:0] add_533635;
  wire [11:0] sel_533637;
  wire [11:0] add_533639;
  wire [11:0] sel_533641;
  wire [11:0] add_533653;
  wire [11:0] sel_533655;
  wire [11:0] add_533657;
  wire [11:0] sel_533659;
  wire [8:0] add_533671;
  wire [11:0] sel_533673;
  wire [8:0] add_533675;
  wire [11:0] sel_533677;
  wire [11:0] add_533687;
  wire [11:0] sel_533689;
  wire [11:0] add_533691;
  wire [11:0] sel_533693;
  wire [11:0] add_533705;
  wire [11:0] sel_533707;
  wire [11:0] add_533709;
  wire [11:0] sel_533711;
  wire [10:0] add_533723;
  wire [11:0] sel_533725;
  wire [10:0] add_533727;
  wire [11:0] sel_533729;
  wire [11:0] add_533739;
  wire [11:0] sel_533741;
  wire [11:0] add_533743;
  wire [11:0] sel_533745;
  wire [11:0] add_533755;
  wire [11:0] sel_533757;
  wire [11:0] add_533759;
  wire [11:0] sel_533761;
  wire [15:0] add_533765;
  wire [11:0] add_533767;
  wire [11:0] sel_533769;
  wire [11:0] add_533771;
  wire [11:0] sel_533773;
  wire [11:0] add_533785;
  wire [11:0] sel_533787;
  wire [11:0] add_533789;
  wire [11:0] sel_533791;
  wire [10:0] add_533803;
  wire [11:0] sel_533805;
  wire [10:0] add_533807;
  wire [11:0] sel_533809;
  wire [10:0] add_533819;
  wire [11:0] sel_533821;
  wire [10:0] add_533823;
  wire [11:0] sel_533825;
  wire [9:0] add_533837;
  wire [11:0] sel_533839;
  wire [9:0] add_533841;
  wire [11:0] sel_533843;
  wire [11:0] add_533855;
  wire [11:0] sel_533857;
  wire [11:0] add_533859;
  wire [11:0] sel_533861;
  wire [10:0] add_533873;
  wire [11:0] sel_533875;
  wire [10:0] add_533877;
  wire [11:0] sel_533879;
  wire [10:0] add_533889;
  wire [11:0] sel_533891;
  wire [10:0] add_533893;
  wire [11:0] sel_533895;
  wire [11:0] add_533905;
  wire [11:0] sel_533907;
  wire [11:0] add_533909;
  wire [11:0] sel_533911;
  wire [11:0] add_533921;
  wire [11:0] sel_533923;
  wire [11:0] add_533925;
  wire [11:0] sel_533927;
  wire [15:0] sel_533938;
  wire [9:0] add_533945;
  wire [11:0] sel_533947;
  wire [9:0] add_533949;
  wire [11:0] sel_533951;
  wire [7:0] add_533963;
  wire [11:0] sel_533965;
  wire [7:0] add_533967;
  wire [11:0] sel_533969;
  wire [11:0] add_533979;
  wire [11:0] sel_533981;
  wire [11:0] add_533983;
  wire [11:0] sel_533985;
  wire [10:0] add_533995;
  wire [11:0] sel_533997;
  wire [10:0] add_533999;
  wire [11:0] sel_534001;
  wire [8:0] add_534011;
  wire [11:0] sel_534013;
  wire [8:0] add_534015;
  wire [11:0] sel_534017;
  wire [8:0] add_534029;
  wire [11:0] sel_534031;
  wire [8:0] add_534033;
  wire [11:0] sel_534035;
  wire [11:0] add_534045;
  wire [11:0] sel_534047;
  wire [11:0] add_534049;
  wire [11:0] sel_534051;
  wire [11:0] add_534061;
  wire [11:0] sel_534063;
  wire [11:0] add_534065;
  wire [11:0] sel_534067;
  wire [11:0] add_534079;
  wire [11:0] sel_534081;
  wire [11:0] add_534083;
  wire [11:0] sel_534085;
  wire [11:0] add_534095;
  wire [11:0] sel_534097;
  wire [11:0] add_534099;
  wire [11:0] sel_534101;
  wire [15:0] add_534105;
  wire [10:0] add_534115;
  wire [11:0] sel_534117;
  wire [10:0] add_534119;
  wire [11:0] sel_534121;
  wire [11:0] add_534131;
  wire [11:0] sel_534133;
  wire [11:0] add_534135;
  wire [11:0] sel_534137;
  wire [11:0] add_534149;
  wire [11:0] sel_534151;
  wire [11:0] add_534153;
  wire [11:0] sel_534155;
  wire [11:0] add_534167;
  wire [11:0] sel_534169;
  wire [11:0] add_534171;
  wire [11:0] sel_534173;
  wire [8:0] add_534185;
  wire [11:0] sel_534187;
  wire [8:0] add_534189;
  wire [11:0] sel_534191;
  wire [11:0] add_534201;
  wire [11:0] sel_534203;
  wire [11:0] add_534205;
  wire [11:0] sel_534207;
  wire [11:0] add_534219;
  wire [11:0] sel_534221;
  wire [11:0] add_534223;
  wire [11:0] sel_534225;
  wire [10:0] add_534237;
  wire [11:0] sel_534239;
  wire [10:0] add_534241;
  wire [11:0] sel_534243;
  wire [11:0] add_534253;
  wire [11:0] sel_534255;
  wire [11:0] add_534257;
  wire [11:0] sel_534259;
  wire [15:0] sel_534270;
  wire [11:0] add_534273;
  wire [11:0] sel_534275;
  wire [11:0] add_534277;
  wire [11:0] sel_534279;
  wire [11:0] add_534291;
  wire [11:0] sel_534293;
  wire [11:0] add_534295;
  wire [11:0] sel_534297;
  wire [10:0] add_534309;
  wire [11:0] sel_534311;
  wire [10:0] add_534313;
  wire [11:0] sel_534315;
  wire [10:0] add_534325;
  wire [11:0] sel_534327;
  wire [10:0] add_534329;
  wire [11:0] sel_534331;
  wire [9:0] add_534343;
  wire [11:0] sel_534345;
  wire [9:0] add_534347;
  wire [11:0] sel_534349;
  wire [11:0] add_534361;
  wire [11:0] sel_534363;
  wire [11:0] add_534365;
  wire [11:0] sel_534367;
  wire [10:0] add_534379;
  wire [11:0] sel_534381;
  wire [10:0] add_534383;
  wire [11:0] sel_534385;
  wire [10:0] add_534395;
  wire [11:0] sel_534397;
  wire [10:0] add_534399;
  wire [11:0] sel_534401;
  wire [11:0] add_534411;
  wire [11:0] sel_534413;
  wire [11:0] add_534415;
  wire [11:0] sel_534417;
  wire [11:0] add_534427;
  wire [11:0] sel_534429;
  wire [11:0] add_534431;
  wire [11:0] sel_534433;
  wire [15:0] add_534437;
  wire [9:0] add_534443;
  wire [11:0] sel_534445;
  wire [9:0] add_534447;
  wire [11:0] sel_534449;
  wire [7:0] add_534461;
  wire [11:0] sel_534463;
  wire [7:0] add_534465;
  wire [11:0] sel_534467;
  wire [11:0] add_534477;
  wire [11:0] sel_534479;
  wire [11:0] add_534481;
  wire [11:0] sel_534483;
  wire [10:0] add_534493;
  wire [11:0] sel_534495;
  wire [10:0] add_534497;
  wire [11:0] sel_534499;
  wire [8:0] add_534509;
  wire [11:0] sel_534511;
  wire [8:0] add_534513;
  wire [11:0] sel_534515;
  wire [8:0] add_534527;
  wire [11:0] sel_534529;
  wire [8:0] add_534531;
  wire [11:0] sel_534533;
  wire [11:0] add_534543;
  wire [11:0] sel_534545;
  wire [11:0] add_534547;
  wire [11:0] sel_534549;
  wire [11:0] add_534559;
  wire [11:0] sel_534561;
  wire [11:0] add_534563;
  wire [11:0] sel_534565;
  wire [11:0] add_534577;
  wire [11:0] sel_534579;
  wire [11:0] add_534581;
  wire [11:0] sel_534583;
  wire [15:0] sel_534594;
  wire [10:0] add_534605;
  wire [11:0] sel_534607;
  wire [10:0] add_534609;
  wire [11:0] sel_534611;
  wire [11:0] add_534621;
  wire [11:0] sel_534623;
  wire [11:0] add_534625;
  wire [11:0] sel_534627;
  wire [11:0] add_534639;
  wire [11:0] sel_534641;
  wire [11:0] add_534643;
  wire [11:0] sel_534645;
  wire [11:0] add_534657;
  wire [11:0] sel_534659;
  wire [11:0] add_534661;
  wire [11:0] sel_534663;
  wire [8:0] add_534675;
  wire [11:0] sel_534677;
  wire [8:0] add_534679;
  wire [11:0] sel_534681;
  wire [11:0] add_534691;
  wire [11:0] sel_534693;
  wire [11:0] add_534695;
  wire [11:0] sel_534697;
  wire [11:0] add_534709;
  wire [11:0] sel_534711;
  wire [11:0] add_534713;
  wire [11:0] sel_534715;
  wire [10:0] add_534727;
  wire [11:0] sel_534729;
  wire [10:0] add_534731;
  wire [11:0] sel_534733;
  wire [11:0] add_534743;
  wire [11:0] sel_534745;
  wire [11:0] add_534747;
  wire [11:0] sel_534749;
  wire [15:0] add_534753;
  wire [11:0] add_534755;
  wire [11:0] sel_534757;
  wire [11:0] add_534759;
  wire [11:0] sel_534761;
  wire [11:0] add_534773;
  wire [11:0] sel_534775;
  wire [11:0] add_534777;
  wire [11:0] sel_534779;
  wire [10:0] add_534791;
  wire [11:0] sel_534793;
  wire [10:0] add_534795;
  wire [11:0] sel_534797;
  wire [10:0] add_534807;
  wire [11:0] sel_534809;
  wire [10:0] add_534811;
  wire [11:0] sel_534813;
  wire [9:0] add_534825;
  wire [11:0] sel_534827;
  wire [9:0] add_534829;
  wire [11:0] sel_534831;
  wire [11:0] add_534843;
  wire [11:0] sel_534845;
  wire [11:0] add_534847;
  wire [11:0] sel_534849;
  wire [10:0] add_534861;
  wire [11:0] sel_534863;
  wire [10:0] add_534865;
  wire [11:0] sel_534867;
  wire [10:0] add_534877;
  wire [11:0] sel_534879;
  wire [10:0] add_534881;
  wire [11:0] sel_534883;
  wire [11:0] add_534893;
  wire [11:0] sel_534895;
  wire [11:0] add_534897;
  wire [11:0] sel_534899;
  wire [15:0] sel_534910;
  wire [9:0] add_534917;
  wire [11:0] sel_534919;
  wire [9:0] add_534921;
  wire [11:0] sel_534923;
  wire [7:0] add_534935;
  wire [11:0] sel_534937;
  wire [7:0] add_534939;
  wire [11:0] sel_534941;
  wire [11:0] add_534951;
  wire [11:0] sel_534953;
  wire [11:0] add_534955;
  wire [11:0] sel_534957;
  wire [10:0] add_534967;
  wire [11:0] sel_534969;
  wire [10:0] add_534971;
  wire [11:0] sel_534973;
  wire [8:0] add_534983;
  wire [11:0] sel_534985;
  wire [8:0] add_534987;
  wire [11:0] sel_534989;
  wire [8:0] add_535001;
  wire [11:0] sel_535003;
  wire [8:0] add_535005;
  wire [11:0] sel_535007;
  wire [11:0] add_535017;
  wire [11:0] sel_535019;
  wire [11:0] add_535021;
  wire [11:0] sel_535023;
  wire [11:0] add_535033;
  wire [11:0] sel_535035;
  wire [11:0] add_535037;
  wire [11:0] sel_535039;
  wire [11:0] add_535051;
  wire [11:0] sel_535053;
  wire [11:0] add_535055;
  wire [11:0] sel_535057;
  wire [15:0] add_535061;
  wire [10:0] add_535071;
  wire [11:0] sel_535073;
  wire [10:0] add_535075;
  wire [11:0] sel_535077;
  wire [11:0] add_535087;
  wire [11:0] sel_535089;
  wire [11:0] add_535091;
  wire [11:0] sel_535093;
  wire [11:0] add_535105;
  wire [11:0] sel_535107;
  wire [11:0] add_535109;
  wire [11:0] sel_535111;
  wire [11:0] add_535123;
  wire [11:0] sel_535125;
  wire [11:0] add_535127;
  wire [11:0] sel_535129;
  wire [8:0] add_535141;
  wire [11:0] sel_535143;
  wire [8:0] add_535145;
  wire [11:0] sel_535147;
  wire [11:0] add_535157;
  wire [11:0] sel_535159;
  wire [11:0] add_535161;
  wire [11:0] sel_535163;
  wire [11:0] add_535175;
  wire [11:0] sel_535177;
  wire [11:0] add_535179;
  wire [11:0] sel_535181;
  wire [10:0] add_535193;
  wire [11:0] sel_535195;
  wire [10:0] add_535197;
  wire [11:0] sel_535199;
  wire [15:0] sel_535210;
  wire [11:0] add_535213;
  wire [11:0] sel_535215;
  wire [11:0] add_535217;
  wire [11:0] sel_535219;
  wire [11:0] add_535231;
  wire [11:0] sel_535233;
  wire [11:0] add_535235;
  wire [11:0] sel_535237;
  wire [10:0] add_535249;
  wire [11:0] sel_535251;
  wire [10:0] add_535253;
  wire [11:0] sel_535255;
  wire [10:0] add_535265;
  wire [11:0] sel_535267;
  wire [10:0] add_535269;
  wire [11:0] sel_535271;
  wire [9:0] add_535283;
  wire [11:0] sel_535285;
  wire [9:0] add_535287;
  wire [11:0] sel_535289;
  wire [11:0] add_535301;
  wire [11:0] sel_535303;
  wire [11:0] add_535305;
  wire [11:0] sel_535307;
  wire [10:0] add_535319;
  wire [11:0] sel_535321;
  wire [10:0] add_535323;
  wire [11:0] sel_535325;
  wire [10:0] add_535335;
  wire [11:0] sel_535337;
  wire [10:0] add_535339;
  wire [11:0] sel_535341;
  wire [11:0] add_535351;
  wire [11:0] sel_535353;
  wire [11:0] add_535355;
  wire [11:0] sel_535357;
  wire [15:0] add_535361;
  wire [9:0] add_535367;
  wire [11:0] sel_535369;
  wire [9:0] add_535371;
  wire [11:0] sel_535373;
  wire [7:0] add_535385;
  wire [11:0] sel_535387;
  wire [7:0] add_535389;
  wire [11:0] sel_535391;
  wire [11:0] add_535401;
  wire [11:0] sel_535403;
  wire [11:0] add_535405;
  wire [11:0] sel_535407;
  wire [10:0] add_535417;
  wire [11:0] sel_535419;
  wire [10:0] add_535421;
  wire [11:0] sel_535423;
  wire [8:0] add_535433;
  wire [11:0] sel_535435;
  wire [8:0] add_535437;
  wire [11:0] sel_535439;
  wire [8:0] add_535451;
  wire [11:0] sel_535453;
  wire [8:0] add_535455;
  wire [11:0] sel_535457;
  wire [11:0] add_535467;
  wire [11:0] sel_535469;
  wire [11:0] add_535471;
  wire [11:0] sel_535473;
  wire [11:0] add_535483;
  wire [11:0] sel_535485;
  wire [11:0] add_535487;
  wire [11:0] sel_535489;
  wire [15:0] sel_535502;
  wire [10:0] add_535513;
  wire [11:0] sel_535515;
  wire [10:0] add_535517;
  wire [11:0] sel_535519;
  wire [11:0] add_535529;
  wire [11:0] sel_535531;
  wire [11:0] add_535533;
  wire [11:0] sel_535535;
  wire [11:0] add_535547;
  wire [11:0] sel_535549;
  wire [11:0] add_535551;
  wire [11:0] sel_535553;
  wire [11:0] add_535565;
  wire [11:0] sel_535567;
  wire [11:0] add_535569;
  wire [11:0] sel_535571;
  wire [8:0] add_535583;
  wire [11:0] sel_535585;
  wire [8:0] add_535587;
  wire [11:0] sel_535589;
  wire [11:0] add_535599;
  wire [11:0] sel_535601;
  wire [11:0] add_535603;
  wire [11:0] sel_535605;
  wire [11:0] add_535617;
  wire [11:0] sel_535619;
  wire [11:0] add_535621;
  wire [11:0] sel_535623;
  wire [10:0] add_535635;
  wire [11:0] sel_535637;
  wire [10:0] add_535639;
  wire [11:0] sel_535641;
  wire [15:0] add_535645;
  wire [11:0] add_535647;
  wire [11:0] sel_535649;
  wire [11:0] add_535651;
  wire [11:0] sel_535653;
  wire [11:0] add_535665;
  wire [11:0] sel_535667;
  wire [11:0] add_535669;
  wire [11:0] sel_535671;
  wire [10:0] add_535683;
  wire [11:0] sel_535685;
  wire [10:0] add_535687;
  wire [11:0] sel_535689;
  wire [10:0] add_535699;
  wire [11:0] sel_535701;
  wire [10:0] add_535703;
  wire [11:0] sel_535705;
  wire [9:0] add_535717;
  wire [11:0] sel_535719;
  wire [9:0] add_535721;
  wire [11:0] sel_535723;
  wire [11:0] add_535735;
  wire [11:0] sel_535737;
  wire [11:0] add_535739;
  wire [11:0] sel_535741;
  wire [10:0] add_535753;
  wire [11:0] sel_535755;
  wire [10:0] add_535757;
  wire [11:0] sel_535759;
  wire [10:0] add_535769;
  wire [11:0] sel_535771;
  wire [10:0] add_535773;
  wire [11:0] sel_535775;
  wire [15:0] sel_535786;
  wire [9:0] add_535793;
  wire [11:0] sel_535795;
  wire [9:0] add_535797;
  wire [11:0] sel_535799;
  wire [7:0] add_535811;
  wire [11:0] sel_535813;
  wire [7:0] add_535815;
  wire [11:0] sel_535817;
  wire [11:0] add_535827;
  wire [11:0] sel_535829;
  wire [11:0] add_535831;
  wire [11:0] sel_535833;
  wire [10:0] add_535843;
  wire [11:0] sel_535845;
  wire [10:0] add_535847;
  wire [11:0] sel_535849;
  wire [8:0] add_535859;
  wire [11:0] sel_535861;
  wire [8:0] add_535863;
  wire [11:0] sel_535865;
  wire [8:0] add_535877;
  wire [11:0] sel_535879;
  wire [8:0] add_535881;
  wire [11:0] sel_535883;
  wire [11:0] add_535893;
  wire [11:0] sel_535895;
  wire [11:0] add_535897;
  wire [11:0] sel_535899;
  wire [11:0] add_535909;
  wire [11:0] sel_535911;
  wire [11:0] add_535913;
  wire [11:0] sel_535915;
  wire [15:0] add_535921;
  wire [10:0] add_535931;
  wire [11:0] sel_535933;
  wire [10:0] add_535935;
  wire [11:0] sel_535937;
  wire [11:0] add_535947;
  wire [11:0] sel_535949;
  wire [11:0] add_535951;
  wire [11:0] sel_535953;
  wire [11:0] add_535965;
  wire [11:0] sel_535967;
  wire [11:0] add_535969;
  wire [11:0] sel_535971;
  wire [11:0] add_535983;
  wire [11:0] sel_535985;
  wire [11:0] add_535987;
  wire [11:0] sel_535989;
  wire [8:0] add_536001;
  wire [11:0] sel_536003;
  wire [8:0] add_536005;
  wire [11:0] sel_536007;
  wire [11:0] add_536017;
  wire [11:0] sel_536019;
  wire [11:0] add_536021;
  wire [11:0] sel_536023;
  wire [11:0] add_536035;
  wire [11:0] sel_536037;
  wire [11:0] add_536039;
  wire [11:0] sel_536041;
  wire [15:0] sel_536054;
  wire [11:0] add_536057;
  wire [11:0] sel_536059;
  wire [11:0] add_536061;
  wire [11:0] sel_536063;
  wire [11:0] add_536075;
  wire [11:0] sel_536077;
  wire [11:0] add_536079;
  wire [11:0] sel_536081;
  wire [10:0] add_536093;
  wire [11:0] sel_536095;
  wire [10:0] add_536097;
  wire [11:0] sel_536099;
  wire [10:0] add_536109;
  wire [11:0] sel_536111;
  wire [10:0] add_536113;
  wire [11:0] sel_536115;
  wire [9:0] add_536127;
  wire [11:0] sel_536129;
  wire [9:0] add_536131;
  wire [11:0] sel_536133;
  wire [11:0] add_536145;
  wire [11:0] sel_536147;
  wire [11:0] add_536149;
  wire [11:0] sel_536151;
  wire [10:0] add_536163;
  wire [11:0] sel_536165;
  wire [10:0] add_536167;
  wire [11:0] sel_536169;
  wire [10:0] add_536179;
  wire [11:0] sel_536181;
  wire [10:0] add_536183;
  wire [11:0] sel_536185;
  wire [15:0] add_536189;
  wire [9:0] add_536195;
  wire [11:0] sel_536197;
  wire [9:0] add_536199;
  wire [11:0] sel_536201;
  wire [7:0] add_536213;
  wire [11:0] sel_536215;
  wire [7:0] add_536217;
  wire [11:0] sel_536219;
  wire [11:0] add_536229;
  wire [11:0] sel_536231;
  wire [11:0] add_536233;
  wire [11:0] sel_536235;
  wire [10:0] add_536245;
  wire [11:0] sel_536247;
  wire [10:0] add_536249;
  wire [11:0] sel_536251;
  wire [8:0] add_536261;
  wire [11:0] sel_536263;
  wire [8:0] add_536265;
  wire [11:0] sel_536267;
  wire [8:0] add_536279;
  wire [11:0] sel_536281;
  wire [8:0] add_536283;
  wire [11:0] sel_536285;
  wire [11:0] add_536295;
  wire [11:0] sel_536297;
  wire [11:0] add_536299;
  wire [11:0] sel_536301;
  wire [15:0] sel_536312;
  wire [10:0] add_536323;
  wire [11:0] sel_536325;
  wire [10:0] add_536327;
  wire [11:0] sel_536329;
  wire [11:0] add_536339;
  wire [11:0] sel_536341;
  wire [11:0] add_536343;
  wire [11:0] sel_536345;
  wire [11:0] add_536357;
  wire [11:0] sel_536359;
  wire [11:0] add_536361;
  wire [11:0] sel_536363;
  wire [11:0] add_536375;
  wire [11:0] sel_536377;
  wire [11:0] add_536379;
  wire [11:0] sel_536381;
  wire [8:0] add_536393;
  wire [11:0] sel_536395;
  wire [8:0] add_536397;
  wire [11:0] sel_536399;
  wire [11:0] add_536409;
  wire [11:0] sel_536411;
  wire [11:0] add_536413;
  wire [11:0] sel_536415;
  wire [11:0] add_536427;
  wire [11:0] sel_536429;
  wire [11:0] add_536431;
  wire [11:0] sel_536433;
  wire [15:0] add_536439;
  wire [11:0] add_536441;
  wire [11:0] sel_536443;
  wire [11:0] add_536445;
  wire [11:0] sel_536447;
  wire [11:0] add_536459;
  wire [11:0] sel_536461;
  wire [11:0] add_536463;
  wire [11:0] sel_536465;
  wire [10:0] add_536477;
  wire [11:0] sel_536479;
  wire [10:0] add_536481;
  wire [11:0] sel_536483;
  wire [10:0] add_536493;
  wire [11:0] sel_536495;
  wire [10:0] add_536497;
  wire [11:0] sel_536499;
  wire [9:0] add_536511;
  wire [11:0] sel_536513;
  wire [9:0] add_536515;
  wire [11:0] sel_536517;
  wire [11:0] add_536529;
  wire [11:0] sel_536531;
  wire [11:0] add_536533;
  wire [11:0] sel_536535;
  wire [10:0] add_536547;
  wire [11:0] sel_536549;
  wire [10:0] add_536551;
  wire [11:0] sel_536553;
  wire [15:0] sel_536564;
  wire [9:0] add_536571;
  wire [11:0] sel_536573;
  wire [9:0] add_536575;
  wire [11:0] sel_536577;
  wire [7:0] add_536589;
  wire [11:0] sel_536591;
  wire [7:0] add_536593;
  wire [11:0] sel_536595;
  wire [11:0] add_536605;
  wire [11:0] sel_536607;
  wire [11:0] add_536609;
  wire [11:0] sel_536611;
  wire [10:0] add_536621;
  wire [11:0] sel_536623;
  wire [10:0] add_536625;
  wire [11:0] sel_536627;
  wire [8:0] add_536637;
  wire [11:0] sel_536639;
  wire [8:0] add_536641;
  wire [11:0] sel_536643;
  wire [8:0] add_536655;
  wire [11:0] sel_536657;
  wire [8:0] add_536659;
  wire [11:0] sel_536661;
  wire [11:0] add_536671;
  wire [11:0] sel_536673;
  wire [11:0] add_536675;
  wire [11:0] sel_536677;
  wire [15:0] add_536681;
  wire [10:0] add_536691;
  wire [11:0] sel_536693;
  wire [10:0] add_536695;
  wire [11:0] sel_536697;
  wire [11:0] add_536707;
  wire [11:0] sel_536709;
  wire [11:0] add_536711;
  wire [11:0] sel_536713;
  wire [11:0] add_536725;
  wire [11:0] sel_536727;
  wire [11:0] add_536729;
  wire [11:0] sel_536731;
  wire [11:0] add_536743;
  wire [11:0] sel_536745;
  wire [11:0] add_536747;
  wire [11:0] sel_536749;
  wire [8:0] add_536761;
  wire [11:0] sel_536763;
  wire [8:0] add_536765;
  wire [11:0] sel_536767;
  wire [11:0] add_536777;
  wire [11:0] sel_536779;
  wire [11:0] add_536781;
  wire [11:0] sel_536783;
  wire [15:0] sel_536796;
  wire [11:0] add_536799;
  wire [11:0] sel_536801;
  wire [11:0] add_536803;
  wire [11:0] sel_536805;
  wire [11:0] add_536817;
  wire [11:0] sel_536819;
  wire [11:0] add_536821;
  wire [11:0] sel_536823;
  wire [10:0] add_536835;
  wire [11:0] sel_536837;
  wire [10:0] add_536839;
  wire [11:0] sel_536841;
  wire [10:0] add_536851;
  wire [11:0] sel_536853;
  wire [10:0] add_536855;
  wire [11:0] sel_536857;
  wire [9:0] add_536869;
  wire [11:0] sel_536871;
  wire [9:0] add_536873;
  wire [11:0] sel_536875;
  wire [11:0] add_536887;
  wire [11:0] sel_536889;
  wire [11:0] add_536891;
  wire [11:0] sel_536893;
  wire [10:0] add_536905;
  wire [11:0] sel_536907;
  wire [10:0] add_536909;
  wire [11:0] sel_536911;
  wire [15:0] add_536915;
  wire [9:0] add_536921;
  wire [11:0] sel_536923;
  wire [9:0] add_536925;
  wire [11:0] sel_536927;
  wire [7:0] add_536939;
  wire [11:0] sel_536941;
  wire [7:0] add_536943;
  wire [11:0] sel_536945;
  wire [11:0] add_536955;
  wire [11:0] sel_536957;
  wire [11:0] add_536959;
  wire [11:0] sel_536961;
  wire [10:0] add_536971;
  wire [11:0] sel_536973;
  wire [10:0] add_536975;
  wire [11:0] sel_536977;
  wire [8:0] add_536987;
  wire [11:0] sel_536989;
  wire [8:0] add_536991;
  wire [11:0] sel_536993;
  wire [8:0] add_537005;
  wire [11:0] sel_537007;
  wire [8:0] add_537009;
  wire [11:0] sel_537011;
  wire [15:0] sel_537022;
  wire [10:0] add_537033;
  wire [11:0] sel_537035;
  wire [10:0] add_537037;
  wire [11:0] sel_537039;
  wire [11:0] add_537049;
  wire [11:0] sel_537051;
  wire [11:0] add_537053;
  wire [11:0] sel_537055;
  wire [11:0] add_537067;
  wire [11:0] sel_537069;
  wire [11:0] add_537071;
  wire [11:0] sel_537073;
  wire [11:0] add_537085;
  wire [11:0] sel_537087;
  wire [11:0] add_537089;
  wire [11:0] sel_537091;
  wire [8:0] add_537103;
  wire [11:0] sel_537105;
  wire [8:0] add_537107;
  wire [11:0] sel_537109;
  wire [11:0] add_537119;
  wire [11:0] sel_537121;
  wire [11:0] add_537123;
  wire [11:0] sel_537125;
  wire [15:0] add_537131;
  wire [11:0] add_537133;
  wire [11:0] sel_537135;
  wire [11:0] add_537137;
  wire [11:0] sel_537139;
  wire [11:0] add_537151;
  wire [11:0] sel_537153;
  wire [11:0] add_537155;
  wire [11:0] sel_537157;
  wire [10:0] add_537169;
  wire [11:0] sel_537171;
  wire [10:0] add_537173;
  wire [11:0] sel_537175;
  wire [10:0] add_537185;
  wire [11:0] sel_537187;
  wire [10:0] add_537189;
  wire [11:0] sel_537191;
  wire [9:0] add_537203;
  wire [11:0] sel_537205;
  wire [9:0] add_537207;
  wire [11:0] sel_537209;
  wire [11:0] add_537221;
  wire [11:0] sel_537223;
  wire [11:0] add_537225;
  wire [11:0] sel_537227;
  wire [15:0] sel_537240;
  wire [9:0] add_537247;
  wire [11:0] sel_537249;
  wire [9:0] add_537251;
  wire [11:0] sel_537253;
  wire [7:0] add_537265;
  wire [11:0] sel_537267;
  wire [7:0] add_537269;
  wire [11:0] sel_537271;
  wire [11:0] add_537281;
  wire [11:0] sel_537283;
  wire [11:0] add_537285;
  wire [11:0] sel_537287;
  wire [10:0] add_537297;
  wire [11:0] sel_537299;
  wire [10:0] add_537301;
  wire [11:0] sel_537303;
  wire [8:0] add_537313;
  wire [11:0] sel_537315;
  wire [8:0] add_537317;
  wire [11:0] sel_537319;
  wire [8:0] add_537331;
  wire [11:0] sel_537333;
  wire [8:0] add_537335;
  wire [11:0] sel_537337;
  wire [15:0] add_537341;
  wire [10:0] add_537351;
  wire [11:0] sel_537353;
  wire [10:0] add_537355;
  wire [11:0] sel_537357;
  wire [11:0] add_537367;
  wire [11:0] sel_537369;
  wire [11:0] add_537371;
  wire [11:0] sel_537373;
  wire [11:0] add_537385;
  wire [11:0] sel_537387;
  wire [11:0] add_537389;
  wire [11:0] sel_537391;
  wire [11:0] add_537403;
  wire [11:0] sel_537405;
  wire [11:0] add_537407;
  wire [11:0] sel_537409;
  wire [8:0] add_537421;
  wire [11:0] sel_537423;
  wire [8:0] add_537425;
  wire [11:0] sel_537427;
  wire [15:0] sel_537438;
  wire [11:0] add_537441;
  wire [11:0] sel_537443;
  wire [11:0] add_537445;
  wire [11:0] sel_537447;
  wire [11:0] add_537459;
  wire [11:0] sel_537461;
  wire [11:0] add_537463;
  wire [11:0] sel_537465;
  wire [10:0] add_537477;
  wire [11:0] sel_537479;
  wire [10:0] add_537481;
  wire [11:0] sel_537483;
  wire [10:0] add_537493;
  wire [11:0] sel_537495;
  wire [10:0] add_537497;
  wire [11:0] sel_537499;
  wire [9:0] add_537511;
  wire [11:0] sel_537513;
  wire [9:0] add_537515;
  wire [11:0] sel_537517;
  wire [11:0] add_537529;
  wire [11:0] sel_537531;
  wire [11:0] add_537533;
  wire [11:0] sel_537535;
  wire [15:0] add_537541;
  wire [9:0] add_537547;
  wire [11:0] sel_537549;
  wire [9:0] add_537551;
  wire [11:0] sel_537553;
  wire [7:0] add_537565;
  wire [11:0] sel_537567;
  wire [7:0] add_537569;
  wire [11:0] sel_537571;
  wire [11:0] add_537581;
  wire [11:0] sel_537583;
  wire [11:0] add_537585;
  wire [11:0] sel_537587;
  wire [10:0] add_537597;
  wire [11:0] sel_537599;
  wire [10:0] add_537601;
  wire [11:0] sel_537603;
  wire [8:0] add_537613;
  wire [11:0] sel_537615;
  wire [8:0] add_537617;
  wire [11:0] sel_537619;
  wire [15:0] sel_537632;
  wire [10:0] add_537643;
  wire [11:0] sel_537645;
  wire [10:0] add_537647;
  wire [11:0] sel_537649;
  wire [11:0] add_537659;
  wire [11:0] sel_537661;
  wire [11:0] add_537663;
  wire [11:0] sel_537665;
  wire [11:0] add_537677;
  wire [11:0] sel_537679;
  wire [11:0] add_537681;
  wire [11:0] sel_537683;
  wire [11:0] add_537695;
  wire [11:0] sel_537697;
  wire [11:0] add_537699;
  wire [11:0] sel_537701;
  wire [8:0] add_537713;
  wire [11:0] sel_537715;
  wire [8:0] add_537717;
  wire [11:0] sel_537719;
  wire [15:0] add_537723;
  wire [11:0] add_537725;
  wire [11:0] sel_537727;
  wire [11:0] add_537729;
  wire [11:0] sel_537731;
  wire [11:0] add_537743;
  wire [11:0] sel_537745;
  wire [11:0] add_537747;
  wire [11:0] sel_537749;
  wire [10:0] add_537761;
  wire [11:0] sel_537763;
  wire [10:0] add_537765;
  wire [11:0] sel_537767;
  wire [10:0] add_537777;
  wire [11:0] sel_537779;
  wire [10:0] add_537781;
  wire [11:0] sel_537783;
  wire [9:0] add_537795;
  wire [11:0] sel_537797;
  wire [9:0] add_537799;
  wire [11:0] sel_537801;
  wire [15:0] sel_537814;
  wire [9:0] add_537821;
  wire [11:0] sel_537823;
  wire [9:0] add_537825;
  wire [11:0] sel_537827;
  wire [7:0] add_537839;
  wire [11:0] sel_537841;
  wire [7:0] add_537843;
  wire [11:0] sel_537845;
  wire [11:0] add_537855;
  wire [11:0] sel_537857;
  wire [11:0] add_537859;
  wire [11:0] sel_537861;
  wire [10:0] add_537871;
  wire [11:0] sel_537873;
  wire [10:0] add_537875;
  wire [11:0] sel_537877;
  wire [8:0] add_537887;
  wire [11:0] sel_537889;
  wire [8:0] add_537891;
  wire [11:0] sel_537893;
  wire [15:0] add_537899;
  wire [10:0] add_537909;
  wire [11:0] sel_537911;
  wire [10:0] add_537913;
  wire [11:0] sel_537915;
  wire [11:0] add_537925;
  wire [11:0] sel_537927;
  wire [11:0] add_537929;
  wire [11:0] sel_537931;
  wire [11:0] add_537943;
  wire [11:0] sel_537945;
  wire [11:0] add_537947;
  wire [11:0] sel_537949;
  wire [11:0] add_537961;
  wire [11:0] sel_537963;
  wire [11:0] add_537965;
  wire [11:0] sel_537967;
  wire [15:0] sel_537980;
  wire [11:0] add_537983;
  wire [11:0] sel_537985;
  wire [11:0] add_537987;
  wire [11:0] sel_537989;
  wire [11:0] add_538001;
  wire [11:0] sel_538003;
  wire [11:0] add_538005;
  wire [11:0] sel_538007;
  wire [10:0] add_538019;
  wire [11:0] sel_538021;
  wire [10:0] add_538023;
  wire [11:0] sel_538025;
  wire [10:0] add_538035;
  wire [11:0] sel_538037;
  wire [10:0] add_538039;
  wire [11:0] sel_538041;
  wire [9:0] add_538053;
  wire [11:0] sel_538055;
  wire [9:0] add_538057;
  wire [11:0] sel_538059;
  wire [15:0] add_538065;
  wire [9:0] add_538071;
  wire [11:0] sel_538073;
  wire [9:0] add_538075;
  wire [11:0] sel_538077;
  wire [7:0] add_538089;
  wire [11:0] sel_538091;
  wire [7:0] add_538093;
  wire [11:0] sel_538095;
  wire [11:0] add_538105;
  wire [11:0] sel_538107;
  wire [11:0] add_538109;
  wire [11:0] sel_538111;
  wire [10:0] add_538121;
  wire [11:0] sel_538123;
  wire [10:0] add_538125;
  wire [11:0] sel_538127;
  wire [15:0] sel_538138;
  wire [10:0] add_538149;
  wire [11:0] sel_538151;
  wire [10:0] add_538153;
  wire [11:0] sel_538155;
  wire [11:0] add_538165;
  wire [11:0] sel_538167;
  wire [11:0] add_538169;
  wire [11:0] sel_538171;
  wire [11:0] add_538183;
  wire [11:0] sel_538185;
  wire [11:0] add_538187;
  wire [11:0] sel_538189;
  wire [11:0] add_538201;
  wire [11:0] sel_538203;
  wire [11:0] add_538205;
  wire [11:0] sel_538207;
  wire [15:0] add_538213;
  wire [11:0] add_538215;
  wire [11:0] sel_538217;
  wire [11:0] add_538219;
  wire [11:0] sel_538221;
  wire [11:0] add_538233;
  wire [11:0] sel_538235;
  wire [11:0] add_538237;
  wire [11:0] sel_538239;
  wire [10:0] add_538251;
  wire [11:0] sel_538253;
  wire [10:0] add_538255;
  wire [11:0] sel_538257;
  wire [10:0] add_538267;
  wire [11:0] sel_538269;
  wire [10:0] add_538271;
  wire [11:0] sel_538273;
  wire [15:0] sel_538286;
  wire [9:0] add_538293;
  wire [11:0] sel_538295;
  wire [9:0] add_538297;
  wire [11:0] sel_538299;
  wire [7:0] add_538311;
  wire [11:0] sel_538313;
  wire [7:0] add_538315;
  wire [11:0] sel_538317;
  wire [11:0] add_538327;
  wire [11:0] sel_538329;
  wire [11:0] add_538331;
  wire [11:0] sel_538333;
  wire [10:0] add_538343;
  wire [11:0] sel_538345;
  wire [10:0] add_538347;
  wire [11:0] sel_538349;
  wire [15:0] add_538353;
  wire [10:0] add_538363;
  wire [11:0] sel_538365;
  wire [10:0] add_538367;
  wire [11:0] sel_538369;
  wire [11:0] add_538379;
  wire [11:0] sel_538381;
  wire [11:0] add_538383;
  wire [11:0] sel_538385;
  wire [11:0] add_538397;
  wire [11:0] sel_538399;
  wire [11:0] add_538401;
  wire [11:0] sel_538403;
  wire [15:0] sel_538416;
  wire [11:0] add_538419;
  wire [11:0] sel_538421;
  wire [11:0] add_538423;
  wire [11:0] sel_538425;
  wire [11:0] add_538437;
  wire [11:0] sel_538439;
  wire [11:0] add_538441;
  wire [11:0] sel_538443;
  wire [10:0] add_538455;
  wire [11:0] sel_538457;
  wire [10:0] add_538459;
  wire [11:0] sel_538461;
  wire [10:0] add_538471;
  wire [11:0] sel_538473;
  wire [10:0] add_538475;
  wire [11:0] sel_538477;
  wire [15:0] add_538483;
  wire [9:0] add_538489;
  wire [11:0] sel_538491;
  wire [9:0] add_538493;
  wire [11:0] sel_538495;
  wire [7:0] add_538507;
  wire [11:0] sel_538509;
  wire [7:0] add_538511;
  wire [11:0] sel_538513;
  wire [11:0] add_538523;
  wire [11:0] sel_538525;
  wire [11:0] add_538527;
  wire [11:0] sel_538529;
  wire [15:0] sel_538540;
  wire [10:0] add_538551;
  wire [11:0] sel_538553;
  wire [10:0] add_538555;
  wire [11:0] sel_538557;
  wire [11:0] add_538567;
  wire [11:0] sel_538569;
  wire [11:0] add_538571;
  wire [11:0] sel_538573;
  wire [11:0] add_538585;
  wire [11:0] sel_538587;
  wire [11:0] add_538589;
  wire [11:0] sel_538591;
  wire [15:0] add_538597;
  wire [11:0] add_538599;
  wire [11:0] sel_538601;
  wire [11:0] add_538603;
  wire [11:0] sel_538605;
  wire [11:0] add_538617;
  wire [11:0] sel_538619;
  wire [11:0] add_538621;
  wire [11:0] sel_538623;
  wire [10:0] add_538635;
  wire [11:0] sel_538637;
  wire [10:0] add_538639;
  wire [11:0] sel_538641;
  wire [15:0] sel_538652;
  wire [9:0] add_538659;
  wire [11:0] sel_538661;
  wire [9:0] add_538663;
  wire [11:0] sel_538665;
  wire [7:0] add_538677;
  wire [11:0] sel_538679;
  wire [7:0] add_538681;
  wire [11:0] sel_538683;
  wire [11:0] add_538693;
  wire [11:0] sel_538695;
  wire [11:0] add_538697;
  wire [11:0] sel_538699;
  wire [15:0] add_538703;
  wire [10:0] add_538713;
  wire [11:0] sel_538715;
  wire [10:0] add_538717;
  wire [11:0] sel_538719;
  wire [11:0] add_538729;
  wire [11:0] sel_538731;
  wire [11:0] add_538733;
  wire [11:0] sel_538735;
  wire [15:0] sel_538748;
  wire [11:0] add_538751;
  wire [11:0] sel_538753;
  wire [11:0] add_538755;
  wire [11:0] sel_538757;
  wire [11:0] add_538769;
  wire [11:0] sel_538771;
  wire [11:0] add_538773;
  wire [11:0] sel_538775;
  wire [10:0] add_538787;
  wire [11:0] sel_538789;
  wire [10:0] add_538791;
  wire [11:0] sel_538793;
  wire [15:0] add_538797;
  wire [9:0] add_538803;
  wire [11:0] sel_538805;
  wire [9:0] add_538807;
  wire [11:0] sel_538809;
  wire [7:0] add_538821;
  wire [11:0] sel_538823;
  wire [7:0] add_538825;
  wire [11:0] sel_538827;
  wire [15:0] sel_538838;
  wire [10:0] add_538849;
  wire [11:0] sel_538851;
  wire [10:0] add_538853;
  wire [11:0] sel_538855;
  wire [11:0] add_538865;
  wire [11:0] sel_538867;
  wire [11:0] add_538869;
  wire [11:0] sel_538871;
  wire [15:0] add_538877;
  wire [11:0] add_538879;
  wire [11:0] sel_538881;
  wire [11:0] add_538883;
  wire [11:0] sel_538885;
  wire [11:0] add_538897;
  wire [11:0] sel_538899;
  wire [11:0] add_538901;
  wire [11:0] sel_538903;
  wire [15:0] sel_538916;
  wire [9:0] add_538923;
  wire [11:0] sel_538925;
  wire [9:0] add_538927;
  wire [11:0] sel_538929;
  wire [7:0] add_538941;
  wire [11:0] sel_538943;
  wire [7:0] add_538945;
  wire [11:0] sel_538947;
  wire [15:0] add_538951;
  wire [10:0] add_538961;
  wire [11:0] sel_538963;
  wire [10:0] add_538965;
  wire [11:0] sel_538967;
  wire [15:0] sel_538978;
  wire [11:0] add_538981;
  wire [11:0] sel_538983;
  wire [11:0] add_538985;
  wire [11:0] sel_538987;
  wire [11:0] add_538999;
  wire [11:0] sel_539001;
  wire [11:0] add_539003;
  wire [11:0] sel_539005;
  wire [15:0] add_539011;
  wire [9:0] add_539017;
  wire [11:0] sel_539019;
  wire [9:0] add_539021;
  wire [11:0] sel_539023;
  wire [15:0] sel_539036;
  wire [10:0] add_539047;
  wire [11:0] sel_539049;
  wire [10:0] add_539051;
  wire [11:0] sel_539053;
  wire [15:0] add_539057;
  wire [11:0] add_539059;
  wire [11:0] sel_539061;
  wire [11:0] add_539063;
  wire [11:0] sel_539065;
  wire [15:0] sel_539078;
  wire [9:0] add_539085;
  wire [11:0] sel_539087;
  wire [9:0] add_539089;
  wire [11:0] sel_539091;
  wire [15:0] add_539097;
  wire [15:0] sel_539108;
  wire [11:0] add_539111;
  wire [11:0] sel_539113;
  wire [11:0] add_539115;
  wire [11:0] sel_539117;
  wire [15:0] add_539123;
  wire [15:0] sel_539130;
  wire [15:0] add_539135;
  wire [15:0] sel_539138;
  wire [15:0] add_539141;
  assign array_index_512818 = set1_unflattened[5'h00];
  assign array_index_512819 = set2_unflattened[5'h00];
  assign add_512826 = array_index_512818[11:0] + 12'h62b;
  assign add_512829 = array_index_512819[11:0] + 12'h62b;
  assign array_index_512834 = set1_unflattened[5'h01];
  assign array_index_512837 = set2_unflattened[5'h01];
  assign add_512841 = array_index_512818[11:1] + 11'h24f;
  assign add_512844 = array_index_512819[11:1] + 11'h24f;
  assign add_512860 = array_index_512834[11:0] + 12'h62b;
  assign sel_512862 = $signed({1'h0, add_512826}) < $signed(13'h0fff) ? add_512826 : 12'hfff;
  assign add_512865 = array_index_512837[11:0] + 12'h62b;
  assign sel_512867 = $signed({1'h0, add_512829}) < $signed(13'h0fff) ? add_512829 : 12'hfff;
  assign array_index_512880 = set1_unflattened[5'h02];
  assign array_index_512883 = set2_unflattened[5'h02];
  assign add_512887 = array_index_512818[11:1] + 11'h75d;
  assign add_512889 = array_index_512819[11:1] + 11'h75d;
  assign add_512891 = array_index_512834[11:1] + 11'h24f;
  assign sel_512894 = $signed({1'h0, add_512841, array_index_512818[0]}) < $signed(13'h0fff) ? {add_512841, array_index_512818[0]} : 12'hfff;
  assign add_512896 = array_index_512837[11:1] + 11'h24f;
  assign sel_512899 = $signed({1'h0, add_512844, array_index_512819[0]}) < $signed(13'h0fff) ? {add_512844, array_index_512819[0]} : 12'hfff;
  assign add_512916 = array_index_512880[11:0] + 12'h62b;
  assign sel_512918 = $signed({1'h0, add_512860}) < $signed({1'h0, sel_512862}) ? add_512860 : sel_512862;
  assign add_512921 = array_index_512883[11:0] + 12'h62b;
  assign sel_512923 = $signed({1'h0, add_512865}) < $signed({1'h0, sel_512867}) ? add_512865 : sel_512867;
  assign array_index_512942 = set1_unflattened[5'h03];
  assign array_index_512945 = set2_unflattened[5'h03];
  assign add_512949 = array_index_512818[11:1] + 11'h6cb;
  assign add_512951 = array_index_512819[11:1] + 11'h6cb;
  assign add_512953 = array_index_512834[11:1] + 11'h75d;
  assign sel_512955 = $signed({1'h0, add_512887, array_index_512818[0]}) < $signed(13'h0fff) ? {add_512887, array_index_512818[0]} : 12'hfff;
  assign add_512957 = array_index_512837[11:1] + 11'h75d;
  assign sel_512959 = $signed({1'h0, add_512889, array_index_512819[0]}) < $signed(13'h0fff) ? {add_512889, array_index_512819[0]} : 12'hfff;
  assign add_512961 = array_index_512880[11:1] + 11'h24f;
  assign sel_512964 = $signed({1'h0, add_512891, array_index_512834[0]}) < $signed({1'h0, sel_512894}) ? {add_512891, array_index_512834[0]} : sel_512894;
  assign add_512966 = array_index_512883[11:1] + 11'h24f;
  assign sel_512969 = $signed({1'h0, add_512896, array_index_512837[0]}) < $signed({1'h0, sel_512899}) ? {add_512896, array_index_512837[0]} : sel_512899;
  assign add_512990 = array_index_512942[11:0] + 12'h62b;
  assign sel_512992 = $signed({1'h0, add_512916}) < $signed({1'h0, sel_512918}) ? add_512916 : sel_512918;
  assign add_512995 = array_index_512945[11:0] + 12'h62b;
  assign sel_512997 = $signed({1'h0, add_512921}) < $signed({1'h0, sel_512923}) ? add_512921 : sel_512923;
  assign array_index_513022 = set1_unflattened[5'h04];
  assign array_index_513025 = set2_unflattened[5'h04];
  assign add_513029 = array_index_512818[11:0] + 12'ha09;
  assign add_513031 = array_index_512819[11:0] + 12'ha09;
  assign add_513033 = array_index_512834[11:1] + 11'h6cb;
  assign sel_513035 = $signed({1'h0, add_512949, array_index_512818[0]}) < $signed(13'h0fff) ? {add_512949, array_index_512818[0]} : 12'hfff;
  assign add_513037 = array_index_512837[11:1] + 11'h6cb;
  assign sel_513039 = $signed({1'h0, add_512951, array_index_512819[0]}) < $signed(13'h0fff) ? {add_512951, array_index_512819[0]} : 12'hfff;
  assign add_513041 = array_index_512880[11:1] + 11'h75d;
  assign sel_513043 = $signed({1'h0, add_512953, array_index_512834[0]}) < $signed({1'h0, sel_512955}) ? {add_512953, array_index_512834[0]} : sel_512955;
  assign add_513045 = array_index_512883[11:1] + 11'h75d;
  assign sel_513047 = $signed({1'h0, add_512957, array_index_512837[0]}) < $signed({1'h0, sel_512959}) ? {add_512957, array_index_512837[0]} : sel_512959;
  assign add_513049 = array_index_512942[11:1] + 11'h24f;
  assign sel_513052 = $signed({1'h0, add_512961, array_index_512880[0]}) < $signed({1'h0, sel_512964}) ? {add_512961, array_index_512880[0]} : sel_512964;
  assign add_513054 = array_index_512945[11:1] + 11'h24f;
  assign sel_513057 = $signed({1'h0, add_512966, array_index_512883[0]}) < $signed({1'h0, sel_512969}) ? {add_512966, array_index_512883[0]} : sel_512969;
  assign add_513082 = array_index_513022[11:0] + 12'h62b;
  assign sel_513084 = $signed({1'h0, add_512990}) < $signed({1'h0, sel_512992}) ? add_512990 : sel_512992;
  assign add_513087 = array_index_513025[11:0] + 12'h62b;
  assign sel_513089 = $signed({1'h0, add_512995}) < $signed({1'h0, sel_512997}) ? add_512995 : sel_512997;
  assign array_index_513120 = set1_unflattened[5'h05];
  assign array_index_513123 = set2_unflattened[5'h05];
  assign add_513127 = array_index_512818[11:4] + 8'h83;
  assign add_513130 = array_index_512819[11:4] + 8'h83;
  assign add_513133 = array_index_512834[11:0] + 12'ha09;
  assign sel_513135 = $signed({1'h0, add_513029}) < $signed(13'h0fff) ? add_513029 : 12'hfff;
  assign add_513137 = array_index_512837[11:0] + 12'ha09;
  assign sel_513139 = $signed({1'h0, add_513031}) < $signed(13'h0fff) ? add_513031 : 12'hfff;
  assign add_513141 = array_index_512880[11:1] + 11'h6cb;
  assign sel_513143 = $signed({1'h0, add_513033, array_index_512834[0]}) < $signed({1'h0, sel_513035}) ? {add_513033, array_index_512834[0]} : sel_513035;
  assign add_513145 = array_index_512883[11:1] + 11'h6cb;
  assign sel_513147 = $signed({1'h0, add_513037, array_index_512837[0]}) < $signed({1'h0, sel_513039}) ? {add_513037, array_index_512837[0]} : sel_513039;
  assign add_513149 = array_index_512942[11:1] + 11'h75d;
  assign sel_513151 = $signed({1'h0, add_513041, array_index_512880[0]}) < $signed({1'h0, sel_513043}) ? {add_513041, array_index_512880[0]} : sel_513043;
  assign add_513153 = array_index_512945[11:1] + 11'h75d;
  assign sel_513155 = $signed({1'h0, add_513045, array_index_512883[0]}) < $signed({1'h0, sel_513047}) ? {add_513045, array_index_512883[0]} : sel_513047;
  assign add_513157 = array_index_513022[11:1] + 11'h24f;
  assign sel_513160 = $signed({1'h0, add_513049, array_index_512942[0]}) < $signed({1'h0, sel_513052}) ? {add_513049, array_index_512942[0]} : sel_513052;
  assign add_513162 = array_index_513025[11:1] + 11'h24f;
  assign sel_513165 = $signed({1'h0, add_513054, array_index_512945[0]}) < $signed({1'h0, sel_513057}) ? {add_513054, array_index_512945[0]} : sel_513057;
  assign add_513194 = array_index_513120[11:0] + 12'h62b;
  assign sel_513196 = $signed({1'h0, add_513082}) < $signed({1'h0, sel_513084}) ? add_513082 : sel_513084;
  assign add_513199 = array_index_513123[11:0] + 12'h62b;
  assign sel_513201 = $signed({1'h0, add_513087}) < $signed({1'h0, sel_513089}) ? add_513087 : sel_513089;
  assign array_index_513238 = set1_unflattened[5'h06];
  assign array_index_513241 = set2_unflattened[5'h06];
  assign add_513245 = array_index_512818[11:0] + 12'h8e1;
  assign add_513247 = array_index_512819[11:0] + 12'h8e1;
  assign add_513249 = array_index_512834[11:4] + 8'h83;
  assign sel_513252 = $signed({1'h0, add_513127, array_index_512818[3:0]}) < $signed(13'h0fff) ? {add_513127, array_index_512818[3:0]} : 12'hfff;
  assign add_513254 = array_index_512837[11:4] + 8'h83;
  assign sel_513257 = $signed({1'h0, add_513130, array_index_512819[3:0]}) < $signed(13'h0fff) ? {add_513130, array_index_512819[3:0]} : 12'hfff;
  assign add_513259 = array_index_512880[11:0] + 12'ha09;
  assign sel_513261 = $signed({1'h0, add_513133}) < $signed({1'h0, sel_513135}) ? add_513133 : sel_513135;
  assign add_513263 = array_index_512883[11:0] + 12'ha09;
  assign sel_513265 = $signed({1'h0, add_513137}) < $signed({1'h0, sel_513139}) ? add_513137 : sel_513139;
  assign add_513267 = array_index_512942[11:1] + 11'h6cb;
  assign sel_513269 = $signed({1'h0, add_513141, array_index_512880[0]}) < $signed({1'h0, sel_513143}) ? {add_513141, array_index_512880[0]} : sel_513143;
  assign add_513271 = array_index_512945[11:1] + 11'h6cb;
  assign sel_513273 = $signed({1'h0, add_513145, array_index_512883[0]}) < $signed({1'h0, sel_513147}) ? {add_513145, array_index_512883[0]} : sel_513147;
  assign add_513275 = array_index_513022[11:1] + 11'h75d;
  assign sel_513277 = $signed({1'h0, add_513149, array_index_512942[0]}) < $signed({1'h0, sel_513151}) ? {add_513149, array_index_512942[0]} : sel_513151;
  assign add_513279 = array_index_513025[11:1] + 11'h75d;
  assign sel_513281 = $signed({1'h0, add_513153, array_index_512945[0]}) < $signed({1'h0, sel_513155}) ? {add_513153, array_index_512945[0]} : sel_513155;
  assign add_513283 = array_index_513120[11:1] + 11'h24f;
  assign sel_513286 = $signed({1'h0, add_513157, array_index_513022[0]}) < $signed({1'h0, sel_513160}) ? {add_513157, array_index_513022[0]} : sel_513160;
  assign add_513288 = array_index_513123[11:1] + 11'h24f;
  assign sel_513291 = $signed({1'h0, add_513162, array_index_513025[0]}) < $signed({1'h0, sel_513165}) ? {add_513162, array_index_513025[0]} : sel_513165;
  assign add_513324 = array_index_513238[11:0] + 12'h62b;
  assign sel_513326 = $signed({1'h0, add_513194}) < $signed({1'h0, sel_513196}) ? add_513194 : sel_513196;
  assign add_513329 = array_index_513241[11:0] + 12'h62b;
  assign sel_513331 = $signed({1'h0, add_513199}) < $signed({1'h0, sel_513201}) ? add_513199 : sel_513201;
  assign array_index_513374 = set1_unflattened[5'h07];
  assign array_index_513377 = set2_unflattened[5'h07];
  assign add_513381 = array_index_512818[11:2] + 10'h2bb;
  assign add_513384 = array_index_512819[11:2] + 10'h2bb;
  assign add_513387 = array_index_512834[11:0] + 12'h8e1;
  assign sel_513389 = $signed({1'h0, add_513245}) < $signed(13'h0fff) ? add_513245 : 12'hfff;
  assign add_513391 = array_index_512837[11:0] + 12'h8e1;
  assign sel_513393 = $signed({1'h0, add_513247}) < $signed(13'h0fff) ? add_513247 : 12'hfff;
  assign add_513395 = array_index_512880[11:4] + 8'h83;
  assign sel_513398 = $signed({1'h0, add_513249, array_index_512834[3:0]}) < $signed({1'h0, sel_513252}) ? {add_513249, array_index_512834[3:0]} : sel_513252;
  assign add_513400 = array_index_512883[11:4] + 8'h83;
  assign sel_513403 = $signed({1'h0, add_513254, array_index_512837[3:0]}) < $signed({1'h0, sel_513257}) ? {add_513254, array_index_512837[3:0]} : sel_513257;
  assign add_513405 = array_index_512942[11:0] + 12'ha09;
  assign sel_513407 = $signed({1'h0, add_513259}) < $signed({1'h0, sel_513261}) ? add_513259 : sel_513261;
  assign add_513409 = array_index_512945[11:0] + 12'ha09;
  assign sel_513411 = $signed({1'h0, add_513263}) < $signed({1'h0, sel_513265}) ? add_513263 : sel_513265;
  assign add_513413 = array_index_513022[11:1] + 11'h6cb;
  assign sel_513415 = $signed({1'h0, add_513267, array_index_512942[0]}) < $signed({1'h0, sel_513269}) ? {add_513267, array_index_512942[0]} : sel_513269;
  assign add_513417 = array_index_513025[11:1] + 11'h6cb;
  assign sel_513419 = $signed({1'h0, add_513271, array_index_512945[0]}) < $signed({1'h0, sel_513273}) ? {add_513271, array_index_512945[0]} : sel_513273;
  assign add_513421 = array_index_513120[11:1] + 11'h75d;
  assign sel_513423 = $signed({1'h0, add_513275, array_index_513022[0]}) < $signed({1'h0, sel_513277}) ? {add_513275, array_index_513022[0]} : sel_513277;
  assign add_513425 = array_index_513123[11:1] + 11'h75d;
  assign sel_513427 = $signed({1'h0, add_513279, array_index_513025[0]}) < $signed({1'h0, sel_513281}) ? {add_513279, array_index_513025[0]} : sel_513281;
  assign add_513429 = array_index_513238[11:1] + 11'h24f;
  assign sel_513432 = $signed({1'h0, add_513283, array_index_513120[0]}) < $signed({1'h0, sel_513286}) ? {add_513283, array_index_513120[0]} : sel_513286;
  assign add_513434 = array_index_513241[11:1] + 11'h24f;
  assign sel_513437 = $signed({1'h0, add_513288, array_index_513123[0]}) < $signed({1'h0, sel_513291}) ? {add_513288, array_index_513123[0]} : sel_513291;
  assign add_513474 = array_index_513374[11:0] + 12'h62b;
  assign sel_513476 = $signed({1'h0, add_513324}) < $signed({1'h0, sel_513326}) ? add_513324 : sel_513326;
  assign add_513479 = array_index_513377[11:0] + 12'h62b;
  assign sel_513481 = $signed({1'h0, add_513329}) < $signed({1'h0, sel_513331}) ? add_513329 : sel_513331;
  assign array_index_513530 = set1_unflattened[5'h08];
  assign array_index_513533 = set2_unflattened[5'h08];
  assign add_513537 = array_index_512818[11:0] + 12'h97d;
  assign add_513539 = array_index_512819[11:0] + 12'h97d;
  assign add_513541 = array_index_512834[11:2] + 10'h2bb;
  assign sel_513544 = $signed({1'h0, add_513381, array_index_512818[1:0]}) < $signed(13'h0fff) ? {add_513381, array_index_512818[1:0]} : 12'hfff;
  assign add_513546 = array_index_512837[11:2] + 10'h2bb;
  assign sel_513549 = $signed({1'h0, add_513384, array_index_512819[1:0]}) < $signed(13'h0fff) ? {add_513384, array_index_512819[1:0]} : 12'hfff;
  assign add_513551 = array_index_512880[11:0] + 12'h8e1;
  assign sel_513553 = $signed({1'h0, add_513387}) < $signed({1'h0, sel_513389}) ? add_513387 : sel_513389;
  assign add_513555 = array_index_512883[11:0] + 12'h8e1;
  assign sel_513557 = $signed({1'h0, add_513391}) < $signed({1'h0, sel_513393}) ? add_513391 : sel_513393;
  assign add_513559 = array_index_512942[11:4] + 8'h83;
  assign sel_513562 = $signed({1'h0, add_513395, array_index_512880[3:0]}) < $signed({1'h0, sel_513398}) ? {add_513395, array_index_512880[3:0]} : sel_513398;
  assign add_513564 = array_index_512945[11:4] + 8'h83;
  assign sel_513567 = $signed({1'h0, add_513400, array_index_512883[3:0]}) < $signed({1'h0, sel_513403}) ? {add_513400, array_index_512883[3:0]} : sel_513403;
  assign add_513569 = array_index_513022[11:0] + 12'ha09;
  assign sel_513571 = $signed({1'h0, add_513405}) < $signed({1'h0, sel_513407}) ? add_513405 : sel_513407;
  assign add_513573 = array_index_513025[11:0] + 12'ha09;
  assign sel_513575 = $signed({1'h0, add_513409}) < $signed({1'h0, sel_513411}) ? add_513409 : sel_513411;
  assign add_513577 = array_index_513120[11:1] + 11'h6cb;
  assign sel_513579 = $signed({1'h0, add_513413, array_index_513022[0]}) < $signed({1'h0, sel_513415}) ? {add_513413, array_index_513022[0]} : sel_513415;
  assign add_513581 = array_index_513123[11:1] + 11'h6cb;
  assign sel_513583 = $signed({1'h0, add_513417, array_index_513025[0]}) < $signed({1'h0, sel_513419}) ? {add_513417, array_index_513025[0]} : sel_513419;
  assign add_513585 = array_index_513238[11:1] + 11'h75d;
  assign sel_513587 = $signed({1'h0, add_513421, array_index_513120[0]}) < $signed({1'h0, sel_513423}) ? {add_513421, array_index_513120[0]} : sel_513423;
  assign add_513589 = array_index_513241[11:1] + 11'h75d;
  assign sel_513591 = $signed({1'h0, add_513425, array_index_513123[0]}) < $signed({1'h0, sel_513427}) ? {add_513425, array_index_513123[0]} : sel_513427;
  assign add_513593 = array_index_513374[11:1] + 11'h24f;
  assign sel_513596 = $signed({1'h0, add_513429, array_index_513238[0]}) < $signed({1'h0, sel_513432}) ? {add_513429, array_index_513238[0]} : sel_513432;
  assign add_513598 = array_index_513377[11:1] + 11'h24f;
  assign sel_513601 = $signed({1'h0, add_513434, array_index_513241[0]}) < $signed({1'h0, sel_513437}) ? {add_513434, array_index_513241[0]} : sel_513437;
  assign add_513642 = array_index_513530[11:0] + 12'h62b;
  assign sel_513644 = $signed({1'h0, add_513474}) < $signed({1'h0, sel_513476}) ? add_513474 : sel_513476;
  assign add_513647 = array_index_513533[11:0] + 12'h62b;
  assign sel_513649 = $signed({1'h0, add_513479}) < $signed({1'h0, sel_513481}) ? add_513479 : sel_513481;
  assign array_index_513702 = set1_unflattened[5'h09];
  assign array_index_513705 = set2_unflattened[5'h09];
  assign add_513709 = array_index_512818[11:0] + 12'hfe9;
  assign add_513711 = array_index_512819[11:0] + 12'hfe9;
  assign add_513713 = array_index_512834[11:0] + 12'h97d;
  assign sel_513715 = $signed({1'h0, add_513537}) < $signed(13'h0fff) ? add_513537 : 12'hfff;
  assign add_513717 = array_index_512837[11:0] + 12'h97d;
  assign sel_513719 = $signed({1'h0, add_513539}) < $signed(13'h0fff) ? add_513539 : 12'hfff;
  assign add_513721 = array_index_512880[11:2] + 10'h2bb;
  assign sel_513724 = $signed({1'h0, add_513541, array_index_512834[1:0]}) < $signed({1'h0, sel_513544}) ? {add_513541, array_index_512834[1:0]} : sel_513544;
  assign add_513726 = array_index_512883[11:2] + 10'h2bb;
  assign sel_513729 = $signed({1'h0, add_513546, array_index_512837[1:0]}) < $signed({1'h0, sel_513549}) ? {add_513546, array_index_512837[1:0]} : sel_513549;
  assign add_513731 = array_index_512942[11:0] + 12'h8e1;
  assign sel_513733 = $signed({1'h0, add_513551}) < $signed({1'h0, sel_513553}) ? add_513551 : sel_513553;
  assign add_513735 = array_index_512945[11:0] + 12'h8e1;
  assign sel_513737 = $signed({1'h0, add_513555}) < $signed({1'h0, sel_513557}) ? add_513555 : sel_513557;
  assign add_513739 = array_index_513022[11:4] + 8'h83;
  assign sel_513742 = $signed({1'h0, add_513559, array_index_512942[3:0]}) < $signed({1'h0, sel_513562}) ? {add_513559, array_index_512942[3:0]} : sel_513562;
  assign add_513744 = array_index_513025[11:4] + 8'h83;
  assign sel_513747 = $signed({1'h0, add_513564, array_index_512945[3:0]}) < $signed({1'h0, sel_513567}) ? {add_513564, array_index_512945[3:0]} : sel_513567;
  assign add_513749 = array_index_513120[11:0] + 12'ha09;
  assign sel_513751 = $signed({1'h0, add_513569}) < $signed({1'h0, sel_513571}) ? add_513569 : sel_513571;
  assign add_513753 = array_index_513123[11:0] + 12'ha09;
  assign sel_513755 = $signed({1'h0, add_513573}) < $signed({1'h0, sel_513575}) ? add_513573 : sel_513575;
  assign add_513757 = array_index_513238[11:1] + 11'h6cb;
  assign sel_513759 = $signed({1'h0, add_513577, array_index_513120[0]}) < $signed({1'h0, sel_513579}) ? {add_513577, array_index_513120[0]} : sel_513579;
  assign add_513761 = array_index_513241[11:1] + 11'h6cb;
  assign sel_513763 = $signed({1'h0, add_513581, array_index_513123[0]}) < $signed({1'h0, sel_513583}) ? {add_513581, array_index_513123[0]} : sel_513583;
  assign add_513765 = array_index_513374[11:1] + 11'h75d;
  assign sel_513767 = $signed({1'h0, add_513585, array_index_513238[0]}) < $signed({1'h0, sel_513587}) ? {add_513585, array_index_513238[0]} : sel_513587;
  assign add_513769 = array_index_513377[11:1] + 11'h75d;
  assign sel_513771 = $signed({1'h0, add_513589, array_index_513241[0]}) < $signed({1'h0, sel_513591}) ? {add_513589, array_index_513241[0]} : sel_513591;
  assign add_513773 = array_index_513530[11:1] + 11'h24f;
  assign sel_513776 = $signed({1'h0, add_513593, array_index_513374[0]}) < $signed({1'h0, sel_513596}) ? {add_513593, array_index_513374[0]} : sel_513596;
  assign add_513778 = array_index_513533[11:1] + 11'h24f;
  assign sel_513781 = $signed({1'h0, add_513598, array_index_513377[0]}) < $signed({1'h0, sel_513601}) ? {add_513598, array_index_513377[0]} : sel_513601;
  assign add_513826 = array_index_513702[11:0] + 12'h62b;
  assign sel_513828 = $signed({1'h0, add_513642}) < $signed({1'h0, sel_513644}) ? add_513642 : sel_513644;
  assign add_513831 = array_index_513705[11:0] + 12'h62b;
  assign sel_513833 = $signed({1'h0, add_513647}) < $signed({1'h0, sel_513649}) ? add_513647 : sel_513649;
  assign array_index_513890 = set1_unflattened[5'h0a];
  assign array_index_513893 = set2_unflattened[5'h0a];
  assign add_513897 = array_index_512818[11:1] + 11'h4cb;
  assign add_513899 = array_index_512819[11:1] + 11'h4cb;
  assign add_513901 = array_index_512834[11:0] + 12'hfe9;
  assign sel_513903 = $signed({1'h0, add_513709}) < $signed(13'h0fff) ? add_513709 : 12'hfff;
  assign add_513905 = array_index_512837[11:0] + 12'hfe9;
  assign sel_513907 = $signed({1'h0, add_513711}) < $signed(13'h0fff) ? add_513711 : 12'hfff;
  assign add_513909 = array_index_512880[11:0] + 12'h97d;
  assign sel_513911 = $signed({1'h0, add_513713}) < $signed({1'h0, sel_513715}) ? add_513713 : sel_513715;
  assign add_513913 = array_index_512883[11:0] + 12'h97d;
  assign sel_513915 = $signed({1'h0, add_513717}) < $signed({1'h0, sel_513719}) ? add_513717 : sel_513719;
  assign add_513917 = array_index_512942[11:2] + 10'h2bb;
  assign sel_513920 = $signed({1'h0, add_513721, array_index_512880[1:0]}) < $signed({1'h0, sel_513724}) ? {add_513721, array_index_512880[1:0]} : sel_513724;
  assign add_513922 = array_index_512945[11:2] + 10'h2bb;
  assign sel_513925 = $signed({1'h0, add_513726, array_index_512883[1:0]}) < $signed({1'h0, sel_513729}) ? {add_513726, array_index_512883[1:0]} : sel_513729;
  assign add_513927 = array_index_513022[11:0] + 12'h8e1;
  assign sel_513929 = $signed({1'h0, add_513731}) < $signed({1'h0, sel_513733}) ? add_513731 : sel_513733;
  assign add_513931 = array_index_513025[11:0] + 12'h8e1;
  assign sel_513933 = $signed({1'h0, add_513735}) < $signed({1'h0, sel_513737}) ? add_513735 : sel_513737;
  assign add_513935 = array_index_513120[11:4] + 8'h83;
  assign sel_513938 = $signed({1'h0, add_513739, array_index_513022[3:0]}) < $signed({1'h0, sel_513742}) ? {add_513739, array_index_513022[3:0]} : sel_513742;
  assign add_513940 = array_index_513123[11:4] + 8'h83;
  assign sel_513943 = $signed({1'h0, add_513744, array_index_513025[3:0]}) < $signed({1'h0, sel_513747}) ? {add_513744, array_index_513025[3:0]} : sel_513747;
  assign add_513945 = array_index_513238[11:0] + 12'ha09;
  assign sel_513947 = $signed({1'h0, add_513749}) < $signed({1'h0, sel_513751}) ? add_513749 : sel_513751;
  assign add_513949 = array_index_513241[11:0] + 12'ha09;
  assign sel_513951 = $signed({1'h0, add_513753}) < $signed({1'h0, sel_513755}) ? add_513753 : sel_513755;
  assign add_513953 = array_index_513374[11:1] + 11'h6cb;
  assign sel_513955 = $signed({1'h0, add_513757, array_index_513238[0]}) < $signed({1'h0, sel_513759}) ? {add_513757, array_index_513238[0]} : sel_513759;
  assign add_513957 = array_index_513377[11:1] + 11'h6cb;
  assign sel_513959 = $signed({1'h0, add_513761, array_index_513241[0]}) < $signed({1'h0, sel_513763}) ? {add_513761, array_index_513241[0]} : sel_513763;
  assign add_513961 = array_index_513530[11:1] + 11'h75d;
  assign sel_513963 = $signed({1'h0, add_513765, array_index_513374[0]}) < $signed({1'h0, sel_513767}) ? {add_513765, array_index_513374[0]} : sel_513767;
  assign add_513965 = array_index_513533[11:1] + 11'h75d;
  assign sel_513967 = $signed({1'h0, add_513769, array_index_513377[0]}) < $signed({1'h0, sel_513771}) ? {add_513769, array_index_513377[0]} : sel_513771;
  assign add_513969 = array_index_513702[11:1] + 11'h24f;
  assign sel_513972 = $signed({1'h0, add_513773, array_index_513530[0]}) < $signed({1'h0, sel_513776}) ? {add_513773, array_index_513530[0]} : sel_513776;
  assign add_513974 = array_index_513705[11:1] + 11'h24f;
  assign sel_513977 = $signed({1'h0, add_513778, array_index_513533[0]}) < $signed({1'h0, sel_513781}) ? {add_513778, array_index_513533[0]} : sel_513781;
  assign add_514026 = array_index_513890[11:0] + 12'h62b;
  assign sel_514028 = $signed({1'h0, add_513826}) < $signed({1'h0, sel_513828}) ? add_513826 : sel_513828;
  assign add_514031 = array_index_513893[11:0] + 12'h62b;
  assign sel_514033 = $signed({1'h0, add_513831}) < $signed({1'h0, sel_513833}) ? add_513831 : sel_513833;
  assign array_index_514096 = set1_unflattened[5'h0b];
  assign array_index_514099 = set2_unflattened[5'h0b];
  assign add_514103 = array_index_512818[11:0] + 12'h0a7;
  assign add_514105 = array_index_512819[11:0] + 12'h0a7;
  assign add_514107 = array_index_512834[11:1] + 11'h4cb;
  assign sel_514109 = $signed({1'h0, add_513897, array_index_512818[0]}) < $signed(13'h0fff) ? {add_513897, array_index_512818[0]} : 12'hfff;
  assign add_514111 = array_index_512837[11:1] + 11'h4cb;
  assign sel_514113 = $signed({1'h0, add_513899, array_index_512819[0]}) < $signed(13'h0fff) ? {add_513899, array_index_512819[0]} : 12'hfff;
  assign add_514115 = array_index_512880[11:0] + 12'hfe9;
  assign sel_514117 = $signed({1'h0, add_513901}) < $signed({1'h0, sel_513903}) ? add_513901 : sel_513903;
  assign add_514119 = array_index_512883[11:0] + 12'hfe9;
  assign sel_514121 = $signed({1'h0, add_513905}) < $signed({1'h0, sel_513907}) ? add_513905 : sel_513907;
  assign add_514123 = array_index_512942[11:0] + 12'h97d;
  assign sel_514125 = $signed({1'h0, add_513909}) < $signed({1'h0, sel_513911}) ? add_513909 : sel_513911;
  assign add_514127 = array_index_512945[11:0] + 12'h97d;
  assign sel_514129 = $signed({1'h0, add_513913}) < $signed({1'h0, sel_513915}) ? add_513913 : sel_513915;
  assign add_514131 = array_index_513022[11:2] + 10'h2bb;
  assign sel_514134 = $signed({1'h0, add_513917, array_index_512942[1:0]}) < $signed({1'h0, sel_513920}) ? {add_513917, array_index_512942[1:0]} : sel_513920;
  assign add_514136 = array_index_513025[11:2] + 10'h2bb;
  assign sel_514139 = $signed({1'h0, add_513922, array_index_512945[1:0]}) < $signed({1'h0, sel_513925}) ? {add_513922, array_index_512945[1:0]} : sel_513925;
  assign add_514141 = array_index_513120[11:0] + 12'h8e1;
  assign sel_514143 = $signed({1'h0, add_513927}) < $signed({1'h0, sel_513929}) ? add_513927 : sel_513929;
  assign add_514145 = array_index_513123[11:0] + 12'h8e1;
  assign sel_514147 = $signed({1'h0, add_513931}) < $signed({1'h0, sel_513933}) ? add_513931 : sel_513933;
  assign add_514149 = array_index_513238[11:4] + 8'h83;
  assign sel_514152 = $signed({1'h0, add_513935, array_index_513120[3:0]}) < $signed({1'h0, sel_513938}) ? {add_513935, array_index_513120[3:0]} : sel_513938;
  assign add_514154 = array_index_513241[11:4] + 8'h83;
  assign sel_514157 = $signed({1'h0, add_513940, array_index_513123[3:0]}) < $signed({1'h0, sel_513943}) ? {add_513940, array_index_513123[3:0]} : sel_513943;
  assign add_514159 = array_index_513374[11:0] + 12'ha09;
  assign sel_514161 = $signed({1'h0, add_513945}) < $signed({1'h0, sel_513947}) ? add_513945 : sel_513947;
  assign add_514163 = array_index_513377[11:0] + 12'ha09;
  assign sel_514165 = $signed({1'h0, add_513949}) < $signed({1'h0, sel_513951}) ? add_513949 : sel_513951;
  assign add_514167 = array_index_513530[11:1] + 11'h6cb;
  assign sel_514169 = $signed({1'h0, add_513953, array_index_513374[0]}) < $signed({1'h0, sel_513955}) ? {add_513953, array_index_513374[0]} : sel_513955;
  assign add_514171 = array_index_513533[11:1] + 11'h6cb;
  assign sel_514173 = $signed({1'h0, add_513957, array_index_513377[0]}) < $signed({1'h0, sel_513959}) ? {add_513957, array_index_513377[0]} : sel_513959;
  assign add_514175 = array_index_513702[11:1] + 11'h75d;
  assign sel_514177 = $signed({1'h0, add_513961, array_index_513530[0]}) < $signed({1'h0, sel_513963}) ? {add_513961, array_index_513530[0]} : sel_513963;
  assign add_514179 = array_index_513705[11:1] + 11'h75d;
  assign sel_514181 = $signed({1'h0, add_513965, array_index_513533[0]}) < $signed({1'h0, sel_513967}) ? {add_513965, array_index_513533[0]} : sel_513967;
  assign add_514183 = array_index_513890[11:1] + 11'h24f;
  assign sel_514186 = $signed({1'h0, add_513969, array_index_513702[0]}) < $signed({1'h0, sel_513972}) ? {add_513969, array_index_513702[0]} : sel_513972;
  assign add_514188 = array_index_513893[11:1] + 11'h24f;
  assign sel_514191 = $signed({1'h0, add_513974, array_index_513705[0]}) < $signed({1'h0, sel_513977}) ? {add_513974, array_index_513705[0]} : sel_513977;
  assign add_514244 = array_index_514096[11:0] + 12'h62b;
  assign sel_514246 = $signed({1'h0, add_514026}) < $signed({1'h0, sel_514028}) ? add_514026 : sel_514028;
  assign add_514249 = array_index_514099[11:0] + 12'h62b;
  assign sel_514251 = $signed({1'h0, add_514031}) < $signed({1'h0, sel_514033}) ? add_514031 : sel_514033;
  assign array_index_514318 = set1_unflattened[5'h0c];
  assign array_index_514321 = set2_unflattened[5'h0c];
  assign add_514325 = array_index_512818[11:2] + 10'h353;
  assign add_514327 = array_index_512819[11:2] + 10'h353;
  assign add_514329 = array_index_512834[11:0] + 12'h0a7;
  assign sel_514331 = $signed({1'h0, add_514103}) < $signed(13'h0fff) ? add_514103 : 12'hfff;
  assign add_514333 = array_index_512837[11:0] + 12'h0a7;
  assign sel_514335 = $signed({1'h0, add_514105}) < $signed(13'h0fff) ? add_514105 : 12'hfff;
  assign add_514337 = array_index_512880[11:1] + 11'h4cb;
  assign sel_514339 = $signed({1'h0, add_514107, array_index_512834[0]}) < $signed({1'h0, sel_514109}) ? {add_514107, array_index_512834[0]} : sel_514109;
  assign add_514341 = array_index_512883[11:1] + 11'h4cb;
  assign sel_514343 = $signed({1'h0, add_514111, array_index_512837[0]}) < $signed({1'h0, sel_514113}) ? {add_514111, array_index_512837[0]} : sel_514113;
  assign add_514345 = array_index_512942[11:0] + 12'hfe9;
  assign sel_514347 = $signed({1'h0, add_514115}) < $signed({1'h0, sel_514117}) ? add_514115 : sel_514117;
  assign add_514349 = array_index_512945[11:0] + 12'hfe9;
  assign sel_514351 = $signed({1'h0, add_514119}) < $signed({1'h0, sel_514121}) ? add_514119 : sel_514121;
  assign add_514353 = array_index_513022[11:0] + 12'h97d;
  assign sel_514355 = $signed({1'h0, add_514123}) < $signed({1'h0, sel_514125}) ? add_514123 : sel_514125;
  assign add_514357 = array_index_513025[11:0] + 12'h97d;
  assign sel_514359 = $signed({1'h0, add_514127}) < $signed({1'h0, sel_514129}) ? add_514127 : sel_514129;
  assign add_514361 = array_index_513120[11:2] + 10'h2bb;
  assign sel_514364 = $signed({1'h0, add_514131, array_index_513022[1:0]}) < $signed({1'h0, sel_514134}) ? {add_514131, array_index_513022[1:0]} : sel_514134;
  assign add_514366 = array_index_513123[11:2] + 10'h2bb;
  assign sel_514369 = $signed({1'h0, add_514136, array_index_513025[1:0]}) < $signed({1'h0, sel_514139}) ? {add_514136, array_index_513025[1:0]} : sel_514139;
  assign add_514371 = array_index_513238[11:0] + 12'h8e1;
  assign sel_514373 = $signed({1'h0, add_514141}) < $signed({1'h0, sel_514143}) ? add_514141 : sel_514143;
  assign add_514375 = array_index_513241[11:0] + 12'h8e1;
  assign sel_514377 = $signed({1'h0, add_514145}) < $signed({1'h0, sel_514147}) ? add_514145 : sel_514147;
  assign add_514379 = array_index_513374[11:4] + 8'h83;
  assign sel_514382 = $signed({1'h0, add_514149, array_index_513238[3:0]}) < $signed({1'h0, sel_514152}) ? {add_514149, array_index_513238[3:0]} : sel_514152;
  assign add_514384 = array_index_513377[11:4] + 8'h83;
  assign sel_514387 = $signed({1'h0, add_514154, array_index_513241[3:0]}) < $signed({1'h0, sel_514157}) ? {add_514154, array_index_513241[3:0]} : sel_514157;
  assign add_514389 = array_index_513530[11:0] + 12'ha09;
  assign sel_514391 = $signed({1'h0, add_514159}) < $signed({1'h0, sel_514161}) ? add_514159 : sel_514161;
  assign add_514393 = array_index_513533[11:0] + 12'ha09;
  assign sel_514395 = $signed({1'h0, add_514163}) < $signed({1'h0, sel_514165}) ? add_514163 : sel_514165;
  assign add_514397 = array_index_513702[11:1] + 11'h6cb;
  assign sel_514399 = $signed({1'h0, add_514167, array_index_513530[0]}) < $signed({1'h0, sel_514169}) ? {add_514167, array_index_513530[0]} : sel_514169;
  assign add_514401 = array_index_513705[11:1] + 11'h6cb;
  assign sel_514403 = $signed({1'h0, add_514171, array_index_513533[0]}) < $signed({1'h0, sel_514173}) ? {add_514171, array_index_513533[0]} : sel_514173;
  assign add_514405 = array_index_513890[11:1] + 11'h75d;
  assign sel_514407 = $signed({1'h0, add_514175, array_index_513702[0]}) < $signed({1'h0, sel_514177}) ? {add_514175, array_index_513702[0]} : sel_514177;
  assign add_514409 = array_index_513893[11:1] + 11'h75d;
  assign sel_514411 = $signed({1'h0, add_514179, array_index_513705[0]}) < $signed({1'h0, sel_514181}) ? {add_514179, array_index_513705[0]} : sel_514181;
  assign add_514413 = array_index_514096[11:1] + 11'h24f;
  assign sel_514416 = $signed({1'h0, add_514183, array_index_513890[0]}) < $signed({1'h0, sel_514186}) ? {add_514183, array_index_513890[0]} : sel_514186;
  assign add_514418 = array_index_514099[11:1] + 11'h24f;
  assign sel_514421 = $signed({1'h0, add_514188, array_index_513893[0]}) < $signed({1'h0, sel_514191}) ? {add_514188, array_index_513893[0]} : sel_514191;
  assign add_514478 = array_index_514318[11:0] + 12'h62b;
  assign sel_514480 = $signed({1'h0, add_514244}) < $signed({1'h0, sel_514246}) ? add_514244 : sel_514246;
  assign add_514483 = array_index_514321[11:0] + 12'h62b;
  assign sel_514485 = $signed({1'h0, add_514249}) < $signed({1'h0, sel_514251}) ? add_514249 : sel_514251;
  assign array_index_514558 = set1_unflattened[5'h0d];
  assign array_index_514561 = set2_unflattened[5'h0d];
  assign add_514565 = array_index_512818[11:1] + 11'h2d5;
  assign add_514567 = array_index_512819[11:1] + 11'h2d5;
  assign add_514569 = array_index_512834[11:2] + 10'h353;
  assign sel_514571 = $signed({1'h0, add_514325, array_index_512818[1:0]}) < $signed(13'h0fff) ? {add_514325, array_index_512818[1:0]} : 12'hfff;
  assign add_514573 = array_index_512837[11:2] + 10'h353;
  assign sel_514575 = $signed({1'h0, add_514327, array_index_512819[1:0]}) < $signed(13'h0fff) ? {add_514327, array_index_512819[1:0]} : 12'hfff;
  assign add_514577 = array_index_512880[11:0] + 12'h0a7;
  assign sel_514579 = $signed({1'h0, add_514329}) < $signed({1'h0, sel_514331}) ? add_514329 : sel_514331;
  assign add_514581 = array_index_512883[11:0] + 12'h0a7;
  assign sel_514583 = $signed({1'h0, add_514333}) < $signed({1'h0, sel_514335}) ? add_514333 : sel_514335;
  assign add_514585 = array_index_512942[11:1] + 11'h4cb;
  assign sel_514587 = $signed({1'h0, add_514337, array_index_512880[0]}) < $signed({1'h0, sel_514339}) ? {add_514337, array_index_512880[0]} : sel_514339;
  assign add_514589 = array_index_512945[11:1] + 11'h4cb;
  assign sel_514591 = $signed({1'h0, add_514341, array_index_512883[0]}) < $signed({1'h0, sel_514343}) ? {add_514341, array_index_512883[0]} : sel_514343;
  assign add_514593 = array_index_513022[11:0] + 12'hfe9;
  assign sel_514595 = $signed({1'h0, add_514345}) < $signed({1'h0, sel_514347}) ? add_514345 : sel_514347;
  assign add_514597 = array_index_513025[11:0] + 12'hfe9;
  assign sel_514599 = $signed({1'h0, add_514349}) < $signed({1'h0, sel_514351}) ? add_514349 : sel_514351;
  assign add_514601 = array_index_513120[11:0] + 12'h97d;
  assign sel_514603 = $signed({1'h0, add_514353}) < $signed({1'h0, sel_514355}) ? add_514353 : sel_514355;
  assign add_514605 = array_index_513123[11:0] + 12'h97d;
  assign sel_514607 = $signed({1'h0, add_514357}) < $signed({1'h0, sel_514359}) ? add_514357 : sel_514359;
  assign add_514609 = array_index_513238[11:2] + 10'h2bb;
  assign sel_514612 = $signed({1'h0, add_514361, array_index_513120[1:0]}) < $signed({1'h0, sel_514364}) ? {add_514361, array_index_513120[1:0]} : sel_514364;
  assign add_514614 = array_index_513241[11:2] + 10'h2bb;
  assign sel_514617 = $signed({1'h0, add_514366, array_index_513123[1:0]}) < $signed({1'h0, sel_514369}) ? {add_514366, array_index_513123[1:0]} : sel_514369;
  assign add_514619 = array_index_513374[11:0] + 12'h8e1;
  assign sel_514621 = $signed({1'h0, add_514371}) < $signed({1'h0, sel_514373}) ? add_514371 : sel_514373;
  assign add_514623 = array_index_513377[11:0] + 12'h8e1;
  assign sel_514625 = $signed({1'h0, add_514375}) < $signed({1'h0, sel_514377}) ? add_514375 : sel_514377;
  assign add_514627 = array_index_513530[11:4] + 8'h83;
  assign sel_514630 = $signed({1'h0, add_514379, array_index_513374[3:0]}) < $signed({1'h0, sel_514382}) ? {add_514379, array_index_513374[3:0]} : sel_514382;
  assign add_514632 = array_index_513533[11:4] + 8'h83;
  assign sel_514635 = $signed({1'h0, add_514384, array_index_513377[3:0]}) < $signed({1'h0, sel_514387}) ? {add_514384, array_index_513377[3:0]} : sel_514387;
  assign add_514637 = array_index_513702[11:0] + 12'ha09;
  assign sel_514639 = $signed({1'h0, add_514389}) < $signed({1'h0, sel_514391}) ? add_514389 : sel_514391;
  assign add_514641 = array_index_513705[11:0] + 12'ha09;
  assign sel_514643 = $signed({1'h0, add_514393}) < $signed({1'h0, sel_514395}) ? add_514393 : sel_514395;
  assign add_514645 = array_index_513890[11:1] + 11'h6cb;
  assign sel_514647 = $signed({1'h0, add_514397, array_index_513702[0]}) < $signed({1'h0, sel_514399}) ? {add_514397, array_index_513702[0]} : sel_514399;
  assign add_514649 = array_index_513893[11:1] + 11'h6cb;
  assign sel_514651 = $signed({1'h0, add_514401, array_index_513705[0]}) < $signed({1'h0, sel_514403}) ? {add_514401, array_index_513705[0]} : sel_514403;
  assign add_514653 = array_index_514096[11:1] + 11'h75d;
  assign sel_514655 = $signed({1'h0, add_514405, array_index_513890[0]}) < $signed({1'h0, sel_514407}) ? {add_514405, array_index_513890[0]} : sel_514407;
  assign add_514657 = array_index_514099[11:1] + 11'h75d;
  assign sel_514659 = $signed({1'h0, add_514409, array_index_513893[0]}) < $signed({1'h0, sel_514411}) ? {add_514409, array_index_513893[0]} : sel_514411;
  assign add_514661 = array_index_514318[11:1] + 11'h24f;
  assign sel_514664 = $signed({1'h0, add_514413, array_index_514096[0]}) < $signed({1'h0, sel_514416}) ? {add_514413, array_index_514096[0]} : sel_514416;
  assign add_514666 = array_index_514321[11:1] + 11'h24f;
  assign sel_514669 = $signed({1'h0, add_514418, array_index_514099[0]}) < $signed({1'h0, sel_514421}) ? {add_514418, array_index_514099[0]} : sel_514421;
  assign add_514730 = array_index_514558[11:0] + 12'h62b;
  assign sel_514732 = $signed({1'h0, add_514478}) < $signed({1'h0, sel_514480}) ? add_514478 : sel_514480;
  assign add_514735 = array_index_514561[11:0] + 12'h62b;
  assign sel_514737 = $signed({1'h0, add_514483}) < $signed({1'h0, sel_514485}) ? add_514483 : sel_514485;
  assign array_index_514818 = set1_unflattened[5'h0e];
  assign array_index_514821 = set2_unflattened[5'h0e];
  assign add_514825 = array_index_512818[11:3] + 9'h1ef;
  assign add_514828 = array_index_512819[11:3] + 9'h1ef;
  assign add_514831 = array_index_512834[11:1] + 11'h2d5;
  assign sel_514833 = $signed({1'h0, add_514565, array_index_512818[0]}) < $signed(13'h0fff) ? {add_514565, array_index_512818[0]} : 12'hfff;
  assign add_514835 = array_index_512837[11:1] + 11'h2d5;
  assign sel_514837 = $signed({1'h0, add_514567, array_index_512819[0]}) < $signed(13'h0fff) ? {add_514567, array_index_512819[0]} : 12'hfff;
  assign add_514839 = array_index_512880[11:2] + 10'h353;
  assign sel_514841 = $signed({1'h0, add_514569, array_index_512834[1:0]}) < $signed({1'h0, sel_514571}) ? {add_514569, array_index_512834[1:0]} : sel_514571;
  assign add_514843 = array_index_512883[11:2] + 10'h353;
  assign sel_514845 = $signed({1'h0, add_514573, array_index_512837[1:0]}) < $signed({1'h0, sel_514575}) ? {add_514573, array_index_512837[1:0]} : sel_514575;
  assign add_514847 = array_index_512942[11:0] + 12'h0a7;
  assign sel_514849 = $signed({1'h0, add_514577}) < $signed({1'h0, sel_514579}) ? add_514577 : sel_514579;
  assign add_514851 = array_index_512945[11:0] + 12'h0a7;
  assign sel_514853 = $signed({1'h0, add_514581}) < $signed({1'h0, sel_514583}) ? add_514581 : sel_514583;
  assign add_514855 = array_index_513022[11:1] + 11'h4cb;
  assign sel_514857 = $signed({1'h0, add_514585, array_index_512942[0]}) < $signed({1'h0, sel_514587}) ? {add_514585, array_index_512942[0]} : sel_514587;
  assign add_514859 = array_index_513025[11:1] + 11'h4cb;
  assign sel_514861 = $signed({1'h0, add_514589, array_index_512945[0]}) < $signed({1'h0, sel_514591}) ? {add_514589, array_index_512945[0]} : sel_514591;
  assign add_514863 = array_index_513120[11:0] + 12'hfe9;
  assign sel_514865 = $signed({1'h0, add_514593}) < $signed({1'h0, sel_514595}) ? add_514593 : sel_514595;
  assign add_514867 = array_index_513123[11:0] + 12'hfe9;
  assign sel_514869 = $signed({1'h0, add_514597}) < $signed({1'h0, sel_514599}) ? add_514597 : sel_514599;
  assign add_514871 = array_index_513238[11:0] + 12'h97d;
  assign sel_514873 = $signed({1'h0, add_514601}) < $signed({1'h0, sel_514603}) ? add_514601 : sel_514603;
  assign add_514875 = array_index_513241[11:0] + 12'h97d;
  assign sel_514877 = $signed({1'h0, add_514605}) < $signed({1'h0, sel_514607}) ? add_514605 : sel_514607;
  assign add_514879 = array_index_513374[11:2] + 10'h2bb;
  assign sel_514882 = $signed({1'h0, add_514609, array_index_513238[1:0]}) < $signed({1'h0, sel_514612}) ? {add_514609, array_index_513238[1:0]} : sel_514612;
  assign add_514884 = array_index_513377[11:2] + 10'h2bb;
  assign sel_514887 = $signed({1'h0, add_514614, array_index_513241[1:0]}) < $signed({1'h0, sel_514617}) ? {add_514614, array_index_513241[1:0]} : sel_514617;
  assign add_514889 = array_index_513530[11:0] + 12'h8e1;
  assign sel_514891 = $signed({1'h0, add_514619}) < $signed({1'h0, sel_514621}) ? add_514619 : sel_514621;
  assign add_514893 = array_index_513533[11:0] + 12'h8e1;
  assign sel_514895 = $signed({1'h0, add_514623}) < $signed({1'h0, sel_514625}) ? add_514623 : sel_514625;
  assign add_514897 = array_index_513702[11:4] + 8'h83;
  assign sel_514900 = $signed({1'h0, add_514627, array_index_513530[3:0]}) < $signed({1'h0, sel_514630}) ? {add_514627, array_index_513530[3:0]} : sel_514630;
  assign add_514902 = array_index_513705[11:4] + 8'h83;
  assign sel_514905 = $signed({1'h0, add_514632, array_index_513533[3:0]}) < $signed({1'h0, sel_514635}) ? {add_514632, array_index_513533[3:0]} : sel_514635;
  assign add_514907 = array_index_513890[11:0] + 12'ha09;
  assign sel_514909 = $signed({1'h0, add_514637}) < $signed({1'h0, sel_514639}) ? add_514637 : sel_514639;
  assign add_514911 = array_index_513893[11:0] + 12'ha09;
  assign sel_514913 = $signed({1'h0, add_514641}) < $signed({1'h0, sel_514643}) ? add_514641 : sel_514643;
  assign add_514915 = array_index_514096[11:1] + 11'h6cb;
  assign sel_514917 = $signed({1'h0, add_514645, array_index_513890[0]}) < $signed({1'h0, sel_514647}) ? {add_514645, array_index_513890[0]} : sel_514647;
  assign add_514919 = array_index_514099[11:1] + 11'h6cb;
  assign sel_514921 = $signed({1'h0, add_514649, array_index_513893[0]}) < $signed({1'h0, sel_514651}) ? {add_514649, array_index_513893[0]} : sel_514651;
  assign add_514923 = array_index_514318[11:1] + 11'h75d;
  assign sel_514925 = $signed({1'h0, add_514653, array_index_514096[0]}) < $signed({1'h0, sel_514655}) ? {add_514653, array_index_514096[0]} : sel_514655;
  assign add_514927 = array_index_514321[11:1] + 11'h75d;
  assign sel_514929 = $signed({1'h0, add_514657, array_index_514099[0]}) < $signed({1'h0, sel_514659}) ? {add_514657, array_index_514099[0]} : sel_514659;
  assign add_514931 = array_index_514558[11:1] + 11'h24f;
  assign sel_514934 = $signed({1'h0, add_514661, array_index_514318[0]}) < $signed({1'h0, sel_514664}) ? {add_514661, array_index_514318[0]} : sel_514664;
  assign add_514936 = array_index_514561[11:1] + 11'h24f;
  assign sel_514939 = $signed({1'h0, add_514666, array_index_514321[0]}) < $signed({1'h0, sel_514669}) ? {add_514666, array_index_514321[0]} : sel_514669;
  assign add_515004 = array_index_514818[11:0] + 12'h62b;
  assign sel_515006 = $signed({1'h0, add_514730}) < $signed({1'h0, sel_514732}) ? add_514730 : sel_514732;
  assign add_515009 = array_index_514821[11:0] + 12'h62b;
  assign sel_515011 = $signed({1'h0, add_514735}) < $signed({1'h0, sel_514737}) ? add_514735 : sel_514737;
  assign array_index_515098 = set1_unflattened[5'h0f];
  assign array_index_515101 = set2_unflattened[5'h0f];
  assign add_515105 = array_index_512818[11:0] + 12'h067;
  assign add_515107 = array_index_512819[11:0] + 12'h067;
  assign add_515109 = array_index_512834[11:3] + 9'h1ef;
  assign sel_515112 = $signed({1'h0, add_514825, array_index_512818[2:0]}) < $signed(13'h0fff) ? {add_514825, array_index_512818[2:0]} : 12'hfff;
  assign add_515114 = array_index_512837[11:3] + 9'h1ef;
  assign sel_515117 = $signed({1'h0, add_514828, array_index_512819[2:0]}) < $signed(13'h0fff) ? {add_514828, array_index_512819[2:0]} : 12'hfff;
  assign add_515119 = array_index_512880[11:1] + 11'h2d5;
  assign sel_515121 = $signed({1'h0, add_514831, array_index_512834[0]}) < $signed({1'h0, sel_514833}) ? {add_514831, array_index_512834[0]} : sel_514833;
  assign add_515123 = array_index_512883[11:1] + 11'h2d5;
  assign sel_515125 = $signed({1'h0, add_514835, array_index_512837[0]}) < $signed({1'h0, sel_514837}) ? {add_514835, array_index_512837[0]} : sel_514837;
  assign add_515127 = array_index_512942[11:2] + 10'h353;
  assign sel_515129 = $signed({1'h0, add_514839, array_index_512880[1:0]}) < $signed({1'h0, sel_514841}) ? {add_514839, array_index_512880[1:0]} : sel_514841;
  assign add_515131 = array_index_512945[11:2] + 10'h353;
  assign sel_515133 = $signed({1'h0, add_514843, array_index_512883[1:0]}) < $signed({1'h0, sel_514845}) ? {add_514843, array_index_512883[1:0]} : sel_514845;
  assign add_515135 = array_index_513022[11:0] + 12'h0a7;
  assign sel_515137 = $signed({1'h0, add_514847}) < $signed({1'h0, sel_514849}) ? add_514847 : sel_514849;
  assign add_515139 = array_index_513025[11:0] + 12'h0a7;
  assign sel_515141 = $signed({1'h0, add_514851}) < $signed({1'h0, sel_514853}) ? add_514851 : sel_514853;
  assign add_515143 = array_index_513120[11:1] + 11'h4cb;
  assign sel_515145 = $signed({1'h0, add_514855, array_index_513022[0]}) < $signed({1'h0, sel_514857}) ? {add_514855, array_index_513022[0]} : sel_514857;
  assign add_515147 = array_index_513123[11:1] + 11'h4cb;
  assign sel_515149 = $signed({1'h0, add_514859, array_index_513025[0]}) < $signed({1'h0, sel_514861}) ? {add_514859, array_index_513025[0]} : sel_514861;
  assign add_515151 = array_index_513238[11:0] + 12'hfe9;
  assign sel_515153 = $signed({1'h0, add_514863}) < $signed({1'h0, sel_514865}) ? add_514863 : sel_514865;
  assign add_515155 = array_index_513241[11:0] + 12'hfe9;
  assign sel_515157 = $signed({1'h0, add_514867}) < $signed({1'h0, sel_514869}) ? add_514867 : sel_514869;
  assign add_515159 = array_index_513374[11:0] + 12'h97d;
  assign sel_515161 = $signed({1'h0, add_514871}) < $signed({1'h0, sel_514873}) ? add_514871 : sel_514873;
  assign add_515163 = array_index_513377[11:0] + 12'h97d;
  assign sel_515165 = $signed({1'h0, add_514875}) < $signed({1'h0, sel_514877}) ? add_514875 : sel_514877;
  assign add_515167 = array_index_513530[11:2] + 10'h2bb;
  assign sel_515170 = $signed({1'h0, add_514879, array_index_513374[1:0]}) < $signed({1'h0, sel_514882}) ? {add_514879, array_index_513374[1:0]} : sel_514882;
  assign add_515172 = array_index_513533[11:2] + 10'h2bb;
  assign sel_515175 = $signed({1'h0, add_514884, array_index_513377[1:0]}) < $signed({1'h0, sel_514887}) ? {add_514884, array_index_513377[1:0]} : sel_514887;
  assign add_515177 = array_index_513702[11:0] + 12'h8e1;
  assign sel_515179 = $signed({1'h0, add_514889}) < $signed({1'h0, sel_514891}) ? add_514889 : sel_514891;
  assign add_515181 = array_index_513705[11:0] + 12'h8e1;
  assign sel_515183 = $signed({1'h0, add_514893}) < $signed({1'h0, sel_514895}) ? add_514893 : sel_514895;
  assign add_515185 = array_index_513890[11:4] + 8'h83;
  assign sel_515188 = $signed({1'h0, add_514897, array_index_513702[3:0]}) < $signed({1'h0, sel_514900}) ? {add_514897, array_index_513702[3:0]} : sel_514900;
  assign add_515190 = array_index_513893[11:4] + 8'h83;
  assign sel_515193 = $signed({1'h0, add_514902, array_index_513705[3:0]}) < $signed({1'h0, sel_514905}) ? {add_514902, array_index_513705[3:0]} : sel_514905;
  assign add_515195 = array_index_514096[11:0] + 12'ha09;
  assign sel_515197 = $signed({1'h0, add_514907}) < $signed({1'h0, sel_514909}) ? add_514907 : sel_514909;
  assign add_515199 = array_index_514099[11:0] + 12'ha09;
  assign sel_515201 = $signed({1'h0, add_514911}) < $signed({1'h0, sel_514913}) ? add_514911 : sel_514913;
  assign add_515203 = array_index_514318[11:1] + 11'h6cb;
  assign sel_515205 = $signed({1'h0, add_514915, array_index_514096[0]}) < $signed({1'h0, sel_514917}) ? {add_514915, array_index_514096[0]} : sel_514917;
  assign add_515207 = array_index_514321[11:1] + 11'h6cb;
  assign sel_515209 = $signed({1'h0, add_514919, array_index_514099[0]}) < $signed({1'h0, sel_514921}) ? {add_514919, array_index_514099[0]} : sel_514921;
  assign add_515211 = array_index_514558[11:1] + 11'h75d;
  assign sel_515213 = $signed({1'h0, add_514923, array_index_514318[0]}) < $signed({1'h0, sel_514925}) ? {add_514923, array_index_514318[0]} : sel_514925;
  assign add_515215 = array_index_514561[11:1] + 11'h75d;
  assign sel_515217 = $signed({1'h0, add_514927, array_index_514321[0]}) < $signed({1'h0, sel_514929}) ? {add_514927, array_index_514321[0]} : sel_514929;
  assign add_515219 = array_index_514818[11:1] + 11'h24f;
  assign sel_515222 = $signed({1'h0, add_514931, array_index_514558[0]}) < $signed({1'h0, sel_514934}) ? {add_514931, array_index_514558[0]} : sel_514934;
  assign add_515224 = array_index_514821[11:1] + 11'h24f;
  assign sel_515227 = $signed({1'h0, add_514936, array_index_514561[0]}) < $signed({1'h0, sel_514939}) ? {add_514936, array_index_514561[0]} : sel_514939;
  assign add_515298 = array_index_515098[11:0] + 12'h62b;
  assign sel_515300 = $signed({1'h0, add_515004}) < $signed({1'h0, sel_515006}) ? add_515004 : sel_515006;
  assign add_515303 = array_index_515101[11:0] + 12'h62b;
  assign sel_515305 = $signed({1'h0, add_515009}) < $signed({1'h0, sel_515011}) ? add_515009 : sel_515011;
  assign add_515307 = array_index_512818[11:3] + 9'h0f5;
  assign add_515309 = array_index_512819[11:3] + 9'h0f5;
  assign array_index_515398 = set1_unflattened[5'h10];
  assign array_index_515401 = set2_unflattened[5'h10];
  assign add_515411 = array_index_512834[11:0] + 12'h067;
  assign sel_515413 = $signed({1'h0, add_515105}) < $signed(13'h0fff) ? add_515105 : 12'hfff;
  assign add_515415 = array_index_512837[11:0] + 12'h067;
  assign sel_515417 = $signed({1'h0, add_515107}) < $signed(13'h0fff) ? add_515107 : 12'hfff;
  assign add_515419 = array_index_512880[11:3] + 9'h1ef;
  assign sel_515422 = $signed({1'h0, add_515109, array_index_512834[2:0]}) < $signed({1'h0, sel_515112}) ? {add_515109, array_index_512834[2:0]} : sel_515112;
  assign add_515424 = array_index_512883[11:3] + 9'h1ef;
  assign sel_515427 = $signed({1'h0, add_515114, array_index_512837[2:0]}) < $signed({1'h0, sel_515117}) ? {add_515114, array_index_512837[2:0]} : sel_515117;
  assign add_515429 = array_index_512942[11:1] + 11'h2d5;
  assign sel_515431 = $signed({1'h0, add_515119, array_index_512880[0]}) < $signed({1'h0, sel_515121}) ? {add_515119, array_index_512880[0]} : sel_515121;
  assign add_515433 = array_index_512945[11:1] + 11'h2d5;
  assign sel_515435 = $signed({1'h0, add_515123, array_index_512883[0]}) < $signed({1'h0, sel_515125}) ? {add_515123, array_index_512883[0]} : sel_515125;
  assign add_515437 = array_index_513022[11:2] + 10'h353;
  assign sel_515439 = $signed({1'h0, add_515127, array_index_512942[1:0]}) < $signed({1'h0, sel_515129}) ? {add_515127, array_index_512942[1:0]} : sel_515129;
  assign add_515441 = array_index_513025[11:2] + 10'h353;
  assign sel_515443 = $signed({1'h0, add_515131, array_index_512945[1:0]}) < $signed({1'h0, sel_515133}) ? {add_515131, array_index_512945[1:0]} : sel_515133;
  assign add_515445 = array_index_513120[11:0] + 12'h0a7;
  assign sel_515447 = $signed({1'h0, add_515135}) < $signed({1'h0, sel_515137}) ? add_515135 : sel_515137;
  assign add_515449 = array_index_513123[11:0] + 12'h0a7;
  assign sel_515451 = $signed({1'h0, add_515139}) < $signed({1'h0, sel_515141}) ? add_515139 : sel_515141;
  assign add_515453 = array_index_513238[11:1] + 11'h4cb;
  assign sel_515455 = $signed({1'h0, add_515143, array_index_513120[0]}) < $signed({1'h0, sel_515145}) ? {add_515143, array_index_513120[0]} : sel_515145;
  assign add_515457 = array_index_513241[11:1] + 11'h4cb;
  assign sel_515459 = $signed({1'h0, add_515147, array_index_513123[0]}) < $signed({1'h0, sel_515149}) ? {add_515147, array_index_513123[0]} : sel_515149;
  assign add_515461 = array_index_513374[11:0] + 12'hfe9;
  assign sel_515463 = $signed({1'h0, add_515151}) < $signed({1'h0, sel_515153}) ? add_515151 : sel_515153;
  assign add_515465 = array_index_513377[11:0] + 12'hfe9;
  assign sel_515467 = $signed({1'h0, add_515155}) < $signed({1'h0, sel_515157}) ? add_515155 : sel_515157;
  assign add_515469 = array_index_513530[11:0] + 12'h97d;
  assign sel_515471 = $signed({1'h0, add_515159}) < $signed({1'h0, sel_515161}) ? add_515159 : sel_515161;
  assign add_515473 = array_index_513533[11:0] + 12'h97d;
  assign sel_515475 = $signed({1'h0, add_515163}) < $signed({1'h0, sel_515165}) ? add_515163 : sel_515165;
  assign add_515477 = array_index_513702[11:2] + 10'h2bb;
  assign sel_515480 = $signed({1'h0, add_515167, array_index_513530[1:0]}) < $signed({1'h0, sel_515170}) ? {add_515167, array_index_513530[1:0]} : sel_515170;
  assign add_515482 = array_index_513705[11:2] + 10'h2bb;
  assign sel_515485 = $signed({1'h0, add_515172, array_index_513533[1:0]}) < $signed({1'h0, sel_515175}) ? {add_515172, array_index_513533[1:0]} : sel_515175;
  assign add_515487 = array_index_513890[11:0] + 12'h8e1;
  assign sel_515489 = $signed({1'h0, add_515177}) < $signed({1'h0, sel_515179}) ? add_515177 : sel_515179;
  assign add_515491 = array_index_513893[11:0] + 12'h8e1;
  assign sel_515493 = $signed({1'h0, add_515181}) < $signed({1'h0, sel_515183}) ? add_515181 : sel_515183;
  assign add_515495 = array_index_514096[11:4] + 8'h83;
  assign sel_515498 = $signed({1'h0, add_515185, array_index_513890[3:0]}) < $signed({1'h0, sel_515188}) ? {add_515185, array_index_513890[3:0]} : sel_515188;
  assign add_515500 = array_index_514099[11:4] + 8'h83;
  assign sel_515503 = $signed({1'h0, add_515190, array_index_513893[3:0]}) < $signed({1'h0, sel_515193}) ? {add_515190, array_index_513893[3:0]} : sel_515193;
  assign add_515505 = array_index_514318[11:0] + 12'ha09;
  assign sel_515507 = $signed({1'h0, add_515195}) < $signed({1'h0, sel_515197}) ? add_515195 : sel_515197;
  assign add_515509 = array_index_514321[11:0] + 12'ha09;
  assign sel_515511 = $signed({1'h0, add_515199}) < $signed({1'h0, sel_515201}) ? add_515199 : sel_515201;
  assign add_515513 = array_index_514558[11:1] + 11'h6cb;
  assign sel_515515 = $signed({1'h0, add_515203, array_index_514318[0]}) < $signed({1'h0, sel_515205}) ? {add_515203, array_index_514318[0]} : sel_515205;
  assign add_515517 = array_index_514561[11:1] + 11'h6cb;
  assign sel_515519 = $signed({1'h0, add_515207, array_index_514321[0]}) < $signed({1'h0, sel_515209}) ? {add_515207, array_index_514321[0]} : sel_515209;
  assign add_515521 = array_index_514818[11:1] + 11'h75d;
  assign sel_515523 = $signed({1'h0, add_515211, array_index_514558[0]}) < $signed({1'h0, sel_515213}) ? {add_515211, array_index_514558[0]} : sel_515213;
  assign add_515525 = array_index_514821[11:1] + 11'h75d;
  assign sel_515527 = $signed({1'h0, add_515215, array_index_514561[0]}) < $signed({1'h0, sel_515217}) ? {add_515215, array_index_514561[0]} : sel_515217;
  assign add_515529 = array_index_515098[11:1] + 11'h24f;
  assign sel_515532 = $signed({1'h0, add_515219, array_index_514818[0]}) < $signed({1'h0, sel_515222}) ? {add_515219, array_index_514818[0]} : sel_515222;
  assign add_515534 = array_index_515101[11:1] + 11'h24f;
  assign sel_515537 = $signed({1'h0, add_515224, array_index_514821[0]}) < $signed({1'h0, sel_515227}) ? {add_515224, array_index_514821[0]} : sel_515227;
  assign add_515545 = array_index_512818[11:0] + 12'h7d5;
  assign add_515547 = array_index_512819[11:0] + 12'h7d5;
  assign add_515618 = array_index_515398[11:0] + 12'h62b;
  assign sel_515620 = $signed({1'h0, add_515298}) < $signed({1'h0, sel_515300}) ? add_515298 : sel_515300;
  assign add_515623 = array_index_515401[11:0] + 12'h62b;
  assign sel_515625 = $signed({1'h0, add_515303}) < $signed({1'h0, sel_515305}) ? add_515303 : sel_515305;
  assign add_515633 = array_index_512834[11:3] + 9'h0f5;
  assign sel_515635 = $signed({1'h0, add_515307, array_index_512818[2:0]}) < $signed(13'h0fff) ? {add_515307, array_index_512818[2:0]} : 12'hfff;
  assign add_515637 = array_index_512837[11:3] + 9'h0f5;
  assign sel_515639 = $signed({1'h0, add_515309, array_index_512819[2:0]}) < $signed(13'h0fff) ? {add_515309, array_index_512819[2:0]} : 12'hfff;
  assign array_index_515726 = set1_unflattened[5'h11];
  assign array_index_515729 = set2_unflattened[5'h11];
  assign add_515733 = array_index_512818[11:1] + 11'h179;
  assign add_515735 = array_index_512819[11:1] + 11'h179;
  assign add_515747 = array_index_512880[11:0] + 12'h067;
  assign sel_515749 = $signed({1'h0, add_515411}) < $signed({1'h0, sel_515413}) ? add_515411 : sel_515413;
  assign add_515751 = array_index_512883[11:0] + 12'h067;
  assign sel_515753 = $signed({1'h0, add_515415}) < $signed({1'h0, sel_515417}) ? add_515415 : sel_515417;
  assign add_515755 = array_index_512942[11:3] + 9'h1ef;
  assign sel_515758 = $signed({1'h0, add_515419, array_index_512880[2:0]}) < $signed({1'h0, sel_515422}) ? {add_515419, array_index_512880[2:0]} : sel_515422;
  assign add_515760 = array_index_512945[11:3] + 9'h1ef;
  assign sel_515763 = $signed({1'h0, add_515424, array_index_512883[2:0]}) < $signed({1'h0, sel_515427}) ? {add_515424, array_index_512883[2:0]} : sel_515427;
  assign add_515765 = array_index_513022[11:1] + 11'h2d5;
  assign sel_515767 = $signed({1'h0, add_515429, array_index_512942[0]}) < $signed({1'h0, sel_515431}) ? {add_515429, array_index_512942[0]} : sel_515431;
  assign add_515769 = array_index_513025[11:1] + 11'h2d5;
  assign sel_515771 = $signed({1'h0, add_515433, array_index_512945[0]}) < $signed({1'h0, sel_515435}) ? {add_515433, array_index_512945[0]} : sel_515435;
  assign add_515773 = array_index_513120[11:2] + 10'h353;
  assign sel_515775 = $signed({1'h0, add_515437, array_index_513022[1:0]}) < $signed({1'h0, sel_515439}) ? {add_515437, array_index_513022[1:0]} : sel_515439;
  assign add_515777 = array_index_513123[11:2] + 10'h353;
  assign sel_515779 = $signed({1'h0, add_515441, array_index_513025[1:0]}) < $signed({1'h0, sel_515443}) ? {add_515441, array_index_513025[1:0]} : sel_515443;
  assign add_515781 = array_index_513238[11:0] + 12'h0a7;
  assign sel_515783 = $signed({1'h0, add_515445}) < $signed({1'h0, sel_515447}) ? add_515445 : sel_515447;
  assign add_515785 = array_index_513241[11:0] + 12'h0a7;
  assign sel_515787 = $signed({1'h0, add_515449}) < $signed({1'h0, sel_515451}) ? add_515449 : sel_515451;
  assign add_515789 = array_index_513374[11:1] + 11'h4cb;
  assign sel_515791 = $signed({1'h0, add_515453, array_index_513238[0]}) < $signed({1'h0, sel_515455}) ? {add_515453, array_index_513238[0]} : sel_515455;
  assign add_515793 = array_index_513377[11:1] + 11'h4cb;
  assign sel_515795 = $signed({1'h0, add_515457, array_index_513241[0]}) < $signed({1'h0, sel_515459}) ? {add_515457, array_index_513241[0]} : sel_515459;
  assign add_515797 = array_index_513530[11:0] + 12'hfe9;
  assign sel_515799 = $signed({1'h0, add_515461}) < $signed({1'h0, sel_515463}) ? add_515461 : sel_515463;
  assign add_515801 = array_index_513533[11:0] + 12'hfe9;
  assign sel_515803 = $signed({1'h0, add_515465}) < $signed({1'h0, sel_515467}) ? add_515465 : sel_515467;
  assign add_515805 = array_index_513702[11:0] + 12'h97d;
  assign sel_515807 = $signed({1'h0, add_515469}) < $signed({1'h0, sel_515471}) ? add_515469 : sel_515471;
  assign add_515809 = array_index_513705[11:0] + 12'h97d;
  assign sel_515811 = $signed({1'h0, add_515473}) < $signed({1'h0, sel_515475}) ? add_515473 : sel_515475;
  assign add_515813 = array_index_513890[11:2] + 10'h2bb;
  assign sel_515816 = $signed({1'h0, add_515477, array_index_513702[1:0]}) < $signed({1'h0, sel_515480}) ? {add_515477, array_index_513702[1:0]} : sel_515480;
  assign add_515818 = array_index_513893[11:2] + 10'h2bb;
  assign sel_515821 = $signed({1'h0, add_515482, array_index_513705[1:0]}) < $signed({1'h0, sel_515485}) ? {add_515482, array_index_513705[1:0]} : sel_515485;
  assign add_515823 = array_index_514096[11:0] + 12'h8e1;
  assign sel_515825 = $signed({1'h0, add_515487}) < $signed({1'h0, sel_515489}) ? add_515487 : sel_515489;
  assign add_515827 = array_index_514099[11:0] + 12'h8e1;
  assign sel_515829 = $signed({1'h0, add_515491}) < $signed({1'h0, sel_515493}) ? add_515491 : sel_515493;
  assign add_515831 = array_index_514318[11:4] + 8'h83;
  assign sel_515834 = $signed({1'h0, add_515495, array_index_514096[3:0]}) < $signed({1'h0, sel_515498}) ? {add_515495, array_index_514096[3:0]} : sel_515498;
  assign add_515836 = array_index_514321[11:4] + 8'h83;
  assign sel_515839 = $signed({1'h0, add_515500, array_index_514099[3:0]}) < $signed({1'h0, sel_515503}) ? {add_515500, array_index_514099[3:0]} : sel_515503;
  assign add_515841 = array_index_514558[11:0] + 12'ha09;
  assign sel_515843 = $signed({1'h0, add_515505}) < $signed({1'h0, sel_515507}) ? add_515505 : sel_515507;
  assign add_515845 = array_index_514561[11:0] + 12'ha09;
  assign sel_515847 = $signed({1'h0, add_515509}) < $signed({1'h0, sel_515511}) ? add_515509 : sel_515511;
  assign add_515849 = array_index_514818[11:1] + 11'h6cb;
  assign sel_515851 = $signed({1'h0, add_515513, array_index_514558[0]}) < $signed({1'h0, sel_515515}) ? {add_515513, array_index_514558[0]} : sel_515515;
  assign add_515853 = array_index_514821[11:1] + 11'h6cb;
  assign sel_515855 = $signed({1'h0, add_515517, array_index_514561[0]}) < $signed({1'h0, sel_515519}) ? {add_515517, array_index_514561[0]} : sel_515519;
  assign add_515857 = array_index_515098[11:1] + 11'h75d;
  assign sel_515859 = $signed({1'h0, add_515521, array_index_514818[0]}) < $signed({1'h0, sel_515523}) ? {add_515521, array_index_514818[0]} : sel_515523;
  assign add_515861 = array_index_515101[11:1] + 11'h75d;
  assign sel_515863 = $signed({1'h0, add_515525, array_index_514821[0]}) < $signed({1'h0, sel_515527}) ? {add_515525, array_index_514821[0]} : sel_515527;
  assign add_515865 = array_index_515398[11:1] + 11'h24f;
  assign sel_515868 = $signed({1'h0, add_515529, array_index_515098[0]}) < $signed({1'h0, sel_515532}) ? {add_515529, array_index_515098[0]} : sel_515532;
  assign add_515870 = array_index_515401[11:1] + 11'h24f;
  assign sel_515873 = $signed({1'h0, add_515534, array_index_515101[0]}) < $signed({1'h0, sel_515537}) ? {add_515534, array_index_515101[0]} : sel_515537;
  assign add_515887 = array_index_512834[11:0] + 12'h7d5;
  assign sel_515889 = $signed({1'h0, add_515545}) < $signed(13'h0fff) ? add_515545 : 12'hfff;
  assign add_515891 = array_index_512837[11:0] + 12'h7d5;
  assign sel_515893 = $signed({1'h0, add_515547}) < $signed(13'h0fff) ? add_515547 : 12'hfff;
  assign add_515962 = array_index_515726[11:0] + 12'h62b;
  assign sel_515964 = $signed({1'h0, add_515618}) < $signed({1'h0, sel_515620}) ? add_515618 : sel_515620;
  assign add_515967 = array_index_515729[11:0] + 12'h62b;
  assign sel_515969 = $signed({1'h0, add_515623}) < $signed({1'h0, sel_515625}) ? add_515623 : sel_515625;
  assign add_515971 = array_index_512818[11:0] + 12'h45b;
  assign add_515973 = array_index_512819[11:0] + 12'h45b;
  assign add_515987 = array_index_512880[11:3] + 9'h0f5;
  assign sel_515989 = $signed({1'h0, add_515633, array_index_512834[2:0]}) < $signed({1'h0, sel_515635}) ? {add_515633, array_index_512834[2:0]} : sel_515635;
  assign add_515991 = array_index_512883[11:3] + 9'h0f5;
  assign sel_515993 = $signed({1'h0, add_515637, array_index_512837[2:0]}) < $signed({1'h0, sel_515639}) ? {add_515637, array_index_512837[2:0]} : sel_515639;
  assign array_index_516080 = set1_unflattened[5'h12];
  assign array_index_516083 = set2_unflattened[5'h12];
  assign add_516093 = array_index_512834[11:1] + 11'h179;
  assign sel_516095 = $signed({1'h0, add_515733, array_index_512818[0]}) < $signed(13'h0fff) ? {add_515733, array_index_512818[0]} : 12'hfff;
  assign add_516097 = array_index_512837[11:1] + 11'h179;
  assign sel_516099 = $signed({1'h0, add_515735, array_index_512819[0]}) < $signed(13'h0fff) ? {add_515735, array_index_512819[0]} : 12'hfff;
  assign add_516109 = array_index_512942[11:0] + 12'h067;
  assign sel_516111 = $signed({1'h0, add_515747}) < $signed({1'h0, sel_515749}) ? add_515747 : sel_515749;
  assign add_516113 = array_index_512945[11:0] + 12'h067;
  assign sel_516115 = $signed({1'h0, add_515751}) < $signed({1'h0, sel_515753}) ? add_515751 : sel_515753;
  assign add_516117 = array_index_513022[11:3] + 9'h1ef;
  assign sel_516120 = $signed({1'h0, add_515755, array_index_512942[2:0]}) < $signed({1'h0, sel_515758}) ? {add_515755, array_index_512942[2:0]} : sel_515758;
  assign add_516122 = array_index_513025[11:3] + 9'h1ef;
  assign sel_516125 = $signed({1'h0, add_515760, array_index_512945[2:0]}) < $signed({1'h0, sel_515763}) ? {add_515760, array_index_512945[2:0]} : sel_515763;
  assign add_516127 = array_index_513120[11:1] + 11'h2d5;
  assign sel_516129 = $signed({1'h0, add_515765, array_index_513022[0]}) < $signed({1'h0, sel_515767}) ? {add_515765, array_index_513022[0]} : sel_515767;
  assign add_516131 = array_index_513123[11:1] + 11'h2d5;
  assign sel_516133 = $signed({1'h0, add_515769, array_index_513025[0]}) < $signed({1'h0, sel_515771}) ? {add_515769, array_index_513025[0]} : sel_515771;
  assign add_516135 = array_index_513238[11:2] + 10'h353;
  assign sel_516137 = $signed({1'h0, add_515773, array_index_513120[1:0]}) < $signed({1'h0, sel_515775}) ? {add_515773, array_index_513120[1:0]} : sel_515775;
  assign add_516139 = array_index_513241[11:2] + 10'h353;
  assign sel_516141 = $signed({1'h0, add_515777, array_index_513123[1:0]}) < $signed({1'h0, sel_515779}) ? {add_515777, array_index_513123[1:0]} : sel_515779;
  assign add_516143 = array_index_513374[11:0] + 12'h0a7;
  assign sel_516145 = $signed({1'h0, add_515781}) < $signed({1'h0, sel_515783}) ? add_515781 : sel_515783;
  assign add_516147 = array_index_513377[11:0] + 12'h0a7;
  assign sel_516149 = $signed({1'h0, add_515785}) < $signed({1'h0, sel_515787}) ? add_515785 : sel_515787;
  assign add_516151 = array_index_513530[11:1] + 11'h4cb;
  assign sel_516153 = $signed({1'h0, add_515789, array_index_513374[0]}) < $signed({1'h0, sel_515791}) ? {add_515789, array_index_513374[0]} : sel_515791;
  assign add_516155 = array_index_513533[11:1] + 11'h4cb;
  assign sel_516157 = $signed({1'h0, add_515793, array_index_513377[0]}) < $signed({1'h0, sel_515795}) ? {add_515793, array_index_513377[0]} : sel_515795;
  assign add_516159 = array_index_513702[11:0] + 12'hfe9;
  assign sel_516161 = $signed({1'h0, add_515797}) < $signed({1'h0, sel_515799}) ? add_515797 : sel_515799;
  assign add_516163 = array_index_513705[11:0] + 12'hfe9;
  assign sel_516165 = $signed({1'h0, add_515801}) < $signed({1'h0, sel_515803}) ? add_515801 : sel_515803;
  assign add_516167 = array_index_513890[11:0] + 12'h97d;
  assign sel_516169 = $signed({1'h0, add_515805}) < $signed({1'h0, sel_515807}) ? add_515805 : sel_515807;
  assign add_516171 = array_index_513893[11:0] + 12'h97d;
  assign sel_516173 = $signed({1'h0, add_515809}) < $signed({1'h0, sel_515811}) ? add_515809 : sel_515811;
  assign add_516175 = array_index_514096[11:2] + 10'h2bb;
  assign sel_516178 = $signed({1'h0, add_515813, array_index_513890[1:0]}) < $signed({1'h0, sel_515816}) ? {add_515813, array_index_513890[1:0]} : sel_515816;
  assign add_516180 = array_index_514099[11:2] + 10'h2bb;
  assign sel_516183 = $signed({1'h0, add_515818, array_index_513893[1:0]}) < $signed({1'h0, sel_515821}) ? {add_515818, array_index_513893[1:0]} : sel_515821;
  assign add_516185 = array_index_514318[11:0] + 12'h8e1;
  assign sel_516187 = $signed({1'h0, add_515823}) < $signed({1'h0, sel_515825}) ? add_515823 : sel_515825;
  assign add_516189 = array_index_514321[11:0] + 12'h8e1;
  assign sel_516191 = $signed({1'h0, add_515827}) < $signed({1'h0, sel_515829}) ? add_515827 : sel_515829;
  assign add_516193 = array_index_514558[11:4] + 8'h83;
  assign sel_516196 = $signed({1'h0, add_515831, array_index_514318[3:0]}) < $signed({1'h0, sel_515834}) ? {add_515831, array_index_514318[3:0]} : sel_515834;
  assign add_516198 = array_index_514561[11:4] + 8'h83;
  assign sel_516201 = $signed({1'h0, add_515836, array_index_514321[3:0]}) < $signed({1'h0, sel_515839}) ? {add_515836, array_index_514321[3:0]} : sel_515839;
  assign add_516203 = array_index_514818[11:0] + 12'ha09;
  assign sel_516205 = $signed({1'h0, add_515841}) < $signed({1'h0, sel_515843}) ? add_515841 : sel_515843;
  assign add_516207 = array_index_514821[11:0] + 12'ha09;
  assign sel_516209 = $signed({1'h0, add_515845}) < $signed({1'h0, sel_515847}) ? add_515845 : sel_515847;
  assign add_516211 = array_index_515098[11:1] + 11'h6cb;
  assign sel_516213 = $signed({1'h0, add_515849, array_index_514818[0]}) < $signed({1'h0, sel_515851}) ? {add_515849, array_index_514818[0]} : sel_515851;
  assign add_516215 = array_index_515101[11:1] + 11'h6cb;
  assign sel_516217 = $signed({1'h0, add_515853, array_index_514821[0]}) < $signed({1'h0, sel_515855}) ? {add_515853, array_index_514821[0]} : sel_515855;
  assign add_516219 = array_index_515398[11:1] + 11'h75d;
  assign sel_516221 = $signed({1'h0, add_515857, array_index_515098[0]}) < $signed({1'h0, sel_515859}) ? {add_515857, array_index_515098[0]} : sel_515859;
  assign add_516223 = array_index_515401[11:1] + 11'h75d;
  assign sel_516225 = $signed({1'h0, add_515861, array_index_515101[0]}) < $signed({1'h0, sel_515863}) ? {add_515861, array_index_515101[0]} : sel_515863;
  assign add_516227 = array_index_515726[11:1] + 11'h24f;
  assign sel_516230 = $signed({1'h0, add_515865, array_index_515398[0]}) < $signed({1'h0, sel_515868}) ? {add_515865, array_index_515398[0]} : sel_515868;
  assign add_516232 = array_index_515729[11:1] + 11'h24f;
  assign sel_516235 = $signed({1'h0, add_515870, array_index_515401[0]}) < $signed({1'h0, sel_515873}) ? {add_515870, array_index_515401[0]} : sel_515873;
  assign add_516243 = array_index_512818[11:0] + 12'h6ab;
  assign add_516245 = array_index_512819[11:0] + 12'h6ab;
  assign add_516257 = array_index_512880[11:0] + 12'h7d5;
  assign sel_516259 = $signed({1'h0, add_515887}) < $signed({1'h0, sel_515889}) ? add_515887 : sel_515889;
  assign add_516261 = array_index_512883[11:0] + 12'h7d5;
  assign sel_516263 = $signed({1'h0, add_515891}) < $signed({1'h0, sel_515893}) ? add_515891 : sel_515893;
  assign add_516332 = array_index_516080[11:0] + 12'h62b;
  assign sel_516334 = $signed({1'h0, add_515962}) < $signed({1'h0, sel_515964}) ? add_515962 : sel_515964;
  assign add_516337 = array_index_516083[11:0] + 12'h62b;
  assign sel_516339 = $signed({1'h0, add_515967}) < $signed({1'h0, sel_515969}) ? add_515967 : sel_515969;
  assign add_516347 = array_index_512834[11:0] + 12'h45b;
  assign sel_516349 = $signed({1'h0, add_515971}) < $signed(13'h0fff) ? add_515971 : 12'hfff;
  assign add_516351 = array_index_512837[11:0] + 12'h45b;
  assign sel_516353 = $signed({1'h0, add_515973}) < $signed(13'h0fff) ? add_515973 : 12'hfff;
  assign add_516365 = array_index_512942[11:3] + 9'h0f5;
  assign sel_516367 = $signed({1'h0, add_515987, array_index_512880[2:0]}) < $signed({1'h0, sel_515989}) ? {add_515987, array_index_512880[2:0]} : sel_515989;
  assign add_516369 = array_index_512945[11:3] + 9'h0f5;
  assign sel_516371 = $signed({1'h0, add_515991, array_index_512883[2:0]}) < $signed({1'h0, sel_515993}) ? {add_515991, array_index_512883[2:0]} : sel_515993;
  assign array_index_516458 = set1_unflattened[5'h13];
  assign array_index_516461 = set2_unflattened[5'h13];
  assign add_516465 = array_index_512818[11:0] + 12'hee1;
  assign add_516467 = array_index_512819[11:0] + 12'hee1;
  assign add_516479 = array_index_512880[11:1] + 11'h179;
  assign sel_516481 = $signed({1'h0, add_516093, array_index_512834[0]}) < $signed({1'h0, sel_516095}) ? {add_516093, array_index_512834[0]} : sel_516095;
  assign add_516483 = array_index_512883[11:1] + 11'h179;
  assign sel_516485 = $signed({1'h0, add_516097, array_index_512837[0]}) < $signed({1'h0, sel_516099}) ? {add_516097, array_index_512837[0]} : sel_516099;
  assign add_516495 = array_index_513022[11:0] + 12'h067;
  assign sel_516497 = $signed({1'h0, add_516109}) < $signed({1'h0, sel_516111}) ? add_516109 : sel_516111;
  assign add_516499 = array_index_513025[11:0] + 12'h067;
  assign sel_516501 = $signed({1'h0, add_516113}) < $signed({1'h0, sel_516115}) ? add_516113 : sel_516115;
  assign add_516503 = array_index_513120[11:3] + 9'h1ef;
  assign sel_516506 = $signed({1'h0, add_516117, array_index_513022[2:0]}) < $signed({1'h0, sel_516120}) ? {add_516117, array_index_513022[2:0]} : sel_516120;
  assign add_516508 = array_index_513123[11:3] + 9'h1ef;
  assign sel_516511 = $signed({1'h0, add_516122, array_index_513025[2:0]}) < $signed({1'h0, sel_516125}) ? {add_516122, array_index_513025[2:0]} : sel_516125;
  assign add_516513 = array_index_513238[11:1] + 11'h2d5;
  assign sel_516515 = $signed({1'h0, add_516127, array_index_513120[0]}) < $signed({1'h0, sel_516129}) ? {add_516127, array_index_513120[0]} : sel_516129;
  assign add_516517 = array_index_513241[11:1] + 11'h2d5;
  assign sel_516519 = $signed({1'h0, add_516131, array_index_513123[0]}) < $signed({1'h0, sel_516133}) ? {add_516131, array_index_513123[0]} : sel_516133;
  assign add_516521 = array_index_513374[11:2] + 10'h353;
  assign sel_516523 = $signed({1'h0, add_516135, array_index_513238[1:0]}) < $signed({1'h0, sel_516137}) ? {add_516135, array_index_513238[1:0]} : sel_516137;
  assign add_516525 = array_index_513377[11:2] + 10'h353;
  assign sel_516527 = $signed({1'h0, add_516139, array_index_513241[1:0]}) < $signed({1'h0, sel_516141}) ? {add_516139, array_index_513241[1:0]} : sel_516141;
  assign add_516529 = array_index_513530[11:0] + 12'h0a7;
  assign sel_516531 = $signed({1'h0, add_516143}) < $signed({1'h0, sel_516145}) ? add_516143 : sel_516145;
  assign add_516533 = array_index_513533[11:0] + 12'h0a7;
  assign sel_516535 = $signed({1'h0, add_516147}) < $signed({1'h0, sel_516149}) ? add_516147 : sel_516149;
  assign add_516537 = array_index_513702[11:1] + 11'h4cb;
  assign sel_516539 = $signed({1'h0, add_516151, array_index_513530[0]}) < $signed({1'h0, sel_516153}) ? {add_516151, array_index_513530[0]} : sel_516153;
  assign add_516541 = array_index_513705[11:1] + 11'h4cb;
  assign sel_516543 = $signed({1'h0, add_516155, array_index_513533[0]}) < $signed({1'h0, sel_516157}) ? {add_516155, array_index_513533[0]} : sel_516157;
  assign add_516545 = array_index_513890[11:0] + 12'hfe9;
  assign sel_516547 = $signed({1'h0, add_516159}) < $signed({1'h0, sel_516161}) ? add_516159 : sel_516161;
  assign add_516549 = array_index_513893[11:0] + 12'hfe9;
  assign sel_516551 = $signed({1'h0, add_516163}) < $signed({1'h0, sel_516165}) ? add_516163 : sel_516165;
  assign add_516553 = array_index_514096[11:0] + 12'h97d;
  assign sel_516555 = $signed({1'h0, add_516167}) < $signed({1'h0, sel_516169}) ? add_516167 : sel_516169;
  assign add_516557 = array_index_514099[11:0] + 12'h97d;
  assign sel_516559 = $signed({1'h0, add_516171}) < $signed({1'h0, sel_516173}) ? add_516171 : sel_516173;
  assign add_516561 = array_index_514318[11:2] + 10'h2bb;
  assign sel_516564 = $signed({1'h0, add_516175, array_index_514096[1:0]}) < $signed({1'h0, sel_516178}) ? {add_516175, array_index_514096[1:0]} : sel_516178;
  assign add_516566 = array_index_514321[11:2] + 10'h2bb;
  assign sel_516569 = $signed({1'h0, add_516180, array_index_514099[1:0]}) < $signed({1'h0, sel_516183}) ? {add_516180, array_index_514099[1:0]} : sel_516183;
  assign add_516571 = array_index_514558[11:0] + 12'h8e1;
  assign sel_516573 = $signed({1'h0, add_516185}) < $signed({1'h0, sel_516187}) ? add_516185 : sel_516187;
  assign add_516575 = array_index_514561[11:0] + 12'h8e1;
  assign sel_516577 = $signed({1'h0, add_516189}) < $signed({1'h0, sel_516191}) ? add_516189 : sel_516191;
  assign add_516579 = array_index_514818[11:4] + 8'h83;
  assign sel_516582 = $signed({1'h0, add_516193, array_index_514558[3:0]}) < $signed({1'h0, sel_516196}) ? {add_516193, array_index_514558[3:0]} : sel_516196;
  assign add_516584 = array_index_514821[11:4] + 8'h83;
  assign sel_516587 = $signed({1'h0, add_516198, array_index_514561[3:0]}) < $signed({1'h0, sel_516201}) ? {add_516198, array_index_514561[3:0]} : sel_516201;
  assign add_516589 = array_index_515098[11:0] + 12'ha09;
  assign sel_516591 = $signed({1'h0, add_516203}) < $signed({1'h0, sel_516205}) ? add_516203 : sel_516205;
  assign add_516593 = array_index_515101[11:0] + 12'ha09;
  assign sel_516595 = $signed({1'h0, add_516207}) < $signed({1'h0, sel_516209}) ? add_516207 : sel_516209;
  assign add_516597 = array_index_515398[11:1] + 11'h6cb;
  assign sel_516599 = $signed({1'h0, add_516211, array_index_515098[0]}) < $signed({1'h0, sel_516213}) ? {add_516211, array_index_515098[0]} : sel_516213;
  assign add_516601 = array_index_515401[11:1] + 11'h6cb;
  assign sel_516603 = $signed({1'h0, add_516215, array_index_515101[0]}) < $signed({1'h0, sel_516217}) ? {add_516215, array_index_515101[0]} : sel_516217;
  assign add_516605 = array_index_515726[11:1] + 11'h75d;
  assign sel_516607 = $signed({1'h0, add_516219, array_index_515398[0]}) < $signed({1'h0, sel_516221}) ? {add_516219, array_index_515398[0]} : sel_516221;
  assign add_516609 = array_index_515729[11:1] + 11'h75d;
  assign sel_516611 = $signed({1'h0, add_516223, array_index_515401[0]}) < $signed({1'h0, sel_516225}) ? {add_516223, array_index_515401[0]} : sel_516225;
  assign add_516613 = array_index_516080[11:1] + 11'h24f;
  assign sel_516616 = $signed({1'h0, add_516227, array_index_515726[0]}) < $signed({1'h0, sel_516230}) ? {add_516227, array_index_515726[0]} : sel_516230;
  assign add_516618 = array_index_516083[11:1] + 11'h24f;
  assign sel_516621 = $signed({1'h0, add_516232, array_index_515729[0]}) < $signed({1'h0, sel_516235}) ? {add_516232, array_index_515729[0]} : sel_516235;
  assign add_516635 = array_index_512834[11:0] + 12'h6ab;
  assign sel_516637 = $signed({1'h0, add_516243}) < $signed(13'h0fff) ? add_516243 : 12'hfff;
  assign add_516639 = array_index_512837[11:0] + 12'h6ab;
  assign sel_516641 = $signed({1'h0, add_516245}) < $signed(13'h0fff) ? add_516245 : 12'hfff;
  assign add_516651 = array_index_512942[11:0] + 12'h7d5;
  assign sel_516653 = $signed({1'h0, add_516257}) < $signed({1'h0, sel_516259}) ? add_516257 : sel_516259;
  assign add_516655 = array_index_512945[11:0] + 12'h7d5;
  assign sel_516657 = $signed({1'h0, add_516261}) < $signed({1'h0, sel_516263}) ? add_516261 : sel_516263;
  assign add_516726 = array_index_516458[11:0] + 12'h62b;
  assign sel_516728 = $signed({1'h0, add_516332}) < $signed({1'h0, sel_516334}) ? add_516332 : sel_516334;
  assign add_516731 = array_index_516461[11:0] + 12'h62b;
  assign sel_516733 = $signed({1'h0, add_516337}) < $signed({1'h0, sel_516339}) ? add_516337 : sel_516339;
  assign add_516735 = array_index_512818[11:0] + 12'h81f;
  assign add_516737 = array_index_512819[11:0] + 12'h81f;
  assign add_516749 = array_index_512880[11:0] + 12'h45b;
  assign sel_516751 = $signed({1'h0, add_516347}) < $signed({1'h0, sel_516349}) ? add_516347 : sel_516349;
  assign add_516753 = array_index_512883[11:0] + 12'h45b;
  assign sel_516755 = $signed({1'h0, add_516351}) < $signed({1'h0, sel_516353}) ? add_516351 : sel_516353;
  assign add_516767 = array_index_513022[11:3] + 9'h0f5;
  assign sel_516769 = $signed({1'h0, add_516365, array_index_512942[2:0]}) < $signed({1'h0, sel_516367}) ? {add_516365, array_index_512942[2:0]} : sel_516367;
  assign add_516771 = array_index_513025[11:3] + 9'h0f5;
  assign sel_516773 = $signed({1'h0, add_516369, array_index_512945[2:0]}) < $signed({1'h0, sel_516371}) ? {add_516369, array_index_512945[2:0]} : sel_516371;
  assign array_index_516860 = set1_unflattened[5'h14];
  assign array_index_516863 = set2_unflattened[5'h14];
  assign add_516873 = array_index_512834[11:0] + 12'hee1;
  assign sel_516875 = $signed({1'h0, add_516465}) < $signed(13'h0fff) ? add_516465 : 12'hfff;
  assign add_516877 = array_index_512837[11:0] + 12'hee1;
  assign sel_516879 = $signed({1'h0, add_516467}) < $signed(13'h0fff) ? add_516467 : 12'hfff;
  assign add_516889 = array_index_512942[11:1] + 11'h179;
  assign sel_516891 = $signed({1'h0, add_516479, array_index_512880[0]}) < $signed({1'h0, sel_516481}) ? {add_516479, array_index_512880[0]} : sel_516481;
  assign add_516893 = array_index_512945[11:1] + 11'h179;
  assign sel_516895 = $signed({1'h0, add_516483, array_index_512883[0]}) < $signed({1'h0, sel_516485}) ? {add_516483, array_index_512883[0]} : sel_516485;
  assign add_516905 = array_index_513120[11:0] + 12'h067;
  assign sel_516907 = $signed({1'h0, add_516495}) < $signed({1'h0, sel_516497}) ? add_516495 : sel_516497;
  assign add_516909 = array_index_513123[11:0] + 12'h067;
  assign sel_516911 = $signed({1'h0, add_516499}) < $signed({1'h0, sel_516501}) ? add_516499 : sel_516501;
  assign add_516913 = array_index_513238[11:3] + 9'h1ef;
  assign sel_516916 = $signed({1'h0, add_516503, array_index_513120[2:0]}) < $signed({1'h0, sel_516506}) ? {add_516503, array_index_513120[2:0]} : sel_516506;
  assign add_516918 = array_index_513241[11:3] + 9'h1ef;
  assign sel_516921 = $signed({1'h0, add_516508, array_index_513123[2:0]}) < $signed({1'h0, sel_516511}) ? {add_516508, array_index_513123[2:0]} : sel_516511;
  assign add_516923 = array_index_513374[11:1] + 11'h2d5;
  assign sel_516925 = $signed({1'h0, add_516513, array_index_513238[0]}) < $signed({1'h0, sel_516515}) ? {add_516513, array_index_513238[0]} : sel_516515;
  assign add_516927 = array_index_513377[11:1] + 11'h2d5;
  assign sel_516929 = $signed({1'h0, add_516517, array_index_513241[0]}) < $signed({1'h0, sel_516519}) ? {add_516517, array_index_513241[0]} : sel_516519;
  assign add_516931 = array_index_513530[11:2] + 10'h353;
  assign sel_516933 = $signed({1'h0, add_516521, array_index_513374[1:0]}) < $signed({1'h0, sel_516523}) ? {add_516521, array_index_513374[1:0]} : sel_516523;
  assign add_516935 = array_index_513533[11:2] + 10'h353;
  assign sel_516937 = $signed({1'h0, add_516525, array_index_513377[1:0]}) < $signed({1'h0, sel_516527}) ? {add_516525, array_index_513377[1:0]} : sel_516527;
  assign add_516939 = array_index_513702[11:0] + 12'h0a7;
  assign sel_516941 = $signed({1'h0, add_516529}) < $signed({1'h0, sel_516531}) ? add_516529 : sel_516531;
  assign add_516943 = array_index_513705[11:0] + 12'h0a7;
  assign sel_516945 = $signed({1'h0, add_516533}) < $signed({1'h0, sel_516535}) ? add_516533 : sel_516535;
  assign add_516947 = array_index_513890[11:1] + 11'h4cb;
  assign sel_516949 = $signed({1'h0, add_516537, array_index_513702[0]}) < $signed({1'h0, sel_516539}) ? {add_516537, array_index_513702[0]} : sel_516539;
  assign add_516951 = array_index_513893[11:1] + 11'h4cb;
  assign sel_516953 = $signed({1'h0, add_516541, array_index_513705[0]}) < $signed({1'h0, sel_516543}) ? {add_516541, array_index_513705[0]} : sel_516543;
  assign add_516955 = array_index_514096[11:0] + 12'hfe9;
  assign sel_516957 = $signed({1'h0, add_516545}) < $signed({1'h0, sel_516547}) ? add_516545 : sel_516547;
  assign add_516959 = array_index_514099[11:0] + 12'hfe9;
  assign sel_516961 = $signed({1'h0, add_516549}) < $signed({1'h0, sel_516551}) ? add_516549 : sel_516551;
  assign add_516963 = array_index_514318[11:0] + 12'h97d;
  assign sel_516965 = $signed({1'h0, add_516553}) < $signed({1'h0, sel_516555}) ? add_516553 : sel_516555;
  assign add_516967 = array_index_514321[11:0] + 12'h97d;
  assign sel_516969 = $signed({1'h0, add_516557}) < $signed({1'h0, sel_516559}) ? add_516557 : sel_516559;
  assign add_516971 = array_index_514558[11:2] + 10'h2bb;
  assign sel_516974 = $signed({1'h0, add_516561, array_index_514318[1:0]}) < $signed({1'h0, sel_516564}) ? {add_516561, array_index_514318[1:0]} : sel_516564;
  assign add_516976 = array_index_514561[11:2] + 10'h2bb;
  assign sel_516979 = $signed({1'h0, add_516566, array_index_514321[1:0]}) < $signed({1'h0, sel_516569}) ? {add_516566, array_index_514321[1:0]} : sel_516569;
  assign add_516981 = array_index_514818[11:0] + 12'h8e1;
  assign sel_516983 = $signed({1'h0, add_516571}) < $signed({1'h0, sel_516573}) ? add_516571 : sel_516573;
  assign add_516985 = array_index_514821[11:0] + 12'h8e1;
  assign sel_516987 = $signed({1'h0, add_516575}) < $signed({1'h0, sel_516577}) ? add_516575 : sel_516577;
  assign add_516989 = array_index_515098[11:4] + 8'h83;
  assign sel_516992 = $signed({1'h0, add_516579, array_index_514818[3:0]}) < $signed({1'h0, sel_516582}) ? {add_516579, array_index_514818[3:0]} : sel_516582;
  assign add_516994 = array_index_515101[11:4] + 8'h83;
  assign sel_516997 = $signed({1'h0, add_516584, array_index_514821[3:0]}) < $signed({1'h0, sel_516587}) ? {add_516584, array_index_514821[3:0]} : sel_516587;
  assign add_516999 = array_index_515398[11:0] + 12'ha09;
  assign sel_517001 = $signed({1'h0, add_516589}) < $signed({1'h0, sel_516591}) ? add_516589 : sel_516591;
  assign add_517003 = array_index_515401[11:0] + 12'ha09;
  assign sel_517005 = $signed({1'h0, add_516593}) < $signed({1'h0, sel_516595}) ? add_516593 : sel_516595;
  assign add_517007 = array_index_515726[11:1] + 11'h6cb;
  assign sel_517009 = $signed({1'h0, add_516597, array_index_515398[0]}) < $signed({1'h0, sel_516599}) ? {add_516597, array_index_515398[0]} : sel_516599;
  assign add_517011 = array_index_515729[11:1] + 11'h6cb;
  assign sel_517013 = $signed({1'h0, add_516601, array_index_515401[0]}) < $signed({1'h0, sel_516603}) ? {add_516601, array_index_515401[0]} : sel_516603;
  assign add_517015 = array_index_516080[11:1] + 11'h75d;
  assign sel_517017 = $signed({1'h0, add_516605, array_index_515726[0]}) < $signed({1'h0, sel_516607}) ? {add_516605, array_index_515726[0]} : sel_516607;
  assign add_517019 = array_index_516083[11:1] + 11'h75d;
  assign sel_517021 = $signed({1'h0, add_516609, array_index_515729[0]}) < $signed({1'h0, sel_516611}) ? {add_516609, array_index_515729[0]} : sel_516611;
  assign add_517023 = array_index_516458[11:1] + 11'h24f;
  assign sel_517026 = $signed({1'h0, add_516613, array_index_516080[0]}) < $signed({1'h0, sel_516616}) ? {add_516613, array_index_516080[0]} : sel_516616;
  assign add_517028 = array_index_516461[11:1] + 11'h24f;
  assign sel_517031 = $signed({1'h0, add_516618, array_index_516083[0]}) < $signed({1'h0, sel_516621}) ? {add_516618, array_index_516083[0]} : sel_516621;
  assign add_517039 = array_index_512818[11:0] + 12'hbb1;
  assign add_517041 = array_index_512819[11:0] + 12'hbb1;
  assign add_517053 = array_index_512880[11:0] + 12'h6ab;
  assign sel_517055 = $signed({1'h0, add_516635}) < $signed({1'h0, sel_516637}) ? add_516635 : sel_516637;
  assign add_517057 = array_index_512883[11:0] + 12'h6ab;
  assign sel_517059 = $signed({1'h0, add_516639}) < $signed({1'h0, sel_516641}) ? add_516639 : sel_516641;
  assign add_517069 = array_index_513022[11:0] + 12'h7d5;
  assign sel_517071 = $signed({1'h0, add_516651}) < $signed({1'h0, sel_516653}) ? add_516651 : sel_516653;
  assign add_517073 = array_index_513025[11:0] + 12'h7d5;
  assign sel_517075 = $signed({1'h0, add_516655}) < $signed({1'h0, sel_516657}) ? add_516655 : sel_516657;
  assign add_517144 = array_index_516860[11:0] + 12'h62b;
  assign sel_517146 = $signed({1'h0, add_516726}) < $signed({1'h0, sel_516728}) ? add_516726 : sel_516728;
  assign add_517149 = array_index_516863[11:0] + 12'h62b;
  assign sel_517151 = $signed({1'h0, add_516731}) < $signed({1'h0, sel_516733}) ? add_516731 : sel_516733;
  assign add_517159 = array_index_512834[11:0] + 12'h81f;
  assign sel_517161 = $signed({1'h0, add_516735}) < $signed(13'h0fff) ? add_516735 : 12'hfff;
  assign add_517163 = array_index_512837[11:0] + 12'h81f;
  assign sel_517165 = $signed({1'h0, add_516737}) < $signed(13'h0fff) ? add_516737 : 12'hfff;
  assign add_517175 = array_index_512942[11:0] + 12'h45b;
  assign sel_517177 = $signed({1'h0, add_516749}) < $signed({1'h0, sel_516751}) ? add_516749 : sel_516751;
  assign add_517179 = array_index_512945[11:0] + 12'h45b;
  assign sel_517181 = $signed({1'h0, add_516753}) < $signed({1'h0, sel_516755}) ? add_516753 : sel_516755;
  assign add_517193 = array_index_513120[11:3] + 9'h0f5;
  assign sel_517195 = $signed({1'h0, add_516767, array_index_513022[2:0]}) < $signed({1'h0, sel_516769}) ? {add_516767, array_index_513022[2:0]} : sel_516769;
  assign add_517197 = array_index_513123[11:3] + 9'h0f5;
  assign sel_517199 = $signed({1'h0, add_516771, array_index_513025[2:0]}) < $signed({1'h0, sel_516773}) ? {add_516771, array_index_513025[2:0]} : sel_516773;
  assign array_index_517286 = set1_unflattened[5'h15];
  assign array_index_517289 = set2_unflattened[5'h15];
  assign add_517293 = array_index_512818[11:0] + 12'h437;
  assign add_517295 = array_index_512819[11:0] + 12'h437;
  assign add_517307 = array_index_512880[11:0] + 12'hee1;
  assign sel_517309 = $signed({1'h0, add_516873}) < $signed({1'h0, sel_516875}) ? add_516873 : sel_516875;
  assign add_517311 = array_index_512883[11:0] + 12'hee1;
  assign sel_517313 = $signed({1'h0, add_516877}) < $signed({1'h0, sel_516879}) ? add_516877 : sel_516879;
  assign add_517323 = array_index_513022[11:1] + 11'h179;
  assign sel_517325 = $signed({1'h0, add_516889, array_index_512942[0]}) < $signed({1'h0, sel_516891}) ? {add_516889, array_index_512942[0]} : sel_516891;
  assign add_517327 = array_index_513025[11:1] + 11'h179;
  assign sel_517329 = $signed({1'h0, add_516893, array_index_512945[0]}) < $signed({1'h0, sel_516895}) ? {add_516893, array_index_512945[0]} : sel_516895;
  assign add_517339 = array_index_513238[11:0] + 12'h067;
  assign sel_517341 = $signed({1'h0, add_516905}) < $signed({1'h0, sel_516907}) ? add_516905 : sel_516907;
  assign add_517343 = array_index_513241[11:0] + 12'h067;
  assign sel_517345 = $signed({1'h0, add_516909}) < $signed({1'h0, sel_516911}) ? add_516909 : sel_516911;
  assign add_517347 = array_index_513374[11:3] + 9'h1ef;
  assign sel_517350 = $signed({1'h0, add_516913, array_index_513238[2:0]}) < $signed({1'h0, sel_516916}) ? {add_516913, array_index_513238[2:0]} : sel_516916;
  assign add_517352 = array_index_513377[11:3] + 9'h1ef;
  assign sel_517355 = $signed({1'h0, add_516918, array_index_513241[2:0]}) < $signed({1'h0, sel_516921}) ? {add_516918, array_index_513241[2:0]} : sel_516921;
  assign add_517357 = array_index_513530[11:1] + 11'h2d5;
  assign sel_517359 = $signed({1'h0, add_516923, array_index_513374[0]}) < $signed({1'h0, sel_516925}) ? {add_516923, array_index_513374[0]} : sel_516925;
  assign add_517361 = array_index_513533[11:1] + 11'h2d5;
  assign sel_517363 = $signed({1'h0, add_516927, array_index_513377[0]}) < $signed({1'h0, sel_516929}) ? {add_516927, array_index_513377[0]} : sel_516929;
  assign add_517365 = array_index_513702[11:2] + 10'h353;
  assign sel_517367 = $signed({1'h0, add_516931, array_index_513530[1:0]}) < $signed({1'h0, sel_516933}) ? {add_516931, array_index_513530[1:0]} : sel_516933;
  assign add_517369 = array_index_513705[11:2] + 10'h353;
  assign sel_517371 = $signed({1'h0, add_516935, array_index_513533[1:0]}) < $signed({1'h0, sel_516937}) ? {add_516935, array_index_513533[1:0]} : sel_516937;
  assign add_517373 = array_index_513890[11:0] + 12'h0a7;
  assign sel_517375 = $signed({1'h0, add_516939}) < $signed({1'h0, sel_516941}) ? add_516939 : sel_516941;
  assign add_517377 = array_index_513893[11:0] + 12'h0a7;
  assign sel_517379 = $signed({1'h0, add_516943}) < $signed({1'h0, sel_516945}) ? add_516943 : sel_516945;
  assign add_517381 = array_index_514096[11:1] + 11'h4cb;
  assign sel_517383 = $signed({1'h0, add_516947, array_index_513890[0]}) < $signed({1'h0, sel_516949}) ? {add_516947, array_index_513890[0]} : sel_516949;
  assign add_517385 = array_index_514099[11:1] + 11'h4cb;
  assign sel_517387 = $signed({1'h0, add_516951, array_index_513893[0]}) < $signed({1'h0, sel_516953}) ? {add_516951, array_index_513893[0]} : sel_516953;
  assign add_517389 = array_index_514318[11:0] + 12'hfe9;
  assign sel_517391 = $signed({1'h0, add_516955}) < $signed({1'h0, sel_516957}) ? add_516955 : sel_516957;
  assign add_517393 = array_index_514321[11:0] + 12'hfe9;
  assign sel_517395 = $signed({1'h0, add_516959}) < $signed({1'h0, sel_516961}) ? add_516959 : sel_516961;
  assign add_517397 = array_index_514558[11:0] + 12'h97d;
  assign sel_517399 = $signed({1'h0, add_516963}) < $signed({1'h0, sel_516965}) ? add_516963 : sel_516965;
  assign add_517401 = array_index_514561[11:0] + 12'h97d;
  assign sel_517403 = $signed({1'h0, add_516967}) < $signed({1'h0, sel_516969}) ? add_516967 : sel_516969;
  assign add_517405 = array_index_514818[11:2] + 10'h2bb;
  assign sel_517408 = $signed({1'h0, add_516971, array_index_514558[1:0]}) < $signed({1'h0, sel_516974}) ? {add_516971, array_index_514558[1:0]} : sel_516974;
  assign add_517410 = array_index_514821[11:2] + 10'h2bb;
  assign sel_517413 = $signed({1'h0, add_516976, array_index_514561[1:0]}) < $signed({1'h0, sel_516979}) ? {add_516976, array_index_514561[1:0]} : sel_516979;
  assign add_517415 = array_index_515098[11:0] + 12'h8e1;
  assign sel_517417 = $signed({1'h0, add_516981}) < $signed({1'h0, sel_516983}) ? add_516981 : sel_516983;
  assign add_517419 = array_index_515101[11:0] + 12'h8e1;
  assign sel_517421 = $signed({1'h0, add_516985}) < $signed({1'h0, sel_516987}) ? add_516985 : sel_516987;
  assign add_517423 = array_index_515398[11:4] + 8'h83;
  assign sel_517426 = $signed({1'h0, add_516989, array_index_515098[3:0]}) < $signed({1'h0, sel_516992}) ? {add_516989, array_index_515098[3:0]} : sel_516992;
  assign add_517428 = array_index_515401[11:4] + 8'h83;
  assign sel_517431 = $signed({1'h0, add_516994, array_index_515101[3:0]}) < $signed({1'h0, sel_516997}) ? {add_516994, array_index_515101[3:0]} : sel_516997;
  assign add_517433 = array_index_515726[11:0] + 12'ha09;
  assign sel_517435 = $signed({1'h0, add_516999}) < $signed({1'h0, sel_517001}) ? add_516999 : sel_517001;
  assign add_517437 = array_index_515729[11:0] + 12'ha09;
  assign sel_517439 = $signed({1'h0, add_517003}) < $signed({1'h0, sel_517005}) ? add_517003 : sel_517005;
  assign add_517441 = array_index_516080[11:1] + 11'h6cb;
  assign sel_517443 = $signed({1'h0, add_517007, array_index_515726[0]}) < $signed({1'h0, sel_517009}) ? {add_517007, array_index_515726[0]} : sel_517009;
  assign add_517445 = array_index_516083[11:1] + 11'h6cb;
  assign sel_517447 = $signed({1'h0, add_517011, array_index_515729[0]}) < $signed({1'h0, sel_517013}) ? {add_517011, array_index_515729[0]} : sel_517013;
  assign add_517449 = array_index_516458[11:1] + 11'h75d;
  assign sel_517451 = $signed({1'h0, add_517015, array_index_516080[0]}) < $signed({1'h0, sel_517017}) ? {add_517015, array_index_516080[0]} : sel_517017;
  assign add_517453 = array_index_516461[11:1] + 11'h75d;
  assign sel_517455 = $signed({1'h0, add_517019, array_index_516083[0]}) < $signed({1'h0, sel_517021}) ? {add_517019, array_index_516083[0]} : sel_517021;
  assign add_517457 = array_index_516860[11:1] + 11'h24f;
  assign sel_517460 = $signed({1'h0, add_517023, array_index_516458[0]}) < $signed({1'h0, sel_517026}) ? {add_517023, array_index_516458[0]} : sel_517026;
  assign add_517462 = array_index_516863[11:1] + 11'h24f;
  assign sel_517465 = $signed({1'h0, add_517028, array_index_516461[0]}) < $signed({1'h0, sel_517031}) ? {add_517028, array_index_516461[0]} : sel_517031;
  assign add_517479 = array_index_512834[11:0] + 12'hbb1;
  assign sel_517481 = $signed({1'h0, add_517039}) < $signed(13'h0fff) ? add_517039 : 12'hfff;
  assign add_517483 = array_index_512837[11:0] + 12'hbb1;
  assign sel_517485 = $signed({1'h0, add_517041}) < $signed(13'h0fff) ? add_517041 : 12'hfff;
  assign add_517495 = array_index_512942[11:0] + 12'h6ab;
  assign sel_517497 = $signed({1'h0, add_517053}) < $signed({1'h0, sel_517055}) ? add_517053 : sel_517055;
  assign add_517499 = array_index_512945[11:0] + 12'h6ab;
  assign sel_517501 = $signed({1'h0, add_517057}) < $signed({1'h0, sel_517059}) ? add_517057 : sel_517059;
  assign add_517511 = array_index_513120[11:0] + 12'h7d5;
  assign sel_517513 = $signed({1'h0, add_517069}) < $signed({1'h0, sel_517071}) ? add_517069 : sel_517071;
  assign add_517515 = array_index_513123[11:0] + 12'h7d5;
  assign sel_517517 = $signed({1'h0, add_517073}) < $signed({1'h0, sel_517075}) ? add_517073 : sel_517075;
  assign add_517586 = array_index_517286[11:0] + 12'h62b;
  assign sel_517588 = $signed({1'h0, add_517144}) < $signed({1'h0, sel_517146}) ? add_517144 : sel_517146;
  assign add_517591 = array_index_517289[11:0] + 12'h62b;
  assign sel_517593 = $signed({1'h0, add_517149}) < $signed({1'h0, sel_517151}) ? add_517149 : sel_517151;
  assign add_517595 = array_index_512818[11:0] + 12'hcb1;
  assign add_517597 = array_index_512819[11:0] + 12'hcb1;
  assign add_517609 = array_index_512880[11:0] + 12'h81f;
  assign sel_517611 = $signed({1'h0, add_517159}) < $signed({1'h0, sel_517161}) ? add_517159 : sel_517161;
  assign add_517613 = array_index_512883[11:0] + 12'h81f;
  assign sel_517615 = $signed({1'h0, add_517163}) < $signed({1'h0, sel_517165}) ? add_517163 : sel_517165;
  assign add_517625 = array_index_513022[11:0] + 12'h45b;
  assign sel_517627 = $signed({1'h0, add_517175}) < $signed({1'h0, sel_517177}) ? add_517175 : sel_517177;
  assign add_517629 = array_index_513025[11:0] + 12'h45b;
  assign sel_517631 = $signed({1'h0, add_517179}) < $signed({1'h0, sel_517181}) ? add_517179 : sel_517181;
  assign add_517643 = array_index_513238[11:3] + 9'h0f5;
  assign sel_517645 = $signed({1'h0, add_517193, array_index_513120[2:0]}) < $signed({1'h0, sel_517195}) ? {add_517193, array_index_513120[2:0]} : sel_517195;
  assign add_517647 = array_index_513241[11:3] + 9'h0f5;
  assign sel_517649 = $signed({1'h0, add_517197, array_index_513123[2:0]}) < $signed({1'h0, sel_517199}) ? {add_517197, array_index_513123[2:0]} : sel_517199;
  assign array_index_517736 = set1_unflattened[5'h16];
  assign array_index_517739 = set2_unflattened[5'h16];
  assign add_517749 = array_index_512834[11:0] + 12'h437;
  assign sel_517751 = $signed({1'h0, add_517293}) < $signed(13'h0fff) ? add_517293 : 12'hfff;
  assign add_517753 = array_index_512837[11:0] + 12'h437;
  assign sel_517755 = $signed({1'h0, add_517295}) < $signed(13'h0fff) ? add_517295 : 12'hfff;
  assign add_517765 = array_index_512942[11:0] + 12'hee1;
  assign sel_517767 = $signed({1'h0, add_517307}) < $signed({1'h0, sel_517309}) ? add_517307 : sel_517309;
  assign add_517769 = array_index_512945[11:0] + 12'hee1;
  assign sel_517771 = $signed({1'h0, add_517311}) < $signed({1'h0, sel_517313}) ? add_517311 : sel_517313;
  assign add_517781 = array_index_513120[11:1] + 11'h179;
  assign sel_517783 = $signed({1'h0, add_517323, array_index_513022[0]}) < $signed({1'h0, sel_517325}) ? {add_517323, array_index_513022[0]} : sel_517325;
  assign add_517785 = array_index_513123[11:1] + 11'h179;
  assign sel_517787 = $signed({1'h0, add_517327, array_index_513025[0]}) < $signed({1'h0, sel_517329}) ? {add_517327, array_index_513025[0]} : sel_517329;
  assign add_517797 = array_index_513374[11:0] + 12'h067;
  assign sel_517799 = $signed({1'h0, add_517339}) < $signed({1'h0, sel_517341}) ? add_517339 : sel_517341;
  assign add_517801 = array_index_513377[11:0] + 12'h067;
  assign sel_517803 = $signed({1'h0, add_517343}) < $signed({1'h0, sel_517345}) ? add_517343 : sel_517345;
  assign add_517805 = array_index_513530[11:3] + 9'h1ef;
  assign sel_517808 = $signed({1'h0, add_517347, array_index_513374[2:0]}) < $signed({1'h0, sel_517350}) ? {add_517347, array_index_513374[2:0]} : sel_517350;
  assign add_517810 = array_index_513533[11:3] + 9'h1ef;
  assign sel_517813 = $signed({1'h0, add_517352, array_index_513377[2:0]}) < $signed({1'h0, sel_517355}) ? {add_517352, array_index_513377[2:0]} : sel_517355;
  assign add_517815 = array_index_513702[11:1] + 11'h2d5;
  assign sel_517817 = $signed({1'h0, add_517357, array_index_513530[0]}) < $signed({1'h0, sel_517359}) ? {add_517357, array_index_513530[0]} : sel_517359;
  assign add_517819 = array_index_513705[11:1] + 11'h2d5;
  assign sel_517821 = $signed({1'h0, add_517361, array_index_513533[0]}) < $signed({1'h0, sel_517363}) ? {add_517361, array_index_513533[0]} : sel_517363;
  assign add_517823 = array_index_513890[11:2] + 10'h353;
  assign sel_517825 = $signed({1'h0, add_517365, array_index_513702[1:0]}) < $signed({1'h0, sel_517367}) ? {add_517365, array_index_513702[1:0]} : sel_517367;
  assign add_517827 = array_index_513893[11:2] + 10'h353;
  assign sel_517829 = $signed({1'h0, add_517369, array_index_513705[1:0]}) < $signed({1'h0, sel_517371}) ? {add_517369, array_index_513705[1:0]} : sel_517371;
  assign add_517831 = array_index_514096[11:0] + 12'h0a7;
  assign sel_517833 = $signed({1'h0, add_517373}) < $signed({1'h0, sel_517375}) ? add_517373 : sel_517375;
  assign add_517835 = array_index_514099[11:0] + 12'h0a7;
  assign sel_517837 = $signed({1'h0, add_517377}) < $signed({1'h0, sel_517379}) ? add_517377 : sel_517379;
  assign add_517839 = array_index_514318[11:1] + 11'h4cb;
  assign sel_517841 = $signed({1'h0, add_517381, array_index_514096[0]}) < $signed({1'h0, sel_517383}) ? {add_517381, array_index_514096[0]} : sel_517383;
  assign add_517843 = array_index_514321[11:1] + 11'h4cb;
  assign sel_517845 = $signed({1'h0, add_517385, array_index_514099[0]}) < $signed({1'h0, sel_517387}) ? {add_517385, array_index_514099[0]} : sel_517387;
  assign add_517847 = array_index_514558[11:0] + 12'hfe9;
  assign sel_517849 = $signed({1'h0, add_517389}) < $signed({1'h0, sel_517391}) ? add_517389 : sel_517391;
  assign add_517851 = array_index_514561[11:0] + 12'hfe9;
  assign sel_517853 = $signed({1'h0, add_517393}) < $signed({1'h0, sel_517395}) ? add_517393 : sel_517395;
  assign add_517855 = array_index_514818[11:0] + 12'h97d;
  assign sel_517857 = $signed({1'h0, add_517397}) < $signed({1'h0, sel_517399}) ? add_517397 : sel_517399;
  assign add_517859 = array_index_514821[11:0] + 12'h97d;
  assign sel_517861 = $signed({1'h0, add_517401}) < $signed({1'h0, sel_517403}) ? add_517401 : sel_517403;
  assign add_517863 = array_index_515098[11:2] + 10'h2bb;
  assign sel_517866 = $signed({1'h0, add_517405, array_index_514818[1:0]}) < $signed({1'h0, sel_517408}) ? {add_517405, array_index_514818[1:0]} : sel_517408;
  assign add_517868 = array_index_515101[11:2] + 10'h2bb;
  assign sel_517871 = $signed({1'h0, add_517410, array_index_514821[1:0]}) < $signed({1'h0, sel_517413}) ? {add_517410, array_index_514821[1:0]} : sel_517413;
  assign add_517873 = array_index_515398[11:0] + 12'h8e1;
  assign sel_517875 = $signed({1'h0, add_517415}) < $signed({1'h0, sel_517417}) ? add_517415 : sel_517417;
  assign add_517877 = array_index_515401[11:0] + 12'h8e1;
  assign sel_517879 = $signed({1'h0, add_517419}) < $signed({1'h0, sel_517421}) ? add_517419 : sel_517421;
  assign add_517881 = array_index_515726[11:4] + 8'h83;
  assign sel_517884 = $signed({1'h0, add_517423, array_index_515398[3:0]}) < $signed({1'h0, sel_517426}) ? {add_517423, array_index_515398[3:0]} : sel_517426;
  assign add_517886 = array_index_515729[11:4] + 8'h83;
  assign sel_517889 = $signed({1'h0, add_517428, array_index_515401[3:0]}) < $signed({1'h0, sel_517431}) ? {add_517428, array_index_515401[3:0]} : sel_517431;
  assign add_517891 = array_index_516080[11:0] + 12'ha09;
  assign sel_517893 = $signed({1'h0, add_517433}) < $signed({1'h0, sel_517435}) ? add_517433 : sel_517435;
  assign add_517895 = array_index_516083[11:0] + 12'ha09;
  assign sel_517897 = $signed({1'h0, add_517437}) < $signed({1'h0, sel_517439}) ? add_517437 : sel_517439;
  assign add_517899 = array_index_516458[11:1] + 11'h6cb;
  assign sel_517901 = $signed({1'h0, add_517441, array_index_516080[0]}) < $signed({1'h0, sel_517443}) ? {add_517441, array_index_516080[0]} : sel_517443;
  assign add_517903 = array_index_516461[11:1] + 11'h6cb;
  assign sel_517905 = $signed({1'h0, add_517445, array_index_516083[0]}) < $signed({1'h0, sel_517447}) ? {add_517445, array_index_516083[0]} : sel_517447;
  assign add_517907 = array_index_516860[11:1] + 11'h75d;
  assign sel_517909 = $signed({1'h0, add_517449, array_index_516458[0]}) < $signed({1'h0, sel_517451}) ? {add_517449, array_index_516458[0]} : sel_517451;
  assign add_517911 = array_index_516863[11:1] + 11'h75d;
  assign sel_517913 = $signed({1'h0, add_517453, array_index_516461[0]}) < $signed({1'h0, sel_517455}) ? {add_517453, array_index_516461[0]} : sel_517455;
  assign add_517915 = array_index_517286[11:1] + 11'h24f;
  assign sel_517918 = $signed({1'h0, add_517457, array_index_516860[0]}) < $signed({1'h0, sel_517460}) ? {add_517457, array_index_516860[0]} : sel_517460;
  assign add_517920 = array_index_517289[11:1] + 11'h24f;
  assign sel_517923 = $signed({1'h0, add_517462, array_index_516863[0]}) < $signed({1'h0, sel_517465}) ? {add_517462, array_index_516863[0]} : sel_517465;
  assign add_517931 = array_index_512818[11:1] + 11'h4c1;
  assign add_517933 = array_index_512819[11:1] + 11'h4c1;
  assign add_517945 = array_index_512880[11:0] + 12'hbb1;
  assign sel_517947 = $signed({1'h0, add_517479}) < $signed({1'h0, sel_517481}) ? add_517479 : sel_517481;
  assign add_517949 = array_index_512883[11:0] + 12'hbb1;
  assign sel_517951 = $signed({1'h0, add_517483}) < $signed({1'h0, sel_517485}) ? add_517483 : sel_517485;
  assign add_517961 = array_index_513022[11:0] + 12'h6ab;
  assign sel_517963 = $signed({1'h0, add_517495}) < $signed({1'h0, sel_517497}) ? add_517495 : sel_517497;
  assign add_517965 = array_index_513025[11:0] + 12'h6ab;
  assign sel_517967 = $signed({1'h0, add_517499}) < $signed({1'h0, sel_517501}) ? add_517499 : sel_517501;
  assign add_517977 = array_index_513238[11:0] + 12'h7d5;
  assign sel_517979 = $signed({1'h0, add_517511}) < $signed({1'h0, sel_517513}) ? add_517511 : sel_517513;
  assign add_517981 = array_index_513241[11:0] + 12'h7d5;
  assign sel_517983 = $signed({1'h0, add_517515}) < $signed({1'h0, sel_517517}) ? add_517515 : sel_517517;
  assign add_518052 = array_index_517736[11:0] + 12'h62b;
  assign sel_518054 = $signed({1'h0, add_517586}) < $signed({1'h0, sel_517588}) ? add_517586 : sel_517588;
  assign add_518057 = array_index_517739[11:0] + 12'h62b;
  assign sel_518059 = $signed({1'h0, add_517591}) < $signed({1'h0, sel_517593}) ? add_517591 : sel_517593;
  assign add_518067 = array_index_512834[11:0] + 12'hcb1;
  assign sel_518069 = $signed({1'h0, add_517595}) < $signed(13'h0fff) ? add_517595 : 12'hfff;
  assign add_518071 = array_index_512837[11:0] + 12'hcb1;
  assign sel_518073 = $signed({1'h0, add_517597}) < $signed(13'h0fff) ? add_517597 : 12'hfff;
  assign add_518083 = array_index_512942[11:0] + 12'h81f;
  assign sel_518085 = $signed({1'h0, add_517609}) < $signed({1'h0, sel_517611}) ? add_517609 : sel_517611;
  assign add_518087 = array_index_512945[11:0] + 12'h81f;
  assign sel_518089 = $signed({1'h0, add_517613}) < $signed({1'h0, sel_517615}) ? add_517613 : sel_517615;
  assign add_518099 = array_index_513120[11:0] + 12'h45b;
  assign sel_518101 = $signed({1'h0, add_517625}) < $signed({1'h0, sel_517627}) ? add_517625 : sel_517627;
  assign add_518103 = array_index_513123[11:0] + 12'h45b;
  assign sel_518105 = $signed({1'h0, add_517629}) < $signed({1'h0, sel_517631}) ? add_517629 : sel_517631;
  assign add_518117 = array_index_513374[11:3] + 9'h0f5;
  assign sel_518119 = $signed({1'h0, add_517643, array_index_513238[2:0]}) < $signed({1'h0, sel_517645}) ? {add_517643, array_index_513238[2:0]} : sel_517645;
  assign add_518121 = array_index_513377[11:3] + 9'h0f5;
  assign sel_518123 = $signed({1'h0, add_517647, array_index_513241[2:0]}) < $signed({1'h0, sel_517649}) ? {add_517647, array_index_513241[2:0]} : sel_517649;
  assign array_index_518210 = set1_unflattened[5'h17];
  assign array_index_518213 = set2_unflattened[5'h17];
  assign add_518217 = array_index_512818[11:0] + 12'hf59;
  assign add_518219 = array_index_512819[11:0] + 12'hf59;
  assign add_518233 = array_index_512880[11:0] + 12'h437;
  assign sel_518235 = $signed({1'h0, add_517749}) < $signed({1'h0, sel_517751}) ? add_517749 : sel_517751;
  assign add_518237 = array_index_512883[11:0] + 12'h437;
  assign sel_518239 = $signed({1'h0, add_517753}) < $signed({1'h0, sel_517755}) ? add_517753 : sel_517755;
  assign add_518249 = array_index_513022[11:0] + 12'hee1;
  assign sel_518251 = $signed({1'h0, add_517765}) < $signed({1'h0, sel_517767}) ? add_517765 : sel_517767;
  assign add_518253 = array_index_513025[11:0] + 12'hee1;
  assign sel_518255 = $signed({1'h0, add_517769}) < $signed({1'h0, sel_517771}) ? add_517769 : sel_517771;
  assign add_518265 = array_index_513238[11:1] + 11'h179;
  assign sel_518267 = $signed({1'h0, add_517781, array_index_513120[0]}) < $signed({1'h0, sel_517783}) ? {add_517781, array_index_513120[0]} : sel_517783;
  assign add_518269 = array_index_513241[11:1] + 11'h179;
  assign sel_518271 = $signed({1'h0, add_517785, array_index_513123[0]}) < $signed({1'h0, sel_517787}) ? {add_517785, array_index_513123[0]} : sel_517787;
  assign add_518281 = array_index_513530[11:0] + 12'h067;
  assign sel_518283 = $signed({1'h0, add_517797}) < $signed({1'h0, sel_517799}) ? add_517797 : sel_517799;
  assign add_518285 = array_index_513533[11:0] + 12'h067;
  assign sel_518287 = $signed({1'h0, add_517801}) < $signed({1'h0, sel_517803}) ? add_517801 : sel_517803;
  assign add_518289 = array_index_513702[11:3] + 9'h1ef;
  assign sel_518292 = $signed({1'h0, add_517805, array_index_513530[2:0]}) < $signed({1'h0, sel_517808}) ? {add_517805, array_index_513530[2:0]} : sel_517808;
  assign add_518294 = array_index_513705[11:3] + 9'h1ef;
  assign sel_518297 = $signed({1'h0, add_517810, array_index_513533[2:0]}) < $signed({1'h0, sel_517813}) ? {add_517810, array_index_513533[2:0]} : sel_517813;
  assign add_518299 = array_index_513890[11:1] + 11'h2d5;
  assign sel_518301 = $signed({1'h0, add_517815, array_index_513702[0]}) < $signed({1'h0, sel_517817}) ? {add_517815, array_index_513702[0]} : sel_517817;
  assign add_518303 = array_index_513893[11:1] + 11'h2d5;
  assign sel_518305 = $signed({1'h0, add_517819, array_index_513705[0]}) < $signed({1'h0, sel_517821}) ? {add_517819, array_index_513705[0]} : sel_517821;
  assign add_518307 = array_index_514096[11:2] + 10'h353;
  assign sel_518309 = $signed({1'h0, add_517823, array_index_513890[1:0]}) < $signed({1'h0, sel_517825}) ? {add_517823, array_index_513890[1:0]} : sel_517825;
  assign add_518311 = array_index_514099[11:2] + 10'h353;
  assign sel_518313 = $signed({1'h0, add_517827, array_index_513893[1:0]}) < $signed({1'h0, sel_517829}) ? {add_517827, array_index_513893[1:0]} : sel_517829;
  assign add_518315 = array_index_514318[11:0] + 12'h0a7;
  assign sel_518317 = $signed({1'h0, add_517831}) < $signed({1'h0, sel_517833}) ? add_517831 : sel_517833;
  assign add_518319 = array_index_514321[11:0] + 12'h0a7;
  assign sel_518321 = $signed({1'h0, add_517835}) < $signed({1'h0, sel_517837}) ? add_517835 : sel_517837;
  assign add_518323 = array_index_514558[11:1] + 11'h4cb;
  assign sel_518325 = $signed({1'h0, add_517839, array_index_514318[0]}) < $signed({1'h0, sel_517841}) ? {add_517839, array_index_514318[0]} : sel_517841;
  assign add_518327 = array_index_514561[11:1] + 11'h4cb;
  assign sel_518329 = $signed({1'h0, add_517843, array_index_514321[0]}) < $signed({1'h0, sel_517845}) ? {add_517843, array_index_514321[0]} : sel_517845;
  assign add_518331 = array_index_514818[11:0] + 12'hfe9;
  assign sel_518333 = $signed({1'h0, add_517847}) < $signed({1'h0, sel_517849}) ? add_517847 : sel_517849;
  assign add_518335 = array_index_514821[11:0] + 12'hfe9;
  assign sel_518337 = $signed({1'h0, add_517851}) < $signed({1'h0, sel_517853}) ? add_517851 : sel_517853;
  assign add_518339 = array_index_515098[11:0] + 12'h97d;
  assign sel_518341 = $signed({1'h0, add_517855}) < $signed({1'h0, sel_517857}) ? add_517855 : sel_517857;
  assign add_518343 = array_index_515101[11:0] + 12'h97d;
  assign sel_518345 = $signed({1'h0, add_517859}) < $signed({1'h0, sel_517861}) ? add_517859 : sel_517861;
  assign add_518347 = array_index_515398[11:2] + 10'h2bb;
  assign sel_518350 = $signed({1'h0, add_517863, array_index_515098[1:0]}) < $signed({1'h0, sel_517866}) ? {add_517863, array_index_515098[1:0]} : sel_517866;
  assign add_518352 = array_index_515401[11:2] + 10'h2bb;
  assign sel_518355 = $signed({1'h0, add_517868, array_index_515101[1:0]}) < $signed({1'h0, sel_517871}) ? {add_517868, array_index_515101[1:0]} : sel_517871;
  assign add_518357 = array_index_515726[11:0] + 12'h8e1;
  assign sel_518359 = $signed({1'h0, add_517873}) < $signed({1'h0, sel_517875}) ? add_517873 : sel_517875;
  assign add_518361 = array_index_515729[11:0] + 12'h8e1;
  assign sel_518363 = $signed({1'h0, add_517877}) < $signed({1'h0, sel_517879}) ? add_517877 : sel_517879;
  assign add_518365 = array_index_516080[11:4] + 8'h83;
  assign sel_518368 = $signed({1'h0, add_517881, array_index_515726[3:0]}) < $signed({1'h0, sel_517884}) ? {add_517881, array_index_515726[3:0]} : sel_517884;
  assign add_518370 = array_index_516083[11:4] + 8'h83;
  assign sel_518373 = $signed({1'h0, add_517886, array_index_515729[3:0]}) < $signed({1'h0, sel_517889}) ? {add_517886, array_index_515729[3:0]} : sel_517889;
  assign add_518375 = array_index_516458[11:0] + 12'ha09;
  assign sel_518377 = $signed({1'h0, add_517891}) < $signed({1'h0, sel_517893}) ? add_517891 : sel_517893;
  assign add_518379 = array_index_516461[11:0] + 12'ha09;
  assign sel_518381 = $signed({1'h0, add_517895}) < $signed({1'h0, sel_517897}) ? add_517895 : sel_517897;
  assign add_518383 = array_index_516860[11:1] + 11'h6cb;
  assign sel_518385 = $signed({1'h0, add_517899, array_index_516458[0]}) < $signed({1'h0, sel_517901}) ? {add_517899, array_index_516458[0]} : sel_517901;
  assign add_518387 = array_index_516863[11:1] + 11'h6cb;
  assign sel_518389 = $signed({1'h0, add_517903, array_index_516461[0]}) < $signed({1'h0, sel_517905}) ? {add_517903, array_index_516461[0]} : sel_517905;
  assign add_518391 = array_index_517286[11:1] + 11'h75d;
  assign sel_518393 = $signed({1'h0, add_517907, array_index_516860[0]}) < $signed({1'h0, sel_517909}) ? {add_517907, array_index_516860[0]} : sel_517909;
  assign add_518395 = array_index_517289[11:1] + 11'h75d;
  assign sel_518397 = $signed({1'h0, add_517911, array_index_516863[0]}) < $signed({1'h0, sel_517913}) ? {add_517911, array_index_516863[0]} : sel_517913;
  assign add_518399 = array_index_517736[11:1] + 11'h24f;
  assign sel_518402 = $signed({1'h0, add_517915, array_index_517286[0]}) < $signed({1'h0, sel_517918}) ? {add_517915, array_index_517286[0]} : sel_517918;
  assign add_518404 = array_index_517739[11:1] + 11'h24f;
  assign sel_518407 = $signed({1'h0, add_517920, array_index_517289[0]}) < $signed({1'h0, sel_517923}) ? {add_517920, array_index_517289[0]} : sel_517923;
  assign add_518421 = array_index_512834[11:1] + 11'h4c1;
  assign sel_518423 = $signed({1'h0, add_517931, array_index_512818[0]}) < $signed(13'h0fff) ? {add_517931, array_index_512818[0]} : 12'hfff;
  assign add_518425 = array_index_512837[11:1] + 11'h4c1;
  assign sel_518427 = $signed({1'h0, add_517933, array_index_512819[0]}) < $signed(13'h0fff) ? {add_517933, array_index_512819[0]} : 12'hfff;
  assign add_518437 = array_index_512942[11:0] + 12'hbb1;
  assign sel_518439 = $signed({1'h0, add_517945}) < $signed({1'h0, sel_517947}) ? add_517945 : sel_517947;
  assign add_518441 = array_index_512945[11:0] + 12'hbb1;
  assign sel_518443 = $signed({1'h0, add_517949}) < $signed({1'h0, sel_517951}) ? add_517949 : sel_517951;
  assign add_518453 = array_index_513120[11:0] + 12'h6ab;
  assign sel_518455 = $signed({1'h0, add_517961}) < $signed({1'h0, sel_517963}) ? add_517961 : sel_517963;
  assign add_518457 = array_index_513123[11:0] + 12'h6ab;
  assign sel_518459 = $signed({1'h0, add_517965}) < $signed({1'h0, sel_517967}) ? add_517965 : sel_517967;
  assign add_518469 = array_index_513374[11:0] + 12'h7d5;
  assign sel_518471 = $signed({1'h0, add_517977}) < $signed({1'h0, sel_517979}) ? add_517977 : sel_517979;
  assign add_518473 = array_index_513377[11:0] + 12'h7d5;
  assign sel_518475 = $signed({1'h0, add_517981}) < $signed({1'h0, sel_517983}) ? add_517981 : sel_517983;
  assign add_518544 = array_index_518210[11:0] + 12'h62b;
  assign sel_518546 = $signed({1'h0, add_518052}) < $signed({1'h0, sel_518054}) ? add_518052 : sel_518054;
  assign add_518549 = array_index_518213[11:0] + 12'h62b;
  assign sel_518551 = $signed({1'h0, add_518057}) < $signed({1'h0, sel_518059}) ? add_518057 : sel_518059;
  assign add_518553 = array_index_512818[11:1] + 11'h44d;
  assign add_518555 = array_index_512819[11:1] + 11'h44d;
  assign add_518567 = array_index_512880[11:0] + 12'hcb1;
  assign sel_518569 = $signed({1'h0, add_518067}) < $signed({1'h0, sel_518069}) ? add_518067 : sel_518069;
  assign add_518571 = array_index_512883[11:0] + 12'hcb1;
  assign sel_518573 = $signed({1'h0, add_518071}) < $signed({1'h0, sel_518073}) ? add_518071 : sel_518073;
  assign add_518583 = array_index_513022[11:0] + 12'h81f;
  assign sel_518585 = $signed({1'h0, add_518083}) < $signed({1'h0, sel_518085}) ? add_518083 : sel_518085;
  assign add_518587 = array_index_513025[11:0] + 12'h81f;
  assign sel_518589 = $signed({1'h0, add_518087}) < $signed({1'h0, sel_518089}) ? add_518087 : sel_518089;
  assign add_518599 = array_index_513238[11:0] + 12'h45b;
  assign sel_518601 = $signed({1'h0, add_518099}) < $signed({1'h0, sel_518101}) ? add_518099 : sel_518101;
  assign add_518603 = array_index_513241[11:0] + 12'h45b;
  assign sel_518605 = $signed({1'h0, add_518103}) < $signed({1'h0, sel_518105}) ? add_518103 : sel_518105;
  assign add_518617 = array_index_513530[11:3] + 9'h0f5;
  assign sel_518619 = $signed({1'h0, add_518117, array_index_513374[2:0]}) < $signed({1'h0, sel_518119}) ? {add_518117, array_index_513374[2:0]} : sel_518119;
  assign add_518621 = array_index_513533[11:3] + 9'h0f5;
  assign sel_518623 = $signed({1'h0, add_518121, array_index_513377[2:0]}) < $signed({1'h0, sel_518123}) ? {add_518121, array_index_513377[2:0]} : sel_518123;
  assign array_index_518710 = set1_unflattened[5'h18];
  assign array_index_518713 = set2_unflattened[5'h18];
  assign add_518723 = array_index_512834[11:0] + 12'hf59;
  assign sel_518725 = $signed({1'h0, add_518217}) < $signed(13'h0fff) ? add_518217 : 12'hfff;
  assign add_518727 = array_index_512837[11:0] + 12'hf59;
  assign sel_518729 = $signed({1'h0, add_518219}) < $signed(13'h0fff) ? add_518219 : 12'hfff;
  assign add_518741 = array_index_512942[11:0] + 12'h437;
  assign sel_518743 = $signed({1'h0, add_518233}) < $signed({1'h0, sel_518235}) ? add_518233 : sel_518235;
  assign add_518745 = array_index_512945[11:0] + 12'h437;
  assign sel_518747 = $signed({1'h0, add_518237}) < $signed({1'h0, sel_518239}) ? add_518237 : sel_518239;
  assign add_518757 = array_index_513120[11:0] + 12'hee1;
  assign sel_518759 = $signed({1'h0, add_518249}) < $signed({1'h0, sel_518251}) ? add_518249 : sel_518251;
  assign add_518761 = array_index_513123[11:0] + 12'hee1;
  assign sel_518763 = $signed({1'h0, add_518253}) < $signed({1'h0, sel_518255}) ? add_518253 : sel_518255;
  assign add_518773 = array_index_513374[11:1] + 11'h179;
  assign sel_518775 = $signed({1'h0, add_518265, array_index_513238[0]}) < $signed({1'h0, sel_518267}) ? {add_518265, array_index_513238[0]} : sel_518267;
  assign add_518777 = array_index_513377[11:1] + 11'h179;
  assign sel_518779 = $signed({1'h0, add_518269, array_index_513241[0]}) < $signed({1'h0, sel_518271}) ? {add_518269, array_index_513241[0]} : sel_518271;
  assign add_518789 = array_index_513702[11:0] + 12'h067;
  assign sel_518791 = $signed({1'h0, add_518281}) < $signed({1'h0, sel_518283}) ? add_518281 : sel_518283;
  assign add_518793 = array_index_513705[11:0] + 12'h067;
  assign sel_518795 = $signed({1'h0, add_518285}) < $signed({1'h0, sel_518287}) ? add_518285 : sel_518287;
  assign add_518797 = array_index_513890[11:3] + 9'h1ef;
  assign sel_518800 = $signed({1'h0, add_518289, array_index_513702[2:0]}) < $signed({1'h0, sel_518292}) ? {add_518289, array_index_513702[2:0]} : sel_518292;
  assign add_518802 = array_index_513893[11:3] + 9'h1ef;
  assign sel_518805 = $signed({1'h0, add_518294, array_index_513705[2:0]}) < $signed({1'h0, sel_518297}) ? {add_518294, array_index_513705[2:0]} : sel_518297;
  assign add_518807 = array_index_514096[11:1] + 11'h2d5;
  assign sel_518809 = $signed({1'h0, add_518299, array_index_513890[0]}) < $signed({1'h0, sel_518301}) ? {add_518299, array_index_513890[0]} : sel_518301;
  assign add_518811 = array_index_514099[11:1] + 11'h2d5;
  assign sel_518813 = $signed({1'h0, add_518303, array_index_513893[0]}) < $signed({1'h0, sel_518305}) ? {add_518303, array_index_513893[0]} : sel_518305;
  assign add_518815 = array_index_514318[11:2] + 10'h353;
  assign sel_518817 = $signed({1'h0, add_518307, array_index_514096[1:0]}) < $signed({1'h0, sel_518309}) ? {add_518307, array_index_514096[1:0]} : sel_518309;
  assign add_518819 = array_index_514321[11:2] + 10'h353;
  assign sel_518821 = $signed({1'h0, add_518311, array_index_514099[1:0]}) < $signed({1'h0, sel_518313}) ? {add_518311, array_index_514099[1:0]} : sel_518313;
  assign add_518823 = array_index_514558[11:0] + 12'h0a7;
  assign sel_518825 = $signed({1'h0, add_518315}) < $signed({1'h0, sel_518317}) ? add_518315 : sel_518317;
  assign add_518827 = array_index_514561[11:0] + 12'h0a7;
  assign sel_518829 = $signed({1'h0, add_518319}) < $signed({1'h0, sel_518321}) ? add_518319 : sel_518321;
  assign add_518831 = array_index_514818[11:1] + 11'h4cb;
  assign sel_518833 = $signed({1'h0, add_518323, array_index_514558[0]}) < $signed({1'h0, sel_518325}) ? {add_518323, array_index_514558[0]} : sel_518325;
  assign add_518835 = array_index_514821[11:1] + 11'h4cb;
  assign sel_518837 = $signed({1'h0, add_518327, array_index_514561[0]}) < $signed({1'h0, sel_518329}) ? {add_518327, array_index_514561[0]} : sel_518329;
  assign add_518839 = array_index_515098[11:0] + 12'hfe9;
  assign sel_518841 = $signed({1'h0, add_518331}) < $signed({1'h0, sel_518333}) ? add_518331 : sel_518333;
  assign add_518843 = array_index_515101[11:0] + 12'hfe9;
  assign sel_518845 = $signed({1'h0, add_518335}) < $signed({1'h0, sel_518337}) ? add_518335 : sel_518337;
  assign add_518847 = array_index_515398[11:0] + 12'h97d;
  assign sel_518849 = $signed({1'h0, add_518339}) < $signed({1'h0, sel_518341}) ? add_518339 : sel_518341;
  assign add_518851 = array_index_515401[11:0] + 12'h97d;
  assign sel_518853 = $signed({1'h0, add_518343}) < $signed({1'h0, sel_518345}) ? add_518343 : sel_518345;
  assign add_518855 = array_index_515726[11:2] + 10'h2bb;
  assign sel_518858 = $signed({1'h0, add_518347, array_index_515398[1:0]}) < $signed({1'h0, sel_518350}) ? {add_518347, array_index_515398[1:0]} : sel_518350;
  assign add_518860 = array_index_515729[11:2] + 10'h2bb;
  assign sel_518863 = $signed({1'h0, add_518352, array_index_515401[1:0]}) < $signed({1'h0, sel_518355}) ? {add_518352, array_index_515401[1:0]} : sel_518355;
  assign add_518865 = array_index_516080[11:0] + 12'h8e1;
  assign sel_518867 = $signed({1'h0, add_518357}) < $signed({1'h0, sel_518359}) ? add_518357 : sel_518359;
  assign add_518869 = array_index_516083[11:0] + 12'h8e1;
  assign sel_518871 = $signed({1'h0, add_518361}) < $signed({1'h0, sel_518363}) ? add_518361 : sel_518363;
  assign add_518873 = array_index_516458[11:4] + 8'h83;
  assign sel_518876 = $signed({1'h0, add_518365, array_index_516080[3:0]}) < $signed({1'h0, sel_518368}) ? {add_518365, array_index_516080[3:0]} : sel_518368;
  assign add_518878 = array_index_516461[11:4] + 8'h83;
  assign sel_518881 = $signed({1'h0, add_518370, array_index_516083[3:0]}) < $signed({1'h0, sel_518373}) ? {add_518370, array_index_516083[3:0]} : sel_518373;
  assign add_518883 = array_index_516860[11:0] + 12'ha09;
  assign sel_518885 = $signed({1'h0, add_518375}) < $signed({1'h0, sel_518377}) ? add_518375 : sel_518377;
  assign add_518887 = array_index_516863[11:0] + 12'ha09;
  assign sel_518889 = $signed({1'h0, add_518379}) < $signed({1'h0, sel_518381}) ? add_518379 : sel_518381;
  assign add_518891 = array_index_517286[11:1] + 11'h6cb;
  assign sel_518893 = $signed({1'h0, add_518383, array_index_516860[0]}) < $signed({1'h0, sel_518385}) ? {add_518383, array_index_516860[0]} : sel_518385;
  assign add_518895 = array_index_517289[11:1] + 11'h6cb;
  assign sel_518897 = $signed({1'h0, add_518387, array_index_516863[0]}) < $signed({1'h0, sel_518389}) ? {add_518387, array_index_516863[0]} : sel_518389;
  assign add_518899 = array_index_517736[11:1] + 11'h75d;
  assign sel_518901 = $signed({1'h0, add_518391, array_index_517286[0]}) < $signed({1'h0, sel_518393}) ? {add_518391, array_index_517286[0]} : sel_518393;
  assign add_518903 = array_index_517739[11:1] + 11'h75d;
  assign sel_518905 = $signed({1'h0, add_518395, array_index_517289[0]}) < $signed({1'h0, sel_518397}) ? {add_518395, array_index_517289[0]} : sel_518397;
  assign add_518907 = array_index_518210[11:1] + 11'h24f;
  assign sel_518910 = $signed({1'h0, add_518399, array_index_517736[0]}) < $signed({1'h0, sel_518402}) ? {add_518399, array_index_517736[0]} : sel_518402;
  assign add_518912 = array_index_518213[11:1] + 11'h24f;
  assign sel_518915 = $signed({1'h0, add_518404, array_index_517739[0]}) < $signed({1'h0, sel_518407}) ? {add_518404, array_index_517739[0]} : sel_518407;
  assign add_518923 = array_index_512818[11:0] + 12'h0b1;
  assign add_518925 = array_index_512819[11:0] + 12'h0b1;
  assign add_518939 = array_index_512880[11:1] + 11'h4c1;
  assign sel_518941 = $signed({1'h0, add_518421, array_index_512834[0]}) < $signed({1'h0, sel_518423}) ? {add_518421, array_index_512834[0]} : sel_518423;
  assign add_518943 = array_index_512883[11:1] + 11'h4c1;
  assign sel_518945 = $signed({1'h0, add_518425, array_index_512837[0]}) < $signed({1'h0, sel_518427}) ? {add_518425, array_index_512837[0]} : sel_518427;
  assign add_518955 = array_index_513022[11:0] + 12'hbb1;
  assign sel_518957 = $signed({1'h0, add_518437}) < $signed({1'h0, sel_518439}) ? add_518437 : sel_518439;
  assign add_518959 = array_index_513025[11:0] + 12'hbb1;
  assign sel_518961 = $signed({1'h0, add_518441}) < $signed({1'h0, sel_518443}) ? add_518441 : sel_518443;
  assign add_518971 = array_index_513238[11:0] + 12'h6ab;
  assign sel_518973 = $signed({1'h0, add_518453}) < $signed({1'h0, sel_518455}) ? add_518453 : sel_518455;
  assign add_518975 = array_index_513241[11:0] + 12'h6ab;
  assign sel_518977 = $signed({1'h0, add_518457}) < $signed({1'h0, sel_518459}) ? add_518457 : sel_518459;
  assign add_518987 = array_index_513530[11:0] + 12'h7d5;
  assign sel_518989 = $signed({1'h0, add_518469}) < $signed({1'h0, sel_518471}) ? add_518469 : sel_518471;
  assign add_518991 = array_index_513533[11:0] + 12'h7d5;
  assign sel_518993 = $signed({1'h0, add_518473}) < $signed({1'h0, sel_518475}) ? add_518473 : sel_518475;
  assign add_519062 = array_index_518710[11:0] + 12'h62b;
  assign sel_519064 = $signed({1'h0, add_518544}) < $signed({1'h0, sel_518546}) ? add_518544 : sel_518546;
  assign add_519067 = array_index_518713[11:0] + 12'h62b;
  assign sel_519069 = $signed({1'h0, add_518549}) < $signed({1'h0, sel_518551}) ? add_518549 : sel_518551;
  assign add_519077 = array_index_512834[11:1] + 11'h44d;
  assign sel_519079 = $signed({1'h0, add_518553, array_index_512818[0]}) < $signed(13'h0fff) ? {add_518553, array_index_512818[0]} : 12'hfff;
  assign add_519081 = array_index_512837[11:1] + 11'h44d;
  assign sel_519083 = $signed({1'h0, add_518555, array_index_512819[0]}) < $signed(13'h0fff) ? {add_518555, array_index_512819[0]} : 12'hfff;
  assign add_519093 = array_index_512942[11:0] + 12'hcb1;
  assign sel_519095 = $signed({1'h0, add_518567}) < $signed({1'h0, sel_518569}) ? add_518567 : sel_518569;
  assign add_519097 = array_index_512945[11:0] + 12'hcb1;
  assign sel_519099 = $signed({1'h0, add_518571}) < $signed({1'h0, sel_518573}) ? add_518571 : sel_518573;
  assign add_519109 = array_index_513120[11:0] + 12'h81f;
  assign sel_519111 = $signed({1'h0, add_518583}) < $signed({1'h0, sel_518585}) ? add_518583 : sel_518585;
  assign add_519113 = array_index_513123[11:0] + 12'h81f;
  assign sel_519115 = $signed({1'h0, add_518587}) < $signed({1'h0, sel_518589}) ? add_518587 : sel_518589;
  assign add_519125 = array_index_513374[11:0] + 12'h45b;
  assign sel_519127 = $signed({1'h0, add_518599}) < $signed({1'h0, sel_518601}) ? add_518599 : sel_518601;
  assign add_519129 = array_index_513377[11:0] + 12'h45b;
  assign sel_519131 = $signed({1'h0, add_518603}) < $signed({1'h0, sel_518605}) ? add_518603 : sel_518605;
  assign add_519143 = array_index_513702[11:3] + 9'h0f5;
  assign sel_519145 = $signed({1'h0, add_518617, array_index_513530[2:0]}) < $signed({1'h0, sel_518619}) ? {add_518617, array_index_513530[2:0]} : sel_518619;
  assign add_519147 = array_index_513705[11:3] + 9'h0f5;
  assign sel_519149 = $signed({1'h0, add_518621, array_index_513533[2:0]}) < $signed({1'h0, sel_518623}) ? {add_518621, array_index_513533[2:0]} : sel_518623;
  assign array_index_519236 = set1_unflattened[5'h19];
  assign array_index_519239 = set2_unflattened[5'h19];
  assign add_519243 = array_index_512818[11:0] + 12'h091;
  assign add_519245 = array_index_512819[11:0] + 12'h091;
  assign add_519257 = array_index_512880[11:0] + 12'hf59;
  assign sel_519259 = $signed({1'h0, add_518723}) < $signed({1'h0, sel_518725}) ? add_518723 : sel_518725;
  assign add_519261 = array_index_512883[11:0] + 12'hf59;
  assign sel_519263 = $signed({1'h0, add_518727}) < $signed({1'h0, sel_518729}) ? add_518727 : sel_518729;
  assign add_519275 = array_index_513022[11:0] + 12'h437;
  assign sel_519277 = $signed({1'h0, add_518741}) < $signed({1'h0, sel_518743}) ? add_518741 : sel_518743;
  assign add_519279 = array_index_513025[11:0] + 12'h437;
  assign sel_519281 = $signed({1'h0, add_518745}) < $signed({1'h0, sel_518747}) ? add_518745 : sel_518747;
  assign add_519291 = array_index_513238[11:0] + 12'hee1;
  assign sel_519293 = $signed({1'h0, add_518757}) < $signed({1'h0, sel_518759}) ? add_518757 : sel_518759;
  assign add_519295 = array_index_513241[11:0] + 12'hee1;
  assign sel_519297 = $signed({1'h0, add_518761}) < $signed({1'h0, sel_518763}) ? add_518761 : sel_518763;
  assign add_519307 = array_index_513530[11:1] + 11'h179;
  assign sel_519309 = $signed({1'h0, add_518773, array_index_513374[0]}) < $signed({1'h0, sel_518775}) ? {add_518773, array_index_513374[0]} : sel_518775;
  assign add_519311 = array_index_513533[11:1] + 11'h179;
  assign sel_519313 = $signed({1'h0, add_518777, array_index_513377[0]}) < $signed({1'h0, sel_518779}) ? {add_518777, array_index_513377[0]} : sel_518779;
  assign add_519323 = array_index_513890[11:0] + 12'h067;
  assign sel_519325 = $signed({1'h0, add_518789}) < $signed({1'h0, sel_518791}) ? add_518789 : sel_518791;
  assign add_519327 = array_index_513893[11:0] + 12'h067;
  assign sel_519329 = $signed({1'h0, add_518793}) < $signed({1'h0, sel_518795}) ? add_518793 : sel_518795;
  assign add_519331 = array_index_514096[11:3] + 9'h1ef;
  assign sel_519334 = $signed({1'h0, add_518797, array_index_513890[2:0]}) < $signed({1'h0, sel_518800}) ? {add_518797, array_index_513890[2:0]} : sel_518800;
  assign add_519336 = array_index_514099[11:3] + 9'h1ef;
  assign sel_519339 = $signed({1'h0, add_518802, array_index_513893[2:0]}) < $signed({1'h0, sel_518805}) ? {add_518802, array_index_513893[2:0]} : sel_518805;
  assign add_519341 = array_index_514318[11:1] + 11'h2d5;
  assign sel_519343 = $signed({1'h0, add_518807, array_index_514096[0]}) < $signed({1'h0, sel_518809}) ? {add_518807, array_index_514096[0]} : sel_518809;
  assign add_519345 = array_index_514321[11:1] + 11'h2d5;
  assign sel_519347 = $signed({1'h0, add_518811, array_index_514099[0]}) < $signed({1'h0, sel_518813}) ? {add_518811, array_index_514099[0]} : sel_518813;
  assign add_519349 = array_index_514558[11:2] + 10'h353;
  assign sel_519351 = $signed({1'h0, add_518815, array_index_514318[1:0]}) < $signed({1'h0, sel_518817}) ? {add_518815, array_index_514318[1:0]} : sel_518817;
  assign add_519353 = array_index_514561[11:2] + 10'h353;
  assign sel_519355 = $signed({1'h0, add_518819, array_index_514321[1:0]}) < $signed({1'h0, sel_518821}) ? {add_518819, array_index_514321[1:0]} : sel_518821;
  assign add_519357 = array_index_514818[11:0] + 12'h0a7;
  assign sel_519359 = $signed({1'h0, add_518823}) < $signed({1'h0, sel_518825}) ? add_518823 : sel_518825;
  assign add_519361 = array_index_514821[11:0] + 12'h0a7;
  assign sel_519363 = $signed({1'h0, add_518827}) < $signed({1'h0, sel_518829}) ? add_518827 : sel_518829;
  assign add_519365 = array_index_515098[11:1] + 11'h4cb;
  assign sel_519367 = $signed({1'h0, add_518831, array_index_514818[0]}) < $signed({1'h0, sel_518833}) ? {add_518831, array_index_514818[0]} : sel_518833;
  assign add_519369 = array_index_515101[11:1] + 11'h4cb;
  assign sel_519371 = $signed({1'h0, add_518835, array_index_514821[0]}) < $signed({1'h0, sel_518837}) ? {add_518835, array_index_514821[0]} : sel_518837;
  assign add_519373 = array_index_515398[11:0] + 12'hfe9;
  assign sel_519375 = $signed({1'h0, add_518839}) < $signed({1'h0, sel_518841}) ? add_518839 : sel_518841;
  assign add_519377 = array_index_515401[11:0] + 12'hfe9;
  assign sel_519379 = $signed({1'h0, add_518843}) < $signed({1'h0, sel_518845}) ? add_518843 : sel_518845;
  assign add_519381 = array_index_515726[11:0] + 12'h97d;
  assign sel_519383 = $signed({1'h0, add_518847}) < $signed({1'h0, sel_518849}) ? add_518847 : sel_518849;
  assign add_519385 = array_index_515729[11:0] + 12'h97d;
  assign sel_519387 = $signed({1'h0, add_518851}) < $signed({1'h0, sel_518853}) ? add_518851 : sel_518853;
  assign add_519389 = array_index_516080[11:2] + 10'h2bb;
  assign sel_519392 = $signed({1'h0, add_518855, array_index_515726[1:0]}) < $signed({1'h0, sel_518858}) ? {add_518855, array_index_515726[1:0]} : sel_518858;
  assign add_519394 = array_index_516083[11:2] + 10'h2bb;
  assign sel_519397 = $signed({1'h0, add_518860, array_index_515729[1:0]}) < $signed({1'h0, sel_518863}) ? {add_518860, array_index_515729[1:0]} : sel_518863;
  assign add_519399 = array_index_516458[11:0] + 12'h8e1;
  assign sel_519401 = $signed({1'h0, add_518865}) < $signed({1'h0, sel_518867}) ? add_518865 : sel_518867;
  assign add_519403 = array_index_516461[11:0] + 12'h8e1;
  assign sel_519405 = $signed({1'h0, add_518869}) < $signed({1'h0, sel_518871}) ? add_518869 : sel_518871;
  assign add_519407 = array_index_516860[11:4] + 8'h83;
  assign sel_519410 = $signed({1'h0, add_518873, array_index_516458[3:0]}) < $signed({1'h0, sel_518876}) ? {add_518873, array_index_516458[3:0]} : sel_518876;
  assign add_519412 = array_index_516863[11:4] + 8'h83;
  assign sel_519415 = $signed({1'h0, add_518878, array_index_516461[3:0]}) < $signed({1'h0, sel_518881}) ? {add_518878, array_index_516461[3:0]} : sel_518881;
  assign add_519417 = array_index_517286[11:0] + 12'ha09;
  assign sel_519419 = $signed({1'h0, add_518883}) < $signed({1'h0, sel_518885}) ? add_518883 : sel_518885;
  assign add_519421 = array_index_517289[11:0] + 12'ha09;
  assign sel_519423 = $signed({1'h0, add_518887}) < $signed({1'h0, sel_518889}) ? add_518887 : sel_518889;
  assign add_519425 = array_index_517736[11:1] + 11'h6cb;
  assign sel_519427 = $signed({1'h0, add_518891, array_index_517286[0]}) < $signed({1'h0, sel_518893}) ? {add_518891, array_index_517286[0]} : sel_518893;
  assign add_519429 = array_index_517739[11:1] + 11'h6cb;
  assign sel_519431 = $signed({1'h0, add_518895, array_index_517289[0]}) < $signed({1'h0, sel_518897}) ? {add_518895, array_index_517289[0]} : sel_518897;
  assign add_519433 = array_index_518210[11:1] + 11'h75d;
  assign sel_519435 = $signed({1'h0, add_518899, array_index_517736[0]}) < $signed({1'h0, sel_518901}) ? {add_518899, array_index_517736[0]} : sel_518901;
  assign add_519437 = array_index_518213[11:1] + 11'h75d;
  assign sel_519439 = $signed({1'h0, add_518903, array_index_517739[0]}) < $signed({1'h0, sel_518905}) ? {add_518903, array_index_517739[0]} : sel_518905;
  assign add_519441 = array_index_518710[11:1] + 11'h24f;
  assign sel_519444 = $signed({1'h0, add_518907, array_index_518210[0]}) < $signed({1'h0, sel_518910}) ? {add_518907, array_index_518210[0]} : sel_518910;
  assign add_519446 = array_index_518713[11:1] + 11'h24f;
  assign sel_519449 = $signed({1'h0, add_518912, array_index_518213[0]}) < $signed({1'h0, sel_518915}) ? {add_518912, array_index_518213[0]} : sel_518915;
  assign add_519463 = array_index_512834[11:0] + 12'h0b1;
  assign sel_519465 = $signed({1'h0, add_518923}) < $signed(13'h0fff) ? add_518923 : 12'hfff;
  assign add_519467 = array_index_512837[11:0] + 12'h0b1;
  assign sel_519469 = $signed({1'h0, add_518925}) < $signed(13'h0fff) ? add_518925 : 12'hfff;
  assign add_519481 = array_index_512942[11:1] + 11'h4c1;
  assign sel_519483 = $signed({1'h0, add_518939, array_index_512880[0]}) < $signed({1'h0, sel_518941}) ? {add_518939, array_index_512880[0]} : sel_518941;
  assign add_519485 = array_index_512945[11:1] + 11'h4c1;
  assign sel_519487 = $signed({1'h0, add_518943, array_index_512883[0]}) < $signed({1'h0, sel_518945}) ? {add_518943, array_index_512883[0]} : sel_518945;
  assign add_519497 = array_index_513120[11:0] + 12'hbb1;
  assign sel_519499 = $signed({1'h0, add_518955}) < $signed({1'h0, sel_518957}) ? add_518955 : sel_518957;
  assign add_519501 = array_index_513123[11:0] + 12'hbb1;
  assign sel_519503 = $signed({1'h0, add_518959}) < $signed({1'h0, sel_518961}) ? add_518959 : sel_518961;
  assign add_519513 = array_index_513374[11:0] + 12'h6ab;
  assign sel_519515 = $signed({1'h0, add_518971}) < $signed({1'h0, sel_518973}) ? add_518971 : sel_518973;
  assign add_519517 = array_index_513377[11:0] + 12'h6ab;
  assign sel_519519 = $signed({1'h0, add_518975}) < $signed({1'h0, sel_518977}) ? add_518975 : sel_518977;
  assign add_519529 = array_index_513702[11:0] + 12'h7d5;
  assign sel_519531 = $signed({1'h0, add_518987}) < $signed({1'h0, sel_518989}) ? add_518987 : sel_518989;
  assign add_519533 = array_index_513705[11:0] + 12'h7d5;
  assign sel_519535 = $signed({1'h0, add_518991}) < $signed({1'h0, sel_518993}) ? add_518991 : sel_518993;
  assign add_519604 = array_index_519236[11:0] + 12'h62b;
  assign sel_519606 = $signed({1'h0, add_519062}) < $signed({1'h0, sel_519064}) ? add_519062 : sel_519064;
  assign add_519609 = array_index_519239[11:0] + 12'h62b;
  assign sel_519611 = $signed({1'h0, add_519067}) < $signed({1'h0, sel_519069}) ? add_519067 : sel_519069;
  assign add_519613 = array_index_512818[11:1] + 11'h283;
  assign add_519615 = array_index_512819[11:1] + 11'h283;
  assign add_519627 = array_index_512880[11:1] + 11'h44d;
  assign sel_519629 = $signed({1'h0, add_519077, array_index_512834[0]}) < $signed({1'h0, sel_519079}) ? {add_519077, array_index_512834[0]} : sel_519079;
  assign add_519631 = array_index_512883[11:1] + 11'h44d;
  assign sel_519633 = $signed({1'h0, add_519081, array_index_512837[0]}) < $signed({1'h0, sel_519083}) ? {add_519081, array_index_512837[0]} : sel_519083;
  assign add_519643 = array_index_513022[11:0] + 12'hcb1;
  assign sel_519645 = $signed({1'h0, add_519093}) < $signed({1'h0, sel_519095}) ? add_519093 : sel_519095;
  assign add_519647 = array_index_513025[11:0] + 12'hcb1;
  assign sel_519649 = $signed({1'h0, add_519097}) < $signed({1'h0, sel_519099}) ? add_519097 : sel_519099;
  assign add_519659 = array_index_513238[11:0] + 12'h81f;
  assign sel_519661 = $signed({1'h0, add_519109}) < $signed({1'h0, sel_519111}) ? add_519109 : sel_519111;
  assign add_519663 = array_index_513241[11:0] + 12'h81f;
  assign sel_519665 = $signed({1'h0, add_519113}) < $signed({1'h0, sel_519115}) ? add_519113 : sel_519115;
  assign add_519675 = array_index_513530[11:0] + 12'h45b;
  assign sel_519677 = $signed({1'h0, add_519125}) < $signed({1'h0, sel_519127}) ? add_519125 : sel_519127;
  assign add_519679 = array_index_513533[11:0] + 12'h45b;
  assign sel_519681 = $signed({1'h0, add_519129}) < $signed({1'h0, sel_519131}) ? add_519129 : sel_519131;
  assign add_519693 = array_index_513890[11:3] + 9'h0f5;
  assign sel_519695 = $signed({1'h0, add_519143, array_index_513702[2:0]}) < $signed({1'h0, sel_519145}) ? {add_519143, array_index_513702[2:0]} : sel_519145;
  assign add_519697 = array_index_513893[11:3] + 9'h0f5;
  assign sel_519699 = $signed({1'h0, add_519147, array_index_513705[2:0]}) < $signed({1'h0, sel_519149}) ? {add_519147, array_index_513705[2:0]} : sel_519149;
  assign array_index_519786 = set1_unflattened[5'h1a];
  assign array_index_519789 = set2_unflattened[5'h1a];
  assign add_519799 = array_index_512834[11:0] + 12'h091;
  assign sel_519801 = $signed({1'h0, add_519243}) < $signed(13'h0fff) ? add_519243 : 12'hfff;
  assign add_519803 = array_index_512837[11:0] + 12'h091;
  assign sel_519805 = $signed({1'h0, add_519245}) < $signed(13'h0fff) ? add_519245 : 12'hfff;
  assign add_519815 = array_index_512942[11:0] + 12'hf59;
  assign sel_519817 = $signed({1'h0, add_519257}) < $signed({1'h0, sel_519259}) ? add_519257 : sel_519259;
  assign add_519819 = array_index_512945[11:0] + 12'hf59;
  assign sel_519821 = $signed({1'h0, add_519261}) < $signed({1'h0, sel_519263}) ? add_519261 : sel_519263;
  assign add_519833 = array_index_513120[11:0] + 12'h437;
  assign sel_519835 = $signed({1'h0, add_519275}) < $signed({1'h0, sel_519277}) ? add_519275 : sel_519277;
  assign add_519837 = array_index_513123[11:0] + 12'h437;
  assign sel_519839 = $signed({1'h0, add_519279}) < $signed({1'h0, sel_519281}) ? add_519279 : sel_519281;
  assign add_519849 = array_index_513374[11:0] + 12'hee1;
  assign sel_519851 = $signed({1'h0, add_519291}) < $signed({1'h0, sel_519293}) ? add_519291 : sel_519293;
  assign add_519853 = array_index_513377[11:0] + 12'hee1;
  assign sel_519855 = $signed({1'h0, add_519295}) < $signed({1'h0, sel_519297}) ? add_519295 : sel_519297;
  assign add_519865 = array_index_513702[11:1] + 11'h179;
  assign sel_519867 = $signed({1'h0, add_519307, array_index_513530[0]}) < $signed({1'h0, sel_519309}) ? {add_519307, array_index_513530[0]} : sel_519309;
  assign add_519869 = array_index_513705[11:1] + 11'h179;
  assign sel_519871 = $signed({1'h0, add_519311, array_index_513533[0]}) < $signed({1'h0, sel_519313}) ? {add_519311, array_index_513533[0]} : sel_519313;
  assign add_519881 = array_index_514096[11:0] + 12'h067;
  assign sel_519883 = $signed({1'h0, add_519323}) < $signed({1'h0, sel_519325}) ? add_519323 : sel_519325;
  assign add_519885 = array_index_514099[11:0] + 12'h067;
  assign sel_519887 = $signed({1'h0, add_519327}) < $signed({1'h0, sel_519329}) ? add_519327 : sel_519329;
  assign add_519889 = array_index_514318[11:3] + 9'h1ef;
  assign sel_519892 = $signed({1'h0, add_519331, array_index_514096[2:0]}) < $signed({1'h0, sel_519334}) ? {add_519331, array_index_514096[2:0]} : sel_519334;
  assign add_519894 = array_index_514321[11:3] + 9'h1ef;
  assign sel_519897 = $signed({1'h0, add_519336, array_index_514099[2:0]}) < $signed({1'h0, sel_519339}) ? {add_519336, array_index_514099[2:0]} : sel_519339;
  assign add_519899 = array_index_514558[11:1] + 11'h2d5;
  assign sel_519901 = $signed({1'h0, add_519341, array_index_514318[0]}) < $signed({1'h0, sel_519343}) ? {add_519341, array_index_514318[0]} : sel_519343;
  assign add_519903 = array_index_514561[11:1] + 11'h2d5;
  assign sel_519905 = $signed({1'h0, add_519345, array_index_514321[0]}) < $signed({1'h0, sel_519347}) ? {add_519345, array_index_514321[0]} : sel_519347;
  assign add_519907 = array_index_514818[11:2] + 10'h353;
  assign sel_519909 = $signed({1'h0, add_519349, array_index_514558[1:0]}) < $signed({1'h0, sel_519351}) ? {add_519349, array_index_514558[1:0]} : sel_519351;
  assign add_519911 = array_index_514821[11:2] + 10'h353;
  assign sel_519913 = $signed({1'h0, add_519353, array_index_514561[1:0]}) < $signed({1'h0, sel_519355}) ? {add_519353, array_index_514561[1:0]} : sel_519355;
  assign add_519915 = array_index_515098[11:0] + 12'h0a7;
  assign sel_519917 = $signed({1'h0, add_519357}) < $signed({1'h0, sel_519359}) ? add_519357 : sel_519359;
  assign add_519919 = array_index_515101[11:0] + 12'h0a7;
  assign sel_519921 = $signed({1'h0, add_519361}) < $signed({1'h0, sel_519363}) ? add_519361 : sel_519363;
  assign add_519923 = array_index_515398[11:1] + 11'h4cb;
  assign sel_519925 = $signed({1'h0, add_519365, array_index_515098[0]}) < $signed({1'h0, sel_519367}) ? {add_519365, array_index_515098[0]} : sel_519367;
  assign add_519927 = array_index_515401[11:1] + 11'h4cb;
  assign sel_519929 = $signed({1'h0, add_519369, array_index_515101[0]}) < $signed({1'h0, sel_519371}) ? {add_519369, array_index_515101[0]} : sel_519371;
  assign add_519931 = array_index_515726[11:0] + 12'hfe9;
  assign sel_519933 = $signed({1'h0, add_519373}) < $signed({1'h0, sel_519375}) ? add_519373 : sel_519375;
  assign add_519935 = array_index_515729[11:0] + 12'hfe9;
  assign sel_519937 = $signed({1'h0, add_519377}) < $signed({1'h0, sel_519379}) ? add_519377 : sel_519379;
  assign add_519939 = array_index_516080[11:0] + 12'h97d;
  assign sel_519941 = $signed({1'h0, add_519381}) < $signed({1'h0, sel_519383}) ? add_519381 : sel_519383;
  assign add_519943 = array_index_516083[11:0] + 12'h97d;
  assign sel_519945 = $signed({1'h0, add_519385}) < $signed({1'h0, sel_519387}) ? add_519385 : sel_519387;
  assign add_519947 = array_index_516458[11:2] + 10'h2bb;
  assign sel_519950 = $signed({1'h0, add_519389, array_index_516080[1:0]}) < $signed({1'h0, sel_519392}) ? {add_519389, array_index_516080[1:0]} : sel_519392;
  assign add_519952 = array_index_516461[11:2] + 10'h2bb;
  assign sel_519955 = $signed({1'h0, add_519394, array_index_516083[1:0]}) < $signed({1'h0, sel_519397}) ? {add_519394, array_index_516083[1:0]} : sel_519397;
  assign add_519957 = array_index_516860[11:0] + 12'h8e1;
  assign sel_519959 = $signed({1'h0, add_519399}) < $signed({1'h0, sel_519401}) ? add_519399 : sel_519401;
  assign add_519961 = array_index_516863[11:0] + 12'h8e1;
  assign sel_519963 = $signed({1'h0, add_519403}) < $signed({1'h0, sel_519405}) ? add_519403 : sel_519405;
  assign add_519965 = array_index_517286[11:4] + 8'h83;
  assign sel_519968 = $signed({1'h0, add_519407, array_index_516860[3:0]}) < $signed({1'h0, sel_519410}) ? {add_519407, array_index_516860[3:0]} : sel_519410;
  assign add_519970 = array_index_517289[11:4] + 8'h83;
  assign sel_519973 = $signed({1'h0, add_519412, array_index_516863[3:0]}) < $signed({1'h0, sel_519415}) ? {add_519412, array_index_516863[3:0]} : sel_519415;
  assign add_519975 = array_index_517736[11:0] + 12'ha09;
  assign sel_519977 = $signed({1'h0, add_519417}) < $signed({1'h0, sel_519419}) ? add_519417 : sel_519419;
  assign add_519979 = array_index_517739[11:0] + 12'ha09;
  assign sel_519981 = $signed({1'h0, add_519421}) < $signed({1'h0, sel_519423}) ? add_519421 : sel_519423;
  assign add_519983 = array_index_518210[11:1] + 11'h6cb;
  assign sel_519985 = $signed({1'h0, add_519425, array_index_517736[0]}) < $signed({1'h0, sel_519427}) ? {add_519425, array_index_517736[0]} : sel_519427;
  assign add_519987 = array_index_518213[11:1] + 11'h6cb;
  assign sel_519989 = $signed({1'h0, add_519429, array_index_517739[0]}) < $signed({1'h0, sel_519431}) ? {add_519429, array_index_517739[0]} : sel_519431;
  assign add_519991 = array_index_518710[11:1] + 11'h75d;
  assign sel_519993 = $signed({1'h0, add_519433, array_index_518210[0]}) < $signed({1'h0, sel_519435}) ? {add_519433, array_index_518210[0]} : sel_519435;
  assign add_519995 = array_index_518713[11:1] + 11'h75d;
  assign sel_519997 = $signed({1'h0, add_519437, array_index_518213[0]}) < $signed({1'h0, sel_519439}) ? {add_519437, array_index_518213[0]} : sel_519439;
  assign add_519999 = array_index_519236[11:1] + 11'h24f;
  assign sel_520002 = $signed({1'h0, add_519441, array_index_518710[0]}) < $signed({1'h0, sel_519444}) ? {add_519441, array_index_518710[0]} : sel_519444;
  assign add_520004 = array_index_519239[11:1] + 11'h24f;
  assign sel_520007 = $signed({1'h0, add_519446, array_index_518713[0]}) < $signed({1'h0, sel_519449}) ? {add_519446, array_index_518713[0]} : sel_519449;
  assign add_520015 = array_index_512818[11:0] + 12'h081;
  assign add_520017 = array_index_512819[11:0] + 12'h081;
  assign add_520031 = array_index_512880[11:0] + 12'h0b1;
  assign sel_520033 = $signed({1'h0, add_519463}) < $signed({1'h0, sel_519465}) ? add_519463 : sel_519465;
  assign add_520035 = array_index_512883[11:0] + 12'h0b1;
  assign sel_520037 = $signed({1'h0, add_519467}) < $signed({1'h0, sel_519469}) ? add_519467 : sel_519469;
  assign add_520049 = array_index_513022[11:1] + 11'h4c1;
  assign sel_520051 = $signed({1'h0, add_519481, array_index_512942[0]}) < $signed({1'h0, sel_519483}) ? {add_519481, array_index_512942[0]} : sel_519483;
  assign add_520053 = array_index_513025[11:1] + 11'h4c1;
  assign sel_520055 = $signed({1'h0, add_519485, array_index_512945[0]}) < $signed({1'h0, sel_519487}) ? {add_519485, array_index_512945[0]} : sel_519487;
  assign add_520065 = array_index_513238[11:0] + 12'hbb1;
  assign sel_520067 = $signed({1'h0, add_519497}) < $signed({1'h0, sel_519499}) ? add_519497 : sel_519499;
  assign add_520069 = array_index_513241[11:0] + 12'hbb1;
  assign sel_520071 = $signed({1'h0, add_519501}) < $signed({1'h0, sel_519503}) ? add_519501 : sel_519503;
  assign add_520081 = array_index_513530[11:0] + 12'h6ab;
  assign sel_520083 = $signed({1'h0, add_519513}) < $signed({1'h0, sel_519515}) ? add_519513 : sel_519515;
  assign add_520085 = array_index_513533[11:0] + 12'h6ab;
  assign sel_520087 = $signed({1'h0, add_519517}) < $signed({1'h0, sel_519519}) ? add_519517 : sel_519519;
  assign add_520097 = array_index_513890[11:0] + 12'h7d5;
  assign sel_520099 = $signed({1'h0, add_519529}) < $signed({1'h0, sel_519531}) ? add_519529 : sel_519531;
  assign add_520101 = array_index_513893[11:0] + 12'h7d5;
  assign sel_520103 = $signed({1'h0, add_519533}) < $signed({1'h0, sel_519535}) ? add_519533 : sel_519535;
  assign add_520172 = array_index_519786[11:0] + 12'h62b;
  assign sel_520174 = $signed({1'h0, add_519604}) < $signed({1'h0, sel_519606}) ? add_519604 : sel_519606;
  assign add_520177 = array_index_519789[11:0] + 12'h62b;
  assign sel_520179 = $signed({1'h0, add_519609}) < $signed({1'h0, sel_519611}) ? add_519609 : sel_519611;
  assign add_520187 = array_index_512834[11:1] + 11'h283;
  assign sel_520189 = $signed({1'h0, add_519613, array_index_512818[0]}) < $signed(13'h0fff) ? {add_519613, array_index_512818[0]} : 12'hfff;
  assign add_520191 = array_index_512837[11:1] + 11'h283;
  assign sel_520193 = $signed({1'h0, add_519615, array_index_512819[0]}) < $signed(13'h0fff) ? {add_519615, array_index_512819[0]} : 12'hfff;
  assign add_520203 = array_index_512942[11:1] + 11'h44d;
  assign sel_520205 = $signed({1'h0, add_519627, array_index_512880[0]}) < $signed({1'h0, sel_519629}) ? {add_519627, array_index_512880[0]} : sel_519629;
  assign add_520207 = array_index_512945[11:1] + 11'h44d;
  assign sel_520209 = $signed({1'h0, add_519631, array_index_512883[0]}) < $signed({1'h0, sel_519633}) ? {add_519631, array_index_512883[0]} : sel_519633;
  assign add_520219 = array_index_513120[11:0] + 12'hcb1;
  assign sel_520221 = $signed({1'h0, add_519643}) < $signed({1'h0, sel_519645}) ? add_519643 : sel_519645;
  assign add_520223 = array_index_513123[11:0] + 12'hcb1;
  assign sel_520225 = $signed({1'h0, add_519647}) < $signed({1'h0, sel_519649}) ? add_519647 : sel_519649;
  assign add_520235 = array_index_513374[11:0] + 12'h81f;
  assign sel_520237 = $signed({1'h0, add_519659}) < $signed({1'h0, sel_519661}) ? add_519659 : sel_519661;
  assign add_520239 = array_index_513377[11:0] + 12'h81f;
  assign sel_520241 = $signed({1'h0, add_519663}) < $signed({1'h0, sel_519665}) ? add_519663 : sel_519665;
  assign add_520251 = array_index_513702[11:0] + 12'h45b;
  assign sel_520253 = $signed({1'h0, add_519675}) < $signed({1'h0, sel_519677}) ? add_519675 : sel_519677;
  assign add_520255 = array_index_513705[11:0] + 12'h45b;
  assign sel_520257 = $signed({1'h0, add_519679}) < $signed({1'h0, sel_519681}) ? add_519679 : sel_519681;
  assign add_520269 = array_index_514096[11:3] + 9'h0f5;
  assign sel_520271 = $signed({1'h0, add_519693, array_index_513890[2:0]}) < $signed({1'h0, sel_519695}) ? {add_519693, array_index_513890[2:0]} : sel_519695;
  assign add_520273 = array_index_514099[11:3] + 9'h0f5;
  assign sel_520275 = $signed({1'h0, add_519697, array_index_513893[2:0]}) < $signed({1'h0, sel_519699}) ? {add_519697, array_index_513893[2:0]} : sel_519699;
  assign array_index_520362 = set1_unflattened[5'h1b];
  assign array_index_520365 = set2_unflattened[5'h1b];
  assign add_520369 = array_index_512818[11:3] + 9'h171;
  assign add_520371 = array_index_512819[11:3] + 9'h171;
  assign add_520383 = array_index_512880[11:0] + 12'h091;
  assign sel_520385 = $signed({1'h0, add_519799}) < $signed({1'h0, sel_519801}) ? add_519799 : sel_519801;
  assign add_520387 = array_index_512883[11:0] + 12'h091;
  assign sel_520389 = $signed({1'h0, add_519803}) < $signed({1'h0, sel_519805}) ? add_519803 : sel_519805;
  assign add_520399 = array_index_513022[11:0] + 12'hf59;
  assign sel_520401 = $signed({1'h0, add_519815}) < $signed({1'h0, sel_519817}) ? add_519815 : sel_519817;
  assign add_520403 = array_index_513025[11:0] + 12'hf59;
  assign sel_520405 = $signed({1'h0, add_519819}) < $signed({1'h0, sel_519821}) ? add_519819 : sel_519821;
  assign add_520417 = array_index_513238[11:0] + 12'h437;
  assign sel_520419 = $signed({1'h0, add_519833}) < $signed({1'h0, sel_519835}) ? add_519833 : sel_519835;
  assign add_520421 = array_index_513241[11:0] + 12'h437;
  assign sel_520423 = $signed({1'h0, add_519837}) < $signed({1'h0, sel_519839}) ? add_519837 : sel_519839;
  assign add_520433 = array_index_513530[11:0] + 12'hee1;
  assign sel_520435 = $signed({1'h0, add_519849}) < $signed({1'h0, sel_519851}) ? add_519849 : sel_519851;
  assign add_520437 = array_index_513533[11:0] + 12'hee1;
  assign sel_520439 = $signed({1'h0, add_519853}) < $signed({1'h0, sel_519855}) ? add_519853 : sel_519855;
  assign add_520449 = array_index_513890[11:1] + 11'h179;
  assign sel_520451 = $signed({1'h0, add_519865, array_index_513702[0]}) < $signed({1'h0, sel_519867}) ? {add_519865, array_index_513702[0]} : sel_519867;
  assign add_520453 = array_index_513893[11:1] + 11'h179;
  assign sel_520455 = $signed({1'h0, add_519869, array_index_513705[0]}) < $signed({1'h0, sel_519871}) ? {add_519869, array_index_513705[0]} : sel_519871;
  assign add_520465 = array_index_514318[11:0] + 12'h067;
  assign sel_520467 = $signed({1'h0, add_519881}) < $signed({1'h0, sel_519883}) ? add_519881 : sel_519883;
  assign add_520469 = array_index_514321[11:0] + 12'h067;
  assign sel_520471 = $signed({1'h0, add_519885}) < $signed({1'h0, sel_519887}) ? add_519885 : sel_519887;
  assign add_520473 = array_index_514558[11:3] + 9'h1ef;
  assign sel_520476 = $signed({1'h0, add_519889, array_index_514318[2:0]}) < $signed({1'h0, sel_519892}) ? {add_519889, array_index_514318[2:0]} : sel_519892;
  assign add_520478 = array_index_514561[11:3] + 9'h1ef;
  assign sel_520481 = $signed({1'h0, add_519894, array_index_514321[2:0]}) < $signed({1'h0, sel_519897}) ? {add_519894, array_index_514321[2:0]} : sel_519897;
  assign add_520483 = array_index_514818[11:1] + 11'h2d5;
  assign sel_520485 = $signed({1'h0, add_519899, array_index_514558[0]}) < $signed({1'h0, sel_519901}) ? {add_519899, array_index_514558[0]} : sel_519901;
  assign add_520487 = array_index_514821[11:1] + 11'h2d5;
  assign sel_520489 = $signed({1'h0, add_519903, array_index_514561[0]}) < $signed({1'h0, sel_519905}) ? {add_519903, array_index_514561[0]} : sel_519905;
  assign add_520491 = array_index_515098[11:2] + 10'h353;
  assign sel_520493 = $signed({1'h0, add_519907, array_index_514818[1:0]}) < $signed({1'h0, sel_519909}) ? {add_519907, array_index_514818[1:0]} : sel_519909;
  assign add_520495 = array_index_515101[11:2] + 10'h353;
  assign sel_520497 = $signed({1'h0, add_519911, array_index_514821[1:0]}) < $signed({1'h0, sel_519913}) ? {add_519911, array_index_514821[1:0]} : sel_519913;
  assign add_520499 = array_index_515398[11:0] + 12'h0a7;
  assign sel_520501 = $signed({1'h0, add_519915}) < $signed({1'h0, sel_519917}) ? add_519915 : sel_519917;
  assign add_520503 = array_index_515401[11:0] + 12'h0a7;
  assign sel_520505 = $signed({1'h0, add_519919}) < $signed({1'h0, sel_519921}) ? add_519919 : sel_519921;
  assign add_520507 = array_index_515726[11:1] + 11'h4cb;
  assign sel_520509 = $signed({1'h0, add_519923, array_index_515398[0]}) < $signed({1'h0, sel_519925}) ? {add_519923, array_index_515398[0]} : sel_519925;
  assign add_520511 = array_index_515729[11:1] + 11'h4cb;
  assign sel_520513 = $signed({1'h0, add_519927, array_index_515401[0]}) < $signed({1'h0, sel_519929}) ? {add_519927, array_index_515401[0]} : sel_519929;
  assign add_520515 = array_index_516080[11:0] + 12'hfe9;
  assign sel_520517 = $signed({1'h0, add_519931}) < $signed({1'h0, sel_519933}) ? add_519931 : sel_519933;
  assign add_520519 = array_index_516083[11:0] + 12'hfe9;
  assign sel_520521 = $signed({1'h0, add_519935}) < $signed({1'h0, sel_519937}) ? add_519935 : sel_519937;
  assign add_520523 = array_index_516458[11:0] + 12'h97d;
  assign sel_520525 = $signed({1'h0, add_519939}) < $signed({1'h0, sel_519941}) ? add_519939 : sel_519941;
  assign add_520527 = array_index_516461[11:0] + 12'h97d;
  assign sel_520529 = $signed({1'h0, add_519943}) < $signed({1'h0, sel_519945}) ? add_519943 : sel_519945;
  assign add_520531 = array_index_516860[11:2] + 10'h2bb;
  assign sel_520534 = $signed({1'h0, add_519947, array_index_516458[1:0]}) < $signed({1'h0, sel_519950}) ? {add_519947, array_index_516458[1:0]} : sel_519950;
  assign add_520536 = array_index_516863[11:2] + 10'h2bb;
  assign sel_520539 = $signed({1'h0, add_519952, array_index_516461[1:0]}) < $signed({1'h0, sel_519955}) ? {add_519952, array_index_516461[1:0]} : sel_519955;
  assign add_520541 = array_index_517286[11:0] + 12'h8e1;
  assign sel_520543 = $signed({1'h0, add_519957}) < $signed({1'h0, sel_519959}) ? add_519957 : sel_519959;
  assign add_520545 = array_index_517289[11:0] + 12'h8e1;
  assign sel_520547 = $signed({1'h0, add_519961}) < $signed({1'h0, sel_519963}) ? add_519961 : sel_519963;
  assign add_520549 = array_index_517736[11:4] + 8'h83;
  assign sel_520552 = $signed({1'h0, add_519965, array_index_517286[3:0]}) < $signed({1'h0, sel_519968}) ? {add_519965, array_index_517286[3:0]} : sel_519968;
  assign add_520554 = array_index_517739[11:4] + 8'h83;
  assign sel_520557 = $signed({1'h0, add_519970, array_index_517289[3:0]}) < $signed({1'h0, sel_519973}) ? {add_519970, array_index_517289[3:0]} : sel_519973;
  assign add_520559 = array_index_518210[11:0] + 12'ha09;
  assign sel_520561 = $signed({1'h0, add_519975}) < $signed({1'h0, sel_519977}) ? add_519975 : sel_519977;
  assign add_520563 = array_index_518213[11:0] + 12'ha09;
  assign sel_520565 = $signed({1'h0, add_519979}) < $signed({1'h0, sel_519981}) ? add_519979 : sel_519981;
  assign add_520567 = array_index_518710[11:1] + 11'h6cb;
  assign sel_520569 = $signed({1'h0, add_519983, array_index_518210[0]}) < $signed({1'h0, sel_519985}) ? {add_519983, array_index_518210[0]} : sel_519985;
  assign add_520571 = array_index_518713[11:1] + 11'h6cb;
  assign sel_520573 = $signed({1'h0, add_519987, array_index_518213[0]}) < $signed({1'h0, sel_519989}) ? {add_519987, array_index_518213[0]} : sel_519989;
  assign add_520575 = array_index_519236[11:1] + 11'h75d;
  assign sel_520577 = $signed({1'h0, add_519991, array_index_518710[0]}) < $signed({1'h0, sel_519993}) ? {add_519991, array_index_518710[0]} : sel_519993;
  assign add_520579 = array_index_519239[11:1] + 11'h75d;
  assign sel_520581 = $signed({1'h0, add_519995, array_index_518713[0]}) < $signed({1'h0, sel_519997}) ? {add_519995, array_index_518713[0]} : sel_519997;
  assign add_520583 = array_index_519786[11:1] + 11'h24f;
  assign sel_520586 = $signed({1'h0, add_519999, array_index_519236[0]}) < $signed({1'h0, sel_520002}) ? {add_519999, array_index_519236[0]} : sel_520002;
  assign add_520588 = array_index_519789[11:1] + 11'h24f;
  assign sel_520591 = $signed({1'h0, add_520004, array_index_519239[0]}) < $signed({1'h0, sel_520007}) ? {add_520004, array_index_519239[0]} : sel_520007;
  assign add_520605 = array_index_512834[11:0] + 12'h081;
  assign sel_520607 = $signed({1'h0, add_520015}) < $signed(13'h0fff) ? add_520015 : 12'hfff;
  assign add_520609 = array_index_512837[11:0] + 12'h081;
  assign sel_520611 = $signed({1'h0, add_520017}) < $signed(13'h0fff) ? add_520017 : 12'hfff;
  assign add_520623 = array_index_512942[11:0] + 12'h0b1;
  assign sel_520625 = $signed({1'h0, add_520031}) < $signed({1'h0, sel_520033}) ? add_520031 : sel_520033;
  assign add_520627 = array_index_512945[11:0] + 12'h0b1;
  assign sel_520629 = $signed({1'h0, add_520035}) < $signed({1'h0, sel_520037}) ? add_520035 : sel_520037;
  assign add_520641 = array_index_513120[11:1] + 11'h4c1;
  assign sel_520643 = $signed({1'h0, add_520049, array_index_513022[0]}) < $signed({1'h0, sel_520051}) ? {add_520049, array_index_513022[0]} : sel_520051;
  assign add_520645 = array_index_513123[11:1] + 11'h4c1;
  assign sel_520647 = $signed({1'h0, add_520053, array_index_513025[0]}) < $signed({1'h0, sel_520055}) ? {add_520053, array_index_513025[0]} : sel_520055;
  assign add_520657 = array_index_513374[11:0] + 12'hbb1;
  assign sel_520659 = $signed({1'h0, add_520065}) < $signed({1'h0, sel_520067}) ? add_520065 : sel_520067;
  assign add_520661 = array_index_513377[11:0] + 12'hbb1;
  assign sel_520663 = $signed({1'h0, add_520069}) < $signed({1'h0, sel_520071}) ? add_520069 : sel_520071;
  assign add_520673 = array_index_513702[11:0] + 12'h6ab;
  assign sel_520675 = $signed({1'h0, add_520081}) < $signed({1'h0, sel_520083}) ? add_520081 : sel_520083;
  assign add_520677 = array_index_513705[11:0] + 12'h6ab;
  assign sel_520679 = $signed({1'h0, add_520085}) < $signed({1'h0, sel_520087}) ? add_520085 : sel_520087;
  assign add_520689 = array_index_514096[11:0] + 12'h7d5;
  assign sel_520691 = $signed({1'h0, add_520097}) < $signed({1'h0, sel_520099}) ? add_520097 : sel_520099;
  assign add_520693 = array_index_514099[11:0] + 12'h7d5;
  assign sel_520695 = $signed({1'h0, add_520101}) < $signed({1'h0, sel_520103}) ? add_520101 : sel_520103;
  assign add_520764 = array_index_520362[11:0] + 12'h62b;
  assign sel_520766 = $signed({1'h0, add_520172}) < $signed({1'h0, sel_520174}) ? add_520172 : sel_520174;
  assign add_520769 = array_index_520365[11:0] + 12'h62b;
  assign sel_520771 = $signed({1'h0, add_520177}) < $signed({1'h0, sel_520179}) ? add_520177 : sel_520179;
  assign add_520773 = array_index_512818[11:0] + 12'h8a7;
  assign add_520775 = array_index_512819[11:0] + 12'h8a7;
  assign add_520789 = array_index_512880[11:1] + 11'h283;
  assign sel_520791 = $signed({1'h0, add_520187, array_index_512834[0]}) < $signed({1'h0, sel_520189}) ? {add_520187, array_index_512834[0]} : sel_520189;
  assign add_520793 = array_index_512883[11:1] + 11'h283;
  assign sel_520795 = $signed({1'h0, add_520191, array_index_512837[0]}) < $signed({1'h0, sel_520193}) ? {add_520191, array_index_512837[0]} : sel_520193;
  assign add_520805 = array_index_513022[11:1] + 11'h44d;
  assign sel_520807 = $signed({1'h0, add_520203, array_index_512942[0]}) < $signed({1'h0, sel_520205}) ? {add_520203, array_index_512942[0]} : sel_520205;
  assign add_520809 = array_index_513025[11:1] + 11'h44d;
  assign sel_520811 = $signed({1'h0, add_520207, array_index_512945[0]}) < $signed({1'h0, sel_520209}) ? {add_520207, array_index_512945[0]} : sel_520209;
  assign add_520821 = array_index_513238[11:0] + 12'hcb1;
  assign sel_520823 = $signed({1'h0, add_520219}) < $signed({1'h0, sel_520221}) ? add_520219 : sel_520221;
  assign add_520825 = array_index_513241[11:0] + 12'hcb1;
  assign sel_520827 = $signed({1'h0, add_520223}) < $signed({1'h0, sel_520225}) ? add_520223 : sel_520225;
  assign add_520837 = array_index_513530[11:0] + 12'h81f;
  assign sel_520839 = $signed({1'h0, add_520235}) < $signed({1'h0, sel_520237}) ? add_520235 : sel_520237;
  assign add_520841 = array_index_513533[11:0] + 12'h81f;
  assign sel_520843 = $signed({1'h0, add_520239}) < $signed({1'h0, sel_520241}) ? add_520239 : sel_520241;
  assign add_520853 = array_index_513890[11:0] + 12'h45b;
  assign sel_520855 = $signed({1'h0, add_520251}) < $signed({1'h0, sel_520253}) ? add_520251 : sel_520253;
  assign add_520857 = array_index_513893[11:0] + 12'h45b;
  assign sel_520859 = $signed({1'h0, add_520255}) < $signed({1'h0, sel_520257}) ? add_520255 : sel_520257;
  assign add_520871 = array_index_514318[11:3] + 9'h0f5;
  assign sel_520873 = $signed({1'h0, add_520269, array_index_514096[2:0]}) < $signed({1'h0, sel_520271}) ? {add_520269, array_index_514096[2:0]} : sel_520271;
  assign add_520875 = array_index_514321[11:3] + 9'h0f5;
  assign sel_520877 = $signed({1'h0, add_520273, array_index_514099[2:0]}) < $signed({1'h0, sel_520275}) ? {add_520273, array_index_514099[2:0]} : sel_520275;
  assign array_index_520964 = set1_unflattened[5'h1c];
  assign array_index_520967 = set2_unflattened[5'h1c];
  assign add_520977 = array_index_512834[11:3] + 9'h171;
  assign sel_520979 = $signed({1'h0, add_520369, array_index_512818[2:0]}) < $signed(13'h0fff) ? {add_520369, array_index_512818[2:0]} : 12'hfff;
  assign add_520981 = array_index_512837[11:3] + 9'h171;
  assign sel_520983 = $signed({1'h0, add_520371, array_index_512819[2:0]}) < $signed(13'h0fff) ? {add_520371, array_index_512819[2:0]} : 12'hfff;
  assign add_520993 = array_index_512942[11:0] + 12'h091;
  assign sel_520995 = $signed({1'h0, add_520383}) < $signed({1'h0, sel_520385}) ? add_520383 : sel_520385;
  assign add_520997 = array_index_512945[11:0] + 12'h091;
  assign sel_520999 = $signed({1'h0, add_520387}) < $signed({1'h0, sel_520389}) ? add_520387 : sel_520389;
  assign add_521009 = array_index_513120[11:0] + 12'hf59;
  assign sel_521011 = $signed({1'h0, add_520399}) < $signed({1'h0, sel_520401}) ? add_520399 : sel_520401;
  assign add_521013 = array_index_513123[11:0] + 12'hf59;
  assign sel_521015 = $signed({1'h0, add_520403}) < $signed({1'h0, sel_520405}) ? add_520403 : sel_520405;
  assign add_521027 = array_index_513374[11:0] + 12'h437;
  assign sel_521029 = $signed({1'h0, add_520417}) < $signed({1'h0, sel_520419}) ? add_520417 : sel_520419;
  assign add_521031 = array_index_513377[11:0] + 12'h437;
  assign sel_521033 = $signed({1'h0, add_520421}) < $signed({1'h0, sel_520423}) ? add_520421 : sel_520423;
  assign add_521043 = array_index_513702[11:0] + 12'hee1;
  assign sel_521045 = $signed({1'h0, add_520433}) < $signed({1'h0, sel_520435}) ? add_520433 : sel_520435;
  assign add_521047 = array_index_513705[11:0] + 12'hee1;
  assign sel_521049 = $signed({1'h0, add_520437}) < $signed({1'h0, sel_520439}) ? add_520437 : sel_520439;
  assign add_521059 = array_index_514096[11:1] + 11'h179;
  assign sel_521061 = $signed({1'h0, add_520449, array_index_513890[0]}) < $signed({1'h0, sel_520451}) ? {add_520449, array_index_513890[0]} : sel_520451;
  assign add_521063 = array_index_514099[11:1] + 11'h179;
  assign sel_521065 = $signed({1'h0, add_520453, array_index_513893[0]}) < $signed({1'h0, sel_520455}) ? {add_520453, array_index_513893[0]} : sel_520455;
  assign add_521075 = array_index_514558[11:0] + 12'h067;
  assign sel_521077 = $signed({1'h0, add_520465}) < $signed({1'h0, sel_520467}) ? add_520465 : sel_520467;
  assign add_521079 = array_index_514561[11:0] + 12'h067;
  assign sel_521081 = $signed({1'h0, add_520469}) < $signed({1'h0, sel_520471}) ? add_520469 : sel_520471;
  assign add_521083 = array_index_514818[11:3] + 9'h1ef;
  assign sel_521086 = $signed({1'h0, add_520473, array_index_514558[2:0]}) < $signed({1'h0, sel_520476}) ? {add_520473, array_index_514558[2:0]} : sel_520476;
  assign add_521088 = array_index_514821[11:3] + 9'h1ef;
  assign sel_521091 = $signed({1'h0, add_520478, array_index_514561[2:0]}) < $signed({1'h0, sel_520481}) ? {add_520478, array_index_514561[2:0]} : sel_520481;
  assign add_521093 = array_index_515098[11:1] + 11'h2d5;
  assign sel_521095 = $signed({1'h0, add_520483, array_index_514818[0]}) < $signed({1'h0, sel_520485}) ? {add_520483, array_index_514818[0]} : sel_520485;
  assign add_521097 = array_index_515101[11:1] + 11'h2d5;
  assign sel_521099 = $signed({1'h0, add_520487, array_index_514821[0]}) < $signed({1'h0, sel_520489}) ? {add_520487, array_index_514821[0]} : sel_520489;
  assign add_521101 = array_index_515398[11:2] + 10'h353;
  assign sel_521103 = $signed({1'h0, add_520491, array_index_515098[1:0]}) < $signed({1'h0, sel_520493}) ? {add_520491, array_index_515098[1:0]} : sel_520493;
  assign add_521105 = array_index_515401[11:2] + 10'h353;
  assign sel_521107 = $signed({1'h0, add_520495, array_index_515101[1:0]}) < $signed({1'h0, sel_520497}) ? {add_520495, array_index_515101[1:0]} : sel_520497;
  assign add_521109 = array_index_515726[11:0] + 12'h0a7;
  assign sel_521111 = $signed({1'h0, add_520499}) < $signed({1'h0, sel_520501}) ? add_520499 : sel_520501;
  assign add_521113 = array_index_515729[11:0] + 12'h0a7;
  assign sel_521115 = $signed({1'h0, add_520503}) < $signed({1'h0, sel_520505}) ? add_520503 : sel_520505;
  assign add_521117 = array_index_516080[11:1] + 11'h4cb;
  assign sel_521119 = $signed({1'h0, add_520507, array_index_515726[0]}) < $signed({1'h0, sel_520509}) ? {add_520507, array_index_515726[0]} : sel_520509;
  assign add_521121 = array_index_516083[11:1] + 11'h4cb;
  assign sel_521123 = $signed({1'h0, add_520511, array_index_515729[0]}) < $signed({1'h0, sel_520513}) ? {add_520511, array_index_515729[0]} : sel_520513;
  assign add_521125 = array_index_516458[11:0] + 12'hfe9;
  assign sel_521127 = $signed({1'h0, add_520515}) < $signed({1'h0, sel_520517}) ? add_520515 : sel_520517;
  assign add_521129 = array_index_516461[11:0] + 12'hfe9;
  assign sel_521131 = $signed({1'h0, add_520519}) < $signed({1'h0, sel_520521}) ? add_520519 : sel_520521;
  assign add_521133 = array_index_516860[11:0] + 12'h97d;
  assign sel_521135 = $signed({1'h0, add_520523}) < $signed({1'h0, sel_520525}) ? add_520523 : sel_520525;
  assign add_521137 = array_index_516863[11:0] + 12'h97d;
  assign sel_521139 = $signed({1'h0, add_520527}) < $signed({1'h0, sel_520529}) ? add_520527 : sel_520529;
  assign add_521141 = array_index_517286[11:2] + 10'h2bb;
  assign sel_521144 = $signed({1'h0, add_520531, array_index_516860[1:0]}) < $signed({1'h0, sel_520534}) ? {add_520531, array_index_516860[1:0]} : sel_520534;
  assign add_521146 = array_index_517289[11:2] + 10'h2bb;
  assign sel_521149 = $signed({1'h0, add_520536, array_index_516863[1:0]}) < $signed({1'h0, sel_520539}) ? {add_520536, array_index_516863[1:0]} : sel_520539;
  assign add_521151 = array_index_517736[11:0] + 12'h8e1;
  assign sel_521153 = $signed({1'h0, add_520541}) < $signed({1'h0, sel_520543}) ? add_520541 : sel_520543;
  assign add_521155 = array_index_517739[11:0] + 12'h8e1;
  assign sel_521157 = $signed({1'h0, add_520545}) < $signed({1'h0, sel_520547}) ? add_520545 : sel_520547;
  assign add_521159 = array_index_518210[11:4] + 8'h83;
  assign sel_521162 = $signed({1'h0, add_520549, array_index_517736[3:0]}) < $signed({1'h0, sel_520552}) ? {add_520549, array_index_517736[3:0]} : sel_520552;
  assign add_521164 = array_index_518213[11:4] + 8'h83;
  assign sel_521167 = $signed({1'h0, add_520554, array_index_517739[3:0]}) < $signed({1'h0, sel_520557}) ? {add_520554, array_index_517739[3:0]} : sel_520557;
  assign add_521169 = array_index_518710[11:0] + 12'ha09;
  assign sel_521171 = $signed({1'h0, add_520559}) < $signed({1'h0, sel_520561}) ? add_520559 : sel_520561;
  assign add_521173 = array_index_518713[11:0] + 12'ha09;
  assign sel_521175 = $signed({1'h0, add_520563}) < $signed({1'h0, sel_520565}) ? add_520563 : sel_520565;
  assign add_521177 = array_index_519236[11:1] + 11'h6cb;
  assign sel_521179 = $signed({1'h0, add_520567, array_index_518710[0]}) < $signed({1'h0, sel_520569}) ? {add_520567, array_index_518710[0]} : sel_520569;
  assign add_521181 = array_index_519239[11:1] + 11'h6cb;
  assign sel_521183 = $signed({1'h0, add_520571, array_index_518713[0]}) < $signed({1'h0, sel_520573}) ? {add_520571, array_index_518713[0]} : sel_520573;
  assign add_521185 = array_index_519786[11:1] + 11'h75d;
  assign sel_521187 = $signed({1'h0, add_520575, array_index_519236[0]}) < $signed({1'h0, sel_520577}) ? {add_520575, array_index_519236[0]} : sel_520577;
  assign add_521189 = array_index_519789[11:1] + 11'h75d;
  assign sel_521191 = $signed({1'h0, add_520579, array_index_519239[0]}) < $signed({1'h0, sel_520581}) ? {add_520579, array_index_519239[0]} : sel_520581;
  assign add_521193 = array_index_520362[11:1] + 11'h24f;
  assign sel_521196 = $signed({1'h0, add_520583, array_index_519786[0]}) < $signed({1'h0, sel_520586}) ? {add_520583, array_index_519786[0]} : sel_520586;
  assign add_521198 = array_index_520365[11:1] + 11'h24f;
  assign sel_521201 = $signed({1'h0, add_520588, array_index_519789[0]}) < $signed({1'h0, sel_520591}) ? {add_520588, array_index_519789[0]} : sel_520591;
  assign add_521209 = array_index_512818[11:3] + 9'h1f1;
  assign add_521211 = array_index_512819[11:3] + 9'h1f1;
  assign add_521223 = array_index_512880[11:0] + 12'h081;
  assign sel_521225 = $signed({1'h0, add_520605}) < $signed({1'h0, sel_520607}) ? add_520605 : sel_520607;
  assign add_521227 = array_index_512883[11:0] + 12'h081;
  assign sel_521229 = $signed({1'h0, add_520609}) < $signed({1'h0, sel_520611}) ? add_520609 : sel_520611;
  assign add_521241 = array_index_513022[11:0] + 12'h0b1;
  assign sel_521243 = $signed({1'h0, add_520623}) < $signed({1'h0, sel_520625}) ? add_520623 : sel_520625;
  assign add_521245 = array_index_513025[11:0] + 12'h0b1;
  assign sel_521247 = $signed({1'h0, add_520627}) < $signed({1'h0, sel_520629}) ? add_520627 : sel_520629;
  assign add_521259 = array_index_513238[11:1] + 11'h4c1;
  assign sel_521261 = $signed({1'h0, add_520641, array_index_513120[0]}) < $signed({1'h0, sel_520643}) ? {add_520641, array_index_513120[0]} : sel_520643;
  assign add_521263 = array_index_513241[11:1] + 11'h4c1;
  assign sel_521265 = $signed({1'h0, add_520645, array_index_513123[0]}) < $signed({1'h0, sel_520647}) ? {add_520645, array_index_513123[0]} : sel_520647;
  assign add_521275 = array_index_513530[11:0] + 12'hbb1;
  assign sel_521277 = $signed({1'h0, add_520657}) < $signed({1'h0, sel_520659}) ? add_520657 : sel_520659;
  assign add_521279 = array_index_513533[11:0] + 12'hbb1;
  assign sel_521281 = $signed({1'h0, add_520661}) < $signed({1'h0, sel_520663}) ? add_520661 : sel_520663;
  assign add_521291 = array_index_513890[11:0] + 12'h6ab;
  assign sel_521293 = $signed({1'h0, add_520673}) < $signed({1'h0, sel_520675}) ? add_520673 : sel_520675;
  assign add_521295 = array_index_513893[11:0] + 12'h6ab;
  assign sel_521297 = $signed({1'h0, add_520677}) < $signed({1'h0, sel_520679}) ? add_520677 : sel_520679;
  assign add_521307 = array_index_514318[11:0] + 12'h7d5;
  assign sel_521309 = $signed({1'h0, add_520689}) < $signed({1'h0, sel_520691}) ? add_520689 : sel_520691;
  assign add_521311 = array_index_514321[11:0] + 12'h7d5;
  assign sel_521313 = $signed({1'h0, add_520693}) < $signed({1'h0, sel_520695}) ? add_520693 : sel_520695;
  assign add_521382 = array_index_520964[11:0] + 12'h62b;
  assign sel_521384 = $signed({1'h0, add_520764}) < $signed({1'h0, sel_520766}) ? add_520764 : sel_520766;
  assign add_521387 = array_index_520967[11:0] + 12'h62b;
  assign sel_521389 = $signed({1'h0, add_520769}) < $signed({1'h0, sel_520771}) ? add_520769 : sel_520771;
  assign add_521397 = array_index_512834[11:0] + 12'h8a7;
  assign sel_521399 = $signed({1'h0, add_520773}) < $signed(13'h0fff) ? add_520773 : 12'hfff;
  assign add_521401 = array_index_512837[11:0] + 12'h8a7;
  assign sel_521403 = $signed({1'h0, add_520775}) < $signed(13'h0fff) ? add_520775 : 12'hfff;
  assign add_521415 = array_index_512942[11:1] + 11'h283;
  assign sel_521417 = $signed({1'h0, add_520789, array_index_512880[0]}) < $signed({1'h0, sel_520791}) ? {add_520789, array_index_512880[0]} : sel_520791;
  assign add_521419 = array_index_512945[11:1] + 11'h283;
  assign sel_521421 = $signed({1'h0, add_520793, array_index_512883[0]}) < $signed({1'h0, sel_520795}) ? {add_520793, array_index_512883[0]} : sel_520795;
  assign add_521431 = array_index_513120[11:1] + 11'h44d;
  assign sel_521433 = $signed({1'h0, add_520805, array_index_513022[0]}) < $signed({1'h0, sel_520807}) ? {add_520805, array_index_513022[0]} : sel_520807;
  assign add_521435 = array_index_513123[11:1] + 11'h44d;
  assign sel_521437 = $signed({1'h0, add_520809, array_index_513025[0]}) < $signed({1'h0, sel_520811}) ? {add_520809, array_index_513025[0]} : sel_520811;
  assign add_521447 = array_index_513374[11:0] + 12'hcb1;
  assign sel_521449 = $signed({1'h0, add_520821}) < $signed({1'h0, sel_520823}) ? add_520821 : sel_520823;
  assign add_521451 = array_index_513377[11:0] + 12'hcb1;
  assign sel_521453 = $signed({1'h0, add_520825}) < $signed({1'h0, sel_520827}) ? add_520825 : sel_520827;
  assign add_521463 = array_index_513702[11:0] + 12'h81f;
  assign sel_521465 = $signed({1'h0, add_520837}) < $signed({1'h0, sel_520839}) ? add_520837 : sel_520839;
  assign add_521467 = array_index_513705[11:0] + 12'h81f;
  assign sel_521469 = $signed({1'h0, add_520841}) < $signed({1'h0, sel_520843}) ? add_520841 : sel_520843;
  assign add_521479 = array_index_514096[11:0] + 12'h45b;
  assign sel_521481 = $signed({1'h0, add_520853}) < $signed({1'h0, sel_520855}) ? add_520853 : sel_520855;
  assign add_521483 = array_index_514099[11:0] + 12'h45b;
  assign sel_521485 = $signed({1'h0, add_520857}) < $signed({1'h0, sel_520859}) ? add_520857 : sel_520859;
  assign add_521497 = array_index_514558[11:3] + 9'h0f5;
  assign sel_521499 = $signed({1'h0, add_520871, array_index_514318[2:0]}) < $signed({1'h0, sel_520873}) ? {add_520871, array_index_514318[2:0]} : sel_520873;
  assign add_521501 = array_index_514561[11:3] + 9'h0f5;
  assign sel_521503 = $signed({1'h0, add_520875, array_index_514321[2:0]}) < $signed({1'h0, sel_520877}) ? {add_520875, array_index_514321[2:0]} : sel_520877;
  assign array_index_521590 = set1_unflattened[5'h1d];
  assign array_index_521593 = set2_unflattened[5'h1d];
  assign add_521597 = array_index_512818[11:3] + 9'h12f;
  assign add_521599 = array_index_512819[11:3] + 9'h12f;
  assign add_521613 = array_index_512880[11:3] + 9'h171;
  assign sel_521615 = $signed({1'h0, add_520977, array_index_512834[2:0]}) < $signed({1'h0, sel_520979}) ? {add_520977, array_index_512834[2:0]} : sel_520979;
  assign add_521617 = array_index_512883[11:3] + 9'h171;
  assign sel_521619 = $signed({1'h0, add_520981, array_index_512837[2:0]}) < $signed({1'h0, sel_520983}) ? {add_520981, array_index_512837[2:0]} : sel_520983;
  assign add_521629 = array_index_513022[11:0] + 12'h091;
  assign sel_521631 = $signed({1'h0, add_520993}) < $signed({1'h0, sel_520995}) ? add_520993 : sel_520995;
  assign add_521633 = array_index_513025[11:0] + 12'h091;
  assign sel_521635 = $signed({1'h0, add_520997}) < $signed({1'h0, sel_520999}) ? add_520997 : sel_520999;
  assign add_521645 = array_index_513238[11:0] + 12'hf59;
  assign sel_521647 = $signed({1'h0, add_521009}) < $signed({1'h0, sel_521011}) ? add_521009 : sel_521011;
  assign add_521649 = array_index_513241[11:0] + 12'hf59;
  assign sel_521651 = $signed({1'h0, add_521013}) < $signed({1'h0, sel_521015}) ? add_521013 : sel_521015;
  assign add_521663 = array_index_513530[11:0] + 12'h437;
  assign sel_521665 = $signed({1'h0, add_521027}) < $signed({1'h0, sel_521029}) ? add_521027 : sel_521029;
  assign add_521667 = array_index_513533[11:0] + 12'h437;
  assign sel_521669 = $signed({1'h0, add_521031}) < $signed({1'h0, sel_521033}) ? add_521031 : sel_521033;
  assign add_521679 = array_index_513890[11:0] + 12'hee1;
  assign sel_521681 = $signed({1'h0, add_521043}) < $signed({1'h0, sel_521045}) ? add_521043 : sel_521045;
  assign add_521683 = array_index_513893[11:0] + 12'hee1;
  assign sel_521685 = $signed({1'h0, add_521047}) < $signed({1'h0, sel_521049}) ? add_521047 : sel_521049;
  assign add_521695 = array_index_514318[11:1] + 11'h179;
  assign sel_521697 = $signed({1'h0, add_521059, array_index_514096[0]}) < $signed({1'h0, sel_521061}) ? {add_521059, array_index_514096[0]} : sel_521061;
  assign add_521699 = array_index_514321[11:1] + 11'h179;
  assign sel_521701 = $signed({1'h0, add_521063, array_index_514099[0]}) < $signed({1'h0, sel_521065}) ? {add_521063, array_index_514099[0]} : sel_521065;
  assign add_521711 = array_index_514818[11:0] + 12'h067;
  assign sel_521713 = $signed({1'h0, add_521075}) < $signed({1'h0, sel_521077}) ? add_521075 : sel_521077;
  assign add_521715 = array_index_514821[11:0] + 12'h067;
  assign sel_521717 = $signed({1'h0, add_521079}) < $signed({1'h0, sel_521081}) ? add_521079 : sel_521081;
  assign add_521719 = array_index_515098[11:3] + 9'h1ef;
  assign sel_521722 = $signed({1'h0, add_521083, array_index_514818[2:0]}) < $signed({1'h0, sel_521086}) ? {add_521083, array_index_514818[2:0]} : sel_521086;
  assign add_521724 = array_index_515101[11:3] + 9'h1ef;
  assign sel_521727 = $signed({1'h0, add_521088, array_index_514821[2:0]}) < $signed({1'h0, sel_521091}) ? {add_521088, array_index_514821[2:0]} : sel_521091;
  assign add_521729 = array_index_515398[11:1] + 11'h2d5;
  assign sel_521731 = $signed({1'h0, add_521093, array_index_515098[0]}) < $signed({1'h0, sel_521095}) ? {add_521093, array_index_515098[0]} : sel_521095;
  assign add_521733 = array_index_515401[11:1] + 11'h2d5;
  assign sel_521735 = $signed({1'h0, add_521097, array_index_515101[0]}) < $signed({1'h0, sel_521099}) ? {add_521097, array_index_515101[0]} : sel_521099;
  assign add_521737 = array_index_515726[11:2] + 10'h353;
  assign sel_521739 = $signed({1'h0, add_521101, array_index_515398[1:0]}) < $signed({1'h0, sel_521103}) ? {add_521101, array_index_515398[1:0]} : sel_521103;
  assign add_521741 = array_index_515729[11:2] + 10'h353;
  assign sel_521743 = $signed({1'h0, add_521105, array_index_515401[1:0]}) < $signed({1'h0, sel_521107}) ? {add_521105, array_index_515401[1:0]} : sel_521107;
  assign add_521745 = array_index_516080[11:0] + 12'h0a7;
  assign sel_521747 = $signed({1'h0, add_521109}) < $signed({1'h0, sel_521111}) ? add_521109 : sel_521111;
  assign add_521749 = array_index_516083[11:0] + 12'h0a7;
  assign sel_521751 = $signed({1'h0, add_521113}) < $signed({1'h0, sel_521115}) ? add_521113 : sel_521115;
  assign add_521753 = array_index_516458[11:1] + 11'h4cb;
  assign sel_521755 = $signed({1'h0, add_521117, array_index_516080[0]}) < $signed({1'h0, sel_521119}) ? {add_521117, array_index_516080[0]} : sel_521119;
  assign add_521757 = array_index_516461[11:1] + 11'h4cb;
  assign sel_521759 = $signed({1'h0, add_521121, array_index_516083[0]}) < $signed({1'h0, sel_521123}) ? {add_521121, array_index_516083[0]} : sel_521123;
  assign add_521761 = array_index_516860[11:0] + 12'hfe9;
  assign sel_521763 = $signed({1'h0, add_521125}) < $signed({1'h0, sel_521127}) ? add_521125 : sel_521127;
  assign add_521765 = array_index_516863[11:0] + 12'hfe9;
  assign sel_521767 = $signed({1'h0, add_521129}) < $signed({1'h0, sel_521131}) ? add_521129 : sel_521131;
  assign add_521769 = array_index_517286[11:0] + 12'h97d;
  assign sel_521771 = $signed({1'h0, add_521133}) < $signed({1'h0, sel_521135}) ? add_521133 : sel_521135;
  assign add_521773 = array_index_517289[11:0] + 12'h97d;
  assign sel_521775 = $signed({1'h0, add_521137}) < $signed({1'h0, sel_521139}) ? add_521137 : sel_521139;
  assign add_521777 = array_index_517736[11:2] + 10'h2bb;
  assign sel_521780 = $signed({1'h0, add_521141, array_index_517286[1:0]}) < $signed({1'h0, sel_521144}) ? {add_521141, array_index_517286[1:0]} : sel_521144;
  assign add_521782 = array_index_517739[11:2] + 10'h2bb;
  assign sel_521785 = $signed({1'h0, add_521146, array_index_517289[1:0]}) < $signed({1'h0, sel_521149}) ? {add_521146, array_index_517289[1:0]} : sel_521149;
  assign add_521787 = array_index_518210[11:0] + 12'h8e1;
  assign sel_521789 = $signed({1'h0, add_521151}) < $signed({1'h0, sel_521153}) ? add_521151 : sel_521153;
  assign add_521791 = array_index_518213[11:0] + 12'h8e1;
  assign sel_521793 = $signed({1'h0, add_521155}) < $signed({1'h0, sel_521157}) ? add_521155 : sel_521157;
  assign add_521795 = array_index_518710[11:4] + 8'h83;
  assign sel_521798 = $signed({1'h0, add_521159, array_index_518210[3:0]}) < $signed({1'h0, sel_521162}) ? {add_521159, array_index_518210[3:0]} : sel_521162;
  assign add_521800 = array_index_518713[11:4] + 8'h83;
  assign sel_521803 = $signed({1'h0, add_521164, array_index_518213[3:0]}) < $signed({1'h0, sel_521167}) ? {add_521164, array_index_518213[3:0]} : sel_521167;
  assign add_521805 = array_index_519236[11:0] + 12'ha09;
  assign sel_521807 = $signed({1'h0, add_521169}) < $signed({1'h0, sel_521171}) ? add_521169 : sel_521171;
  assign add_521809 = array_index_519239[11:0] + 12'ha09;
  assign sel_521811 = $signed({1'h0, add_521173}) < $signed({1'h0, sel_521175}) ? add_521173 : sel_521175;
  assign add_521813 = array_index_519786[11:1] + 11'h6cb;
  assign sel_521815 = $signed({1'h0, add_521177, array_index_519236[0]}) < $signed({1'h0, sel_521179}) ? {add_521177, array_index_519236[0]} : sel_521179;
  assign add_521817 = array_index_519789[11:1] + 11'h6cb;
  assign sel_521819 = $signed({1'h0, add_521181, array_index_519239[0]}) < $signed({1'h0, sel_521183}) ? {add_521181, array_index_519239[0]} : sel_521183;
  assign add_521821 = array_index_520362[11:1] + 11'h75d;
  assign sel_521823 = $signed({1'h0, add_521185, array_index_519786[0]}) < $signed({1'h0, sel_521187}) ? {add_521185, array_index_519786[0]} : sel_521187;
  assign add_521825 = array_index_520365[11:1] + 11'h75d;
  assign sel_521827 = $signed({1'h0, add_521189, array_index_519789[0]}) < $signed({1'h0, sel_521191}) ? {add_521189, array_index_519789[0]} : sel_521191;
  assign add_521829 = array_index_520964[11:1] + 11'h24f;
  assign sel_521832 = $signed({1'h0, add_521193, array_index_520362[0]}) < $signed({1'h0, sel_521196}) ? {add_521193, array_index_520362[0]} : sel_521196;
  assign add_521834 = array_index_520967[11:1] + 11'h24f;
  assign sel_521837 = $signed({1'h0, add_521198, array_index_520365[0]}) < $signed({1'h0, sel_521201}) ? {add_521198, array_index_520365[0]} : sel_521201;
  assign add_521851 = array_index_512834[11:3] + 9'h1f1;
  assign sel_521853 = $signed({1'h0, add_521209, array_index_512818[2:0]}) < $signed(13'h0fff) ? {add_521209, array_index_512818[2:0]} : 12'hfff;
  assign add_521855 = array_index_512837[11:3] + 9'h1f1;
  assign sel_521857 = $signed({1'h0, add_521211, array_index_512819[2:0]}) < $signed(13'h0fff) ? {add_521211, array_index_512819[2:0]} : 12'hfff;
  assign add_521867 = array_index_512942[11:0] + 12'h081;
  assign sel_521869 = $signed({1'h0, add_521223}) < $signed({1'h0, sel_521225}) ? add_521223 : sel_521225;
  assign add_521871 = array_index_512945[11:0] + 12'h081;
  assign sel_521873 = $signed({1'h0, add_521227}) < $signed({1'h0, sel_521229}) ? add_521227 : sel_521229;
  assign add_521885 = array_index_513120[11:0] + 12'h0b1;
  assign sel_521887 = $signed({1'h0, add_521241}) < $signed({1'h0, sel_521243}) ? add_521241 : sel_521243;
  assign add_521889 = array_index_513123[11:0] + 12'h0b1;
  assign sel_521891 = $signed({1'h0, add_521245}) < $signed({1'h0, sel_521247}) ? add_521245 : sel_521247;
  assign add_521903 = array_index_513374[11:1] + 11'h4c1;
  assign sel_521905 = $signed({1'h0, add_521259, array_index_513238[0]}) < $signed({1'h0, sel_521261}) ? {add_521259, array_index_513238[0]} : sel_521261;
  assign add_521907 = array_index_513377[11:1] + 11'h4c1;
  assign sel_521909 = $signed({1'h0, add_521263, array_index_513241[0]}) < $signed({1'h0, sel_521265}) ? {add_521263, array_index_513241[0]} : sel_521265;
  assign add_521919 = array_index_513702[11:0] + 12'hbb1;
  assign sel_521921 = $signed({1'h0, add_521275}) < $signed({1'h0, sel_521277}) ? add_521275 : sel_521277;
  assign add_521923 = array_index_513705[11:0] + 12'hbb1;
  assign sel_521925 = $signed({1'h0, add_521279}) < $signed({1'h0, sel_521281}) ? add_521279 : sel_521281;
  assign add_521935 = array_index_514096[11:0] + 12'h6ab;
  assign sel_521937 = $signed({1'h0, add_521291}) < $signed({1'h0, sel_521293}) ? add_521291 : sel_521293;
  assign add_521939 = array_index_514099[11:0] + 12'h6ab;
  assign sel_521941 = $signed({1'h0, add_521295}) < $signed({1'h0, sel_521297}) ? add_521295 : sel_521297;
  assign add_521951 = array_index_514558[11:0] + 12'h7d5;
  assign sel_521953 = $signed({1'h0, add_521307}) < $signed({1'h0, sel_521309}) ? add_521307 : sel_521309;
  assign add_521955 = array_index_514561[11:0] + 12'h7d5;
  assign sel_521957 = $signed({1'h0, add_521311}) < $signed({1'h0, sel_521313}) ? add_521311 : sel_521313;
  assign add_522025 = array_index_521590[11:0] + 12'h62b;
  assign sel_522027 = $signed({1'h0, add_521382}) < $signed({1'h0, sel_521384}) ? add_521382 : sel_521384;
  assign add_522029 = array_index_521593[11:0] + 12'h62b;
  assign sel_522031 = $signed({1'h0, add_521387}) < $signed({1'h0, sel_521389}) ? add_521387 : sel_521389;
  assign add_522033 = array_index_512818[11:2] + 10'h181;
  assign add_522035 = array_index_512819[11:2] + 10'h181;
  assign add_522049 = array_index_512880[11:0] + 12'h8a7;
  assign sel_522051 = $signed({1'h0, add_521397}) < $signed({1'h0, sel_521399}) ? add_521397 : sel_521399;
  assign add_522053 = array_index_512883[11:0] + 12'h8a7;
  assign sel_522055 = $signed({1'h0, add_521401}) < $signed({1'h0, sel_521403}) ? add_521401 : sel_521403;
  assign add_522067 = array_index_513022[11:1] + 11'h283;
  assign sel_522069 = $signed({1'h0, add_521415, array_index_512942[0]}) < $signed({1'h0, sel_521417}) ? {add_521415, array_index_512942[0]} : sel_521417;
  assign add_522071 = array_index_513025[11:1] + 11'h283;
  assign sel_522073 = $signed({1'h0, add_521419, array_index_512945[0]}) < $signed({1'h0, sel_521421}) ? {add_521419, array_index_512945[0]} : sel_521421;
  assign add_522083 = array_index_513238[11:1] + 11'h44d;
  assign sel_522085 = $signed({1'h0, add_521431, array_index_513120[0]}) < $signed({1'h0, sel_521433}) ? {add_521431, array_index_513120[0]} : sel_521433;
  assign add_522087 = array_index_513241[11:1] + 11'h44d;
  assign sel_522089 = $signed({1'h0, add_521435, array_index_513123[0]}) < $signed({1'h0, sel_521437}) ? {add_521435, array_index_513123[0]} : sel_521437;
  assign add_522099 = array_index_513530[11:0] + 12'hcb1;
  assign sel_522101 = $signed({1'h0, add_521447}) < $signed({1'h0, sel_521449}) ? add_521447 : sel_521449;
  assign add_522103 = array_index_513533[11:0] + 12'hcb1;
  assign sel_522105 = $signed({1'h0, add_521451}) < $signed({1'h0, sel_521453}) ? add_521451 : sel_521453;
  assign add_522115 = array_index_513890[11:0] + 12'h81f;
  assign sel_522117 = $signed({1'h0, add_521463}) < $signed({1'h0, sel_521465}) ? add_521463 : sel_521465;
  assign add_522119 = array_index_513893[11:0] + 12'h81f;
  assign sel_522121 = $signed({1'h0, add_521467}) < $signed({1'h0, sel_521469}) ? add_521467 : sel_521469;
  assign add_522131 = array_index_514318[11:0] + 12'h45b;
  assign sel_522133 = $signed({1'h0, add_521479}) < $signed({1'h0, sel_521481}) ? add_521479 : sel_521481;
  assign add_522135 = array_index_514321[11:0] + 12'h45b;
  assign sel_522137 = $signed({1'h0, add_521483}) < $signed({1'h0, sel_521485}) ? add_521483 : sel_521485;
  assign add_522149 = array_index_514818[11:3] + 9'h0f5;
  assign sel_522151 = $signed({1'h0, add_521497, array_index_514558[2:0]}) < $signed({1'h0, sel_521499}) ? {add_521497, array_index_514558[2:0]} : sel_521499;
  assign add_522153 = array_index_514821[11:3] + 9'h0f5;
  assign sel_522155 = $signed({1'h0, add_521501, array_index_514561[2:0]}) < $signed({1'h0, sel_521503}) ? {add_521501, array_index_514561[2:0]} : sel_521503;
  assign add_522253 = array_index_512834[11:3] + 9'h12f;
  assign sel_522255 = $signed({1'h0, add_521597, array_index_512818[2:0]}) < $signed(13'h0fff) ? {add_521597, array_index_512818[2:0]} : 12'hfff;
  assign add_522257 = array_index_512837[11:3] + 9'h12f;
  assign sel_522259 = $signed({1'h0, add_521599, array_index_512819[2:0]}) < $signed(13'h0fff) ? {add_521599, array_index_512819[2:0]} : 12'hfff;
  assign add_522271 = array_index_512942[11:3] + 9'h171;
  assign sel_522273 = $signed({1'h0, add_521613, array_index_512880[2:0]}) < $signed({1'h0, sel_521615}) ? {add_521613, array_index_512880[2:0]} : sel_521615;
  assign add_522275 = array_index_512945[11:3] + 9'h171;
  assign sel_522277 = $signed({1'h0, add_521617, array_index_512883[2:0]}) < $signed({1'h0, sel_521619}) ? {add_521617, array_index_512883[2:0]} : sel_521619;
  assign add_522287 = array_index_513120[11:0] + 12'h091;
  assign sel_522289 = $signed({1'h0, add_521629}) < $signed({1'h0, sel_521631}) ? add_521629 : sel_521631;
  assign add_522291 = array_index_513123[11:0] + 12'h091;
  assign sel_522293 = $signed({1'h0, add_521633}) < $signed({1'h0, sel_521635}) ? add_521633 : sel_521635;
  assign add_522303 = array_index_513374[11:0] + 12'hf59;
  assign sel_522305 = $signed({1'h0, add_521645}) < $signed({1'h0, sel_521647}) ? add_521645 : sel_521647;
  assign add_522307 = array_index_513377[11:0] + 12'hf59;
  assign sel_522309 = $signed({1'h0, add_521649}) < $signed({1'h0, sel_521651}) ? add_521649 : sel_521651;
  assign add_522321 = array_index_513702[11:0] + 12'h437;
  assign sel_522323 = $signed({1'h0, add_521663}) < $signed({1'h0, sel_521665}) ? add_521663 : sel_521665;
  assign add_522325 = array_index_513705[11:0] + 12'h437;
  assign sel_522327 = $signed({1'h0, add_521667}) < $signed({1'h0, sel_521669}) ? add_521667 : sel_521669;
  assign add_522337 = array_index_514096[11:0] + 12'hee1;
  assign sel_522339 = $signed({1'h0, add_521679}) < $signed({1'h0, sel_521681}) ? add_521679 : sel_521681;
  assign add_522341 = array_index_514099[11:0] + 12'hee1;
  assign sel_522343 = $signed({1'h0, add_521683}) < $signed({1'h0, sel_521685}) ? add_521683 : sel_521685;
  assign add_522353 = array_index_514558[11:1] + 11'h179;
  assign sel_522355 = $signed({1'h0, add_521695, array_index_514318[0]}) < $signed({1'h0, sel_521697}) ? {add_521695, array_index_514318[0]} : sel_521697;
  assign add_522357 = array_index_514561[11:1] + 11'h179;
  assign sel_522359 = $signed({1'h0, add_521699, array_index_514321[0]}) < $signed({1'h0, sel_521701}) ? {add_521699, array_index_514321[0]} : sel_521701;
  assign add_522369 = array_index_515098[11:0] + 12'h067;
  assign sel_522371 = $signed({1'h0, add_521711}) < $signed({1'h0, sel_521713}) ? add_521711 : sel_521713;
  assign add_522373 = array_index_515101[11:0] + 12'h067;
  assign sel_522375 = $signed({1'h0, add_521715}) < $signed({1'h0, sel_521717}) ? add_521715 : sel_521717;
  assign add_522377 = array_index_515398[11:3] + 9'h1ef;
  assign sel_522380 = $signed({1'h0, add_521719, array_index_515098[2:0]}) < $signed({1'h0, sel_521722}) ? {add_521719, array_index_515098[2:0]} : sel_521722;
  assign add_522382 = array_index_515401[11:3] + 9'h1ef;
  assign sel_522385 = $signed({1'h0, add_521724, array_index_515101[2:0]}) < $signed({1'h0, sel_521727}) ? {add_521724, array_index_515101[2:0]} : sel_521727;
  assign add_522387 = array_index_515726[11:1] + 11'h2d5;
  assign sel_522389 = $signed({1'h0, add_521729, array_index_515398[0]}) < $signed({1'h0, sel_521731}) ? {add_521729, array_index_515398[0]} : sel_521731;
  assign add_522391 = array_index_515729[11:1] + 11'h2d5;
  assign sel_522393 = $signed({1'h0, add_521733, array_index_515401[0]}) < $signed({1'h0, sel_521735}) ? {add_521733, array_index_515401[0]} : sel_521735;
  assign add_522395 = array_index_516080[11:2] + 10'h353;
  assign sel_522397 = $signed({1'h0, add_521737, array_index_515726[1:0]}) < $signed({1'h0, sel_521739}) ? {add_521737, array_index_515726[1:0]} : sel_521739;
  assign add_522399 = array_index_516083[11:2] + 10'h353;
  assign sel_522401 = $signed({1'h0, add_521741, array_index_515729[1:0]}) < $signed({1'h0, sel_521743}) ? {add_521741, array_index_515729[1:0]} : sel_521743;
  assign add_522403 = array_index_516458[11:0] + 12'h0a7;
  assign sel_522405 = $signed({1'h0, add_521745}) < $signed({1'h0, sel_521747}) ? add_521745 : sel_521747;
  assign add_522407 = array_index_516461[11:0] + 12'h0a7;
  assign sel_522409 = $signed({1'h0, add_521749}) < $signed({1'h0, sel_521751}) ? add_521749 : sel_521751;
  assign add_522411 = array_index_516860[11:1] + 11'h4cb;
  assign sel_522413 = $signed({1'h0, add_521753, array_index_516458[0]}) < $signed({1'h0, sel_521755}) ? {add_521753, array_index_516458[0]} : sel_521755;
  assign add_522415 = array_index_516863[11:1] + 11'h4cb;
  assign sel_522417 = $signed({1'h0, add_521757, array_index_516461[0]}) < $signed({1'h0, sel_521759}) ? {add_521757, array_index_516461[0]} : sel_521759;
  assign add_522419 = array_index_517286[11:0] + 12'hfe9;
  assign sel_522421 = $signed({1'h0, add_521761}) < $signed({1'h0, sel_521763}) ? add_521761 : sel_521763;
  assign add_522423 = array_index_517289[11:0] + 12'hfe9;
  assign sel_522425 = $signed({1'h0, add_521765}) < $signed({1'h0, sel_521767}) ? add_521765 : sel_521767;
  assign add_522427 = array_index_517736[11:0] + 12'h97d;
  assign sel_522429 = $signed({1'h0, add_521769}) < $signed({1'h0, sel_521771}) ? add_521769 : sel_521771;
  assign add_522431 = array_index_517739[11:0] + 12'h97d;
  assign sel_522433 = $signed({1'h0, add_521773}) < $signed({1'h0, sel_521775}) ? add_521773 : sel_521775;
  assign add_522435 = array_index_518210[11:2] + 10'h2bb;
  assign sel_522438 = $signed({1'h0, add_521777, array_index_517736[1:0]}) < $signed({1'h0, sel_521780}) ? {add_521777, array_index_517736[1:0]} : sel_521780;
  assign add_522440 = array_index_518213[11:2] + 10'h2bb;
  assign sel_522443 = $signed({1'h0, add_521782, array_index_517739[1:0]}) < $signed({1'h0, sel_521785}) ? {add_521782, array_index_517739[1:0]} : sel_521785;
  assign add_522445 = array_index_518710[11:0] + 12'h8e1;
  assign sel_522447 = $signed({1'h0, add_521787}) < $signed({1'h0, sel_521789}) ? add_521787 : sel_521789;
  assign add_522449 = array_index_518713[11:0] + 12'h8e1;
  assign sel_522451 = $signed({1'h0, add_521791}) < $signed({1'h0, sel_521793}) ? add_521791 : sel_521793;
  assign add_522453 = array_index_519236[11:4] + 8'h83;
  assign sel_522456 = $signed({1'h0, add_521795, array_index_518710[3:0]}) < $signed({1'h0, sel_521798}) ? {add_521795, array_index_518710[3:0]} : sel_521798;
  assign add_522458 = array_index_519239[11:4] + 8'h83;
  assign sel_522461 = $signed({1'h0, add_521800, array_index_518713[3:0]}) < $signed({1'h0, sel_521803}) ? {add_521800, array_index_518713[3:0]} : sel_521803;
  assign add_522463 = array_index_519786[11:0] + 12'ha09;
  assign sel_522465 = $signed({1'h0, add_521805}) < $signed({1'h0, sel_521807}) ? add_521805 : sel_521807;
  assign add_522467 = array_index_519789[11:0] + 12'ha09;
  assign sel_522469 = $signed({1'h0, add_521809}) < $signed({1'h0, sel_521811}) ? add_521809 : sel_521811;
  assign add_522471 = array_index_520362[11:1] + 11'h6cb;
  assign sel_522473 = $signed({1'h0, add_521813, array_index_519786[0]}) < $signed({1'h0, sel_521815}) ? {add_521813, array_index_519786[0]} : sel_521815;
  assign add_522475 = array_index_520365[11:1] + 11'h6cb;
  assign sel_522477 = $signed({1'h0, add_521817, array_index_519789[0]}) < $signed({1'h0, sel_521819}) ? {add_521817, array_index_519789[0]} : sel_521819;
  assign add_522479 = array_index_520964[11:1] + 11'h75d;
  assign sel_522481 = $signed({1'h0, add_521821, array_index_520362[0]}) < $signed({1'h0, sel_521823}) ? {add_521821, array_index_520362[0]} : sel_521823;
  assign add_522483 = array_index_520967[11:1] + 11'h75d;
  assign sel_522485 = $signed({1'h0, add_521825, array_index_520365[0]}) < $signed({1'h0, sel_521827}) ? {add_521825, array_index_520365[0]} : sel_521827;
  assign add_522487 = array_index_521590[11:1] + 11'h24f;
  assign sel_522490 = $signed({1'h0, add_521829, array_index_520964[0]}) < $signed({1'h0, sel_521832}) ? {add_521829, array_index_520964[0]} : sel_521832;
  assign add_522492 = array_index_521593[11:1] + 11'h24f;
  assign sel_522495 = $signed({1'h0, add_521834, array_index_520967[0]}) < $signed({1'h0, sel_521837}) ? {add_521834, array_index_520967[0]} : sel_521837;
  assign add_522499 = array_index_512818[11:0] + 12'h70f;
  assign add_522501 = array_index_512819[11:0] + 12'h70f;
  assign add_522515 = array_index_512880[11:3] + 9'h1f1;
  assign sel_522517 = $signed({1'h0, add_521851, array_index_512834[2:0]}) < $signed({1'h0, sel_521853}) ? {add_521851, array_index_512834[2:0]} : sel_521853;
  assign add_522519 = array_index_512883[11:3] + 9'h1f1;
  assign sel_522521 = $signed({1'h0, add_521855, array_index_512837[2:0]}) < $signed({1'h0, sel_521857}) ? {add_521855, array_index_512837[2:0]} : sel_521857;
  assign add_522531 = array_index_513022[11:0] + 12'h081;
  assign sel_522533 = $signed({1'h0, add_521867}) < $signed({1'h0, sel_521869}) ? add_521867 : sel_521869;
  assign add_522535 = array_index_513025[11:0] + 12'h081;
  assign sel_522537 = $signed({1'h0, add_521871}) < $signed({1'h0, sel_521873}) ? add_521871 : sel_521873;
  assign add_522549 = array_index_513238[11:0] + 12'h0b1;
  assign sel_522551 = $signed({1'h0, add_521885}) < $signed({1'h0, sel_521887}) ? add_521885 : sel_521887;
  assign add_522553 = array_index_513241[11:0] + 12'h0b1;
  assign sel_522555 = $signed({1'h0, add_521889}) < $signed({1'h0, sel_521891}) ? add_521889 : sel_521891;
  assign add_522567 = array_index_513530[11:1] + 11'h4c1;
  assign sel_522569 = $signed({1'h0, add_521903, array_index_513374[0]}) < $signed({1'h0, sel_521905}) ? {add_521903, array_index_513374[0]} : sel_521905;
  assign add_522571 = array_index_513533[11:1] + 11'h4c1;
  assign sel_522573 = $signed({1'h0, add_521907, array_index_513377[0]}) < $signed({1'h0, sel_521909}) ? {add_521907, array_index_513377[0]} : sel_521909;
  assign add_522583 = array_index_513890[11:0] + 12'hbb1;
  assign sel_522585 = $signed({1'h0, add_521919}) < $signed({1'h0, sel_521921}) ? add_521919 : sel_521921;
  assign add_522587 = array_index_513893[11:0] + 12'hbb1;
  assign sel_522589 = $signed({1'h0, add_521923}) < $signed({1'h0, sel_521925}) ? add_521923 : sel_521925;
  assign add_522599 = array_index_514318[11:0] + 12'h6ab;
  assign sel_522601 = $signed({1'h0, add_521935}) < $signed({1'h0, sel_521937}) ? add_521935 : sel_521937;
  assign add_522603 = array_index_514321[11:0] + 12'h6ab;
  assign sel_522605 = $signed({1'h0, add_521939}) < $signed({1'h0, sel_521941}) ? add_521939 : sel_521941;
  assign add_522615 = array_index_514818[11:0] + 12'h7d5;
  assign sel_522617 = $signed({1'h0, add_521951}) < $signed({1'h0, sel_521953}) ? add_521951 : sel_521953;
  assign add_522619 = array_index_514821[11:0] + 12'h7d5;
  assign sel_522621 = $signed({1'h0, add_521955}) < $signed({1'h0, sel_521957}) ? add_521955 : sel_521957;
  assign add_522697 = array_index_512834[11:2] + 10'h181;
  assign sel_522699 = $signed({1'h0, add_522033, array_index_512818[1:0]}) < $signed(13'h0fff) ? {add_522033, array_index_512818[1:0]} : 12'hfff;
  assign add_522701 = array_index_512837[11:2] + 10'h181;
  assign sel_522703 = $signed({1'h0, add_522035, array_index_512819[1:0]}) < $signed(13'h0fff) ? {add_522035, array_index_512819[1:0]} : 12'hfff;
  assign add_522715 = array_index_512942[11:0] + 12'h8a7;
  assign sel_522717 = $signed({1'h0, add_522049}) < $signed({1'h0, sel_522051}) ? add_522049 : sel_522051;
  assign add_522719 = array_index_512945[11:0] + 12'h8a7;
  assign sel_522721 = $signed({1'h0, add_522053}) < $signed({1'h0, sel_522055}) ? add_522053 : sel_522055;
  assign add_522733 = array_index_513120[11:1] + 11'h283;
  assign sel_522735 = $signed({1'h0, add_522067, array_index_513022[0]}) < $signed({1'h0, sel_522069}) ? {add_522067, array_index_513022[0]} : sel_522069;
  assign add_522737 = array_index_513123[11:1] + 11'h283;
  assign sel_522739 = $signed({1'h0, add_522071, array_index_513025[0]}) < $signed({1'h0, sel_522073}) ? {add_522071, array_index_513025[0]} : sel_522073;
  assign add_522749 = array_index_513374[11:1] + 11'h44d;
  assign sel_522751 = $signed({1'h0, add_522083, array_index_513238[0]}) < $signed({1'h0, sel_522085}) ? {add_522083, array_index_513238[0]} : sel_522085;
  assign add_522753 = array_index_513377[11:1] + 11'h44d;
  assign sel_522755 = $signed({1'h0, add_522087, array_index_513241[0]}) < $signed({1'h0, sel_522089}) ? {add_522087, array_index_513241[0]} : sel_522089;
  assign add_522765 = array_index_513702[11:0] + 12'hcb1;
  assign sel_522767 = $signed({1'h0, add_522099}) < $signed({1'h0, sel_522101}) ? add_522099 : sel_522101;
  assign add_522769 = array_index_513705[11:0] + 12'hcb1;
  assign sel_522771 = $signed({1'h0, add_522103}) < $signed({1'h0, sel_522105}) ? add_522103 : sel_522105;
  assign add_522781 = array_index_514096[11:0] + 12'h81f;
  assign sel_522783 = $signed({1'h0, add_522115}) < $signed({1'h0, sel_522117}) ? add_522115 : sel_522117;
  assign add_522785 = array_index_514099[11:0] + 12'h81f;
  assign sel_522787 = $signed({1'h0, add_522119}) < $signed({1'h0, sel_522121}) ? add_522119 : sel_522121;
  assign add_522797 = array_index_514558[11:0] + 12'h45b;
  assign sel_522799 = $signed({1'h0, add_522131}) < $signed({1'h0, sel_522133}) ? add_522131 : sel_522133;
  assign add_522801 = array_index_514561[11:0] + 12'h45b;
  assign sel_522803 = $signed({1'h0, add_522135}) < $signed({1'h0, sel_522137}) ? add_522135 : sel_522137;
  assign add_522815 = array_index_515098[11:3] + 9'h0f5;
  assign sel_522817 = $signed({1'h0, add_522149, array_index_514818[2:0]}) < $signed({1'h0, sel_522151}) ? {add_522149, array_index_514818[2:0]} : sel_522151;
  assign add_522819 = array_index_515101[11:3] + 9'h0f5;
  assign sel_522821 = $signed({1'h0, add_522153, array_index_514821[2:0]}) < $signed({1'h0, sel_522155}) ? {add_522153, array_index_514821[2:0]} : sel_522155;
  assign add_522907 = array_index_512818[11:1] + 11'h109;
  assign add_522909 = array_index_512819[11:1] + 11'h109;
  assign add_522921 = array_index_512880[11:3] + 9'h12f;
  assign sel_522923 = $signed({1'h0, add_522253, array_index_512834[2:0]}) < $signed({1'h0, sel_522255}) ? {add_522253, array_index_512834[2:0]} : sel_522255;
  assign add_522925 = array_index_512883[11:3] + 9'h12f;
  assign sel_522927 = $signed({1'h0, add_522257, array_index_512837[2:0]}) < $signed({1'h0, sel_522259}) ? {add_522257, array_index_512837[2:0]} : sel_522259;
  assign add_522939 = array_index_513022[11:3] + 9'h171;
  assign sel_522941 = $signed({1'h0, add_522271, array_index_512942[2:0]}) < $signed({1'h0, sel_522273}) ? {add_522271, array_index_512942[2:0]} : sel_522273;
  assign add_522943 = array_index_513025[11:3] + 9'h171;
  assign sel_522945 = $signed({1'h0, add_522275, array_index_512945[2:0]}) < $signed({1'h0, sel_522277}) ? {add_522275, array_index_512945[2:0]} : sel_522277;
  assign add_522955 = array_index_513238[11:0] + 12'h091;
  assign sel_522957 = $signed({1'h0, add_522287}) < $signed({1'h0, sel_522289}) ? add_522287 : sel_522289;
  assign add_522959 = array_index_513241[11:0] + 12'h091;
  assign sel_522961 = $signed({1'h0, add_522291}) < $signed({1'h0, sel_522293}) ? add_522291 : sel_522293;
  assign add_522971 = array_index_513530[11:0] + 12'hf59;
  assign sel_522973 = $signed({1'h0, add_522303}) < $signed({1'h0, sel_522305}) ? add_522303 : sel_522305;
  assign add_522975 = array_index_513533[11:0] + 12'hf59;
  assign sel_522977 = $signed({1'h0, add_522307}) < $signed({1'h0, sel_522309}) ? add_522307 : sel_522309;
  assign add_522989 = array_index_513890[11:0] + 12'h437;
  assign sel_522991 = $signed({1'h0, add_522321}) < $signed({1'h0, sel_522323}) ? add_522321 : sel_522323;
  assign add_522993 = array_index_513893[11:0] + 12'h437;
  assign sel_522995 = $signed({1'h0, add_522325}) < $signed({1'h0, sel_522327}) ? add_522325 : sel_522327;
  assign add_523005 = array_index_514318[11:0] + 12'hee1;
  assign sel_523007 = $signed({1'h0, add_522337}) < $signed({1'h0, sel_522339}) ? add_522337 : sel_522339;
  assign add_523009 = array_index_514321[11:0] + 12'hee1;
  assign sel_523011 = $signed({1'h0, add_522341}) < $signed({1'h0, sel_522343}) ? add_522341 : sel_522343;
  assign add_523021 = array_index_514818[11:1] + 11'h179;
  assign sel_523023 = $signed({1'h0, add_522353, array_index_514558[0]}) < $signed({1'h0, sel_522355}) ? {add_522353, array_index_514558[0]} : sel_522355;
  assign add_523025 = array_index_514821[11:1] + 11'h179;
  assign sel_523027 = $signed({1'h0, add_522357, array_index_514561[0]}) < $signed({1'h0, sel_522359}) ? {add_522357, array_index_514561[0]} : sel_522359;
  assign add_523037 = array_index_515398[11:0] + 12'h067;
  assign sel_523039 = $signed({1'h0, add_522369}) < $signed({1'h0, sel_522371}) ? add_522369 : sel_522371;
  assign add_523041 = array_index_515401[11:0] + 12'h067;
  assign sel_523043 = $signed({1'h0, add_522373}) < $signed({1'h0, sel_522375}) ? add_522373 : sel_522375;
  assign add_523045 = array_index_515726[11:3] + 9'h1ef;
  assign sel_523048 = $signed({1'h0, add_522377, array_index_515398[2:0]}) < $signed({1'h0, sel_522380}) ? {add_522377, array_index_515398[2:0]} : sel_522380;
  assign add_523050 = array_index_515729[11:3] + 9'h1ef;
  assign sel_523053 = $signed({1'h0, add_522382, array_index_515401[2:0]}) < $signed({1'h0, sel_522385}) ? {add_522382, array_index_515401[2:0]} : sel_522385;
  assign add_523055 = array_index_516080[11:1] + 11'h2d5;
  assign sel_523057 = $signed({1'h0, add_522387, array_index_515726[0]}) < $signed({1'h0, sel_522389}) ? {add_522387, array_index_515726[0]} : sel_522389;
  assign add_523059 = array_index_516083[11:1] + 11'h2d5;
  assign sel_523061 = $signed({1'h0, add_522391, array_index_515729[0]}) < $signed({1'h0, sel_522393}) ? {add_522391, array_index_515729[0]} : sel_522393;
  assign add_523063 = array_index_516458[11:2] + 10'h353;
  assign sel_523065 = $signed({1'h0, add_522395, array_index_516080[1:0]}) < $signed({1'h0, sel_522397}) ? {add_522395, array_index_516080[1:0]} : sel_522397;
  assign add_523067 = array_index_516461[11:2] + 10'h353;
  assign sel_523069 = $signed({1'h0, add_522399, array_index_516083[1:0]}) < $signed({1'h0, sel_522401}) ? {add_522399, array_index_516083[1:0]} : sel_522401;
  assign add_523071 = array_index_516860[11:0] + 12'h0a7;
  assign sel_523073 = $signed({1'h0, add_522403}) < $signed({1'h0, sel_522405}) ? add_522403 : sel_522405;
  assign add_523075 = array_index_516863[11:0] + 12'h0a7;
  assign sel_523077 = $signed({1'h0, add_522407}) < $signed({1'h0, sel_522409}) ? add_522407 : sel_522409;
  assign add_523079 = array_index_517286[11:1] + 11'h4cb;
  assign sel_523081 = $signed({1'h0, add_522411, array_index_516860[0]}) < $signed({1'h0, sel_522413}) ? {add_522411, array_index_516860[0]} : sel_522413;
  assign add_523083 = array_index_517289[11:1] + 11'h4cb;
  assign sel_523085 = $signed({1'h0, add_522415, array_index_516863[0]}) < $signed({1'h0, sel_522417}) ? {add_522415, array_index_516863[0]} : sel_522417;
  assign add_523087 = array_index_517736[11:0] + 12'hfe9;
  assign sel_523089 = $signed({1'h0, add_522419}) < $signed({1'h0, sel_522421}) ? add_522419 : sel_522421;
  assign add_523091 = array_index_517739[11:0] + 12'hfe9;
  assign sel_523093 = $signed({1'h0, add_522423}) < $signed({1'h0, sel_522425}) ? add_522423 : sel_522425;
  assign add_523095 = array_index_518210[11:0] + 12'h97d;
  assign sel_523097 = $signed({1'h0, add_522427}) < $signed({1'h0, sel_522429}) ? add_522427 : sel_522429;
  assign add_523099 = array_index_518213[11:0] + 12'h97d;
  assign sel_523101 = $signed({1'h0, add_522431}) < $signed({1'h0, sel_522433}) ? add_522431 : sel_522433;
  assign add_523103 = array_index_518710[11:2] + 10'h2bb;
  assign sel_523106 = $signed({1'h0, add_522435, array_index_518210[1:0]}) < $signed({1'h0, sel_522438}) ? {add_522435, array_index_518210[1:0]} : sel_522438;
  assign add_523108 = array_index_518713[11:2] + 10'h2bb;
  assign sel_523111 = $signed({1'h0, add_522440, array_index_518213[1:0]}) < $signed({1'h0, sel_522443}) ? {add_522440, array_index_518213[1:0]} : sel_522443;
  assign add_523113 = array_index_519236[11:0] + 12'h8e1;
  assign sel_523115 = $signed({1'h0, add_522445}) < $signed({1'h0, sel_522447}) ? add_522445 : sel_522447;
  assign add_523117 = array_index_519239[11:0] + 12'h8e1;
  assign sel_523119 = $signed({1'h0, add_522449}) < $signed({1'h0, sel_522451}) ? add_522449 : sel_522451;
  assign add_523121 = array_index_519786[11:4] + 8'h83;
  assign sel_523124 = $signed({1'h0, add_522453, array_index_519236[3:0]}) < $signed({1'h0, sel_522456}) ? {add_522453, array_index_519236[3:0]} : sel_522456;
  assign add_523126 = array_index_519789[11:4] + 8'h83;
  assign sel_523129 = $signed({1'h0, add_522458, array_index_519239[3:0]}) < $signed({1'h0, sel_522461}) ? {add_522458, array_index_519239[3:0]} : sel_522461;
  assign add_523131 = array_index_520362[11:0] + 12'ha09;
  assign sel_523133 = $signed({1'h0, add_522463}) < $signed({1'h0, sel_522465}) ? add_522463 : sel_522465;
  assign add_523135 = array_index_520365[11:0] + 12'ha09;
  assign sel_523137 = $signed({1'h0, add_522467}) < $signed({1'h0, sel_522469}) ? add_522467 : sel_522469;
  assign add_523139 = array_index_520964[11:1] + 11'h6cb;
  assign sel_523141 = $signed({1'h0, add_522471, array_index_520362[0]}) < $signed({1'h0, sel_522473}) ? {add_522471, array_index_520362[0]} : sel_522473;
  assign add_523143 = array_index_520967[11:1] + 11'h6cb;
  assign sel_523145 = $signed({1'h0, add_522475, array_index_520365[0]}) < $signed({1'h0, sel_522477}) ? {add_522475, array_index_520365[0]} : sel_522477;
  assign add_523147 = array_index_521590[11:1] + 11'h75d;
  assign sel_523149 = $signed({1'h0, add_522479, array_index_520964[0]}) < $signed({1'h0, sel_522481}) ? {add_522479, array_index_520964[0]} : sel_522481;
  assign add_523151 = array_index_521593[11:1] + 11'h75d;
  assign sel_523153 = $signed({1'h0, add_522483, array_index_520967[0]}) < $signed({1'h0, sel_522485}) ? {add_522483, array_index_520967[0]} : sel_522485;
  assign concat_523156 = {1'h0, ($signed({1'h0, add_522025}) < $signed({1'h0, sel_522027}) ? add_522025 : sel_522027) == ($signed({1'h0, add_522029}) < $signed({1'h0, sel_522031}) ? add_522029 : sel_522031)};
  assign add_523165 = array_index_512834[11:0] + 12'h70f;
  assign sel_523167 = $signed({1'h0, add_522499}) < $signed(13'h0fff) ? add_522499 : 12'hfff;
  assign add_523169 = array_index_512837[11:0] + 12'h70f;
  assign sel_523171 = $signed({1'h0, add_522501}) < $signed(13'h0fff) ? add_522501 : 12'hfff;
  assign add_523183 = array_index_512942[11:3] + 9'h1f1;
  assign sel_523185 = $signed({1'h0, add_522515, array_index_512880[2:0]}) < $signed({1'h0, sel_522517}) ? {add_522515, array_index_512880[2:0]} : sel_522517;
  assign add_523187 = array_index_512945[11:3] + 9'h1f1;
  assign sel_523189 = $signed({1'h0, add_522519, array_index_512883[2:0]}) < $signed({1'h0, sel_522521}) ? {add_522519, array_index_512883[2:0]} : sel_522521;
  assign add_523199 = array_index_513120[11:0] + 12'h081;
  assign sel_523201 = $signed({1'h0, add_522531}) < $signed({1'h0, sel_522533}) ? add_522531 : sel_522533;
  assign add_523203 = array_index_513123[11:0] + 12'h081;
  assign sel_523205 = $signed({1'h0, add_522535}) < $signed({1'h0, sel_522537}) ? add_522535 : sel_522537;
  assign add_523217 = array_index_513374[11:0] + 12'h0b1;
  assign sel_523219 = $signed({1'h0, add_522549}) < $signed({1'h0, sel_522551}) ? add_522549 : sel_522551;
  assign add_523221 = array_index_513377[11:0] + 12'h0b1;
  assign sel_523223 = $signed({1'h0, add_522553}) < $signed({1'h0, sel_522555}) ? add_522553 : sel_522555;
  assign add_523235 = array_index_513702[11:1] + 11'h4c1;
  assign sel_523237 = $signed({1'h0, add_522567, array_index_513530[0]}) < $signed({1'h0, sel_522569}) ? {add_522567, array_index_513530[0]} : sel_522569;
  assign add_523239 = array_index_513705[11:1] + 11'h4c1;
  assign sel_523241 = $signed({1'h0, add_522571, array_index_513533[0]}) < $signed({1'h0, sel_522573}) ? {add_522571, array_index_513533[0]} : sel_522573;
  assign add_523251 = array_index_514096[11:0] + 12'hbb1;
  assign sel_523253 = $signed({1'h0, add_522583}) < $signed({1'h0, sel_522585}) ? add_522583 : sel_522585;
  assign add_523255 = array_index_514099[11:0] + 12'hbb1;
  assign sel_523257 = $signed({1'h0, add_522587}) < $signed({1'h0, sel_522589}) ? add_522587 : sel_522589;
  assign add_523267 = array_index_514558[11:0] + 12'h6ab;
  assign sel_523269 = $signed({1'h0, add_522599}) < $signed({1'h0, sel_522601}) ? add_522599 : sel_522601;
  assign add_523271 = array_index_514561[11:0] + 12'h6ab;
  assign sel_523273 = $signed({1'h0, add_522603}) < $signed({1'h0, sel_522605}) ? add_522603 : sel_522605;
  assign add_523283 = array_index_515098[11:0] + 12'h7d5;
  assign sel_523285 = $signed({1'h0, add_522615}) < $signed({1'h0, sel_522617}) ? add_522615 : sel_522617;
  assign add_523287 = array_index_515101[11:0] + 12'h7d5;
  assign sel_523289 = $signed({1'h0, add_522619}) < $signed({1'h0, sel_522621}) ? add_522619 : sel_522621;
  assign add_523353 = concat_523156 + 2'h1;
  assign add_523355 = array_index_512818[11:1] + 11'h075;
  assign add_523357 = array_index_512819[11:1] + 11'h075;
  assign add_523371 = array_index_512880[11:2] + 10'h181;
  assign sel_523373 = $signed({1'h0, add_522697, array_index_512834[1:0]}) < $signed({1'h0, sel_522699}) ? {add_522697, array_index_512834[1:0]} : sel_522699;
  assign add_523375 = array_index_512883[11:2] + 10'h181;
  assign sel_523377 = $signed({1'h0, add_522701, array_index_512837[1:0]}) < $signed({1'h0, sel_522703}) ? {add_522701, array_index_512837[1:0]} : sel_522703;
  assign add_523389 = array_index_513022[11:0] + 12'h8a7;
  assign sel_523391 = $signed({1'h0, add_522715}) < $signed({1'h0, sel_522717}) ? add_522715 : sel_522717;
  assign add_523393 = array_index_513025[11:0] + 12'h8a7;
  assign sel_523395 = $signed({1'h0, add_522719}) < $signed({1'h0, sel_522721}) ? add_522719 : sel_522721;
  assign add_523407 = array_index_513238[11:1] + 11'h283;
  assign sel_523409 = $signed({1'h0, add_522733, array_index_513120[0]}) < $signed({1'h0, sel_522735}) ? {add_522733, array_index_513120[0]} : sel_522735;
  assign add_523411 = array_index_513241[11:1] + 11'h283;
  assign sel_523413 = $signed({1'h0, add_522737, array_index_513123[0]}) < $signed({1'h0, sel_522739}) ? {add_522737, array_index_513123[0]} : sel_522739;
  assign add_523423 = array_index_513530[11:1] + 11'h44d;
  assign sel_523425 = $signed({1'h0, add_522749, array_index_513374[0]}) < $signed({1'h0, sel_522751}) ? {add_522749, array_index_513374[0]} : sel_522751;
  assign add_523427 = array_index_513533[11:1] + 11'h44d;
  assign sel_523429 = $signed({1'h0, add_522753, array_index_513377[0]}) < $signed({1'h0, sel_522755}) ? {add_522753, array_index_513377[0]} : sel_522755;
  assign add_523439 = array_index_513890[11:0] + 12'hcb1;
  assign sel_523441 = $signed({1'h0, add_522765}) < $signed({1'h0, sel_522767}) ? add_522765 : sel_522767;
  assign add_523443 = array_index_513893[11:0] + 12'hcb1;
  assign sel_523445 = $signed({1'h0, add_522769}) < $signed({1'h0, sel_522771}) ? add_522769 : sel_522771;
  assign add_523455 = array_index_514318[11:0] + 12'h81f;
  assign sel_523457 = $signed({1'h0, add_522781}) < $signed({1'h0, sel_522783}) ? add_522781 : sel_522783;
  assign add_523459 = array_index_514321[11:0] + 12'h81f;
  assign sel_523461 = $signed({1'h0, add_522785}) < $signed({1'h0, sel_522787}) ? add_522785 : sel_522787;
  assign add_523471 = array_index_514818[11:0] + 12'h45b;
  assign sel_523473 = $signed({1'h0, add_522797}) < $signed({1'h0, sel_522799}) ? add_522797 : sel_522799;
  assign add_523475 = array_index_514821[11:0] + 12'h45b;
  assign sel_523477 = $signed({1'h0, add_522801}) < $signed({1'h0, sel_522803}) ? add_522801 : sel_522803;
  assign add_523489 = array_index_515398[11:3] + 9'h0f5;
  assign sel_523491 = $signed({1'h0, add_522815, array_index_515098[2:0]}) < $signed({1'h0, sel_522817}) ? {add_522815, array_index_515098[2:0]} : sel_522817;
  assign add_523493 = array_index_515401[11:3] + 9'h0f5;
  assign sel_523495 = $signed({1'h0, add_522819, array_index_515101[2:0]}) < $signed({1'h0, sel_522821}) ? {add_522819, array_index_515101[2:0]} : sel_522821;
  assign add_523581 = array_index_512834[11:1] + 11'h109;
  assign sel_523583 = $signed({1'h0, add_522907, array_index_512818[0]}) < $signed(13'h0fff) ? {add_522907, array_index_512818[0]} : 12'hfff;
  assign add_523585 = array_index_512837[11:1] + 11'h109;
  assign sel_523587 = $signed({1'h0, add_522909, array_index_512819[0]}) < $signed(13'h0fff) ? {add_522909, array_index_512819[0]} : 12'hfff;
  assign add_523597 = array_index_512942[11:3] + 9'h12f;
  assign sel_523599 = $signed({1'h0, add_522921, array_index_512880[2:0]}) < $signed({1'h0, sel_522923}) ? {add_522921, array_index_512880[2:0]} : sel_522923;
  assign add_523601 = array_index_512945[11:3] + 9'h12f;
  assign sel_523603 = $signed({1'h0, add_522925, array_index_512883[2:0]}) < $signed({1'h0, sel_522927}) ? {add_522925, array_index_512883[2:0]} : sel_522927;
  assign add_523615 = array_index_513120[11:3] + 9'h171;
  assign sel_523617 = $signed({1'h0, add_522939, array_index_513022[2:0]}) < $signed({1'h0, sel_522941}) ? {add_522939, array_index_513022[2:0]} : sel_522941;
  assign add_523619 = array_index_513123[11:3] + 9'h171;
  assign sel_523621 = $signed({1'h0, add_522943, array_index_513025[2:0]}) < $signed({1'h0, sel_522945}) ? {add_522943, array_index_513025[2:0]} : sel_522945;
  assign add_523631 = array_index_513374[11:0] + 12'h091;
  assign sel_523633 = $signed({1'h0, add_522955}) < $signed({1'h0, sel_522957}) ? add_522955 : sel_522957;
  assign add_523635 = array_index_513377[11:0] + 12'h091;
  assign sel_523637 = $signed({1'h0, add_522959}) < $signed({1'h0, sel_522961}) ? add_522959 : sel_522961;
  assign add_523647 = array_index_513702[11:0] + 12'hf59;
  assign sel_523649 = $signed({1'h0, add_522971}) < $signed({1'h0, sel_522973}) ? add_522971 : sel_522973;
  assign add_523651 = array_index_513705[11:0] + 12'hf59;
  assign sel_523653 = $signed({1'h0, add_522975}) < $signed({1'h0, sel_522977}) ? add_522975 : sel_522977;
  assign add_523665 = array_index_514096[11:0] + 12'h437;
  assign sel_523667 = $signed({1'h0, add_522989}) < $signed({1'h0, sel_522991}) ? add_522989 : sel_522991;
  assign add_523669 = array_index_514099[11:0] + 12'h437;
  assign sel_523671 = $signed({1'h0, add_522993}) < $signed({1'h0, sel_522995}) ? add_522993 : sel_522995;
  assign add_523681 = array_index_514558[11:0] + 12'hee1;
  assign sel_523683 = $signed({1'h0, add_523005}) < $signed({1'h0, sel_523007}) ? add_523005 : sel_523007;
  assign add_523685 = array_index_514561[11:0] + 12'hee1;
  assign sel_523687 = $signed({1'h0, add_523009}) < $signed({1'h0, sel_523011}) ? add_523009 : sel_523011;
  assign add_523697 = array_index_515098[11:1] + 11'h179;
  assign sel_523699 = $signed({1'h0, add_523021, array_index_514818[0]}) < $signed({1'h0, sel_523023}) ? {add_523021, array_index_514818[0]} : sel_523023;
  assign add_523701 = array_index_515101[11:1] + 11'h179;
  assign sel_523703 = $signed({1'h0, add_523025, array_index_514821[0]}) < $signed({1'h0, sel_523027}) ? {add_523025, array_index_514821[0]} : sel_523027;
  assign add_523713 = array_index_515726[11:0] + 12'h067;
  assign sel_523715 = $signed({1'h0, add_523037}) < $signed({1'h0, sel_523039}) ? add_523037 : sel_523039;
  assign add_523717 = array_index_515729[11:0] + 12'h067;
  assign sel_523719 = $signed({1'h0, add_523041}) < $signed({1'h0, sel_523043}) ? add_523041 : sel_523043;
  assign add_523721 = array_index_516080[11:3] + 9'h1ef;
  assign sel_523724 = $signed({1'h0, add_523045, array_index_515726[2:0]}) < $signed({1'h0, sel_523048}) ? {add_523045, array_index_515726[2:0]} : sel_523048;
  assign add_523726 = array_index_516083[11:3] + 9'h1ef;
  assign sel_523729 = $signed({1'h0, add_523050, array_index_515729[2:0]}) < $signed({1'h0, sel_523053}) ? {add_523050, array_index_515729[2:0]} : sel_523053;
  assign add_523731 = array_index_516458[11:1] + 11'h2d5;
  assign sel_523733 = $signed({1'h0, add_523055, array_index_516080[0]}) < $signed({1'h0, sel_523057}) ? {add_523055, array_index_516080[0]} : sel_523057;
  assign add_523735 = array_index_516461[11:1] + 11'h2d5;
  assign sel_523737 = $signed({1'h0, add_523059, array_index_516083[0]}) < $signed({1'h0, sel_523061}) ? {add_523059, array_index_516083[0]} : sel_523061;
  assign add_523739 = array_index_516860[11:2] + 10'h353;
  assign sel_523741 = $signed({1'h0, add_523063, array_index_516458[1:0]}) < $signed({1'h0, sel_523065}) ? {add_523063, array_index_516458[1:0]} : sel_523065;
  assign add_523743 = array_index_516863[11:2] + 10'h353;
  assign sel_523745 = $signed({1'h0, add_523067, array_index_516461[1:0]}) < $signed({1'h0, sel_523069}) ? {add_523067, array_index_516461[1:0]} : sel_523069;
  assign add_523747 = array_index_517286[11:0] + 12'h0a7;
  assign sel_523749 = $signed({1'h0, add_523071}) < $signed({1'h0, sel_523073}) ? add_523071 : sel_523073;
  assign add_523751 = array_index_517289[11:0] + 12'h0a7;
  assign sel_523753 = $signed({1'h0, add_523075}) < $signed({1'h0, sel_523077}) ? add_523075 : sel_523077;
  assign add_523755 = array_index_517736[11:1] + 11'h4cb;
  assign sel_523757 = $signed({1'h0, add_523079, array_index_517286[0]}) < $signed({1'h0, sel_523081}) ? {add_523079, array_index_517286[0]} : sel_523081;
  assign add_523759 = array_index_517739[11:1] + 11'h4cb;
  assign sel_523761 = $signed({1'h0, add_523083, array_index_517289[0]}) < $signed({1'h0, sel_523085}) ? {add_523083, array_index_517289[0]} : sel_523085;
  assign add_523763 = array_index_518210[11:0] + 12'hfe9;
  assign sel_523765 = $signed({1'h0, add_523087}) < $signed({1'h0, sel_523089}) ? add_523087 : sel_523089;
  assign add_523767 = array_index_518213[11:0] + 12'hfe9;
  assign sel_523769 = $signed({1'h0, add_523091}) < $signed({1'h0, sel_523093}) ? add_523091 : sel_523093;
  assign add_523771 = array_index_518710[11:0] + 12'h97d;
  assign sel_523773 = $signed({1'h0, add_523095}) < $signed({1'h0, sel_523097}) ? add_523095 : sel_523097;
  assign add_523775 = array_index_518713[11:0] + 12'h97d;
  assign sel_523777 = $signed({1'h0, add_523099}) < $signed({1'h0, sel_523101}) ? add_523099 : sel_523101;
  assign add_523779 = array_index_519236[11:2] + 10'h2bb;
  assign sel_523782 = $signed({1'h0, add_523103, array_index_518710[1:0]}) < $signed({1'h0, sel_523106}) ? {add_523103, array_index_518710[1:0]} : sel_523106;
  assign add_523784 = array_index_519239[11:2] + 10'h2bb;
  assign sel_523787 = $signed({1'h0, add_523108, array_index_518713[1:0]}) < $signed({1'h0, sel_523111}) ? {add_523108, array_index_518713[1:0]} : sel_523111;
  assign add_523789 = array_index_519786[11:0] + 12'h8e1;
  assign sel_523791 = $signed({1'h0, add_523113}) < $signed({1'h0, sel_523115}) ? add_523113 : sel_523115;
  assign add_523793 = array_index_519789[11:0] + 12'h8e1;
  assign sel_523795 = $signed({1'h0, add_523117}) < $signed({1'h0, sel_523119}) ? add_523117 : sel_523119;
  assign add_523797 = array_index_520362[11:4] + 8'h83;
  assign sel_523800 = $signed({1'h0, add_523121, array_index_519786[3:0]}) < $signed({1'h0, sel_523124}) ? {add_523121, array_index_519786[3:0]} : sel_523124;
  assign add_523802 = array_index_520365[11:4] + 8'h83;
  assign sel_523805 = $signed({1'h0, add_523126, array_index_519789[3:0]}) < $signed({1'h0, sel_523129}) ? {add_523126, array_index_519789[3:0]} : sel_523129;
  assign add_523807 = array_index_520964[11:0] + 12'ha09;
  assign sel_523809 = $signed({1'h0, add_523131}) < $signed({1'h0, sel_523133}) ? add_523131 : sel_523133;
  assign add_523811 = array_index_520967[11:0] + 12'ha09;
  assign sel_523813 = $signed({1'h0, add_523135}) < $signed({1'h0, sel_523137}) ? add_523135 : sel_523137;
  assign add_523815 = array_index_521590[11:1] + 11'h6cb;
  assign sel_523817 = $signed({1'h0, add_523139, array_index_520964[0]}) < $signed({1'h0, sel_523141}) ? {add_523139, array_index_520964[0]} : sel_523141;
  assign add_523819 = array_index_521593[11:1] + 11'h6cb;
  assign sel_523821 = $signed({1'h0, add_523143, array_index_520967[0]}) < $signed({1'h0, sel_523145}) ? {add_523143, array_index_520967[0]} : sel_523145;
  assign concat_523824 = {1'h0, ($signed({1'h0, add_522487, array_index_521590[0]}) < $signed({1'h0, sel_522490}) ? {add_522487, array_index_521590[0]} : sel_522490) == ($signed({1'h0, add_522492, array_index_521593[0]}) < $signed({1'h0, sel_522495}) ? {add_522492, array_index_521593[0]} : sel_522495) ? add_523353 : concat_523156};
  assign add_523827 = array_index_512818[11:0] + 12'h811;
  assign add_523829 = array_index_512819[11:0] + 12'h811;
  assign add_523843 = array_index_512880[11:0] + 12'h70f;
  assign sel_523845 = $signed({1'h0, add_523165}) < $signed({1'h0, sel_523167}) ? add_523165 : sel_523167;
  assign add_523847 = array_index_512883[11:0] + 12'h70f;
  assign sel_523849 = $signed({1'h0, add_523169}) < $signed({1'h0, sel_523171}) ? add_523169 : sel_523171;
  assign add_523861 = array_index_513022[11:3] + 9'h1f1;
  assign sel_523863 = $signed({1'h0, add_523183, array_index_512942[2:0]}) < $signed({1'h0, sel_523185}) ? {add_523183, array_index_512942[2:0]} : sel_523185;
  assign add_523865 = array_index_513025[11:3] + 9'h1f1;
  assign sel_523867 = $signed({1'h0, add_523187, array_index_512945[2:0]}) < $signed({1'h0, sel_523189}) ? {add_523187, array_index_512945[2:0]} : sel_523189;
  assign add_523877 = array_index_513238[11:0] + 12'h081;
  assign sel_523879 = $signed({1'h0, add_523199}) < $signed({1'h0, sel_523201}) ? add_523199 : sel_523201;
  assign add_523881 = array_index_513241[11:0] + 12'h081;
  assign sel_523883 = $signed({1'h0, add_523203}) < $signed({1'h0, sel_523205}) ? add_523203 : sel_523205;
  assign add_523895 = array_index_513530[11:0] + 12'h0b1;
  assign sel_523897 = $signed({1'h0, add_523217}) < $signed({1'h0, sel_523219}) ? add_523217 : sel_523219;
  assign add_523899 = array_index_513533[11:0] + 12'h0b1;
  assign sel_523901 = $signed({1'h0, add_523221}) < $signed({1'h0, sel_523223}) ? add_523221 : sel_523223;
  assign add_523913 = array_index_513890[11:1] + 11'h4c1;
  assign sel_523915 = $signed({1'h0, add_523235, array_index_513702[0]}) < $signed({1'h0, sel_523237}) ? {add_523235, array_index_513702[0]} : sel_523237;
  assign add_523917 = array_index_513893[11:1] + 11'h4c1;
  assign sel_523919 = $signed({1'h0, add_523239, array_index_513705[0]}) < $signed({1'h0, sel_523241}) ? {add_523239, array_index_513705[0]} : sel_523241;
  assign add_523929 = array_index_514318[11:0] + 12'hbb1;
  assign sel_523931 = $signed({1'h0, add_523251}) < $signed({1'h0, sel_523253}) ? add_523251 : sel_523253;
  assign add_523933 = array_index_514321[11:0] + 12'hbb1;
  assign sel_523935 = $signed({1'h0, add_523255}) < $signed({1'h0, sel_523257}) ? add_523255 : sel_523257;
  assign add_523945 = array_index_514818[11:0] + 12'h6ab;
  assign sel_523947 = $signed({1'h0, add_523267}) < $signed({1'h0, sel_523269}) ? add_523267 : sel_523269;
  assign add_523949 = array_index_514821[11:0] + 12'h6ab;
  assign sel_523951 = $signed({1'h0, add_523271}) < $signed({1'h0, sel_523273}) ? add_523271 : sel_523273;
  assign add_523961 = array_index_515398[11:0] + 12'h7d5;
  assign sel_523963 = $signed({1'h0, add_523283}) < $signed({1'h0, sel_523285}) ? add_523283 : sel_523285;
  assign add_523965 = array_index_515401[11:0] + 12'h7d5;
  assign sel_523967 = $signed({1'h0, add_523287}) < $signed({1'h0, sel_523289}) ? add_523287 : sel_523289;
  assign add_524027 = concat_523824 + 3'h1;
  assign add_524035 = array_index_512834[11:1] + 11'h075;
  assign sel_524037 = $signed({1'h0, add_523355, array_index_512818[0]}) < $signed(13'h0fff) ? {add_523355, array_index_512818[0]} : 12'hfff;
  assign add_524039 = array_index_512837[11:1] + 11'h075;
  assign sel_524041 = $signed({1'h0, add_523357, array_index_512819[0]}) < $signed(13'h0fff) ? {add_523357, array_index_512819[0]} : 12'hfff;
  assign add_524053 = array_index_512942[11:2] + 10'h181;
  assign sel_524055 = $signed({1'h0, add_523371, array_index_512880[1:0]}) < $signed({1'h0, sel_523373}) ? {add_523371, array_index_512880[1:0]} : sel_523373;
  assign add_524057 = array_index_512945[11:2] + 10'h181;
  assign sel_524059 = $signed({1'h0, add_523375, array_index_512883[1:0]}) < $signed({1'h0, sel_523377}) ? {add_523375, array_index_512883[1:0]} : sel_523377;
  assign add_524071 = array_index_513120[11:0] + 12'h8a7;
  assign sel_524073 = $signed({1'h0, add_523389}) < $signed({1'h0, sel_523391}) ? add_523389 : sel_523391;
  assign add_524075 = array_index_513123[11:0] + 12'h8a7;
  assign sel_524077 = $signed({1'h0, add_523393}) < $signed({1'h0, sel_523395}) ? add_523393 : sel_523395;
  assign add_524089 = array_index_513374[11:1] + 11'h283;
  assign sel_524091 = $signed({1'h0, add_523407, array_index_513238[0]}) < $signed({1'h0, sel_523409}) ? {add_523407, array_index_513238[0]} : sel_523409;
  assign add_524093 = array_index_513377[11:1] + 11'h283;
  assign sel_524095 = $signed({1'h0, add_523411, array_index_513241[0]}) < $signed({1'h0, sel_523413}) ? {add_523411, array_index_513241[0]} : sel_523413;
  assign add_524105 = array_index_513702[11:1] + 11'h44d;
  assign sel_524107 = $signed({1'h0, add_523423, array_index_513530[0]}) < $signed({1'h0, sel_523425}) ? {add_523423, array_index_513530[0]} : sel_523425;
  assign add_524109 = array_index_513705[11:1] + 11'h44d;
  assign sel_524111 = $signed({1'h0, add_523427, array_index_513533[0]}) < $signed({1'h0, sel_523429}) ? {add_523427, array_index_513533[0]} : sel_523429;
  assign add_524121 = array_index_514096[11:0] + 12'hcb1;
  assign sel_524123 = $signed({1'h0, add_523439}) < $signed({1'h0, sel_523441}) ? add_523439 : sel_523441;
  assign add_524125 = array_index_514099[11:0] + 12'hcb1;
  assign sel_524127 = $signed({1'h0, add_523443}) < $signed({1'h0, sel_523445}) ? add_523443 : sel_523445;
  assign add_524137 = array_index_514558[11:0] + 12'h81f;
  assign sel_524139 = $signed({1'h0, add_523455}) < $signed({1'h0, sel_523457}) ? add_523455 : sel_523457;
  assign add_524141 = array_index_514561[11:0] + 12'h81f;
  assign sel_524143 = $signed({1'h0, add_523459}) < $signed({1'h0, sel_523461}) ? add_523459 : sel_523461;
  assign add_524153 = array_index_515098[11:0] + 12'h45b;
  assign sel_524155 = $signed({1'h0, add_523471}) < $signed({1'h0, sel_523473}) ? add_523471 : sel_523473;
  assign add_524157 = array_index_515101[11:0] + 12'h45b;
  assign sel_524159 = $signed({1'h0, add_523475}) < $signed({1'h0, sel_523477}) ? add_523475 : sel_523477;
  assign add_524171 = array_index_515726[11:3] + 9'h0f5;
  assign sel_524173 = $signed({1'h0, add_523489, array_index_515398[2:0]}) < $signed({1'h0, sel_523491}) ? {add_523489, array_index_515398[2:0]} : sel_523491;
  assign add_524175 = array_index_515729[11:3] + 9'h0f5;
  assign sel_524177 = $signed({1'h0, add_523493, array_index_515401[2:0]}) < $signed({1'h0, sel_523495}) ? {add_523493, array_index_515401[2:0]} : sel_523495;
  assign add_524251 = array_index_512818[11:0] + 12'h263;
  assign add_524253 = array_index_512819[11:0] + 12'h263;
  assign add_524265 = array_index_512880[11:1] + 11'h109;
  assign sel_524267 = $signed({1'h0, add_523581, array_index_512834[0]}) < $signed({1'h0, sel_523583}) ? {add_523581, array_index_512834[0]} : sel_523583;
  assign add_524269 = array_index_512883[11:1] + 11'h109;
  assign sel_524271 = $signed({1'h0, add_523585, array_index_512837[0]}) < $signed({1'h0, sel_523587}) ? {add_523585, array_index_512837[0]} : sel_523587;
  assign add_524281 = array_index_513022[11:3] + 9'h12f;
  assign sel_524283 = $signed({1'h0, add_523597, array_index_512942[2:0]}) < $signed({1'h0, sel_523599}) ? {add_523597, array_index_512942[2:0]} : sel_523599;
  assign add_524285 = array_index_513025[11:3] + 9'h12f;
  assign sel_524287 = $signed({1'h0, add_523601, array_index_512945[2:0]}) < $signed({1'h0, sel_523603}) ? {add_523601, array_index_512945[2:0]} : sel_523603;
  assign add_524299 = array_index_513238[11:3] + 9'h171;
  assign sel_524301 = $signed({1'h0, add_523615, array_index_513120[2:0]}) < $signed({1'h0, sel_523617}) ? {add_523615, array_index_513120[2:0]} : sel_523617;
  assign add_524303 = array_index_513241[11:3] + 9'h171;
  assign sel_524305 = $signed({1'h0, add_523619, array_index_513123[2:0]}) < $signed({1'h0, sel_523621}) ? {add_523619, array_index_513123[2:0]} : sel_523621;
  assign add_524315 = array_index_513530[11:0] + 12'h091;
  assign sel_524317 = $signed({1'h0, add_523631}) < $signed({1'h0, sel_523633}) ? add_523631 : sel_523633;
  assign add_524319 = array_index_513533[11:0] + 12'h091;
  assign sel_524321 = $signed({1'h0, add_523635}) < $signed({1'h0, sel_523637}) ? add_523635 : sel_523637;
  assign add_524331 = array_index_513890[11:0] + 12'hf59;
  assign sel_524333 = $signed({1'h0, add_523647}) < $signed({1'h0, sel_523649}) ? add_523647 : sel_523649;
  assign add_524335 = array_index_513893[11:0] + 12'hf59;
  assign sel_524337 = $signed({1'h0, add_523651}) < $signed({1'h0, sel_523653}) ? add_523651 : sel_523653;
  assign add_524349 = array_index_514318[11:0] + 12'h437;
  assign sel_524351 = $signed({1'h0, add_523665}) < $signed({1'h0, sel_523667}) ? add_523665 : sel_523667;
  assign add_524353 = array_index_514321[11:0] + 12'h437;
  assign sel_524355 = $signed({1'h0, add_523669}) < $signed({1'h0, sel_523671}) ? add_523669 : sel_523671;
  assign add_524365 = array_index_514818[11:0] + 12'hee1;
  assign sel_524367 = $signed({1'h0, add_523681}) < $signed({1'h0, sel_523683}) ? add_523681 : sel_523683;
  assign add_524369 = array_index_514821[11:0] + 12'hee1;
  assign sel_524371 = $signed({1'h0, add_523685}) < $signed({1'h0, sel_523687}) ? add_523685 : sel_523687;
  assign add_524381 = array_index_515398[11:1] + 11'h179;
  assign sel_524383 = $signed({1'h0, add_523697, array_index_515098[0]}) < $signed({1'h0, sel_523699}) ? {add_523697, array_index_515098[0]} : sel_523699;
  assign add_524385 = array_index_515401[11:1] + 11'h179;
  assign sel_524387 = $signed({1'h0, add_523701, array_index_515101[0]}) < $signed({1'h0, sel_523703}) ? {add_523701, array_index_515101[0]} : sel_523703;
  assign add_524397 = array_index_516080[11:0] + 12'h067;
  assign sel_524399 = $signed({1'h0, add_523713}) < $signed({1'h0, sel_523715}) ? add_523713 : sel_523715;
  assign add_524401 = array_index_516083[11:0] + 12'h067;
  assign sel_524403 = $signed({1'h0, add_523717}) < $signed({1'h0, sel_523719}) ? add_523717 : sel_523719;
  assign add_524405 = array_index_516458[11:3] + 9'h1ef;
  assign sel_524408 = $signed({1'h0, add_523721, array_index_516080[2:0]}) < $signed({1'h0, sel_523724}) ? {add_523721, array_index_516080[2:0]} : sel_523724;
  assign add_524410 = array_index_516461[11:3] + 9'h1ef;
  assign sel_524413 = $signed({1'h0, add_523726, array_index_516083[2:0]}) < $signed({1'h0, sel_523729}) ? {add_523726, array_index_516083[2:0]} : sel_523729;
  assign add_524415 = array_index_516860[11:1] + 11'h2d5;
  assign sel_524417 = $signed({1'h0, add_523731, array_index_516458[0]}) < $signed({1'h0, sel_523733}) ? {add_523731, array_index_516458[0]} : sel_523733;
  assign add_524419 = array_index_516863[11:1] + 11'h2d5;
  assign sel_524421 = $signed({1'h0, add_523735, array_index_516461[0]}) < $signed({1'h0, sel_523737}) ? {add_523735, array_index_516461[0]} : sel_523737;
  assign add_524423 = array_index_517286[11:2] + 10'h353;
  assign sel_524425 = $signed({1'h0, add_523739, array_index_516860[1:0]}) < $signed({1'h0, sel_523741}) ? {add_523739, array_index_516860[1:0]} : sel_523741;
  assign add_524427 = array_index_517289[11:2] + 10'h353;
  assign sel_524429 = $signed({1'h0, add_523743, array_index_516863[1:0]}) < $signed({1'h0, sel_523745}) ? {add_523743, array_index_516863[1:0]} : sel_523745;
  assign add_524431 = array_index_517736[11:0] + 12'h0a7;
  assign sel_524433 = $signed({1'h0, add_523747}) < $signed({1'h0, sel_523749}) ? add_523747 : sel_523749;
  assign add_524435 = array_index_517739[11:0] + 12'h0a7;
  assign sel_524437 = $signed({1'h0, add_523751}) < $signed({1'h0, sel_523753}) ? add_523751 : sel_523753;
  assign add_524439 = array_index_518210[11:1] + 11'h4cb;
  assign sel_524441 = $signed({1'h0, add_523755, array_index_517736[0]}) < $signed({1'h0, sel_523757}) ? {add_523755, array_index_517736[0]} : sel_523757;
  assign add_524443 = array_index_518213[11:1] + 11'h4cb;
  assign sel_524445 = $signed({1'h0, add_523759, array_index_517739[0]}) < $signed({1'h0, sel_523761}) ? {add_523759, array_index_517739[0]} : sel_523761;
  assign add_524447 = array_index_518710[11:0] + 12'hfe9;
  assign sel_524449 = $signed({1'h0, add_523763}) < $signed({1'h0, sel_523765}) ? add_523763 : sel_523765;
  assign add_524451 = array_index_518713[11:0] + 12'hfe9;
  assign sel_524453 = $signed({1'h0, add_523767}) < $signed({1'h0, sel_523769}) ? add_523767 : sel_523769;
  assign add_524455 = array_index_519236[11:0] + 12'h97d;
  assign sel_524457 = $signed({1'h0, add_523771}) < $signed({1'h0, sel_523773}) ? add_523771 : sel_523773;
  assign add_524459 = array_index_519239[11:0] + 12'h97d;
  assign sel_524461 = $signed({1'h0, add_523775}) < $signed({1'h0, sel_523777}) ? add_523775 : sel_523777;
  assign add_524463 = array_index_519786[11:2] + 10'h2bb;
  assign sel_524466 = $signed({1'h0, add_523779, array_index_519236[1:0]}) < $signed({1'h0, sel_523782}) ? {add_523779, array_index_519236[1:0]} : sel_523782;
  assign add_524468 = array_index_519789[11:2] + 10'h2bb;
  assign sel_524471 = $signed({1'h0, add_523784, array_index_519239[1:0]}) < $signed({1'h0, sel_523787}) ? {add_523784, array_index_519239[1:0]} : sel_523787;
  assign add_524473 = array_index_520362[11:0] + 12'h8e1;
  assign sel_524475 = $signed({1'h0, add_523789}) < $signed({1'h0, sel_523791}) ? add_523789 : sel_523791;
  assign add_524477 = array_index_520365[11:0] + 12'h8e1;
  assign sel_524479 = $signed({1'h0, add_523793}) < $signed({1'h0, sel_523795}) ? add_523793 : sel_523795;
  assign add_524481 = array_index_520964[11:4] + 8'h83;
  assign sel_524484 = $signed({1'h0, add_523797, array_index_520362[3:0]}) < $signed({1'h0, sel_523800}) ? {add_523797, array_index_520362[3:0]} : sel_523800;
  assign add_524486 = array_index_520967[11:4] + 8'h83;
  assign sel_524489 = $signed({1'h0, add_523802, array_index_520365[3:0]}) < $signed({1'h0, sel_523805}) ? {add_523802, array_index_520365[3:0]} : sel_523805;
  assign add_524491 = array_index_521590[11:0] + 12'ha09;
  assign sel_524493 = $signed({1'h0, add_523807}) < $signed({1'h0, sel_523809}) ? add_523807 : sel_523809;
  assign add_524495 = array_index_521593[11:0] + 12'ha09;
  assign sel_524497 = $signed({1'h0, add_523811}) < $signed({1'h0, sel_523813}) ? add_523811 : sel_523813;
  assign concat_524500 = {1'h0, ($signed({1'h0, add_523147, array_index_521590[0]}) < $signed({1'h0, sel_523149}) ? {add_523147, array_index_521590[0]} : sel_523149) == ($signed({1'h0, add_523151, array_index_521593[0]}) < $signed({1'h0, sel_523153}) ? {add_523151, array_index_521593[0]} : sel_523153) ? add_524027 : concat_523824};
  assign add_524509 = array_index_512834[11:0] + 12'h811;
  assign sel_524511 = $signed({1'h0, add_523827}) < $signed(13'h0fff) ? add_523827 : 12'hfff;
  assign add_524513 = array_index_512837[11:0] + 12'h811;
  assign sel_524515 = $signed({1'h0, add_523829}) < $signed(13'h0fff) ? add_523829 : 12'hfff;
  assign add_524527 = array_index_512942[11:0] + 12'h70f;
  assign sel_524529 = $signed({1'h0, add_523843}) < $signed({1'h0, sel_523845}) ? add_523843 : sel_523845;
  assign add_524531 = array_index_512945[11:0] + 12'h70f;
  assign sel_524533 = $signed({1'h0, add_523847}) < $signed({1'h0, sel_523849}) ? add_523847 : sel_523849;
  assign add_524545 = array_index_513120[11:3] + 9'h1f1;
  assign sel_524547 = $signed({1'h0, add_523861, array_index_513022[2:0]}) < $signed({1'h0, sel_523863}) ? {add_523861, array_index_513022[2:0]} : sel_523863;
  assign add_524549 = array_index_513123[11:3] + 9'h1f1;
  assign sel_524551 = $signed({1'h0, add_523865, array_index_513025[2:0]}) < $signed({1'h0, sel_523867}) ? {add_523865, array_index_513025[2:0]} : sel_523867;
  assign add_524561 = array_index_513374[11:0] + 12'h081;
  assign sel_524563 = $signed({1'h0, add_523877}) < $signed({1'h0, sel_523879}) ? add_523877 : sel_523879;
  assign add_524565 = array_index_513377[11:0] + 12'h081;
  assign sel_524567 = $signed({1'h0, add_523881}) < $signed({1'h0, sel_523883}) ? add_523881 : sel_523883;
  assign add_524579 = array_index_513702[11:0] + 12'h0b1;
  assign sel_524581 = $signed({1'h0, add_523895}) < $signed({1'h0, sel_523897}) ? add_523895 : sel_523897;
  assign add_524583 = array_index_513705[11:0] + 12'h0b1;
  assign sel_524585 = $signed({1'h0, add_523899}) < $signed({1'h0, sel_523901}) ? add_523899 : sel_523901;
  assign add_524597 = array_index_514096[11:1] + 11'h4c1;
  assign sel_524599 = $signed({1'h0, add_523913, array_index_513890[0]}) < $signed({1'h0, sel_523915}) ? {add_523913, array_index_513890[0]} : sel_523915;
  assign add_524601 = array_index_514099[11:1] + 11'h4c1;
  assign sel_524603 = $signed({1'h0, add_523917, array_index_513893[0]}) < $signed({1'h0, sel_523919}) ? {add_523917, array_index_513893[0]} : sel_523919;
  assign add_524613 = array_index_514558[11:0] + 12'hbb1;
  assign sel_524615 = $signed({1'h0, add_523929}) < $signed({1'h0, sel_523931}) ? add_523929 : sel_523931;
  assign add_524617 = array_index_514561[11:0] + 12'hbb1;
  assign sel_524619 = $signed({1'h0, add_523933}) < $signed({1'h0, sel_523935}) ? add_523933 : sel_523935;
  assign add_524629 = array_index_515098[11:0] + 12'h6ab;
  assign sel_524631 = $signed({1'h0, add_523945}) < $signed({1'h0, sel_523947}) ? add_523945 : sel_523947;
  assign add_524633 = array_index_515101[11:0] + 12'h6ab;
  assign sel_524635 = $signed({1'h0, add_523949}) < $signed({1'h0, sel_523951}) ? add_523949 : sel_523951;
  assign add_524645 = array_index_515726[11:0] + 12'h7d5;
  assign sel_524647 = $signed({1'h0, add_523961}) < $signed({1'h0, sel_523963}) ? add_523961 : sel_523963;
  assign add_524649 = array_index_515729[11:0] + 12'h7d5;
  assign sel_524651 = $signed({1'h0, add_523965}) < $signed({1'h0, sel_523967}) ? add_523965 : sel_523967;
  assign add_524707 = concat_524500 + 4'h1;
  assign add_524709 = array_index_512818[11:1] + 11'h663;
  assign add_524711 = array_index_512819[11:1] + 11'h663;
  assign add_524723 = array_index_512880[11:1] + 11'h075;
  assign sel_524725 = $signed({1'h0, add_524035, array_index_512834[0]}) < $signed({1'h0, sel_524037}) ? {add_524035, array_index_512834[0]} : sel_524037;
  assign add_524727 = array_index_512883[11:1] + 11'h075;
  assign sel_524729 = $signed({1'h0, add_524039, array_index_512837[0]}) < $signed({1'h0, sel_524041}) ? {add_524039, array_index_512837[0]} : sel_524041;
  assign add_524741 = array_index_513022[11:2] + 10'h181;
  assign sel_524743 = $signed({1'h0, add_524053, array_index_512942[1:0]}) < $signed({1'h0, sel_524055}) ? {add_524053, array_index_512942[1:0]} : sel_524055;
  assign add_524745 = array_index_513025[11:2] + 10'h181;
  assign sel_524747 = $signed({1'h0, add_524057, array_index_512945[1:0]}) < $signed({1'h0, sel_524059}) ? {add_524057, array_index_512945[1:0]} : sel_524059;
  assign add_524759 = array_index_513238[11:0] + 12'h8a7;
  assign sel_524761 = $signed({1'h0, add_524071}) < $signed({1'h0, sel_524073}) ? add_524071 : sel_524073;
  assign add_524763 = array_index_513241[11:0] + 12'h8a7;
  assign sel_524765 = $signed({1'h0, add_524075}) < $signed({1'h0, sel_524077}) ? add_524075 : sel_524077;
  assign add_524777 = array_index_513530[11:1] + 11'h283;
  assign sel_524779 = $signed({1'h0, add_524089, array_index_513374[0]}) < $signed({1'h0, sel_524091}) ? {add_524089, array_index_513374[0]} : sel_524091;
  assign add_524781 = array_index_513533[11:1] + 11'h283;
  assign sel_524783 = $signed({1'h0, add_524093, array_index_513377[0]}) < $signed({1'h0, sel_524095}) ? {add_524093, array_index_513377[0]} : sel_524095;
  assign add_524793 = array_index_513890[11:1] + 11'h44d;
  assign sel_524795 = $signed({1'h0, add_524105, array_index_513702[0]}) < $signed({1'h0, sel_524107}) ? {add_524105, array_index_513702[0]} : sel_524107;
  assign add_524797 = array_index_513893[11:1] + 11'h44d;
  assign sel_524799 = $signed({1'h0, add_524109, array_index_513705[0]}) < $signed({1'h0, sel_524111}) ? {add_524109, array_index_513705[0]} : sel_524111;
  assign add_524809 = array_index_514318[11:0] + 12'hcb1;
  assign sel_524811 = $signed({1'h0, add_524121}) < $signed({1'h0, sel_524123}) ? add_524121 : sel_524123;
  assign add_524813 = array_index_514321[11:0] + 12'hcb1;
  assign sel_524815 = $signed({1'h0, add_524125}) < $signed({1'h0, sel_524127}) ? add_524125 : sel_524127;
  assign add_524825 = array_index_514818[11:0] + 12'h81f;
  assign sel_524827 = $signed({1'h0, add_524137}) < $signed({1'h0, sel_524139}) ? add_524137 : sel_524139;
  assign add_524829 = array_index_514821[11:0] + 12'h81f;
  assign sel_524831 = $signed({1'h0, add_524141}) < $signed({1'h0, sel_524143}) ? add_524141 : sel_524143;
  assign add_524841 = array_index_515398[11:0] + 12'h45b;
  assign sel_524843 = $signed({1'h0, add_524153}) < $signed({1'h0, sel_524155}) ? add_524153 : sel_524155;
  assign add_524845 = array_index_515401[11:0] + 12'h45b;
  assign sel_524847 = $signed({1'h0, add_524157}) < $signed({1'h0, sel_524159}) ? add_524157 : sel_524159;
  assign add_524859 = array_index_516080[11:3] + 9'h0f5;
  assign sel_524861 = $signed({1'h0, add_524171, array_index_515726[2:0]}) < $signed({1'h0, sel_524173}) ? {add_524171, array_index_515726[2:0]} : sel_524173;
  assign add_524863 = array_index_516083[11:3] + 9'h0f5;
  assign sel_524865 = $signed({1'h0, add_524175, array_index_515729[2:0]}) < $signed({1'h0, sel_524177}) ? {add_524175, array_index_515729[2:0]} : sel_524177;
  assign add_524939 = array_index_512834[11:0] + 12'h263;
  assign sel_524941 = $signed({1'h0, add_524251}) < $signed(13'h0fff) ? add_524251 : 12'hfff;
  assign add_524943 = array_index_512837[11:0] + 12'h263;
  assign sel_524945 = $signed({1'h0, add_524253}) < $signed(13'h0fff) ? add_524253 : 12'hfff;
  assign add_524955 = array_index_512942[11:1] + 11'h109;
  assign sel_524957 = $signed({1'h0, add_524265, array_index_512880[0]}) < $signed({1'h0, sel_524267}) ? {add_524265, array_index_512880[0]} : sel_524267;
  assign add_524959 = array_index_512945[11:1] + 11'h109;
  assign sel_524961 = $signed({1'h0, add_524269, array_index_512883[0]}) < $signed({1'h0, sel_524271}) ? {add_524269, array_index_512883[0]} : sel_524271;
  assign add_524971 = array_index_513120[11:3] + 9'h12f;
  assign sel_524973 = $signed({1'h0, add_524281, array_index_513022[2:0]}) < $signed({1'h0, sel_524283}) ? {add_524281, array_index_513022[2:0]} : sel_524283;
  assign add_524975 = array_index_513123[11:3] + 9'h12f;
  assign sel_524977 = $signed({1'h0, add_524285, array_index_513025[2:0]}) < $signed({1'h0, sel_524287}) ? {add_524285, array_index_513025[2:0]} : sel_524287;
  assign add_524989 = array_index_513374[11:3] + 9'h171;
  assign sel_524991 = $signed({1'h0, add_524299, array_index_513238[2:0]}) < $signed({1'h0, sel_524301}) ? {add_524299, array_index_513238[2:0]} : sel_524301;
  assign add_524993 = array_index_513377[11:3] + 9'h171;
  assign sel_524995 = $signed({1'h0, add_524303, array_index_513241[2:0]}) < $signed({1'h0, sel_524305}) ? {add_524303, array_index_513241[2:0]} : sel_524305;
  assign add_525005 = array_index_513702[11:0] + 12'h091;
  assign sel_525007 = $signed({1'h0, add_524315}) < $signed({1'h0, sel_524317}) ? add_524315 : sel_524317;
  assign add_525009 = array_index_513705[11:0] + 12'h091;
  assign sel_525011 = $signed({1'h0, add_524319}) < $signed({1'h0, sel_524321}) ? add_524319 : sel_524321;
  assign add_525021 = array_index_514096[11:0] + 12'hf59;
  assign sel_525023 = $signed({1'h0, add_524331}) < $signed({1'h0, sel_524333}) ? add_524331 : sel_524333;
  assign add_525025 = array_index_514099[11:0] + 12'hf59;
  assign sel_525027 = $signed({1'h0, add_524335}) < $signed({1'h0, sel_524337}) ? add_524335 : sel_524337;
  assign add_525039 = array_index_514558[11:0] + 12'h437;
  assign sel_525041 = $signed({1'h0, add_524349}) < $signed({1'h0, sel_524351}) ? add_524349 : sel_524351;
  assign add_525043 = array_index_514561[11:0] + 12'h437;
  assign sel_525045 = $signed({1'h0, add_524353}) < $signed({1'h0, sel_524355}) ? add_524353 : sel_524355;
  assign add_525055 = array_index_515098[11:0] + 12'hee1;
  assign sel_525057 = $signed({1'h0, add_524365}) < $signed({1'h0, sel_524367}) ? add_524365 : sel_524367;
  assign add_525059 = array_index_515101[11:0] + 12'hee1;
  assign sel_525061 = $signed({1'h0, add_524369}) < $signed({1'h0, sel_524371}) ? add_524369 : sel_524371;
  assign add_525071 = array_index_515726[11:1] + 11'h179;
  assign sel_525073 = $signed({1'h0, add_524381, array_index_515398[0]}) < $signed({1'h0, sel_524383}) ? {add_524381, array_index_515398[0]} : sel_524383;
  assign add_525075 = array_index_515729[11:1] + 11'h179;
  assign sel_525077 = $signed({1'h0, add_524385, array_index_515401[0]}) < $signed({1'h0, sel_524387}) ? {add_524385, array_index_515401[0]} : sel_524387;
  assign add_525087 = array_index_516458[11:0] + 12'h067;
  assign sel_525089 = $signed({1'h0, add_524397}) < $signed({1'h0, sel_524399}) ? add_524397 : sel_524399;
  assign add_525091 = array_index_516461[11:0] + 12'h067;
  assign sel_525093 = $signed({1'h0, add_524401}) < $signed({1'h0, sel_524403}) ? add_524401 : sel_524403;
  assign add_525095 = array_index_516860[11:3] + 9'h1ef;
  assign sel_525098 = $signed({1'h0, add_524405, array_index_516458[2:0]}) < $signed({1'h0, sel_524408}) ? {add_524405, array_index_516458[2:0]} : sel_524408;
  assign add_525100 = array_index_516863[11:3] + 9'h1ef;
  assign sel_525103 = $signed({1'h0, add_524410, array_index_516461[2:0]}) < $signed({1'h0, sel_524413}) ? {add_524410, array_index_516461[2:0]} : sel_524413;
  assign add_525105 = array_index_517286[11:1] + 11'h2d5;
  assign sel_525107 = $signed({1'h0, add_524415, array_index_516860[0]}) < $signed({1'h0, sel_524417}) ? {add_524415, array_index_516860[0]} : sel_524417;
  assign add_525109 = array_index_517289[11:1] + 11'h2d5;
  assign sel_525111 = $signed({1'h0, add_524419, array_index_516863[0]}) < $signed({1'h0, sel_524421}) ? {add_524419, array_index_516863[0]} : sel_524421;
  assign add_525113 = array_index_517736[11:2] + 10'h353;
  assign sel_525115 = $signed({1'h0, add_524423, array_index_517286[1:0]}) < $signed({1'h0, sel_524425}) ? {add_524423, array_index_517286[1:0]} : sel_524425;
  assign add_525117 = array_index_517739[11:2] + 10'h353;
  assign sel_525119 = $signed({1'h0, add_524427, array_index_517289[1:0]}) < $signed({1'h0, sel_524429}) ? {add_524427, array_index_517289[1:0]} : sel_524429;
  assign add_525121 = array_index_518210[11:0] + 12'h0a7;
  assign sel_525123 = $signed({1'h0, add_524431}) < $signed({1'h0, sel_524433}) ? add_524431 : sel_524433;
  assign add_525125 = array_index_518213[11:0] + 12'h0a7;
  assign sel_525127 = $signed({1'h0, add_524435}) < $signed({1'h0, sel_524437}) ? add_524435 : sel_524437;
  assign add_525129 = array_index_518710[11:1] + 11'h4cb;
  assign sel_525131 = $signed({1'h0, add_524439, array_index_518210[0]}) < $signed({1'h0, sel_524441}) ? {add_524439, array_index_518210[0]} : sel_524441;
  assign add_525133 = array_index_518713[11:1] + 11'h4cb;
  assign sel_525135 = $signed({1'h0, add_524443, array_index_518213[0]}) < $signed({1'h0, sel_524445}) ? {add_524443, array_index_518213[0]} : sel_524445;
  assign add_525137 = array_index_519236[11:0] + 12'hfe9;
  assign sel_525139 = $signed({1'h0, add_524447}) < $signed({1'h0, sel_524449}) ? add_524447 : sel_524449;
  assign add_525141 = array_index_519239[11:0] + 12'hfe9;
  assign sel_525143 = $signed({1'h0, add_524451}) < $signed({1'h0, sel_524453}) ? add_524451 : sel_524453;
  assign add_525145 = array_index_519786[11:0] + 12'h97d;
  assign sel_525147 = $signed({1'h0, add_524455}) < $signed({1'h0, sel_524457}) ? add_524455 : sel_524457;
  assign add_525149 = array_index_519789[11:0] + 12'h97d;
  assign sel_525151 = $signed({1'h0, add_524459}) < $signed({1'h0, sel_524461}) ? add_524459 : sel_524461;
  assign add_525153 = array_index_520362[11:2] + 10'h2bb;
  assign sel_525156 = $signed({1'h0, add_524463, array_index_519786[1:0]}) < $signed({1'h0, sel_524466}) ? {add_524463, array_index_519786[1:0]} : sel_524466;
  assign add_525158 = array_index_520365[11:2] + 10'h2bb;
  assign sel_525161 = $signed({1'h0, add_524468, array_index_519789[1:0]}) < $signed({1'h0, sel_524471}) ? {add_524468, array_index_519789[1:0]} : sel_524471;
  assign add_525163 = array_index_520964[11:0] + 12'h8e1;
  assign sel_525165 = $signed({1'h0, add_524473}) < $signed({1'h0, sel_524475}) ? add_524473 : sel_524475;
  assign add_525167 = array_index_520967[11:0] + 12'h8e1;
  assign sel_525169 = $signed({1'h0, add_524477}) < $signed({1'h0, sel_524479}) ? add_524477 : sel_524479;
  assign add_525171 = array_index_521590[11:4] + 8'h83;
  assign sel_525174 = $signed({1'h0, add_524481, array_index_520964[3:0]}) < $signed({1'h0, sel_524484}) ? {add_524481, array_index_520964[3:0]} : sel_524484;
  assign add_525176 = array_index_521593[11:4] + 8'h83;
  assign sel_525179 = $signed({1'h0, add_524486, array_index_520967[3:0]}) < $signed({1'h0, sel_524489}) ? {add_524486, array_index_520967[3:0]} : sel_524489;
  assign concat_525182 = {1'h0, ($signed({1'h0, add_523815, array_index_521590[0]}) < $signed({1'h0, sel_523817}) ? {add_523815, array_index_521590[0]} : sel_523817) == ($signed({1'h0, add_523819, array_index_521593[0]}) < $signed({1'h0, sel_523821}) ? {add_523819, array_index_521593[0]} : sel_523821) ? add_524707 : concat_524500};
  assign add_525185 = array_index_512818[11:0] + 12'h37b;
  assign add_525187 = array_index_512819[11:0] + 12'h37b;
  assign add_525201 = array_index_512880[11:0] + 12'h811;
  assign sel_525203 = $signed({1'h0, add_524509}) < $signed({1'h0, sel_524511}) ? add_524509 : sel_524511;
  assign add_525205 = array_index_512883[11:0] + 12'h811;
  assign sel_525207 = $signed({1'h0, add_524513}) < $signed({1'h0, sel_524515}) ? add_524513 : sel_524515;
  assign add_525219 = array_index_513022[11:0] + 12'h70f;
  assign sel_525221 = $signed({1'h0, add_524527}) < $signed({1'h0, sel_524529}) ? add_524527 : sel_524529;
  assign add_525223 = array_index_513025[11:0] + 12'h70f;
  assign sel_525225 = $signed({1'h0, add_524531}) < $signed({1'h0, sel_524533}) ? add_524531 : sel_524533;
  assign add_525237 = array_index_513238[11:3] + 9'h1f1;
  assign sel_525239 = $signed({1'h0, add_524545, array_index_513120[2:0]}) < $signed({1'h0, sel_524547}) ? {add_524545, array_index_513120[2:0]} : sel_524547;
  assign add_525241 = array_index_513241[11:3] + 9'h1f1;
  assign sel_525243 = $signed({1'h0, add_524549, array_index_513123[2:0]}) < $signed({1'h0, sel_524551}) ? {add_524549, array_index_513123[2:0]} : sel_524551;
  assign add_525253 = array_index_513530[11:0] + 12'h081;
  assign sel_525255 = $signed({1'h0, add_524561}) < $signed({1'h0, sel_524563}) ? add_524561 : sel_524563;
  assign add_525257 = array_index_513533[11:0] + 12'h081;
  assign sel_525259 = $signed({1'h0, add_524565}) < $signed({1'h0, sel_524567}) ? add_524565 : sel_524567;
  assign add_525271 = array_index_513890[11:0] + 12'h0b1;
  assign sel_525273 = $signed({1'h0, add_524579}) < $signed({1'h0, sel_524581}) ? add_524579 : sel_524581;
  assign add_525275 = array_index_513893[11:0] + 12'h0b1;
  assign sel_525277 = $signed({1'h0, add_524583}) < $signed({1'h0, sel_524585}) ? add_524583 : sel_524585;
  assign add_525289 = array_index_514318[11:1] + 11'h4c1;
  assign sel_525291 = $signed({1'h0, add_524597, array_index_514096[0]}) < $signed({1'h0, sel_524599}) ? {add_524597, array_index_514096[0]} : sel_524599;
  assign add_525293 = array_index_514321[11:1] + 11'h4c1;
  assign sel_525295 = $signed({1'h0, add_524601, array_index_514099[0]}) < $signed({1'h0, sel_524603}) ? {add_524601, array_index_514099[0]} : sel_524603;
  assign add_525305 = array_index_514818[11:0] + 12'hbb1;
  assign sel_525307 = $signed({1'h0, add_524613}) < $signed({1'h0, sel_524615}) ? add_524613 : sel_524615;
  assign add_525309 = array_index_514821[11:0] + 12'hbb1;
  assign sel_525311 = $signed({1'h0, add_524617}) < $signed({1'h0, sel_524619}) ? add_524617 : sel_524619;
  assign add_525321 = array_index_515398[11:0] + 12'h6ab;
  assign sel_525323 = $signed({1'h0, add_524629}) < $signed({1'h0, sel_524631}) ? add_524629 : sel_524631;
  assign add_525325 = array_index_515401[11:0] + 12'h6ab;
  assign sel_525327 = $signed({1'h0, add_524633}) < $signed({1'h0, sel_524635}) ? add_524633 : sel_524635;
  assign add_525337 = array_index_516080[11:0] + 12'h7d5;
  assign sel_525339 = $signed({1'h0, add_524645}) < $signed({1'h0, sel_524647}) ? add_524645 : sel_524647;
  assign add_525341 = array_index_516083[11:0] + 12'h7d5;
  assign sel_525343 = $signed({1'h0, add_524649}) < $signed({1'h0, sel_524651}) ? add_524649 : sel_524651;
  assign add_525395 = concat_525182 + 5'h01;
  assign add_525403 = array_index_512834[11:1] + 11'h663;
  assign sel_525405 = $signed({1'h0, add_524709, array_index_512818[0]}) < $signed(13'h0fff) ? {add_524709, array_index_512818[0]} : 12'hfff;
  assign add_525407 = array_index_512837[11:1] + 11'h663;
  assign sel_525409 = $signed({1'h0, add_524711, array_index_512819[0]}) < $signed(13'h0fff) ? {add_524711, array_index_512819[0]} : 12'hfff;
  assign add_525419 = array_index_512942[11:1] + 11'h075;
  assign sel_525421 = $signed({1'h0, add_524723, array_index_512880[0]}) < $signed({1'h0, sel_524725}) ? {add_524723, array_index_512880[0]} : sel_524725;
  assign add_525423 = array_index_512945[11:1] + 11'h075;
  assign sel_525425 = $signed({1'h0, add_524727, array_index_512883[0]}) < $signed({1'h0, sel_524729}) ? {add_524727, array_index_512883[0]} : sel_524729;
  assign add_525437 = array_index_513120[11:2] + 10'h181;
  assign sel_525439 = $signed({1'h0, add_524741, array_index_513022[1:0]}) < $signed({1'h0, sel_524743}) ? {add_524741, array_index_513022[1:0]} : sel_524743;
  assign add_525441 = array_index_513123[11:2] + 10'h181;
  assign sel_525443 = $signed({1'h0, add_524745, array_index_513025[1:0]}) < $signed({1'h0, sel_524747}) ? {add_524745, array_index_513025[1:0]} : sel_524747;
  assign add_525455 = array_index_513374[11:0] + 12'h8a7;
  assign sel_525457 = $signed({1'h0, add_524759}) < $signed({1'h0, sel_524761}) ? add_524759 : sel_524761;
  assign add_525459 = array_index_513377[11:0] + 12'h8a7;
  assign sel_525461 = $signed({1'h0, add_524763}) < $signed({1'h0, sel_524765}) ? add_524763 : sel_524765;
  assign add_525473 = array_index_513702[11:1] + 11'h283;
  assign sel_525475 = $signed({1'h0, add_524777, array_index_513530[0]}) < $signed({1'h0, sel_524779}) ? {add_524777, array_index_513530[0]} : sel_524779;
  assign add_525477 = array_index_513705[11:1] + 11'h283;
  assign sel_525479 = $signed({1'h0, add_524781, array_index_513533[0]}) < $signed({1'h0, sel_524783}) ? {add_524781, array_index_513533[0]} : sel_524783;
  assign add_525489 = array_index_514096[11:1] + 11'h44d;
  assign sel_525491 = $signed({1'h0, add_524793, array_index_513890[0]}) < $signed({1'h0, sel_524795}) ? {add_524793, array_index_513890[0]} : sel_524795;
  assign add_525493 = array_index_514099[11:1] + 11'h44d;
  assign sel_525495 = $signed({1'h0, add_524797, array_index_513893[0]}) < $signed({1'h0, sel_524799}) ? {add_524797, array_index_513893[0]} : sel_524799;
  assign add_525505 = array_index_514558[11:0] + 12'hcb1;
  assign sel_525507 = $signed({1'h0, add_524809}) < $signed({1'h0, sel_524811}) ? add_524809 : sel_524811;
  assign add_525509 = array_index_514561[11:0] + 12'hcb1;
  assign sel_525511 = $signed({1'h0, add_524813}) < $signed({1'h0, sel_524815}) ? add_524813 : sel_524815;
  assign add_525521 = array_index_515098[11:0] + 12'h81f;
  assign sel_525523 = $signed({1'h0, add_524825}) < $signed({1'h0, sel_524827}) ? add_524825 : sel_524827;
  assign add_525525 = array_index_515101[11:0] + 12'h81f;
  assign sel_525527 = $signed({1'h0, add_524829}) < $signed({1'h0, sel_524831}) ? add_524829 : sel_524831;
  assign add_525537 = array_index_515726[11:0] + 12'h45b;
  assign sel_525539 = $signed({1'h0, add_524841}) < $signed({1'h0, sel_524843}) ? add_524841 : sel_524843;
  assign add_525541 = array_index_515729[11:0] + 12'h45b;
  assign sel_525543 = $signed({1'h0, add_524845}) < $signed({1'h0, sel_524847}) ? add_524845 : sel_524847;
  assign add_525555 = array_index_516458[11:3] + 9'h0f5;
  assign sel_525557 = $signed({1'h0, add_524859, array_index_516080[2:0]}) < $signed({1'h0, sel_524861}) ? {add_524859, array_index_516080[2:0]} : sel_524861;
  assign add_525559 = array_index_516461[11:3] + 9'h0f5;
  assign sel_525561 = $signed({1'h0, add_524863, array_index_516083[2:0]}) < $signed({1'h0, sel_524865}) ? {add_524863, array_index_516083[2:0]} : sel_524865;
  assign add_525623 = array_index_512818[11:4] + 8'h49;
  assign add_525625 = array_index_512819[11:4] + 8'h49;
  assign add_525637 = array_index_512880[11:0] + 12'h263;
  assign sel_525639 = $signed({1'h0, add_524939}) < $signed({1'h0, sel_524941}) ? add_524939 : sel_524941;
  assign add_525641 = array_index_512883[11:0] + 12'h263;
  assign sel_525643 = $signed({1'h0, add_524943}) < $signed({1'h0, sel_524945}) ? add_524943 : sel_524945;
  assign add_525653 = array_index_513022[11:1] + 11'h109;
  assign sel_525655 = $signed({1'h0, add_524955, array_index_512942[0]}) < $signed({1'h0, sel_524957}) ? {add_524955, array_index_512942[0]} : sel_524957;
  assign add_525657 = array_index_513025[11:1] + 11'h109;
  assign sel_525659 = $signed({1'h0, add_524959, array_index_512945[0]}) < $signed({1'h0, sel_524961}) ? {add_524959, array_index_512945[0]} : sel_524961;
  assign add_525669 = array_index_513238[11:3] + 9'h12f;
  assign sel_525671 = $signed({1'h0, add_524971, array_index_513120[2:0]}) < $signed({1'h0, sel_524973}) ? {add_524971, array_index_513120[2:0]} : sel_524973;
  assign add_525673 = array_index_513241[11:3] + 9'h12f;
  assign sel_525675 = $signed({1'h0, add_524975, array_index_513123[2:0]}) < $signed({1'h0, sel_524977}) ? {add_524975, array_index_513123[2:0]} : sel_524977;
  assign add_525687 = array_index_513530[11:3] + 9'h171;
  assign sel_525689 = $signed({1'h0, add_524989, array_index_513374[2:0]}) < $signed({1'h0, sel_524991}) ? {add_524989, array_index_513374[2:0]} : sel_524991;
  assign add_525691 = array_index_513533[11:3] + 9'h171;
  assign sel_525693 = $signed({1'h0, add_524993, array_index_513377[2:0]}) < $signed({1'h0, sel_524995}) ? {add_524993, array_index_513377[2:0]} : sel_524995;
  assign add_525703 = array_index_513890[11:0] + 12'h091;
  assign sel_525705 = $signed({1'h0, add_525005}) < $signed({1'h0, sel_525007}) ? add_525005 : sel_525007;
  assign add_525707 = array_index_513893[11:0] + 12'h091;
  assign sel_525709 = $signed({1'h0, add_525009}) < $signed({1'h0, sel_525011}) ? add_525009 : sel_525011;
  assign add_525719 = array_index_514318[11:0] + 12'hf59;
  assign sel_525721 = $signed({1'h0, add_525021}) < $signed({1'h0, sel_525023}) ? add_525021 : sel_525023;
  assign add_525723 = array_index_514321[11:0] + 12'hf59;
  assign sel_525725 = $signed({1'h0, add_525025}) < $signed({1'h0, sel_525027}) ? add_525025 : sel_525027;
  assign add_525737 = array_index_514818[11:0] + 12'h437;
  assign sel_525739 = $signed({1'h0, add_525039}) < $signed({1'h0, sel_525041}) ? add_525039 : sel_525041;
  assign add_525741 = array_index_514821[11:0] + 12'h437;
  assign sel_525743 = $signed({1'h0, add_525043}) < $signed({1'h0, sel_525045}) ? add_525043 : sel_525045;
  assign add_525753 = array_index_515398[11:0] + 12'hee1;
  assign sel_525755 = $signed({1'h0, add_525055}) < $signed({1'h0, sel_525057}) ? add_525055 : sel_525057;
  assign add_525757 = array_index_515401[11:0] + 12'hee1;
  assign sel_525759 = $signed({1'h0, add_525059}) < $signed({1'h0, sel_525061}) ? add_525059 : sel_525061;
  assign add_525769 = array_index_516080[11:1] + 11'h179;
  assign sel_525771 = $signed({1'h0, add_525071, array_index_515726[0]}) < $signed({1'h0, sel_525073}) ? {add_525071, array_index_515726[0]} : sel_525073;
  assign add_525773 = array_index_516083[11:1] + 11'h179;
  assign sel_525775 = $signed({1'h0, add_525075, array_index_515729[0]}) < $signed({1'h0, sel_525077}) ? {add_525075, array_index_515729[0]} : sel_525077;
  assign add_525785 = array_index_516860[11:0] + 12'h067;
  assign sel_525787 = $signed({1'h0, add_525087}) < $signed({1'h0, sel_525089}) ? add_525087 : sel_525089;
  assign add_525789 = array_index_516863[11:0] + 12'h067;
  assign sel_525791 = $signed({1'h0, add_525091}) < $signed({1'h0, sel_525093}) ? add_525091 : sel_525093;
  assign add_525793 = array_index_517286[11:3] + 9'h1ef;
  assign sel_525796 = $signed({1'h0, add_525095, array_index_516860[2:0]}) < $signed({1'h0, sel_525098}) ? {add_525095, array_index_516860[2:0]} : sel_525098;
  assign add_525798 = array_index_517289[11:3] + 9'h1ef;
  assign sel_525801 = $signed({1'h0, add_525100, array_index_516863[2:0]}) < $signed({1'h0, sel_525103}) ? {add_525100, array_index_516863[2:0]} : sel_525103;
  assign add_525803 = array_index_517736[11:1] + 11'h2d5;
  assign sel_525805 = $signed({1'h0, add_525105, array_index_517286[0]}) < $signed({1'h0, sel_525107}) ? {add_525105, array_index_517286[0]} : sel_525107;
  assign add_525807 = array_index_517739[11:1] + 11'h2d5;
  assign sel_525809 = $signed({1'h0, add_525109, array_index_517289[0]}) < $signed({1'h0, sel_525111}) ? {add_525109, array_index_517289[0]} : sel_525111;
  assign add_525811 = array_index_518210[11:2] + 10'h353;
  assign sel_525813 = $signed({1'h0, add_525113, array_index_517736[1:0]}) < $signed({1'h0, sel_525115}) ? {add_525113, array_index_517736[1:0]} : sel_525115;
  assign add_525815 = array_index_518213[11:2] + 10'h353;
  assign sel_525817 = $signed({1'h0, add_525117, array_index_517739[1:0]}) < $signed({1'h0, sel_525119}) ? {add_525117, array_index_517739[1:0]} : sel_525119;
  assign add_525819 = array_index_518710[11:0] + 12'h0a7;
  assign sel_525821 = $signed({1'h0, add_525121}) < $signed({1'h0, sel_525123}) ? add_525121 : sel_525123;
  assign add_525823 = array_index_518713[11:0] + 12'h0a7;
  assign sel_525825 = $signed({1'h0, add_525125}) < $signed({1'h0, sel_525127}) ? add_525125 : sel_525127;
  assign add_525827 = array_index_519236[11:1] + 11'h4cb;
  assign sel_525829 = $signed({1'h0, add_525129, array_index_518710[0]}) < $signed({1'h0, sel_525131}) ? {add_525129, array_index_518710[0]} : sel_525131;
  assign add_525831 = array_index_519239[11:1] + 11'h4cb;
  assign sel_525833 = $signed({1'h0, add_525133, array_index_518713[0]}) < $signed({1'h0, sel_525135}) ? {add_525133, array_index_518713[0]} : sel_525135;
  assign add_525835 = array_index_519786[11:0] + 12'hfe9;
  assign sel_525837 = $signed({1'h0, add_525137}) < $signed({1'h0, sel_525139}) ? add_525137 : sel_525139;
  assign add_525839 = array_index_519789[11:0] + 12'hfe9;
  assign sel_525841 = $signed({1'h0, add_525141}) < $signed({1'h0, sel_525143}) ? add_525141 : sel_525143;
  assign add_525843 = array_index_520362[11:0] + 12'h97d;
  assign sel_525845 = $signed({1'h0, add_525145}) < $signed({1'h0, sel_525147}) ? add_525145 : sel_525147;
  assign add_525847 = array_index_520365[11:0] + 12'h97d;
  assign sel_525849 = $signed({1'h0, add_525149}) < $signed({1'h0, sel_525151}) ? add_525149 : sel_525151;
  assign add_525851 = array_index_520964[11:2] + 10'h2bb;
  assign sel_525854 = $signed({1'h0, add_525153, array_index_520362[1:0]}) < $signed({1'h0, sel_525156}) ? {add_525153, array_index_520362[1:0]} : sel_525156;
  assign add_525856 = array_index_520967[11:2] + 10'h2bb;
  assign sel_525859 = $signed({1'h0, add_525158, array_index_520365[1:0]}) < $signed({1'h0, sel_525161}) ? {add_525158, array_index_520365[1:0]} : sel_525161;
  assign add_525861 = array_index_521590[11:0] + 12'h8e1;
  assign sel_525863 = $signed({1'h0, add_525163}) < $signed({1'h0, sel_525165}) ? add_525163 : sel_525165;
  assign add_525865 = array_index_521593[11:0] + 12'h8e1;
  assign sel_525867 = $signed({1'h0, add_525167}) < $signed({1'h0, sel_525169}) ? add_525167 : sel_525169;
  assign concat_525870 = {1'h0, ($signed({1'h0, add_524491}) < $signed({1'h0, sel_524493}) ? add_524491 : sel_524493) == ($signed({1'h0, add_524495}) < $signed({1'h0, sel_524497}) ? add_524495 : sel_524497) ? add_525395 : concat_525182};
  assign add_525879 = array_index_512834[11:0] + 12'h37b;
  assign sel_525881 = $signed({1'h0, add_525185}) < $signed(13'h0fff) ? add_525185 : 12'hfff;
  assign add_525883 = array_index_512837[11:0] + 12'h37b;
  assign sel_525885 = $signed({1'h0, add_525187}) < $signed(13'h0fff) ? add_525187 : 12'hfff;
  assign add_525897 = array_index_512942[11:0] + 12'h811;
  assign sel_525899 = $signed({1'h0, add_525201}) < $signed({1'h0, sel_525203}) ? add_525201 : sel_525203;
  assign add_525901 = array_index_512945[11:0] + 12'h811;
  assign sel_525903 = $signed({1'h0, add_525205}) < $signed({1'h0, sel_525207}) ? add_525205 : sel_525207;
  assign add_525915 = array_index_513120[11:0] + 12'h70f;
  assign sel_525917 = $signed({1'h0, add_525219}) < $signed({1'h0, sel_525221}) ? add_525219 : sel_525221;
  assign add_525919 = array_index_513123[11:0] + 12'h70f;
  assign sel_525921 = $signed({1'h0, add_525223}) < $signed({1'h0, sel_525225}) ? add_525223 : sel_525225;
  assign add_525933 = array_index_513374[11:3] + 9'h1f1;
  assign sel_525935 = $signed({1'h0, add_525237, array_index_513238[2:0]}) < $signed({1'h0, sel_525239}) ? {add_525237, array_index_513238[2:0]} : sel_525239;
  assign add_525937 = array_index_513377[11:3] + 9'h1f1;
  assign sel_525939 = $signed({1'h0, add_525241, array_index_513241[2:0]}) < $signed({1'h0, sel_525243}) ? {add_525241, array_index_513241[2:0]} : sel_525243;
  assign add_525949 = array_index_513702[11:0] + 12'h081;
  assign sel_525951 = $signed({1'h0, add_525253}) < $signed({1'h0, sel_525255}) ? add_525253 : sel_525255;
  assign add_525953 = array_index_513705[11:0] + 12'h081;
  assign sel_525955 = $signed({1'h0, add_525257}) < $signed({1'h0, sel_525259}) ? add_525257 : sel_525259;
  assign add_525967 = array_index_514096[11:0] + 12'h0b1;
  assign sel_525969 = $signed({1'h0, add_525271}) < $signed({1'h0, sel_525273}) ? add_525271 : sel_525273;
  assign add_525971 = array_index_514099[11:0] + 12'h0b1;
  assign sel_525973 = $signed({1'h0, add_525275}) < $signed({1'h0, sel_525277}) ? add_525275 : sel_525277;
  assign add_525985 = array_index_514558[11:1] + 11'h4c1;
  assign sel_525987 = $signed({1'h0, add_525289, array_index_514318[0]}) < $signed({1'h0, sel_525291}) ? {add_525289, array_index_514318[0]} : sel_525291;
  assign add_525989 = array_index_514561[11:1] + 11'h4c1;
  assign sel_525991 = $signed({1'h0, add_525293, array_index_514321[0]}) < $signed({1'h0, sel_525295}) ? {add_525293, array_index_514321[0]} : sel_525295;
  assign add_526001 = array_index_515098[11:0] + 12'hbb1;
  assign sel_526003 = $signed({1'h0, add_525305}) < $signed({1'h0, sel_525307}) ? add_525305 : sel_525307;
  assign add_526005 = array_index_515101[11:0] + 12'hbb1;
  assign sel_526007 = $signed({1'h0, add_525309}) < $signed({1'h0, sel_525311}) ? add_525309 : sel_525311;
  assign add_526017 = array_index_515726[11:0] + 12'h6ab;
  assign sel_526019 = $signed({1'h0, add_525321}) < $signed({1'h0, sel_525323}) ? add_525321 : sel_525323;
  assign add_526021 = array_index_515729[11:0] + 12'h6ab;
  assign sel_526023 = $signed({1'h0, add_525325}) < $signed({1'h0, sel_525327}) ? add_525325 : sel_525327;
  assign add_526033 = array_index_516458[11:0] + 12'h7d5;
  assign sel_526035 = $signed({1'h0, add_525337}) < $signed({1'h0, sel_525339}) ? add_525337 : sel_525339;
  assign add_526037 = array_index_516461[11:0] + 12'h7d5;
  assign sel_526039 = $signed({1'h0, add_525341}) < $signed({1'h0, sel_525343}) ? add_525341 : sel_525343;
  assign add_526087 = concat_525870 + 6'h01;
  assign add_526089 = array_index_512818[11:0] + 12'ha87;
  assign add_526091 = array_index_512819[11:0] + 12'ha87;
  assign add_526105 = array_index_512880[11:1] + 11'h663;
  assign sel_526107 = $signed({1'h0, add_525403, array_index_512834[0]}) < $signed({1'h0, sel_525405}) ? {add_525403, array_index_512834[0]} : sel_525405;
  assign add_526109 = array_index_512883[11:1] + 11'h663;
  assign sel_526111 = $signed({1'h0, add_525407, array_index_512837[0]}) < $signed({1'h0, sel_525409}) ? {add_525407, array_index_512837[0]} : sel_525409;
  assign add_526121 = array_index_513022[11:1] + 11'h075;
  assign sel_526123 = $signed({1'h0, add_525419, array_index_512942[0]}) < $signed({1'h0, sel_525421}) ? {add_525419, array_index_512942[0]} : sel_525421;
  assign add_526125 = array_index_513025[11:1] + 11'h075;
  assign sel_526127 = $signed({1'h0, add_525423, array_index_512945[0]}) < $signed({1'h0, sel_525425}) ? {add_525423, array_index_512945[0]} : sel_525425;
  assign add_526139 = array_index_513238[11:2] + 10'h181;
  assign sel_526141 = $signed({1'h0, add_525437, array_index_513120[1:0]}) < $signed({1'h0, sel_525439}) ? {add_525437, array_index_513120[1:0]} : sel_525439;
  assign add_526143 = array_index_513241[11:2] + 10'h181;
  assign sel_526145 = $signed({1'h0, add_525441, array_index_513123[1:0]}) < $signed({1'h0, sel_525443}) ? {add_525441, array_index_513123[1:0]} : sel_525443;
  assign add_526157 = array_index_513530[11:0] + 12'h8a7;
  assign sel_526159 = $signed({1'h0, add_525455}) < $signed({1'h0, sel_525457}) ? add_525455 : sel_525457;
  assign add_526161 = array_index_513533[11:0] + 12'h8a7;
  assign sel_526163 = $signed({1'h0, add_525459}) < $signed({1'h0, sel_525461}) ? add_525459 : sel_525461;
  assign add_526175 = array_index_513890[11:1] + 11'h283;
  assign sel_526177 = $signed({1'h0, add_525473, array_index_513702[0]}) < $signed({1'h0, sel_525475}) ? {add_525473, array_index_513702[0]} : sel_525475;
  assign add_526179 = array_index_513893[11:1] + 11'h283;
  assign sel_526181 = $signed({1'h0, add_525477, array_index_513705[0]}) < $signed({1'h0, sel_525479}) ? {add_525477, array_index_513705[0]} : sel_525479;
  assign add_526191 = array_index_514318[11:1] + 11'h44d;
  assign sel_526193 = $signed({1'h0, add_525489, array_index_514096[0]}) < $signed({1'h0, sel_525491}) ? {add_525489, array_index_514096[0]} : sel_525491;
  assign add_526195 = array_index_514321[11:1] + 11'h44d;
  assign sel_526197 = $signed({1'h0, add_525493, array_index_514099[0]}) < $signed({1'h0, sel_525495}) ? {add_525493, array_index_514099[0]} : sel_525495;
  assign add_526207 = array_index_514818[11:0] + 12'hcb1;
  assign sel_526209 = $signed({1'h0, add_525505}) < $signed({1'h0, sel_525507}) ? add_525505 : sel_525507;
  assign add_526211 = array_index_514821[11:0] + 12'hcb1;
  assign sel_526213 = $signed({1'h0, add_525509}) < $signed({1'h0, sel_525511}) ? add_525509 : sel_525511;
  assign add_526223 = array_index_515398[11:0] + 12'h81f;
  assign sel_526225 = $signed({1'h0, add_525521}) < $signed({1'h0, sel_525523}) ? add_525521 : sel_525523;
  assign add_526227 = array_index_515401[11:0] + 12'h81f;
  assign sel_526229 = $signed({1'h0, add_525525}) < $signed({1'h0, sel_525527}) ? add_525525 : sel_525527;
  assign add_526239 = array_index_516080[11:0] + 12'h45b;
  assign sel_526241 = $signed({1'h0, add_525537}) < $signed({1'h0, sel_525539}) ? add_525537 : sel_525539;
  assign add_526243 = array_index_516083[11:0] + 12'h45b;
  assign sel_526245 = $signed({1'h0, add_525541}) < $signed({1'h0, sel_525543}) ? add_525541 : sel_525543;
  assign add_526257 = array_index_516860[11:3] + 9'h0f5;
  assign sel_526259 = $signed({1'h0, add_525555, array_index_516458[2:0]}) < $signed({1'h0, sel_525557}) ? {add_525555, array_index_516458[2:0]} : sel_525557;
  assign add_526261 = array_index_516863[11:3] + 9'h0f5;
  assign sel_526263 = $signed({1'h0, add_525559, array_index_516461[2:0]}) < $signed({1'h0, sel_525561}) ? {add_525559, array_index_516461[2:0]} : sel_525561;
  assign add_526325 = array_index_512834[11:4] + 8'h49;
  assign sel_526327 = $signed({1'h0, add_525623, array_index_512818[3:0]}) < $signed(13'h0fff) ? {add_525623, array_index_512818[3:0]} : 12'hfff;
  assign add_526329 = array_index_512837[11:4] + 8'h49;
  assign sel_526331 = $signed({1'h0, add_525625, array_index_512819[3:0]}) < $signed(13'h0fff) ? {add_525625, array_index_512819[3:0]} : 12'hfff;
  assign add_526341 = array_index_512942[11:0] + 12'h263;
  assign sel_526343 = $signed({1'h0, add_525637}) < $signed({1'h0, sel_525639}) ? add_525637 : sel_525639;
  assign add_526345 = array_index_512945[11:0] + 12'h263;
  assign sel_526347 = $signed({1'h0, add_525641}) < $signed({1'h0, sel_525643}) ? add_525641 : sel_525643;
  assign add_526357 = array_index_513120[11:1] + 11'h109;
  assign sel_526359 = $signed({1'h0, add_525653, array_index_513022[0]}) < $signed({1'h0, sel_525655}) ? {add_525653, array_index_513022[0]} : sel_525655;
  assign add_526361 = array_index_513123[11:1] + 11'h109;
  assign sel_526363 = $signed({1'h0, add_525657, array_index_513025[0]}) < $signed({1'h0, sel_525659}) ? {add_525657, array_index_513025[0]} : sel_525659;
  assign add_526373 = array_index_513374[11:3] + 9'h12f;
  assign sel_526375 = $signed({1'h0, add_525669, array_index_513238[2:0]}) < $signed({1'h0, sel_525671}) ? {add_525669, array_index_513238[2:0]} : sel_525671;
  assign add_526377 = array_index_513377[11:3] + 9'h12f;
  assign sel_526379 = $signed({1'h0, add_525673, array_index_513241[2:0]}) < $signed({1'h0, sel_525675}) ? {add_525673, array_index_513241[2:0]} : sel_525675;
  assign add_526391 = array_index_513702[11:3] + 9'h171;
  assign sel_526393 = $signed({1'h0, add_525687, array_index_513530[2:0]}) < $signed({1'h0, sel_525689}) ? {add_525687, array_index_513530[2:0]} : sel_525689;
  assign add_526395 = array_index_513705[11:3] + 9'h171;
  assign sel_526397 = $signed({1'h0, add_525691, array_index_513533[2:0]}) < $signed({1'h0, sel_525693}) ? {add_525691, array_index_513533[2:0]} : sel_525693;
  assign add_526407 = array_index_514096[11:0] + 12'h091;
  assign sel_526409 = $signed({1'h0, add_525703}) < $signed({1'h0, sel_525705}) ? add_525703 : sel_525705;
  assign add_526411 = array_index_514099[11:0] + 12'h091;
  assign sel_526413 = $signed({1'h0, add_525707}) < $signed({1'h0, sel_525709}) ? add_525707 : sel_525709;
  assign add_526423 = array_index_514558[11:0] + 12'hf59;
  assign sel_526425 = $signed({1'h0, add_525719}) < $signed({1'h0, sel_525721}) ? add_525719 : sel_525721;
  assign add_526427 = array_index_514561[11:0] + 12'hf59;
  assign sel_526429 = $signed({1'h0, add_525723}) < $signed({1'h0, sel_525725}) ? add_525723 : sel_525725;
  assign add_526441 = array_index_515098[11:0] + 12'h437;
  assign sel_526443 = $signed({1'h0, add_525737}) < $signed({1'h0, sel_525739}) ? add_525737 : sel_525739;
  assign add_526445 = array_index_515101[11:0] + 12'h437;
  assign sel_526447 = $signed({1'h0, add_525741}) < $signed({1'h0, sel_525743}) ? add_525741 : sel_525743;
  assign add_526457 = array_index_515726[11:0] + 12'hee1;
  assign sel_526459 = $signed({1'h0, add_525753}) < $signed({1'h0, sel_525755}) ? add_525753 : sel_525755;
  assign add_526461 = array_index_515729[11:0] + 12'hee1;
  assign sel_526463 = $signed({1'h0, add_525757}) < $signed({1'h0, sel_525759}) ? add_525757 : sel_525759;
  assign add_526473 = array_index_516458[11:1] + 11'h179;
  assign sel_526475 = $signed({1'h0, add_525769, array_index_516080[0]}) < $signed({1'h0, sel_525771}) ? {add_525769, array_index_516080[0]} : sel_525771;
  assign add_526477 = array_index_516461[11:1] + 11'h179;
  assign sel_526479 = $signed({1'h0, add_525773, array_index_516083[0]}) < $signed({1'h0, sel_525775}) ? {add_525773, array_index_516083[0]} : sel_525775;
  assign add_526489 = array_index_517286[11:0] + 12'h067;
  assign sel_526491 = $signed({1'h0, add_525785}) < $signed({1'h0, sel_525787}) ? add_525785 : sel_525787;
  assign add_526493 = array_index_517289[11:0] + 12'h067;
  assign sel_526495 = $signed({1'h0, add_525789}) < $signed({1'h0, sel_525791}) ? add_525789 : sel_525791;
  assign add_526497 = array_index_517736[11:3] + 9'h1ef;
  assign sel_526500 = $signed({1'h0, add_525793, array_index_517286[2:0]}) < $signed({1'h0, sel_525796}) ? {add_525793, array_index_517286[2:0]} : sel_525796;
  assign add_526502 = array_index_517739[11:3] + 9'h1ef;
  assign sel_526505 = $signed({1'h0, add_525798, array_index_517289[2:0]}) < $signed({1'h0, sel_525801}) ? {add_525798, array_index_517289[2:0]} : sel_525801;
  assign add_526507 = array_index_518210[11:1] + 11'h2d5;
  assign sel_526509 = $signed({1'h0, add_525803, array_index_517736[0]}) < $signed({1'h0, sel_525805}) ? {add_525803, array_index_517736[0]} : sel_525805;
  assign add_526511 = array_index_518213[11:1] + 11'h2d5;
  assign sel_526513 = $signed({1'h0, add_525807, array_index_517739[0]}) < $signed({1'h0, sel_525809}) ? {add_525807, array_index_517739[0]} : sel_525809;
  assign add_526515 = array_index_518710[11:2] + 10'h353;
  assign sel_526517 = $signed({1'h0, add_525811, array_index_518210[1:0]}) < $signed({1'h0, sel_525813}) ? {add_525811, array_index_518210[1:0]} : sel_525813;
  assign add_526519 = array_index_518713[11:2] + 10'h353;
  assign sel_526521 = $signed({1'h0, add_525815, array_index_518213[1:0]}) < $signed({1'h0, sel_525817}) ? {add_525815, array_index_518213[1:0]} : sel_525817;
  assign add_526523 = array_index_519236[11:0] + 12'h0a7;
  assign sel_526525 = $signed({1'h0, add_525819}) < $signed({1'h0, sel_525821}) ? add_525819 : sel_525821;
  assign add_526527 = array_index_519239[11:0] + 12'h0a7;
  assign sel_526529 = $signed({1'h0, add_525823}) < $signed({1'h0, sel_525825}) ? add_525823 : sel_525825;
  assign add_526531 = array_index_519786[11:1] + 11'h4cb;
  assign sel_526533 = $signed({1'h0, add_525827, array_index_519236[0]}) < $signed({1'h0, sel_525829}) ? {add_525827, array_index_519236[0]} : sel_525829;
  assign add_526535 = array_index_519789[11:1] + 11'h4cb;
  assign sel_526537 = $signed({1'h0, add_525831, array_index_519239[0]}) < $signed({1'h0, sel_525833}) ? {add_525831, array_index_519239[0]} : sel_525833;
  assign add_526539 = array_index_520362[11:0] + 12'hfe9;
  assign sel_526541 = $signed({1'h0, add_525835}) < $signed({1'h0, sel_525837}) ? add_525835 : sel_525837;
  assign add_526543 = array_index_520365[11:0] + 12'hfe9;
  assign sel_526545 = $signed({1'h0, add_525839}) < $signed({1'h0, sel_525841}) ? add_525839 : sel_525841;
  assign add_526547 = array_index_520964[11:0] + 12'h97d;
  assign sel_526549 = $signed({1'h0, add_525843}) < $signed({1'h0, sel_525845}) ? add_525843 : sel_525845;
  assign add_526551 = array_index_520967[11:0] + 12'h97d;
  assign sel_526553 = $signed({1'h0, add_525847}) < $signed({1'h0, sel_525849}) ? add_525847 : sel_525849;
  assign add_526555 = array_index_521590[11:2] + 10'h2bb;
  assign sel_526558 = $signed({1'h0, add_525851, array_index_520964[1:0]}) < $signed({1'h0, sel_525854}) ? {add_525851, array_index_520964[1:0]} : sel_525854;
  assign add_526560 = array_index_521593[11:2] + 10'h2bb;
  assign sel_526563 = $signed({1'h0, add_525856, array_index_520967[1:0]}) < $signed({1'h0, sel_525859}) ? {add_525856, array_index_520967[1:0]} : sel_525859;
  assign concat_526566 = {1'h0, ($signed({1'h0, add_525171, array_index_521590[3:0]}) < $signed({1'h0, sel_525174}) ? {add_525171, array_index_521590[3:0]} : sel_525174) == ($signed({1'h0, add_525176, array_index_521593[3:0]}) < $signed({1'h0, sel_525179}) ? {add_525176, array_index_521593[3:0]} : sel_525179) ? add_526087 : concat_525870};
  assign add_526569 = array_index_512818[11:1] + 11'h5b9;
  assign add_526571 = array_index_512819[11:1] + 11'h5b9;
  assign add_526583 = array_index_512880[11:0] + 12'h37b;
  assign sel_526585 = $signed({1'h0, add_525879}) < $signed({1'h0, sel_525881}) ? add_525879 : sel_525881;
  assign add_526587 = array_index_512883[11:0] + 12'h37b;
  assign sel_526589 = $signed({1'h0, add_525883}) < $signed({1'h0, sel_525885}) ? add_525883 : sel_525885;
  assign add_526601 = array_index_513022[11:0] + 12'h811;
  assign sel_526603 = $signed({1'h0, add_525897}) < $signed({1'h0, sel_525899}) ? add_525897 : sel_525899;
  assign add_526605 = array_index_513025[11:0] + 12'h811;
  assign sel_526607 = $signed({1'h0, add_525901}) < $signed({1'h0, sel_525903}) ? add_525901 : sel_525903;
  assign add_526619 = array_index_513238[11:0] + 12'h70f;
  assign sel_526621 = $signed({1'h0, add_525915}) < $signed({1'h0, sel_525917}) ? add_525915 : sel_525917;
  assign add_526623 = array_index_513241[11:0] + 12'h70f;
  assign sel_526625 = $signed({1'h0, add_525919}) < $signed({1'h0, sel_525921}) ? add_525919 : sel_525921;
  assign add_526637 = array_index_513530[11:3] + 9'h1f1;
  assign sel_526639 = $signed({1'h0, add_525933, array_index_513374[2:0]}) < $signed({1'h0, sel_525935}) ? {add_525933, array_index_513374[2:0]} : sel_525935;
  assign add_526641 = array_index_513533[11:3] + 9'h1f1;
  assign sel_526643 = $signed({1'h0, add_525937, array_index_513377[2:0]}) < $signed({1'h0, sel_525939}) ? {add_525937, array_index_513377[2:0]} : sel_525939;
  assign add_526653 = array_index_513890[11:0] + 12'h081;
  assign sel_526655 = $signed({1'h0, add_525949}) < $signed({1'h0, sel_525951}) ? add_525949 : sel_525951;
  assign add_526657 = array_index_513893[11:0] + 12'h081;
  assign sel_526659 = $signed({1'h0, add_525953}) < $signed({1'h0, sel_525955}) ? add_525953 : sel_525955;
  assign add_526671 = array_index_514318[11:0] + 12'h0b1;
  assign sel_526673 = $signed({1'h0, add_525967}) < $signed({1'h0, sel_525969}) ? add_525967 : sel_525969;
  assign add_526675 = array_index_514321[11:0] + 12'h0b1;
  assign sel_526677 = $signed({1'h0, add_525971}) < $signed({1'h0, sel_525973}) ? add_525971 : sel_525973;
  assign add_526689 = array_index_514818[11:1] + 11'h4c1;
  assign sel_526691 = $signed({1'h0, add_525985, array_index_514558[0]}) < $signed({1'h0, sel_525987}) ? {add_525985, array_index_514558[0]} : sel_525987;
  assign add_526693 = array_index_514821[11:1] + 11'h4c1;
  assign sel_526695 = $signed({1'h0, add_525989, array_index_514561[0]}) < $signed({1'h0, sel_525991}) ? {add_525989, array_index_514561[0]} : sel_525991;
  assign add_526705 = array_index_515398[11:0] + 12'hbb1;
  assign sel_526707 = $signed({1'h0, add_526001}) < $signed({1'h0, sel_526003}) ? add_526001 : sel_526003;
  assign add_526709 = array_index_515401[11:0] + 12'hbb1;
  assign sel_526711 = $signed({1'h0, add_526005}) < $signed({1'h0, sel_526007}) ? add_526005 : sel_526007;
  assign add_526721 = array_index_516080[11:0] + 12'h6ab;
  assign sel_526723 = $signed({1'h0, add_526017}) < $signed({1'h0, sel_526019}) ? add_526017 : sel_526019;
  assign add_526725 = array_index_516083[11:0] + 12'h6ab;
  assign sel_526727 = $signed({1'h0, add_526021}) < $signed({1'h0, sel_526023}) ? add_526021 : sel_526023;
  assign add_526737 = array_index_516860[11:0] + 12'h7d5;
  assign sel_526739 = $signed({1'h0, add_526033}) < $signed({1'h0, sel_526035}) ? add_526033 : sel_526035;
  assign add_526741 = array_index_516863[11:0] + 12'h7d5;
  assign sel_526743 = $signed({1'h0, add_526037}) < $signed({1'h0, sel_526039}) ? add_526037 : sel_526039;
  assign add_526787 = concat_526566 + 7'h01;
  assign add_526795 = array_index_512834[11:0] + 12'ha87;
  assign sel_526797 = $signed({1'h0, add_526089}) < $signed(13'h0fff) ? add_526089 : 12'hfff;
  assign add_526799 = array_index_512837[11:0] + 12'ha87;
  assign sel_526801 = $signed({1'h0, add_526091}) < $signed(13'h0fff) ? add_526091 : 12'hfff;
  assign add_526813 = array_index_512942[11:1] + 11'h663;
  assign sel_526815 = $signed({1'h0, add_526105, array_index_512880[0]}) < $signed({1'h0, sel_526107}) ? {add_526105, array_index_512880[0]} : sel_526107;
  assign add_526817 = array_index_512945[11:1] + 11'h663;
  assign sel_526819 = $signed({1'h0, add_526109, array_index_512883[0]}) < $signed({1'h0, sel_526111}) ? {add_526109, array_index_512883[0]} : sel_526111;
  assign add_526829 = array_index_513120[11:1] + 11'h075;
  assign sel_526831 = $signed({1'h0, add_526121, array_index_513022[0]}) < $signed({1'h0, sel_526123}) ? {add_526121, array_index_513022[0]} : sel_526123;
  assign add_526833 = array_index_513123[11:1] + 11'h075;
  assign sel_526835 = $signed({1'h0, add_526125, array_index_513025[0]}) < $signed({1'h0, sel_526127}) ? {add_526125, array_index_513025[0]} : sel_526127;
  assign add_526847 = array_index_513374[11:2] + 10'h181;
  assign sel_526849 = $signed({1'h0, add_526139, array_index_513238[1:0]}) < $signed({1'h0, sel_526141}) ? {add_526139, array_index_513238[1:0]} : sel_526141;
  assign add_526851 = array_index_513377[11:2] + 10'h181;
  assign sel_526853 = $signed({1'h0, add_526143, array_index_513241[1:0]}) < $signed({1'h0, sel_526145}) ? {add_526143, array_index_513241[1:0]} : sel_526145;
  assign add_526865 = array_index_513702[11:0] + 12'h8a7;
  assign sel_526867 = $signed({1'h0, add_526157}) < $signed({1'h0, sel_526159}) ? add_526157 : sel_526159;
  assign add_526869 = array_index_513705[11:0] + 12'h8a7;
  assign sel_526871 = $signed({1'h0, add_526161}) < $signed({1'h0, sel_526163}) ? add_526161 : sel_526163;
  assign add_526883 = array_index_514096[11:1] + 11'h283;
  assign sel_526885 = $signed({1'h0, add_526175, array_index_513890[0]}) < $signed({1'h0, sel_526177}) ? {add_526175, array_index_513890[0]} : sel_526177;
  assign add_526887 = array_index_514099[11:1] + 11'h283;
  assign sel_526889 = $signed({1'h0, add_526179, array_index_513893[0]}) < $signed({1'h0, sel_526181}) ? {add_526179, array_index_513893[0]} : sel_526181;
  assign add_526899 = array_index_514558[11:1] + 11'h44d;
  assign sel_526901 = $signed({1'h0, add_526191, array_index_514318[0]}) < $signed({1'h0, sel_526193}) ? {add_526191, array_index_514318[0]} : sel_526193;
  assign add_526903 = array_index_514561[11:1] + 11'h44d;
  assign sel_526905 = $signed({1'h0, add_526195, array_index_514321[0]}) < $signed({1'h0, sel_526197}) ? {add_526195, array_index_514321[0]} : sel_526197;
  assign add_526915 = array_index_515098[11:0] + 12'hcb1;
  assign sel_526917 = $signed({1'h0, add_526207}) < $signed({1'h0, sel_526209}) ? add_526207 : sel_526209;
  assign add_526919 = array_index_515101[11:0] + 12'hcb1;
  assign sel_526921 = $signed({1'h0, add_526211}) < $signed({1'h0, sel_526213}) ? add_526211 : sel_526213;
  assign add_526931 = array_index_515726[11:0] + 12'h81f;
  assign sel_526933 = $signed({1'h0, add_526223}) < $signed({1'h0, sel_526225}) ? add_526223 : sel_526225;
  assign add_526935 = array_index_515729[11:0] + 12'h81f;
  assign sel_526937 = $signed({1'h0, add_526227}) < $signed({1'h0, sel_526229}) ? add_526227 : sel_526229;
  assign add_526947 = array_index_516458[11:0] + 12'h45b;
  assign sel_526949 = $signed({1'h0, add_526239}) < $signed({1'h0, sel_526241}) ? add_526239 : sel_526241;
  assign add_526951 = array_index_516461[11:0] + 12'h45b;
  assign sel_526953 = $signed({1'h0, add_526243}) < $signed({1'h0, sel_526245}) ? add_526243 : sel_526245;
  assign add_526965 = array_index_517286[11:3] + 9'h0f5;
  assign sel_526967 = $signed({1'h0, add_526257, array_index_516860[2:0]}) < $signed({1'h0, sel_526259}) ? {add_526257, array_index_516860[2:0]} : sel_526259;
  assign add_526969 = array_index_517289[11:3] + 9'h0f5;
  assign sel_526971 = $signed({1'h0, add_526261, array_index_516863[2:0]}) < $signed({1'h0, sel_526263}) ? {add_526261, array_index_516863[2:0]} : sel_526263;
  assign add_527021 = array_index_512818[11:2] + 10'h113;
  assign add_527023 = array_index_512819[11:2] + 10'h113;
  assign add_527037 = array_index_512880[11:4] + 8'h49;
  assign sel_527039 = $signed({1'h0, add_526325, array_index_512834[3:0]}) < $signed({1'h0, sel_526327}) ? {add_526325, array_index_512834[3:0]} : sel_526327;
  assign add_527041 = array_index_512883[11:4] + 8'h49;
  assign sel_527043 = $signed({1'h0, add_526329, array_index_512837[3:0]}) < $signed({1'h0, sel_526331}) ? {add_526329, array_index_512837[3:0]} : sel_526331;
  assign add_527053 = array_index_513022[11:0] + 12'h263;
  assign sel_527055 = $signed({1'h0, add_526341}) < $signed({1'h0, sel_526343}) ? add_526341 : sel_526343;
  assign add_527057 = array_index_513025[11:0] + 12'h263;
  assign sel_527059 = $signed({1'h0, add_526345}) < $signed({1'h0, sel_526347}) ? add_526345 : sel_526347;
  assign add_527069 = array_index_513238[11:1] + 11'h109;
  assign sel_527071 = $signed({1'h0, add_526357, array_index_513120[0]}) < $signed({1'h0, sel_526359}) ? {add_526357, array_index_513120[0]} : sel_526359;
  assign add_527073 = array_index_513241[11:1] + 11'h109;
  assign sel_527075 = $signed({1'h0, add_526361, array_index_513123[0]}) < $signed({1'h0, sel_526363}) ? {add_526361, array_index_513123[0]} : sel_526363;
  assign add_527085 = array_index_513530[11:3] + 9'h12f;
  assign sel_527087 = $signed({1'h0, add_526373, array_index_513374[2:0]}) < $signed({1'h0, sel_526375}) ? {add_526373, array_index_513374[2:0]} : sel_526375;
  assign add_527089 = array_index_513533[11:3] + 9'h12f;
  assign sel_527091 = $signed({1'h0, add_526377, array_index_513377[2:0]}) < $signed({1'h0, sel_526379}) ? {add_526377, array_index_513377[2:0]} : sel_526379;
  assign add_527103 = array_index_513890[11:3] + 9'h171;
  assign sel_527105 = $signed({1'h0, add_526391, array_index_513702[2:0]}) < $signed({1'h0, sel_526393}) ? {add_526391, array_index_513702[2:0]} : sel_526393;
  assign add_527107 = array_index_513893[11:3] + 9'h171;
  assign sel_527109 = $signed({1'h0, add_526395, array_index_513705[2:0]}) < $signed({1'h0, sel_526397}) ? {add_526395, array_index_513705[2:0]} : sel_526397;
  assign add_527119 = array_index_514318[11:0] + 12'h091;
  assign sel_527121 = $signed({1'h0, add_526407}) < $signed({1'h0, sel_526409}) ? add_526407 : sel_526409;
  assign add_527123 = array_index_514321[11:0] + 12'h091;
  assign sel_527125 = $signed({1'h0, add_526411}) < $signed({1'h0, sel_526413}) ? add_526411 : sel_526413;
  assign add_527135 = array_index_514818[11:0] + 12'hf59;
  assign sel_527137 = $signed({1'h0, add_526423}) < $signed({1'h0, sel_526425}) ? add_526423 : sel_526425;
  assign add_527139 = array_index_514821[11:0] + 12'hf59;
  assign sel_527141 = $signed({1'h0, add_526427}) < $signed({1'h0, sel_526429}) ? add_526427 : sel_526429;
  assign add_527153 = array_index_515398[11:0] + 12'h437;
  assign sel_527155 = $signed({1'h0, add_526441}) < $signed({1'h0, sel_526443}) ? add_526441 : sel_526443;
  assign add_527157 = array_index_515401[11:0] + 12'h437;
  assign sel_527159 = $signed({1'h0, add_526445}) < $signed({1'h0, sel_526447}) ? add_526445 : sel_526447;
  assign add_527169 = array_index_516080[11:0] + 12'hee1;
  assign sel_527171 = $signed({1'h0, add_526457}) < $signed({1'h0, sel_526459}) ? add_526457 : sel_526459;
  assign add_527173 = array_index_516083[11:0] + 12'hee1;
  assign sel_527175 = $signed({1'h0, add_526461}) < $signed({1'h0, sel_526463}) ? add_526461 : sel_526463;
  assign add_527185 = array_index_516860[11:1] + 11'h179;
  assign sel_527187 = $signed({1'h0, add_526473, array_index_516458[0]}) < $signed({1'h0, sel_526475}) ? {add_526473, array_index_516458[0]} : sel_526475;
  assign add_527189 = array_index_516863[11:1] + 11'h179;
  assign sel_527191 = $signed({1'h0, add_526477, array_index_516461[0]}) < $signed({1'h0, sel_526479}) ? {add_526477, array_index_516461[0]} : sel_526479;
  assign add_527201 = array_index_517736[11:0] + 12'h067;
  assign sel_527203 = $signed({1'h0, add_526489}) < $signed({1'h0, sel_526491}) ? add_526489 : sel_526491;
  assign add_527205 = array_index_517739[11:0] + 12'h067;
  assign sel_527207 = $signed({1'h0, add_526493}) < $signed({1'h0, sel_526495}) ? add_526493 : sel_526495;
  assign add_527209 = array_index_518210[11:3] + 9'h1ef;
  assign sel_527212 = $signed({1'h0, add_526497, array_index_517736[2:0]}) < $signed({1'h0, sel_526500}) ? {add_526497, array_index_517736[2:0]} : sel_526500;
  assign add_527214 = array_index_518213[11:3] + 9'h1ef;
  assign sel_527217 = $signed({1'h0, add_526502, array_index_517739[2:0]}) < $signed({1'h0, sel_526505}) ? {add_526502, array_index_517739[2:0]} : sel_526505;
  assign add_527219 = array_index_518710[11:1] + 11'h2d5;
  assign sel_527221 = $signed({1'h0, add_526507, array_index_518210[0]}) < $signed({1'h0, sel_526509}) ? {add_526507, array_index_518210[0]} : sel_526509;
  assign add_527223 = array_index_518713[11:1] + 11'h2d5;
  assign sel_527225 = $signed({1'h0, add_526511, array_index_518213[0]}) < $signed({1'h0, sel_526513}) ? {add_526511, array_index_518213[0]} : sel_526513;
  assign add_527227 = array_index_519236[11:2] + 10'h353;
  assign sel_527229 = $signed({1'h0, add_526515, array_index_518710[1:0]}) < $signed({1'h0, sel_526517}) ? {add_526515, array_index_518710[1:0]} : sel_526517;
  assign add_527231 = array_index_519239[11:2] + 10'h353;
  assign sel_527233 = $signed({1'h0, add_526519, array_index_518713[1:0]}) < $signed({1'h0, sel_526521}) ? {add_526519, array_index_518713[1:0]} : sel_526521;
  assign add_527235 = array_index_519786[11:0] + 12'h0a7;
  assign sel_527237 = $signed({1'h0, add_526523}) < $signed({1'h0, sel_526525}) ? add_526523 : sel_526525;
  assign add_527239 = array_index_519789[11:0] + 12'h0a7;
  assign sel_527241 = $signed({1'h0, add_526527}) < $signed({1'h0, sel_526529}) ? add_526527 : sel_526529;
  assign add_527243 = array_index_520362[11:1] + 11'h4cb;
  assign sel_527245 = $signed({1'h0, add_526531, array_index_519786[0]}) < $signed({1'h0, sel_526533}) ? {add_526531, array_index_519786[0]} : sel_526533;
  assign add_527247 = array_index_520365[11:1] + 11'h4cb;
  assign sel_527249 = $signed({1'h0, add_526535, array_index_519789[0]}) < $signed({1'h0, sel_526537}) ? {add_526535, array_index_519789[0]} : sel_526537;
  assign add_527251 = array_index_520964[11:0] + 12'hfe9;
  assign sel_527253 = $signed({1'h0, add_526539}) < $signed({1'h0, sel_526541}) ? add_526539 : sel_526541;
  assign add_527255 = array_index_520967[11:0] + 12'hfe9;
  assign sel_527257 = $signed({1'h0, add_526543}) < $signed({1'h0, sel_526545}) ? add_526543 : sel_526545;
  assign add_527259 = array_index_521590[11:0] + 12'h97d;
  assign sel_527261 = $signed({1'h0, add_526547}) < $signed({1'h0, sel_526549}) ? add_526547 : sel_526549;
  assign add_527263 = array_index_521593[11:0] + 12'h97d;
  assign sel_527265 = $signed({1'h0, add_526551}) < $signed({1'h0, sel_526553}) ? add_526551 : sel_526553;
  assign concat_527268 = {1'h0, ($signed({1'h0, add_525861}) < $signed({1'h0, sel_525863}) ? add_525861 : sel_525863) == ($signed({1'h0, add_525865}) < $signed({1'h0, sel_525867}) ? add_525865 : sel_525867) ? add_526787 : concat_526566};
  assign add_527277 = array_index_512834[11:1] + 11'h5b9;
  assign sel_527279 = $signed({1'h0, add_526569, array_index_512818[0]}) < $signed(13'h0fff) ? {add_526569, array_index_512818[0]} : 12'hfff;
  assign add_527281 = array_index_512837[11:1] + 11'h5b9;
  assign sel_527283 = $signed({1'h0, add_526571, array_index_512819[0]}) < $signed(13'h0fff) ? {add_526571, array_index_512819[0]} : 12'hfff;
  assign add_527293 = array_index_512942[11:0] + 12'h37b;
  assign sel_527295 = $signed({1'h0, add_526583}) < $signed({1'h0, sel_526585}) ? add_526583 : sel_526585;
  assign add_527297 = array_index_512945[11:0] + 12'h37b;
  assign sel_527299 = $signed({1'h0, add_526587}) < $signed({1'h0, sel_526589}) ? add_526587 : sel_526589;
  assign add_527311 = array_index_513120[11:0] + 12'h811;
  assign sel_527313 = $signed({1'h0, add_526601}) < $signed({1'h0, sel_526603}) ? add_526601 : sel_526603;
  assign add_527315 = array_index_513123[11:0] + 12'h811;
  assign sel_527317 = $signed({1'h0, add_526605}) < $signed({1'h0, sel_526607}) ? add_526605 : sel_526607;
  assign add_527329 = array_index_513374[11:0] + 12'h70f;
  assign sel_527331 = $signed({1'h0, add_526619}) < $signed({1'h0, sel_526621}) ? add_526619 : sel_526621;
  assign add_527333 = array_index_513377[11:0] + 12'h70f;
  assign sel_527335 = $signed({1'h0, add_526623}) < $signed({1'h0, sel_526625}) ? add_526623 : sel_526625;
  assign add_527347 = array_index_513702[11:3] + 9'h1f1;
  assign sel_527349 = $signed({1'h0, add_526637, array_index_513530[2:0]}) < $signed({1'h0, sel_526639}) ? {add_526637, array_index_513530[2:0]} : sel_526639;
  assign add_527351 = array_index_513705[11:3] + 9'h1f1;
  assign sel_527353 = $signed({1'h0, add_526641, array_index_513533[2:0]}) < $signed({1'h0, sel_526643}) ? {add_526641, array_index_513533[2:0]} : sel_526643;
  assign add_527363 = array_index_514096[11:0] + 12'h081;
  assign sel_527365 = $signed({1'h0, add_526653}) < $signed({1'h0, sel_526655}) ? add_526653 : sel_526655;
  assign add_527367 = array_index_514099[11:0] + 12'h081;
  assign sel_527369 = $signed({1'h0, add_526657}) < $signed({1'h0, sel_526659}) ? add_526657 : sel_526659;
  assign add_527381 = array_index_514558[11:0] + 12'h0b1;
  assign sel_527383 = $signed({1'h0, add_526671}) < $signed({1'h0, sel_526673}) ? add_526671 : sel_526673;
  assign add_527385 = array_index_514561[11:0] + 12'h0b1;
  assign sel_527387 = $signed({1'h0, add_526675}) < $signed({1'h0, sel_526677}) ? add_526675 : sel_526677;
  assign add_527399 = array_index_515098[11:1] + 11'h4c1;
  assign sel_527401 = $signed({1'h0, add_526689, array_index_514818[0]}) < $signed({1'h0, sel_526691}) ? {add_526689, array_index_514818[0]} : sel_526691;
  assign add_527403 = array_index_515101[11:1] + 11'h4c1;
  assign sel_527405 = $signed({1'h0, add_526693, array_index_514821[0]}) < $signed({1'h0, sel_526695}) ? {add_526693, array_index_514821[0]} : sel_526695;
  assign add_527415 = array_index_515726[11:0] + 12'hbb1;
  assign sel_527417 = $signed({1'h0, add_526705}) < $signed({1'h0, sel_526707}) ? add_526705 : sel_526707;
  assign add_527419 = array_index_515729[11:0] + 12'hbb1;
  assign sel_527421 = $signed({1'h0, add_526709}) < $signed({1'h0, sel_526711}) ? add_526709 : sel_526711;
  assign add_527431 = array_index_516458[11:0] + 12'h6ab;
  assign sel_527433 = $signed({1'h0, add_526721}) < $signed({1'h0, sel_526723}) ? add_526721 : sel_526723;
  assign add_527435 = array_index_516461[11:0] + 12'h6ab;
  assign sel_527437 = $signed({1'h0, add_526725}) < $signed({1'h0, sel_526727}) ? add_526725 : sel_526727;
  assign add_527447 = array_index_517286[11:0] + 12'h7d5;
  assign sel_527449 = $signed({1'h0, add_526737}) < $signed({1'h0, sel_526739}) ? add_526737 : sel_526739;
  assign add_527451 = array_index_517289[11:0] + 12'h7d5;
  assign sel_527453 = $signed({1'h0, add_526741}) < $signed({1'h0, sel_526743}) ? add_526741 : sel_526743;
  assign add_527493 = concat_527268 + 8'h01;
  assign add_527495 = array_index_512818[11:0] + 12'hcc1;
  assign add_527497 = array_index_512819[11:0] + 12'hcc1;
  assign add_527511 = array_index_512880[11:0] + 12'ha87;
  assign sel_527513 = $signed({1'h0, add_526795}) < $signed({1'h0, sel_526797}) ? add_526795 : sel_526797;
  assign add_527515 = array_index_512883[11:0] + 12'ha87;
  assign sel_527517 = $signed({1'h0, add_526799}) < $signed({1'h0, sel_526801}) ? add_526799 : sel_526801;
  assign add_527529 = array_index_513022[11:1] + 11'h663;
  assign sel_527531 = $signed({1'h0, add_526813, array_index_512942[0]}) < $signed({1'h0, sel_526815}) ? {add_526813, array_index_512942[0]} : sel_526815;
  assign add_527533 = array_index_513025[11:1] + 11'h663;
  assign sel_527535 = $signed({1'h0, add_526817, array_index_512945[0]}) < $signed({1'h0, sel_526819}) ? {add_526817, array_index_512945[0]} : sel_526819;
  assign add_527545 = array_index_513238[11:1] + 11'h075;
  assign sel_527547 = $signed({1'h0, add_526829, array_index_513120[0]}) < $signed({1'h0, sel_526831}) ? {add_526829, array_index_513120[0]} : sel_526831;
  assign add_527549 = array_index_513241[11:1] + 11'h075;
  assign sel_527551 = $signed({1'h0, add_526833, array_index_513123[0]}) < $signed({1'h0, sel_526835}) ? {add_526833, array_index_513123[0]} : sel_526835;
  assign add_527563 = array_index_513530[11:2] + 10'h181;
  assign sel_527565 = $signed({1'h0, add_526847, array_index_513374[1:0]}) < $signed({1'h0, sel_526849}) ? {add_526847, array_index_513374[1:0]} : sel_526849;
  assign add_527567 = array_index_513533[11:2] + 10'h181;
  assign sel_527569 = $signed({1'h0, add_526851, array_index_513377[1:0]}) < $signed({1'h0, sel_526853}) ? {add_526851, array_index_513377[1:0]} : sel_526853;
  assign add_527581 = array_index_513890[11:0] + 12'h8a7;
  assign sel_527583 = $signed({1'h0, add_526865}) < $signed({1'h0, sel_526867}) ? add_526865 : sel_526867;
  assign add_527585 = array_index_513893[11:0] + 12'h8a7;
  assign sel_527587 = $signed({1'h0, add_526869}) < $signed({1'h0, sel_526871}) ? add_526869 : sel_526871;
  assign add_527599 = array_index_514318[11:1] + 11'h283;
  assign sel_527601 = $signed({1'h0, add_526883, array_index_514096[0]}) < $signed({1'h0, sel_526885}) ? {add_526883, array_index_514096[0]} : sel_526885;
  assign add_527603 = array_index_514321[11:1] + 11'h283;
  assign sel_527605 = $signed({1'h0, add_526887, array_index_514099[0]}) < $signed({1'h0, sel_526889}) ? {add_526887, array_index_514099[0]} : sel_526889;
  assign add_527615 = array_index_514818[11:1] + 11'h44d;
  assign sel_527617 = $signed({1'h0, add_526899, array_index_514558[0]}) < $signed({1'h0, sel_526901}) ? {add_526899, array_index_514558[0]} : sel_526901;
  assign add_527619 = array_index_514821[11:1] + 11'h44d;
  assign sel_527621 = $signed({1'h0, add_526903, array_index_514561[0]}) < $signed({1'h0, sel_526905}) ? {add_526903, array_index_514561[0]} : sel_526905;
  assign add_527631 = array_index_515398[11:0] + 12'hcb1;
  assign sel_527633 = $signed({1'h0, add_526915}) < $signed({1'h0, sel_526917}) ? add_526915 : sel_526917;
  assign add_527635 = array_index_515401[11:0] + 12'hcb1;
  assign sel_527637 = $signed({1'h0, add_526919}) < $signed({1'h0, sel_526921}) ? add_526919 : sel_526921;
  assign add_527647 = array_index_516080[11:0] + 12'h81f;
  assign sel_527649 = $signed({1'h0, add_526931}) < $signed({1'h0, sel_526933}) ? add_526931 : sel_526933;
  assign add_527651 = array_index_516083[11:0] + 12'h81f;
  assign sel_527653 = $signed({1'h0, add_526935}) < $signed({1'h0, sel_526937}) ? add_526935 : sel_526937;
  assign add_527663 = array_index_516860[11:0] + 12'h45b;
  assign sel_527665 = $signed({1'h0, add_526947}) < $signed({1'h0, sel_526949}) ? add_526947 : sel_526949;
  assign add_527667 = array_index_516863[11:0] + 12'h45b;
  assign sel_527669 = $signed({1'h0, add_526951}) < $signed({1'h0, sel_526953}) ? add_526951 : sel_526953;
  assign add_527681 = array_index_517736[11:3] + 9'h0f5;
  assign sel_527683 = $signed({1'h0, add_526965, array_index_517286[2:0]}) < $signed({1'h0, sel_526967}) ? {add_526965, array_index_517286[2:0]} : sel_526967;
  assign add_527685 = array_index_517739[11:3] + 9'h0f5;
  assign sel_527687 = $signed({1'h0, add_526969, array_index_517289[2:0]}) < $signed({1'h0, sel_526971}) ? {add_526969, array_index_517289[2:0]} : sel_526971;
  assign add_527735 = array_index_512834[11:2] + 10'h113;
  assign sel_527737 = $signed({1'h0, add_527021, array_index_512818[1:0]}) < $signed(13'h0fff) ? {add_527021, array_index_512818[1:0]} : 12'hfff;
  assign add_527739 = array_index_512837[11:2] + 10'h113;
  assign sel_527741 = $signed({1'h0, add_527023, array_index_512819[1:0]}) < $signed(13'h0fff) ? {add_527023, array_index_512819[1:0]} : 12'hfff;
  assign add_527753 = array_index_512942[11:4] + 8'h49;
  assign sel_527755 = $signed({1'h0, add_527037, array_index_512880[3:0]}) < $signed({1'h0, sel_527039}) ? {add_527037, array_index_512880[3:0]} : sel_527039;
  assign add_527757 = array_index_512945[11:4] + 8'h49;
  assign sel_527759 = $signed({1'h0, add_527041, array_index_512883[3:0]}) < $signed({1'h0, sel_527043}) ? {add_527041, array_index_512883[3:0]} : sel_527043;
  assign add_527769 = array_index_513120[11:0] + 12'h263;
  assign sel_527771 = $signed({1'h0, add_527053}) < $signed({1'h0, sel_527055}) ? add_527053 : sel_527055;
  assign add_527773 = array_index_513123[11:0] + 12'h263;
  assign sel_527775 = $signed({1'h0, add_527057}) < $signed({1'h0, sel_527059}) ? add_527057 : sel_527059;
  assign add_527785 = array_index_513374[11:1] + 11'h109;
  assign sel_527787 = $signed({1'h0, add_527069, array_index_513238[0]}) < $signed({1'h0, sel_527071}) ? {add_527069, array_index_513238[0]} : sel_527071;
  assign add_527789 = array_index_513377[11:1] + 11'h109;
  assign sel_527791 = $signed({1'h0, add_527073, array_index_513241[0]}) < $signed({1'h0, sel_527075}) ? {add_527073, array_index_513241[0]} : sel_527075;
  assign add_527801 = array_index_513702[11:3] + 9'h12f;
  assign sel_527803 = $signed({1'h0, add_527085, array_index_513530[2:0]}) < $signed({1'h0, sel_527087}) ? {add_527085, array_index_513530[2:0]} : sel_527087;
  assign add_527805 = array_index_513705[11:3] + 9'h12f;
  assign sel_527807 = $signed({1'h0, add_527089, array_index_513533[2:0]}) < $signed({1'h0, sel_527091}) ? {add_527089, array_index_513533[2:0]} : sel_527091;
  assign add_527819 = array_index_514096[11:3] + 9'h171;
  assign sel_527821 = $signed({1'h0, add_527103, array_index_513890[2:0]}) < $signed({1'h0, sel_527105}) ? {add_527103, array_index_513890[2:0]} : sel_527105;
  assign add_527823 = array_index_514099[11:3] + 9'h171;
  assign sel_527825 = $signed({1'h0, add_527107, array_index_513893[2:0]}) < $signed({1'h0, sel_527109}) ? {add_527107, array_index_513893[2:0]} : sel_527109;
  assign add_527835 = array_index_514558[11:0] + 12'h091;
  assign sel_527837 = $signed({1'h0, add_527119}) < $signed({1'h0, sel_527121}) ? add_527119 : sel_527121;
  assign add_527839 = array_index_514561[11:0] + 12'h091;
  assign sel_527841 = $signed({1'h0, add_527123}) < $signed({1'h0, sel_527125}) ? add_527123 : sel_527125;
  assign add_527851 = array_index_515098[11:0] + 12'hf59;
  assign sel_527853 = $signed({1'h0, add_527135}) < $signed({1'h0, sel_527137}) ? add_527135 : sel_527137;
  assign add_527855 = array_index_515101[11:0] + 12'hf59;
  assign sel_527857 = $signed({1'h0, add_527139}) < $signed({1'h0, sel_527141}) ? add_527139 : sel_527141;
  assign add_527869 = array_index_515726[11:0] + 12'h437;
  assign sel_527871 = $signed({1'h0, add_527153}) < $signed({1'h0, sel_527155}) ? add_527153 : sel_527155;
  assign add_527873 = array_index_515729[11:0] + 12'h437;
  assign sel_527875 = $signed({1'h0, add_527157}) < $signed({1'h0, sel_527159}) ? add_527157 : sel_527159;
  assign add_527885 = array_index_516458[11:0] + 12'hee1;
  assign sel_527887 = $signed({1'h0, add_527169}) < $signed({1'h0, sel_527171}) ? add_527169 : sel_527171;
  assign add_527889 = array_index_516461[11:0] + 12'hee1;
  assign sel_527891 = $signed({1'h0, add_527173}) < $signed({1'h0, sel_527175}) ? add_527173 : sel_527175;
  assign add_527901 = array_index_517286[11:1] + 11'h179;
  assign sel_527903 = $signed({1'h0, add_527185, array_index_516860[0]}) < $signed({1'h0, sel_527187}) ? {add_527185, array_index_516860[0]} : sel_527187;
  assign add_527905 = array_index_517289[11:1] + 11'h179;
  assign sel_527907 = $signed({1'h0, add_527189, array_index_516863[0]}) < $signed({1'h0, sel_527191}) ? {add_527189, array_index_516863[0]} : sel_527191;
  assign add_527917 = array_index_518210[11:0] + 12'h067;
  assign sel_527919 = $signed({1'h0, add_527201}) < $signed({1'h0, sel_527203}) ? add_527201 : sel_527203;
  assign add_527921 = array_index_518213[11:0] + 12'h067;
  assign sel_527923 = $signed({1'h0, add_527205}) < $signed({1'h0, sel_527207}) ? add_527205 : sel_527207;
  assign add_527925 = array_index_518710[11:3] + 9'h1ef;
  assign sel_527928 = $signed({1'h0, add_527209, array_index_518210[2:0]}) < $signed({1'h0, sel_527212}) ? {add_527209, array_index_518210[2:0]} : sel_527212;
  assign add_527930 = array_index_518713[11:3] + 9'h1ef;
  assign sel_527933 = $signed({1'h0, add_527214, array_index_518213[2:0]}) < $signed({1'h0, sel_527217}) ? {add_527214, array_index_518213[2:0]} : sel_527217;
  assign add_527935 = array_index_519236[11:1] + 11'h2d5;
  assign sel_527937 = $signed({1'h0, add_527219, array_index_518710[0]}) < $signed({1'h0, sel_527221}) ? {add_527219, array_index_518710[0]} : sel_527221;
  assign add_527939 = array_index_519239[11:1] + 11'h2d5;
  assign sel_527941 = $signed({1'h0, add_527223, array_index_518713[0]}) < $signed({1'h0, sel_527225}) ? {add_527223, array_index_518713[0]} : sel_527225;
  assign add_527943 = array_index_519786[11:2] + 10'h353;
  assign sel_527945 = $signed({1'h0, add_527227, array_index_519236[1:0]}) < $signed({1'h0, sel_527229}) ? {add_527227, array_index_519236[1:0]} : sel_527229;
  assign add_527947 = array_index_519789[11:2] + 10'h353;
  assign sel_527949 = $signed({1'h0, add_527231, array_index_519239[1:0]}) < $signed({1'h0, sel_527233}) ? {add_527231, array_index_519239[1:0]} : sel_527233;
  assign add_527951 = array_index_520362[11:0] + 12'h0a7;
  assign sel_527953 = $signed({1'h0, add_527235}) < $signed({1'h0, sel_527237}) ? add_527235 : sel_527237;
  assign add_527955 = array_index_520365[11:0] + 12'h0a7;
  assign sel_527957 = $signed({1'h0, add_527239}) < $signed({1'h0, sel_527241}) ? add_527239 : sel_527241;
  assign add_527959 = array_index_520964[11:1] + 11'h4cb;
  assign sel_527961 = $signed({1'h0, add_527243, array_index_520362[0]}) < $signed({1'h0, sel_527245}) ? {add_527243, array_index_520362[0]} : sel_527245;
  assign add_527963 = array_index_520967[11:1] + 11'h4cb;
  assign sel_527965 = $signed({1'h0, add_527247, array_index_520365[0]}) < $signed({1'h0, sel_527249}) ? {add_527247, array_index_520365[0]} : sel_527249;
  assign add_527967 = array_index_521590[11:0] + 12'hfe9;
  assign sel_527969 = $signed({1'h0, add_527251}) < $signed({1'h0, sel_527253}) ? add_527251 : sel_527253;
  assign add_527971 = array_index_521593[11:0] + 12'hfe9;
  assign sel_527973 = $signed({1'h0, add_527255}) < $signed({1'h0, sel_527257}) ? add_527255 : sel_527257;
  assign concat_527976 = {1'h0, ($signed({1'h0, add_526555, array_index_521590[1:0]}) < $signed({1'h0, sel_526558}) ? {add_526555, array_index_521590[1:0]} : sel_526558) == ($signed({1'h0, add_526560, array_index_521593[1:0]}) < $signed({1'h0, sel_526563}) ? {add_526560, array_index_521593[1:0]} : sel_526563) ? add_527493 : concat_527268};
  assign add_527989 = array_index_512880[11:1] + 11'h5b9;
  assign sel_527991 = $signed({1'h0, add_527277, array_index_512834[0]}) < $signed({1'h0, sel_527279}) ? {add_527277, array_index_512834[0]} : sel_527279;
  assign add_527993 = array_index_512883[11:1] + 11'h5b9;
  assign sel_527995 = $signed({1'h0, add_527281, array_index_512837[0]}) < $signed({1'h0, sel_527283}) ? {add_527281, array_index_512837[0]} : sel_527283;
  assign add_528005 = array_index_513022[11:0] + 12'h37b;
  assign sel_528007 = $signed({1'h0, add_527293}) < $signed({1'h0, sel_527295}) ? add_527293 : sel_527295;
  assign add_528009 = array_index_513025[11:0] + 12'h37b;
  assign sel_528011 = $signed({1'h0, add_527297}) < $signed({1'h0, sel_527299}) ? add_527297 : sel_527299;
  assign add_528023 = array_index_513238[11:0] + 12'h811;
  assign sel_528025 = $signed({1'h0, add_527311}) < $signed({1'h0, sel_527313}) ? add_527311 : sel_527313;
  assign add_528027 = array_index_513241[11:0] + 12'h811;
  assign sel_528029 = $signed({1'h0, add_527315}) < $signed({1'h0, sel_527317}) ? add_527315 : sel_527317;
  assign add_528041 = array_index_513530[11:0] + 12'h70f;
  assign sel_528043 = $signed({1'h0, add_527329}) < $signed({1'h0, sel_527331}) ? add_527329 : sel_527331;
  assign add_528045 = array_index_513533[11:0] + 12'h70f;
  assign sel_528047 = $signed({1'h0, add_527333}) < $signed({1'h0, sel_527335}) ? add_527333 : sel_527335;
  assign add_528059 = array_index_513890[11:3] + 9'h1f1;
  assign sel_528061 = $signed({1'h0, add_527347, array_index_513702[2:0]}) < $signed({1'h0, sel_527349}) ? {add_527347, array_index_513702[2:0]} : sel_527349;
  assign add_528063 = array_index_513893[11:3] + 9'h1f1;
  assign sel_528065 = $signed({1'h0, add_527351, array_index_513705[2:0]}) < $signed({1'h0, sel_527353}) ? {add_527351, array_index_513705[2:0]} : sel_527353;
  assign add_528075 = array_index_514318[11:0] + 12'h081;
  assign sel_528077 = $signed({1'h0, add_527363}) < $signed({1'h0, sel_527365}) ? add_527363 : sel_527365;
  assign add_528079 = array_index_514321[11:0] + 12'h081;
  assign sel_528081 = $signed({1'h0, add_527367}) < $signed({1'h0, sel_527369}) ? add_527367 : sel_527369;
  assign add_528093 = array_index_514818[11:0] + 12'h0b1;
  assign sel_528095 = $signed({1'h0, add_527381}) < $signed({1'h0, sel_527383}) ? add_527381 : sel_527383;
  assign add_528097 = array_index_514821[11:0] + 12'h0b1;
  assign sel_528099 = $signed({1'h0, add_527385}) < $signed({1'h0, sel_527387}) ? add_527385 : sel_527387;
  assign add_528111 = array_index_515398[11:1] + 11'h4c1;
  assign sel_528113 = $signed({1'h0, add_527399, array_index_515098[0]}) < $signed({1'h0, sel_527401}) ? {add_527399, array_index_515098[0]} : sel_527401;
  assign add_528115 = array_index_515401[11:1] + 11'h4c1;
  assign sel_528117 = $signed({1'h0, add_527403, array_index_515101[0]}) < $signed({1'h0, sel_527405}) ? {add_527403, array_index_515101[0]} : sel_527405;
  assign add_528127 = array_index_516080[11:0] + 12'hbb1;
  assign sel_528129 = $signed({1'h0, add_527415}) < $signed({1'h0, sel_527417}) ? add_527415 : sel_527417;
  assign add_528131 = array_index_516083[11:0] + 12'hbb1;
  assign sel_528133 = $signed({1'h0, add_527419}) < $signed({1'h0, sel_527421}) ? add_527419 : sel_527421;
  assign add_528143 = array_index_516860[11:0] + 12'h6ab;
  assign sel_528145 = $signed({1'h0, add_527431}) < $signed({1'h0, sel_527433}) ? add_527431 : sel_527433;
  assign add_528147 = array_index_516863[11:0] + 12'h6ab;
  assign sel_528149 = $signed({1'h0, add_527435}) < $signed({1'h0, sel_527437}) ? add_527435 : sel_527437;
  assign add_528159 = array_index_517736[11:0] + 12'h7d5;
  assign sel_528161 = $signed({1'h0, add_527447}) < $signed({1'h0, sel_527449}) ? add_527447 : sel_527449;
  assign add_528163 = array_index_517739[11:0] + 12'h7d5;
  assign sel_528165 = $signed({1'h0, add_527451}) < $signed({1'h0, sel_527453}) ? add_527451 : sel_527453;
  assign add_528201 = concat_527976 + 9'h001;
  assign add_528203 = array_index_512834[11:0] + 12'hcc1;
  assign sel_528205 = $signed({1'h0, add_527495}) < $signed(13'h0fff) ? add_527495 : 12'hfff;
  assign add_528207 = array_index_512837[11:0] + 12'hcc1;
  assign sel_528209 = $signed({1'h0, add_527497}) < $signed(13'h0fff) ? add_527497 : 12'hfff;
  assign add_528221 = array_index_512942[11:0] + 12'ha87;
  assign sel_528223 = $signed({1'h0, add_527511}) < $signed({1'h0, sel_527513}) ? add_527511 : sel_527513;
  assign add_528225 = array_index_512945[11:0] + 12'ha87;
  assign sel_528227 = $signed({1'h0, add_527515}) < $signed({1'h0, sel_527517}) ? add_527515 : sel_527517;
  assign add_528239 = array_index_513120[11:1] + 11'h663;
  assign sel_528241 = $signed({1'h0, add_527529, array_index_513022[0]}) < $signed({1'h0, sel_527531}) ? {add_527529, array_index_513022[0]} : sel_527531;
  assign add_528243 = array_index_513123[11:1] + 11'h663;
  assign sel_528245 = $signed({1'h0, add_527533, array_index_513025[0]}) < $signed({1'h0, sel_527535}) ? {add_527533, array_index_513025[0]} : sel_527535;
  assign add_528255 = array_index_513374[11:1] + 11'h075;
  assign sel_528257 = $signed({1'h0, add_527545, array_index_513238[0]}) < $signed({1'h0, sel_527547}) ? {add_527545, array_index_513238[0]} : sel_527547;
  assign add_528259 = array_index_513377[11:1] + 11'h075;
  assign sel_528261 = $signed({1'h0, add_527549, array_index_513241[0]}) < $signed({1'h0, sel_527551}) ? {add_527549, array_index_513241[0]} : sel_527551;
  assign add_528273 = array_index_513702[11:2] + 10'h181;
  assign sel_528275 = $signed({1'h0, add_527563, array_index_513530[1:0]}) < $signed({1'h0, sel_527565}) ? {add_527563, array_index_513530[1:0]} : sel_527565;
  assign add_528277 = array_index_513705[11:2] + 10'h181;
  assign sel_528279 = $signed({1'h0, add_527567, array_index_513533[1:0]}) < $signed({1'h0, sel_527569}) ? {add_527567, array_index_513533[1:0]} : sel_527569;
  assign add_528291 = array_index_514096[11:0] + 12'h8a7;
  assign sel_528293 = $signed({1'h0, add_527581}) < $signed({1'h0, sel_527583}) ? add_527581 : sel_527583;
  assign add_528295 = array_index_514099[11:0] + 12'h8a7;
  assign sel_528297 = $signed({1'h0, add_527585}) < $signed({1'h0, sel_527587}) ? add_527585 : sel_527587;
  assign add_528309 = array_index_514558[11:1] + 11'h283;
  assign sel_528311 = $signed({1'h0, add_527599, array_index_514318[0]}) < $signed({1'h0, sel_527601}) ? {add_527599, array_index_514318[0]} : sel_527601;
  assign add_528313 = array_index_514561[11:1] + 11'h283;
  assign sel_528315 = $signed({1'h0, add_527603, array_index_514321[0]}) < $signed({1'h0, sel_527605}) ? {add_527603, array_index_514321[0]} : sel_527605;
  assign add_528325 = array_index_515098[11:1] + 11'h44d;
  assign sel_528327 = $signed({1'h0, add_527615, array_index_514818[0]}) < $signed({1'h0, sel_527617}) ? {add_527615, array_index_514818[0]} : sel_527617;
  assign add_528329 = array_index_515101[11:1] + 11'h44d;
  assign sel_528331 = $signed({1'h0, add_527619, array_index_514821[0]}) < $signed({1'h0, sel_527621}) ? {add_527619, array_index_514821[0]} : sel_527621;
  assign add_528341 = array_index_515726[11:0] + 12'hcb1;
  assign sel_528343 = $signed({1'h0, add_527631}) < $signed({1'h0, sel_527633}) ? add_527631 : sel_527633;
  assign add_528345 = array_index_515729[11:0] + 12'hcb1;
  assign sel_528347 = $signed({1'h0, add_527635}) < $signed({1'h0, sel_527637}) ? add_527635 : sel_527637;
  assign add_528357 = array_index_516458[11:0] + 12'h81f;
  assign sel_528359 = $signed({1'h0, add_527647}) < $signed({1'h0, sel_527649}) ? add_527647 : sel_527649;
  assign add_528361 = array_index_516461[11:0] + 12'h81f;
  assign sel_528363 = $signed({1'h0, add_527651}) < $signed({1'h0, sel_527653}) ? add_527651 : sel_527653;
  assign add_528373 = array_index_517286[11:0] + 12'h45b;
  assign sel_528375 = $signed({1'h0, add_527663}) < $signed({1'h0, sel_527665}) ? add_527663 : sel_527665;
  assign add_528377 = array_index_517289[11:0] + 12'h45b;
  assign sel_528379 = $signed({1'h0, add_527667}) < $signed({1'h0, sel_527669}) ? add_527667 : sel_527669;
  assign add_528391 = array_index_518210[11:3] + 9'h0f5;
  assign sel_528393 = $signed({1'h0, add_527681, array_index_517736[2:0]}) < $signed({1'h0, sel_527683}) ? {add_527681, array_index_517736[2:0]} : sel_527683;
  assign add_528395 = array_index_518213[11:3] + 9'h0f5;
  assign sel_528397 = $signed({1'h0, add_527685, array_index_517739[2:0]}) < $signed({1'h0, sel_527687}) ? {add_527685, array_index_517739[2:0]} : sel_527687;
  assign add_528441 = array_index_512880[11:2] + 10'h113;
  assign sel_528443 = $signed({1'h0, add_527735, array_index_512834[1:0]}) < $signed({1'h0, sel_527737}) ? {add_527735, array_index_512834[1:0]} : sel_527737;
  assign add_528445 = array_index_512883[11:2] + 10'h113;
  assign sel_528447 = $signed({1'h0, add_527739, array_index_512837[1:0]}) < $signed({1'h0, sel_527741}) ? {add_527739, array_index_512837[1:0]} : sel_527741;
  assign add_528459 = array_index_513022[11:4] + 8'h49;
  assign sel_528461 = $signed({1'h0, add_527753, array_index_512942[3:0]}) < $signed({1'h0, sel_527755}) ? {add_527753, array_index_512942[3:0]} : sel_527755;
  assign add_528463 = array_index_513025[11:4] + 8'h49;
  assign sel_528465 = $signed({1'h0, add_527757, array_index_512945[3:0]}) < $signed({1'h0, sel_527759}) ? {add_527757, array_index_512945[3:0]} : sel_527759;
  assign add_528475 = array_index_513238[11:0] + 12'h263;
  assign sel_528477 = $signed({1'h0, add_527769}) < $signed({1'h0, sel_527771}) ? add_527769 : sel_527771;
  assign add_528479 = array_index_513241[11:0] + 12'h263;
  assign sel_528481 = $signed({1'h0, add_527773}) < $signed({1'h0, sel_527775}) ? add_527773 : sel_527775;
  assign add_528491 = array_index_513530[11:1] + 11'h109;
  assign sel_528493 = $signed({1'h0, add_527785, array_index_513374[0]}) < $signed({1'h0, sel_527787}) ? {add_527785, array_index_513374[0]} : sel_527787;
  assign add_528495 = array_index_513533[11:1] + 11'h109;
  assign sel_528497 = $signed({1'h0, add_527789, array_index_513377[0]}) < $signed({1'h0, sel_527791}) ? {add_527789, array_index_513377[0]} : sel_527791;
  assign add_528507 = array_index_513890[11:3] + 9'h12f;
  assign sel_528509 = $signed({1'h0, add_527801, array_index_513702[2:0]}) < $signed({1'h0, sel_527803}) ? {add_527801, array_index_513702[2:0]} : sel_527803;
  assign add_528511 = array_index_513893[11:3] + 9'h12f;
  assign sel_528513 = $signed({1'h0, add_527805, array_index_513705[2:0]}) < $signed({1'h0, sel_527807}) ? {add_527805, array_index_513705[2:0]} : sel_527807;
  assign add_528525 = array_index_514318[11:3] + 9'h171;
  assign sel_528527 = $signed({1'h0, add_527819, array_index_514096[2:0]}) < $signed({1'h0, sel_527821}) ? {add_527819, array_index_514096[2:0]} : sel_527821;
  assign add_528529 = array_index_514321[11:3] + 9'h171;
  assign sel_528531 = $signed({1'h0, add_527823, array_index_514099[2:0]}) < $signed({1'h0, sel_527825}) ? {add_527823, array_index_514099[2:0]} : sel_527825;
  assign add_528541 = array_index_514818[11:0] + 12'h091;
  assign sel_528543 = $signed({1'h0, add_527835}) < $signed({1'h0, sel_527837}) ? add_527835 : sel_527837;
  assign add_528545 = array_index_514821[11:0] + 12'h091;
  assign sel_528547 = $signed({1'h0, add_527839}) < $signed({1'h0, sel_527841}) ? add_527839 : sel_527841;
  assign add_528557 = array_index_515398[11:0] + 12'hf59;
  assign sel_528559 = $signed({1'h0, add_527851}) < $signed({1'h0, sel_527853}) ? add_527851 : sel_527853;
  assign add_528561 = array_index_515401[11:0] + 12'hf59;
  assign sel_528563 = $signed({1'h0, add_527855}) < $signed({1'h0, sel_527857}) ? add_527855 : sel_527857;
  assign add_528575 = array_index_516080[11:0] + 12'h437;
  assign sel_528577 = $signed({1'h0, add_527869}) < $signed({1'h0, sel_527871}) ? add_527869 : sel_527871;
  assign add_528579 = array_index_516083[11:0] + 12'h437;
  assign sel_528581 = $signed({1'h0, add_527873}) < $signed({1'h0, sel_527875}) ? add_527873 : sel_527875;
  assign add_528591 = array_index_516860[11:0] + 12'hee1;
  assign sel_528593 = $signed({1'h0, add_527885}) < $signed({1'h0, sel_527887}) ? add_527885 : sel_527887;
  assign add_528595 = array_index_516863[11:0] + 12'hee1;
  assign sel_528597 = $signed({1'h0, add_527889}) < $signed({1'h0, sel_527891}) ? add_527889 : sel_527891;
  assign add_528607 = array_index_517736[11:1] + 11'h179;
  assign sel_528609 = $signed({1'h0, add_527901, array_index_517286[0]}) < $signed({1'h0, sel_527903}) ? {add_527901, array_index_517286[0]} : sel_527903;
  assign add_528611 = array_index_517739[11:1] + 11'h179;
  assign sel_528613 = $signed({1'h0, add_527905, array_index_517289[0]}) < $signed({1'h0, sel_527907}) ? {add_527905, array_index_517289[0]} : sel_527907;
  assign add_528623 = array_index_518710[11:0] + 12'h067;
  assign sel_528625 = $signed({1'h0, add_527917}) < $signed({1'h0, sel_527919}) ? add_527917 : sel_527919;
  assign add_528627 = array_index_518713[11:0] + 12'h067;
  assign sel_528629 = $signed({1'h0, add_527921}) < $signed({1'h0, sel_527923}) ? add_527921 : sel_527923;
  assign add_528631 = array_index_519236[11:3] + 9'h1ef;
  assign sel_528634 = $signed({1'h0, add_527925, array_index_518710[2:0]}) < $signed({1'h0, sel_527928}) ? {add_527925, array_index_518710[2:0]} : sel_527928;
  assign add_528636 = array_index_519239[11:3] + 9'h1ef;
  assign sel_528639 = $signed({1'h0, add_527930, array_index_518713[2:0]}) < $signed({1'h0, sel_527933}) ? {add_527930, array_index_518713[2:0]} : sel_527933;
  assign add_528641 = array_index_519786[11:1] + 11'h2d5;
  assign sel_528643 = $signed({1'h0, add_527935, array_index_519236[0]}) < $signed({1'h0, sel_527937}) ? {add_527935, array_index_519236[0]} : sel_527937;
  assign add_528645 = array_index_519789[11:1] + 11'h2d5;
  assign sel_528647 = $signed({1'h0, add_527939, array_index_519239[0]}) < $signed({1'h0, sel_527941}) ? {add_527939, array_index_519239[0]} : sel_527941;
  assign add_528649 = array_index_520362[11:2] + 10'h353;
  assign sel_528651 = $signed({1'h0, add_527943, array_index_519786[1:0]}) < $signed({1'h0, sel_527945}) ? {add_527943, array_index_519786[1:0]} : sel_527945;
  assign add_528653 = array_index_520365[11:2] + 10'h353;
  assign sel_528655 = $signed({1'h0, add_527947, array_index_519789[1:0]}) < $signed({1'h0, sel_527949}) ? {add_527947, array_index_519789[1:0]} : sel_527949;
  assign add_528657 = array_index_520964[11:0] + 12'h0a7;
  assign sel_528659 = $signed({1'h0, add_527951}) < $signed({1'h0, sel_527953}) ? add_527951 : sel_527953;
  assign add_528661 = array_index_520967[11:0] + 12'h0a7;
  assign sel_528663 = $signed({1'h0, add_527955}) < $signed({1'h0, sel_527957}) ? add_527955 : sel_527957;
  assign add_528665 = array_index_521590[11:1] + 11'h4cb;
  assign sel_528667 = $signed({1'h0, add_527959, array_index_520964[0]}) < $signed({1'h0, sel_527961}) ? {add_527959, array_index_520964[0]} : sel_527961;
  assign add_528669 = array_index_521593[11:1] + 11'h4cb;
  assign sel_528671 = $signed({1'h0, add_527963, array_index_520967[0]}) < $signed({1'h0, sel_527965}) ? {add_527963, array_index_520967[0]} : sel_527965;
  assign concat_528674 = {1'h0, ($signed({1'h0, add_527259}) < $signed({1'h0, sel_527261}) ? add_527259 : sel_527261) == ($signed({1'h0, add_527263}) < $signed({1'h0, sel_527265}) ? add_527263 : sel_527265) ? add_528201 : concat_527976};
  assign add_528685 = array_index_512942[11:1] + 11'h5b9;
  assign sel_528687 = $signed({1'h0, add_527989, array_index_512880[0]}) < $signed({1'h0, sel_527991}) ? {add_527989, array_index_512880[0]} : sel_527991;
  assign add_528689 = array_index_512945[11:1] + 11'h5b9;
  assign sel_528691 = $signed({1'h0, add_527993, array_index_512883[0]}) < $signed({1'h0, sel_527995}) ? {add_527993, array_index_512883[0]} : sel_527995;
  assign add_528701 = array_index_513120[11:0] + 12'h37b;
  assign sel_528703 = $signed({1'h0, add_528005}) < $signed({1'h0, sel_528007}) ? add_528005 : sel_528007;
  assign add_528705 = array_index_513123[11:0] + 12'h37b;
  assign sel_528707 = $signed({1'h0, add_528009}) < $signed({1'h0, sel_528011}) ? add_528009 : sel_528011;
  assign add_528719 = array_index_513374[11:0] + 12'h811;
  assign sel_528721 = $signed({1'h0, add_528023}) < $signed({1'h0, sel_528025}) ? add_528023 : sel_528025;
  assign add_528723 = array_index_513377[11:0] + 12'h811;
  assign sel_528725 = $signed({1'h0, add_528027}) < $signed({1'h0, sel_528029}) ? add_528027 : sel_528029;
  assign add_528737 = array_index_513702[11:0] + 12'h70f;
  assign sel_528739 = $signed({1'h0, add_528041}) < $signed({1'h0, sel_528043}) ? add_528041 : sel_528043;
  assign add_528741 = array_index_513705[11:0] + 12'h70f;
  assign sel_528743 = $signed({1'h0, add_528045}) < $signed({1'h0, sel_528047}) ? add_528045 : sel_528047;
  assign add_528755 = array_index_514096[11:3] + 9'h1f1;
  assign sel_528757 = $signed({1'h0, add_528059, array_index_513890[2:0]}) < $signed({1'h0, sel_528061}) ? {add_528059, array_index_513890[2:0]} : sel_528061;
  assign add_528759 = array_index_514099[11:3] + 9'h1f1;
  assign sel_528761 = $signed({1'h0, add_528063, array_index_513893[2:0]}) < $signed({1'h0, sel_528065}) ? {add_528063, array_index_513893[2:0]} : sel_528065;
  assign add_528771 = array_index_514558[11:0] + 12'h081;
  assign sel_528773 = $signed({1'h0, add_528075}) < $signed({1'h0, sel_528077}) ? add_528075 : sel_528077;
  assign add_528775 = array_index_514561[11:0] + 12'h081;
  assign sel_528777 = $signed({1'h0, add_528079}) < $signed({1'h0, sel_528081}) ? add_528079 : sel_528081;
  assign add_528789 = array_index_515098[11:0] + 12'h0b1;
  assign sel_528791 = $signed({1'h0, add_528093}) < $signed({1'h0, sel_528095}) ? add_528093 : sel_528095;
  assign add_528793 = array_index_515101[11:0] + 12'h0b1;
  assign sel_528795 = $signed({1'h0, add_528097}) < $signed({1'h0, sel_528099}) ? add_528097 : sel_528099;
  assign add_528807 = array_index_515726[11:1] + 11'h4c1;
  assign sel_528809 = $signed({1'h0, add_528111, array_index_515398[0]}) < $signed({1'h0, sel_528113}) ? {add_528111, array_index_515398[0]} : sel_528113;
  assign add_528811 = array_index_515729[11:1] + 11'h4c1;
  assign sel_528813 = $signed({1'h0, add_528115, array_index_515401[0]}) < $signed({1'h0, sel_528117}) ? {add_528115, array_index_515401[0]} : sel_528117;
  assign add_528823 = array_index_516458[11:0] + 12'hbb1;
  assign sel_528825 = $signed({1'h0, add_528127}) < $signed({1'h0, sel_528129}) ? add_528127 : sel_528129;
  assign add_528827 = array_index_516461[11:0] + 12'hbb1;
  assign sel_528829 = $signed({1'h0, add_528131}) < $signed({1'h0, sel_528133}) ? add_528131 : sel_528133;
  assign add_528839 = array_index_517286[11:0] + 12'h6ab;
  assign sel_528841 = $signed({1'h0, add_528143}) < $signed({1'h0, sel_528145}) ? add_528143 : sel_528145;
  assign add_528843 = array_index_517289[11:0] + 12'h6ab;
  assign sel_528845 = $signed({1'h0, add_528147}) < $signed({1'h0, sel_528149}) ? add_528147 : sel_528149;
  assign add_528855 = array_index_518210[11:0] + 12'h7d5;
  assign sel_528857 = $signed({1'h0, add_528159}) < $signed({1'h0, sel_528161}) ? add_528159 : sel_528161;
  assign add_528859 = array_index_518213[11:0] + 12'h7d5;
  assign sel_528861 = $signed({1'h0, add_528163}) < $signed({1'h0, sel_528165}) ? add_528163 : sel_528165;
  assign add_528893 = concat_528674 + 10'h001;
  assign add_528895 = array_index_512880[11:0] + 12'hcc1;
  assign sel_528897 = $signed({1'h0, add_528203}) < $signed({1'h0, sel_528205}) ? add_528203 : sel_528205;
  assign add_528899 = array_index_512883[11:0] + 12'hcc1;
  assign sel_528901 = $signed({1'h0, add_528207}) < $signed({1'h0, sel_528209}) ? add_528207 : sel_528209;
  assign add_528913 = array_index_513022[11:0] + 12'ha87;
  assign sel_528915 = $signed({1'h0, add_528221}) < $signed({1'h0, sel_528223}) ? add_528221 : sel_528223;
  assign add_528917 = array_index_513025[11:0] + 12'ha87;
  assign sel_528919 = $signed({1'h0, add_528225}) < $signed({1'h0, sel_528227}) ? add_528225 : sel_528227;
  assign add_528931 = array_index_513238[11:1] + 11'h663;
  assign sel_528933 = $signed({1'h0, add_528239, array_index_513120[0]}) < $signed({1'h0, sel_528241}) ? {add_528239, array_index_513120[0]} : sel_528241;
  assign add_528935 = array_index_513241[11:1] + 11'h663;
  assign sel_528937 = $signed({1'h0, add_528243, array_index_513123[0]}) < $signed({1'h0, sel_528245}) ? {add_528243, array_index_513123[0]} : sel_528245;
  assign add_528947 = array_index_513530[11:1] + 11'h075;
  assign sel_528949 = $signed({1'h0, add_528255, array_index_513374[0]}) < $signed({1'h0, sel_528257}) ? {add_528255, array_index_513374[0]} : sel_528257;
  assign add_528951 = array_index_513533[11:1] + 11'h075;
  assign sel_528953 = $signed({1'h0, add_528259, array_index_513377[0]}) < $signed({1'h0, sel_528261}) ? {add_528259, array_index_513377[0]} : sel_528261;
  assign add_528965 = array_index_513890[11:2] + 10'h181;
  assign sel_528967 = $signed({1'h0, add_528273, array_index_513702[1:0]}) < $signed({1'h0, sel_528275}) ? {add_528273, array_index_513702[1:0]} : sel_528275;
  assign add_528969 = array_index_513893[11:2] + 10'h181;
  assign sel_528971 = $signed({1'h0, add_528277, array_index_513705[1:0]}) < $signed({1'h0, sel_528279}) ? {add_528277, array_index_513705[1:0]} : sel_528279;
  assign add_528983 = array_index_514318[11:0] + 12'h8a7;
  assign sel_528985 = $signed({1'h0, add_528291}) < $signed({1'h0, sel_528293}) ? add_528291 : sel_528293;
  assign add_528987 = array_index_514321[11:0] + 12'h8a7;
  assign sel_528989 = $signed({1'h0, add_528295}) < $signed({1'h0, sel_528297}) ? add_528295 : sel_528297;
  assign add_529001 = array_index_514818[11:1] + 11'h283;
  assign sel_529003 = $signed({1'h0, add_528309, array_index_514558[0]}) < $signed({1'h0, sel_528311}) ? {add_528309, array_index_514558[0]} : sel_528311;
  assign add_529005 = array_index_514821[11:1] + 11'h283;
  assign sel_529007 = $signed({1'h0, add_528313, array_index_514561[0]}) < $signed({1'h0, sel_528315}) ? {add_528313, array_index_514561[0]} : sel_528315;
  assign add_529017 = array_index_515398[11:1] + 11'h44d;
  assign sel_529019 = $signed({1'h0, add_528325, array_index_515098[0]}) < $signed({1'h0, sel_528327}) ? {add_528325, array_index_515098[0]} : sel_528327;
  assign add_529021 = array_index_515401[11:1] + 11'h44d;
  assign sel_529023 = $signed({1'h0, add_528329, array_index_515101[0]}) < $signed({1'h0, sel_528331}) ? {add_528329, array_index_515101[0]} : sel_528331;
  assign add_529033 = array_index_516080[11:0] + 12'hcb1;
  assign sel_529035 = $signed({1'h0, add_528341}) < $signed({1'h0, sel_528343}) ? add_528341 : sel_528343;
  assign add_529037 = array_index_516083[11:0] + 12'hcb1;
  assign sel_529039 = $signed({1'h0, add_528345}) < $signed({1'h0, sel_528347}) ? add_528345 : sel_528347;
  assign add_529049 = array_index_516860[11:0] + 12'h81f;
  assign sel_529051 = $signed({1'h0, add_528357}) < $signed({1'h0, sel_528359}) ? add_528357 : sel_528359;
  assign add_529053 = array_index_516863[11:0] + 12'h81f;
  assign sel_529055 = $signed({1'h0, add_528361}) < $signed({1'h0, sel_528363}) ? add_528361 : sel_528363;
  assign add_529065 = array_index_517736[11:0] + 12'h45b;
  assign sel_529067 = $signed({1'h0, add_528373}) < $signed({1'h0, sel_528375}) ? add_528373 : sel_528375;
  assign add_529069 = array_index_517739[11:0] + 12'h45b;
  assign sel_529071 = $signed({1'h0, add_528377}) < $signed({1'h0, sel_528379}) ? add_528377 : sel_528379;
  assign add_529083 = array_index_518710[11:3] + 9'h0f5;
  assign sel_529085 = $signed({1'h0, add_528391, array_index_518210[2:0]}) < $signed({1'h0, sel_528393}) ? {add_528391, array_index_518210[2:0]} : sel_528393;
  assign add_529087 = array_index_518713[11:3] + 9'h0f5;
  assign sel_529089 = $signed({1'h0, add_528395, array_index_518213[2:0]}) < $signed({1'h0, sel_528397}) ? {add_528395, array_index_518213[2:0]} : sel_528397;
  assign add_529129 = array_index_512942[11:2] + 10'h113;
  assign sel_529131 = $signed({1'h0, add_528441, array_index_512880[1:0]}) < $signed({1'h0, sel_528443}) ? {add_528441, array_index_512880[1:0]} : sel_528443;
  assign add_529133 = array_index_512945[11:2] + 10'h113;
  assign sel_529135 = $signed({1'h0, add_528445, array_index_512883[1:0]}) < $signed({1'h0, sel_528447}) ? {add_528445, array_index_512883[1:0]} : sel_528447;
  assign add_529147 = array_index_513120[11:4] + 8'h49;
  assign sel_529149 = $signed({1'h0, add_528459, array_index_513022[3:0]}) < $signed({1'h0, sel_528461}) ? {add_528459, array_index_513022[3:0]} : sel_528461;
  assign add_529151 = array_index_513123[11:4] + 8'h49;
  assign sel_529153 = $signed({1'h0, add_528463, array_index_513025[3:0]}) < $signed({1'h0, sel_528465}) ? {add_528463, array_index_513025[3:0]} : sel_528465;
  assign add_529163 = array_index_513374[11:0] + 12'h263;
  assign sel_529165 = $signed({1'h0, add_528475}) < $signed({1'h0, sel_528477}) ? add_528475 : sel_528477;
  assign add_529167 = array_index_513377[11:0] + 12'h263;
  assign sel_529169 = $signed({1'h0, add_528479}) < $signed({1'h0, sel_528481}) ? add_528479 : sel_528481;
  assign add_529179 = array_index_513702[11:1] + 11'h109;
  assign sel_529181 = $signed({1'h0, add_528491, array_index_513530[0]}) < $signed({1'h0, sel_528493}) ? {add_528491, array_index_513530[0]} : sel_528493;
  assign add_529183 = array_index_513705[11:1] + 11'h109;
  assign sel_529185 = $signed({1'h0, add_528495, array_index_513533[0]}) < $signed({1'h0, sel_528497}) ? {add_528495, array_index_513533[0]} : sel_528497;
  assign add_529195 = array_index_514096[11:3] + 9'h12f;
  assign sel_529197 = $signed({1'h0, add_528507, array_index_513890[2:0]}) < $signed({1'h0, sel_528509}) ? {add_528507, array_index_513890[2:0]} : sel_528509;
  assign add_529199 = array_index_514099[11:3] + 9'h12f;
  assign sel_529201 = $signed({1'h0, add_528511, array_index_513893[2:0]}) < $signed({1'h0, sel_528513}) ? {add_528511, array_index_513893[2:0]} : sel_528513;
  assign add_529213 = array_index_514558[11:3] + 9'h171;
  assign sel_529215 = $signed({1'h0, add_528525, array_index_514318[2:0]}) < $signed({1'h0, sel_528527}) ? {add_528525, array_index_514318[2:0]} : sel_528527;
  assign add_529217 = array_index_514561[11:3] + 9'h171;
  assign sel_529219 = $signed({1'h0, add_528529, array_index_514321[2:0]}) < $signed({1'h0, sel_528531}) ? {add_528529, array_index_514321[2:0]} : sel_528531;
  assign add_529229 = array_index_515098[11:0] + 12'h091;
  assign sel_529231 = $signed({1'h0, add_528541}) < $signed({1'h0, sel_528543}) ? add_528541 : sel_528543;
  assign add_529233 = array_index_515101[11:0] + 12'h091;
  assign sel_529235 = $signed({1'h0, add_528545}) < $signed({1'h0, sel_528547}) ? add_528545 : sel_528547;
  assign add_529245 = array_index_515726[11:0] + 12'hf59;
  assign sel_529247 = $signed({1'h0, add_528557}) < $signed({1'h0, sel_528559}) ? add_528557 : sel_528559;
  assign add_529249 = array_index_515729[11:0] + 12'hf59;
  assign sel_529251 = $signed({1'h0, add_528561}) < $signed({1'h0, sel_528563}) ? add_528561 : sel_528563;
  assign add_529263 = array_index_516458[11:0] + 12'h437;
  assign sel_529265 = $signed({1'h0, add_528575}) < $signed({1'h0, sel_528577}) ? add_528575 : sel_528577;
  assign add_529267 = array_index_516461[11:0] + 12'h437;
  assign sel_529269 = $signed({1'h0, add_528579}) < $signed({1'h0, sel_528581}) ? add_528579 : sel_528581;
  assign add_529279 = array_index_517286[11:0] + 12'hee1;
  assign sel_529281 = $signed({1'h0, add_528591}) < $signed({1'h0, sel_528593}) ? add_528591 : sel_528593;
  assign add_529283 = array_index_517289[11:0] + 12'hee1;
  assign sel_529285 = $signed({1'h0, add_528595}) < $signed({1'h0, sel_528597}) ? add_528595 : sel_528597;
  assign add_529295 = array_index_518210[11:1] + 11'h179;
  assign sel_529297 = $signed({1'h0, add_528607, array_index_517736[0]}) < $signed({1'h0, sel_528609}) ? {add_528607, array_index_517736[0]} : sel_528609;
  assign add_529299 = array_index_518213[11:1] + 11'h179;
  assign sel_529301 = $signed({1'h0, add_528611, array_index_517739[0]}) < $signed({1'h0, sel_528613}) ? {add_528611, array_index_517739[0]} : sel_528613;
  assign add_529311 = array_index_519236[11:0] + 12'h067;
  assign sel_529313 = $signed({1'h0, add_528623}) < $signed({1'h0, sel_528625}) ? add_528623 : sel_528625;
  assign add_529315 = array_index_519239[11:0] + 12'h067;
  assign sel_529317 = $signed({1'h0, add_528627}) < $signed({1'h0, sel_528629}) ? add_528627 : sel_528629;
  assign add_529319 = array_index_519786[11:3] + 9'h1ef;
  assign sel_529322 = $signed({1'h0, add_528631, array_index_519236[2:0]}) < $signed({1'h0, sel_528634}) ? {add_528631, array_index_519236[2:0]} : sel_528634;
  assign add_529324 = array_index_519789[11:3] + 9'h1ef;
  assign sel_529327 = $signed({1'h0, add_528636, array_index_519239[2:0]}) < $signed({1'h0, sel_528639}) ? {add_528636, array_index_519239[2:0]} : sel_528639;
  assign add_529329 = array_index_520362[11:1] + 11'h2d5;
  assign sel_529331 = $signed({1'h0, add_528641, array_index_519786[0]}) < $signed({1'h0, sel_528643}) ? {add_528641, array_index_519786[0]} : sel_528643;
  assign add_529333 = array_index_520365[11:1] + 11'h2d5;
  assign sel_529335 = $signed({1'h0, add_528645, array_index_519789[0]}) < $signed({1'h0, sel_528647}) ? {add_528645, array_index_519789[0]} : sel_528647;
  assign add_529337 = array_index_520964[11:2] + 10'h353;
  assign sel_529339 = $signed({1'h0, add_528649, array_index_520362[1:0]}) < $signed({1'h0, sel_528651}) ? {add_528649, array_index_520362[1:0]} : sel_528651;
  assign add_529341 = array_index_520967[11:2] + 10'h353;
  assign sel_529343 = $signed({1'h0, add_528653, array_index_520365[1:0]}) < $signed({1'h0, sel_528655}) ? {add_528653, array_index_520365[1:0]} : sel_528655;
  assign add_529345 = array_index_521590[11:0] + 12'h0a7;
  assign sel_529347 = $signed({1'h0, add_528657}) < $signed({1'h0, sel_528659}) ? add_528657 : sel_528659;
  assign add_529349 = array_index_521593[11:0] + 12'h0a7;
  assign sel_529351 = $signed({1'h0, add_528661}) < $signed({1'h0, sel_528663}) ? add_528661 : sel_528663;
  assign concat_529354 = {1'h0, ($signed({1'h0, add_527967}) < $signed({1'h0, sel_527969}) ? add_527967 : sel_527969) == ($signed({1'h0, add_527971}) < $signed({1'h0, sel_527973}) ? add_527971 : sel_527973) ? add_528893 : concat_528674};
  assign add_529365 = array_index_513022[11:1] + 11'h5b9;
  assign sel_529367 = $signed({1'h0, add_528685, array_index_512942[0]}) < $signed({1'h0, sel_528687}) ? {add_528685, array_index_512942[0]} : sel_528687;
  assign add_529369 = array_index_513025[11:1] + 11'h5b9;
  assign sel_529371 = $signed({1'h0, add_528689, array_index_512945[0]}) < $signed({1'h0, sel_528691}) ? {add_528689, array_index_512945[0]} : sel_528691;
  assign add_529381 = array_index_513238[11:0] + 12'h37b;
  assign sel_529383 = $signed({1'h0, add_528701}) < $signed({1'h0, sel_528703}) ? add_528701 : sel_528703;
  assign add_529385 = array_index_513241[11:0] + 12'h37b;
  assign sel_529387 = $signed({1'h0, add_528705}) < $signed({1'h0, sel_528707}) ? add_528705 : sel_528707;
  assign add_529399 = array_index_513530[11:0] + 12'h811;
  assign sel_529401 = $signed({1'h0, add_528719}) < $signed({1'h0, sel_528721}) ? add_528719 : sel_528721;
  assign add_529403 = array_index_513533[11:0] + 12'h811;
  assign sel_529405 = $signed({1'h0, add_528723}) < $signed({1'h0, sel_528725}) ? add_528723 : sel_528725;
  assign add_529417 = array_index_513890[11:0] + 12'h70f;
  assign sel_529419 = $signed({1'h0, add_528737}) < $signed({1'h0, sel_528739}) ? add_528737 : sel_528739;
  assign add_529421 = array_index_513893[11:0] + 12'h70f;
  assign sel_529423 = $signed({1'h0, add_528741}) < $signed({1'h0, sel_528743}) ? add_528741 : sel_528743;
  assign add_529435 = array_index_514318[11:3] + 9'h1f1;
  assign sel_529437 = $signed({1'h0, add_528755, array_index_514096[2:0]}) < $signed({1'h0, sel_528757}) ? {add_528755, array_index_514096[2:0]} : sel_528757;
  assign add_529439 = array_index_514321[11:3] + 9'h1f1;
  assign sel_529441 = $signed({1'h0, add_528759, array_index_514099[2:0]}) < $signed({1'h0, sel_528761}) ? {add_528759, array_index_514099[2:0]} : sel_528761;
  assign add_529451 = array_index_514818[11:0] + 12'h081;
  assign sel_529453 = $signed({1'h0, add_528771}) < $signed({1'h0, sel_528773}) ? add_528771 : sel_528773;
  assign add_529455 = array_index_514821[11:0] + 12'h081;
  assign sel_529457 = $signed({1'h0, add_528775}) < $signed({1'h0, sel_528777}) ? add_528775 : sel_528777;
  assign add_529469 = array_index_515398[11:0] + 12'h0b1;
  assign sel_529471 = $signed({1'h0, add_528789}) < $signed({1'h0, sel_528791}) ? add_528789 : sel_528791;
  assign add_529473 = array_index_515401[11:0] + 12'h0b1;
  assign sel_529475 = $signed({1'h0, add_528793}) < $signed({1'h0, sel_528795}) ? add_528793 : sel_528795;
  assign add_529487 = array_index_516080[11:1] + 11'h4c1;
  assign sel_529489 = $signed({1'h0, add_528807, array_index_515726[0]}) < $signed({1'h0, sel_528809}) ? {add_528807, array_index_515726[0]} : sel_528809;
  assign add_529491 = array_index_516083[11:1] + 11'h4c1;
  assign sel_529493 = $signed({1'h0, add_528811, array_index_515729[0]}) < $signed({1'h0, sel_528813}) ? {add_528811, array_index_515729[0]} : sel_528813;
  assign add_529503 = array_index_516860[11:0] + 12'hbb1;
  assign sel_529505 = $signed({1'h0, add_528823}) < $signed({1'h0, sel_528825}) ? add_528823 : sel_528825;
  assign add_529507 = array_index_516863[11:0] + 12'hbb1;
  assign sel_529509 = $signed({1'h0, add_528827}) < $signed({1'h0, sel_528829}) ? add_528827 : sel_528829;
  assign add_529519 = array_index_517736[11:0] + 12'h6ab;
  assign sel_529521 = $signed({1'h0, add_528839}) < $signed({1'h0, sel_528841}) ? add_528839 : sel_528841;
  assign add_529523 = array_index_517739[11:0] + 12'h6ab;
  assign sel_529525 = $signed({1'h0, add_528843}) < $signed({1'h0, sel_528845}) ? add_528843 : sel_528845;
  assign add_529535 = array_index_518710[11:0] + 12'h7d5;
  assign sel_529537 = $signed({1'h0, add_528855}) < $signed({1'h0, sel_528857}) ? add_528855 : sel_528857;
  assign add_529539 = array_index_518713[11:0] + 12'h7d5;
  assign sel_529541 = $signed({1'h0, add_528859}) < $signed({1'h0, sel_528861}) ? add_528859 : sel_528861;
  assign add_529569 = concat_529354 + 11'h001;
  assign add_529571 = array_index_512942[11:0] + 12'hcc1;
  assign sel_529573 = $signed({1'h0, add_528895}) < $signed({1'h0, sel_528897}) ? add_528895 : sel_528897;
  assign add_529575 = array_index_512945[11:0] + 12'hcc1;
  assign sel_529577 = $signed({1'h0, add_528899}) < $signed({1'h0, sel_528901}) ? add_528899 : sel_528901;
  assign add_529589 = array_index_513120[11:0] + 12'ha87;
  assign sel_529591 = $signed({1'h0, add_528913}) < $signed({1'h0, sel_528915}) ? add_528913 : sel_528915;
  assign add_529593 = array_index_513123[11:0] + 12'ha87;
  assign sel_529595 = $signed({1'h0, add_528917}) < $signed({1'h0, sel_528919}) ? add_528917 : sel_528919;
  assign add_529607 = array_index_513374[11:1] + 11'h663;
  assign sel_529609 = $signed({1'h0, add_528931, array_index_513238[0]}) < $signed({1'h0, sel_528933}) ? {add_528931, array_index_513238[0]} : sel_528933;
  assign add_529611 = array_index_513377[11:1] + 11'h663;
  assign sel_529613 = $signed({1'h0, add_528935, array_index_513241[0]}) < $signed({1'h0, sel_528937}) ? {add_528935, array_index_513241[0]} : sel_528937;
  assign add_529623 = array_index_513702[11:1] + 11'h075;
  assign sel_529625 = $signed({1'h0, add_528947, array_index_513530[0]}) < $signed({1'h0, sel_528949}) ? {add_528947, array_index_513530[0]} : sel_528949;
  assign add_529627 = array_index_513705[11:1] + 11'h075;
  assign sel_529629 = $signed({1'h0, add_528951, array_index_513533[0]}) < $signed({1'h0, sel_528953}) ? {add_528951, array_index_513533[0]} : sel_528953;
  assign add_529641 = array_index_514096[11:2] + 10'h181;
  assign sel_529643 = $signed({1'h0, add_528965, array_index_513890[1:0]}) < $signed({1'h0, sel_528967}) ? {add_528965, array_index_513890[1:0]} : sel_528967;
  assign add_529645 = array_index_514099[11:2] + 10'h181;
  assign sel_529647 = $signed({1'h0, add_528969, array_index_513893[1:0]}) < $signed({1'h0, sel_528971}) ? {add_528969, array_index_513893[1:0]} : sel_528971;
  assign add_529659 = array_index_514558[11:0] + 12'h8a7;
  assign sel_529661 = $signed({1'h0, add_528983}) < $signed({1'h0, sel_528985}) ? add_528983 : sel_528985;
  assign add_529663 = array_index_514561[11:0] + 12'h8a7;
  assign sel_529665 = $signed({1'h0, add_528987}) < $signed({1'h0, sel_528989}) ? add_528987 : sel_528989;
  assign add_529677 = array_index_515098[11:1] + 11'h283;
  assign sel_529679 = $signed({1'h0, add_529001, array_index_514818[0]}) < $signed({1'h0, sel_529003}) ? {add_529001, array_index_514818[0]} : sel_529003;
  assign add_529681 = array_index_515101[11:1] + 11'h283;
  assign sel_529683 = $signed({1'h0, add_529005, array_index_514821[0]}) < $signed({1'h0, sel_529007}) ? {add_529005, array_index_514821[0]} : sel_529007;
  assign add_529693 = array_index_515726[11:1] + 11'h44d;
  assign sel_529695 = $signed({1'h0, add_529017, array_index_515398[0]}) < $signed({1'h0, sel_529019}) ? {add_529017, array_index_515398[0]} : sel_529019;
  assign add_529697 = array_index_515729[11:1] + 11'h44d;
  assign sel_529699 = $signed({1'h0, add_529021, array_index_515401[0]}) < $signed({1'h0, sel_529023}) ? {add_529021, array_index_515401[0]} : sel_529023;
  assign add_529709 = array_index_516458[11:0] + 12'hcb1;
  assign sel_529711 = $signed({1'h0, add_529033}) < $signed({1'h0, sel_529035}) ? add_529033 : sel_529035;
  assign add_529713 = array_index_516461[11:0] + 12'hcb1;
  assign sel_529715 = $signed({1'h0, add_529037}) < $signed({1'h0, sel_529039}) ? add_529037 : sel_529039;
  assign add_529725 = array_index_517286[11:0] + 12'h81f;
  assign sel_529727 = $signed({1'h0, add_529049}) < $signed({1'h0, sel_529051}) ? add_529049 : sel_529051;
  assign add_529729 = array_index_517289[11:0] + 12'h81f;
  assign sel_529731 = $signed({1'h0, add_529053}) < $signed({1'h0, sel_529055}) ? add_529053 : sel_529055;
  assign add_529741 = array_index_518210[11:0] + 12'h45b;
  assign sel_529743 = $signed({1'h0, add_529065}) < $signed({1'h0, sel_529067}) ? add_529065 : sel_529067;
  assign add_529745 = array_index_518213[11:0] + 12'h45b;
  assign sel_529747 = $signed({1'h0, add_529069}) < $signed({1'h0, sel_529071}) ? add_529069 : sel_529071;
  assign add_529759 = array_index_519236[11:3] + 9'h0f5;
  assign sel_529761 = $signed({1'h0, add_529083, array_index_518710[2:0]}) < $signed({1'h0, sel_529085}) ? {add_529083, array_index_518710[2:0]} : sel_529085;
  assign add_529763 = array_index_519239[11:3] + 9'h0f5;
  assign sel_529765 = $signed({1'h0, add_529087, array_index_518713[2:0]}) < $signed({1'h0, sel_529089}) ? {add_529087, array_index_518713[2:0]} : sel_529089;
  assign add_529799 = array_index_513022[11:2] + 10'h113;
  assign sel_529801 = $signed({1'h0, add_529129, array_index_512942[1:0]}) < $signed({1'h0, sel_529131}) ? {add_529129, array_index_512942[1:0]} : sel_529131;
  assign add_529803 = array_index_513025[11:2] + 10'h113;
  assign sel_529805 = $signed({1'h0, add_529133, array_index_512945[1:0]}) < $signed({1'h0, sel_529135}) ? {add_529133, array_index_512945[1:0]} : sel_529135;
  assign add_529817 = array_index_513238[11:4] + 8'h49;
  assign sel_529819 = $signed({1'h0, add_529147, array_index_513120[3:0]}) < $signed({1'h0, sel_529149}) ? {add_529147, array_index_513120[3:0]} : sel_529149;
  assign add_529821 = array_index_513241[11:4] + 8'h49;
  assign sel_529823 = $signed({1'h0, add_529151, array_index_513123[3:0]}) < $signed({1'h0, sel_529153}) ? {add_529151, array_index_513123[3:0]} : sel_529153;
  assign add_529833 = array_index_513530[11:0] + 12'h263;
  assign sel_529835 = $signed({1'h0, add_529163}) < $signed({1'h0, sel_529165}) ? add_529163 : sel_529165;
  assign add_529837 = array_index_513533[11:0] + 12'h263;
  assign sel_529839 = $signed({1'h0, add_529167}) < $signed({1'h0, sel_529169}) ? add_529167 : sel_529169;
  assign add_529849 = array_index_513890[11:1] + 11'h109;
  assign sel_529851 = $signed({1'h0, add_529179, array_index_513702[0]}) < $signed({1'h0, sel_529181}) ? {add_529179, array_index_513702[0]} : sel_529181;
  assign add_529853 = array_index_513893[11:1] + 11'h109;
  assign sel_529855 = $signed({1'h0, add_529183, array_index_513705[0]}) < $signed({1'h0, sel_529185}) ? {add_529183, array_index_513705[0]} : sel_529185;
  assign add_529865 = array_index_514318[11:3] + 9'h12f;
  assign sel_529867 = $signed({1'h0, add_529195, array_index_514096[2:0]}) < $signed({1'h0, sel_529197}) ? {add_529195, array_index_514096[2:0]} : sel_529197;
  assign add_529869 = array_index_514321[11:3] + 9'h12f;
  assign sel_529871 = $signed({1'h0, add_529199, array_index_514099[2:0]}) < $signed({1'h0, sel_529201}) ? {add_529199, array_index_514099[2:0]} : sel_529201;
  assign add_529883 = array_index_514818[11:3] + 9'h171;
  assign sel_529885 = $signed({1'h0, add_529213, array_index_514558[2:0]}) < $signed({1'h0, sel_529215}) ? {add_529213, array_index_514558[2:0]} : sel_529215;
  assign add_529887 = array_index_514821[11:3] + 9'h171;
  assign sel_529889 = $signed({1'h0, add_529217, array_index_514561[2:0]}) < $signed({1'h0, sel_529219}) ? {add_529217, array_index_514561[2:0]} : sel_529219;
  assign add_529899 = array_index_515398[11:0] + 12'h091;
  assign sel_529901 = $signed({1'h0, add_529229}) < $signed({1'h0, sel_529231}) ? add_529229 : sel_529231;
  assign add_529903 = array_index_515401[11:0] + 12'h091;
  assign sel_529905 = $signed({1'h0, add_529233}) < $signed({1'h0, sel_529235}) ? add_529233 : sel_529235;
  assign add_529915 = array_index_516080[11:0] + 12'hf59;
  assign sel_529917 = $signed({1'h0, add_529245}) < $signed({1'h0, sel_529247}) ? add_529245 : sel_529247;
  assign add_529919 = array_index_516083[11:0] + 12'hf59;
  assign sel_529921 = $signed({1'h0, add_529249}) < $signed({1'h0, sel_529251}) ? add_529249 : sel_529251;
  assign add_529933 = array_index_516860[11:0] + 12'h437;
  assign sel_529935 = $signed({1'h0, add_529263}) < $signed({1'h0, sel_529265}) ? add_529263 : sel_529265;
  assign add_529937 = array_index_516863[11:0] + 12'h437;
  assign sel_529939 = $signed({1'h0, add_529267}) < $signed({1'h0, sel_529269}) ? add_529267 : sel_529269;
  assign add_529949 = array_index_517736[11:0] + 12'hee1;
  assign sel_529951 = $signed({1'h0, add_529279}) < $signed({1'h0, sel_529281}) ? add_529279 : sel_529281;
  assign add_529953 = array_index_517739[11:0] + 12'hee1;
  assign sel_529955 = $signed({1'h0, add_529283}) < $signed({1'h0, sel_529285}) ? add_529283 : sel_529285;
  assign add_529965 = array_index_518710[11:1] + 11'h179;
  assign sel_529967 = $signed({1'h0, add_529295, array_index_518210[0]}) < $signed({1'h0, sel_529297}) ? {add_529295, array_index_518210[0]} : sel_529297;
  assign add_529969 = array_index_518713[11:1] + 11'h179;
  assign sel_529971 = $signed({1'h0, add_529299, array_index_518213[0]}) < $signed({1'h0, sel_529301}) ? {add_529299, array_index_518213[0]} : sel_529301;
  assign add_529981 = array_index_519786[11:0] + 12'h067;
  assign sel_529983 = $signed({1'h0, add_529311}) < $signed({1'h0, sel_529313}) ? add_529311 : sel_529313;
  assign add_529985 = array_index_519789[11:0] + 12'h067;
  assign sel_529987 = $signed({1'h0, add_529315}) < $signed({1'h0, sel_529317}) ? add_529315 : sel_529317;
  assign add_529989 = array_index_520362[11:3] + 9'h1ef;
  assign sel_529992 = $signed({1'h0, add_529319, array_index_519786[2:0]}) < $signed({1'h0, sel_529322}) ? {add_529319, array_index_519786[2:0]} : sel_529322;
  assign add_529994 = array_index_520365[11:3] + 9'h1ef;
  assign sel_529997 = $signed({1'h0, add_529324, array_index_519789[2:0]}) < $signed({1'h0, sel_529327}) ? {add_529324, array_index_519789[2:0]} : sel_529327;
  assign add_529999 = array_index_520964[11:1] + 11'h2d5;
  assign sel_530001 = $signed({1'h0, add_529329, array_index_520362[0]}) < $signed({1'h0, sel_529331}) ? {add_529329, array_index_520362[0]} : sel_529331;
  assign add_530003 = array_index_520967[11:1] + 11'h2d5;
  assign sel_530005 = $signed({1'h0, add_529333, array_index_520365[0]}) < $signed({1'h0, sel_529335}) ? {add_529333, array_index_520365[0]} : sel_529335;
  assign add_530007 = array_index_521590[11:2] + 10'h353;
  assign sel_530009 = $signed({1'h0, add_529337, array_index_520964[1:0]}) < $signed({1'h0, sel_529339}) ? {add_529337, array_index_520964[1:0]} : sel_529339;
  assign add_530011 = array_index_521593[11:2] + 10'h353;
  assign sel_530013 = $signed({1'h0, add_529341, array_index_520967[1:0]}) < $signed({1'h0, sel_529343}) ? {add_529341, array_index_520967[1:0]} : sel_529343;
  assign concat_530016 = {1'h0, ($signed({1'h0, add_528665, array_index_521590[0]}) < $signed({1'h0, sel_528667}) ? {add_528665, array_index_521590[0]} : sel_528667) == ($signed({1'h0, add_528669, array_index_521593[0]}) < $signed({1'h0, sel_528671}) ? {add_528669, array_index_521593[0]} : sel_528671) ? add_529569 : concat_529354};
  assign add_530027 = array_index_513120[11:1] + 11'h5b9;
  assign sel_530029 = $signed({1'h0, add_529365, array_index_513022[0]}) < $signed({1'h0, sel_529367}) ? {add_529365, array_index_513022[0]} : sel_529367;
  assign add_530031 = array_index_513123[11:1] + 11'h5b9;
  assign sel_530033 = $signed({1'h0, add_529369, array_index_513025[0]}) < $signed({1'h0, sel_529371}) ? {add_529369, array_index_513025[0]} : sel_529371;
  assign add_530043 = array_index_513374[11:0] + 12'h37b;
  assign sel_530045 = $signed({1'h0, add_529381}) < $signed({1'h0, sel_529383}) ? add_529381 : sel_529383;
  assign add_530047 = array_index_513377[11:0] + 12'h37b;
  assign sel_530049 = $signed({1'h0, add_529385}) < $signed({1'h0, sel_529387}) ? add_529385 : sel_529387;
  assign add_530061 = array_index_513702[11:0] + 12'h811;
  assign sel_530063 = $signed({1'h0, add_529399}) < $signed({1'h0, sel_529401}) ? add_529399 : sel_529401;
  assign add_530065 = array_index_513705[11:0] + 12'h811;
  assign sel_530067 = $signed({1'h0, add_529403}) < $signed({1'h0, sel_529405}) ? add_529403 : sel_529405;
  assign add_530079 = array_index_514096[11:0] + 12'h70f;
  assign sel_530081 = $signed({1'h0, add_529417}) < $signed({1'h0, sel_529419}) ? add_529417 : sel_529419;
  assign add_530083 = array_index_514099[11:0] + 12'h70f;
  assign sel_530085 = $signed({1'h0, add_529421}) < $signed({1'h0, sel_529423}) ? add_529421 : sel_529423;
  assign add_530097 = array_index_514558[11:3] + 9'h1f1;
  assign sel_530099 = $signed({1'h0, add_529435, array_index_514318[2:0]}) < $signed({1'h0, sel_529437}) ? {add_529435, array_index_514318[2:0]} : sel_529437;
  assign add_530101 = array_index_514561[11:3] + 9'h1f1;
  assign sel_530103 = $signed({1'h0, add_529439, array_index_514321[2:0]}) < $signed({1'h0, sel_529441}) ? {add_529439, array_index_514321[2:0]} : sel_529441;
  assign add_530113 = array_index_515098[11:0] + 12'h081;
  assign sel_530115 = $signed({1'h0, add_529451}) < $signed({1'h0, sel_529453}) ? add_529451 : sel_529453;
  assign add_530117 = array_index_515101[11:0] + 12'h081;
  assign sel_530119 = $signed({1'h0, add_529455}) < $signed({1'h0, sel_529457}) ? add_529455 : sel_529457;
  assign add_530131 = array_index_515726[11:0] + 12'h0b1;
  assign sel_530133 = $signed({1'h0, add_529469}) < $signed({1'h0, sel_529471}) ? add_529469 : sel_529471;
  assign add_530135 = array_index_515729[11:0] + 12'h0b1;
  assign sel_530137 = $signed({1'h0, add_529473}) < $signed({1'h0, sel_529475}) ? add_529473 : sel_529475;
  assign add_530149 = array_index_516458[11:1] + 11'h4c1;
  assign sel_530151 = $signed({1'h0, add_529487, array_index_516080[0]}) < $signed({1'h0, sel_529489}) ? {add_529487, array_index_516080[0]} : sel_529489;
  assign add_530153 = array_index_516461[11:1] + 11'h4c1;
  assign sel_530155 = $signed({1'h0, add_529491, array_index_516083[0]}) < $signed({1'h0, sel_529493}) ? {add_529491, array_index_516083[0]} : sel_529493;
  assign add_530165 = array_index_517286[11:0] + 12'hbb1;
  assign sel_530167 = $signed({1'h0, add_529503}) < $signed({1'h0, sel_529505}) ? add_529503 : sel_529505;
  assign add_530169 = array_index_517289[11:0] + 12'hbb1;
  assign sel_530171 = $signed({1'h0, add_529507}) < $signed({1'h0, sel_529509}) ? add_529507 : sel_529509;
  assign add_530181 = array_index_518210[11:0] + 12'h6ab;
  assign sel_530183 = $signed({1'h0, add_529519}) < $signed({1'h0, sel_529521}) ? add_529519 : sel_529521;
  assign add_530185 = array_index_518213[11:0] + 12'h6ab;
  assign sel_530187 = $signed({1'h0, add_529523}) < $signed({1'h0, sel_529525}) ? add_529523 : sel_529525;
  assign add_530197 = array_index_519236[11:0] + 12'h7d5;
  assign sel_530199 = $signed({1'h0, add_529535}) < $signed({1'h0, sel_529537}) ? add_529535 : sel_529537;
  assign add_530201 = array_index_519239[11:0] + 12'h7d5;
  assign sel_530203 = $signed({1'h0, add_529539}) < $signed({1'h0, sel_529541}) ? add_529539 : sel_529541;
  assign add_530227 = concat_530016 + 12'h001;
  assign add_530229 = array_index_513022[11:0] + 12'hcc1;
  assign sel_530231 = $signed({1'h0, add_529571}) < $signed({1'h0, sel_529573}) ? add_529571 : sel_529573;
  assign add_530233 = array_index_513025[11:0] + 12'hcc1;
  assign sel_530235 = $signed({1'h0, add_529575}) < $signed({1'h0, sel_529577}) ? add_529575 : sel_529577;
  assign add_530247 = array_index_513238[11:0] + 12'ha87;
  assign sel_530249 = $signed({1'h0, add_529589}) < $signed({1'h0, sel_529591}) ? add_529589 : sel_529591;
  assign add_530251 = array_index_513241[11:0] + 12'ha87;
  assign sel_530253 = $signed({1'h0, add_529593}) < $signed({1'h0, sel_529595}) ? add_529593 : sel_529595;
  assign add_530265 = array_index_513530[11:1] + 11'h663;
  assign sel_530267 = $signed({1'h0, add_529607, array_index_513374[0]}) < $signed({1'h0, sel_529609}) ? {add_529607, array_index_513374[0]} : sel_529609;
  assign add_530269 = array_index_513533[11:1] + 11'h663;
  assign sel_530271 = $signed({1'h0, add_529611, array_index_513377[0]}) < $signed({1'h0, sel_529613}) ? {add_529611, array_index_513377[0]} : sel_529613;
  assign add_530281 = array_index_513890[11:1] + 11'h075;
  assign sel_530283 = $signed({1'h0, add_529623, array_index_513702[0]}) < $signed({1'h0, sel_529625}) ? {add_529623, array_index_513702[0]} : sel_529625;
  assign add_530285 = array_index_513893[11:1] + 11'h075;
  assign sel_530287 = $signed({1'h0, add_529627, array_index_513705[0]}) < $signed({1'h0, sel_529629}) ? {add_529627, array_index_513705[0]} : sel_529629;
  assign add_530299 = array_index_514318[11:2] + 10'h181;
  assign sel_530301 = $signed({1'h0, add_529641, array_index_514096[1:0]}) < $signed({1'h0, sel_529643}) ? {add_529641, array_index_514096[1:0]} : sel_529643;
  assign add_530303 = array_index_514321[11:2] + 10'h181;
  assign sel_530305 = $signed({1'h0, add_529645, array_index_514099[1:0]}) < $signed({1'h0, sel_529647}) ? {add_529645, array_index_514099[1:0]} : sel_529647;
  assign add_530317 = array_index_514818[11:0] + 12'h8a7;
  assign sel_530319 = $signed({1'h0, add_529659}) < $signed({1'h0, sel_529661}) ? add_529659 : sel_529661;
  assign add_530321 = array_index_514821[11:0] + 12'h8a7;
  assign sel_530323 = $signed({1'h0, add_529663}) < $signed({1'h0, sel_529665}) ? add_529663 : sel_529665;
  assign add_530335 = array_index_515398[11:1] + 11'h283;
  assign sel_530337 = $signed({1'h0, add_529677, array_index_515098[0]}) < $signed({1'h0, sel_529679}) ? {add_529677, array_index_515098[0]} : sel_529679;
  assign add_530339 = array_index_515401[11:1] + 11'h283;
  assign sel_530341 = $signed({1'h0, add_529681, array_index_515101[0]}) < $signed({1'h0, sel_529683}) ? {add_529681, array_index_515101[0]} : sel_529683;
  assign add_530351 = array_index_516080[11:1] + 11'h44d;
  assign sel_530353 = $signed({1'h0, add_529693, array_index_515726[0]}) < $signed({1'h0, sel_529695}) ? {add_529693, array_index_515726[0]} : sel_529695;
  assign add_530355 = array_index_516083[11:1] + 11'h44d;
  assign sel_530357 = $signed({1'h0, add_529697, array_index_515729[0]}) < $signed({1'h0, sel_529699}) ? {add_529697, array_index_515729[0]} : sel_529699;
  assign add_530367 = array_index_516860[11:0] + 12'hcb1;
  assign sel_530369 = $signed({1'h0, add_529709}) < $signed({1'h0, sel_529711}) ? add_529709 : sel_529711;
  assign add_530371 = array_index_516863[11:0] + 12'hcb1;
  assign sel_530373 = $signed({1'h0, add_529713}) < $signed({1'h0, sel_529715}) ? add_529713 : sel_529715;
  assign add_530383 = array_index_517736[11:0] + 12'h81f;
  assign sel_530385 = $signed({1'h0, add_529725}) < $signed({1'h0, sel_529727}) ? add_529725 : sel_529727;
  assign add_530387 = array_index_517739[11:0] + 12'h81f;
  assign sel_530389 = $signed({1'h0, add_529729}) < $signed({1'h0, sel_529731}) ? add_529729 : sel_529731;
  assign add_530399 = array_index_518710[11:0] + 12'h45b;
  assign sel_530401 = $signed({1'h0, add_529741}) < $signed({1'h0, sel_529743}) ? add_529741 : sel_529743;
  assign add_530403 = array_index_518713[11:0] + 12'h45b;
  assign sel_530405 = $signed({1'h0, add_529745}) < $signed({1'h0, sel_529747}) ? add_529745 : sel_529747;
  assign add_530417 = array_index_519786[11:3] + 9'h0f5;
  assign sel_530419 = $signed({1'h0, add_529759, array_index_519236[2:0]}) < $signed({1'h0, sel_529761}) ? {add_529759, array_index_519236[2:0]} : sel_529761;
  assign add_530421 = array_index_519789[11:3] + 9'h0f5;
  assign sel_530423 = $signed({1'h0, add_529763, array_index_519239[2:0]}) < $signed({1'h0, sel_529765}) ? {add_529763, array_index_519239[2:0]} : sel_529765;
  assign add_530453 = array_index_513120[11:2] + 10'h113;
  assign sel_530455 = $signed({1'h0, add_529799, array_index_513022[1:0]}) < $signed({1'h0, sel_529801}) ? {add_529799, array_index_513022[1:0]} : sel_529801;
  assign add_530457 = array_index_513123[11:2] + 10'h113;
  assign sel_530459 = $signed({1'h0, add_529803, array_index_513025[1:0]}) < $signed({1'h0, sel_529805}) ? {add_529803, array_index_513025[1:0]} : sel_529805;
  assign add_530471 = array_index_513374[11:4] + 8'h49;
  assign sel_530473 = $signed({1'h0, add_529817, array_index_513238[3:0]}) < $signed({1'h0, sel_529819}) ? {add_529817, array_index_513238[3:0]} : sel_529819;
  assign add_530475 = array_index_513377[11:4] + 8'h49;
  assign sel_530477 = $signed({1'h0, add_529821, array_index_513241[3:0]}) < $signed({1'h0, sel_529823}) ? {add_529821, array_index_513241[3:0]} : sel_529823;
  assign add_530487 = array_index_513702[11:0] + 12'h263;
  assign sel_530489 = $signed({1'h0, add_529833}) < $signed({1'h0, sel_529835}) ? add_529833 : sel_529835;
  assign add_530491 = array_index_513705[11:0] + 12'h263;
  assign sel_530493 = $signed({1'h0, add_529837}) < $signed({1'h0, sel_529839}) ? add_529837 : sel_529839;
  assign add_530503 = array_index_514096[11:1] + 11'h109;
  assign sel_530505 = $signed({1'h0, add_529849, array_index_513890[0]}) < $signed({1'h0, sel_529851}) ? {add_529849, array_index_513890[0]} : sel_529851;
  assign add_530507 = array_index_514099[11:1] + 11'h109;
  assign sel_530509 = $signed({1'h0, add_529853, array_index_513893[0]}) < $signed({1'h0, sel_529855}) ? {add_529853, array_index_513893[0]} : sel_529855;
  assign add_530519 = array_index_514558[11:3] + 9'h12f;
  assign sel_530521 = $signed({1'h0, add_529865, array_index_514318[2:0]}) < $signed({1'h0, sel_529867}) ? {add_529865, array_index_514318[2:0]} : sel_529867;
  assign add_530523 = array_index_514561[11:3] + 9'h12f;
  assign sel_530525 = $signed({1'h0, add_529869, array_index_514321[2:0]}) < $signed({1'h0, sel_529871}) ? {add_529869, array_index_514321[2:0]} : sel_529871;
  assign add_530537 = array_index_515098[11:3] + 9'h171;
  assign sel_530539 = $signed({1'h0, add_529883, array_index_514818[2:0]}) < $signed({1'h0, sel_529885}) ? {add_529883, array_index_514818[2:0]} : sel_529885;
  assign add_530541 = array_index_515101[11:3] + 9'h171;
  assign sel_530543 = $signed({1'h0, add_529887, array_index_514821[2:0]}) < $signed({1'h0, sel_529889}) ? {add_529887, array_index_514821[2:0]} : sel_529889;
  assign add_530553 = array_index_515726[11:0] + 12'h091;
  assign sel_530555 = $signed({1'h0, add_529899}) < $signed({1'h0, sel_529901}) ? add_529899 : sel_529901;
  assign add_530557 = array_index_515729[11:0] + 12'h091;
  assign sel_530559 = $signed({1'h0, add_529903}) < $signed({1'h0, sel_529905}) ? add_529903 : sel_529905;
  assign add_530569 = array_index_516458[11:0] + 12'hf59;
  assign sel_530571 = $signed({1'h0, add_529915}) < $signed({1'h0, sel_529917}) ? add_529915 : sel_529917;
  assign add_530573 = array_index_516461[11:0] + 12'hf59;
  assign sel_530575 = $signed({1'h0, add_529919}) < $signed({1'h0, sel_529921}) ? add_529919 : sel_529921;
  assign add_530587 = array_index_517286[11:0] + 12'h437;
  assign sel_530589 = $signed({1'h0, add_529933}) < $signed({1'h0, sel_529935}) ? add_529933 : sel_529935;
  assign add_530591 = array_index_517289[11:0] + 12'h437;
  assign sel_530593 = $signed({1'h0, add_529937}) < $signed({1'h0, sel_529939}) ? add_529937 : sel_529939;
  assign add_530603 = array_index_518210[11:0] + 12'hee1;
  assign sel_530605 = $signed({1'h0, add_529949}) < $signed({1'h0, sel_529951}) ? add_529949 : sel_529951;
  assign add_530607 = array_index_518213[11:0] + 12'hee1;
  assign sel_530609 = $signed({1'h0, add_529953}) < $signed({1'h0, sel_529955}) ? add_529953 : sel_529955;
  assign add_530619 = array_index_519236[11:1] + 11'h179;
  assign sel_530621 = $signed({1'h0, add_529965, array_index_518710[0]}) < $signed({1'h0, sel_529967}) ? {add_529965, array_index_518710[0]} : sel_529967;
  assign add_530623 = array_index_519239[11:1] + 11'h179;
  assign sel_530625 = $signed({1'h0, add_529969, array_index_518713[0]}) < $signed({1'h0, sel_529971}) ? {add_529969, array_index_518713[0]} : sel_529971;
  assign add_530635 = array_index_520362[11:0] + 12'h067;
  assign sel_530637 = $signed({1'h0, add_529981}) < $signed({1'h0, sel_529983}) ? add_529981 : sel_529983;
  assign add_530639 = array_index_520365[11:0] + 12'h067;
  assign sel_530641 = $signed({1'h0, add_529985}) < $signed({1'h0, sel_529987}) ? add_529985 : sel_529987;
  assign add_530643 = array_index_520964[11:3] + 9'h1ef;
  assign sel_530646 = $signed({1'h0, add_529989, array_index_520362[2:0]}) < $signed({1'h0, sel_529992}) ? {add_529989, array_index_520362[2:0]} : sel_529992;
  assign add_530648 = array_index_520967[11:3] + 9'h1ef;
  assign sel_530651 = $signed({1'h0, add_529994, array_index_520365[2:0]}) < $signed({1'h0, sel_529997}) ? {add_529994, array_index_520365[2:0]} : sel_529997;
  assign add_530653 = array_index_521590[11:1] + 11'h2d5;
  assign sel_530655 = $signed({1'h0, add_529999, array_index_520964[0]}) < $signed({1'h0, sel_530001}) ? {add_529999, array_index_520964[0]} : sel_530001;
  assign add_530657 = array_index_521593[11:1] + 11'h2d5;
  assign sel_530659 = $signed({1'h0, add_530003, array_index_520967[0]}) < $signed({1'h0, sel_530005}) ? {add_530003, array_index_520967[0]} : sel_530005;
  assign concat_530662 = {1'h0, ($signed({1'h0, add_529345}) < $signed({1'h0, sel_529347}) ? add_529345 : sel_529347) == ($signed({1'h0, add_529349}) < $signed({1'h0, sel_529351}) ? add_529349 : sel_529351) ? add_530227 : concat_530016};
  assign add_530673 = array_index_513238[11:1] + 11'h5b9;
  assign sel_530675 = $signed({1'h0, add_530027, array_index_513120[0]}) < $signed({1'h0, sel_530029}) ? {add_530027, array_index_513120[0]} : sel_530029;
  assign add_530677 = array_index_513241[11:1] + 11'h5b9;
  assign sel_530679 = $signed({1'h0, add_530031, array_index_513123[0]}) < $signed({1'h0, sel_530033}) ? {add_530031, array_index_513123[0]} : sel_530033;
  assign add_530689 = array_index_513530[11:0] + 12'h37b;
  assign sel_530691 = $signed({1'h0, add_530043}) < $signed({1'h0, sel_530045}) ? add_530043 : sel_530045;
  assign add_530693 = array_index_513533[11:0] + 12'h37b;
  assign sel_530695 = $signed({1'h0, add_530047}) < $signed({1'h0, sel_530049}) ? add_530047 : sel_530049;
  assign add_530707 = array_index_513890[11:0] + 12'h811;
  assign sel_530709 = $signed({1'h0, add_530061}) < $signed({1'h0, sel_530063}) ? add_530061 : sel_530063;
  assign add_530711 = array_index_513893[11:0] + 12'h811;
  assign sel_530713 = $signed({1'h0, add_530065}) < $signed({1'h0, sel_530067}) ? add_530065 : sel_530067;
  assign add_530725 = array_index_514318[11:0] + 12'h70f;
  assign sel_530727 = $signed({1'h0, add_530079}) < $signed({1'h0, sel_530081}) ? add_530079 : sel_530081;
  assign add_530729 = array_index_514321[11:0] + 12'h70f;
  assign sel_530731 = $signed({1'h0, add_530083}) < $signed({1'h0, sel_530085}) ? add_530083 : sel_530085;
  assign add_530743 = array_index_514818[11:3] + 9'h1f1;
  assign sel_530745 = $signed({1'h0, add_530097, array_index_514558[2:0]}) < $signed({1'h0, sel_530099}) ? {add_530097, array_index_514558[2:0]} : sel_530099;
  assign add_530747 = array_index_514821[11:3] + 9'h1f1;
  assign sel_530749 = $signed({1'h0, add_530101, array_index_514561[2:0]}) < $signed({1'h0, sel_530103}) ? {add_530101, array_index_514561[2:0]} : sel_530103;
  assign add_530759 = array_index_515398[11:0] + 12'h081;
  assign sel_530761 = $signed({1'h0, add_530113}) < $signed({1'h0, sel_530115}) ? add_530113 : sel_530115;
  assign add_530763 = array_index_515401[11:0] + 12'h081;
  assign sel_530765 = $signed({1'h0, add_530117}) < $signed({1'h0, sel_530119}) ? add_530117 : sel_530119;
  assign add_530777 = array_index_516080[11:0] + 12'h0b1;
  assign sel_530779 = $signed({1'h0, add_530131}) < $signed({1'h0, sel_530133}) ? add_530131 : sel_530133;
  assign add_530781 = array_index_516083[11:0] + 12'h0b1;
  assign sel_530783 = $signed({1'h0, add_530135}) < $signed({1'h0, sel_530137}) ? add_530135 : sel_530137;
  assign add_530795 = array_index_516860[11:1] + 11'h4c1;
  assign sel_530797 = $signed({1'h0, add_530149, array_index_516458[0]}) < $signed({1'h0, sel_530151}) ? {add_530149, array_index_516458[0]} : sel_530151;
  assign add_530799 = array_index_516863[11:1] + 11'h4c1;
  assign sel_530801 = $signed({1'h0, add_530153, array_index_516461[0]}) < $signed({1'h0, sel_530155}) ? {add_530153, array_index_516461[0]} : sel_530155;
  assign add_530811 = array_index_517736[11:0] + 12'hbb1;
  assign sel_530813 = $signed({1'h0, add_530165}) < $signed({1'h0, sel_530167}) ? add_530165 : sel_530167;
  assign add_530815 = array_index_517739[11:0] + 12'hbb1;
  assign sel_530817 = $signed({1'h0, add_530169}) < $signed({1'h0, sel_530171}) ? add_530169 : sel_530171;
  assign add_530827 = array_index_518710[11:0] + 12'h6ab;
  assign sel_530829 = $signed({1'h0, add_530181}) < $signed({1'h0, sel_530183}) ? add_530181 : sel_530183;
  assign add_530831 = array_index_518713[11:0] + 12'h6ab;
  assign sel_530833 = $signed({1'h0, add_530185}) < $signed({1'h0, sel_530187}) ? add_530185 : sel_530187;
  assign add_530843 = array_index_519786[11:0] + 12'h7d5;
  assign sel_530845 = $signed({1'h0, add_530197}) < $signed({1'h0, sel_530199}) ? add_530197 : sel_530199;
  assign add_530847 = array_index_519789[11:0] + 12'h7d5;
  assign sel_530849 = $signed({1'h0, add_530201}) < $signed({1'h0, sel_530203}) ? add_530201 : sel_530203;
  assign add_530869 = concat_530662 + 13'h0001;
  assign add_530871 = array_index_513120[11:0] + 12'hcc1;
  assign sel_530873 = $signed({1'h0, add_530229}) < $signed({1'h0, sel_530231}) ? add_530229 : sel_530231;
  assign add_530875 = array_index_513123[11:0] + 12'hcc1;
  assign sel_530877 = $signed({1'h0, add_530233}) < $signed({1'h0, sel_530235}) ? add_530233 : sel_530235;
  assign add_530889 = array_index_513374[11:0] + 12'ha87;
  assign sel_530891 = $signed({1'h0, add_530247}) < $signed({1'h0, sel_530249}) ? add_530247 : sel_530249;
  assign add_530893 = array_index_513377[11:0] + 12'ha87;
  assign sel_530895 = $signed({1'h0, add_530251}) < $signed({1'h0, sel_530253}) ? add_530251 : sel_530253;
  assign add_530907 = array_index_513702[11:1] + 11'h663;
  assign sel_530909 = $signed({1'h0, add_530265, array_index_513530[0]}) < $signed({1'h0, sel_530267}) ? {add_530265, array_index_513530[0]} : sel_530267;
  assign add_530911 = array_index_513705[11:1] + 11'h663;
  assign sel_530913 = $signed({1'h0, add_530269, array_index_513533[0]}) < $signed({1'h0, sel_530271}) ? {add_530269, array_index_513533[0]} : sel_530271;
  assign add_530923 = array_index_514096[11:1] + 11'h075;
  assign sel_530925 = $signed({1'h0, add_530281, array_index_513890[0]}) < $signed({1'h0, sel_530283}) ? {add_530281, array_index_513890[0]} : sel_530283;
  assign add_530927 = array_index_514099[11:1] + 11'h075;
  assign sel_530929 = $signed({1'h0, add_530285, array_index_513893[0]}) < $signed({1'h0, sel_530287}) ? {add_530285, array_index_513893[0]} : sel_530287;
  assign add_530941 = array_index_514558[11:2] + 10'h181;
  assign sel_530943 = $signed({1'h0, add_530299, array_index_514318[1:0]}) < $signed({1'h0, sel_530301}) ? {add_530299, array_index_514318[1:0]} : sel_530301;
  assign add_530945 = array_index_514561[11:2] + 10'h181;
  assign sel_530947 = $signed({1'h0, add_530303, array_index_514321[1:0]}) < $signed({1'h0, sel_530305}) ? {add_530303, array_index_514321[1:0]} : sel_530305;
  assign add_530959 = array_index_515098[11:0] + 12'h8a7;
  assign sel_530961 = $signed({1'h0, add_530317}) < $signed({1'h0, sel_530319}) ? add_530317 : sel_530319;
  assign add_530963 = array_index_515101[11:0] + 12'h8a7;
  assign sel_530965 = $signed({1'h0, add_530321}) < $signed({1'h0, sel_530323}) ? add_530321 : sel_530323;
  assign add_530977 = array_index_515726[11:1] + 11'h283;
  assign sel_530979 = $signed({1'h0, add_530335, array_index_515398[0]}) < $signed({1'h0, sel_530337}) ? {add_530335, array_index_515398[0]} : sel_530337;
  assign add_530981 = array_index_515729[11:1] + 11'h283;
  assign sel_530983 = $signed({1'h0, add_530339, array_index_515401[0]}) < $signed({1'h0, sel_530341}) ? {add_530339, array_index_515401[0]} : sel_530341;
  assign add_530993 = array_index_516458[11:1] + 11'h44d;
  assign sel_530995 = $signed({1'h0, add_530351, array_index_516080[0]}) < $signed({1'h0, sel_530353}) ? {add_530351, array_index_516080[0]} : sel_530353;
  assign add_530997 = array_index_516461[11:1] + 11'h44d;
  assign sel_530999 = $signed({1'h0, add_530355, array_index_516083[0]}) < $signed({1'h0, sel_530357}) ? {add_530355, array_index_516083[0]} : sel_530357;
  assign add_531009 = array_index_517286[11:0] + 12'hcb1;
  assign sel_531011 = $signed({1'h0, add_530367}) < $signed({1'h0, sel_530369}) ? add_530367 : sel_530369;
  assign add_531013 = array_index_517289[11:0] + 12'hcb1;
  assign sel_531015 = $signed({1'h0, add_530371}) < $signed({1'h0, sel_530373}) ? add_530371 : sel_530373;
  assign add_531025 = array_index_518210[11:0] + 12'h81f;
  assign sel_531027 = $signed({1'h0, add_530383}) < $signed({1'h0, sel_530385}) ? add_530383 : sel_530385;
  assign add_531029 = array_index_518213[11:0] + 12'h81f;
  assign sel_531031 = $signed({1'h0, add_530387}) < $signed({1'h0, sel_530389}) ? add_530387 : sel_530389;
  assign add_531041 = array_index_519236[11:0] + 12'h45b;
  assign sel_531043 = $signed({1'h0, add_530399}) < $signed({1'h0, sel_530401}) ? add_530399 : sel_530401;
  assign add_531045 = array_index_519239[11:0] + 12'h45b;
  assign sel_531047 = $signed({1'h0, add_530403}) < $signed({1'h0, sel_530405}) ? add_530403 : sel_530405;
  assign add_531059 = array_index_520362[11:3] + 9'h0f5;
  assign sel_531061 = $signed({1'h0, add_530417, array_index_519786[2:0]}) < $signed({1'h0, sel_530419}) ? {add_530417, array_index_519786[2:0]} : sel_530419;
  assign add_531063 = array_index_520365[11:3] + 9'h0f5;
  assign sel_531065 = $signed({1'h0, add_530421, array_index_519789[2:0]}) < $signed({1'h0, sel_530423}) ? {add_530421, array_index_519789[2:0]} : sel_530423;
  assign add_531089 = array_index_513238[11:2] + 10'h113;
  assign sel_531091 = $signed({1'h0, add_530453, array_index_513120[1:0]}) < $signed({1'h0, sel_530455}) ? {add_530453, array_index_513120[1:0]} : sel_530455;
  assign add_531093 = array_index_513241[11:2] + 10'h113;
  assign sel_531095 = $signed({1'h0, add_530457, array_index_513123[1:0]}) < $signed({1'h0, sel_530459}) ? {add_530457, array_index_513123[1:0]} : sel_530459;
  assign add_531107 = array_index_513530[11:4] + 8'h49;
  assign sel_531109 = $signed({1'h0, add_530471, array_index_513374[3:0]}) < $signed({1'h0, sel_530473}) ? {add_530471, array_index_513374[3:0]} : sel_530473;
  assign add_531111 = array_index_513533[11:4] + 8'h49;
  assign sel_531113 = $signed({1'h0, add_530475, array_index_513377[3:0]}) < $signed({1'h0, sel_530477}) ? {add_530475, array_index_513377[3:0]} : sel_530477;
  assign add_531123 = array_index_513890[11:0] + 12'h263;
  assign sel_531125 = $signed({1'h0, add_530487}) < $signed({1'h0, sel_530489}) ? add_530487 : sel_530489;
  assign add_531127 = array_index_513893[11:0] + 12'h263;
  assign sel_531129 = $signed({1'h0, add_530491}) < $signed({1'h0, sel_530493}) ? add_530491 : sel_530493;
  assign add_531139 = array_index_514318[11:1] + 11'h109;
  assign sel_531141 = $signed({1'h0, add_530503, array_index_514096[0]}) < $signed({1'h0, sel_530505}) ? {add_530503, array_index_514096[0]} : sel_530505;
  assign add_531143 = array_index_514321[11:1] + 11'h109;
  assign sel_531145 = $signed({1'h0, add_530507, array_index_514099[0]}) < $signed({1'h0, sel_530509}) ? {add_530507, array_index_514099[0]} : sel_530509;
  assign add_531155 = array_index_514818[11:3] + 9'h12f;
  assign sel_531157 = $signed({1'h0, add_530519, array_index_514558[2:0]}) < $signed({1'h0, sel_530521}) ? {add_530519, array_index_514558[2:0]} : sel_530521;
  assign add_531159 = array_index_514821[11:3] + 9'h12f;
  assign sel_531161 = $signed({1'h0, add_530523, array_index_514561[2:0]}) < $signed({1'h0, sel_530525}) ? {add_530523, array_index_514561[2:0]} : sel_530525;
  assign add_531173 = array_index_515398[11:3] + 9'h171;
  assign sel_531175 = $signed({1'h0, add_530537, array_index_515098[2:0]}) < $signed({1'h0, sel_530539}) ? {add_530537, array_index_515098[2:0]} : sel_530539;
  assign add_531177 = array_index_515401[11:3] + 9'h171;
  assign sel_531179 = $signed({1'h0, add_530541, array_index_515101[2:0]}) < $signed({1'h0, sel_530543}) ? {add_530541, array_index_515101[2:0]} : sel_530543;
  assign add_531189 = array_index_516080[11:0] + 12'h091;
  assign sel_531191 = $signed({1'h0, add_530553}) < $signed({1'h0, sel_530555}) ? add_530553 : sel_530555;
  assign add_531193 = array_index_516083[11:0] + 12'h091;
  assign sel_531195 = $signed({1'h0, add_530557}) < $signed({1'h0, sel_530559}) ? add_530557 : sel_530559;
  assign add_531205 = array_index_516860[11:0] + 12'hf59;
  assign sel_531207 = $signed({1'h0, add_530569}) < $signed({1'h0, sel_530571}) ? add_530569 : sel_530571;
  assign add_531209 = array_index_516863[11:0] + 12'hf59;
  assign sel_531211 = $signed({1'h0, add_530573}) < $signed({1'h0, sel_530575}) ? add_530573 : sel_530575;
  assign add_531223 = array_index_517736[11:0] + 12'h437;
  assign sel_531225 = $signed({1'h0, add_530587}) < $signed({1'h0, sel_530589}) ? add_530587 : sel_530589;
  assign add_531227 = array_index_517739[11:0] + 12'h437;
  assign sel_531229 = $signed({1'h0, add_530591}) < $signed({1'h0, sel_530593}) ? add_530591 : sel_530593;
  assign add_531239 = array_index_518710[11:0] + 12'hee1;
  assign sel_531241 = $signed({1'h0, add_530603}) < $signed({1'h0, sel_530605}) ? add_530603 : sel_530605;
  assign add_531243 = array_index_518713[11:0] + 12'hee1;
  assign sel_531245 = $signed({1'h0, add_530607}) < $signed({1'h0, sel_530609}) ? add_530607 : sel_530609;
  assign add_531255 = array_index_519786[11:1] + 11'h179;
  assign sel_531257 = $signed({1'h0, add_530619, array_index_519236[0]}) < $signed({1'h0, sel_530621}) ? {add_530619, array_index_519236[0]} : sel_530621;
  assign add_531259 = array_index_519789[11:1] + 11'h179;
  assign sel_531261 = $signed({1'h0, add_530623, array_index_519239[0]}) < $signed({1'h0, sel_530625}) ? {add_530623, array_index_519239[0]} : sel_530625;
  assign add_531271 = array_index_520964[11:0] + 12'h067;
  assign sel_531273 = $signed({1'h0, add_530635}) < $signed({1'h0, sel_530637}) ? add_530635 : sel_530637;
  assign add_531275 = array_index_520967[11:0] + 12'h067;
  assign sel_531277 = $signed({1'h0, add_530639}) < $signed({1'h0, sel_530641}) ? add_530639 : sel_530641;
  assign add_531279 = array_index_521590[11:3] + 9'h1ef;
  assign sel_531282 = $signed({1'h0, add_530643, array_index_520964[2:0]}) < $signed({1'h0, sel_530646}) ? {add_530643, array_index_520964[2:0]} : sel_530646;
  assign add_531284 = array_index_521593[11:3] + 9'h1ef;
  assign sel_531287 = $signed({1'h0, add_530648, array_index_520967[2:0]}) < $signed({1'h0, sel_530651}) ? {add_530648, array_index_520967[2:0]} : sel_530651;
  assign concat_531290 = {1'h0, ($signed({1'h0, add_530007, array_index_521590[1:0]}) < $signed({1'h0, sel_530009}) ? {add_530007, array_index_521590[1:0]} : sel_530009) == ($signed({1'h0, add_530011, array_index_521593[1:0]}) < $signed({1'h0, sel_530013}) ? {add_530011, array_index_521593[1:0]} : sel_530013) ? add_530869 : concat_530662};
  assign add_531301 = array_index_513374[11:1] + 11'h5b9;
  assign sel_531303 = $signed({1'h0, add_530673, array_index_513238[0]}) < $signed({1'h0, sel_530675}) ? {add_530673, array_index_513238[0]} : sel_530675;
  assign add_531305 = array_index_513377[11:1] + 11'h5b9;
  assign sel_531307 = $signed({1'h0, add_530677, array_index_513241[0]}) < $signed({1'h0, sel_530679}) ? {add_530677, array_index_513241[0]} : sel_530679;
  assign add_531317 = array_index_513702[11:0] + 12'h37b;
  assign sel_531319 = $signed({1'h0, add_530689}) < $signed({1'h0, sel_530691}) ? add_530689 : sel_530691;
  assign add_531321 = array_index_513705[11:0] + 12'h37b;
  assign sel_531323 = $signed({1'h0, add_530693}) < $signed({1'h0, sel_530695}) ? add_530693 : sel_530695;
  assign add_531335 = array_index_514096[11:0] + 12'h811;
  assign sel_531337 = $signed({1'h0, add_530707}) < $signed({1'h0, sel_530709}) ? add_530707 : sel_530709;
  assign add_531339 = array_index_514099[11:0] + 12'h811;
  assign sel_531341 = $signed({1'h0, add_530711}) < $signed({1'h0, sel_530713}) ? add_530711 : sel_530713;
  assign add_531353 = array_index_514558[11:0] + 12'h70f;
  assign sel_531355 = $signed({1'h0, add_530725}) < $signed({1'h0, sel_530727}) ? add_530725 : sel_530727;
  assign add_531357 = array_index_514561[11:0] + 12'h70f;
  assign sel_531359 = $signed({1'h0, add_530729}) < $signed({1'h0, sel_530731}) ? add_530729 : sel_530731;
  assign add_531371 = array_index_515098[11:3] + 9'h1f1;
  assign sel_531373 = $signed({1'h0, add_530743, array_index_514818[2:0]}) < $signed({1'h0, sel_530745}) ? {add_530743, array_index_514818[2:0]} : sel_530745;
  assign add_531375 = array_index_515101[11:3] + 9'h1f1;
  assign sel_531377 = $signed({1'h0, add_530747, array_index_514821[2:0]}) < $signed({1'h0, sel_530749}) ? {add_530747, array_index_514821[2:0]} : sel_530749;
  assign add_531387 = array_index_515726[11:0] + 12'h081;
  assign sel_531389 = $signed({1'h0, add_530759}) < $signed({1'h0, sel_530761}) ? add_530759 : sel_530761;
  assign add_531391 = array_index_515729[11:0] + 12'h081;
  assign sel_531393 = $signed({1'h0, add_530763}) < $signed({1'h0, sel_530765}) ? add_530763 : sel_530765;
  assign add_531405 = array_index_516458[11:0] + 12'h0b1;
  assign sel_531407 = $signed({1'h0, add_530777}) < $signed({1'h0, sel_530779}) ? add_530777 : sel_530779;
  assign add_531409 = array_index_516461[11:0] + 12'h0b1;
  assign sel_531411 = $signed({1'h0, add_530781}) < $signed({1'h0, sel_530783}) ? add_530781 : sel_530783;
  assign add_531423 = array_index_517286[11:1] + 11'h4c1;
  assign sel_531425 = $signed({1'h0, add_530795, array_index_516860[0]}) < $signed({1'h0, sel_530797}) ? {add_530795, array_index_516860[0]} : sel_530797;
  assign add_531427 = array_index_517289[11:1] + 11'h4c1;
  assign sel_531429 = $signed({1'h0, add_530799, array_index_516863[0]}) < $signed({1'h0, sel_530801}) ? {add_530799, array_index_516863[0]} : sel_530801;
  assign add_531439 = array_index_518210[11:0] + 12'hbb1;
  assign sel_531441 = $signed({1'h0, add_530811}) < $signed({1'h0, sel_530813}) ? add_530811 : sel_530813;
  assign add_531443 = array_index_518213[11:0] + 12'hbb1;
  assign sel_531445 = $signed({1'h0, add_530815}) < $signed({1'h0, sel_530817}) ? add_530815 : sel_530817;
  assign add_531455 = array_index_519236[11:0] + 12'h6ab;
  assign sel_531457 = $signed({1'h0, add_530827}) < $signed({1'h0, sel_530829}) ? add_530827 : sel_530829;
  assign add_531459 = array_index_519239[11:0] + 12'h6ab;
  assign sel_531461 = $signed({1'h0, add_530831}) < $signed({1'h0, sel_530833}) ? add_530831 : sel_530833;
  assign add_531471 = array_index_520362[11:0] + 12'h7d5;
  assign sel_531473 = $signed({1'h0, add_530843}) < $signed({1'h0, sel_530845}) ? add_530843 : sel_530845;
  assign add_531475 = array_index_520365[11:0] + 12'h7d5;
  assign sel_531477 = $signed({1'h0, add_530847}) < $signed({1'h0, sel_530849}) ? add_530847 : sel_530849;
  assign add_531493 = concat_531290 + 14'h0001;
  assign add_531495 = array_index_513238[11:0] + 12'hcc1;
  assign sel_531497 = $signed({1'h0, add_530871}) < $signed({1'h0, sel_530873}) ? add_530871 : sel_530873;
  assign add_531499 = array_index_513241[11:0] + 12'hcc1;
  assign sel_531501 = $signed({1'h0, add_530875}) < $signed({1'h0, sel_530877}) ? add_530875 : sel_530877;
  assign add_531513 = array_index_513530[11:0] + 12'ha87;
  assign sel_531515 = $signed({1'h0, add_530889}) < $signed({1'h0, sel_530891}) ? add_530889 : sel_530891;
  assign add_531517 = array_index_513533[11:0] + 12'ha87;
  assign sel_531519 = $signed({1'h0, add_530893}) < $signed({1'h0, sel_530895}) ? add_530893 : sel_530895;
  assign add_531531 = array_index_513890[11:1] + 11'h663;
  assign sel_531533 = $signed({1'h0, add_530907, array_index_513702[0]}) < $signed({1'h0, sel_530909}) ? {add_530907, array_index_513702[0]} : sel_530909;
  assign add_531535 = array_index_513893[11:1] + 11'h663;
  assign sel_531537 = $signed({1'h0, add_530911, array_index_513705[0]}) < $signed({1'h0, sel_530913}) ? {add_530911, array_index_513705[0]} : sel_530913;
  assign add_531547 = array_index_514318[11:1] + 11'h075;
  assign sel_531549 = $signed({1'h0, add_530923, array_index_514096[0]}) < $signed({1'h0, sel_530925}) ? {add_530923, array_index_514096[0]} : sel_530925;
  assign add_531551 = array_index_514321[11:1] + 11'h075;
  assign sel_531553 = $signed({1'h0, add_530927, array_index_514099[0]}) < $signed({1'h0, sel_530929}) ? {add_530927, array_index_514099[0]} : sel_530929;
  assign add_531565 = array_index_514818[11:2] + 10'h181;
  assign sel_531567 = $signed({1'h0, add_530941, array_index_514558[1:0]}) < $signed({1'h0, sel_530943}) ? {add_530941, array_index_514558[1:0]} : sel_530943;
  assign add_531569 = array_index_514821[11:2] + 10'h181;
  assign sel_531571 = $signed({1'h0, add_530945, array_index_514561[1:0]}) < $signed({1'h0, sel_530947}) ? {add_530945, array_index_514561[1:0]} : sel_530947;
  assign add_531583 = array_index_515398[11:0] + 12'h8a7;
  assign sel_531585 = $signed({1'h0, add_530959}) < $signed({1'h0, sel_530961}) ? add_530959 : sel_530961;
  assign add_531587 = array_index_515401[11:0] + 12'h8a7;
  assign sel_531589 = $signed({1'h0, add_530963}) < $signed({1'h0, sel_530965}) ? add_530963 : sel_530965;
  assign add_531601 = array_index_516080[11:1] + 11'h283;
  assign sel_531603 = $signed({1'h0, add_530977, array_index_515726[0]}) < $signed({1'h0, sel_530979}) ? {add_530977, array_index_515726[0]} : sel_530979;
  assign add_531605 = array_index_516083[11:1] + 11'h283;
  assign sel_531607 = $signed({1'h0, add_530981, array_index_515729[0]}) < $signed({1'h0, sel_530983}) ? {add_530981, array_index_515729[0]} : sel_530983;
  assign add_531617 = array_index_516860[11:1] + 11'h44d;
  assign sel_531619 = $signed({1'h0, add_530993, array_index_516458[0]}) < $signed({1'h0, sel_530995}) ? {add_530993, array_index_516458[0]} : sel_530995;
  assign add_531621 = array_index_516863[11:1] + 11'h44d;
  assign sel_531623 = $signed({1'h0, add_530997, array_index_516461[0]}) < $signed({1'h0, sel_530999}) ? {add_530997, array_index_516461[0]} : sel_530999;
  assign add_531633 = array_index_517736[11:0] + 12'hcb1;
  assign sel_531635 = $signed({1'h0, add_531009}) < $signed({1'h0, sel_531011}) ? add_531009 : sel_531011;
  assign add_531637 = array_index_517739[11:0] + 12'hcb1;
  assign sel_531639 = $signed({1'h0, add_531013}) < $signed({1'h0, sel_531015}) ? add_531013 : sel_531015;
  assign add_531649 = array_index_518710[11:0] + 12'h81f;
  assign sel_531651 = $signed({1'h0, add_531025}) < $signed({1'h0, sel_531027}) ? add_531025 : sel_531027;
  assign add_531653 = array_index_518713[11:0] + 12'h81f;
  assign sel_531655 = $signed({1'h0, add_531029}) < $signed({1'h0, sel_531031}) ? add_531029 : sel_531031;
  assign add_531665 = array_index_519786[11:0] + 12'h45b;
  assign sel_531667 = $signed({1'h0, add_531041}) < $signed({1'h0, sel_531043}) ? add_531041 : sel_531043;
  assign add_531669 = array_index_519789[11:0] + 12'h45b;
  assign sel_531671 = $signed({1'h0, add_531045}) < $signed({1'h0, sel_531047}) ? add_531045 : sel_531047;
  assign add_531683 = array_index_520964[11:3] + 9'h0f5;
  assign sel_531685 = $signed({1'h0, add_531059, array_index_520362[2:0]}) < $signed({1'h0, sel_531061}) ? {add_531059, array_index_520362[2:0]} : sel_531061;
  assign add_531687 = array_index_520967[11:3] + 9'h0f5;
  assign sel_531689 = $signed({1'h0, add_531063, array_index_520365[2:0]}) < $signed({1'h0, sel_531065}) ? {add_531063, array_index_520365[2:0]} : sel_531065;
  assign add_531705 = array_index_513374[11:2] + 10'h113;
  assign sel_531707 = $signed({1'h0, add_531089, array_index_513238[1:0]}) < $signed({1'h0, sel_531091}) ? {add_531089, array_index_513238[1:0]} : sel_531091;
  assign add_531709 = array_index_513377[11:2] + 10'h113;
  assign sel_531711 = $signed({1'h0, add_531093, array_index_513241[1:0]}) < $signed({1'h0, sel_531095}) ? {add_531093, array_index_513241[1:0]} : sel_531095;
  assign add_531723 = array_index_513702[11:4] + 8'h49;
  assign sel_531725 = $signed({1'h0, add_531107, array_index_513530[3:0]}) < $signed({1'h0, sel_531109}) ? {add_531107, array_index_513530[3:0]} : sel_531109;
  assign add_531727 = array_index_513705[11:4] + 8'h49;
  assign sel_531729 = $signed({1'h0, add_531111, array_index_513533[3:0]}) < $signed({1'h0, sel_531113}) ? {add_531111, array_index_513533[3:0]} : sel_531113;
  assign add_531739 = array_index_514096[11:0] + 12'h263;
  assign sel_531741 = $signed({1'h0, add_531123}) < $signed({1'h0, sel_531125}) ? add_531123 : sel_531125;
  assign add_531743 = array_index_514099[11:0] + 12'h263;
  assign sel_531745 = $signed({1'h0, add_531127}) < $signed({1'h0, sel_531129}) ? add_531127 : sel_531129;
  assign add_531755 = array_index_514558[11:1] + 11'h109;
  assign sel_531757 = $signed({1'h0, add_531139, array_index_514318[0]}) < $signed({1'h0, sel_531141}) ? {add_531139, array_index_514318[0]} : sel_531141;
  assign add_531759 = array_index_514561[11:1] + 11'h109;
  assign sel_531761 = $signed({1'h0, add_531143, array_index_514321[0]}) < $signed({1'h0, sel_531145}) ? {add_531143, array_index_514321[0]} : sel_531145;
  assign add_531771 = array_index_515098[11:3] + 9'h12f;
  assign sel_531773 = $signed({1'h0, add_531155, array_index_514818[2:0]}) < $signed({1'h0, sel_531157}) ? {add_531155, array_index_514818[2:0]} : sel_531157;
  assign add_531775 = array_index_515101[11:3] + 9'h12f;
  assign sel_531777 = $signed({1'h0, add_531159, array_index_514821[2:0]}) < $signed({1'h0, sel_531161}) ? {add_531159, array_index_514821[2:0]} : sel_531161;
  assign add_531789 = array_index_515726[11:3] + 9'h171;
  assign sel_531791 = $signed({1'h0, add_531173, array_index_515398[2:0]}) < $signed({1'h0, sel_531175}) ? {add_531173, array_index_515398[2:0]} : sel_531175;
  assign add_531793 = array_index_515729[11:3] + 9'h171;
  assign sel_531795 = $signed({1'h0, add_531177, array_index_515401[2:0]}) < $signed({1'h0, sel_531179}) ? {add_531177, array_index_515401[2:0]} : sel_531179;
  assign add_531805 = array_index_516458[11:0] + 12'h091;
  assign sel_531807 = $signed({1'h0, add_531189}) < $signed({1'h0, sel_531191}) ? add_531189 : sel_531191;
  assign add_531809 = array_index_516461[11:0] + 12'h091;
  assign sel_531811 = $signed({1'h0, add_531193}) < $signed({1'h0, sel_531195}) ? add_531193 : sel_531195;
  assign add_531821 = array_index_517286[11:0] + 12'hf59;
  assign sel_531823 = $signed({1'h0, add_531205}) < $signed({1'h0, sel_531207}) ? add_531205 : sel_531207;
  assign add_531825 = array_index_517289[11:0] + 12'hf59;
  assign sel_531827 = $signed({1'h0, add_531209}) < $signed({1'h0, sel_531211}) ? add_531209 : sel_531211;
  assign add_531839 = array_index_518210[11:0] + 12'h437;
  assign sel_531841 = $signed({1'h0, add_531223}) < $signed({1'h0, sel_531225}) ? add_531223 : sel_531225;
  assign add_531843 = array_index_518213[11:0] + 12'h437;
  assign sel_531845 = $signed({1'h0, add_531227}) < $signed({1'h0, sel_531229}) ? add_531227 : sel_531229;
  assign add_531855 = array_index_519236[11:0] + 12'hee1;
  assign sel_531857 = $signed({1'h0, add_531239}) < $signed({1'h0, sel_531241}) ? add_531239 : sel_531241;
  assign add_531859 = array_index_519239[11:0] + 12'hee1;
  assign sel_531861 = $signed({1'h0, add_531243}) < $signed({1'h0, sel_531245}) ? add_531243 : sel_531245;
  assign add_531871 = array_index_520362[11:1] + 11'h179;
  assign sel_531873 = $signed({1'h0, add_531255, array_index_519786[0]}) < $signed({1'h0, sel_531257}) ? {add_531255, array_index_519786[0]} : sel_531257;
  assign add_531875 = array_index_520365[11:1] + 11'h179;
  assign sel_531877 = $signed({1'h0, add_531259, array_index_519789[0]}) < $signed({1'h0, sel_531261}) ? {add_531259, array_index_519789[0]} : sel_531261;
  assign add_531887 = array_index_521590[11:0] + 12'h067;
  assign sel_531889 = $signed({1'h0, add_531271}) < $signed({1'h0, sel_531273}) ? add_531271 : sel_531273;
  assign add_531891 = array_index_521593[11:0] + 12'h067;
  assign sel_531893 = $signed({1'h0, add_531275}) < $signed({1'h0, sel_531277}) ? add_531275 : sel_531277;
  assign concat_531896 = {1'h0, ($signed({1'h0, add_530653, array_index_521590[0]}) < $signed({1'h0, sel_530655}) ? {add_530653, array_index_521590[0]} : sel_530655) == ($signed({1'h0, add_530657, array_index_521593[0]}) < $signed({1'h0, sel_530659}) ? {add_530657, array_index_521593[0]} : sel_530659) ? add_531493 : concat_531290};
  assign add_531907 = array_index_513530[11:1] + 11'h5b9;
  assign sel_531909 = $signed({1'h0, add_531301, array_index_513374[0]}) < $signed({1'h0, sel_531303}) ? {add_531301, array_index_513374[0]} : sel_531303;
  assign add_531911 = array_index_513533[11:1] + 11'h5b9;
  assign sel_531913 = $signed({1'h0, add_531305, array_index_513377[0]}) < $signed({1'h0, sel_531307}) ? {add_531305, array_index_513377[0]} : sel_531307;
  assign add_531923 = array_index_513890[11:0] + 12'h37b;
  assign sel_531925 = $signed({1'h0, add_531317}) < $signed({1'h0, sel_531319}) ? add_531317 : sel_531319;
  assign add_531927 = array_index_513893[11:0] + 12'h37b;
  assign sel_531929 = $signed({1'h0, add_531321}) < $signed({1'h0, sel_531323}) ? add_531321 : sel_531323;
  assign add_531941 = array_index_514318[11:0] + 12'h811;
  assign sel_531943 = $signed({1'h0, add_531335}) < $signed({1'h0, sel_531337}) ? add_531335 : sel_531337;
  assign add_531945 = array_index_514321[11:0] + 12'h811;
  assign sel_531947 = $signed({1'h0, add_531339}) < $signed({1'h0, sel_531341}) ? add_531339 : sel_531341;
  assign add_531959 = array_index_514818[11:0] + 12'h70f;
  assign sel_531961 = $signed({1'h0, add_531353}) < $signed({1'h0, sel_531355}) ? add_531353 : sel_531355;
  assign add_531963 = array_index_514821[11:0] + 12'h70f;
  assign sel_531965 = $signed({1'h0, add_531357}) < $signed({1'h0, sel_531359}) ? add_531357 : sel_531359;
  assign add_531977 = array_index_515398[11:3] + 9'h1f1;
  assign sel_531979 = $signed({1'h0, add_531371, array_index_515098[2:0]}) < $signed({1'h0, sel_531373}) ? {add_531371, array_index_515098[2:0]} : sel_531373;
  assign add_531981 = array_index_515401[11:3] + 9'h1f1;
  assign sel_531983 = $signed({1'h0, add_531375, array_index_515101[2:0]}) < $signed({1'h0, sel_531377}) ? {add_531375, array_index_515101[2:0]} : sel_531377;
  assign add_531993 = array_index_516080[11:0] + 12'h081;
  assign sel_531995 = $signed({1'h0, add_531387}) < $signed({1'h0, sel_531389}) ? add_531387 : sel_531389;
  assign add_531997 = array_index_516083[11:0] + 12'h081;
  assign sel_531999 = $signed({1'h0, add_531391}) < $signed({1'h0, sel_531393}) ? add_531391 : sel_531393;
  assign add_532011 = array_index_516860[11:0] + 12'h0b1;
  assign sel_532013 = $signed({1'h0, add_531405}) < $signed({1'h0, sel_531407}) ? add_531405 : sel_531407;
  assign add_532015 = array_index_516863[11:0] + 12'h0b1;
  assign sel_532017 = $signed({1'h0, add_531409}) < $signed({1'h0, sel_531411}) ? add_531409 : sel_531411;
  assign add_532029 = array_index_517736[11:1] + 11'h4c1;
  assign sel_532031 = $signed({1'h0, add_531423, array_index_517286[0]}) < $signed({1'h0, sel_531425}) ? {add_531423, array_index_517286[0]} : sel_531425;
  assign add_532033 = array_index_517739[11:1] + 11'h4c1;
  assign sel_532035 = $signed({1'h0, add_531427, array_index_517289[0]}) < $signed({1'h0, sel_531429}) ? {add_531427, array_index_517289[0]} : sel_531429;
  assign add_532045 = array_index_518710[11:0] + 12'hbb1;
  assign sel_532047 = $signed({1'h0, add_531439}) < $signed({1'h0, sel_531441}) ? add_531439 : sel_531441;
  assign add_532049 = array_index_518713[11:0] + 12'hbb1;
  assign sel_532051 = $signed({1'h0, add_531443}) < $signed({1'h0, sel_531445}) ? add_531443 : sel_531445;
  assign add_532061 = array_index_519786[11:0] + 12'h6ab;
  assign sel_532063 = $signed({1'h0, add_531455}) < $signed({1'h0, sel_531457}) ? add_531455 : sel_531457;
  assign add_532065 = array_index_519789[11:0] + 12'h6ab;
  assign sel_532067 = $signed({1'h0, add_531459}) < $signed({1'h0, sel_531461}) ? add_531459 : sel_531461;
  assign add_532077 = array_index_520964[11:0] + 12'h7d5;
  assign sel_532079 = $signed({1'h0, add_531471}) < $signed({1'h0, sel_531473}) ? add_531471 : sel_531473;
  assign add_532081 = array_index_520967[11:0] + 12'h7d5;
  assign sel_532083 = $signed({1'h0, add_531475}) < $signed({1'h0, sel_531477}) ? add_531475 : sel_531477;
  assign add_532095 = concat_531896 + 15'h0001;
  assign add_532097 = array_index_513374[11:0] + 12'hcc1;
  assign sel_532099 = $signed({1'h0, add_531495}) < $signed({1'h0, sel_531497}) ? add_531495 : sel_531497;
  assign add_532101 = array_index_513377[11:0] + 12'hcc1;
  assign sel_532103 = $signed({1'h0, add_531499}) < $signed({1'h0, sel_531501}) ? add_531499 : sel_531501;
  assign add_532115 = array_index_513702[11:0] + 12'ha87;
  assign sel_532117 = $signed({1'h0, add_531513}) < $signed({1'h0, sel_531515}) ? add_531513 : sel_531515;
  assign add_532119 = array_index_513705[11:0] + 12'ha87;
  assign sel_532121 = $signed({1'h0, add_531517}) < $signed({1'h0, sel_531519}) ? add_531517 : sel_531519;
  assign add_532133 = array_index_514096[11:1] + 11'h663;
  assign sel_532135 = $signed({1'h0, add_531531, array_index_513890[0]}) < $signed({1'h0, sel_531533}) ? {add_531531, array_index_513890[0]} : sel_531533;
  assign add_532137 = array_index_514099[11:1] + 11'h663;
  assign sel_532139 = $signed({1'h0, add_531535, array_index_513893[0]}) < $signed({1'h0, sel_531537}) ? {add_531535, array_index_513893[0]} : sel_531537;
  assign add_532149 = array_index_514558[11:1] + 11'h075;
  assign sel_532151 = $signed({1'h0, add_531547, array_index_514318[0]}) < $signed({1'h0, sel_531549}) ? {add_531547, array_index_514318[0]} : sel_531549;
  assign add_532153 = array_index_514561[11:1] + 11'h075;
  assign sel_532155 = $signed({1'h0, add_531551, array_index_514321[0]}) < $signed({1'h0, sel_531553}) ? {add_531551, array_index_514321[0]} : sel_531553;
  assign add_532167 = array_index_515098[11:2] + 10'h181;
  assign sel_532169 = $signed({1'h0, add_531565, array_index_514818[1:0]}) < $signed({1'h0, sel_531567}) ? {add_531565, array_index_514818[1:0]} : sel_531567;
  assign add_532171 = array_index_515101[11:2] + 10'h181;
  assign sel_532173 = $signed({1'h0, add_531569, array_index_514821[1:0]}) < $signed({1'h0, sel_531571}) ? {add_531569, array_index_514821[1:0]} : sel_531571;
  assign add_532185 = array_index_515726[11:0] + 12'h8a7;
  assign sel_532187 = $signed({1'h0, add_531583}) < $signed({1'h0, sel_531585}) ? add_531583 : sel_531585;
  assign add_532189 = array_index_515729[11:0] + 12'h8a7;
  assign sel_532191 = $signed({1'h0, add_531587}) < $signed({1'h0, sel_531589}) ? add_531587 : sel_531589;
  assign add_532203 = array_index_516458[11:1] + 11'h283;
  assign sel_532205 = $signed({1'h0, add_531601, array_index_516080[0]}) < $signed({1'h0, sel_531603}) ? {add_531601, array_index_516080[0]} : sel_531603;
  assign add_532207 = array_index_516461[11:1] + 11'h283;
  assign sel_532209 = $signed({1'h0, add_531605, array_index_516083[0]}) < $signed({1'h0, sel_531607}) ? {add_531605, array_index_516083[0]} : sel_531607;
  assign add_532219 = array_index_517286[11:1] + 11'h44d;
  assign sel_532221 = $signed({1'h0, add_531617, array_index_516860[0]}) < $signed({1'h0, sel_531619}) ? {add_531617, array_index_516860[0]} : sel_531619;
  assign add_532223 = array_index_517289[11:1] + 11'h44d;
  assign sel_532225 = $signed({1'h0, add_531621, array_index_516863[0]}) < $signed({1'h0, sel_531623}) ? {add_531621, array_index_516863[0]} : sel_531623;
  assign add_532235 = array_index_518210[11:0] + 12'hcb1;
  assign sel_532237 = $signed({1'h0, add_531633}) < $signed({1'h0, sel_531635}) ? add_531633 : sel_531635;
  assign add_532239 = array_index_518213[11:0] + 12'hcb1;
  assign sel_532241 = $signed({1'h0, add_531637}) < $signed({1'h0, sel_531639}) ? add_531637 : sel_531639;
  assign add_532251 = array_index_519236[11:0] + 12'h81f;
  assign sel_532253 = $signed({1'h0, add_531649}) < $signed({1'h0, sel_531651}) ? add_531649 : sel_531651;
  assign add_532255 = array_index_519239[11:0] + 12'h81f;
  assign sel_532257 = $signed({1'h0, add_531653}) < $signed({1'h0, sel_531655}) ? add_531653 : sel_531655;
  assign add_532267 = array_index_520362[11:0] + 12'h45b;
  assign sel_532269 = $signed({1'h0, add_531665}) < $signed({1'h0, sel_531667}) ? add_531665 : sel_531667;
  assign add_532271 = array_index_520365[11:0] + 12'h45b;
  assign sel_532273 = $signed({1'h0, add_531669}) < $signed({1'h0, sel_531671}) ? add_531669 : sel_531671;
  assign add_532285 = array_index_521590[11:3] + 9'h0f5;
  assign sel_532287 = $signed({1'h0, add_531683, array_index_520964[2:0]}) < $signed({1'h0, sel_531685}) ? {add_531683, array_index_520964[2:0]} : sel_531685;
  assign add_532289 = array_index_521593[11:3] + 9'h0f5;
  assign sel_532291 = $signed({1'h0, add_531687, array_index_520967[2:0]}) < $signed({1'h0, sel_531689}) ? {add_531687, array_index_520967[2:0]} : sel_531689;
  assign add_532301 = array_index_513530[11:2] + 10'h113;
  assign sel_532303 = $signed({1'h0, add_531705, array_index_513374[1:0]}) < $signed({1'h0, sel_531707}) ? {add_531705, array_index_513374[1:0]} : sel_531707;
  assign add_532305 = array_index_513533[11:2] + 10'h113;
  assign sel_532307 = $signed({1'h0, add_531709, array_index_513377[1:0]}) < $signed({1'h0, sel_531711}) ? {add_531709, array_index_513377[1:0]} : sel_531711;
  assign add_532319 = array_index_513890[11:4] + 8'h49;
  assign sel_532321 = $signed({1'h0, add_531723, array_index_513702[3:0]}) < $signed({1'h0, sel_531725}) ? {add_531723, array_index_513702[3:0]} : sel_531725;
  assign add_532323 = array_index_513893[11:4] + 8'h49;
  assign sel_532325 = $signed({1'h0, add_531727, array_index_513705[3:0]}) < $signed({1'h0, sel_531729}) ? {add_531727, array_index_513705[3:0]} : sel_531729;
  assign add_532335 = array_index_514318[11:0] + 12'h263;
  assign sel_532337 = $signed({1'h0, add_531739}) < $signed({1'h0, sel_531741}) ? add_531739 : sel_531741;
  assign add_532339 = array_index_514321[11:0] + 12'h263;
  assign sel_532341 = $signed({1'h0, add_531743}) < $signed({1'h0, sel_531745}) ? add_531743 : sel_531745;
  assign add_532351 = array_index_514818[11:1] + 11'h109;
  assign sel_532353 = $signed({1'h0, add_531755, array_index_514558[0]}) < $signed({1'h0, sel_531757}) ? {add_531755, array_index_514558[0]} : sel_531757;
  assign add_532355 = array_index_514821[11:1] + 11'h109;
  assign sel_532357 = $signed({1'h0, add_531759, array_index_514561[0]}) < $signed({1'h0, sel_531761}) ? {add_531759, array_index_514561[0]} : sel_531761;
  assign add_532367 = array_index_515398[11:3] + 9'h12f;
  assign sel_532369 = $signed({1'h0, add_531771, array_index_515098[2:0]}) < $signed({1'h0, sel_531773}) ? {add_531771, array_index_515098[2:0]} : sel_531773;
  assign add_532371 = array_index_515401[11:3] + 9'h12f;
  assign sel_532373 = $signed({1'h0, add_531775, array_index_515101[2:0]}) < $signed({1'h0, sel_531777}) ? {add_531775, array_index_515101[2:0]} : sel_531777;
  assign add_532385 = array_index_516080[11:3] + 9'h171;
  assign sel_532387 = $signed({1'h0, add_531789, array_index_515726[2:0]}) < $signed({1'h0, sel_531791}) ? {add_531789, array_index_515726[2:0]} : sel_531791;
  assign add_532389 = array_index_516083[11:3] + 9'h171;
  assign sel_532391 = $signed({1'h0, add_531793, array_index_515729[2:0]}) < $signed({1'h0, sel_531795}) ? {add_531793, array_index_515729[2:0]} : sel_531795;
  assign add_532401 = array_index_516860[11:0] + 12'h091;
  assign sel_532403 = $signed({1'h0, add_531805}) < $signed({1'h0, sel_531807}) ? add_531805 : sel_531807;
  assign add_532405 = array_index_516863[11:0] + 12'h091;
  assign sel_532407 = $signed({1'h0, add_531809}) < $signed({1'h0, sel_531811}) ? add_531809 : sel_531811;
  assign add_532417 = array_index_517736[11:0] + 12'hf59;
  assign sel_532419 = $signed({1'h0, add_531821}) < $signed({1'h0, sel_531823}) ? add_531821 : sel_531823;
  assign add_532421 = array_index_517739[11:0] + 12'hf59;
  assign sel_532423 = $signed({1'h0, add_531825}) < $signed({1'h0, sel_531827}) ? add_531825 : sel_531827;
  assign add_532435 = array_index_518710[11:0] + 12'h437;
  assign sel_532437 = $signed({1'h0, add_531839}) < $signed({1'h0, sel_531841}) ? add_531839 : sel_531841;
  assign add_532439 = array_index_518713[11:0] + 12'h437;
  assign sel_532441 = $signed({1'h0, add_531843}) < $signed({1'h0, sel_531845}) ? add_531843 : sel_531845;
  assign add_532451 = array_index_519786[11:0] + 12'hee1;
  assign sel_532453 = $signed({1'h0, add_531855}) < $signed({1'h0, sel_531857}) ? add_531855 : sel_531857;
  assign add_532455 = array_index_519789[11:0] + 12'hee1;
  assign sel_532457 = $signed({1'h0, add_531859}) < $signed({1'h0, sel_531861}) ? add_531859 : sel_531861;
  assign add_532467 = array_index_520964[11:1] + 11'h179;
  assign sel_532469 = $signed({1'h0, add_531871, array_index_520362[0]}) < $signed({1'h0, sel_531873}) ? {add_531871, array_index_520362[0]} : sel_531873;
  assign add_532471 = array_index_520967[11:1] + 11'h179;
  assign sel_532473 = $signed({1'h0, add_531875, array_index_520365[0]}) < $signed({1'h0, sel_531877}) ? {add_531875, array_index_520365[0]} : sel_531877;
  assign concat_532484 = {1'h0, ($signed({1'h0, add_531279, array_index_521590[2:0]}) < $signed({1'h0, sel_531282}) ? {add_531279, array_index_521590[2:0]} : sel_531282) == ($signed({1'h0, add_531284, array_index_521593[2:0]}) < $signed({1'h0, sel_531287}) ? {add_531284, array_index_521593[2:0]} : sel_531287) ? add_532095 : concat_531896};
  assign add_532495 = array_index_513702[11:1] + 11'h5b9;
  assign sel_532497 = $signed({1'h0, add_531907, array_index_513530[0]}) < $signed({1'h0, sel_531909}) ? {add_531907, array_index_513530[0]} : sel_531909;
  assign add_532499 = array_index_513705[11:1] + 11'h5b9;
  assign sel_532501 = $signed({1'h0, add_531911, array_index_513533[0]}) < $signed({1'h0, sel_531913}) ? {add_531911, array_index_513533[0]} : sel_531913;
  assign add_532511 = array_index_514096[11:0] + 12'h37b;
  assign sel_532513 = $signed({1'h0, add_531923}) < $signed({1'h0, sel_531925}) ? add_531923 : sel_531925;
  assign add_532515 = array_index_514099[11:0] + 12'h37b;
  assign sel_532517 = $signed({1'h0, add_531927}) < $signed({1'h0, sel_531929}) ? add_531927 : sel_531929;
  assign add_532529 = array_index_514558[11:0] + 12'h811;
  assign sel_532531 = $signed({1'h0, add_531941}) < $signed({1'h0, sel_531943}) ? add_531941 : sel_531943;
  assign add_532533 = array_index_514561[11:0] + 12'h811;
  assign sel_532535 = $signed({1'h0, add_531945}) < $signed({1'h0, sel_531947}) ? add_531945 : sel_531947;
  assign add_532547 = array_index_515098[11:0] + 12'h70f;
  assign sel_532549 = $signed({1'h0, add_531959}) < $signed({1'h0, sel_531961}) ? add_531959 : sel_531961;
  assign add_532551 = array_index_515101[11:0] + 12'h70f;
  assign sel_532553 = $signed({1'h0, add_531963}) < $signed({1'h0, sel_531965}) ? add_531963 : sel_531965;
  assign add_532565 = array_index_515726[11:3] + 9'h1f1;
  assign sel_532567 = $signed({1'h0, add_531977, array_index_515398[2:0]}) < $signed({1'h0, sel_531979}) ? {add_531977, array_index_515398[2:0]} : sel_531979;
  assign add_532569 = array_index_515729[11:3] + 9'h1f1;
  assign sel_532571 = $signed({1'h0, add_531981, array_index_515401[2:0]}) < $signed({1'h0, sel_531983}) ? {add_531981, array_index_515401[2:0]} : sel_531983;
  assign add_532581 = array_index_516458[11:0] + 12'h081;
  assign sel_532583 = $signed({1'h0, add_531993}) < $signed({1'h0, sel_531995}) ? add_531993 : sel_531995;
  assign add_532585 = array_index_516461[11:0] + 12'h081;
  assign sel_532587 = $signed({1'h0, add_531997}) < $signed({1'h0, sel_531999}) ? add_531997 : sel_531999;
  assign add_532599 = array_index_517286[11:0] + 12'h0b1;
  assign sel_532601 = $signed({1'h0, add_532011}) < $signed({1'h0, sel_532013}) ? add_532011 : sel_532013;
  assign add_532603 = array_index_517289[11:0] + 12'h0b1;
  assign sel_532605 = $signed({1'h0, add_532015}) < $signed({1'h0, sel_532017}) ? add_532015 : sel_532017;
  assign add_532617 = array_index_518210[11:1] + 11'h4c1;
  assign sel_532619 = $signed({1'h0, add_532029, array_index_517736[0]}) < $signed({1'h0, sel_532031}) ? {add_532029, array_index_517736[0]} : sel_532031;
  assign add_532621 = array_index_518213[11:1] + 11'h4c1;
  assign sel_532623 = $signed({1'h0, add_532033, array_index_517739[0]}) < $signed({1'h0, sel_532035}) ? {add_532033, array_index_517739[0]} : sel_532035;
  assign add_532633 = array_index_519236[11:0] + 12'hbb1;
  assign sel_532635 = $signed({1'h0, add_532045}) < $signed({1'h0, sel_532047}) ? add_532045 : sel_532047;
  assign add_532637 = array_index_519239[11:0] + 12'hbb1;
  assign sel_532639 = $signed({1'h0, add_532049}) < $signed({1'h0, sel_532051}) ? add_532049 : sel_532051;
  assign add_532649 = array_index_520362[11:0] + 12'h6ab;
  assign sel_532651 = $signed({1'h0, add_532061}) < $signed({1'h0, sel_532063}) ? add_532061 : sel_532063;
  assign add_532653 = array_index_520365[11:0] + 12'h6ab;
  assign sel_532655 = $signed({1'h0, add_532065}) < $signed({1'h0, sel_532067}) ? add_532065 : sel_532067;
  assign add_532665 = array_index_521590[11:0] + 12'h7d5;
  assign sel_532667 = $signed({1'h0, add_532077}) < $signed({1'h0, sel_532079}) ? add_532077 : sel_532079;
  assign add_532669 = array_index_521593[11:0] + 12'h7d5;
  assign sel_532671 = $signed({1'h0, add_532081}) < $signed({1'h0, sel_532083}) ? add_532081 : sel_532083;
  assign add_532677 = concat_532484 + 16'h0001;
  assign add_532679 = array_index_513530[11:0] + 12'hcc1;
  assign sel_532681 = $signed({1'h0, add_532097}) < $signed({1'h0, sel_532099}) ? add_532097 : sel_532099;
  assign add_532683 = array_index_513533[11:0] + 12'hcc1;
  assign sel_532685 = $signed({1'h0, add_532101}) < $signed({1'h0, sel_532103}) ? add_532101 : sel_532103;
  assign add_532697 = array_index_513890[11:0] + 12'ha87;
  assign sel_532699 = $signed({1'h0, add_532115}) < $signed({1'h0, sel_532117}) ? add_532115 : sel_532117;
  assign add_532701 = array_index_513893[11:0] + 12'ha87;
  assign sel_532703 = $signed({1'h0, add_532119}) < $signed({1'h0, sel_532121}) ? add_532119 : sel_532121;
  assign add_532715 = array_index_514318[11:1] + 11'h663;
  assign sel_532717 = $signed({1'h0, add_532133, array_index_514096[0]}) < $signed({1'h0, sel_532135}) ? {add_532133, array_index_514096[0]} : sel_532135;
  assign add_532719 = array_index_514321[11:1] + 11'h663;
  assign sel_532721 = $signed({1'h0, add_532137, array_index_514099[0]}) < $signed({1'h0, sel_532139}) ? {add_532137, array_index_514099[0]} : sel_532139;
  assign add_532731 = array_index_514818[11:1] + 11'h075;
  assign sel_532733 = $signed({1'h0, add_532149, array_index_514558[0]}) < $signed({1'h0, sel_532151}) ? {add_532149, array_index_514558[0]} : sel_532151;
  assign add_532735 = array_index_514821[11:1] + 11'h075;
  assign sel_532737 = $signed({1'h0, add_532153, array_index_514561[0]}) < $signed({1'h0, sel_532155}) ? {add_532153, array_index_514561[0]} : sel_532155;
  assign add_532749 = array_index_515398[11:2] + 10'h181;
  assign sel_532751 = $signed({1'h0, add_532167, array_index_515098[1:0]}) < $signed({1'h0, sel_532169}) ? {add_532167, array_index_515098[1:0]} : sel_532169;
  assign add_532753 = array_index_515401[11:2] + 10'h181;
  assign sel_532755 = $signed({1'h0, add_532171, array_index_515101[1:0]}) < $signed({1'h0, sel_532173}) ? {add_532171, array_index_515101[1:0]} : sel_532173;
  assign add_532767 = array_index_516080[11:0] + 12'h8a7;
  assign sel_532769 = $signed({1'h0, add_532185}) < $signed({1'h0, sel_532187}) ? add_532185 : sel_532187;
  assign add_532771 = array_index_516083[11:0] + 12'h8a7;
  assign sel_532773 = $signed({1'h0, add_532189}) < $signed({1'h0, sel_532191}) ? add_532189 : sel_532191;
  assign add_532785 = array_index_516860[11:1] + 11'h283;
  assign sel_532787 = $signed({1'h0, add_532203, array_index_516458[0]}) < $signed({1'h0, sel_532205}) ? {add_532203, array_index_516458[0]} : sel_532205;
  assign add_532789 = array_index_516863[11:1] + 11'h283;
  assign sel_532791 = $signed({1'h0, add_532207, array_index_516461[0]}) < $signed({1'h0, sel_532209}) ? {add_532207, array_index_516461[0]} : sel_532209;
  assign add_532801 = array_index_517736[11:1] + 11'h44d;
  assign sel_532803 = $signed({1'h0, add_532219, array_index_517286[0]}) < $signed({1'h0, sel_532221}) ? {add_532219, array_index_517286[0]} : sel_532221;
  assign add_532805 = array_index_517739[11:1] + 11'h44d;
  assign sel_532807 = $signed({1'h0, add_532223, array_index_517289[0]}) < $signed({1'h0, sel_532225}) ? {add_532223, array_index_517289[0]} : sel_532225;
  assign add_532817 = array_index_518710[11:0] + 12'hcb1;
  assign sel_532819 = $signed({1'h0, add_532235}) < $signed({1'h0, sel_532237}) ? add_532235 : sel_532237;
  assign add_532821 = array_index_518713[11:0] + 12'hcb1;
  assign sel_532823 = $signed({1'h0, add_532239}) < $signed({1'h0, sel_532241}) ? add_532239 : sel_532241;
  assign add_532833 = array_index_519786[11:0] + 12'h81f;
  assign sel_532835 = $signed({1'h0, add_532251}) < $signed({1'h0, sel_532253}) ? add_532251 : sel_532253;
  assign add_532837 = array_index_519789[11:0] + 12'h81f;
  assign sel_532839 = $signed({1'h0, add_532255}) < $signed({1'h0, sel_532257}) ? add_532255 : sel_532257;
  assign add_532849 = array_index_520964[11:0] + 12'h45b;
  assign sel_532851 = $signed({1'h0, add_532267}) < $signed({1'h0, sel_532269}) ? add_532267 : sel_532269;
  assign add_532853 = array_index_520967[11:0] + 12'h45b;
  assign sel_532855 = $signed({1'h0, add_532271}) < $signed({1'h0, sel_532273}) ? add_532271 : sel_532273;
  assign sel_532868 = ($signed({1'h0, add_531887}) < $signed({1'h0, sel_531889}) ? add_531887 : sel_531889) == ($signed({1'h0, add_531891}) < $signed({1'h0, sel_531893}) ? add_531891 : sel_531893) ? add_532677 : concat_532484;
  assign add_532875 = array_index_513702[11:2] + 10'h113;
  assign sel_532877 = $signed({1'h0, add_532301, array_index_513530[1:0]}) < $signed({1'h0, sel_532303}) ? {add_532301, array_index_513530[1:0]} : sel_532303;
  assign add_532879 = array_index_513705[11:2] + 10'h113;
  assign sel_532881 = $signed({1'h0, add_532305, array_index_513533[1:0]}) < $signed({1'h0, sel_532307}) ? {add_532305, array_index_513533[1:0]} : sel_532307;
  assign add_532893 = array_index_514096[11:4] + 8'h49;
  assign sel_532895 = $signed({1'h0, add_532319, array_index_513890[3:0]}) < $signed({1'h0, sel_532321}) ? {add_532319, array_index_513890[3:0]} : sel_532321;
  assign add_532897 = array_index_514099[11:4] + 8'h49;
  assign sel_532899 = $signed({1'h0, add_532323, array_index_513893[3:0]}) < $signed({1'h0, sel_532325}) ? {add_532323, array_index_513893[3:0]} : sel_532325;
  assign add_532909 = array_index_514558[11:0] + 12'h263;
  assign sel_532911 = $signed({1'h0, add_532335}) < $signed({1'h0, sel_532337}) ? add_532335 : sel_532337;
  assign add_532913 = array_index_514561[11:0] + 12'h263;
  assign sel_532915 = $signed({1'h0, add_532339}) < $signed({1'h0, sel_532341}) ? add_532339 : sel_532341;
  assign add_532925 = array_index_515098[11:1] + 11'h109;
  assign sel_532927 = $signed({1'h0, add_532351, array_index_514818[0]}) < $signed({1'h0, sel_532353}) ? {add_532351, array_index_514818[0]} : sel_532353;
  assign add_532929 = array_index_515101[11:1] + 11'h109;
  assign sel_532931 = $signed({1'h0, add_532355, array_index_514821[0]}) < $signed({1'h0, sel_532357}) ? {add_532355, array_index_514821[0]} : sel_532357;
  assign add_532941 = array_index_515726[11:3] + 9'h12f;
  assign sel_532943 = $signed({1'h0, add_532367, array_index_515398[2:0]}) < $signed({1'h0, sel_532369}) ? {add_532367, array_index_515398[2:0]} : sel_532369;
  assign add_532945 = array_index_515729[11:3] + 9'h12f;
  assign sel_532947 = $signed({1'h0, add_532371, array_index_515401[2:0]}) < $signed({1'h0, sel_532373}) ? {add_532371, array_index_515401[2:0]} : sel_532373;
  assign add_532959 = array_index_516458[11:3] + 9'h171;
  assign sel_532961 = $signed({1'h0, add_532385, array_index_516080[2:0]}) < $signed({1'h0, sel_532387}) ? {add_532385, array_index_516080[2:0]} : sel_532387;
  assign add_532963 = array_index_516461[11:3] + 9'h171;
  assign sel_532965 = $signed({1'h0, add_532389, array_index_516083[2:0]}) < $signed({1'h0, sel_532391}) ? {add_532389, array_index_516083[2:0]} : sel_532391;
  assign add_532975 = array_index_517286[11:0] + 12'h091;
  assign sel_532977 = $signed({1'h0, add_532401}) < $signed({1'h0, sel_532403}) ? add_532401 : sel_532403;
  assign add_532979 = array_index_517289[11:0] + 12'h091;
  assign sel_532981 = $signed({1'h0, add_532405}) < $signed({1'h0, sel_532407}) ? add_532405 : sel_532407;
  assign add_532991 = array_index_518210[11:0] + 12'hf59;
  assign sel_532993 = $signed({1'h0, add_532417}) < $signed({1'h0, sel_532419}) ? add_532417 : sel_532419;
  assign add_532995 = array_index_518213[11:0] + 12'hf59;
  assign sel_532997 = $signed({1'h0, add_532421}) < $signed({1'h0, sel_532423}) ? add_532421 : sel_532423;
  assign add_533009 = array_index_519236[11:0] + 12'h437;
  assign sel_533011 = $signed({1'h0, add_532435}) < $signed({1'h0, sel_532437}) ? add_532435 : sel_532437;
  assign add_533013 = array_index_519239[11:0] + 12'h437;
  assign sel_533015 = $signed({1'h0, add_532439}) < $signed({1'h0, sel_532441}) ? add_532439 : sel_532441;
  assign add_533025 = array_index_520362[11:0] + 12'hee1;
  assign sel_533027 = $signed({1'h0, add_532451}) < $signed({1'h0, sel_532453}) ? add_532451 : sel_532453;
  assign add_533029 = array_index_520365[11:0] + 12'hee1;
  assign sel_533031 = $signed({1'h0, add_532455}) < $signed({1'h0, sel_532457}) ? add_532455 : sel_532457;
  assign add_533041 = array_index_521590[11:1] + 11'h179;
  assign sel_533043 = $signed({1'h0, add_532467, array_index_520964[0]}) < $signed({1'h0, sel_532469}) ? {add_532467, array_index_520964[0]} : sel_532469;
  assign add_533045 = array_index_521593[11:1] + 11'h179;
  assign sel_533047 = $signed({1'h0, add_532471, array_index_520967[0]}) < $signed({1'h0, sel_532473}) ? {add_532471, array_index_520967[0]} : sel_532473;
  assign add_533051 = sel_532868 + 16'h0001;
  assign add_533061 = array_index_513890[11:1] + 11'h5b9;
  assign sel_533063 = $signed({1'h0, add_532495, array_index_513702[0]}) < $signed({1'h0, sel_532497}) ? {add_532495, array_index_513702[0]} : sel_532497;
  assign add_533065 = array_index_513893[11:1] + 11'h5b9;
  assign sel_533067 = $signed({1'h0, add_532499, array_index_513705[0]}) < $signed({1'h0, sel_532501}) ? {add_532499, array_index_513705[0]} : sel_532501;
  assign add_533077 = array_index_514318[11:0] + 12'h37b;
  assign sel_533079 = $signed({1'h0, add_532511}) < $signed({1'h0, sel_532513}) ? add_532511 : sel_532513;
  assign add_533081 = array_index_514321[11:0] + 12'h37b;
  assign sel_533083 = $signed({1'h0, add_532515}) < $signed({1'h0, sel_532517}) ? add_532515 : sel_532517;
  assign add_533095 = array_index_514818[11:0] + 12'h811;
  assign sel_533097 = $signed({1'h0, add_532529}) < $signed({1'h0, sel_532531}) ? add_532529 : sel_532531;
  assign add_533099 = array_index_514821[11:0] + 12'h811;
  assign sel_533101 = $signed({1'h0, add_532533}) < $signed({1'h0, sel_532535}) ? add_532533 : sel_532535;
  assign add_533113 = array_index_515398[11:0] + 12'h70f;
  assign sel_533115 = $signed({1'h0, add_532547}) < $signed({1'h0, sel_532549}) ? add_532547 : sel_532549;
  assign add_533117 = array_index_515401[11:0] + 12'h70f;
  assign sel_533119 = $signed({1'h0, add_532551}) < $signed({1'h0, sel_532553}) ? add_532551 : sel_532553;
  assign add_533131 = array_index_516080[11:3] + 9'h1f1;
  assign sel_533133 = $signed({1'h0, add_532565, array_index_515726[2:0]}) < $signed({1'h0, sel_532567}) ? {add_532565, array_index_515726[2:0]} : sel_532567;
  assign add_533135 = array_index_516083[11:3] + 9'h1f1;
  assign sel_533137 = $signed({1'h0, add_532569, array_index_515729[2:0]}) < $signed({1'h0, sel_532571}) ? {add_532569, array_index_515729[2:0]} : sel_532571;
  assign add_533147 = array_index_516860[11:0] + 12'h081;
  assign sel_533149 = $signed({1'h0, add_532581}) < $signed({1'h0, sel_532583}) ? add_532581 : sel_532583;
  assign add_533151 = array_index_516863[11:0] + 12'h081;
  assign sel_533153 = $signed({1'h0, add_532585}) < $signed({1'h0, sel_532587}) ? add_532585 : sel_532587;
  assign add_533165 = array_index_517736[11:0] + 12'h0b1;
  assign sel_533167 = $signed({1'h0, add_532599}) < $signed({1'h0, sel_532601}) ? add_532599 : sel_532601;
  assign add_533169 = array_index_517739[11:0] + 12'h0b1;
  assign sel_533171 = $signed({1'h0, add_532603}) < $signed({1'h0, sel_532605}) ? add_532603 : sel_532605;
  assign add_533183 = array_index_518710[11:1] + 11'h4c1;
  assign sel_533185 = $signed({1'h0, add_532617, array_index_518210[0]}) < $signed({1'h0, sel_532619}) ? {add_532617, array_index_518210[0]} : sel_532619;
  assign add_533187 = array_index_518713[11:1] + 11'h4c1;
  assign sel_533189 = $signed({1'h0, add_532621, array_index_518213[0]}) < $signed({1'h0, sel_532623}) ? {add_532621, array_index_518213[0]} : sel_532623;
  assign add_533199 = array_index_519786[11:0] + 12'hbb1;
  assign sel_533201 = $signed({1'h0, add_532633}) < $signed({1'h0, sel_532635}) ? add_532633 : sel_532635;
  assign add_533203 = array_index_519789[11:0] + 12'hbb1;
  assign sel_533205 = $signed({1'h0, add_532637}) < $signed({1'h0, sel_532639}) ? add_532637 : sel_532639;
  assign add_533215 = array_index_520964[11:0] + 12'h6ab;
  assign sel_533217 = $signed({1'h0, add_532649}) < $signed({1'h0, sel_532651}) ? add_532649 : sel_532651;
  assign add_533219 = array_index_520967[11:0] + 12'h6ab;
  assign sel_533221 = $signed({1'h0, add_532653}) < $signed({1'h0, sel_532655}) ? add_532653 : sel_532655;
  assign sel_533232 = ($signed({1'h0, add_532285, array_index_521590[2:0]}) < $signed({1'h0, sel_532287}) ? {add_532285, array_index_521590[2:0]} : sel_532287) == ($signed({1'h0, add_532289, array_index_521593[2:0]}) < $signed({1'h0, sel_532291}) ? {add_532289, array_index_521593[2:0]} : sel_532291) ? add_533051 : sel_532868;
  assign add_533235 = array_index_513702[11:0] + 12'hcc1;
  assign sel_533237 = $signed({1'h0, add_532679}) < $signed({1'h0, sel_532681}) ? add_532679 : sel_532681;
  assign add_533239 = array_index_513705[11:0] + 12'hcc1;
  assign sel_533241 = $signed({1'h0, add_532683}) < $signed({1'h0, sel_532685}) ? add_532683 : sel_532685;
  assign add_533253 = array_index_514096[11:0] + 12'ha87;
  assign sel_533255 = $signed({1'h0, add_532697}) < $signed({1'h0, sel_532699}) ? add_532697 : sel_532699;
  assign add_533257 = array_index_514099[11:0] + 12'ha87;
  assign sel_533259 = $signed({1'h0, add_532701}) < $signed({1'h0, sel_532703}) ? add_532701 : sel_532703;
  assign add_533271 = array_index_514558[11:1] + 11'h663;
  assign sel_533273 = $signed({1'h0, add_532715, array_index_514318[0]}) < $signed({1'h0, sel_532717}) ? {add_532715, array_index_514318[0]} : sel_532717;
  assign add_533275 = array_index_514561[11:1] + 11'h663;
  assign sel_533277 = $signed({1'h0, add_532719, array_index_514321[0]}) < $signed({1'h0, sel_532721}) ? {add_532719, array_index_514321[0]} : sel_532721;
  assign add_533287 = array_index_515098[11:1] + 11'h075;
  assign sel_533289 = $signed({1'h0, add_532731, array_index_514818[0]}) < $signed({1'h0, sel_532733}) ? {add_532731, array_index_514818[0]} : sel_532733;
  assign add_533291 = array_index_515101[11:1] + 11'h075;
  assign sel_533293 = $signed({1'h0, add_532735, array_index_514821[0]}) < $signed({1'h0, sel_532737}) ? {add_532735, array_index_514821[0]} : sel_532737;
  assign add_533305 = array_index_515726[11:2] + 10'h181;
  assign sel_533307 = $signed({1'h0, add_532749, array_index_515398[1:0]}) < $signed({1'h0, sel_532751}) ? {add_532749, array_index_515398[1:0]} : sel_532751;
  assign add_533309 = array_index_515729[11:2] + 10'h181;
  assign sel_533311 = $signed({1'h0, add_532753, array_index_515401[1:0]}) < $signed({1'h0, sel_532755}) ? {add_532753, array_index_515401[1:0]} : sel_532755;
  assign add_533323 = array_index_516458[11:0] + 12'h8a7;
  assign sel_533325 = $signed({1'h0, add_532767}) < $signed({1'h0, sel_532769}) ? add_532767 : sel_532769;
  assign add_533327 = array_index_516461[11:0] + 12'h8a7;
  assign sel_533329 = $signed({1'h0, add_532771}) < $signed({1'h0, sel_532773}) ? add_532771 : sel_532773;
  assign add_533341 = array_index_517286[11:1] + 11'h283;
  assign sel_533343 = $signed({1'h0, add_532785, array_index_516860[0]}) < $signed({1'h0, sel_532787}) ? {add_532785, array_index_516860[0]} : sel_532787;
  assign add_533345 = array_index_517289[11:1] + 11'h283;
  assign sel_533347 = $signed({1'h0, add_532789, array_index_516863[0]}) < $signed({1'h0, sel_532791}) ? {add_532789, array_index_516863[0]} : sel_532791;
  assign add_533357 = array_index_518210[11:1] + 11'h44d;
  assign sel_533359 = $signed({1'h0, add_532801, array_index_517736[0]}) < $signed({1'h0, sel_532803}) ? {add_532801, array_index_517736[0]} : sel_532803;
  assign add_533361 = array_index_518213[11:1] + 11'h44d;
  assign sel_533363 = $signed({1'h0, add_532805, array_index_517739[0]}) < $signed({1'h0, sel_532807}) ? {add_532805, array_index_517739[0]} : sel_532807;
  assign add_533373 = array_index_519236[11:0] + 12'hcb1;
  assign sel_533375 = $signed({1'h0, add_532817}) < $signed({1'h0, sel_532819}) ? add_532817 : sel_532819;
  assign add_533377 = array_index_519239[11:0] + 12'hcb1;
  assign sel_533379 = $signed({1'h0, add_532821}) < $signed({1'h0, sel_532823}) ? add_532821 : sel_532823;
  assign add_533389 = array_index_520362[11:0] + 12'h81f;
  assign sel_533391 = $signed({1'h0, add_532833}) < $signed({1'h0, sel_532835}) ? add_532833 : sel_532835;
  assign add_533393 = array_index_520365[11:0] + 12'h81f;
  assign sel_533395 = $signed({1'h0, add_532837}) < $signed({1'h0, sel_532839}) ? add_532837 : sel_532839;
  assign add_533405 = array_index_521590[11:0] + 12'h45b;
  assign sel_533407 = $signed({1'h0, add_532849}) < $signed({1'h0, sel_532851}) ? add_532849 : sel_532851;
  assign add_533409 = array_index_521593[11:0] + 12'h45b;
  assign sel_533411 = $signed({1'h0, add_532853}) < $signed({1'h0, sel_532855}) ? add_532853 : sel_532855;
  assign add_533417 = sel_533232 + 16'h0001;
  assign add_533423 = array_index_513890[11:2] + 10'h113;
  assign sel_533425 = $signed({1'h0, add_532875, array_index_513702[1:0]}) < $signed({1'h0, sel_532877}) ? {add_532875, array_index_513702[1:0]} : sel_532877;
  assign add_533427 = array_index_513893[11:2] + 10'h113;
  assign sel_533429 = $signed({1'h0, add_532879, array_index_513705[1:0]}) < $signed({1'h0, sel_532881}) ? {add_532879, array_index_513705[1:0]} : sel_532881;
  assign add_533441 = array_index_514318[11:4] + 8'h49;
  assign sel_533443 = $signed({1'h0, add_532893, array_index_514096[3:0]}) < $signed({1'h0, sel_532895}) ? {add_532893, array_index_514096[3:0]} : sel_532895;
  assign add_533445 = array_index_514321[11:4] + 8'h49;
  assign sel_533447 = $signed({1'h0, add_532897, array_index_514099[3:0]}) < $signed({1'h0, sel_532899}) ? {add_532897, array_index_514099[3:0]} : sel_532899;
  assign add_533457 = array_index_514818[11:0] + 12'h263;
  assign sel_533459 = $signed({1'h0, add_532909}) < $signed({1'h0, sel_532911}) ? add_532909 : sel_532911;
  assign add_533461 = array_index_514821[11:0] + 12'h263;
  assign sel_533463 = $signed({1'h0, add_532913}) < $signed({1'h0, sel_532915}) ? add_532913 : sel_532915;
  assign add_533473 = array_index_515398[11:1] + 11'h109;
  assign sel_533475 = $signed({1'h0, add_532925, array_index_515098[0]}) < $signed({1'h0, sel_532927}) ? {add_532925, array_index_515098[0]} : sel_532927;
  assign add_533477 = array_index_515401[11:1] + 11'h109;
  assign sel_533479 = $signed({1'h0, add_532929, array_index_515101[0]}) < $signed({1'h0, sel_532931}) ? {add_532929, array_index_515101[0]} : sel_532931;
  assign add_533489 = array_index_516080[11:3] + 9'h12f;
  assign sel_533491 = $signed({1'h0, add_532941, array_index_515726[2:0]}) < $signed({1'h0, sel_532943}) ? {add_532941, array_index_515726[2:0]} : sel_532943;
  assign add_533493 = array_index_516083[11:3] + 9'h12f;
  assign sel_533495 = $signed({1'h0, add_532945, array_index_515729[2:0]}) < $signed({1'h0, sel_532947}) ? {add_532945, array_index_515729[2:0]} : sel_532947;
  assign add_533507 = array_index_516860[11:3] + 9'h171;
  assign sel_533509 = $signed({1'h0, add_532959, array_index_516458[2:0]}) < $signed({1'h0, sel_532961}) ? {add_532959, array_index_516458[2:0]} : sel_532961;
  assign add_533511 = array_index_516863[11:3] + 9'h171;
  assign sel_533513 = $signed({1'h0, add_532963, array_index_516461[2:0]}) < $signed({1'h0, sel_532965}) ? {add_532963, array_index_516461[2:0]} : sel_532965;
  assign add_533523 = array_index_517736[11:0] + 12'h091;
  assign sel_533525 = $signed({1'h0, add_532975}) < $signed({1'h0, sel_532977}) ? add_532975 : sel_532977;
  assign add_533527 = array_index_517739[11:0] + 12'h091;
  assign sel_533529 = $signed({1'h0, add_532979}) < $signed({1'h0, sel_532981}) ? add_532979 : sel_532981;
  assign add_533539 = array_index_518710[11:0] + 12'hf59;
  assign sel_533541 = $signed({1'h0, add_532991}) < $signed({1'h0, sel_532993}) ? add_532991 : sel_532993;
  assign add_533543 = array_index_518713[11:0] + 12'hf59;
  assign sel_533545 = $signed({1'h0, add_532995}) < $signed({1'h0, sel_532997}) ? add_532995 : sel_532997;
  assign add_533557 = array_index_519786[11:0] + 12'h437;
  assign sel_533559 = $signed({1'h0, add_533009}) < $signed({1'h0, sel_533011}) ? add_533009 : sel_533011;
  assign add_533561 = array_index_519789[11:0] + 12'h437;
  assign sel_533563 = $signed({1'h0, add_533013}) < $signed({1'h0, sel_533015}) ? add_533013 : sel_533015;
  assign add_533573 = array_index_520964[11:0] + 12'hee1;
  assign sel_533575 = $signed({1'h0, add_533025}) < $signed({1'h0, sel_533027}) ? add_533025 : sel_533027;
  assign add_533577 = array_index_520967[11:0] + 12'hee1;
  assign sel_533579 = $signed({1'h0, add_533029}) < $signed({1'h0, sel_533031}) ? add_533029 : sel_533031;
  assign sel_533590 = ($signed({1'h0, add_532665}) < $signed({1'h0, sel_532667}) ? add_532665 : sel_532667) == ($signed({1'h0, add_532669}) < $signed({1'h0, sel_532671}) ? add_532669 : sel_532671) ? add_533417 : sel_533232;
  assign add_533601 = array_index_514096[11:1] + 11'h5b9;
  assign sel_533603 = $signed({1'h0, add_533061, array_index_513890[0]}) < $signed({1'h0, sel_533063}) ? {add_533061, array_index_513890[0]} : sel_533063;
  assign add_533605 = array_index_514099[11:1] + 11'h5b9;
  assign sel_533607 = $signed({1'h0, add_533065, array_index_513893[0]}) < $signed({1'h0, sel_533067}) ? {add_533065, array_index_513893[0]} : sel_533067;
  assign add_533617 = array_index_514558[11:0] + 12'h37b;
  assign sel_533619 = $signed({1'h0, add_533077}) < $signed({1'h0, sel_533079}) ? add_533077 : sel_533079;
  assign add_533621 = array_index_514561[11:0] + 12'h37b;
  assign sel_533623 = $signed({1'h0, add_533081}) < $signed({1'h0, sel_533083}) ? add_533081 : sel_533083;
  assign add_533635 = array_index_515098[11:0] + 12'h811;
  assign sel_533637 = $signed({1'h0, add_533095}) < $signed({1'h0, sel_533097}) ? add_533095 : sel_533097;
  assign add_533639 = array_index_515101[11:0] + 12'h811;
  assign sel_533641 = $signed({1'h0, add_533099}) < $signed({1'h0, sel_533101}) ? add_533099 : sel_533101;
  assign add_533653 = array_index_515726[11:0] + 12'h70f;
  assign sel_533655 = $signed({1'h0, add_533113}) < $signed({1'h0, sel_533115}) ? add_533113 : sel_533115;
  assign add_533657 = array_index_515729[11:0] + 12'h70f;
  assign sel_533659 = $signed({1'h0, add_533117}) < $signed({1'h0, sel_533119}) ? add_533117 : sel_533119;
  assign add_533671 = array_index_516458[11:3] + 9'h1f1;
  assign sel_533673 = $signed({1'h0, add_533131, array_index_516080[2:0]}) < $signed({1'h0, sel_533133}) ? {add_533131, array_index_516080[2:0]} : sel_533133;
  assign add_533675 = array_index_516461[11:3] + 9'h1f1;
  assign sel_533677 = $signed({1'h0, add_533135, array_index_516083[2:0]}) < $signed({1'h0, sel_533137}) ? {add_533135, array_index_516083[2:0]} : sel_533137;
  assign add_533687 = array_index_517286[11:0] + 12'h081;
  assign sel_533689 = $signed({1'h0, add_533147}) < $signed({1'h0, sel_533149}) ? add_533147 : sel_533149;
  assign add_533691 = array_index_517289[11:0] + 12'h081;
  assign sel_533693 = $signed({1'h0, add_533151}) < $signed({1'h0, sel_533153}) ? add_533151 : sel_533153;
  assign add_533705 = array_index_518210[11:0] + 12'h0b1;
  assign sel_533707 = $signed({1'h0, add_533165}) < $signed({1'h0, sel_533167}) ? add_533165 : sel_533167;
  assign add_533709 = array_index_518213[11:0] + 12'h0b1;
  assign sel_533711 = $signed({1'h0, add_533169}) < $signed({1'h0, sel_533171}) ? add_533169 : sel_533171;
  assign add_533723 = array_index_519236[11:1] + 11'h4c1;
  assign sel_533725 = $signed({1'h0, add_533183, array_index_518710[0]}) < $signed({1'h0, sel_533185}) ? {add_533183, array_index_518710[0]} : sel_533185;
  assign add_533727 = array_index_519239[11:1] + 11'h4c1;
  assign sel_533729 = $signed({1'h0, add_533187, array_index_518713[0]}) < $signed({1'h0, sel_533189}) ? {add_533187, array_index_518713[0]} : sel_533189;
  assign add_533739 = array_index_520362[11:0] + 12'hbb1;
  assign sel_533741 = $signed({1'h0, add_533199}) < $signed({1'h0, sel_533201}) ? add_533199 : sel_533201;
  assign add_533743 = array_index_520365[11:0] + 12'hbb1;
  assign sel_533745 = $signed({1'h0, add_533203}) < $signed({1'h0, sel_533205}) ? add_533203 : sel_533205;
  assign add_533755 = array_index_521590[11:0] + 12'h6ab;
  assign sel_533757 = $signed({1'h0, add_533215}) < $signed({1'h0, sel_533217}) ? add_533215 : sel_533217;
  assign add_533759 = array_index_521593[11:0] + 12'h6ab;
  assign sel_533761 = $signed({1'h0, add_533219}) < $signed({1'h0, sel_533221}) ? add_533219 : sel_533221;
  assign add_533765 = sel_533590 + 16'h0001;
  assign add_533767 = array_index_513890[11:0] + 12'hcc1;
  assign sel_533769 = $signed({1'h0, add_533235}) < $signed({1'h0, sel_533237}) ? add_533235 : sel_533237;
  assign add_533771 = array_index_513893[11:0] + 12'hcc1;
  assign sel_533773 = $signed({1'h0, add_533239}) < $signed({1'h0, sel_533241}) ? add_533239 : sel_533241;
  assign add_533785 = array_index_514318[11:0] + 12'ha87;
  assign sel_533787 = $signed({1'h0, add_533253}) < $signed({1'h0, sel_533255}) ? add_533253 : sel_533255;
  assign add_533789 = array_index_514321[11:0] + 12'ha87;
  assign sel_533791 = $signed({1'h0, add_533257}) < $signed({1'h0, sel_533259}) ? add_533257 : sel_533259;
  assign add_533803 = array_index_514818[11:1] + 11'h663;
  assign sel_533805 = $signed({1'h0, add_533271, array_index_514558[0]}) < $signed({1'h0, sel_533273}) ? {add_533271, array_index_514558[0]} : sel_533273;
  assign add_533807 = array_index_514821[11:1] + 11'h663;
  assign sel_533809 = $signed({1'h0, add_533275, array_index_514561[0]}) < $signed({1'h0, sel_533277}) ? {add_533275, array_index_514561[0]} : sel_533277;
  assign add_533819 = array_index_515398[11:1] + 11'h075;
  assign sel_533821 = $signed({1'h0, add_533287, array_index_515098[0]}) < $signed({1'h0, sel_533289}) ? {add_533287, array_index_515098[0]} : sel_533289;
  assign add_533823 = array_index_515401[11:1] + 11'h075;
  assign sel_533825 = $signed({1'h0, add_533291, array_index_515101[0]}) < $signed({1'h0, sel_533293}) ? {add_533291, array_index_515101[0]} : sel_533293;
  assign add_533837 = array_index_516080[11:2] + 10'h181;
  assign sel_533839 = $signed({1'h0, add_533305, array_index_515726[1:0]}) < $signed({1'h0, sel_533307}) ? {add_533305, array_index_515726[1:0]} : sel_533307;
  assign add_533841 = array_index_516083[11:2] + 10'h181;
  assign sel_533843 = $signed({1'h0, add_533309, array_index_515729[1:0]}) < $signed({1'h0, sel_533311}) ? {add_533309, array_index_515729[1:0]} : sel_533311;
  assign add_533855 = array_index_516860[11:0] + 12'h8a7;
  assign sel_533857 = $signed({1'h0, add_533323}) < $signed({1'h0, sel_533325}) ? add_533323 : sel_533325;
  assign add_533859 = array_index_516863[11:0] + 12'h8a7;
  assign sel_533861 = $signed({1'h0, add_533327}) < $signed({1'h0, sel_533329}) ? add_533327 : sel_533329;
  assign add_533873 = array_index_517736[11:1] + 11'h283;
  assign sel_533875 = $signed({1'h0, add_533341, array_index_517286[0]}) < $signed({1'h0, sel_533343}) ? {add_533341, array_index_517286[0]} : sel_533343;
  assign add_533877 = array_index_517739[11:1] + 11'h283;
  assign sel_533879 = $signed({1'h0, add_533345, array_index_517289[0]}) < $signed({1'h0, sel_533347}) ? {add_533345, array_index_517289[0]} : sel_533347;
  assign add_533889 = array_index_518710[11:1] + 11'h44d;
  assign sel_533891 = $signed({1'h0, add_533357, array_index_518210[0]}) < $signed({1'h0, sel_533359}) ? {add_533357, array_index_518210[0]} : sel_533359;
  assign add_533893 = array_index_518713[11:1] + 11'h44d;
  assign sel_533895 = $signed({1'h0, add_533361, array_index_518213[0]}) < $signed({1'h0, sel_533363}) ? {add_533361, array_index_518213[0]} : sel_533363;
  assign add_533905 = array_index_519786[11:0] + 12'hcb1;
  assign sel_533907 = $signed({1'h0, add_533373}) < $signed({1'h0, sel_533375}) ? add_533373 : sel_533375;
  assign add_533909 = array_index_519789[11:0] + 12'hcb1;
  assign sel_533911 = $signed({1'h0, add_533377}) < $signed({1'h0, sel_533379}) ? add_533377 : sel_533379;
  assign add_533921 = array_index_520964[11:0] + 12'h81f;
  assign sel_533923 = $signed({1'h0, add_533389}) < $signed({1'h0, sel_533391}) ? add_533389 : sel_533391;
  assign add_533925 = array_index_520967[11:0] + 12'h81f;
  assign sel_533927 = $signed({1'h0, add_533393}) < $signed({1'h0, sel_533395}) ? add_533393 : sel_533395;
  assign sel_533938 = ($signed({1'h0, add_533041, array_index_521590[0]}) < $signed({1'h0, sel_533043}) ? {add_533041, array_index_521590[0]} : sel_533043) == ($signed({1'h0, add_533045, array_index_521593[0]}) < $signed({1'h0, sel_533047}) ? {add_533045, array_index_521593[0]} : sel_533047) ? add_533765 : sel_533590;
  assign add_533945 = array_index_514096[11:2] + 10'h113;
  assign sel_533947 = $signed({1'h0, add_533423, array_index_513890[1:0]}) < $signed({1'h0, sel_533425}) ? {add_533423, array_index_513890[1:0]} : sel_533425;
  assign add_533949 = array_index_514099[11:2] + 10'h113;
  assign sel_533951 = $signed({1'h0, add_533427, array_index_513893[1:0]}) < $signed({1'h0, sel_533429}) ? {add_533427, array_index_513893[1:0]} : sel_533429;
  assign add_533963 = array_index_514558[11:4] + 8'h49;
  assign sel_533965 = $signed({1'h0, add_533441, array_index_514318[3:0]}) < $signed({1'h0, sel_533443}) ? {add_533441, array_index_514318[3:0]} : sel_533443;
  assign add_533967 = array_index_514561[11:4] + 8'h49;
  assign sel_533969 = $signed({1'h0, add_533445, array_index_514321[3:0]}) < $signed({1'h0, sel_533447}) ? {add_533445, array_index_514321[3:0]} : sel_533447;
  assign add_533979 = array_index_515098[11:0] + 12'h263;
  assign sel_533981 = $signed({1'h0, add_533457}) < $signed({1'h0, sel_533459}) ? add_533457 : sel_533459;
  assign add_533983 = array_index_515101[11:0] + 12'h263;
  assign sel_533985 = $signed({1'h0, add_533461}) < $signed({1'h0, sel_533463}) ? add_533461 : sel_533463;
  assign add_533995 = array_index_515726[11:1] + 11'h109;
  assign sel_533997 = $signed({1'h0, add_533473, array_index_515398[0]}) < $signed({1'h0, sel_533475}) ? {add_533473, array_index_515398[0]} : sel_533475;
  assign add_533999 = array_index_515729[11:1] + 11'h109;
  assign sel_534001 = $signed({1'h0, add_533477, array_index_515401[0]}) < $signed({1'h0, sel_533479}) ? {add_533477, array_index_515401[0]} : sel_533479;
  assign add_534011 = array_index_516458[11:3] + 9'h12f;
  assign sel_534013 = $signed({1'h0, add_533489, array_index_516080[2:0]}) < $signed({1'h0, sel_533491}) ? {add_533489, array_index_516080[2:0]} : sel_533491;
  assign add_534015 = array_index_516461[11:3] + 9'h12f;
  assign sel_534017 = $signed({1'h0, add_533493, array_index_516083[2:0]}) < $signed({1'h0, sel_533495}) ? {add_533493, array_index_516083[2:0]} : sel_533495;
  assign add_534029 = array_index_517286[11:3] + 9'h171;
  assign sel_534031 = $signed({1'h0, add_533507, array_index_516860[2:0]}) < $signed({1'h0, sel_533509}) ? {add_533507, array_index_516860[2:0]} : sel_533509;
  assign add_534033 = array_index_517289[11:3] + 9'h171;
  assign sel_534035 = $signed({1'h0, add_533511, array_index_516863[2:0]}) < $signed({1'h0, sel_533513}) ? {add_533511, array_index_516863[2:0]} : sel_533513;
  assign add_534045 = array_index_518210[11:0] + 12'h091;
  assign sel_534047 = $signed({1'h0, add_533523}) < $signed({1'h0, sel_533525}) ? add_533523 : sel_533525;
  assign add_534049 = array_index_518213[11:0] + 12'h091;
  assign sel_534051 = $signed({1'h0, add_533527}) < $signed({1'h0, sel_533529}) ? add_533527 : sel_533529;
  assign add_534061 = array_index_519236[11:0] + 12'hf59;
  assign sel_534063 = $signed({1'h0, add_533539}) < $signed({1'h0, sel_533541}) ? add_533539 : sel_533541;
  assign add_534065 = array_index_519239[11:0] + 12'hf59;
  assign sel_534067 = $signed({1'h0, add_533543}) < $signed({1'h0, sel_533545}) ? add_533543 : sel_533545;
  assign add_534079 = array_index_520362[11:0] + 12'h437;
  assign sel_534081 = $signed({1'h0, add_533557}) < $signed({1'h0, sel_533559}) ? add_533557 : sel_533559;
  assign add_534083 = array_index_520365[11:0] + 12'h437;
  assign sel_534085 = $signed({1'h0, add_533561}) < $signed({1'h0, sel_533563}) ? add_533561 : sel_533563;
  assign add_534095 = array_index_521590[11:0] + 12'hee1;
  assign sel_534097 = $signed({1'h0, add_533573}) < $signed({1'h0, sel_533575}) ? add_533573 : sel_533575;
  assign add_534099 = array_index_521593[11:0] + 12'hee1;
  assign sel_534101 = $signed({1'h0, add_533577}) < $signed({1'h0, sel_533579}) ? add_533577 : sel_533579;
  assign add_534105 = sel_533938 + 16'h0001;
  assign add_534115 = array_index_514318[11:1] + 11'h5b9;
  assign sel_534117 = $signed({1'h0, add_533601, array_index_514096[0]}) < $signed({1'h0, sel_533603}) ? {add_533601, array_index_514096[0]} : sel_533603;
  assign add_534119 = array_index_514321[11:1] + 11'h5b9;
  assign sel_534121 = $signed({1'h0, add_533605, array_index_514099[0]}) < $signed({1'h0, sel_533607}) ? {add_533605, array_index_514099[0]} : sel_533607;
  assign add_534131 = array_index_514818[11:0] + 12'h37b;
  assign sel_534133 = $signed({1'h0, add_533617}) < $signed({1'h0, sel_533619}) ? add_533617 : sel_533619;
  assign add_534135 = array_index_514821[11:0] + 12'h37b;
  assign sel_534137 = $signed({1'h0, add_533621}) < $signed({1'h0, sel_533623}) ? add_533621 : sel_533623;
  assign add_534149 = array_index_515398[11:0] + 12'h811;
  assign sel_534151 = $signed({1'h0, add_533635}) < $signed({1'h0, sel_533637}) ? add_533635 : sel_533637;
  assign add_534153 = array_index_515401[11:0] + 12'h811;
  assign sel_534155 = $signed({1'h0, add_533639}) < $signed({1'h0, sel_533641}) ? add_533639 : sel_533641;
  assign add_534167 = array_index_516080[11:0] + 12'h70f;
  assign sel_534169 = $signed({1'h0, add_533653}) < $signed({1'h0, sel_533655}) ? add_533653 : sel_533655;
  assign add_534171 = array_index_516083[11:0] + 12'h70f;
  assign sel_534173 = $signed({1'h0, add_533657}) < $signed({1'h0, sel_533659}) ? add_533657 : sel_533659;
  assign add_534185 = array_index_516860[11:3] + 9'h1f1;
  assign sel_534187 = $signed({1'h0, add_533671, array_index_516458[2:0]}) < $signed({1'h0, sel_533673}) ? {add_533671, array_index_516458[2:0]} : sel_533673;
  assign add_534189 = array_index_516863[11:3] + 9'h1f1;
  assign sel_534191 = $signed({1'h0, add_533675, array_index_516461[2:0]}) < $signed({1'h0, sel_533677}) ? {add_533675, array_index_516461[2:0]} : sel_533677;
  assign add_534201 = array_index_517736[11:0] + 12'h081;
  assign sel_534203 = $signed({1'h0, add_533687}) < $signed({1'h0, sel_533689}) ? add_533687 : sel_533689;
  assign add_534205 = array_index_517739[11:0] + 12'h081;
  assign sel_534207 = $signed({1'h0, add_533691}) < $signed({1'h0, sel_533693}) ? add_533691 : sel_533693;
  assign add_534219 = array_index_518710[11:0] + 12'h0b1;
  assign sel_534221 = $signed({1'h0, add_533705}) < $signed({1'h0, sel_533707}) ? add_533705 : sel_533707;
  assign add_534223 = array_index_518713[11:0] + 12'h0b1;
  assign sel_534225 = $signed({1'h0, add_533709}) < $signed({1'h0, sel_533711}) ? add_533709 : sel_533711;
  assign add_534237 = array_index_519786[11:1] + 11'h4c1;
  assign sel_534239 = $signed({1'h0, add_533723, array_index_519236[0]}) < $signed({1'h0, sel_533725}) ? {add_533723, array_index_519236[0]} : sel_533725;
  assign add_534241 = array_index_519789[11:1] + 11'h4c1;
  assign sel_534243 = $signed({1'h0, add_533727, array_index_519239[0]}) < $signed({1'h0, sel_533729}) ? {add_533727, array_index_519239[0]} : sel_533729;
  assign add_534253 = array_index_520964[11:0] + 12'hbb1;
  assign sel_534255 = $signed({1'h0, add_533739}) < $signed({1'h0, sel_533741}) ? add_533739 : sel_533741;
  assign add_534257 = array_index_520967[11:0] + 12'hbb1;
  assign sel_534259 = $signed({1'h0, add_533743}) < $signed({1'h0, sel_533745}) ? add_533743 : sel_533745;
  assign sel_534270 = ($signed({1'h0, add_533405}) < $signed({1'h0, sel_533407}) ? add_533405 : sel_533407) == ($signed({1'h0, add_533409}) < $signed({1'h0, sel_533411}) ? add_533409 : sel_533411) ? add_534105 : sel_533938;
  assign add_534273 = array_index_514096[11:0] + 12'hcc1;
  assign sel_534275 = $signed({1'h0, add_533767}) < $signed({1'h0, sel_533769}) ? add_533767 : sel_533769;
  assign add_534277 = array_index_514099[11:0] + 12'hcc1;
  assign sel_534279 = $signed({1'h0, add_533771}) < $signed({1'h0, sel_533773}) ? add_533771 : sel_533773;
  assign add_534291 = array_index_514558[11:0] + 12'ha87;
  assign sel_534293 = $signed({1'h0, add_533785}) < $signed({1'h0, sel_533787}) ? add_533785 : sel_533787;
  assign add_534295 = array_index_514561[11:0] + 12'ha87;
  assign sel_534297 = $signed({1'h0, add_533789}) < $signed({1'h0, sel_533791}) ? add_533789 : sel_533791;
  assign add_534309 = array_index_515098[11:1] + 11'h663;
  assign sel_534311 = $signed({1'h0, add_533803, array_index_514818[0]}) < $signed({1'h0, sel_533805}) ? {add_533803, array_index_514818[0]} : sel_533805;
  assign add_534313 = array_index_515101[11:1] + 11'h663;
  assign sel_534315 = $signed({1'h0, add_533807, array_index_514821[0]}) < $signed({1'h0, sel_533809}) ? {add_533807, array_index_514821[0]} : sel_533809;
  assign add_534325 = array_index_515726[11:1] + 11'h075;
  assign sel_534327 = $signed({1'h0, add_533819, array_index_515398[0]}) < $signed({1'h0, sel_533821}) ? {add_533819, array_index_515398[0]} : sel_533821;
  assign add_534329 = array_index_515729[11:1] + 11'h075;
  assign sel_534331 = $signed({1'h0, add_533823, array_index_515401[0]}) < $signed({1'h0, sel_533825}) ? {add_533823, array_index_515401[0]} : sel_533825;
  assign add_534343 = array_index_516458[11:2] + 10'h181;
  assign sel_534345 = $signed({1'h0, add_533837, array_index_516080[1:0]}) < $signed({1'h0, sel_533839}) ? {add_533837, array_index_516080[1:0]} : sel_533839;
  assign add_534347 = array_index_516461[11:2] + 10'h181;
  assign sel_534349 = $signed({1'h0, add_533841, array_index_516083[1:0]}) < $signed({1'h0, sel_533843}) ? {add_533841, array_index_516083[1:0]} : sel_533843;
  assign add_534361 = array_index_517286[11:0] + 12'h8a7;
  assign sel_534363 = $signed({1'h0, add_533855}) < $signed({1'h0, sel_533857}) ? add_533855 : sel_533857;
  assign add_534365 = array_index_517289[11:0] + 12'h8a7;
  assign sel_534367 = $signed({1'h0, add_533859}) < $signed({1'h0, sel_533861}) ? add_533859 : sel_533861;
  assign add_534379 = array_index_518210[11:1] + 11'h283;
  assign sel_534381 = $signed({1'h0, add_533873, array_index_517736[0]}) < $signed({1'h0, sel_533875}) ? {add_533873, array_index_517736[0]} : sel_533875;
  assign add_534383 = array_index_518213[11:1] + 11'h283;
  assign sel_534385 = $signed({1'h0, add_533877, array_index_517739[0]}) < $signed({1'h0, sel_533879}) ? {add_533877, array_index_517739[0]} : sel_533879;
  assign add_534395 = array_index_519236[11:1] + 11'h44d;
  assign sel_534397 = $signed({1'h0, add_533889, array_index_518710[0]}) < $signed({1'h0, sel_533891}) ? {add_533889, array_index_518710[0]} : sel_533891;
  assign add_534399 = array_index_519239[11:1] + 11'h44d;
  assign sel_534401 = $signed({1'h0, add_533893, array_index_518713[0]}) < $signed({1'h0, sel_533895}) ? {add_533893, array_index_518713[0]} : sel_533895;
  assign add_534411 = array_index_520362[11:0] + 12'hcb1;
  assign sel_534413 = $signed({1'h0, add_533905}) < $signed({1'h0, sel_533907}) ? add_533905 : sel_533907;
  assign add_534415 = array_index_520365[11:0] + 12'hcb1;
  assign sel_534417 = $signed({1'h0, add_533909}) < $signed({1'h0, sel_533911}) ? add_533909 : sel_533911;
  assign add_534427 = array_index_521590[11:0] + 12'h81f;
  assign sel_534429 = $signed({1'h0, add_533921}) < $signed({1'h0, sel_533923}) ? add_533921 : sel_533923;
  assign add_534431 = array_index_521593[11:0] + 12'h81f;
  assign sel_534433 = $signed({1'h0, add_533925}) < $signed({1'h0, sel_533927}) ? add_533925 : sel_533927;
  assign add_534437 = sel_534270 + 16'h0001;
  assign add_534443 = array_index_514318[11:2] + 10'h113;
  assign sel_534445 = $signed({1'h0, add_533945, array_index_514096[1:0]}) < $signed({1'h0, sel_533947}) ? {add_533945, array_index_514096[1:0]} : sel_533947;
  assign add_534447 = array_index_514321[11:2] + 10'h113;
  assign sel_534449 = $signed({1'h0, add_533949, array_index_514099[1:0]}) < $signed({1'h0, sel_533951}) ? {add_533949, array_index_514099[1:0]} : sel_533951;
  assign add_534461 = array_index_514818[11:4] + 8'h49;
  assign sel_534463 = $signed({1'h0, add_533963, array_index_514558[3:0]}) < $signed({1'h0, sel_533965}) ? {add_533963, array_index_514558[3:0]} : sel_533965;
  assign add_534465 = array_index_514821[11:4] + 8'h49;
  assign sel_534467 = $signed({1'h0, add_533967, array_index_514561[3:0]}) < $signed({1'h0, sel_533969}) ? {add_533967, array_index_514561[3:0]} : sel_533969;
  assign add_534477 = array_index_515398[11:0] + 12'h263;
  assign sel_534479 = $signed({1'h0, add_533979}) < $signed({1'h0, sel_533981}) ? add_533979 : sel_533981;
  assign add_534481 = array_index_515401[11:0] + 12'h263;
  assign sel_534483 = $signed({1'h0, add_533983}) < $signed({1'h0, sel_533985}) ? add_533983 : sel_533985;
  assign add_534493 = array_index_516080[11:1] + 11'h109;
  assign sel_534495 = $signed({1'h0, add_533995, array_index_515726[0]}) < $signed({1'h0, sel_533997}) ? {add_533995, array_index_515726[0]} : sel_533997;
  assign add_534497 = array_index_516083[11:1] + 11'h109;
  assign sel_534499 = $signed({1'h0, add_533999, array_index_515729[0]}) < $signed({1'h0, sel_534001}) ? {add_533999, array_index_515729[0]} : sel_534001;
  assign add_534509 = array_index_516860[11:3] + 9'h12f;
  assign sel_534511 = $signed({1'h0, add_534011, array_index_516458[2:0]}) < $signed({1'h0, sel_534013}) ? {add_534011, array_index_516458[2:0]} : sel_534013;
  assign add_534513 = array_index_516863[11:3] + 9'h12f;
  assign sel_534515 = $signed({1'h0, add_534015, array_index_516461[2:0]}) < $signed({1'h0, sel_534017}) ? {add_534015, array_index_516461[2:0]} : sel_534017;
  assign add_534527 = array_index_517736[11:3] + 9'h171;
  assign sel_534529 = $signed({1'h0, add_534029, array_index_517286[2:0]}) < $signed({1'h0, sel_534031}) ? {add_534029, array_index_517286[2:0]} : sel_534031;
  assign add_534531 = array_index_517739[11:3] + 9'h171;
  assign sel_534533 = $signed({1'h0, add_534033, array_index_517289[2:0]}) < $signed({1'h0, sel_534035}) ? {add_534033, array_index_517289[2:0]} : sel_534035;
  assign add_534543 = array_index_518710[11:0] + 12'h091;
  assign sel_534545 = $signed({1'h0, add_534045}) < $signed({1'h0, sel_534047}) ? add_534045 : sel_534047;
  assign add_534547 = array_index_518713[11:0] + 12'h091;
  assign sel_534549 = $signed({1'h0, add_534049}) < $signed({1'h0, sel_534051}) ? add_534049 : sel_534051;
  assign add_534559 = array_index_519786[11:0] + 12'hf59;
  assign sel_534561 = $signed({1'h0, add_534061}) < $signed({1'h0, sel_534063}) ? add_534061 : sel_534063;
  assign add_534563 = array_index_519789[11:0] + 12'hf59;
  assign sel_534565 = $signed({1'h0, add_534065}) < $signed({1'h0, sel_534067}) ? add_534065 : sel_534067;
  assign add_534577 = array_index_520964[11:0] + 12'h437;
  assign sel_534579 = $signed({1'h0, add_534079}) < $signed({1'h0, sel_534081}) ? add_534079 : sel_534081;
  assign add_534581 = array_index_520967[11:0] + 12'h437;
  assign sel_534583 = $signed({1'h0, add_534083}) < $signed({1'h0, sel_534085}) ? add_534083 : sel_534085;
  assign sel_534594 = ($signed({1'h0, add_533755}) < $signed({1'h0, sel_533757}) ? add_533755 : sel_533757) == ($signed({1'h0, add_533759}) < $signed({1'h0, sel_533761}) ? add_533759 : sel_533761) ? add_534437 : sel_534270;
  assign add_534605 = array_index_514558[11:1] + 11'h5b9;
  assign sel_534607 = $signed({1'h0, add_534115, array_index_514318[0]}) < $signed({1'h0, sel_534117}) ? {add_534115, array_index_514318[0]} : sel_534117;
  assign add_534609 = array_index_514561[11:1] + 11'h5b9;
  assign sel_534611 = $signed({1'h0, add_534119, array_index_514321[0]}) < $signed({1'h0, sel_534121}) ? {add_534119, array_index_514321[0]} : sel_534121;
  assign add_534621 = array_index_515098[11:0] + 12'h37b;
  assign sel_534623 = $signed({1'h0, add_534131}) < $signed({1'h0, sel_534133}) ? add_534131 : sel_534133;
  assign add_534625 = array_index_515101[11:0] + 12'h37b;
  assign sel_534627 = $signed({1'h0, add_534135}) < $signed({1'h0, sel_534137}) ? add_534135 : sel_534137;
  assign add_534639 = array_index_515726[11:0] + 12'h811;
  assign sel_534641 = $signed({1'h0, add_534149}) < $signed({1'h0, sel_534151}) ? add_534149 : sel_534151;
  assign add_534643 = array_index_515729[11:0] + 12'h811;
  assign sel_534645 = $signed({1'h0, add_534153}) < $signed({1'h0, sel_534155}) ? add_534153 : sel_534155;
  assign add_534657 = array_index_516458[11:0] + 12'h70f;
  assign sel_534659 = $signed({1'h0, add_534167}) < $signed({1'h0, sel_534169}) ? add_534167 : sel_534169;
  assign add_534661 = array_index_516461[11:0] + 12'h70f;
  assign sel_534663 = $signed({1'h0, add_534171}) < $signed({1'h0, sel_534173}) ? add_534171 : sel_534173;
  assign add_534675 = array_index_517286[11:3] + 9'h1f1;
  assign sel_534677 = $signed({1'h0, add_534185, array_index_516860[2:0]}) < $signed({1'h0, sel_534187}) ? {add_534185, array_index_516860[2:0]} : sel_534187;
  assign add_534679 = array_index_517289[11:3] + 9'h1f1;
  assign sel_534681 = $signed({1'h0, add_534189, array_index_516863[2:0]}) < $signed({1'h0, sel_534191}) ? {add_534189, array_index_516863[2:0]} : sel_534191;
  assign add_534691 = array_index_518210[11:0] + 12'h081;
  assign sel_534693 = $signed({1'h0, add_534201}) < $signed({1'h0, sel_534203}) ? add_534201 : sel_534203;
  assign add_534695 = array_index_518213[11:0] + 12'h081;
  assign sel_534697 = $signed({1'h0, add_534205}) < $signed({1'h0, sel_534207}) ? add_534205 : sel_534207;
  assign add_534709 = array_index_519236[11:0] + 12'h0b1;
  assign sel_534711 = $signed({1'h0, add_534219}) < $signed({1'h0, sel_534221}) ? add_534219 : sel_534221;
  assign add_534713 = array_index_519239[11:0] + 12'h0b1;
  assign sel_534715 = $signed({1'h0, add_534223}) < $signed({1'h0, sel_534225}) ? add_534223 : sel_534225;
  assign add_534727 = array_index_520362[11:1] + 11'h4c1;
  assign sel_534729 = $signed({1'h0, add_534237, array_index_519786[0]}) < $signed({1'h0, sel_534239}) ? {add_534237, array_index_519786[0]} : sel_534239;
  assign add_534731 = array_index_520365[11:1] + 11'h4c1;
  assign sel_534733 = $signed({1'h0, add_534241, array_index_519789[0]}) < $signed({1'h0, sel_534243}) ? {add_534241, array_index_519789[0]} : sel_534243;
  assign add_534743 = array_index_521590[11:0] + 12'hbb1;
  assign sel_534745 = $signed({1'h0, add_534253}) < $signed({1'h0, sel_534255}) ? add_534253 : sel_534255;
  assign add_534747 = array_index_521593[11:0] + 12'hbb1;
  assign sel_534749 = $signed({1'h0, add_534257}) < $signed({1'h0, sel_534259}) ? add_534257 : sel_534259;
  assign add_534753 = sel_534594 + 16'h0001;
  assign add_534755 = array_index_514318[11:0] + 12'hcc1;
  assign sel_534757 = $signed({1'h0, add_534273}) < $signed({1'h0, sel_534275}) ? add_534273 : sel_534275;
  assign add_534759 = array_index_514321[11:0] + 12'hcc1;
  assign sel_534761 = $signed({1'h0, add_534277}) < $signed({1'h0, sel_534279}) ? add_534277 : sel_534279;
  assign add_534773 = array_index_514818[11:0] + 12'ha87;
  assign sel_534775 = $signed({1'h0, add_534291}) < $signed({1'h0, sel_534293}) ? add_534291 : sel_534293;
  assign add_534777 = array_index_514821[11:0] + 12'ha87;
  assign sel_534779 = $signed({1'h0, add_534295}) < $signed({1'h0, sel_534297}) ? add_534295 : sel_534297;
  assign add_534791 = array_index_515398[11:1] + 11'h663;
  assign sel_534793 = $signed({1'h0, add_534309, array_index_515098[0]}) < $signed({1'h0, sel_534311}) ? {add_534309, array_index_515098[0]} : sel_534311;
  assign add_534795 = array_index_515401[11:1] + 11'h663;
  assign sel_534797 = $signed({1'h0, add_534313, array_index_515101[0]}) < $signed({1'h0, sel_534315}) ? {add_534313, array_index_515101[0]} : sel_534315;
  assign add_534807 = array_index_516080[11:1] + 11'h075;
  assign sel_534809 = $signed({1'h0, add_534325, array_index_515726[0]}) < $signed({1'h0, sel_534327}) ? {add_534325, array_index_515726[0]} : sel_534327;
  assign add_534811 = array_index_516083[11:1] + 11'h075;
  assign sel_534813 = $signed({1'h0, add_534329, array_index_515729[0]}) < $signed({1'h0, sel_534331}) ? {add_534329, array_index_515729[0]} : sel_534331;
  assign add_534825 = array_index_516860[11:2] + 10'h181;
  assign sel_534827 = $signed({1'h0, add_534343, array_index_516458[1:0]}) < $signed({1'h0, sel_534345}) ? {add_534343, array_index_516458[1:0]} : sel_534345;
  assign add_534829 = array_index_516863[11:2] + 10'h181;
  assign sel_534831 = $signed({1'h0, add_534347, array_index_516461[1:0]}) < $signed({1'h0, sel_534349}) ? {add_534347, array_index_516461[1:0]} : sel_534349;
  assign add_534843 = array_index_517736[11:0] + 12'h8a7;
  assign sel_534845 = $signed({1'h0, add_534361}) < $signed({1'h0, sel_534363}) ? add_534361 : sel_534363;
  assign add_534847 = array_index_517739[11:0] + 12'h8a7;
  assign sel_534849 = $signed({1'h0, add_534365}) < $signed({1'h0, sel_534367}) ? add_534365 : sel_534367;
  assign add_534861 = array_index_518710[11:1] + 11'h283;
  assign sel_534863 = $signed({1'h0, add_534379, array_index_518210[0]}) < $signed({1'h0, sel_534381}) ? {add_534379, array_index_518210[0]} : sel_534381;
  assign add_534865 = array_index_518713[11:1] + 11'h283;
  assign sel_534867 = $signed({1'h0, add_534383, array_index_518213[0]}) < $signed({1'h0, sel_534385}) ? {add_534383, array_index_518213[0]} : sel_534385;
  assign add_534877 = array_index_519786[11:1] + 11'h44d;
  assign sel_534879 = $signed({1'h0, add_534395, array_index_519236[0]}) < $signed({1'h0, sel_534397}) ? {add_534395, array_index_519236[0]} : sel_534397;
  assign add_534881 = array_index_519789[11:1] + 11'h44d;
  assign sel_534883 = $signed({1'h0, add_534399, array_index_519239[0]}) < $signed({1'h0, sel_534401}) ? {add_534399, array_index_519239[0]} : sel_534401;
  assign add_534893 = array_index_520964[11:0] + 12'hcb1;
  assign sel_534895 = $signed({1'h0, add_534411}) < $signed({1'h0, sel_534413}) ? add_534411 : sel_534413;
  assign add_534897 = array_index_520967[11:0] + 12'hcb1;
  assign sel_534899 = $signed({1'h0, add_534415}) < $signed({1'h0, sel_534417}) ? add_534415 : sel_534417;
  assign sel_534910 = ($signed({1'h0, add_534095}) < $signed({1'h0, sel_534097}) ? add_534095 : sel_534097) == ($signed({1'h0, add_534099}) < $signed({1'h0, sel_534101}) ? add_534099 : sel_534101) ? add_534753 : sel_534594;
  assign add_534917 = array_index_514558[11:2] + 10'h113;
  assign sel_534919 = $signed({1'h0, add_534443, array_index_514318[1:0]}) < $signed({1'h0, sel_534445}) ? {add_534443, array_index_514318[1:0]} : sel_534445;
  assign add_534921 = array_index_514561[11:2] + 10'h113;
  assign sel_534923 = $signed({1'h0, add_534447, array_index_514321[1:0]}) < $signed({1'h0, sel_534449}) ? {add_534447, array_index_514321[1:0]} : sel_534449;
  assign add_534935 = array_index_515098[11:4] + 8'h49;
  assign sel_534937 = $signed({1'h0, add_534461, array_index_514818[3:0]}) < $signed({1'h0, sel_534463}) ? {add_534461, array_index_514818[3:0]} : sel_534463;
  assign add_534939 = array_index_515101[11:4] + 8'h49;
  assign sel_534941 = $signed({1'h0, add_534465, array_index_514821[3:0]}) < $signed({1'h0, sel_534467}) ? {add_534465, array_index_514821[3:0]} : sel_534467;
  assign add_534951 = array_index_515726[11:0] + 12'h263;
  assign sel_534953 = $signed({1'h0, add_534477}) < $signed({1'h0, sel_534479}) ? add_534477 : sel_534479;
  assign add_534955 = array_index_515729[11:0] + 12'h263;
  assign sel_534957 = $signed({1'h0, add_534481}) < $signed({1'h0, sel_534483}) ? add_534481 : sel_534483;
  assign add_534967 = array_index_516458[11:1] + 11'h109;
  assign sel_534969 = $signed({1'h0, add_534493, array_index_516080[0]}) < $signed({1'h0, sel_534495}) ? {add_534493, array_index_516080[0]} : sel_534495;
  assign add_534971 = array_index_516461[11:1] + 11'h109;
  assign sel_534973 = $signed({1'h0, add_534497, array_index_516083[0]}) < $signed({1'h0, sel_534499}) ? {add_534497, array_index_516083[0]} : sel_534499;
  assign add_534983 = array_index_517286[11:3] + 9'h12f;
  assign sel_534985 = $signed({1'h0, add_534509, array_index_516860[2:0]}) < $signed({1'h0, sel_534511}) ? {add_534509, array_index_516860[2:0]} : sel_534511;
  assign add_534987 = array_index_517289[11:3] + 9'h12f;
  assign sel_534989 = $signed({1'h0, add_534513, array_index_516863[2:0]}) < $signed({1'h0, sel_534515}) ? {add_534513, array_index_516863[2:0]} : sel_534515;
  assign add_535001 = array_index_518210[11:3] + 9'h171;
  assign sel_535003 = $signed({1'h0, add_534527, array_index_517736[2:0]}) < $signed({1'h0, sel_534529}) ? {add_534527, array_index_517736[2:0]} : sel_534529;
  assign add_535005 = array_index_518213[11:3] + 9'h171;
  assign sel_535007 = $signed({1'h0, add_534531, array_index_517739[2:0]}) < $signed({1'h0, sel_534533}) ? {add_534531, array_index_517739[2:0]} : sel_534533;
  assign add_535017 = array_index_519236[11:0] + 12'h091;
  assign sel_535019 = $signed({1'h0, add_534543}) < $signed({1'h0, sel_534545}) ? add_534543 : sel_534545;
  assign add_535021 = array_index_519239[11:0] + 12'h091;
  assign sel_535023 = $signed({1'h0, add_534547}) < $signed({1'h0, sel_534549}) ? add_534547 : sel_534549;
  assign add_535033 = array_index_520362[11:0] + 12'hf59;
  assign sel_535035 = $signed({1'h0, add_534559}) < $signed({1'h0, sel_534561}) ? add_534559 : sel_534561;
  assign add_535037 = array_index_520365[11:0] + 12'hf59;
  assign sel_535039 = $signed({1'h0, add_534563}) < $signed({1'h0, sel_534565}) ? add_534563 : sel_534565;
  assign add_535051 = array_index_521590[11:0] + 12'h437;
  assign sel_535053 = $signed({1'h0, add_534577}) < $signed({1'h0, sel_534579}) ? add_534577 : sel_534579;
  assign add_535055 = array_index_521593[11:0] + 12'h437;
  assign sel_535057 = $signed({1'h0, add_534581}) < $signed({1'h0, sel_534583}) ? add_534581 : sel_534583;
  assign add_535061 = sel_534910 + 16'h0001;
  assign add_535071 = array_index_514818[11:1] + 11'h5b9;
  assign sel_535073 = $signed({1'h0, add_534605, array_index_514558[0]}) < $signed({1'h0, sel_534607}) ? {add_534605, array_index_514558[0]} : sel_534607;
  assign add_535075 = array_index_514821[11:1] + 11'h5b9;
  assign sel_535077 = $signed({1'h0, add_534609, array_index_514561[0]}) < $signed({1'h0, sel_534611}) ? {add_534609, array_index_514561[0]} : sel_534611;
  assign add_535087 = array_index_515398[11:0] + 12'h37b;
  assign sel_535089 = $signed({1'h0, add_534621}) < $signed({1'h0, sel_534623}) ? add_534621 : sel_534623;
  assign add_535091 = array_index_515401[11:0] + 12'h37b;
  assign sel_535093 = $signed({1'h0, add_534625}) < $signed({1'h0, sel_534627}) ? add_534625 : sel_534627;
  assign add_535105 = array_index_516080[11:0] + 12'h811;
  assign sel_535107 = $signed({1'h0, add_534639}) < $signed({1'h0, sel_534641}) ? add_534639 : sel_534641;
  assign add_535109 = array_index_516083[11:0] + 12'h811;
  assign sel_535111 = $signed({1'h0, add_534643}) < $signed({1'h0, sel_534645}) ? add_534643 : sel_534645;
  assign add_535123 = array_index_516860[11:0] + 12'h70f;
  assign sel_535125 = $signed({1'h0, add_534657}) < $signed({1'h0, sel_534659}) ? add_534657 : sel_534659;
  assign add_535127 = array_index_516863[11:0] + 12'h70f;
  assign sel_535129 = $signed({1'h0, add_534661}) < $signed({1'h0, sel_534663}) ? add_534661 : sel_534663;
  assign add_535141 = array_index_517736[11:3] + 9'h1f1;
  assign sel_535143 = $signed({1'h0, add_534675, array_index_517286[2:0]}) < $signed({1'h0, sel_534677}) ? {add_534675, array_index_517286[2:0]} : sel_534677;
  assign add_535145 = array_index_517739[11:3] + 9'h1f1;
  assign sel_535147 = $signed({1'h0, add_534679, array_index_517289[2:0]}) < $signed({1'h0, sel_534681}) ? {add_534679, array_index_517289[2:0]} : sel_534681;
  assign add_535157 = array_index_518710[11:0] + 12'h081;
  assign sel_535159 = $signed({1'h0, add_534691}) < $signed({1'h0, sel_534693}) ? add_534691 : sel_534693;
  assign add_535161 = array_index_518713[11:0] + 12'h081;
  assign sel_535163 = $signed({1'h0, add_534695}) < $signed({1'h0, sel_534697}) ? add_534695 : sel_534697;
  assign add_535175 = array_index_519786[11:0] + 12'h0b1;
  assign sel_535177 = $signed({1'h0, add_534709}) < $signed({1'h0, sel_534711}) ? add_534709 : sel_534711;
  assign add_535179 = array_index_519789[11:0] + 12'h0b1;
  assign sel_535181 = $signed({1'h0, add_534713}) < $signed({1'h0, sel_534715}) ? add_534713 : sel_534715;
  assign add_535193 = array_index_520964[11:1] + 11'h4c1;
  assign sel_535195 = $signed({1'h0, add_534727, array_index_520362[0]}) < $signed({1'h0, sel_534729}) ? {add_534727, array_index_520362[0]} : sel_534729;
  assign add_535197 = array_index_520967[11:1] + 11'h4c1;
  assign sel_535199 = $signed({1'h0, add_534731, array_index_520365[0]}) < $signed({1'h0, sel_534733}) ? {add_534731, array_index_520365[0]} : sel_534733;
  assign sel_535210 = ($signed({1'h0, add_534427}) < $signed({1'h0, sel_534429}) ? add_534427 : sel_534429) == ($signed({1'h0, add_534431}) < $signed({1'h0, sel_534433}) ? add_534431 : sel_534433) ? add_535061 : sel_534910;
  assign add_535213 = array_index_514558[11:0] + 12'hcc1;
  assign sel_535215 = $signed({1'h0, add_534755}) < $signed({1'h0, sel_534757}) ? add_534755 : sel_534757;
  assign add_535217 = array_index_514561[11:0] + 12'hcc1;
  assign sel_535219 = $signed({1'h0, add_534759}) < $signed({1'h0, sel_534761}) ? add_534759 : sel_534761;
  assign add_535231 = array_index_515098[11:0] + 12'ha87;
  assign sel_535233 = $signed({1'h0, add_534773}) < $signed({1'h0, sel_534775}) ? add_534773 : sel_534775;
  assign add_535235 = array_index_515101[11:0] + 12'ha87;
  assign sel_535237 = $signed({1'h0, add_534777}) < $signed({1'h0, sel_534779}) ? add_534777 : sel_534779;
  assign add_535249 = array_index_515726[11:1] + 11'h663;
  assign sel_535251 = $signed({1'h0, add_534791, array_index_515398[0]}) < $signed({1'h0, sel_534793}) ? {add_534791, array_index_515398[0]} : sel_534793;
  assign add_535253 = array_index_515729[11:1] + 11'h663;
  assign sel_535255 = $signed({1'h0, add_534795, array_index_515401[0]}) < $signed({1'h0, sel_534797}) ? {add_534795, array_index_515401[0]} : sel_534797;
  assign add_535265 = array_index_516458[11:1] + 11'h075;
  assign sel_535267 = $signed({1'h0, add_534807, array_index_516080[0]}) < $signed({1'h0, sel_534809}) ? {add_534807, array_index_516080[0]} : sel_534809;
  assign add_535269 = array_index_516461[11:1] + 11'h075;
  assign sel_535271 = $signed({1'h0, add_534811, array_index_516083[0]}) < $signed({1'h0, sel_534813}) ? {add_534811, array_index_516083[0]} : sel_534813;
  assign add_535283 = array_index_517286[11:2] + 10'h181;
  assign sel_535285 = $signed({1'h0, add_534825, array_index_516860[1:0]}) < $signed({1'h0, sel_534827}) ? {add_534825, array_index_516860[1:0]} : sel_534827;
  assign add_535287 = array_index_517289[11:2] + 10'h181;
  assign sel_535289 = $signed({1'h0, add_534829, array_index_516863[1:0]}) < $signed({1'h0, sel_534831}) ? {add_534829, array_index_516863[1:0]} : sel_534831;
  assign add_535301 = array_index_518210[11:0] + 12'h8a7;
  assign sel_535303 = $signed({1'h0, add_534843}) < $signed({1'h0, sel_534845}) ? add_534843 : sel_534845;
  assign add_535305 = array_index_518213[11:0] + 12'h8a7;
  assign sel_535307 = $signed({1'h0, add_534847}) < $signed({1'h0, sel_534849}) ? add_534847 : sel_534849;
  assign add_535319 = array_index_519236[11:1] + 11'h283;
  assign sel_535321 = $signed({1'h0, add_534861, array_index_518710[0]}) < $signed({1'h0, sel_534863}) ? {add_534861, array_index_518710[0]} : sel_534863;
  assign add_535323 = array_index_519239[11:1] + 11'h283;
  assign sel_535325 = $signed({1'h0, add_534865, array_index_518713[0]}) < $signed({1'h0, sel_534867}) ? {add_534865, array_index_518713[0]} : sel_534867;
  assign add_535335 = array_index_520362[11:1] + 11'h44d;
  assign sel_535337 = $signed({1'h0, add_534877, array_index_519786[0]}) < $signed({1'h0, sel_534879}) ? {add_534877, array_index_519786[0]} : sel_534879;
  assign add_535339 = array_index_520365[11:1] + 11'h44d;
  assign sel_535341 = $signed({1'h0, add_534881, array_index_519789[0]}) < $signed({1'h0, sel_534883}) ? {add_534881, array_index_519789[0]} : sel_534883;
  assign add_535351 = array_index_521590[11:0] + 12'hcb1;
  assign sel_535353 = $signed({1'h0, add_534893}) < $signed({1'h0, sel_534895}) ? add_534893 : sel_534895;
  assign add_535355 = array_index_521593[11:0] + 12'hcb1;
  assign sel_535357 = $signed({1'h0, add_534897}) < $signed({1'h0, sel_534899}) ? add_534897 : sel_534899;
  assign add_535361 = sel_535210 + 16'h0001;
  assign add_535367 = array_index_514818[11:2] + 10'h113;
  assign sel_535369 = $signed({1'h0, add_534917, array_index_514558[1:0]}) < $signed({1'h0, sel_534919}) ? {add_534917, array_index_514558[1:0]} : sel_534919;
  assign add_535371 = array_index_514821[11:2] + 10'h113;
  assign sel_535373 = $signed({1'h0, add_534921, array_index_514561[1:0]}) < $signed({1'h0, sel_534923}) ? {add_534921, array_index_514561[1:0]} : sel_534923;
  assign add_535385 = array_index_515398[11:4] + 8'h49;
  assign sel_535387 = $signed({1'h0, add_534935, array_index_515098[3:0]}) < $signed({1'h0, sel_534937}) ? {add_534935, array_index_515098[3:0]} : sel_534937;
  assign add_535389 = array_index_515401[11:4] + 8'h49;
  assign sel_535391 = $signed({1'h0, add_534939, array_index_515101[3:0]}) < $signed({1'h0, sel_534941}) ? {add_534939, array_index_515101[3:0]} : sel_534941;
  assign add_535401 = array_index_516080[11:0] + 12'h263;
  assign sel_535403 = $signed({1'h0, add_534951}) < $signed({1'h0, sel_534953}) ? add_534951 : sel_534953;
  assign add_535405 = array_index_516083[11:0] + 12'h263;
  assign sel_535407 = $signed({1'h0, add_534955}) < $signed({1'h0, sel_534957}) ? add_534955 : sel_534957;
  assign add_535417 = array_index_516860[11:1] + 11'h109;
  assign sel_535419 = $signed({1'h0, add_534967, array_index_516458[0]}) < $signed({1'h0, sel_534969}) ? {add_534967, array_index_516458[0]} : sel_534969;
  assign add_535421 = array_index_516863[11:1] + 11'h109;
  assign sel_535423 = $signed({1'h0, add_534971, array_index_516461[0]}) < $signed({1'h0, sel_534973}) ? {add_534971, array_index_516461[0]} : sel_534973;
  assign add_535433 = array_index_517736[11:3] + 9'h12f;
  assign sel_535435 = $signed({1'h0, add_534983, array_index_517286[2:0]}) < $signed({1'h0, sel_534985}) ? {add_534983, array_index_517286[2:0]} : sel_534985;
  assign add_535437 = array_index_517739[11:3] + 9'h12f;
  assign sel_535439 = $signed({1'h0, add_534987, array_index_517289[2:0]}) < $signed({1'h0, sel_534989}) ? {add_534987, array_index_517289[2:0]} : sel_534989;
  assign add_535451 = array_index_518710[11:3] + 9'h171;
  assign sel_535453 = $signed({1'h0, add_535001, array_index_518210[2:0]}) < $signed({1'h0, sel_535003}) ? {add_535001, array_index_518210[2:0]} : sel_535003;
  assign add_535455 = array_index_518713[11:3] + 9'h171;
  assign sel_535457 = $signed({1'h0, add_535005, array_index_518213[2:0]}) < $signed({1'h0, sel_535007}) ? {add_535005, array_index_518213[2:0]} : sel_535007;
  assign add_535467 = array_index_519786[11:0] + 12'h091;
  assign sel_535469 = $signed({1'h0, add_535017}) < $signed({1'h0, sel_535019}) ? add_535017 : sel_535019;
  assign add_535471 = array_index_519789[11:0] + 12'h091;
  assign sel_535473 = $signed({1'h0, add_535021}) < $signed({1'h0, sel_535023}) ? add_535021 : sel_535023;
  assign add_535483 = array_index_520964[11:0] + 12'hf59;
  assign sel_535485 = $signed({1'h0, add_535033}) < $signed({1'h0, sel_535035}) ? add_535033 : sel_535035;
  assign add_535487 = array_index_520967[11:0] + 12'hf59;
  assign sel_535489 = $signed({1'h0, add_535037}) < $signed({1'h0, sel_535039}) ? add_535037 : sel_535039;
  assign sel_535502 = ($signed({1'h0, add_534743}) < $signed({1'h0, sel_534745}) ? add_534743 : sel_534745) == ($signed({1'h0, add_534747}) < $signed({1'h0, sel_534749}) ? add_534747 : sel_534749) ? add_535361 : sel_535210;
  assign add_535513 = array_index_515098[11:1] + 11'h5b9;
  assign sel_535515 = $signed({1'h0, add_535071, array_index_514818[0]}) < $signed({1'h0, sel_535073}) ? {add_535071, array_index_514818[0]} : sel_535073;
  assign add_535517 = array_index_515101[11:1] + 11'h5b9;
  assign sel_535519 = $signed({1'h0, add_535075, array_index_514821[0]}) < $signed({1'h0, sel_535077}) ? {add_535075, array_index_514821[0]} : sel_535077;
  assign add_535529 = array_index_515726[11:0] + 12'h37b;
  assign sel_535531 = $signed({1'h0, add_535087}) < $signed({1'h0, sel_535089}) ? add_535087 : sel_535089;
  assign add_535533 = array_index_515729[11:0] + 12'h37b;
  assign sel_535535 = $signed({1'h0, add_535091}) < $signed({1'h0, sel_535093}) ? add_535091 : sel_535093;
  assign add_535547 = array_index_516458[11:0] + 12'h811;
  assign sel_535549 = $signed({1'h0, add_535105}) < $signed({1'h0, sel_535107}) ? add_535105 : sel_535107;
  assign add_535551 = array_index_516461[11:0] + 12'h811;
  assign sel_535553 = $signed({1'h0, add_535109}) < $signed({1'h0, sel_535111}) ? add_535109 : sel_535111;
  assign add_535565 = array_index_517286[11:0] + 12'h70f;
  assign sel_535567 = $signed({1'h0, add_535123}) < $signed({1'h0, sel_535125}) ? add_535123 : sel_535125;
  assign add_535569 = array_index_517289[11:0] + 12'h70f;
  assign sel_535571 = $signed({1'h0, add_535127}) < $signed({1'h0, sel_535129}) ? add_535127 : sel_535129;
  assign add_535583 = array_index_518210[11:3] + 9'h1f1;
  assign sel_535585 = $signed({1'h0, add_535141, array_index_517736[2:0]}) < $signed({1'h0, sel_535143}) ? {add_535141, array_index_517736[2:0]} : sel_535143;
  assign add_535587 = array_index_518213[11:3] + 9'h1f1;
  assign sel_535589 = $signed({1'h0, add_535145, array_index_517739[2:0]}) < $signed({1'h0, sel_535147}) ? {add_535145, array_index_517739[2:0]} : sel_535147;
  assign add_535599 = array_index_519236[11:0] + 12'h081;
  assign sel_535601 = $signed({1'h0, add_535157}) < $signed({1'h0, sel_535159}) ? add_535157 : sel_535159;
  assign add_535603 = array_index_519239[11:0] + 12'h081;
  assign sel_535605 = $signed({1'h0, add_535161}) < $signed({1'h0, sel_535163}) ? add_535161 : sel_535163;
  assign add_535617 = array_index_520362[11:0] + 12'h0b1;
  assign sel_535619 = $signed({1'h0, add_535175}) < $signed({1'h0, sel_535177}) ? add_535175 : sel_535177;
  assign add_535621 = array_index_520365[11:0] + 12'h0b1;
  assign sel_535623 = $signed({1'h0, add_535179}) < $signed({1'h0, sel_535181}) ? add_535179 : sel_535181;
  assign add_535635 = array_index_521590[11:1] + 11'h4c1;
  assign sel_535637 = $signed({1'h0, add_535193, array_index_520964[0]}) < $signed({1'h0, sel_535195}) ? {add_535193, array_index_520964[0]} : sel_535195;
  assign add_535639 = array_index_521593[11:1] + 11'h4c1;
  assign sel_535641 = $signed({1'h0, add_535197, array_index_520967[0]}) < $signed({1'h0, sel_535199}) ? {add_535197, array_index_520967[0]} : sel_535199;
  assign add_535645 = sel_535502 + 16'h0001;
  assign add_535647 = array_index_514818[11:0] + 12'hcc1;
  assign sel_535649 = $signed({1'h0, add_535213}) < $signed({1'h0, sel_535215}) ? add_535213 : sel_535215;
  assign add_535651 = array_index_514821[11:0] + 12'hcc1;
  assign sel_535653 = $signed({1'h0, add_535217}) < $signed({1'h0, sel_535219}) ? add_535217 : sel_535219;
  assign add_535665 = array_index_515398[11:0] + 12'ha87;
  assign sel_535667 = $signed({1'h0, add_535231}) < $signed({1'h0, sel_535233}) ? add_535231 : sel_535233;
  assign add_535669 = array_index_515401[11:0] + 12'ha87;
  assign sel_535671 = $signed({1'h0, add_535235}) < $signed({1'h0, sel_535237}) ? add_535235 : sel_535237;
  assign add_535683 = array_index_516080[11:1] + 11'h663;
  assign sel_535685 = $signed({1'h0, add_535249, array_index_515726[0]}) < $signed({1'h0, sel_535251}) ? {add_535249, array_index_515726[0]} : sel_535251;
  assign add_535687 = array_index_516083[11:1] + 11'h663;
  assign sel_535689 = $signed({1'h0, add_535253, array_index_515729[0]}) < $signed({1'h0, sel_535255}) ? {add_535253, array_index_515729[0]} : sel_535255;
  assign add_535699 = array_index_516860[11:1] + 11'h075;
  assign sel_535701 = $signed({1'h0, add_535265, array_index_516458[0]}) < $signed({1'h0, sel_535267}) ? {add_535265, array_index_516458[0]} : sel_535267;
  assign add_535703 = array_index_516863[11:1] + 11'h075;
  assign sel_535705 = $signed({1'h0, add_535269, array_index_516461[0]}) < $signed({1'h0, sel_535271}) ? {add_535269, array_index_516461[0]} : sel_535271;
  assign add_535717 = array_index_517736[11:2] + 10'h181;
  assign sel_535719 = $signed({1'h0, add_535283, array_index_517286[1:0]}) < $signed({1'h0, sel_535285}) ? {add_535283, array_index_517286[1:0]} : sel_535285;
  assign add_535721 = array_index_517739[11:2] + 10'h181;
  assign sel_535723 = $signed({1'h0, add_535287, array_index_517289[1:0]}) < $signed({1'h0, sel_535289}) ? {add_535287, array_index_517289[1:0]} : sel_535289;
  assign add_535735 = array_index_518710[11:0] + 12'h8a7;
  assign sel_535737 = $signed({1'h0, add_535301}) < $signed({1'h0, sel_535303}) ? add_535301 : sel_535303;
  assign add_535739 = array_index_518713[11:0] + 12'h8a7;
  assign sel_535741 = $signed({1'h0, add_535305}) < $signed({1'h0, sel_535307}) ? add_535305 : sel_535307;
  assign add_535753 = array_index_519786[11:1] + 11'h283;
  assign sel_535755 = $signed({1'h0, add_535319, array_index_519236[0]}) < $signed({1'h0, sel_535321}) ? {add_535319, array_index_519236[0]} : sel_535321;
  assign add_535757 = array_index_519789[11:1] + 11'h283;
  assign sel_535759 = $signed({1'h0, add_535323, array_index_519239[0]}) < $signed({1'h0, sel_535325}) ? {add_535323, array_index_519239[0]} : sel_535325;
  assign add_535769 = array_index_520964[11:1] + 11'h44d;
  assign sel_535771 = $signed({1'h0, add_535335, array_index_520362[0]}) < $signed({1'h0, sel_535337}) ? {add_535335, array_index_520362[0]} : sel_535337;
  assign add_535773 = array_index_520967[11:1] + 11'h44d;
  assign sel_535775 = $signed({1'h0, add_535339, array_index_520365[0]}) < $signed({1'h0, sel_535341}) ? {add_535339, array_index_520365[0]} : sel_535341;
  assign sel_535786 = ($signed({1'h0, add_535051}) < $signed({1'h0, sel_535053}) ? add_535051 : sel_535053) == ($signed({1'h0, add_535055}) < $signed({1'h0, sel_535057}) ? add_535055 : sel_535057) ? add_535645 : sel_535502;
  assign add_535793 = array_index_515098[11:2] + 10'h113;
  assign sel_535795 = $signed({1'h0, add_535367, array_index_514818[1:0]}) < $signed({1'h0, sel_535369}) ? {add_535367, array_index_514818[1:0]} : sel_535369;
  assign add_535797 = array_index_515101[11:2] + 10'h113;
  assign sel_535799 = $signed({1'h0, add_535371, array_index_514821[1:0]}) < $signed({1'h0, sel_535373}) ? {add_535371, array_index_514821[1:0]} : sel_535373;
  assign add_535811 = array_index_515726[11:4] + 8'h49;
  assign sel_535813 = $signed({1'h0, add_535385, array_index_515398[3:0]}) < $signed({1'h0, sel_535387}) ? {add_535385, array_index_515398[3:0]} : sel_535387;
  assign add_535815 = array_index_515729[11:4] + 8'h49;
  assign sel_535817 = $signed({1'h0, add_535389, array_index_515401[3:0]}) < $signed({1'h0, sel_535391}) ? {add_535389, array_index_515401[3:0]} : sel_535391;
  assign add_535827 = array_index_516458[11:0] + 12'h263;
  assign sel_535829 = $signed({1'h0, add_535401}) < $signed({1'h0, sel_535403}) ? add_535401 : sel_535403;
  assign add_535831 = array_index_516461[11:0] + 12'h263;
  assign sel_535833 = $signed({1'h0, add_535405}) < $signed({1'h0, sel_535407}) ? add_535405 : sel_535407;
  assign add_535843 = array_index_517286[11:1] + 11'h109;
  assign sel_535845 = $signed({1'h0, add_535417, array_index_516860[0]}) < $signed({1'h0, sel_535419}) ? {add_535417, array_index_516860[0]} : sel_535419;
  assign add_535847 = array_index_517289[11:1] + 11'h109;
  assign sel_535849 = $signed({1'h0, add_535421, array_index_516863[0]}) < $signed({1'h0, sel_535423}) ? {add_535421, array_index_516863[0]} : sel_535423;
  assign add_535859 = array_index_518210[11:3] + 9'h12f;
  assign sel_535861 = $signed({1'h0, add_535433, array_index_517736[2:0]}) < $signed({1'h0, sel_535435}) ? {add_535433, array_index_517736[2:0]} : sel_535435;
  assign add_535863 = array_index_518213[11:3] + 9'h12f;
  assign sel_535865 = $signed({1'h0, add_535437, array_index_517739[2:0]}) < $signed({1'h0, sel_535439}) ? {add_535437, array_index_517739[2:0]} : sel_535439;
  assign add_535877 = array_index_519236[11:3] + 9'h171;
  assign sel_535879 = $signed({1'h0, add_535451, array_index_518710[2:0]}) < $signed({1'h0, sel_535453}) ? {add_535451, array_index_518710[2:0]} : sel_535453;
  assign add_535881 = array_index_519239[11:3] + 9'h171;
  assign sel_535883 = $signed({1'h0, add_535455, array_index_518713[2:0]}) < $signed({1'h0, sel_535457}) ? {add_535455, array_index_518713[2:0]} : sel_535457;
  assign add_535893 = array_index_520362[11:0] + 12'h091;
  assign sel_535895 = $signed({1'h0, add_535467}) < $signed({1'h0, sel_535469}) ? add_535467 : sel_535469;
  assign add_535897 = array_index_520365[11:0] + 12'h091;
  assign sel_535899 = $signed({1'h0, add_535471}) < $signed({1'h0, sel_535473}) ? add_535471 : sel_535473;
  assign add_535909 = array_index_521590[11:0] + 12'hf59;
  assign sel_535911 = $signed({1'h0, add_535483}) < $signed({1'h0, sel_535485}) ? add_535483 : sel_535485;
  assign add_535913 = array_index_521593[11:0] + 12'hf59;
  assign sel_535915 = $signed({1'h0, add_535487}) < $signed({1'h0, sel_535489}) ? add_535487 : sel_535489;
  assign add_535921 = sel_535786 + 16'h0001;
  assign add_535931 = array_index_515398[11:1] + 11'h5b9;
  assign sel_535933 = $signed({1'h0, add_535513, array_index_515098[0]}) < $signed({1'h0, sel_535515}) ? {add_535513, array_index_515098[0]} : sel_535515;
  assign add_535935 = array_index_515401[11:1] + 11'h5b9;
  assign sel_535937 = $signed({1'h0, add_535517, array_index_515101[0]}) < $signed({1'h0, sel_535519}) ? {add_535517, array_index_515101[0]} : sel_535519;
  assign add_535947 = array_index_516080[11:0] + 12'h37b;
  assign sel_535949 = $signed({1'h0, add_535529}) < $signed({1'h0, sel_535531}) ? add_535529 : sel_535531;
  assign add_535951 = array_index_516083[11:0] + 12'h37b;
  assign sel_535953 = $signed({1'h0, add_535533}) < $signed({1'h0, sel_535535}) ? add_535533 : sel_535535;
  assign add_535965 = array_index_516860[11:0] + 12'h811;
  assign sel_535967 = $signed({1'h0, add_535547}) < $signed({1'h0, sel_535549}) ? add_535547 : sel_535549;
  assign add_535969 = array_index_516863[11:0] + 12'h811;
  assign sel_535971 = $signed({1'h0, add_535551}) < $signed({1'h0, sel_535553}) ? add_535551 : sel_535553;
  assign add_535983 = array_index_517736[11:0] + 12'h70f;
  assign sel_535985 = $signed({1'h0, add_535565}) < $signed({1'h0, sel_535567}) ? add_535565 : sel_535567;
  assign add_535987 = array_index_517739[11:0] + 12'h70f;
  assign sel_535989 = $signed({1'h0, add_535569}) < $signed({1'h0, sel_535571}) ? add_535569 : sel_535571;
  assign add_536001 = array_index_518710[11:3] + 9'h1f1;
  assign sel_536003 = $signed({1'h0, add_535583, array_index_518210[2:0]}) < $signed({1'h0, sel_535585}) ? {add_535583, array_index_518210[2:0]} : sel_535585;
  assign add_536005 = array_index_518713[11:3] + 9'h1f1;
  assign sel_536007 = $signed({1'h0, add_535587, array_index_518213[2:0]}) < $signed({1'h0, sel_535589}) ? {add_535587, array_index_518213[2:0]} : sel_535589;
  assign add_536017 = array_index_519786[11:0] + 12'h081;
  assign sel_536019 = $signed({1'h0, add_535599}) < $signed({1'h0, sel_535601}) ? add_535599 : sel_535601;
  assign add_536021 = array_index_519789[11:0] + 12'h081;
  assign sel_536023 = $signed({1'h0, add_535603}) < $signed({1'h0, sel_535605}) ? add_535603 : sel_535605;
  assign add_536035 = array_index_520964[11:0] + 12'h0b1;
  assign sel_536037 = $signed({1'h0, add_535617}) < $signed({1'h0, sel_535619}) ? add_535617 : sel_535619;
  assign add_536039 = array_index_520967[11:0] + 12'h0b1;
  assign sel_536041 = $signed({1'h0, add_535621}) < $signed({1'h0, sel_535623}) ? add_535621 : sel_535623;
  assign sel_536054 = ($signed({1'h0, add_535351}) < $signed({1'h0, sel_535353}) ? add_535351 : sel_535353) == ($signed({1'h0, add_535355}) < $signed({1'h0, sel_535357}) ? add_535355 : sel_535357) ? add_535921 : sel_535786;
  assign add_536057 = array_index_515098[11:0] + 12'hcc1;
  assign sel_536059 = $signed({1'h0, add_535647}) < $signed({1'h0, sel_535649}) ? add_535647 : sel_535649;
  assign add_536061 = array_index_515101[11:0] + 12'hcc1;
  assign sel_536063 = $signed({1'h0, add_535651}) < $signed({1'h0, sel_535653}) ? add_535651 : sel_535653;
  assign add_536075 = array_index_515726[11:0] + 12'ha87;
  assign sel_536077 = $signed({1'h0, add_535665}) < $signed({1'h0, sel_535667}) ? add_535665 : sel_535667;
  assign add_536079 = array_index_515729[11:0] + 12'ha87;
  assign sel_536081 = $signed({1'h0, add_535669}) < $signed({1'h0, sel_535671}) ? add_535669 : sel_535671;
  assign add_536093 = array_index_516458[11:1] + 11'h663;
  assign sel_536095 = $signed({1'h0, add_535683, array_index_516080[0]}) < $signed({1'h0, sel_535685}) ? {add_535683, array_index_516080[0]} : sel_535685;
  assign add_536097 = array_index_516461[11:1] + 11'h663;
  assign sel_536099 = $signed({1'h0, add_535687, array_index_516083[0]}) < $signed({1'h0, sel_535689}) ? {add_535687, array_index_516083[0]} : sel_535689;
  assign add_536109 = array_index_517286[11:1] + 11'h075;
  assign sel_536111 = $signed({1'h0, add_535699, array_index_516860[0]}) < $signed({1'h0, sel_535701}) ? {add_535699, array_index_516860[0]} : sel_535701;
  assign add_536113 = array_index_517289[11:1] + 11'h075;
  assign sel_536115 = $signed({1'h0, add_535703, array_index_516863[0]}) < $signed({1'h0, sel_535705}) ? {add_535703, array_index_516863[0]} : sel_535705;
  assign add_536127 = array_index_518210[11:2] + 10'h181;
  assign sel_536129 = $signed({1'h0, add_535717, array_index_517736[1:0]}) < $signed({1'h0, sel_535719}) ? {add_535717, array_index_517736[1:0]} : sel_535719;
  assign add_536131 = array_index_518213[11:2] + 10'h181;
  assign sel_536133 = $signed({1'h0, add_535721, array_index_517739[1:0]}) < $signed({1'h0, sel_535723}) ? {add_535721, array_index_517739[1:0]} : sel_535723;
  assign add_536145 = array_index_519236[11:0] + 12'h8a7;
  assign sel_536147 = $signed({1'h0, add_535735}) < $signed({1'h0, sel_535737}) ? add_535735 : sel_535737;
  assign add_536149 = array_index_519239[11:0] + 12'h8a7;
  assign sel_536151 = $signed({1'h0, add_535739}) < $signed({1'h0, sel_535741}) ? add_535739 : sel_535741;
  assign add_536163 = array_index_520362[11:1] + 11'h283;
  assign sel_536165 = $signed({1'h0, add_535753, array_index_519786[0]}) < $signed({1'h0, sel_535755}) ? {add_535753, array_index_519786[0]} : sel_535755;
  assign add_536167 = array_index_520365[11:1] + 11'h283;
  assign sel_536169 = $signed({1'h0, add_535757, array_index_519789[0]}) < $signed({1'h0, sel_535759}) ? {add_535757, array_index_519789[0]} : sel_535759;
  assign add_536179 = array_index_521590[11:1] + 11'h44d;
  assign sel_536181 = $signed({1'h0, add_535769, array_index_520964[0]}) < $signed({1'h0, sel_535771}) ? {add_535769, array_index_520964[0]} : sel_535771;
  assign add_536183 = array_index_521593[11:1] + 11'h44d;
  assign sel_536185 = $signed({1'h0, add_535773, array_index_520967[0]}) < $signed({1'h0, sel_535775}) ? {add_535773, array_index_520967[0]} : sel_535775;
  assign add_536189 = sel_536054 + 16'h0001;
  assign add_536195 = array_index_515398[11:2] + 10'h113;
  assign sel_536197 = $signed({1'h0, add_535793, array_index_515098[1:0]}) < $signed({1'h0, sel_535795}) ? {add_535793, array_index_515098[1:0]} : sel_535795;
  assign add_536199 = array_index_515401[11:2] + 10'h113;
  assign sel_536201 = $signed({1'h0, add_535797, array_index_515101[1:0]}) < $signed({1'h0, sel_535799}) ? {add_535797, array_index_515101[1:0]} : sel_535799;
  assign add_536213 = array_index_516080[11:4] + 8'h49;
  assign sel_536215 = $signed({1'h0, add_535811, array_index_515726[3:0]}) < $signed({1'h0, sel_535813}) ? {add_535811, array_index_515726[3:0]} : sel_535813;
  assign add_536217 = array_index_516083[11:4] + 8'h49;
  assign sel_536219 = $signed({1'h0, add_535815, array_index_515729[3:0]}) < $signed({1'h0, sel_535817}) ? {add_535815, array_index_515729[3:0]} : sel_535817;
  assign add_536229 = array_index_516860[11:0] + 12'h263;
  assign sel_536231 = $signed({1'h0, add_535827}) < $signed({1'h0, sel_535829}) ? add_535827 : sel_535829;
  assign add_536233 = array_index_516863[11:0] + 12'h263;
  assign sel_536235 = $signed({1'h0, add_535831}) < $signed({1'h0, sel_535833}) ? add_535831 : sel_535833;
  assign add_536245 = array_index_517736[11:1] + 11'h109;
  assign sel_536247 = $signed({1'h0, add_535843, array_index_517286[0]}) < $signed({1'h0, sel_535845}) ? {add_535843, array_index_517286[0]} : sel_535845;
  assign add_536249 = array_index_517739[11:1] + 11'h109;
  assign sel_536251 = $signed({1'h0, add_535847, array_index_517289[0]}) < $signed({1'h0, sel_535849}) ? {add_535847, array_index_517289[0]} : sel_535849;
  assign add_536261 = array_index_518710[11:3] + 9'h12f;
  assign sel_536263 = $signed({1'h0, add_535859, array_index_518210[2:0]}) < $signed({1'h0, sel_535861}) ? {add_535859, array_index_518210[2:0]} : sel_535861;
  assign add_536265 = array_index_518713[11:3] + 9'h12f;
  assign sel_536267 = $signed({1'h0, add_535863, array_index_518213[2:0]}) < $signed({1'h0, sel_535865}) ? {add_535863, array_index_518213[2:0]} : sel_535865;
  assign add_536279 = array_index_519786[11:3] + 9'h171;
  assign sel_536281 = $signed({1'h0, add_535877, array_index_519236[2:0]}) < $signed({1'h0, sel_535879}) ? {add_535877, array_index_519236[2:0]} : sel_535879;
  assign add_536283 = array_index_519789[11:3] + 9'h171;
  assign sel_536285 = $signed({1'h0, add_535881, array_index_519239[2:0]}) < $signed({1'h0, sel_535883}) ? {add_535881, array_index_519239[2:0]} : sel_535883;
  assign add_536295 = array_index_520964[11:0] + 12'h091;
  assign sel_536297 = $signed({1'h0, add_535893}) < $signed({1'h0, sel_535895}) ? add_535893 : sel_535895;
  assign add_536299 = array_index_520967[11:0] + 12'h091;
  assign sel_536301 = $signed({1'h0, add_535897}) < $signed({1'h0, sel_535899}) ? add_535897 : sel_535899;
  assign sel_536312 = ($signed({1'h0, add_535635, array_index_521590[0]}) < $signed({1'h0, sel_535637}) ? {add_535635, array_index_521590[0]} : sel_535637) == ($signed({1'h0, add_535639, array_index_521593[0]}) < $signed({1'h0, sel_535641}) ? {add_535639, array_index_521593[0]} : sel_535641) ? add_536189 : sel_536054;
  assign add_536323 = array_index_515726[11:1] + 11'h5b9;
  assign sel_536325 = $signed({1'h0, add_535931, array_index_515398[0]}) < $signed({1'h0, sel_535933}) ? {add_535931, array_index_515398[0]} : sel_535933;
  assign add_536327 = array_index_515729[11:1] + 11'h5b9;
  assign sel_536329 = $signed({1'h0, add_535935, array_index_515401[0]}) < $signed({1'h0, sel_535937}) ? {add_535935, array_index_515401[0]} : sel_535937;
  assign add_536339 = array_index_516458[11:0] + 12'h37b;
  assign sel_536341 = $signed({1'h0, add_535947}) < $signed({1'h0, sel_535949}) ? add_535947 : sel_535949;
  assign add_536343 = array_index_516461[11:0] + 12'h37b;
  assign sel_536345 = $signed({1'h0, add_535951}) < $signed({1'h0, sel_535953}) ? add_535951 : sel_535953;
  assign add_536357 = array_index_517286[11:0] + 12'h811;
  assign sel_536359 = $signed({1'h0, add_535965}) < $signed({1'h0, sel_535967}) ? add_535965 : sel_535967;
  assign add_536361 = array_index_517289[11:0] + 12'h811;
  assign sel_536363 = $signed({1'h0, add_535969}) < $signed({1'h0, sel_535971}) ? add_535969 : sel_535971;
  assign add_536375 = array_index_518210[11:0] + 12'h70f;
  assign sel_536377 = $signed({1'h0, add_535983}) < $signed({1'h0, sel_535985}) ? add_535983 : sel_535985;
  assign add_536379 = array_index_518213[11:0] + 12'h70f;
  assign sel_536381 = $signed({1'h0, add_535987}) < $signed({1'h0, sel_535989}) ? add_535987 : sel_535989;
  assign add_536393 = array_index_519236[11:3] + 9'h1f1;
  assign sel_536395 = $signed({1'h0, add_536001, array_index_518710[2:0]}) < $signed({1'h0, sel_536003}) ? {add_536001, array_index_518710[2:0]} : sel_536003;
  assign add_536397 = array_index_519239[11:3] + 9'h1f1;
  assign sel_536399 = $signed({1'h0, add_536005, array_index_518713[2:0]}) < $signed({1'h0, sel_536007}) ? {add_536005, array_index_518713[2:0]} : sel_536007;
  assign add_536409 = array_index_520362[11:0] + 12'h081;
  assign sel_536411 = $signed({1'h0, add_536017}) < $signed({1'h0, sel_536019}) ? add_536017 : sel_536019;
  assign add_536413 = array_index_520365[11:0] + 12'h081;
  assign sel_536415 = $signed({1'h0, add_536021}) < $signed({1'h0, sel_536023}) ? add_536021 : sel_536023;
  assign add_536427 = array_index_521590[11:0] + 12'h0b1;
  assign sel_536429 = $signed({1'h0, add_536035}) < $signed({1'h0, sel_536037}) ? add_536035 : sel_536037;
  assign add_536431 = array_index_521593[11:0] + 12'h0b1;
  assign sel_536433 = $signed({1'h0, add_536039}) < $signed({1'h0, sel_536041}) ? add_536039 : sel_536041;
  assign add_536439 = sel_536312 + 16'h0001;
  assign add_536441 = array_index_515398[11:0] + 12'hcc1;
  assign sel_536443 = $signed({1'h0, add_536057}) < $signed({1'h0, sel_536059}) ? add_536057 : sel_536059;
  assign add_536445 = array_index_515401[11:0] + 12'hcc1;
  assign sel_536447 = $signed({1'h0, add_536061}) < $signed({1'h0, sel_536063}) ? add_536061 : sel_536063;
  assign add_536459 = array_index_516080[11:0] + 12'ha87;
  assign sel_536461 = $signed({1'h0, add_536075}) < $signed({1'h0, sel_536077}) ? add_536075 : sel_536077;
  assign add_536463 = array_index_516083[11:0] + 12'ha87;
  assign sel_536465 = $signed({1'h0, add_536079}) < $signed({1'h0, sel_536081}) ? add_536079 : sel_536081;
  assign add_536477 = array_index_516860[11:1] + 11'h663;
  assign sel_536479 = $signed({1'h0, add_536093, array_index_516458[0]}) < $signed({1'h0, sel_536095}) ? {add_536093, array_index_516458[0]} : sel_536095;
  assign add_536481 = array_index_516863[11:1] + 11'h663;
  assign sel_536483 = $signed({1'h0, add_536097, array_index_516461[0]}) < $signed({1'h0, sel_536099}) ? {add_536097, array_index_516461[0]} : sel_536099;
  assign add_536493 = array_index_517736[11:1] + 11'h075;
  assign sel_536495 = $signed({1'h0, add_536109, array_index_517286[0]}) < $signed({1'h0, sel_536111}) ? {add_536109, array_index_517286[0]} : sel_536111;
  assign add_536497 = array_index_517739[11:1] + 11'h075;
  assign sel_536499 = $signed({1'h0, add_536113, array_index_517289[0]}) < $signed({1'h0, sel_536115}) ? {add_536113, array_index_517289[0]} : sel_536115;
  assign add_536511 = array_index_518710[11:2] + 10'h181;
  assign sel_536513 = $signed({1'h0, add_536127, array_index_518210[1:0]}) < $signed({1'h0, sel_536129}) ? {add_536127, array_index_518210[1:0]} : sel_536129;
  assign add_536515 = array_index_518713[11:2] + 10'h181;
  assign sel_536517 = $signed({1'h0, add_536131, array_index_518213[1:0]}) < $signed({1'h0, sel_536133}) ? {add_536131, array_index_518213[1:0]} : sel_536133;
  assign add_536529 = array_index_519786[11:0] + 12'h8a7;
  assign sel_536531 = $signed({1'h0, add_536145}) < $signed({1'h0, sel_536147}) ? add_536145 : sel_536147;
  assign add_536533 = array_index_519789[11:0] + 12'h8a7;
  assign sel_536535 = $signed({1'h0, add_536149}) < $signed({1'h0, sel_536151}) ? add_536149 : sel_536151;
  assign add_536547 = array_index_520964[11:1] + 11'h283;
  assign sel_536549 = $signed({1'h0, add_536163, array_index_520362[0]}) < $signed({1'h0, sel_536165}) ? {add_536163, array_index_520362[0]} : sel_536165;
  assign add_536551 = array_index_520967[11:1] + 11'h283;
  assign sel_536553 = $signed({1'h0, add_536167, array_index_520365[0]}) < $signed({1'h0, sel_536169}) ? {add_536167, array_index_520365[0]} : sel_536169;
  assign sel_536564 = ($signed({1'h0, add_535909}) < $signed({1'h0, sel_535911}) ? add_535909 : sel_535911) == ($signed({1'h0, add_535913}) < $signed({1'h0, sel_535915}) ? add_535913 : sel_535915) ? add_536439 : sel_536312;
  assign add_536571 = array_index_515726[11:2] + 10'h113;
  assign sel_536573 = $signed({1'h0, add_536195, array_index_515398[1:0]}) < $signed({1'h0, sel_536197}) ? {add_536195, array_index_515398[1:0]} : sel_536197;
  assign add_536575 = array_index_515729[11:2] + 10'h113;
  assign sel_536577 = $signed({1'h0, add_536199, array_index_515401[1:0]}) < $signed({1'h0, sel_536201}) ? {add_536199, array_index_515401[1:0]} : sel_536201;
  assign add_536589 = array_index_516458[11:4] + 8'h49;
  assign sel_536591 = $signed({1'h0, add_536213, array_index_516080[3:0]}) < $signed({1'h0, sel_536215}) ? {add_536213, array_index_516080[3:0]} : sel_536215;
  assign add_536593 = array_index_516461[11:4] + 8'h49;
  assign sel_536595 = $signed({1'h0, add_536217, array_index_516083[3:0]}) < $signed({1'h0, sel_536219}) ? {add_536217, array_index_516083[3:0]} : sel_536219;
  assign add_536605 = array_index_517286[11:0] + 12'h263;
  assign sel_536607 = $signed({1'h0, add_536229}) < $signed({1'h0, sel_536231}) ? add_536229 : sel_536231;
  assign add_536609 = array_index_517289[11:0] + 12'h263;
  assign sel_536611 = $signed({1'h0, add_536233}) < $signed({1'h0, sel_536235}) ? add_536233 : sel_536235;
  assign add_536621 = array_index_518210[11:1] + 11'h109;
  assign sel_536623 = $signed({1'h0, add_536245, array_index_517736[0]}) < $signed({1'h0, sel_536247}) ? {add_536245, array_index_517736[0]} : sel_536247;
  assign add_536625 = array_index_518213[11:1] + 11'h109;
  assign sel_536627 = $signed({1'h0, add_536249, array_index_517739[0]}) < $signed({1'h0, sel_536251}) ? {add_536249, array_index_517739[0]} : sel_536251;
  assign add_536637 = array_index_519236[11:3] + 9'h12f;
  assign sel_536639 = $signed({1'h0, add_536261, array_index_518710[2:0]}) < $signed({1'h0, sel_536263}) ? {add_536261, array_index_518710[2:0]} : sel_536263;
  assign add_536641 = array_index_519239[11:3] + 9'h12f;
  assign sel_536643 = $signed({1'h0, add_536265, array_index_518713[2:0]}) < $signed({1'h0, sel_536267}) ? {add_536265, array_index_518713[2:0]} : sel_536267;
  assign add_536655 = array_index_520362[11:3] + 9'h171;
  assign sel_536657 = $signed({1'h0, add_536279, array_index_519786[2:0]}) < $signed({1'h0, sel_536281}) ? {add_536279, array_index_519786[2:0]} : sel_536281;
  assign add_536659 = array_index_520365[11:3] + 9'h171;
  assign sel_536661 = $signed({1'h0, add_536283, array_index_519789[2:0]}) < $signed({1'h0, sel_536285}) ? {add_536283, array_index_519789[2:0]} : sel_536285;
  assign add_536671 = array_index_521590[11:0] + 12'h091;
  assign sel_536673 = $signed({1'h0, add_536295}) < $signed({1'h0, sel_536297}) ? add_536295 : sel_536297;
  assign add_536675 = array_index_521593[11:0] + 12'h091;
  assign sel_536677 = $signed({1'h0, add_536299}) < $signed({1'h0, sel_536301}) ? add_536299 : sel_536301;
  assign add_536681 = sel_536564 + 16'h0001;
  assign add_536691 = array_index_516080[11:1] + 11'h5b9;
  assign sel_536693 = $signed({1'h0, add_536323, array_index_515726[0]}) < $signed({1'h0, sel_536325}) ? {add_536323, array_index_515726[0]} : sel_536325;
  assign add_536695 = array_index_516083[11:1] + 11'h5b9;
  assign sel_536697 = $signed({1'h0, add_536327, array_index_515729[0]}) < $signed({1'h0, sel_536329}) ? {add_536327, array_index_515729[0]} : sel_536329;
  assign add_536707 = array_index_516860[11:0] + 12'h37b;
  assign sel_536709 = $signed({1'h0, add_536339}) < $signed({1'h0, sel_536341}) ? add_536339 : sel_536341;
  assign add_536711 = array_index_516863[11:0] + 12'h37b;
  assign sel_536713 = $signed({1'h0, add_536343}) < $signed({1'h0, sel_536345}) ? add_536343 : sel_536345;
  assign add_536725 = array_index_517736[11:0] + 12'h811;
  assign sel_536727 = $signed({1'h0, add_536357}) < $signed({1'h0, sel_536359}) ? add_536357 : sel_536359;
  assign add_536729 = array_index_517739[11:0] + 12'h811;
  assign sel_536731 = $signed({1'h0, add_536361}) < $signed({1'h0, sel_536363}) ? add_536361 : sel_536363;
  assign add_536743 = array_index_518710[11:0] + 12'h70f;
  assign sel_536745 = $signed({1'h0, add_536375}) < $signed({1'h0, sel_536377}) ? add_536375 : sel_536377;
  assign add_536747 = array_index_518713[11:0] + 12'h70f;
  assign sel_536749 = $signed({1'h0, add_536379}) < $signed({1'h0, sel_536381}) ? add_536379 : sel_536381;
  assign add_536761 = array_index_519786[11:3] + 9'h1f1;
  assign sel_536763 = $signed({1'h0, add_536393, array_index_519236[2:0]}) < $signed({1'h0, sel_536395}) ? {add_536393, array_index_519236[2:0]} : sel_536395;
  assign add_536765 = array_index_519789[11:3] + 9'h1f1;
  assign sel_536767 = $signed({1'h0, add_536397, array_index_519239[2:0]}) < $signed({1'h0, sel_536399}) ? {add_536397, array_index_519239[2:0]} : sel_536399;
  assign add_536777 = array_index_520964[11:0] + 12'h081;
  assign sel_536779 = $signed({1'h0, add_536409}) < $signed({1'h0, sel_536411}) ? add_536409 : sel_536411;
  assign add_536781 = array_index_520967[11:0] + 12'h081;
  assign sel_536783 = $signed({1'h0, add_536413}) < $signed({1'h0, sel_536415}) ? add_536413 : sel_536415;
  assign sel_536796 = ($signed({1'h0, add_536179, array_index_521590[0]}) < $signed({1'h0, sel_536181}) ? {add_536179, array_index_521590[0]} : sel_536181) == ($signed({1'h0, add_536183, array_index_521593[0]}) < $signed({1'h0, sel_536185}) ? {add_536183, array_index_521593[0]} : sel_536185) ? add_536681 : sel_536564;
  assign add_536799 = array_index_515726[11:0] + 12'hcc1;
  assign sel_536801 = $signed({1'h0, add_536441}) < $signed({1'h0, sel_536443}) ? add_536441 : sel_536443;
  assign add_536803 = array_index_515729[11:0] + 12'hcc1;
  assign sel_536805 = $signed({1'h0, add_536445}) < $signed({1'h0, sel_536447}) ? add_536445 : sel_536447;
  assign add_536817 = array_index_516458[11:0] + 12'ha87;
  assign sel_536819 = $signed({1'h0, add_536459}) < $signed({1'h0, sel_536461}) ? add_536459 : sel_536461;
  assign add_536821 = array_index_516461[11:0] + 12'ha87;
  assign sel_536823 = $signed({1'h0, add_536463}) < $signed({1'h0, sel_536465}) ? add_536463 : sel_536465;
  assign add_536835 = array_index_517286[11:1] + 11'h663;
  assign sel_536837 = $signed({1'h0, add_536477, array_index_516860[0]}) < $signed({1'h0, sel_536479}) ? {add_536477, array_index_516860[0]} : sel_536479;
  assign add_536839 = array_index_517289[11:1] + 11'h663;
  assign sel_536841 = $signed({1'h0, add_536481, array_index_516863[0]}) < $signed({1'h0, sel_536483}) ? {add_536481, array_index_516863[0]} : sel_536483;
  assign add_536851 = array_index_518210[11:1] + 11'h075;
  assign sel_536853 = $signed({1'h0, add_536493, array_index_517736[0]}) < $signed({1'h0, sel_536495}) ? {add_536493, array_index_517736[0]} : sel_536495;
  assign add_536855 = array_index_518213[11:1] + 11'h075;
  assign sel_536857 = $signed({1'h0, add_536497, array_index_517739[0]}) < $signed({1'h0, sel_536499}) ? {add_536497, array_index_517739[0]} : sel_536499;
  assign add_536869 = array_index_519236[11:2] + 10'h181;
  assign sel_536871 = $signed({1'h0, add_536511, array_index_518710[1:0]}) < $signed({1'h0, sel_536513}) ? {add_536511, array_index_518710[1:0]} : sel_536513;
  assign add_536873 = array_index_519239[11:2] + 10'h181;
  assign sel_536875 = $signed({1'h0, add_536515, array_index_518713[1:0]}) < $signed({1'h0, sel_536517}) ? {add_536515, array_index_518713[1:0]} : sel_536517;
  assign add_536887 = array_index_520362[11:0] + 12'h8a7;
  assign sel_536889 = $signed({1'h0, add_536529}) < $signed({1'h0, sel_536531}) ? add_536529 : sel_536531;
  assign add_536891 = array_index_520365[11:0] + 12'h8a7;
  assign sel_536893 = $signed({1'h0, add_536533}) < $signed({1'h0, sel_536535}) ? add_536533 : sel_536535;
  assign add_536905 = array_index_521590[11:1] + 11'h283;
  assign sel_536907 = $signed({1'h0, add_536547, array_index_520964[0]}) < $signed({1'h0, sel_536549}) ? {add_536547, array_index_520964[0]} : sel_536549;
  assign add_536909 = array_index_521593[11:1] + 11'h283;
  assign sel_536911 = $signed({1'h0, add_536551, array_index_520967[0]}) < $signed({1'h0, sel_536553}) ? {add_536551, array_index_520967[0]} : sel_536553;
  assign add_536915 = sel_536796 + 16'h0001;
  assign add_536921 = array_index_516080[11:2] + 10'h113;
  assign sel_536923 = $signed({1'h0, add_536571, array_index_515726[1:0]}) < $signed({1'h0, sel_536573}) ? {add_536571, array_index_515726[1:0]} : sel_536573;
  assign add_536925 = array_index_516083[11:2] + 10'h113;
  assign sel_536927 = $signed({1'h0, add_536575, array_index_515729[1:0]}) < $signed({1'h0, sel_536577}) ? {add_536575, array_index_515729[1:0]} : sel_536577;
  assign add_536939 = array_index_516860[11:4] + 8'h49;
  assign sel_536941 = $signed({1'h0, add_536589, array_index_516458[3:0]}) < $signed({1'h0, sel_536591}) ? {add_536589, array_index_516458[3:0]} : sel_536591;
  assign add_536943 = array_index_516863[11:4] + 8'h49;
  assign sel_536945 = $signed({1'h0, add_536593, array_index_516461[3:0]}) < $signed({1'h0, sel_536595}) ? {add_536593, array_index_516461[3:0]} : sel_536595;
  assign add_536955 = array_index_517736[11:0] + 12'h263;
  assign sel_536957 = $signed({1'h0, add_536605}) < $signed({1'h0, sel_536607}) ? add_536605 : sel_536607;
  assign add_536959 = array_index_517739[11:0] + 12'h263;
  assign sel_536961 = $signed({1'h0, add_536609}) < $signed({1'h0, sel_536611}) ? add_536609 : sel_536611;
  assign add_536971 = array_index_518710[11:1] + 11'h109;
  assign sel_536973 = $signed({1'h0, add_536621, array_index_518210[0]}) < $signed({1'h0, sel_536623}) ? {add_536621, array_index_518210[0]} : sel_536623;
  assign add_536975 = array_index_518713[11:1] + 11'h109;
  assign sel_536977 = $signed({1'h0, add_536625, array_index_518213[0]}) < $signed({1'h0, sel_536627}) ? {add_536625, array_index_518213[0]} : sel_536627;
  assign add_536987 = array_index_519786[11:3] + 9'h12f;
  assign sel_536989 = $signed({1'h0, add_536637, array_index_519236[2:0]}) < $signed({1'h0, sel_536639}) ? {add_536637, array_index_519236[2:0]} : sel_536639;
  assign add_536991 = array_index_519789[11:3] + 9'h12f;
  assign sel_536993 = $signed({1'h0, add_536641, array_index_519239[2:0]}) < $signed({1'h0, sel_536643}) ? {add_536641, array_index_519239[2:0]} : sel_536643;
  assign add_537005 = array_index_520964[11:3] + 9'h171;
  assign sel_537007 = $signed({1'h0, add_536655, array_index_520362[2:0]}) < $signed({1'h0, sel_536657}) ? {add_536655, array_index_520362[2:0]} : sel_536657;
  assign add_537009 = array_index_520967[11:3] + 9'h171;
  assign sel_537011 = $signed({1'h0, add_536659, array_index_520365[2:0]}) < $signed({1'h0, sel_536661}) ? {add_536659, array_index_520365[2:0]} : sel_536661;
  assign sel_537022 = ($signed({1'h0, add_536427}) < $signed({1'h0, sel_536429}) ? add_536427 : sel_536429) == ($signed({1'h0, add_536431}) < $signed({1'h0, sel_536433}) ? add_536431 : sel_536433) ? add_536915 : sel_536796;
  assign add_537033 = array_index_516458[11:1] + 11'h5b9;
  assign sel_537035 = $signed({1'h0, add_536691, array_index_516080[0]}) < $signed({1'h0, sel_536693}) ? {add_536691, array_index_516080[0]} : sel_536693;
  assign add_537037 = array_index_516461[11:1] + 11'h5b9;
  assign sel_537039 = $signed({1'h0, add_536695, array_index_516083[0]}) < $signed({1'h0, sel_536697}) ? {add_536695, array_index_516083[0]} : sel_536697;
  assign add_537049 = array_index_517286[11:0] + 12'h37b;
  assign sel_537051 = $signed({1'h0, add_536707}) < $signed({1'h0, sel_536709}) ? add_536707 : sel_536709;
  assign add_537053 = array_index_517289[11:0] + 12'h37b;
  assign sel_537055 = $signed({1'h0, add_536711}) < $signed({1'h0, sel_536713}) ? add_536711 : sel_536713;
  assign add_537067 = array_index_518210[11:0] + 12'h811;
  assign sel_537069 = $signed({1'h0, add_536725}) < $signed({1'h0, sel_536727}) ? add_536725 : sel_536727;
  assign add_537071 = array_index_518213[11:0] + 12'h811;
  assign sel_537073 = $signed({1'h0, add_536729}) < $signed({1'h0, sel_536731}) ? add_536729 : sel_536731;
  assign add_537085 = array_index_519236[11:0] + 12'h70f;
  assign sel_537087 = $signed({1'h0, add_536743}) < $signed({1'h0, sel_536745}) ? add_536743 : sel_536745;
  assign add_537089 = array_index_519239[11:0] + 12'h70f;
  assign sel_537091 = $signed({1'h0, add_536747}) < $signed({1'h0, sel_536749}) ? add_536747 : sel_536749;
  assign add_537103 = array_index_520362[11:3] + 9'h1f1;
  assign sel_537105 = $signed({1'h0, add_536761, array_index_519786[2:0]}) < $signed({1'h0, sel_536763}) ? {add_536761, array_index_519786[2:0]} : sel_536763;
  assign add_537107 = array_index_520365[11:3] + 9'h1f1;
  assign sel_537109 = $signed({1'h0, add_536765, array_index_519789[2:0]}) < $signed({1'h0, sel_536767}) ? {add_536765, array_index_519789[2:0]} : sel_536767;
  assign add_537119 = array_index_521590[11:0] + 12'h081;
  assign sel_537121 = $signed({1'h0, add_536777}) < $signed({1'h0, sel_536779}) ? add_536777 : sel_536779;
  assign add_537123 = array_index_521593[11:0] + 12'h081;
  assign sel_537125 = $signed({1'h0, add_536781}) < $signed({1'h0, sel_536783}) ? add_536781 : sel_536783;
  assign add_537131 = sel_537022 + 16'h0001;
  assign add_537133 = array_index_516080[11:0] + 12'hcc1;
  assign sel_537135 = $signed({1'h0, add_536799}) < $signed({1'h0, sel_536801}) ? add_536799 : sel_536801;
  assign add_537137 = array_index_516083[11:0] + 12'hcc1;
  assign sel_537139 = $signed({1'h0, add_536803}) < $signed({1'h0, sel_536805}) ? add_536803 : sel_536805;
  assign add_537151 = array_index_516860[11:0] + 12'ha87;
  assign sel_537153 = $signed({1'h0, add_536817}) < $signed({1'h0, sel_536819}) ? add_536817 : sel_536819;
  assign add_537155 = array_index_516863[11:0] + 12'ha87;
  assign sel_537157 = $signed({1'h0, add_536821}) < $signed({1'h0, sel_536823}) ? add_536821 : sel_536823;
  assign add_537169 = array_index_517736[11:1] + 11'h663;
  assign sel_537171 = $signed({1'h0, add_536835, array_index_517286[0]}) < $signed({1'h0, sel_536837}) ? {add_536835, array_index_517286[0]} : sel_536837;
  assign add_537173 = array_index_517739[11:1] + 11'h663;
  assign sel_537175 = $signed({1'h0, add_536839, array_index_517289[0]}) < $signed({1'h0, sel_536841}) ? {add_536839, array_index_517289[0]} : sel_536841;
  assign add_537185 = array_index_518710[11:1] + 11'h075;
  assign sel_537187 = $signed({1'h0, add_536851, array_index_518210[0]}) < $signed({1'h0, sel_536853}) ? {add_536851, array_index_518210[0]} : sel_536853;
  assign add_537189 = array_index_518713[11:1] + 11'h075;
  assign sel_537191 = $signed({1'h0, add_536855, array_index_518213[0]}) < $signed({1'h0, sel_536857}) ? {add_536855, array_index_518213[0]} : sel_536857;
  assign add_537203 = array_index_519786[11:2] + 10'h181;
  assign sel_537205 = $signed({1'h0, add_536869, array_index_519236[1:0]}) < $signed({1'h0, sel_536871}) ? {add_536869, array_index_519236[1:0]} : sel_536871;
  assign add_537207 = array_index_519789[11:2] + 10'h181;
  assign sel_537209 = $signed({1'h0, add_536873, array_index_519239[1:0]}) < $signed({1'h0, sel_536875}) ? {add_536873, array_index_519239[1:0]} : sel_536875;
  assign add_537221 = array_index_520964[11:0] + 12'h8a7;
  assign sel_537223 = $signed({1'h0, add_536887}) < $signed({1'h0, sel_536889}) ? add_536887 : sel_536889;
  assign add_537225 = array_index_520967[11:0] + 12'h8a7;
  assign sel_537227 = $signed({1'h0, add_536891}) < $signed({1'h0, sel_536893}) ? add_536891 : sel_536893;
  assign sel_537240 = ($signed({1'h0, add_536671}) < $signed({1'h0, sel_536673}) ? add_536671 : sel_536673) == ($signed({1'h0, add_536675}) < $signed({1'h0, sel_536677}) ? add_536675 : sel_536677) ? add_537131 : sel_537022;
  assign add_537247 = array_index_516458[11:2] + 10'h113;
  assign sel_537249 = $signed({1'h0, add_536921, array_index_516080[1:0]}) < $signed({1'h0, sel_536923}) ? {add_536921, array_index_516080[1:0]} : sel_536923;
  assign add_537251 = array_index_516461[11:2] + 10'h113;
  assign sel_537253 = $signed({1'h0, add_536925, array_index_516083[1:0]}) < $signed({1'h0, sel_536927}) ? {add_536925, array_index_516083[1:0]} : sel_536927;
  assign add_537265 = array_index_517286[11:4] + 8'h49;
  assign sel_537267 = $signed({1'h0, add_536939, array_index_516860[3:0]}) < $signed({1'h0, sel_536941}) ? {add_536939, array_index_516860[3:0]} : sel_536941;
  assign add_537269 = array_index_517289[11:4] + 8'h49;
  assign sel_537271 = $signed({1'h0, add_536943, array_index_516863[3:0]}) < $signed({1'h0, sel_536945}) ? {add_536943, array_index_516863[3:0]} : sel_536945;
  assign add_537281 = array_index_518210[11:0] + 12'h263;
  assign sel_537283 = $signed({1'h0, add_536955}) < $signed({1'h0, sel_536957}) ? add_536955 : sel_536957;
  assign add_537285 = array_index_518213[11:0] + 12'h263;
  assign sel_537287 = $signed({1'h0, add_536959}) < $signed({1'h0, sel_536961}) ? add_536959 : sel_536961;
  assign add_537297 = array_index_519236[11:1] + 11'h109;
  assign sel_537299 = $signed({1'h0, add_536971, array_index_518710[0]}) < $signed({1'h0, sel_536973}) ? {add_536971, array_index_518710[0]} : sel_536973;
  assign add_537301 = array_index_519239[11:1] + 11'h109;
  assign sel_537303 = $signed({1'h0, add_536975, array_index_518713[0]}) < $signed({1'h0, sel_536977}) ? {add_536975, array_index_518713[0]} : sel_536977;
  assign add_537313 = array_index_520362[11:3] + 9'h12f;
  assign sel_537315 = $signed({1'h0, add_536987, array_index_519786[2:0]}) < $signed({1'h0, sel_536989}) ? {add_536987, array_index_519786[2:0]} : sel_536989;
  assign add_537317 = array_index_520365[11:3] + 9'h12f;
  assign sel_537319 = $signed({1'h0, add_536991, array_index_519789[2:0]}) < $signed({1'h0, sel_536993}) ? {add_536991, array_index_519789[2:0]} : sel_536993;
  assign add_537331 = array_index_521590[11:3] + 9'h171;
  assign sel_537333 = $signed({1'h0, add_537005, array_index_520964[2:0]}) < $signed({1'h0, sel_537007}) ? {add_537005, array_index_520964[2:0]} : sel_537007;
  assign add_537335 = array_index_521593[11:3] + 9'h171;
  assign sel_537337 = $signed({1'h0, add_537009, array_index_520967[2:0]}) < $signed({1'h0, sel_537011}) ? {add_537009, array_index_520967[2:0]} : sel_537011;
  assign add_537341 = sel_537240 + 16'h0001;
  assign add_537351 = array_index_516860[11:1] + 11'h5b9;
  assign sel_537353 = $signed({1'h0, add_537033, array_index_516458[0]}) < $signed({1'h0, sel_537035}) ? {add_537033, array_index_516458[0]} : sel_537035;
  assign add_537355 = array_index_516863[11:1] + 11'h5b9;
  assign sel_537357 = $signed({1'h0, add_537037, array_index_516461[0]}) < $signed({1'h0, sel_537039}) ? {add_537037, array_index_516461[0]} : sel_537039;
  assign add_537367 = array_index_517736[11:0] + 12'h37b;
  assign sel_537369 = $signed({1'h0, add_537049}) < $signed({1'h0, sel_537051}) ? add_537049 : sel_537051;
  assign add_537371 = array_index_517739[11:0] + 12'h37b;
  assign sel_537373 = $signed({1'h0, add_537053}) < $signed({1'h0, sel_537055}) ? add_537053 : sel_537055;
  assign add_537385 = array_index_518710[11:0] + 12'h811;
  assign sel_537387 = $signed({1'h0, add_537067}) < $signed({1'h0, sel_537069}) ? add_537067 : sel_537069;
  assign add_537389 = array_index_518713[11:0] + 12'h811;
  assign sel_537391 = $signed({1'h0, add_537071}) < $signed({1'h0, sel_537073}) ? add_537071 : sel_537073;
  assign add_537403 = array_index_519786[11:0] + 12'h70f;
  assign sel_537405 = $signed({1'h0, add_537085}) < $signed({1'h0, sel_537087}) ? add_537085 : sel_537087;
  assign add_537407 = array_index_519789[11:0] + 12'h70f;
  assign sel_537409 = $signed({1'h0, add_537089}) < $signed({1'h0, sel_537091}) ? add_537089 : sel_537091;
  assign add_537421 = array_index_520964[11:3] + 9'h1f1;
  assign sel_537423 = $signed({1'h0, add_537103, array_index_520362[2:0]}) < $signed({1'h0, sel_537105}) ? {add_537103, array_index_520362[2:0]} : sel_537105;
  assign add_537425 = array_index_520967[11:3] + 9'h1f1;
  assign sel_537427 = $signed({1'h0, add_537107, array_index_520365[2:0]}) < $signed({1'h0, sel_537109}) ? {add_537107, array_index_520365[2:0]} : sel_537109;
  assign sel_537438 = ($signed({1'h0, add_536905, array_index_521590[0]}) < $signed({1'h0, sel_536907}) ? {add_536905, array_index_521590[0]} : sel_536907) == ($signed({1'h0, add_536909, array_index_521593[0]}) < $signed({1'h0, sel_536911}) ? {add_536909, array_index_521593[0]} : sel_536911) ? add_537341 : sel_537240;
  assign add_537441 = array_index_516458[11:0] + 12'hcc1;
  assign sel_537443 = $signed({1'h0, add_537133}) < $signed({1'h0, sel_537135}) ? add_537133 : sel_537135;
  assign add_537445 = array_index_516461[11:0] + 12'hcc1;
  assign sel_537447 = $signed({1'h0, add_537137}) < $signed({1'h0, sel_537139}) ? add_537137 : sel_537139;
  assign add_537459 = array_index_517286[11:0] + 12'ha87;
  assign sel_537461 = $signed({1'h0, add_537151}) < $signed({1'h0, sel_537153}) ? add_537151 : sel_537153;
  assign add_537463 = array_index_517289[11:0] + 12'ha87;
  assign sel_537465 = $signed({1'h0, add_537155}) < $signed({1'h0, sel_537157}) ? add_537155 : sel_537157;
  assign add_537477 = array_index_518210[11:1] + 11'h663;
  assign sel_537479 = $signed({1'h0, add_537169, array_index_517736[0]}) < $signed({1'h0, sel_537171}) ? {add_537169, array_index_517736[0]} : sel_537171;
  assign add_537481 = array_index_518213[11:1] + 11'h663;
  assign sel_537483 = $signed({1'h0, add_537173, array_index_517739[0]}) < $signed({1'h0, sel_537175}) ? {add_537173, array_index_517739[0]} : sel_537175;
  assign add_537493 = array_index_519236[11:1] + 11'h075;
  assign sel_537495 = $signed({1'h0, add_537185, array_index_518710[0]}) < $signed({1'h0, sel_537187}) ? {add_537185, array_index_518710[0]} : sel_537187;
  assign add_537497 = array_index_519239[11:1] + 11'h075;
  assign sel_537499 = $signed({1'h0, add_537189, array_index_518713[0]}) < $signed({1'h0, sel_537191}) ? {add_537189, array_index_518713[0]} : sel_537191;
  assign add_537511 = array_index_520362[11:2] + 10'h181;
  assign sel_537513 = $signed({1'h0, add_537203, array_index_519786[1:0]}) < $signed({1'h0, sel_537205}) ? {add_537203, array_index_519786[1:0]} : sel_537205;
  assign add_537515 = array_index_520365[11:2] + 10'h181;
  assign sel_537517 = $signed({1'h0, add_537207, array_index_519789[1:0]}) < $signed({1'h0, sel_537209}) ? {add_537207, array_index_519789[1:0]} : sel_537209;
  assign add_537529 = array_index_521590[11:0] + 12'h8a7;
  assign sel_537531 = $signed({1'h0, add_537221}) < $signed({1'h0, sel_537223}) ? add_537221 : sel_537223;
  assign add_537533 = array_index_521593[11:0] + 12'h8a7;
  assign sel_537535 = $signed({1'h0, add_537225}) < $signed({1'h0, sel_537227}) ? add_537225 : sel_537227;
  assign add_537541 = sel_537438 + 16'h0001;
  assign add_537547 = array_index_516860[11:2] + 10'h113;
  assign sel_537549 = $signed({1'h0, add_537247, array_index_516458[1:0]}) < $signed({1'h0, sel_537249}) ? {add_537247, array_index_516458[1:0]} : sel_537249;
  assign add_537551 = array_index_516863[11:2] + 10'h113;
  assign sel_537553 = $signed({1'h0, add_537251, array_index_516461[1:0]}) < $signed({1'h0, sel_537253}) ? {add_537251, array_index_516461[1:0]} : sel_537253;
  assign add_537565 = array_index_517736[11:4] + 8'h49;
  assign sel_537567 = $signed({1'h0, add_537265, array_index_517286[3:0]}) < $signed({1'h0, sel_537267}) ? {add_537265, array_index_517286[3:0]} : sel_537267;
  assign add_537569 = array_index_517739[11:4] + 8'h49;
  assign sel_537571 = $signed({1'h0, add_537269, array_index_517289[3:0]}) < $signed({1'h0, sel_537271}) ? {add_537269, array_index_517289[3:0]} : sel_537271;
  assign add_537581 = array_index_518710[11:0] + 12'h263;
  assign sel_537583 = $signed({1'h0, add_537281}) < $signed({1'h0, sel_537283}) ? add_537281 : sel_537283;
  assign add_537585 = array_index_518713[11:0] + 12'h263;
  assign sel_537587 = $signed({1'h0, add_537285}) < $signed({1'h0, sel_537287}) ? add_537285 : sel_537287;
  assign add_537597 = array_index_519786[11:1] + 11'h109;
  assign sel_537599 = $signed({1'h0, add_537297, array_index_519236[0]}) < $signed({1'h0, sel_537299}) ? {add_537297, array_index_519236[0]} : sel_537299;
  assign add_537601 = array_index_519789[11:1] + 11'h109;
  assign sel_537603 = $signed({1'h0, add_537301, array_index_519239[0]}) < $signed({1'h0, sel_537303}) ? {add_537301, array_index_519239[0]} : sel_537303;
  assign add_537613 = array_index_520964[11:3] + 9'h12f;
  assign sel_537615 = $signed({1'h0, add_537313, array_index_520362[2:0]}) < $signed({1'h0, sel_537315}) ? {add_537313, array_index_520362[2:0]} : sel_537315;
  assign add_537617 = array_index_520967[11:3] + 9'h12f;
  assign sel_537619 = $signed({1'h0, add_537317, array_index_520365[2:0]}) < $signed({1'h0, sel_537319}) ? {add_537317, array_index_520365[2:0]} : sel_537319;
  assign sel_537632 = ($signed({1'h0, add_537119}) < $signed({1'h0, sel_537121}) ? add_537119 : sel_537121) == ($signed({1'h0, add_537123}) < $signed({1'h0, sel_537125}) ? add_537123 : sel_537125) ? add_537541 : sel_537438;
  assign add_537643 = array_index_517286[11:1] + 11'h5b9;
  assign sel_537645 = $signed({1'h0, add_537351, array_index_516860[0]}) < $signed({1'h0, sel_537353}) ? {add_537351, array_index_516860[0]} : sel_537353;
  assign add_537647 = array_index_517289[11:1] + 11'h5b9;
  assign sel_537649 = $signed({1'h0, add_537355, array_index_516863[0]}) < $signed({1'h0, sel_537357}) ? {add_537355, array_index_516863[0]} : sel_537357;
  assign add_537659 = array_index_518210[11:0] + 12'h37b;
  assign sel_537661 = $signed({1'h0, add_537367}) < $signed({1'h0, sel_537369}) ? add_537367 : sel_537369;
  assign add_537663 = array_index_518213[11:0] + 12'h37b;
  assign sel_537665 = $signed({1'h0, add_537371}) < $signed({1'h0, sel_537373}) ? add_537371 : sel_537373;
  assign add_537677 = array_index_519236[11:0] + 12'h811;
  assign sel_537679 = $signed({1'h0, add_537385}) < $signed({1'h0, sel_537387}) ? add_537385 : sel_537387;
  assign add_537681 = array_index_519239[11:0] + 12'h811;
  assign sel_537683 = $signed({1'h0, add_537389}) < $signed({1'h0, sel_537391}) ? add_537389 : sel_537391;
  assign add_537695 = array_index_520362[11:0] + 12'h70f;
  assign sel_537697 = $signed({1'h0, add_537403}) < $signed({1'h0, sel_537405}) ? add_537403 : sel_537405;
  assign add_537699 = array_index_520365[11:0] + 12'h70f;
  assign sel_537701 = $signed({1'h0, add_537407}) < $signed({1'h0, sel_537409}) ? add_537407 : sel_537409;
  assign add_537713 = array_index_521590[11:3] + 9'h1f1;
  assign sel_537715 = $signed({1'h0, add_537421, array_index_520964[2:0]}) < $signed({1'h0, sel_537423}) ? {add_537421, array_index_520964[2:0]} : sel_537423;
  assign add_537717 = array_index_521593[11:3] + 9'h1f1;
  assign sel_537719 = $signed({1'h0, add_537425, array_index_520967[2:0]}) < $signed({1'h0, sel_537427}) ? {add_537425, array_index_520967[2:0]} : sel_537427;
  assign add_537723 = sel_537632 + 16'h0001;
  assign add_537725 = array_index_516860[11:0] + 12'hcc1;
  assign sel_537727 = $signed({1'h0, add_537441}) < $signed({1'h0, sel_537443}) ? add_537441 : sel_537443;
  assign add_537729 = array_index_516863[11:0] + 12'hcc1;
  assign sel_537731 = $signed({1'h0, add_537445}) < $signed({1'h0, sel_537447}) ? add_537445 : sel_537447;
  assign add_537743 = array_index_517736[11:0] + 12'ha87;
  assign sel_537745 = $signed({1'h0, add_537459}) < $signed({1'h0, sel_537461}) ? add_537459 : sel_537461;
  assign add_537747 = array_index_517739[11:0] + 12'ha87;
  assign sel_537749 = $signed({1'h0, add_537463}) < $signed({1'h0, sel_537465}) ? add_537463 : sel_537465;
  assign add_537761 = array_index_518710[11:1] + 11'h663;
  assign sel_537763 = $signed({1'h0, add_537477, array_index_518210[0]}) < $signed({1'h0, sel_537479}) ? {add_537477, array_index_518210[0]} : sel_537479;
  assign add_537765 = array_index_518713[11:1] + 11'h663;
  assign sel_537767 = $signed({1'h0, add_537481, array_index_518213[0]}) < $signed({1'h0, sel_537483}) ? {add_537481, array_index_518213[0]} : sel_537483;
  assign add_537777 = array_index_519786[11:1] + 11'h075;
  assign sel_537779 = $signed({1'h0, add_537493, array_index_519236[0]}) < $signed({1'h0, sel_537495}) ? {add_537493, array_index_519236[0]} : sel_537495;
  assign add_537781 = array_index_519789[11:1] + 11'h075;
  assign sel_537783 = $signed({1'h0, add_537497, array_index_519239[0]}) < $signed({1'h0, sel_537499}) ? {add_537497, array_index_519239[0]} : sel_537499;
  assign add_537795 = array_index_520964[11:2] + 10'h181;
  assign sel_537797 = $signed({1'h0, add_537511, array_index_520362[1:0]}) < $signed({1'h0, sel_537513}) ? {add_537511, array_index_520362[1:0]} : sel_537513;
  assign add_537799 = array_index_520967[11:2] + 10'h181;
  assign sel_537801 = $signed({1'h0, add_537515, array_index_520365[1:0]}) < $signed({1'h0, sel_537517}) ? {add_537515, array_index_520365[1:0]} : sel_537517;
  assign sel_537814 = ($signed({1'h0, add_537331, array_index_521590[2:0]}) < $signed({1'h0, sel_537333}) ? {add_537331, array_index_521590[2:0]} : sel_537333) == ($signed({1'h0, add_537335, array_index_521593[2:0]}) < $signed({1'h0, sel_537337}) ? {add_537335, array_index_521593[2:0]} : sel_537337) ? add_537723 : sel_537632;
  assign add_537821 = array_index_517286[11:2] + 10'h113;
  assign sel_537823 = $signed({1'h0, add_537547, array_index_516860[1:0]}) < $signed({1'h0, sel_537549}) ? {add_537547, array_index_516860[1:0]} : sel_537549;
  assign add_537825 = array_index_517289[11:2] + 10'h113;
  assign sel_537827 = $signed({1'h0, add_537551, array_index_516863[1:0]}) < $signed({1'h0, sel_537553}) ? {add_537551, array_index_516863[1:0]} : sel_537553;
  assign add_537839 = array_index_518210[11:4] + 8'h49;
  assign sel_537841 = $signed({1'h0, add_537565, array_index_517736[3:0]}) < $signed({1'h0, sel_537567}) ? {add_537565, array_index_517736[3:0]} : sel_537567;
  assign add_537843 = array_index_518213[11:4] + 8'h49;
  assign sel_537845 = $signed({1'h0, add_537569, array_index_517739[3:0]}) < $signed({1'h0, sel_537571}) ? {add_537569, array_index_517739[3:0]} : sel_537571;
  assign add_537855 = array_index_519236[11:0] + 12'h263;
  assign sel_537857 = $signed({1'h0, add_537581}) < $signed({1'h0, sel_537583}) ? add_537581 : sel_537583;
  assign add_537859 = array_index_519239[11:0] + 12'h263;
  assign sel_537861 = $signed({1'h0, add_537585}) < $signed({1'h0, sel_537587}) ? add_537585 : sel_537587;
  assign add_537871 = array_index_520362[11:1] + 11'h109;
  assign sel_537873 = $signed({1'h0, add_537597, array_index_519786[0]}) < $signed({1'h0, sel_537599}) ? {add_537597, array_index_519786[0]} : sel_537599;
  assign add_537875 = array_index_520365[11:1] + 11'h109;
  assign sel_537877 = $signed({1'h0, add_537601, array_index_519789[0]}) < $signed({1'h0, sel_537603}) ? {add_537601, array_index_519789[0]} : sel_537603;
  assign add_537887 = array_index_521590[11:3] + 9'h12f;
  assign sel_537889 = $signed({1'h0, add_537613, array_index_520964[2:0]}) < $signed({1'h0, sel_537615}) ? {add_537613, array_index_520964[2:0]} : sel_537615;
  assign add_537891 = array_index_521593[11:3] + 9'h12f;
  assign sel_537893 = $signed({1'h0, add_537617, array_index_520967[2:0]}) < $signed({1'h0, sel_537619}) ? {add_537617, array_index_520967[2:0]} : sel_537619;
  assign add_537899 = sel_537814 + 16'h0001;
  assign add_537909 = array_index_517736[11:1] + 11'h5b9;
  assign sel_537911 = $signed({1'h0, add_537643, array_index_517286[0]}) < $signed({1'h0, sel_537645}) ? {add_537643, array_index_517286[0]} : sel_537645;
  assign add_537913 = array_index_517739[11:1] + 11'h5b9;
  assign sel_537915 = $signed({1'h0, add_537647, array_index_517289[0]}) < $signed({1'h0, sel_537649}) ? {add_537647, array_index_517289[0]} : sel_537649;
  assign add_537925 = array_index_518710[11:0] + 12'h37b;
  assign sel_537927 = $signed({1'h0, add_537659}) < $signed({1'h0, sel_537661}) ? add_537659 : sel_537661;
  assign add_537929 = array_index_518713[11:0] + 12'h37b;
  assign sel_537931 = $signed({1'h0, add_537663}) < $signed({1'h0, sel_537665}) ? add_537663 : sel_537665;
  assign add_537943 = array_index_519786[11:0] + 12'h811;
  assign sel_537945 = $signed({1'h0, add_537677}) < $signed({1'h0, sel_537679}) ? add_537677 : sel_537679;
  assign add_537947 = array_index_519789[11:0] + 12'h811;
  assign sel_537949 = $signed({1'h0, add_537681}) < $signed({1'h0, sel_537683}) ? add_537681 : sel_537683;
  assign add_537961 = array_index_520964[11:0] + 12'h70f;
  assign sel_537963 = $signed({1'h0, add_537695}) < $signed({1'h0, sel_537697}) ? add_537695 : sel_537697;
  assign add_537965 = array_index_520967[11:0] + 12'h70f;
  assign sel_537967 = $signed({1'h0, add_537699}) < $signed({1'h0, sel_537701}) ? add_537699 : sel_537701;
  assign sel_537980 = ($signed({1'h0, add_537529}) < $signed({1'h0, sel_537531}) ? add_537529 : sel_537531) == ($signed({1'h0, add_537533}) < $signed({1'h0, sel_537535}) ? add_537533 : sel_537535) ? add_537899 : sel_537814;
  assign add_537983 = array_index_517286[11:0] + 12'hcc1;
  assign sel_537985 = $signed({1'h0, add_537725}) < $signed({1'h0, sel_537727}) ? add_537725 : sel_537727;
  assign add_537987 = array_index_517289[11:0] + 12'hcc1;
  assign sel_537989 = $signed({1'h0, add_537729}) < $signed({1'h0, sel_537731}) ? add_537729 : sel_537731;
  assign add_538001 = array_index_518210[11:0] + 12'ha87;
  assign sel_538003 = $signed({1'h0, add_537743}) < $signed({1'h0, sel_537745}) ? add_537743 : sel_537745;
  assign add_538005 = array_index_518213[11:0] + 12'ha87;
  assign sel_538007 = $signed({1'h0, add_537747}) < $signed({1'h0, sel_537749}) ? add_537747 : sel_537749;
  assign add_538019 = array_index_519236[11:1] + 11'h663;
  assign sel_538021 = $signed({1'h0, add_537761, array_index_518710[0]}) < $signed({1'h0, sel_537763}) ? {add_537761, array_index_518710[0]} : sel_537763;
  assign add_538023 = array_index_519239[11:1] + 11'h663;
  assign sel_538025 = $signed({1'h0, add_537765, array_index_518713[0]}) < $signed({1'h0, sel_537767}) ? {add_537765, array_index_518713[0]} : sel_537767;
  assign add_538035 = array_index_520362[11:1] + 11'h075;
  assign sel_538037 = $signed({1'h0, add_537777, array_index_519786[0]}) < $signed({1'h0, sel_537779}) ? {add_537777, array_index_519786[0]} : sel_537779;
  assign add_538039 = array_index_520365[11:1] + 11'h075;
  assign sel_538041 = $signed({1'h0, add_537781, array_index_519789[0]}) < $signed({1'h0, sel_537783}) ? {add_537781, array_index_519789[0]} : sel_537783;
  assign add_538053 = array_index_521590[11:2] + 10'h181;
  assign sel_538055 = $signed({1'h0, add_537795, array_index_520964[1:0]}) < $signed({1'h0, sel_537797}) ? {add_537795, array_index_520964[1:0]} : sel_537797;
  assign add_538057 = array_index_521593[11:2] + 10'h181;
  assign sel_538059 = $signed({1'h0, add_537799, array_index_520967[1:0]}) < $signed({1'h0, sel_537801}) ? {add_537799, array_index_520967[1:0]} : sel_537801;
  assign add_538065 = sel_537980 + 16'h0001;
  assign add_538071 = array_index_517736[11:2] + 10'h113;
  assign sel_538073 = $signed({1'h0, add_537821, array_index_517286[1:0]}) < $signed({1'h0, sel_537823}) ? {add_537821, array_index_517286[1:0]} : sel_537823;
  assign add_538075 = array_index_517739[11:2] + 10'h113;
  assign sel_538077 = $signed({1'h0, add_537825, array_index_517289[1:0]}) < $signed({1'h0, sel_537827}) ? {add_537825, array_index_517289[1:0]} : sel_537827;
  assign add_538089 = array_index_518710[11:4] + 8'h49;
  assign sel_538091 = $signed({1'h0, add_537839, array_index_518210[3:0]}) < $signed({1'h0, sel_537841}) ? {add_537839, array_index_518210[3:0]} : sel_537841;
  assign add_538093 = array_index_518713[11:4] + 8'h49;
  assign sel_538095 = $signed({1'h0, add_537843, array_index_518213[3:0]}) < $signed({1'h0, sel_537845}) ? {add_537843, array_index_518213[3:0]} : sel_537845;
  assign add_538105 = array_index_519786[11:0] + 12'h263;
  assign sel_538107 = $signed({1'h0, add_537855}) < $signed({1'h0, sel_537857}) ? add_537855 : sel_537857;
  assign add_538109 = array_index_519789[11:0] + 12'h263;
  assign sel_538111 = $signed({1'h0, add_537859}) < $signed({1'h0, sel_537861}) ? add_537859 : sel_537861;
  assign add_538121 = array_index_520964[11:1] + 11'h109;
  assign sel_538123 = $signed({1'h0, add_537871, array_index_520362[0]}) < $signed({1'h0, sel_537873}) ? {add_537871, array_index_520362[0]} : sel_537873;
  assign add_538125 = array_index_520967[11:1] + 11'h109;
  assign sel_538127 = $signed({1'h0, add_537875, array_index_520365[0]}) < $signed({1'h0, sel_537877}) ? {add_537875, array_index_520365[0]} : sel_537877;
  assign sel_538138 = ($signed({1'h0, add_537713, array_index_521590[2:0]}) < $signed({1'h0, sel_537715}) ? {add_537713, array_index_521590[2:0]} : sel_537715) == ($signed({1'h0, add_537717, array_index_521593[2:0]}) < $signed({1'h0, sel_537719}) ? {add_537717, array_index_521593[2:0]} : sel_537719) ? add_538065 : sel_537980;
  assign add_538149 = array_index_518210[11:1] + 11'h5b9;
  assign sel_538151 = $signed({1'h0, add_537909, array_index_517736[0]}) < $signed({1'h0, sel_537911}) ? {add_537909, array_index_517736[0]} : sel_537911;
  assign add_538153 = array_index_518213[11:1] + 11'h5b9;
  assign sel_538155 = $signed({1'h0, add_537913, array_index_517739[0]}) < $signed({1'h0, sel_537915}) ? {add_537913, array_index_517739[0]} : sel_537915;
  assign add_538165 = array_index_519236[11:0] + 12'h37b;
  assign sel_538167 = $signed({1'h0, add_537925}) < $signed({1'h0, sel_537927}) ? add_537925 : sel_537927;
  assign add_538169 = array_index_519239[11:0] + 12'h37b;
  assign sel_538171 = $signed({1'h0, add_537929}) < $signed({1'h0, sel_537931}) ? add_537929 : sel_537931;
  assign add_538183 = array_index_520362[11:0] + 12'h811;
  assign sel_538185 = $signed({1'h0, add_537943}) < $signed({1'h0, sel_537945}) ? add_537943 : sel_537945;
  assign add_538187 = array_index_520365[11:0] + 12'h811;
  assign sel_538189 = $signed({1'h0, add_537947}) < $signed({1'h0, sel_537949}) ? add_537947 : sel_537949;
  assign add_538201 = array_index_521590[11:0] + 12'h70f;
  assign sel_538203 = $signed({1'h0, add_537961}) < $signed({1'h0, sel_537963}) ? add_537961 : sel_537963;
  assign add_538205 = array_index_521593[11:0] + 12'h70f;
  assign sel_538207 = $signed({1'h0, add_537965}) < $signed({1'h0, sel_537967}) ? add_537965 : sel_537967;
  assign add_538213 = sel_538138 + 16'h0001;
  assign add_538215 = array_index_517736[11:0] + 12'hcc1;
  assign sel_538217 = $signed({1'h0, add_537983}) < $signed({1'h0, sel_537985}) ? add_537983 : sel_537985;
  assign add_538219 = array_index_517739[11:0] + 12'hcc1;
  assign sel_538221 = $signed({1'h0, add_537987}) < $signed({1'h0, sel_537989}) ? add_537987 : sel_537989;
  assign add_538233 = array_index_518710[11:0] + 12'ha87;
  assign sel_538235 = $signed({1'h0, add_538001}) < $signed({1'h0, sel_538003}) ? add_538001 : sel_538003;
  assign add_538237 = array_index_518713[11:0] + 12'ha87;
  assign sel_538239 = $signed({1'h0, add_538005}) < $signed({1'h0, sel_538007}) ? add_538005 : sel_538007;
  assign add_538251 = array_index_519786[11:1] + 11'h663;
  assign sel_538253 = $signed({1'h0, add_538019, array_index_519236[0]}) < $signed({1'h0, sel_538021}) ? {add_538019, array_index_519236[0]} : sel_538021;
  assign add_538255 = array_index_519789[11:1] + 11'h663;
  assign sel_538257 = $signed({1'h0, add_538023, array_index_519239[0]}) < $signed({1'h0, sel_538025}) ? {add_538023, array_index_519239[0]} : sel_538025;
  assign add_538267 = array_index_520964[11:1] + 11'h075;
  assign sel_538269 = $signed({1'h0, add_538035, array_index_520362[0]}) < $signed({1'h0, sel_538037}) ? {add_538035, array_index_520362[0]} : sel_538037;
  assign add_538271 = array_index_520967[11:1] + 11'h075;
  assign sel_538273 = $signed({1'h0, add_538039, array_index_520365[0]}) < $signed({1'h0, sel_538041}) ? {add_538039, array_index_520365[0]} : sel_538041;
  assign sel_538286 = ($signed({1'h0, add_537887, array_index_521590[2:0]}) < $signed({1'h0, sel_537889}) ? {add_537887, array_index_521590[2:0]} : sel_537889) == ($signed({1'h0, add_537891, array_index_521593[2:0]}) < $signed({1'h0, sel_537893}) ? {add_537891, array_index_521593[2:0]} : sel_537893) ? add_538213 : sel_538138;
  assign add_538293 = array_index_518210[11:2] + 10'h113;
  assign sel_538295 = $signed({1'h0, add_538071, array_index_517736[1:0]}) < $signed({1'h0, sel_538073}) ? {add_538071, array_index_517736[1:0]} : sel_538073;
  assign add_538297 = array_index_518213[11:2] + 10'h113;
  assign sel_538299 = $signed({1'h0, add_538075, array_index_517739[1:0]}) < $signed({1'h0, sel_538077}) ? {add_538075, array_index_517739[1:0]} : sel_538077;
  assign add_538311 = array_index_519236[11:4] + 8'h49;
  assign sel_538313 = $signed({1'h0, add_538089, array_index_518710[3:0]}) < $signed({1'h0, sel_538091}) ? {add_538089, array_index_518710[3:0]} : sel_538091;
  assign add_538315 = array_index_519239[11:4] + 8'h49;
  assign sel_538317 = $signed({1'h0, add_538093, array_index_518713[3:0]}) < $signed({1'h0, sel_538095}) ? {add_538093, array_index_518713[3:0]} : sel_538095;
  assign add_538327 = array_index_520362[11:0] + 12'h263;
  assign sel_538329 = $signed({1'h0, add_538105}) < $signed({1'h0, sel_538107}) ? add_538105 : sel_538107;
  assign add_538331 = array_index_520365[11:0] + 12'h263;
  assign sel_538333 = $signed({1'h0, add_538109}) < $signed({1'h0, sel_538111}) ? add_538109 : sel_538111;
  assign add_538343 = array_index_521590[11:1] + 11'h109;
  assign sel_538345 = $signed({1'h0, add_538121, array_index_520964[0]}) < $signed({1'h0, sel_538123}) ? {add_538121, array_index_520964[0]} : sel_538123;
  assign add_538347 = array_index_521593[11:1] + 11'h109;
  assign sel_538349 = $signed({1'h0, add_538125, array_index_520967[0]}) < $signed({1'h0, sel_538127}) ? {add_538125, array_index_520967[0]} : sel_538127;
  assign add_538353 = sel_538286 + 16'h0001;
  assign add_538363 = array_index_518710[11:1] + 11'h5b9;
  assign sel_538365 = $signed({1'h0, add_538149, array_index_518210[0]}) < $signed({1'h0, sel_538151}) ? {add_538149, array_index_518210[0]} : sel_538151;
  assign add_538367 = array_index_518713[11:1] + 11'h5b9;
  assign sel_538369 = $signed({1'h0, add_538153, array_index_518213[0]}) < $signed({1'h0, sel_538155}) ? {add_538153, array_index_518213[0]} : sel_538155;
  assign add_538379 = array_index_519786[11:0] + 12'h37b;
  assign sel_538381 = $signed({1'h0, add_538165}) < $signed({1'h0, sel_538167}) ? add_538165 : sel_538167;
  assign add_538383 = array_index_519789[11:0] + 12'h37b;
  assign sel_538385 = $signed({1'h0, add_538169}) < $signed({1'h0, sel_538171}) ? add_538169 : sel_538171;
  assign add_538397 = array_index_520964[11:0] + 12'h811;
  assign sel_538399 = $signed({1'h0, add_538183}) < $signed({1'h0, sel_538185}) ? add_538183 : sel_538185;
  assign add_538401 = array_index_520967[11:0] + 12'h811;
  assign sel_538403 = $signed({1'h0, add_538187}) < $signed({1'h0, sel_538189}) ? add_538187 : sel_538189;
  assign sel_538416 = ($signed({1'h0, add_538053, array_index_521590[1:0]}) < $signed({1'h0, sel_538055}) ? {add_538053, array_index_521590[1:0]} : sel_538055) == ($signed({1'h0, add_538057, array_index_521593[1:0]}) < $signed({1'h0, sel_538059}) ? {add_538057, array_index_521593[1:0]} : sel_538059) ? add_538353 : sel_538286;
  assign add_538419 = array_index_518210[11:0] + 12'hcc1;
  assign sel_538421 = $signed({1'h0, add_538215}) < $signed({1'h0, sel_538217}) ? add_538215 : sel_538217;
  assign add_538423 = array_index_518213[11:0] + 12'hcc1;
  assign sel_538425 = $signed({1'h0, add_538219}) < $signed({1'h0, sel_538221}) ? add_538219 : sel_538221;
  assign add_538437 = array_index_519236[11:0] + 12'ha87;
  assign sel_538439 = $signed({1'h0, add_538233}) < $signed({1'h0, sel_538235}) ? add_538233 : sel_538235;
  assign add_538441 = array_index_519239[11:0] + 12'ha87;
  assign sel_538443 = $signed({1'h0, add_538237}) < $signed({1'h0, sel_538239}) ? add_538237 : sel_538239;
  assign add_538455 = array_index_520362[11:1] + 11'h663;
  assign sel_538457 = $signed({1'h0, add_538251, array_index_519786[0]}) < $signed({1'h0, sel_538253}) ? {add_538251, array_index_519786[0]} : sel_538253;
  assign add_538459 = array_index_520365[11:1] + 11'h663;
  assign sel_538461 = $signed({1'h0, add_538255, array_index_519789[0]}) < $signed({1'h0, sel_538257}) ? {add_538255, array_index_519789[0]} : sel_538257;
  assign add_538471 = array_index_521590[11:1] + 11'h075;
  assign sel_538473 = $signed({1'h0, add_538267, array_index_520964[0]}) < $signed({1'h0, sel_538269}) ? {add_538267, array_index_520964[0]} : sel_538269;
  assign add_538475 = array_index_521593[11:1] + 11'h075;
  assign sel_538477 = $signed({1'h0, add_538271, array_index_520967[0]}) < $signed({1'h0, sel_538273}) ? {add_538271, array_index_520967[0]} : sel_538273;
  assign add_538483 = sel_538416 + 16'h0001;
  assign add_538489 = array_index_518710[11:2] + 10'h113;
  assign sel_538491 = $signed({1'h0, add_538293, array_index_518210[1:0]}) < $signed({1'h0, sel_538295}) ? {add_538293, array_index_518210[1:0]} : sel_538295;
  assign add_538493 = array_index_518713[11:2] + 10'h113;
  assign sel_538495 = $signed({1'h0, add_538297, array_index_518213[1:0]}) < $signed({1'h0, sel_538299}) ? {add_538297, array_index_518213[1:0]} : sel_538299;
  assign add_538507 = array_index_519786[11:4] + 8'h49;
  assign sel_538509 = $signed({1'h0, add_538311, array_index_519236[3:0]}) < $signed({1'h0, sel_538313}) ? {add_538311, array_index_519236[3:0]} : sel_538313;
  assign add_538511 = array_index_519789[11:4] + 8'h49;
  assign sel_538513 = $signed({1'h0, add_538315, array_index_519239[3:0]}) < $signed({1'h0, sel_538317}) ? {add_538315, array_index_519239[3:0]} : sel_538317;
  assign add_538523 = array_index_520964[11:0] + 12'h263;
  assign sel_538525 = $signed({1'h0, add_538327}) < $signed({1'h0, sel_538329}) ? add_538327 : sel_538329;
  assign add_538527 = array_index_520967[11:0] + 12'h263;
  assign sel_538529 = $signed({1'h0, add_538331}) < $signed({1'h0, sel_538333}) ? add_538331 : sel_538333;
  assign sel_538540 = ($signed({1'h0, add_538201}) < $signed({1'h0, sel_538203}) ? add_538201 : sel_538203) == ($signed({1'h0, add_538205}) < $signed({1'h0, sel_538207}) ? add_538205 : sel_538207) ? add_538483 : sel_538416;
  assign add_538551 = array_index_519236[11:1] + 11'h5b9;
  assign sel_538553 = $signed({1'h0, add_538363, array_index_518710[0]}) < $signed({1'h0, sel_538365}) ? {add_538363, array_index_518710[0]} : sel_538365;
  assign add_538555 = array_index_519239[11:1] + 11'h5b9;
  assign sel_538557 = $signed({1'h0, add_538367, array_index_518713[0]}) < $signed({1'h0, sel_538369}) ? {add_538367, array_index_518713[0]} : sel_538369;
  assign add_538567 = array_index_520362[11:0] + 12'h37b;
  assign sel_538569 = $signed({1'h0, add_538379}) < $signed({1'h0, sel_538381}) ? add_538379 : sel_538381;
  assign add_538571 = array_index_520365[11:0] + 12'h37b;
  assign sel_538573 = $signed({1'h0, add_538383}) < $signed({1'h0, sel_538385}) ? add_538383 : sel_538385;
  assign add_538585 = array_index_521590[11:0] + 12'h811;
  assign sel_538587 = $signed({1'h0, add_538397}) < $signed({1'h0, sel_538399}) ? add_538397 : sel_538399;
  assign add_538589 = array_index_521593[11:0] + 12'h811;
  assign sel_538591 = $signed({1'h0, add_538401}) < $signed({1'h0, sel_538403}) ? add_538401 : sel_538403;
  assign add_538597 = sel_538540 + 16'h0001;
  assign add_538599 = array_index_518710[11:0] + 12'hcc1;
  assign sel_538601 = $signed({1'h0, add_538419}) < $signed({1'h0, sel_538421}) ? add_538419 : sel_538421;
  assign add_538603 = array_index_518713[11:0] + 12'hcc1;
  assign sel_538605 = $signed({1'h0, add_538423}) < $signed({1'h0, sel_538425}) ? add_538423 : sel_538425;
  assign add_538617 = array_index_519786[11:0] + 12'ha87;
  assign sel_538619 = $signed({1'h0, add_538437}) < $signed({1'h0, sel_538439}) ? add_538437 : sel_538439;
  assign add_538621 = array_index_519789[11:0] + 12'ha87;
  assign sel_538623 = $signed({1'h0, add_538441}) < $signed({1'h0, sel_538443}) ? add_538441 : sel_538443;
  assign add_538635 = array_index_520964[11:1] + 11'h663;
  assign sel_538637 = $signed({1'h0, add_538455, array_index_520362[0]}) < $signed({1'h0, sel_538457}) ? {add_538455, array_index_520362[0]} : sel_538457;
  assign add_538639 = array_index_520967[11:1] + 11'h663;
  assign sel_538641 = $signed({1'h0, add_538459, array_index_520365[0]}) < $signed({1'h0, sel_538461}) ? {add_538459, array_index_520365[0]} : sel_538461;
  assign sel_538652 = ($signed({1'h0, add_538343, array_index_521590[0]}) < $signed({1'h0, sel_538345}) ? {add_538343, array_index_521590[0]} : sel_538345) == ($signed({1'h0, add_538347, array_index_521593[0]}) < $signed({1'h0, sel_538349}) ? {add_538347, array_index_521593[0]} : sel_538349) ? add_538597 : sel_538540;
  assign add_538659 = array_index_519236[11:2] + 10'h113;
  assign sel_538661 = $signed({1'h0, add_538489, array_index_518710[1:0]}) < $signed({1'h0, sel_538491}) ? {add_538489, array_index_518710[1:0]} : sel_538491;
  assign add_538663 = array_index_519239[11:2] + 10'h113;
  assign sel_538665 = $signed({1'h0, add_538493, array_index_518713[1:0]}) < $signed({1'h0, sel_538495}) ? {add_538493, array_index_518713[1:0]} : sel_538495;
  assign add_538677 = array_index_520362[11:4] + 8'h49;
  assign sel_538679 = $signed({1'h0, add_538507, array_index_519786[3:0]}) < $signed({1'h0, sel_538509}) ? {add_538507, array_index_519786[3:0]} : sel_538509;
  assign add_538681 = array_index_520365[11:4] + 8'h49;
  assign sel_538683 = $signed({1'h0, add_538511, array_index_519789[3:0]}) < $signed({1'h0, sel_538513}) ? {add_538511, array_index_519789[3:0]} : sel_538513;
  assign add_538693 = array_index_521590[11:0] + 12'h263;
  assign sel_538695 = $signed({1'h0, add_538523}) < $signed({1'h0, sel_538525}) ? add_538523 : sel_538525;
  assign add_538697 = array_index_521593[11:0] + 12'h263;
  assign sel_538699 = $signed({1'h0, add_538527}) < $signed({1'h0, sel_538529}) ? add_538527 : sel_538529;
  assign add_538703 = sel_538652 + 16'h0001;
  assign add_538713 = array_index_519786[11:1] + 11'h5b9;
  assign sel_538715 = $signed({1'h0, add_538551, array_index_519236[0]}) < $signed({1'h0, sel_538553}) ? {add_538551, array_index_519236[0]} : sel_538553;
  assign add_538717 = array_index_519789[11:1] + 11'h5b9;
  assign sel_538719 = $signed({1'h0, add_538555, array_index_519239[0]}) < $signed({1'h0, sel_538557}) ? {add_538555, array_index_519239[0]} : sel_538557;
  assign add_538729 = array_index_520964[11:0] + 12'h37b;
  assign sel_538731 = $signed({1'h0, add_538567}) < $signed({1'h0, sel_538569}) ? add_538567 : sel_538569;
  assign add_538733 = array_index_520967[11:0] + 12'h37b;
  assign sel_538735 = $signed({1'h0, add_538571}) < $signed({1'h0, sel_538573}) ? add_538571 : sel_538573;
  assign sel_538748 = ($signed({1'h0, add_538471, array_index_521590[0]}) < $signed({1'h0, sel_538473}) ? {add_538471, array_index_521590[0]} : sel_538473) == ($signed({1'h0, add_538475, array_index_521593[0]}) < $signed({1'h0, sel_538477}) ? {add_538475, array_index_521593[0]} : sel_538477) ? add_538703 : sel_538652;
  assign add_538751 = array_index_519236[11:0] + 12'hcc1;
  assign sel_538753 = $signed({1'h0, add_538599}) < $signed({1'h0, sel_538601}) ? add_538599 : sel_538601;
  assign add_538755 = array_index_519239[11:0] + 12'hcc1;
  assign sel_538757 = $signed({1'h0, add_538603}) < $signed({1'h0, sel_538605}) ? add_538603 : sel_538605;
  assign add_538769 = array_index_520362[11:0] + 12'ha87;
  assign sel_538771 = $signed({1'h0, add_538617}) < $signed({1'h0, sel_538619}) ? add_538617 : sel_538619;
  assign add_538773 = array_index_520365[11:0] + 12'ha87;
  assign sel_538775 = $signed({1'h0, add_538621}) < $signed({1'h0, sel_538623}) ? add_538621 : sel_538623;
  assign add_538787 = array_index_521590[11:1] + 11'h663;
  assign sel_538789 = $signed({1'h0, add_538635, array_index_520964[0]}) < $signed({1'h0, sel_538637}) ? {add_538635, array_index_520964[0]} : sel_538637;
  assign add_538791 = array_index_521593[11:1] + 11'h663;
  assign sel_538793 = $signed({1'h0, add_538639, array_index_520967[0]}) < $signed({1'h0, sel_538641}) ? {add_538639, array_index_520967[0]} : sel_538641;
  assign add_538797 = sel_538748 + 16'h0001;
  assign add_538803 = array_index_519786[11:2] + 10'h113;
  assign sel_538805 = $signed({1'h0, add_538659, array_index_519236[1:0]}) < $signed({1'h0, sel_538661}) ? {add_538659, array_index_519236[1:0]} : sel_538661;
  assign add_538807 = array_index_519789[11:2] + 10'h113;
  assign sel_538809 = $signed({1'h0, add_538663, array_index_519239[1:0]}) < $signed({1'h0, sel_538665}) ? {add_538663, array_index_519239[1:0]} : sel_538665;
  assign add_538821 = array_index_520964[11:4] + 8'h49;
  assign sel_538823 = $signed({1'h0, add_538677, array_index_520362[3:0]}) < $signed({1'h0, sel_538679}) ? {add_538677, array_index_520362[3:0]} : sel_538679;
  assign add_538825 = array_index_520967[11:4] + 8'h49;
  assign sel_538827 = $signed({1'h0, add_538681, array_index_520365[3:0]}) < $signed({1'h0, sel_538683}) ? {add_538681, array_index_520365[3:0]} : sel_538683;
  assign sel_538838 = ($signed({1'h0, add_538585}) < $signed({1'h0, sel_538587}) ? add_538585 : sel_538587) == ($signed({1'h0, add_538589}) < $signed({1'h0, sel_538591}) ? add_538589 : sel_538591) ? add_538797 : sel_538748;
  assign add_538849 = array_index_520362[11:1] + 11'h5b9;
  assign sel_538851 = $signed({1'h0, add_538713, array_index_519786[0]}) < $signed({1'h0, sel_538715}) ? {add_538713, array_index_519786[0]} : sel_538715;
  assign add_538853 = array_index_520365[11:1] + 11'h5b9;
  assign sel_538855 = $signed({1'h0, add_538717, array_index_519789[0]}) < $signed({1'h0, sel_538719}) ? {add_538717, array_index_519789[0]} : sel_538719;
  assign add_538865 = array_index_521590[11:0] + 12'h37b;
  assign sel_538867 = $signed({1'h0, add_538729}) < $signed({1'h0, sel_538731}) ? add_538729 : sel_538731;
  assign add_538869 = array_index_521593[11:0] + 12'h37b;
  assign sel_538871 = $signed({1'h0, add_538733}) < $signed({1'h0, sel_538735}) ? add_538733 : sel_538735;
  assign add_538877 = sel_538838 + 16'h0001;
  assign add_538879 = array_index_519786[11:0] + 12'hcc1;
  assign sel_538881 = $signed({1'h0, add_538751}) < $signed({1'h0, sel_538753}) ? add_538751 : sel_538753;
  assign add_538883 = array_index_519789[11:0] + 12'hcc1;
  assign sel_538885 = $signed({1'h0, add_538755}) < $signed({1'h0, sel_538757}) ? add_538755 : sel_538757;
  assign add_538897 = array_index_520964[11:0] + 12'ha87;
  assign sel_538899 = $signed({1'h0, add_538769}) < $signed({1'h0, sel_538771}) ? add_538769 : sel_538771;
  assign add_538901 = array_index_520967[11:0] + 12'ha87;
  assign sel_538903 = $signed({1'h0, add_538773}) < $signed({1'h0, sel_538775}) ? add_538773 : sel_538775;
  assign sel_538916 = ($signed({1'h0, add_538693}) < $signed({1'h0, sel_538695}) ? add_538693 : sel_538695) == ($signed({1'h0, add_538697}) < $signed({1'h0, sel_538699}) ? add_538697 : sel_538699) ? add_538877 : sel_538838;
  assign add_538923 = array_index_520362[11:2] + 10'h113;
  assign sel_538925 = $signed({1'h0, add_538803, array_index_519786[1:0]}) < $signed({1'h0, sel_538805}) ? {add_538803, array_index_519786[1:0]} : sel_538805;
  assign add_538927 = array_index_520365[11:2] + 10'h113;
  assign sel_538929 = $signed({1'h0, add_538807, array_index_519789[1:0]}) < $signed({1'h0, sel_538809}) ? {add_538807, array_index_519789[1:0]} : sel_538809;
  assign add_538941 = array_index_521590[11:4] + 8'h49;
  assign sel_538943 = $signed({1'h0, add_538821, array_index_520964[3:0]}) < $signed({1'h0, sel_538823}) ? {add_538821, array_index_520964[3:0]} : sel_538823;
  assign add_538945 = array_index_521593[11:4] + 8'h49;
  assign sel_538947 = $signed({1'h0, add_538825, array_index_520967[3:0]}) < $signed({1'h0, sel_538827}) ? {add_538825, array_index_520967[3:0]} : sel_538827;
  assign add_538951 = sel_538916 + 16'h0001;
  assign add_538961 = array_index_520964[11:1] + 11'h5b9;
  assign sel_538963 = $signed({1'h0, add_538849, array_index_520362[0]}) < $signed({1'h0, sel_538851}) ? {add_538849, array_index_520362[0]} : sel_538851;
  assign add_538965 = array_index_520967[11:1] + 11'h5b9;
  assign sel_538967 = $signed({1'h0, add_538853, array_index_520365[0]}) < $signed({1'h0, sel_538855}) ? {add_538853, array_index_520365[0]} : sel_538855;
  assign sel_538978 = ($signed({1'h0, add_538787, array_index_521590[0]}) < $signed({1'h0, sel_538789}) ? {add_538787, array_index_521590[0]} : sel_538789) == ($signed({1'h0, add_538791, array_index_521593[0]}) < $signed({1'h0, sel_538793}) ? {add_538791, array_index_521593[0]} : sel_538793) ? add_538951 : sel_538916;
  assign add_538981 = array_index_520362[11:0] + 12'hcc1;
  assign sel_538983 = $signed({1'h0, add_538879}) < $signed({1'h0, sel_538881}) ? add_538879 : sel_538881;
  assign add_538985 = array_index_520365[11:0] + 12'hcc1;
  assign sel_538987 = $signed({1'h0, add_538883}) < $signed({1'h0, sel_538885}) ? add_538883 : sel_538885;
  assign add_538999 = array_index_521590[11:0] + 12'ha87;
  assign sel_539001 = $signed({1'h0, add_538897}) < $signed({1'h0, sel_538899}) ? add_538897 : sel_538899;
  assign add_539003 = array_index_521593[11:0] + 12'ha87;
  assign sel_539005 = $signed({1'h0, add_538901}) < $signed({1'h0, sel_538903}) ? add_538901 : sel_538903;
  assign add_539011 = sel_538978 + 16'h0001;
  assign add_539017 = array_index_520964[11:2] + 10'h113;
  assign sel_539019 = $signed({1'h0, add_538923, array_index_520362[1:0]}) < $signed({1'h0, sel_538925}) ? {add_538923, array_index_520362[1:0]} : sel_538925;
  assign add_539021 = array_index_520967[11:2] + 10'h113;
  assign sel_539023 = $signed({1'h0, add_538927, array_index_520365[1:0]}) < $signed({1'h0, sel_538929}) ? {add_538927, array_index_520365[1:0]} : sel_538929;
  assign sel_539036 = ($signed({1'h0, add_538865}) < $signed({1'h0, sel_538867}) ? add_538865 : sel_538867) == ($signed({1'h0, add_538869}) < $signed({1'h0, sel_538871}) ? add_538869 : sel_538871) ? add_539011 : sel_538978;
  assign add_539047 = array_index_521590[11:1] + 11'h5b9;
  assign sel_539049 = $signed({1'h0, add_538961, array_index_520964[0]}) < $signed({1'h0, sel_538963}) ? {add_538961, array_index_520964[0]} : sel_538963;
  assign add_539051 = array_index_521593[11:1] + 11'h5b9;
  assign sel_539053 = $signed({1'h0, add_538965, array_index_520967[0]}) < $signed({1'h0, sel_538967}) ? {add_538965, array_index_520967[0]} : sel_538967;
  assign add_539057 = sel_539036 + 16'h0001;
  assign add_539059 = array_index_520964[11:0] + 12'hcc1;
  assign sel_539061 = $signed({1'h0, add_538981}) < $signed({1'h0, sel_538983}) ? add_538981 : sel_538983;
  assign add_539063 = array_index_520967[11:0] + 12'hcc1;
  assign sel_539065 = $signed({1'h0, add_538985}) < $signed({1'h0, sel_538987}) ? add_538985 : sel_538987;
  assign sel_539078 = ($signed({1'h0, add_538941, array_index_521590[3:0]}) < $signed({1'h0, sel_538943}) ? {add_538941, array_index_521590[3:0]} : sel_538943) == ($signed({1'h0, add_538945, array_index_521593[3:0]}) < $signed({1'h0, sel_538947}) ? {add_538945, array_index_521593[3:0]} : sel_538947) ? add_539057 : sel_539036;
  assign add_539085 = array_index_521590[11:2] + 10'h113;
  assign sel_539087 = $signed({1'h0, add_539017, array_index_520964[1:0]}) < $signed({1'h0, sel_539019}) ? {add_539017, array_index_520964[1:0]} : sel_539019;
  assign add_539089 = array_index_521593[11:2] + 10'h113;
  assign sel_539091 = $signed({1'h0, add_539021, array_index_520967[1:0]}) < $signed({1'h0, sel_539023}) ? {add_539021, array_index_520967[1:0]} : sel_539023;
  assign add_539097 = sel_539078 + 16'h0001;
  assign sel_539108 = ($signed({1'h0, add_538999}) < $signed({1'h0, sel_539001}) ? add_538999 : sel_539001) == ($signed({1'h0, add_539003}) < $signed({1'h0, sel_539005}) ? add_539003 : sel_539005) ? add_539097 : sel_539078;
  assign add_539111 = array_index_521590[11:0] + 12'hcc1;
  assign sel_539113 = $signed({1'h0, add_539059}) < $signed({1'h0, sel_539061}) ? add_539059 : sel_539061;
  assign add_539115 = array_index_521593[11:0] + 12'hcc1;
  assign sel_539117 = $signed({1'h0, add_539063}) < $signed({1'h0, sel_539065}) ? add_539063 : sel_539065;
  assign add_539123 = sel_539108 + 16'h0001;
  assign sel_539130 = ($signed({1'h0, add_539047, array_index_521590[0]}) < $signed({1'h0, sel_539049}) ? {add_539047, array_index_521590[0]} : sel_539049) == ($signed({1'h0, add_539051, array_index_521593[0]}) < $signed({1'h0, sel_539053}) ? {add_539051, array_index_521593[0]} : sel_539053) ? add_539123 : sel_539108;
  assign add_539135 = sel_539130 + 16'h0001;
  assign sel_539138 = ($signed({1'h0, add_539085, array_index_521590[1:0]}) < $signed({1'h0, sel_539087}) ? {add_539085, array_index_521590[1:0]} : sel_539087) == ($signed({1'h0, add_539089, array_index_521593[1:0]}) < $signed({1'h0, sel_539091}) ? {add_539089, array_index_521593[1:0]} : sel_539091) ? add_539135 : sel_539130;
  assign add_539141 = sel_539138 + 16'h0001;
  assign out = {($signed({1'h0, add_539111}) < $signed({1'h0, sel_539113}) ? add_539111 : sel_539113) == ($signed({1'h0, add_539115}) < $signed({1'h0, sel_539117}) ? add_539115 : sel_539117) ? add_539141 : sel_539138, {set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
