module min_hash(
  input wire [319:0] set1,
  input wire [319:0] set2,
  output wire [655:0] out
);
  wire [15:0] set1_unflattened[20];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  wire [15:0] set2_unflattened[20];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  wire [15:0] array_index_35342;
  wire [15:0] array_index_35343;
  wire [11:0] add_35350;
  wire [11:0] add_35353;
  wire [15:0] array_index_35358;
  wire [15:0] array_index_35361;
  wire [10:0] add_35365;
  wire [10:0] add_35368;
  wire [11:0] add_35384;
  wire [11:0] sel_35386;
  wire [11:0] add_35389;
  wire [11:0] sel_35391;
  wire [15:0] array_index_35406;
  wire [15:0] array_index_35409;
  wire [8:0] add_35413;
  wire [8:0] add_35416;
  wire [10:0] add_35419;
  wire [11:0] sel_35422;
  wire [10:0] add_35424;
  wire [11:0] sel_35427;
  wire [11:0] add_35444;
  wire [11:0] sel_35446;
  wire [11:0] add_35449;
  wire [11:0] sel_35451;
  wire [15:0] array_index_35472;
  wire [15:0] array_index_35475;
  wire [10:0] add_35479;
  wire [10:0] add_35481;
  wire [8:0] add_35483;
  wire [11:0] sel_35486;
  wire [8:0] add_35488;
  wire [11:0] sel_35491;
  wire [10:0] add_35493;
  wire [11:0] sel_35496;
  wire [10:0] add_35498;
  wire [11:0] sel_35501;
  wire [11:0] add_35522;
  wire [11:0] sel_35524;
  wire [11:0] add_35527;
  wire [11:0] sel_35529;
  wire [15:0] array_index_35556;
  wire [15:0] array_index_35559;
  wire [10:0] add_35563;
  wire [10:0] add_35565;
  wire [10:0] add_35567;
  wire [11:0] sel_35569;
  wire [10:0] add_35571;
  wire [11:0] sel_35573;
  wire [8:0] add_35575;
  wire [11:0] sel_35578;
  wire [8:0] add_35580;
  wire [11:0] sel_35583;
  wire [10:0] add_35585;
  wire [11:0] sel_35588;
  wire [10:0] add_35590;
  wire [11:0] sel_35593;
  wire [11:0] add_35618;
  wire [11:0] sel_35620;
  wire [11:0] add_35623;
  wire [11:0] sel_35625;
  wire [15:0] array_index_35656;
  wire [15:0] array_index_35659;
  wire [10:0] add_35663;
  wire [11:0] sel_35665;
  wire [10:0] add_35667;
  wire [11:0] sel_35669;
  wire [10:0] add_35671;
  wire [11:0] sel_35673;
  wire [10:0] add_35675;
  wire [11:0] sel_35677;
  wire [8:0] add_35679;
  wire [11:0] sel_35682;
  wire [8:0] add_35684;
  wire [11:0] sel_35687;
  wire [10:0] add_35689;
  wire [11:0] sel_35692;
  wire [10:0] add_35694;
  wire [11:0] sel_35697;
  wire [11:0] add_35722;
  wire [11:0] sel_35724;
  wire [11:0] add_35727;
  wire [11:0] sel_35729;
  wire [15:0] array_index_35758;
  wire [15:0] array_index_35761;
  wire [10:0] add_35765;
  wire [11:0] sel_35767;
  wire [10:0] add_35769;
  wire [11:0] sel_35771;
  wire [10:0] add_35773;
  wire [11:0] sel_35775;
  wire [10:0] add_35777;
  wire [11:0] sel_35779;
  wire [8:0] add_35781;
  wire [11:0] sel_35784;
  wire [8:0] add_35786;
  wire [11:0] sel_35789;
  wire [10:0] add_35791;
  wire [11:0] sel_35794;
  wire [10:0] add_35796;
  wire [11:0] sel_35799;
  wire [11:0] add_35824;
  wire [11:0] sel_35826;
  wire [11:0] add_35829;
  wire [11:0] sel_35831;
  wire [15:0] array_index_35860;
  wire [15:0] array_index_35863;
  wire [10:0] add_35867;
  wire [11:0] sel_35869;
  wire [10:0] add_35871;
  wire [11:0] sel_35873;
  wire [10:0] add_35875;
  wire [11:0] sel_35877;
  wire [10:0] add_35879;
  wire [11:0] sel_35881;
  wire [8:0] add_35883;
  wire [11:0] sel_35886;
  wire [8:0] add_35888;
  wire [11:0] sel_35891;
  wire [10:0] add_35893;
  wire [11:0] sel_35896;
  wire [10:0] add_35898;
  wire [11:0] sel_35901;
  wire [11:0] add_35926;
  wire [11:0] sel_35928;
  wire [11:0] add_35931;
  wire [11:0] sel_35933;
  wire [15:0] array_index_35962;
  wire [15:0] array_index_35965;
  wire [10:0] add_35969;
  wire [11:0] sel_35971;
  wire [10:0] add_35973;
  wire [11:0] sel_35975;
  wire [10:0] add_35977;
  wire [11:0] sel_35979;
  wire [10:0] add_35981;
  wire [11:0] sel_35983;
  wire [8:0] add_35985;
  wire [11:0] sel_35988;
  wire [8:0] add_35990;
  wire [11:0] sel_35993;
  wire [10:0] add_35995;
  wire [11:0] sel_35998;
  wire [10:0] add_36000;
  wire [11:0] sel_36003;
  wire [11:0] add_36028;
  wire [11:0] sel_36030;
  wire [11:0] add_36033;
  wire [11:0] sel_36035;
  wire [15:0] array_index_36064;
  wire [15:0] array_index_36067;
  wire [10:0] add_36071;
  wire [11:0] sel_36073;
  wire [10:0] add_36075;
  wire [11:0] sel_36077;
  wire [10:0] add_36079;
  wire [11:0] sel_36081;
  wire [10:0] add_36083;
  wire [11:0] sel_36085;
  wire [8:0] add_36087;
  wire [11:0] sel_36090;
  wire [8:0] add_36092;
  wire [11:0] sel_36095;
  wire [10:0] add_36097;
  wire [11:0] sel_36100;
  wire [10:0] add_36102;
  wire [11:0] sel_36105;
  wire [11:0] add_36130;
  wire [11:0] sel_36132;
  wire [11:0] add_36135;
  wire [11:0] sel_36137;
  wire [15:0] array_index_36166;
  wire [15:0] array_index_36169;
  wire [10:0] add_36173;
  wire [11:0] sel_36175;
  wire [10:0] add_36177;
  wire [11:0] sel_36179;
  wire [10:0] add_36181;
  wire [11:0] sel_36183;
  wire [10:0] add_36185;
  wire [11:0] sel_36187;
  wire [8:0] add_36189;
  wire [11:0] sel_36192;
  wire [8:0] add_36194;
  wire [11:0] sel_36197;
  wire [10:0] add_36199;
  wire [11:0] sel_36202;
  wire [10:0] add_36204;
  wire [11:0] sel_36207;
  wire [11:0] add_36232;
  wire [11:0] sel_36234;
  wire [11:0] add_36237;
  wire [11:0] sel_36239;
  wire [15:0] array_index_36268;
  wire [15:0] array_index_36271;
  wire [10:0] add_36275;
  wire [11:0] sel_36277;
  wire [10:0] add_36279;
  wire [11:0] sel_36281;
  wire [10:0] add_36283;
  wire [11:0] sel_36285;
  wire [10:0] add_36287;
  wire [11:0] sel_36289;
  wire [8:0] add_36291;
  wire [11:0] sel_36294;
  wire [8:0] add_36296;
  wire [11:0] sel_36299;
  wire [10:0] add_36301;
  wire [11:0] sel_36304;
  wire [10:0] add_36306;
  wire [11:0] sel_36309;
  wire [11:0] add_36334;
  wire [11:0] sel_36336;
  wire [11:0] add_36339;
  wire [11:0] sel_36341;
  wire [15:0] array_index_36370;
  wire [15:0] array_index_36373;
  wire [10:0] add_36377;
  wire [11:0] sel_36379;
  wire [10:0] add_36381;
  wire [11:0] sel_36383;
  wire [10:0] add_36385;
  wire [11:0] sel_36387;
  wire [10:0] add_36389;
  wire [11:0] sel_36391;
  wire [8:0] add_36393;
  wire [11:0] sel_36396;
  wire [8:0] add_36398;
  wire [11:0] sel_36401;
  wire [10:0] add_36403;
  wire [11:0] sel_36406;
  wire [10:0] add_36408;
  wire [11:0] sel_36411;
  wire [11:0] add_36436;
  wire [11:0] sel_36438;
  wire [11:0] add_36441;
  wire [11:0] sel_36443;
  wire [15:0] array_index_36472;
  wire [15:0] array_index_36475;
  wire [10:0] add_36479;
  wire [11:0] sel_36481;
  wire [10:0] add_36483;
  wire [11:0] sel_36485;
  wire [10:0] add_36487;
  wire [11:0] sel_36489;
  wire [10:0] add_36491;
  wire [11:0] sel_36493;
  wire [8:0] add_36495;
  wire [11:0] sel_36498;
  wire [8:0] add_36500;
  wire [11:0] sel_36503;
  wire [10:0] add_36505;
  wire [11:0] sel_36508;
  wire [10:0] add_36510;
  wire [11:0] sel_36513;
  wire [11:0] add_36538;
  wire [11:0] sel_36540;
  wire [11:0] add_36543;
  wire [11:0] sel_36545;
  wire [15:0] array_index_36574;
  wire [15:0] array_index_36577;
  wire [10:0] add_36581;
  wire [11:0] sel_36583;
  wire [10:0] add_36585;
  wire [11:0] sel_36587;
  wire [10:0] add_36589;
  wire [11:0] sel_36591;
  wire [10:0] add_36593;
  wire [11:0] sel_36595;
  wire [8:0] add_36597;
  wire [11:0] sel_36600;
  wire [8:0] add_36602;
  wire [11:0] sel_36605;
  wire [10:0] add_36607;
  wire [11:0] sel_36610;
  wire [10:0] add_36612;
  wire [11:0] sel_36615;
  wire [11:0] add_36640;
  wire [11:0] sel_36642;
  wire [11:0] add_36645;
  wire [11:0] sel_36647;
  wire [15:0] array_index_36676;
  wire [15:0] array_index_36679;
  wire [10:0] add_36683;
  wire [11:0] sel_36685;
  wire [10:0] add_36687;
  wire [11:0] sel_36689;
  wire [10:0] add_36691;
  wire [11:0] sel_36693;
  wire [10:0] add_36695;
  wire [11:0] sel_36697;
  wire [8:0] add_36699;
  wire [11:0] sel_36702;
  wire [8:0] add_36704;
  wire [11:0] sel_36707;
  wire [10:0] add_36709;
  wire [11:0] sel_36712;
  wire [10:0] add_36714;
  wire [11:0] sel_36717;
  wire [11:0] add_36742;
  wire [11:0] sel_36744;
  wire [11:0] add_36747;
  wire [11:0] sel_36749;
  wire [15:0] array_index_36778;
  wire [15:0] array_index_36781;
  wire [10:0] add_36785;
  wire [11:0] sel_36787;
  wire [10:0] add_36789;
  wire [11:0] sel_36791;
  wire [10:0] add_36793;
  wire [11:0] sel_36795;
  wire [10:0] add_36797;
  wire [11:0] sel_36799;
  wire [8:0] add_36801;
  wire [11:0] sel_36804;
  wire [8:0] add_36806;
  wire [11:0] sel_36809;
  wire [10:0] add_36811;
  wire [11:0] sel_36814;
  wire [10:0] add_36816;
  wire [11:0] sel_36819;
  wire [11:0] add_36844;
  wire [11:0] sel_36846;
  wire [11:0] add_36849;
  wire [11:0] sel_36851;
  wire [15:0] array_index_36880;
  wire [15:0] array_index_36883;
  wire [10:0] add_36887;
  wire [11:0] sel_36889;
  wire [10:0] add_36891;
  wire [11:0] sel_36893;
  wire [10:0] add_36895;
  wire [11:0] sel_36897;
  wire [10:0] add_36899;
  wire [11:0] sel_36901;
  wire [8:0] add_36903;
  wire [11:0] sel_36906;
  wire [8:0] add_36908;
  wire [11:0] sel_36911;
  wire [10:0] add_36913;
  wire [11:0] sel_36916;
  wire [10:0] add_36918;
  wire [11:0] sel_36921;
  wire [11:0] add_36946;
  wire [11:0] sel_36948;
  wire [11:0] add_36951;
  wire [11:0] sel_36953;
  wire [15:0] array_index_36982;
  wire [15:0] array_index_36985;
  wire [10:0] add_36989;
  wire [11:0] sel_36991;
  wire [10:0] add_36993;
  wire [11:0] sel_36995;
  wire [10:0] add_36997;
  wire [11:0] sel_36999;
  wire [10:0] add_37001;
  wire [11:0] sel_37003;
  wire [8:0] add_37005;
  wire [11:0] sel_37008;
  wire [8:0] add_37010;
  wire [11:0] sel_37013;
  wire [10:0] add_37015;
  wire [11:0] sel_37018;
  wire [10:0] add_37020;
  wire [11:0] sel_37023;
  wire [11:0] add_37048;
  wire [11:0] sel_37050;
  wire [11:0] add_37053;
  wire [11:0] sel_37055;
  wire [15:0] array_index_37084;
  wire [15:0] array_index_37087;
  wire [10:0] add_37091;
  wire [11:0] sel_37093;
  wire [10:0] add_37095;
  wire [11:0] sel_37097;
  wire [10:0] add_37099;
  wire [11:0] sel_37101;
  wire [10:0] add_37103;
  wire [11:0] sel_37105;
  wire [8:0] add_37107;
  wire [11:0] sel_37110;
  wire [8:0] add_37112;
  wire [11:0] sel_37115;
  wire [10:0] add_37117;
  wire [11:0] sel_37120;
  wire [10:0] add_37122;
  wire [11:0] sel_37125;
  wire [11:0] add_37149;
  wire [11:0] sel_37151;
  wire [11:0] add_37153;
  wire [11:0] sel_37155;
  wire [10:0] add_37189;
  wire [11:0] sel_37191;
  wire [10:0] add_37193;
  wire [11:0] sel_37195;
  wire [10:0] add_37197;
  wire [11:0] sel_37199;
  wire [10:0] add_37201;
  wire [11:0] sel_37203;
  wire [8:0] add_37205;
  wire [11:0] sel_37208;
  wire [8:0] add_37210;
  wire [11:0] sel_37213;
  wire [10:0] add_37215;
  wire [11:0] sel_37218;
  wire [10:0] add_37220;
  wire [11:0] sel_37223;
  wire [10:0] add_37271;
  wire [11:0] sel_37273;
  wire [10:0] add_37275;
  wire [11:0] sel_37277;
  wire [10:0] add_37279;
  wire [11:0] sel_37281;
  wire [10:0] add_37283;
  wire [11:0] sel_37285;
  wire [8:0] add_37287;
  wire [11:0] sel_37290;
  wire [8:0] add_37292;
  wire [11:0] sel_37295;
  wire [1:0] concat_37298;
  wire [1:0] add_37313;
  wire [10:0] add_37333;
  wire [11:0] sel_37335;
  wire [10:0] add_37337;
  wire [11:0] sel_37339;
  wire [10:0] add_37341;
  wire [11:0] sel_37343;
  wire [10:0] add_37345;
  wire [11:0] sel_37347;
  wire [2:0] concat_37350;
  wire [2:0] add_37361;
  wire [10:0] add_37375;
  wire [11:0] sel_37377;
  wire [10:0] add_37379;
  wire [11:0] sel_37381;
  wire [3:0] concat_37384;
  wire [3:0] add_37391;
  wire [4:0] concat_37400;
  wire [4:0] add_37403;
  assign array_index_35342 = set1_unflattened[5'h00];
  assign array_index_35343 = set2_unflattened[5'h00];
  assign add_35350 = array_index_35342[11:0] + 12'h247;
  assign add_35353 = array_index_35343[11:0] + 12'h247;
  assign array_index_35358 = set1_unflattened[5'h01];
  assign array_index_35361 = set2_unflattened[5'h01];
  assign add_35365 = array_index_35342[11:1] + 11'h247;
  assign add_35368 = array_index_35343[11:1] + 11'h247;
  assign add_35384 = array_index_35358[11:0] + 12'h247;
  assign sel_35386 = $signed({1'h0, add_35350}) < $signed(13'h0fff) ? add_35350 : 12'hfff;
  assign add_35389 = array_index_35361[11:0] + 12'h247;
  assign sel_35391 = $signed({1'h0, add_35353}) < $signed(13'h0fff) ? add_35353 : 12'hfff;
  assign array_index_35406 = set1_unflattened[5'h02];
  assign array_index_35409 = set2_unflattened[5'h02];
  assign add_35413 = array_index_35342[11:3] + 9'h0bd;
  assign add_35416 = array_index_35343[11:3] + 9'h0bd;
  assign add_35419 = array_index_35358[11:1] + 11'h247;
  assign sel_35422 = $signed({1'h0, add_35365, array_index_35342[0]}) < $signed(13'h0fff) ? {add_35365, array_index_35342[0]} : 12'hfff;
  assign add_35424 = array_index_35361[11:1] + 11'h247;
  assign sel_35427 = $signed({1'h0, add_35368, array_index_35343[0]}) < $signed(13'h0fff) ? {add_35368, array_index_35343[0]} : 12'hfff;
  assign add_35444 = array_index_35406[11:0] + 12'h247;
  assign sel_35446 = $signed({1'h0, add_35384}) < $signed({1'h0, sel_35386}) ? add_35384 : sel_35386;
  assign add_35449 = array_index_35409[11:0] + 12'h247;
  assign sel_35451 = $signed({1'h0, add_35389}) < $signed({1'h0, sel_35391}) ? add_35389 : sel_35391;
  assign array_index_35472 = set1_unflattened[5'h03];
  assign array_index_35475 = set2_unflattened[5'h03];
  assign add_35479 = array_index_35342[11:1] + 11'h347;
  assign add_35481 = array_index_35343[11:1] + 11'h347;
  assign add_35483 = array_index_35358[11:3] + 9'h0bd;
  assign sel_35486 = $signed({1'h0, add_35413, array_index_35342[2:0]}) < $signed(13'h0fff) ? {add_35413, array_index_35342[2:0]} : 12'hfff;
  assign add_35488 = array_index_35361[11:3] + 9'h0bd;
  assign sel_35491 = $signed({1'h0, add_35416, array_index_35343[2:0]}) < $signed(13'h0fff) ? {add_35416, array_index_35343[2:0]} : 12'hfff;
  assign add_35493 = array_index_35406[11:1] + 11'h247;
  assign sel_35496 = $signed({1'h0, add_35419, array_index_35358[0]}) < $signed({1'h0, sel_35422}) ? {add_35419, array_index_35358[0]} : sel_35422;
  assign add_35498 = array_index_35409[11:1] + 11'h247;
  assign sel_35501 = $signed({1'h0, add_35424, array_index_35361[0]}) < $signed({1'h0, sel_35427}) ? {add_35424, array_index_35361[0]} : sel_35427;
  assign add_35522 = array_index_35472[11:0] + 12'h247;
  assign sel_35524 = $signed({1'h0, add_35444}) < $signed({1'h0, sel_35446}) ? add_35444 : sel_35446;
  assign add_35527 = array_index_35475[11:0] + 12'h247;
  assign sel_35529 = $signed({1'h0, add_35449}) < $signed({1'h0, sel_35451}) ? add_35449 : sel_35451;
  assign array_index_35556 = set1_unflattened[5'h04];
  assign array_index_35559 = set2_unflattened[5'h04];
  assign add_35563 = array_index_35342[11:1] + 11'h79d;
  assign add_35565 = array_index_35343[11:1] + 11'h79d;
  assign add_35567 = array_index_35358[11:1] + 11'h347;
  assign sel_35569 = $signed({1'h0, add_35479, array_index_35342[0]}) < $signed(13'h0fff) ? {add_35479, array_index_35342[0]} : 12'hfff;
  assign add_35571 = array_index_35361[11:1] + 11'h347;
  assign sel_35573 = $signed({1'h0, add_35481, array_index_35343[0]}) < $signed(13'h0fff) ? {add_35481, array_index_35343[0]} : 12'hfff;
  assign add_35575 = array_index_35406[11:3] + 9'h0bd;
  assign sel_35578 = $signed({1'h0, add_35483, array_index_35358[2:0]}) < $signed({1'h0, sel_35486}) ? {add_35483, array_index_35358[2:0]} : sel_35486;
  assign add_35580 = array_index_35409[11:3] + 9'h0bd;
  assign sel_35583 = $signed({1'h0, add_35488, array_index_35361[2:0]}) < $signed({1'h0, sel_35491}) ? {add_35488, array_index_35361[2:0]} : sel_35491;
  assign add_35585 = array_index_35472[11:1] + 11'h247;
  assign sel_35588 = $signed({1'h0, add_35493, array_index_35406[0]}) < $signed({1'h0, sel_35496}) ? {add_35493, array_index_35406[0]} : sel_35496;
  assign add_35590 = array_index_35475[11:1] + 11'h247;
  assign sel_35593 = $signed({1'h0, add_35498, array_index_35409[0]}) < $signed({1'h0, sel_35501}) ? {add_35498, array_index_35409[0]} : sel_35501;
  assign add_35618 = array_index_35556[11:0] + 12'h247;
  assign sel_35620 = $signed({1'h0, add_35522}) < $signed({1'h0, sel_35524}) ? add_35522 : sel_35524;
  assign add_35623 = array_index_35559[11:0] + 12'h247;
  assign sel_35625 = $signed({1'h0, add_35527}) < $signed({1'h0, sel_35529}) ? add_35527 : sel_35529;
  assign array_index_35656 = set1_unflattened[5'h05];
  assign array_index_35659 = set2_unflattened[5'h05];
  assign add_35663 = array_index_35358[11:1] + 11'h79d;
  assign sel_35665 = $signed({1'h0, add_35563, array_index_35342[0]}) < $signed(13'h0fff) ? {add_35563, array_index_35342[0]} : 12'hfff;
  assign add_35667 = array_index_35361[11:1] + 11'h79d;
  assign sel_35669 = $signed({1'h0, add_35565, array_index_35343[0]}) < $signed(13'h0fff) ? {add_35565, array_index_35343[0]} : 12'hfff;
  assign add_35671 = array_index_35406[11:1] + 11'h347;
  assign sel_35673 = $signed({1'h0, add_35567, array_index_35358[0]}) < $signed({1'h0, sel_35569}) ? {add_35567, array_index_35358[0]} : sel_35569;
  assign add_35675 = array_index_35409[11:1] + 11'h347;
  assign sel_35677 = $signed({1'h0, add_35571, array_index_35361[0]}) < $signed({1'h0, sel_35573}) ? {add_35571, array_index_35361[0]} : sel_35573;
  assign add_35679 = array_index_35472[11:3] + 9'h0bd;
  assign sel_35682 = $signed({1'h0, add_35575, array_index_35406[2:0]}) < $signed({1'h0, sel_35578}) ? {add_35575, array_index_35406[2:0]} : sel_35578;
  assign add_35684 = array_index_35475[11:3] + 9'h0bd;
  assign sel_35687 = $signed({1'h0, add_35580, array_index_35409[2:0]}) < $signed({1'h0, sel_35583}) ? {add_35580, array_index_35409[2:0]} : sel_35583;
  assign add_35689 = array_index_35556[11:1] + 11'h247;
  assign sel_35692 = $signed({1'h0, add_35585, array_index_35472[0]}) < $signed({1'h0, sel_35588}) ? {add_35585, array_index_35472[0]} : sel_35588;
  assign add_35694 = array_index_35559[11:1] + 11'h247;
  assign sel_35697 = $signed({1'h0, add_35590, array_index_35475[0]}) < $signed({1'h0, sel_35593}) ? {add_35590, array_index_35475[0]} : sel_35593;
  assign add_35722 = array_index_35656[11:0] + 12'h247;
  assign sel_35724 = $signed({1'h0, add_35618}) < $signed({1'h0, sel_35620}) ? add_35618 : sel_35620;
  assign add_35727 = array_index_35659[11:0] + 12'h247;
  assign sel_35729 = $signed({1'h0, add_35623}) < $signed({1'h0, sel_35625}) ? add_35623 : sel_35625;
  assign array_index_35758 = set1_unflattened[5'h06];
  assign array_index_35761 = set2_unflattened[5'h06];
  assign add_35765 = array_index_35406[11:1] + 11'h79d;
  assign sel_35767 = $signed({1'h0, add_35663, array_index_35358[0]}) < $signed({1'h0, sel_35665}) ? {add_35663, array_index_35358[0]} : sel_35665;
  assign add_35769 = array_index_35409[11:1] + 11'h79d;
  assign sel_35771 = $signed({1'h0, add_35667, array_index_35361[0]}) < $signed({1'h0, sel_35669}) ? {add_35667, array_index_35361[0]} : sel_35669;
  assign add_35773 = array_index_35472[11:1] + 11'h347;
  assign sel_35775 = $signed({1'h0, add_35671, array_index_35406[0]}) < $signed({1'h0, sel_35673}) ? {add_35671, array_index_35406[0]} : sel_35673;
  assign add_35777 = array_index_35475[11:1] + 11'h347;
  assign sel_35779 = $signed({1'h0, add_35675, array_index_35409[0]}) < $signed({1'h0, sel_35677}) ? {add_35675, array_index_35409[0]} : sel_35677;
  assign add_35781 = array_index_35556[11:3] + 9'h0bd;
  assign sel_35784 = $signed({1'h0, add_35679, array_index_35472[2:0]}) < $signed({1'h0, sel_35682}) ? {add_35679, array_index_35472[2:0]} : sel_35682;
  assign add_35786 = array_index_35559[11:3] + 9'h0bd;
  assign sel_35789 = $signed({1'h0, add_35684, array_index_35475[2:0]}) < $signed({1'h0, sel_35687}) ? {add_35684, array_index_35475[2:0]} : sel_35687;
  assign add_35791 = array_index_35656[11:1] + 11'h247;
  assign sel_35794 = $signed({1'h0, add_35689, array_index_35556[0]}) < $signed({1'h0, sel_35692}) ? {add_35689, array_index_35556[0]} : sel_35692;
  assign add_35796 = array_index_35659[11:1] + 11'h247;
  assign sel_35799 = $signed({1'h0, add_35694, array_index_35559[0]}) < $signed({1'h0, sel_35697}) ? {add_35694, array_index_35559[0]} : sel_35697;
  assign add_35824 = array_index_35758[11:0] + 12'h247;
  assign sel_35826 = $signed({1'h0, add_35722}) < $signed({1'h0, sel_35724}) ? add_35722 : sel_35724;
  assign add_35829 = array_index_35761[11:0] + 12'h247;
  assign sel_35831 = $signed({1'h0, add_35727}) < $signed({1'h0, sel_35729}) ? add_35727 : sel_35729;
  assign array_index_35860 = set1_unflattened[5'h07];
  assign array_index_35863 = set2_unflattened[5'h07];
  assign add_35867 = array_index_35472[11:1] + 11'h79d;
  assign sel_35869 = $signed({1'h0, add_35765, array_index_35406[0]}) < $signed({1'h0, sel_35767}) ? {add_35765, array_index_35406[0]} : sel_35767;
  assign add_35871 = array_index_35475[11:1] + 11'h79d;
  assign sel_35873 = $signed({1'h0, add_35769, array_index_35409[0]}) < $signed({1'h0, sel_35771}) ? {add_35769, array_index_35409[0]} : sel_35771;
  assign add_35875 = array_index_35556[11:1] + 11'h347;
  assign sel_35877 = $signed({1'h0, add_35773, array_index_35472[0]}) < $signed({1'h0, sel_35775}) ? {add_35773, array_index_35472[0]} : sel_35775;
  assign add_35879 = array_index_35559[11:1] + 11'h347;
  assign sel_35881 = $signed({1'h0, add_35777, array_index_35475[0]}) < $signed({1'h0, sel_35779}) ? {add_35777, array_index_35475[0]} : sel_35779;
  assign add_35883 = array_index_35656[11:3] + 9'h0bd;
  assign sel_35886 = $signed({1'h0, add_35781, array_index_35556[2:0]}) < $signed({1'h0, sel_35784}) ? {add_35781, array_index_35556[2:0]} : sel_35784;
  assign add_35888 = array_index_35659[11:3] + 9'h0bd;
  assign sel_35891 = $signed({1'h0, add_35786, array_index_35559[2:0]}) < $signed({1'h0, sel_35789}) ? {add_35786, array_index_35559[2:0]} : sel_35789;
  assign add_35893 = array_index_35758[11:1] + 11'h247;
  assign sel_35896 = $signed({1'h0, add_35791, array_index_35656[0]}) < $signed({1'h0, sel_35794}) ? {add_35791, array_index_35656[0]} : sel_35794;
  assign add_35898 = array_index_35761[11:1] + 11'h247;
  assign sel_35901 = $signed({1'h0, add_35796, array_index_35659[0]}) < $signed({1'h0, sel_35799}) ? {add_35796, array_index_35659[0]} : sel_35799;
  assign add_35926 = array_index_35860[11:0] + 12'h247;
  assign sel_35928 = $signed({1'h0, add_35824}) < $signed({1'h0, sel_35826}) ? add_35824 : sel_35826;
  assign add_35931 = array_index_35863[11:0] + 12'h247;
  assign sel_35933 = $signed({1'h0, add_35829}) < $signed({1'h0, sel_35831}) ? add_35829 : sel_35831;
  assign array_index_35962 = set1_unflattened[5'h08];
  assign array_index_35965 = set2_unflattened[5'h08];
  assign add_35969 = array_index_35556[11:1] + 11'h79d;
  assign sel_35971 = $signed({1'h0, add_35867, array_index_35472[0]}) < $signed({1'h0, sel_35869}) ? {add_35867, array_index_35472[0]} : sel_35869;
  assign add_35973 = array_index_35559[11:1] + 11'h79d;
  assign sel_35975 = $signed({1'h0, add_35871, array_index_35475[0]}) < $signed({1'h0, sel_35873}) ? {add_35871, array_index_35475[0]} : sel_35873;
  assign add_35977 = array_index_35656[11:1] + 11'h347;
  assign sel_35979 = $signed({1'h0, add_35875, array_index_35556[0]}) < $signed({1'h0, sel_35877}) ? {add_35875, array_index_35556[0]} : sel_35877;
  assign add_35981 = array_index_35659[11:1] + 11'h347;
  assign sel_35983 = $signed({1'h0, add_35879, array_index_35559[0]}) < $signed({1'h0, sel_35881}) ? {add_35879, array_index_35559[0]} : sel_35881;
  assign add_35985 = array_index_35758[11:3] + 9'h0bd;
  assign sel_35988 = $signed({1'h0, add_35883, array_index_35656[2:0]}) < $signed({1'h0, sel_35886}) ? {add_35883, array_index_35656[2:0]} : sel_35886;
  assign add_35990 = array_index_35761[11:3] + 9'h0bd;
  assign sel_35993 = $signed({1'h0, add_35888, array_index_35659[2:0]}) < $signed({1'h0, sel_35891}) ? {add_35888, array_index_35659[2:0]} : sel_35891;
  assign add_35995 = array_index_35860[11:1] + 11'h247;
  assign sel_35998 = $signed({1'h0, add_35893, array_index_35758[0]}) < $signed({1'h0, sel_35896}) ? {add_35893, array_index_35758[0]} : sel_35896;
  assign add_36000 = array_index_35863[11:1] + 11'h247;
  assign sel_36003 = $signed({1'h0, add_35898, array_index_35761[0]}) < $signed({1'h0, sel_35901}) ? {add_35898, array_index_35761[0]} : sel_35901;
  assign add_36028 = array_index_35962[11:0] + 12'h247;
  assign sel_36030 = $signed({1'h0, add_35926}) < $signed({1'h0, sel_35928}) ? add_35926 : sel_35928;
  assign add_36033 = array_index_35965[11:0] + 12'h247;
  assign sel_36035 = $signed({1'h0, add_35931}) < $signed({1'h0, sel_35933}) ? add_35931 : sel_35933;
  assign array_index_36064 = set1_unflattened[5'h09];
  assign array_index_36067 = set2_unflattened[5'h09];
  assign add_36071 = array_index_35656[11:1] + 11'h79d;
  assign sel_36073 = $signed({1'h0, add_35969, array_index_35556[0]}) < $signed({1'h0, sel_35971}) ? {add_35969, array_index_35556[0]} : sel_35971;
  assign add_36075 = array_index_35659[11:1] + 11'h79d;
  assign sel_36077 = $signed({1'h0, add_35973, array_index_35559[0]}) < $signed({1'h0, sel_35975}) ? {add_35973, array_index_35559[0]} : sel_35975;
  assign add_36079 = array_index_35758[11:1] + 11'h347;
  assign sel_36081 = $signed({1'h0, add_35977, array_index_35656[0]}) < $signed({1'h0, sel_35979}) ? {add_35977, array_index_35656[0]} : sel_35979;
  assign add_36083 = array_index_35761[11:1] + 11'h347;
  assign sel_36085 = $signed({1'h0, add_35981, array_index_35659[0]}) < $signed({1'h0, sel_35983}) ? {add_35981, array_index_35659[0]} : sel_35983;
  assign add_36087 = array_index_35860[11:3] + 9'h0bd;
  assign sel_36090 = $signed({1'h0, add_35985, array_index_35758[2:0]}) < $signed({1'h0, sel_35988}) ? {add_35985, array_index_35758[2:0]} : sel_35988;
  assign add_36092 = array_index_35863[11:3] + 9'h0bd;
  assign sel_36095 = $signed({1'h0, add_35990, array_index_35761[2:0]}) < $signed({1'h0, sel_35993}) ? {add_35990, array_index_35761[2:0]} : sel_35993;
  assign add_36097 = array_index_35962[11:1] + 11'h247;
  assign sel_36100 = $signed({1'h0, add_35995, array_index_35860[0]}) < $signed({1'h0, sel_35998}) ? {add_35995, array_index_35860[0]} : sel_35998;
  assign add_36102 = array_index_35965[11:1] + 11'h247;
  assign sel_36105 = $signed({1'h0, add_36000, array_index_35863[0]}) < $signed({1'h0, sel_36003}) ? {add_36000, array_index_35863[0]} : sel_36003;
  assign add_36130 = array_index_36064[11:0] + 12'h247;
  assign sel_36132 = $signed({1'h0, add_36028}) < $signed({1'h0, sel_36030}) ? add_36028 : sel_36030;
  assign add_36135 = array_index_36067[11:0] + 12'h247;
  assign sel_36137 = $signed({1'h0, add_36033}) < $signed({1'h0, sel_36035}) ? add_36033 : sel_36035;
  assign array_index_36166 = set1_unflattened[5'h0a];
  assign array_index_36169 = set2_unflattened[5'h0a];
  assign add_36173 = array_index_35758[11:1] + 11'h79d;
  assign sel_36175 = $signed({1'h0, add_36071, array_index_35656[0]}) < $signed({1'h0, sel_36073}) ? {add_36071, array_index_35656[0]} : sel_36073;
  assign add_36177 = array_index_35761[11:1] + 11'h79d;
  assign sel_36179 = $signed({1'h0, add_36075, array_index_35659[0]}) < $signed({1'h0, sel_36077}) ? {add_36075, array_index_35659[0]} : sel_36077;
  assign add_36181 = array_index_35860[11:1] + 11'h347;
  assign sel_36183 = $signed({1'h0, add_36079, array_index_35758[0]}) < $signed({1'h0, sel_36081}) ? {add_36079, array_index_35758[0]} : sel_36081;
  assign add_36185 = array_index_35863[11:1] + 11'h347;
  assign sel_36187 = $signed({1'h0, add_36083, array_index_35761[0]}) < $signed({1'h0, sel_36085}) ? {add_36083, array_index_35761[0]} : sel_36085;
  assign add_36189 = array_index_35962[11:3] + 9'h0bd;
  assign sel_36192 = $signed({1'h0, add_36087, array_index_35860[2:0]}) < $signed({1'h0, sel_36090}) ? {add_36087, array_index_35860[2:0]} : sel_36090;
  assign add_36194 = array_index_35965[11:3] + 9'h0bd;
  assign sel_36197 = $signed({1'h0, add_36092, array_index_35863[2:0]}) < $signed({1'h0, sel_36095}) ? {add_36092, array_index_35863[2:0]} : sel_36095;
  assign add_36199 = array_index_36064[11:1] + 11'h247;
  assign sel_36202 = $signed({1'h0, add_36097, array_index_35962[0]}) < $signed({1'h0, sel_36100}) ? {add_36097, array_index_35962[0]} : sel_36100;
  assign add_36204 = array_index_36067[11:1] + 11'h247;
  assign sel_36207 = $signed({1'h0, add_36102, array_index_35965[0]}) < $signed({1'h0, sel_36105}) ? {add_36102, array_index_35965[0]} : sel_36105;
  assign add_36232 = array_index_36166[11:0] + 12'h247;
  assign sel_36234 = $signed({1'h0, add_36130}) < $signed({1'h0, sel_36132}) ? add_36130 : sel_36132;
  assign add_36237 = array_index_36169[11:0] + 12'h247;
  assign sel_36239 = $signed({1'h0, add_36135}) < $signed({1'h0, sel_36137}) ? add_36135 : sel_36137;
  assign array_index_36268 = set1_unflattened[5'h0b];
  assign array_index_36271 = set2_unflattened[5'h0b];
  assign add_36275 = array_index_35860[11:1] + 11'h79d;
  assign sel_36277 = $signed({1'h0, add_36173, array_index_35758[0]}) < $signed({1'h0, sel_36175}) ? {add_36173, array_index_35758[0]} : sel_36175;
  assign add_36279 = array_index_35863[11:1] + 11'h79d;
  assign sel_36281 = $signed({1'h0, add_36177, array_index_35761[0]}) < $signed({1'h0, sel_36179}) ? {add_36177, array_index_35761[0]} : sel_36179;
  assign add_36283 = array_index_35962[11:1] + 11'h347;
  assign sel_36285 = $signed({1'h0, add_36181, array_index_35860[0]}) < $signed({1'h0, sel_36183}) ? {add_36181, array_index_35860[0]} : sel_36183;
  assign add_36287 = array_index_35965[11:1] + 11'h347;
  assign sel_36289 = $signed({1'h0, add_36185, array_index_35863[0]}) < $signed({1'h0, sel_36187}) ? {add_36185, array_index_35863[0]} : sel_36187;
  assign add_36291 = array_index_36064[11:3] + 9'h0bd;
  assign sel_36294 = $signed({1'h0, add_36189, array_index_35962[2:0]}) < $signed({1'h0, sel_36192}) ? {add_36189, array_index_35962[2:0]} : sel_36192;
  assign add_36296 = array_index_36067[11:3] + 9'h0bd;
  assign sel_36299 = $signed({1'h0, add_36194, array_index_35965[2:0]}) < $signed({1'h0, sel_36197}) ? {add_36194, array_index_35965[2:0]} : sel_36197;
  assign add_36301 = array_index_36166[11:1] + 11'h247;
  assign sel_36304 = $signed({1'h0, add_36199, array_index_36064[0]}) < $signed({1'h0, sel_36202}) ? {add_36199, array_index_36064[0]} : sel_36202;
  assign add_36306 = array_index_36169[11:1] + 11'h247;
  assign sel_36309 = $signed({1'h0, add_36204, array_index_36067[0]}) < $signed({1'h0, sel_36207}) ? {add_36204, array_index_36067[0]} : sel_36207;
  assign add_36334 = array_index_36268[11:0] + 12'h247;
  assign sel_36336 = $signed({1'h0, add_36232}) < $signed({1'h0, sel_36234}) ? add_36232 : sel_36234;
  assign add_36339 = array_index_36271[11:0] + 12'h247;
  assign sel_36341 = $signed({1'h0, add_36237}) < $signed({1'h0, sel_36239}) ? add_36237 : sel_36239;
  assign array_index_36370 = set1_unflattened[5'h0c];
  assign array_index_36373 = set2_unflattened[5'h0c];
  assign add_36377 = array_index_35962[11:1] + 11'h79d;
  assign sel_36379 = $signed({1'h0, add_36275, array_index_35860[0]}) < $signed({1'h0, sel_36277}) ? {add_36275, array_index_35860[0]} : sel_36277;
  assign add_36381 = array_index_35965[11:1] + 11'h79d;
  assign sel_36383 = $signed({1'h0, add_36279, array_index_35863[0]}) < $signed({1'h0, sel_36281}) ? {add_36279, array_index_35863[0]} : sel_36281;
  assign add_36385 = array_index_36064[11:1] + 11'h347;
  assign sel_36387 = $signed({1'h0, add_36283, array_index_35962[0]}) < $signed({1'h0, sel_36285}) ? {add_36283, array_index_35962[0]} : sel_36285;
  assign add_36389 = array_index_36067[11:1] + 11'h347;
  assign sel_36391 = $signed({1'h0, add_36287, array_index_35965[0]}) < $signed({1'h0, sel_36289}) ? {add_36287, array_index_35965[0]} : sel_36289;
  assign add_36393 = array_index_36166[11:3] + 9'h0bd;
  assign sel_36396 = $signed({1'h0, add_36291, array_index_36064[2:0]}) < $signed({1'h0, sel_36294}) ? {add_36291, array_index_36064[2:0]} : sel_36294;
  assign add_36398 = array_index_36169[11:3] + 9'h0bd;
  assign sel_36401 = $signed({1'h0, add_36296, array_index_36067[2:0]}) < $signed({1'h0, sel_36299}) ? {add_36296, array_index_36067[2:0]} : sel_36299;
  assign add_36403 = array_index_36268[11:1] + 11'h247;
  assign sel_36406 = $signed({1'h0, add_36301, array_index_36166[0]}) < $signed({1'h0, sel_36304}) ? {add_36301, array_index_36166[0]} : sel_36304;
  assign add_36408 = array_index_36271[11:1] + 11'h247;
  assign sel_36411 = $signed({1'h0, add_36306, array_index_36169[0]}) < $signed({1'h0, sel_36309}) ? {add_36306, array_index_36169[0]} : sel_36309;
  assign add_36436 = array_index_36370[11:0] + 12'h247;
  assign sel_36438 = $signed({1'h0, add_36334}) < $signed({1'h0, sel_36336}) ? add_36334 : sel_36336;
  assign add_36441 = array_index_36373[11:0] + 12'h247;
  assign sel_36443 = $signed({1'h0, add_36339}) < $signed({1'h0, sel_36341}) ? add_36339 : sel_36341;
  assign array_index_36472 = set1_unflattened[5'h0d];
  assign array_index_36475 = set2_unflattened[5'h0d];
  assign add_36479 = array_index_36064[11:1] + 11'h79d;
  assign sel_36481 = $signed({1'h0, add_36377, array_index_35962[0]}) < $signed({1'h0, sel_36379}) ? {add_36377, array_index_35962[0]} : sel_36379;
  assign add_36483 = array_index_36067[11:1] + 11'h79d;
  assign sel_36485 = $signed({1'h0, add_36381, array_index_35965[0]}) < $signed({1'h0, sel_36383}) ? {add_36381, array_index_35965[0]} : sel_36383;
  assign add_36487 = array_index_36166[11:1] + 11'h347;
  assign sel_36489 = $signed({1'h0, add_36385, array_index_36064[0]}) < $signed({1'h0, sel_36387}) ? {add_36385, array_index_36064[0]} : sel_36387;
  assign add_36491 = array_index_36169[11:1] + 11'h347;
  assign sel_36493 = $signed({1'h0, add_36389, array_index_36067[0]}) < $signed({1'h0, sel_36391}) ? {add_36389, array_index_36067[0]} : sel_36391;
  assign add_36495 = array_index_36268[11:3] + 9'h0bd;
  assign sel_36498 = $signed({1'h0, add_36393, array_index_36166[2:0]}) < $signed({1'h0, sel_36396}) ? {add_36393, array_index_36166[2:0]} : sel_36396;
  assign add_36500 = array_index_36271[11:3] + 9'h0bd;
  assign sel_36503 = $signed({1'h0, add_36398, array_index_36169[2:0]}) < $signed({1'h0, sel_36401}) ? {add_36398, array_index_36169[2:0]} : sel_36401;
  assign add_36505 = array_index_36370[11:1] + 11'h247;
  assign sel_36508 = $signed({1'h0, add_36403, array_index_36268[0]}) < $signed({1'h0, sel_36406}) ? {add_36403, array_index_36268[0]} : sel_36406;
  assign add_36510 = array_index_36373[11:1] + 11'h247;
  assign sel_36513 = $signed({1'h0, add_36408, array_index_36271[0]}) < $signed({1'h0, sel_36411}) ? {add_36408, array_index_36271[0]} : sel_36411;
  assign add_36538 = array_index_36472[11:0] + 12'h247;
  assign sel_36540 = $signed({1'h0, add_36436}) < $signed({1'h0, sel_36438}) ? add_36436 : sel_36438;
  assign add_36543 = array_index_36475[11:0] + 12'h247;
  assign sel_36545 = $signed({1'h0, add_36441}) < $signed({1'h0, sel_36443}) ? add_36441 : sel_36443;
  assign array_index_36574 = set1_unflattened[5'h0e];
  assign array_index_36577 = set2_unflattened[5'h0e];
  assign add_36581 = array_index_36166[11:1] + 11'h79d;
  assign sel_36583 = $signed({1'h0, add_36479, array_index_36064[0]}) < $signed({1'h0, sel_36481}) ? {add_36479, array_index_36064[0]} : sel_36481;
  assign add_36585 = array_index_36169[11:1] + 11'h79d;
  assign sel_36587 = $signed({1'h0, add_36483, array_index_36067[0]}) < $signed({1'h0, sel_36485}) ? {add_36483, array_index_36067[0]} : sel_36485;
  assign add_36589 = array_index_36268[11:1] + 11'h347;
  assign sel_36591 = $signed({1'h0, add_36487, array_index_36166[0]}) < $signed({1'h0, sel_36489}) ? {add_36487, array_index_36166[0]} : sel_36489;
  assign add_36593 = array_index_36271[11:1] + 11'h347;
  assign sel_36595 = $signed({1'h0, add_36491, array_index_36169[0]}) < $signed({1'h0, sel_36493}) ? {add_36491, array_index_36169[0]} : sel_36493;
  assign add_36597 = array_index_36370[11:3] + 9'h0bd;
  assign sel_36600 = $signed({1'h0, add_36495, array_index_36268[2:0]}) < $signed({1'h0, sel_36498}) ? {add_36495, array_index_36268[2:0]} : sel_36498;
  assign add_36602 = array_index_36373[11:3] + 9'h0bd;
  assign sel_36605 = $signed({1'h0, add_36500, array_index_36271[2:0]}) < $signed({1'h0, sel_36503}) ? {add_36500, array_index_36271[2:0]} : sel_36503;
  assign add_36607 = array_index_36472[11:1] + 11'h247;
  assign sel_36610 = $signed({1'h0, add_36505, array_index_36370[0]}) < $signed({1'h0, sel_36508}) ? {add_36505, array_index_36370[0]} : sel_36508;
  assign add_36612 = array_index_36475[11:1] + 11'h247;
  assign sel_36615 = $signed({1'h0, add_36510, array_index_36373[0]}) < $signed({1'h0, sel_36513}) ? {add_36510, array_index_36373[0]} : sel_36513;
  assign add_36640 = array_index_36574[11:0] + 12'h247;
  assign sel_36642 = $signed({1'h0, add_36538}) < $signed({1'h0, sel_36540}) ? add_36538 : sel_36540;
  assign add_36645 = array_index_36577[11:0] + 12'h247;
  assign sel_36647 = $signed({1'h0, add_36543}) < $signed({1'h0, sel_36545}) ? add_36543 : sel_36545;
  assign array_index_36676 = set1_unflattened[5'h0f];
  assign array_index_36679 = set2_unflattened[5'h0f];
  assign add_36683 = array_index_36268[11:1] + 11'h79d;
  assign sel_36685 = $signed({1'h0, add_36581, array_index_36166[0]}) < $signed({1'h0, sel_36583}) ? {add_36581, array_index_36166[0]} : sel_36583;
  assign add_36687 = array_index_36271[11:1] + 11'h79d;
  assign sel_36689 = $signed({1'h0, add_36585, array_index_36169[0]}) < $signed({1'h0, sel_36587}) ? {add_36585, array_index_36169[0]} : sel_36587;
  assign add_36691 = array_index_36370[11:1] + 11'h347;
  assign sel_36693 = $signed({1'h0, add_36589, array_index_36268[0]}) < $signed({1'h0, sel_36591}) ? {add_36589, array_index_36268[0]} : sel_36591;
  assign add_36695 = array_index_36373[11:1] + 11'h347;
  assign sel_36697 = $signed({1'h0, add_36593, array_index_36271[0]}) < $signed({1'h0, sel_36595}) ? {add_36593, array_index_36271[0]} : sel_36595;
  assign add_36699 = array_index_36472[11:3] + 9'h0bd;
  assign sel_36702 = $signed({1'h0, add_36597, array_index_36370[2:0]}) < $signed({1'h0, sel_36600}) ? {add_36597, array_index_36370[2:0]} : sel_36600;
  assign add_36704 = array_index_36475[11:3] + 9'h0bd;
  assign sel_36707 = $signed({1'h0, add_36602, array_index_36373[2:0]}) < $signed({1'h0, sel_36605}) ? {add_36602, array_index_36373[2:0]} : sel_36605;
  assign add_36709 = array_index_36574[11:1] + 11'h247;
  assign sel_36712 = $signed({1'h0, add_36607, array_index_36472[0]}) < $signed({1'h0, sel_36610}) ? {add_36607, array_index_36472[0]} : sel_36610;
  assign add_36714 = array_index_36577[11:1] + 11'h247;
  assign sel_36717 = $signed({1'h0, add_36612, array_index_36475[0]}) < $signed({1'h0, sel_36615}) ? {add_36612, array_index_36475[0]} : sel_36615;
  assign add_36742 = array_index_36676[11:0] + 12'h247;
  assign sel_36744 = $signed({1'h0, add_36640}) < $signed({1'h0, sel_36642}) ? add_36640 : sel_36642;
  assign add_36747 = array_index_36679[11:0] + 12'h247;
  assign sel_36749 = $signed({1'h0, add_36645}) < $signed({1'h0, sel_36647}) ? add_36645 : sel_36647;
  assign array_index_36778 = set1_unflattened[5'h10];
  assign array_index_36781 = set2_unflattened[5'h10];
  assign add_36785 = array_index_36370[11:1] + 11'h79d;
  assign sel_36787 = $signed({1'h0, add_36683, array_index_36268[0]}) < $signed({1'h0, sel_36685}) ? {add_36683, array_index_36268[0]} : sel_36685;
  assign add_36789 = array_index_36373[11:1] + 11'h79d;
  assign sel_36791 = $signed({1'h0, add_36687, array_index_36271[0]}) < $signed({1'h0, sel_36689}) ? {add_36687, array_index_36271[0]} : sel_36689;
  assign add_36793 = array_index_36472[11:1] + 11'h347;
  assign sel_36795 = $signed({1'h0, add_36691, array_index_36370[0]}) < $signed({1'h0, sel_36693}) ? {add_36691, array_index_36370[0]} : sel_36693;
  assign add_36797 = array_index_36475[11:1] + 11'h347;
  assign sel_36799 = $signed({1'h0, add_36695, array_index_36373[0]}) < $signed({1'h0, sel_36697}) ? {add_36695, array_index_36373[0]} : sel_36697;
  assign add_36801 = array_index_36574[11:3] + 9'h0bd;
  assign sel_36804 = $signed({1'h0, add_36699, array_index_36472[2:0]}) < $signed({1'h0, sel_36702}) ? {add_36699, array_index_36472[2:0]} : sel_36702;
  assign add_36806 = array_index_36577[11:3] + 9'h0bd;
  assign sel_36809 = $signed({1'h0, add_36704, array_index_36475[2:0]}) < $signed({1'h0, sel_36707}) ? {add_36704, array_index_36475[2:0]} : sel_36707;
  assign add_36811 = array_index_36676[11:1] + 11'h247;
  assign sel_36814 = $signed({1'h0, add_36709, array_index_36574[0]}) < $signed({1'h0, sel_36712}) ? {add_36709, array_index_36574[0]} : sel_36712;
  assign add_36816 = array_index_36679[11:1] + 11'h247;
  assign sel_36819 = $signed({1'h0, add_36714, array_index_36577[0]}) < $signed({1'h0, sel_36717}) ? {add_36714, array_index_36577[0]} : sel_36717;
  assign add_36844 = array_index_36778[11:0] + 12'h247;
  assign sel_36846 = $signed({1'h0, add_36742}) < $signed({1'h0, sel_36744}) ? add_36742 : sel_36744;
  assign add_36849 = array_index_36781[11:0] + 12'h247;
  assign sel_36851 = $signed({1'h0, add_36747}) < $signed({1'h0, sel_36749}) ? add_36747 : sel_36749;
  assign array_index_36880 = set1_unflattened[5'h11];
  assign array_index_36883 = set2_unflattened[5'h11];
  assign add_36887 = array_index_36472[11:1] + 11'h79d;
  assign sel_36889 = $signed({1'h0, add_36785, array_index_36370[0]}) < $signed({1'h0, sel_36787}) ? {add_36785, array_index_36370[0]} : sel_36787;
  assign add_36891 = array_index_36475[11:1] + 11'h79d;
  assign sel_36893 = $signed({1'h0, add_36789, array_index_36373[0]}) < $signed({1'h0, sel_36791}) ? {add_36789, array_index_36373[0]} : sel_36791;
  assign add_36895 = array_index_36574[11:1] + 11'h347;
  assign sel_36897 = $signed({1'h0, add_36793, array_index_36472[0]}) < $signed({1'h0, sel_36795}) ? {add_36793, array_index_36472[0]} : sel_36795;
  assign add_36899 = array_index_36577[11:1] + 11'h347;
  assign sel_36901 = $signed({1'h0, add_36797, array_index_36475[0]}) < $signed({1'h0, sel_36799}) ? {add_36797, array_index_36475[0]} : sel_36799;
  assign add_36903 = array_index_36676[11:3] + 9'h0bd;
  assign sel_36906 = $signed({1'h0, add_36801, array_index_36574[2:0]}) < $signed({1'h0, sel_36804}) ? {add_36801, array_index_36574[2:0]} : sel_36804;
  assign add_36908 = array_index_36679[11:3] + 9'h0bd;
  assign sel_36911 = $signed({1'h0, add_36806, array_index_36577[2:0]}) < $signed({1'h0, sel_36809}) ? {add_36806, array_index_36577[2:0]} : sel_36809;
  assign add_36913 = array_index_36778[11:1] + 11'h247;
  assign sel_36916 = $signed({1'h0, add_36811, array_index_36676[0]}) < $signed({1'h0, sel_36814}) ? {add_36811, array_index_36676[0]} : sel_36814;
  assign add_36918 = array_index_36781[11:1] + 11'h247;
  assign sel_36921 = $signed({1'h0, add_36816, array_index_36679[0]}) < $signed({1'h0, sel_36819}) ? {add_36816, array_index_36679[0]} : sel_36819;
  assign add_36946 = array_index_36880[11:0] + 12'h247;
  assign sel_36948 = $signed({1'h0, add_36844}) < $signed({1'h0, sel_36846}) ? add_36844 : sel_36846;
  assign add_36951 = array_index_36883[11:0] + 12'h247;
  assign sel_36953 = $signed({1'h0, add_36849}) < $signed({1'h0, sel_36851}) ? add_36849 : sel_36851;
  assign array_index_36982 = set1_unflattened[5'h12];
  assign array_index_36985 = set2_unflattened[5'h12];
  assign add_36989 = array_index_36574[11:1] + 11'h79d;
  assign sel_36991 = $signed({1'h0, add_36887, array_index_36472[0]}) < $signed({1'h0, sel_36889}) ? {add_36887, array_index_36472[0]} : sel_36889;
  assign add_36993 = array_index_36577[11:1] + 11'h79d;
  assign sel_36995 = $signed({1'h0, add_36891, array_index_36475[0]}) < $signed({1'h0, sel_36893}) ? {add_36891, array_index_36475[0]} : sel_36893;
  assign add_36997 = array_index_36676[11:1] + 11'h347;
  assign sel_36999 = $signed({1'h0, add_36895, array_index_36574[0]}) < $signed({1'h0, sel_36897}) ? {add_36895, array_index_36574[0]} : sel_36897;
  assign add_37001 = array_index_36679[11:1] + 11'h347;
  assign sel_37003 = $signed({1'h0, add_36899, array_index_36577[0]}) < $signed({1'h0, sel_36901}) ? {add_36899, array_index_36577[0]} : sel_36901;
  assign add_37005 = array_index_36778[11:3] + 9'h0bd;
  assign sel_37008 = $signed({1'h0, add_36903, array_index_36676[2:0]}) < $signed({1'h0, sel_36906}) ? {add_36903, array_index_36676[2:0]} : sel_36906;
  assign add_37010 = array_index_36781[11:3] + 9'h0bd;
  assign sel_37013 = $signed({1'h0, add_36908, array_index_36679[2:0]}) < $signed({1'h0, sel_36911}) ? {add_36908, array_index_36679[2:0]} : sel_36911;
  assign add_37015 = array_index_36880[11:1] + 11'h247;
  assign sel_37018 = $signed({1'h0, add_36913, array_index_36778[0]}) < $signed({1'h0, sel_36916}) ? {add_36913, array_index_36778[0]} : sel_36916;
  assign add_37020 = array_index_36883[11:1] + 11'h247;
  assign sel_37023 = $signed({1'h0, add_36918, array_index_36781[0]}) < $signed({1'h0, sel_36921}) ? {add_36918, array_index_36781[0]} : sel_36921;
  assign add_37048 = array_index_36982[11:0] + 12'h247;
  assign sel_37050 = $signed({1'h0, add_36946}) < $signed({1'h0, sel_36948}) ? add_36946 : sel_36948;
  assign add_37053 = array_index_36985[11:0] + 12'h247;
  assign sel_37055 = $signed({1'h0, add_36951}) < $signed({1'h0, sel_36953}) ? add_36951 : sel_36953;
  assign array_index_37084 = set1_unflattened[5'h13];
  assign array_index_37087 = set2_unflattened[5'h13];
  assign add_37091 = array_index_36676[11:1] + 11'h79d;
  assign sel_37093 = $signed({1'h0, add_36989, array_index_36574[0]}) < $signed({1'h0, sel_36991}) ? {add_36989, array_index_36574[0]} : sel_36991;
  assign add_37095 = array_index_36679[11:1] + 11'h79d;
  assign sel_37097 = $signed({1'h0, add_36993, array_index_36577[0]}) < $signed({1'h0, sel_36995}) ? {add_36993, array_index_36577[0]} : sel_36995;
  assign add_37099 = array_index_36778[11:1] + 11'h347;
  assign sel_37101 = $signed({1'h0, add_36997, array_index_36676[0]}) < $signed({1'h0, sel_36999}) ? {add_36997, array_index_36676[0]} : sel_36999;
  assign add_37103 = array_index_36781[11:1] + 11'h347;
  assign sel_37105 = $signed({1'h0, add_37001, array_index_36679[0]}) < $signed({1'h0, sel_37003}) ? {add_37001, array_index_36679[0]} : sel_37003;
  assign add_37107 = array_index_36880[11:3] + 9'h0bd;
  assign sel_37110 = $signed({1'h0, add_37005, array_index_36778[2:0]}) < $signed({1'h0, sel_37008}) ? {add_37005, array_index_36778[2:0]} : sel_37008;
  assign add_37112 = array_index_36883[11:3] + 9'h0bd;
  assign sel_37115 = $signed({1'h0, add_37010, array_index_36781[2:0]}) < $signed({1'h0, sel_37013}) ? {add_37010, array_index_36781[2:0]} : sel_37013;
  assign add_37117 = array_index_36982[11:1] + 11'h247;
  assign sel_37120 = $signed({1'h0, add_37015, array_index_36880[0]}) < $signed({1'h0, sel_37018}) ? {add_37015, array_index_36880[0]} : sel_37018;
  assign add_37122 = array_index_36985[11:1] + 11'h247;
  assign sel_37125 = $signed({1'h0, add_37020, array_index_36883[0]}) < $signed({1'h0, sel_37023}) ? {add_37020, array_index_36883[0]} : sel_37023;
  assign add_37149 = array_index_37084[11:0] + 12'h247;
  assign sel_37151 = $signed({1'h0, add_37048}) < $signed({1'h0, sel_37050}) ? add_37048 : sel_37050;
  assign add_37153 = array_index_37087[11:0] + 12'h247;
  assign sel_37155 = $signed({1'h0, add_37053}) < $signed({1'h0, sel_37055}) ? add_37053 : sel_37055;
  assign add_37189 = array_index_36778[11:1] + 11'h79d;
  assign sel_37191 = $signed({1'h0, add_37091, array_index_36676[0]}) < $signed({1'h0, sel_37093}) ? {add_37091, array_index_36676[0]} : sel_37093;
  assign add_37193 = array_index_36781[11:1] + 11'h79d;
  assign sel_37195 = $signed({1'h0, add_37095, array_index_36679[0]}) < $signed({1'h0, sel_37097}) ? {add_37095, array_index_36679[0]} : sel_37097;
  assign add_37197 = array_index_36880[11:1] + 11'h347;
  assign sel_37199 = $signed({1'h0, add_37099, array_index_36778[0]}) < $signed({1'h0, sel_37101}) ? {add_37099, array_index_36778[0]} : sel_37101;
  assign add_37201 = array_index_36883[11:1] + 11'h347;
  assign sel_37203 = $signed({1'h0, add_37103, array_index_36781[0]}) < $signed({1'h0, sel_37105}) ? {add_37103, array_index_36781[0]} : sel_37105;
  assign add_37205 = array_index_36982[11:3] + 9'h0bd;
  assign sel_37208 = $signed({1'h0, add_37107, array_index_36880[2:0]}) < $signed({1'h0, sel_37110}) ? {add_37107, array_index_36880[2:0]} : sel_37110;
  assign add_37210 = array_index_36985[11:3] + 9'h0bd;
  assign sel_37213 = $signed({1'h0, add_37112, array_index_36883[2:0]}) < $signed({1'h0, sel_37115}) ? {add_37112, array_index_36883[2:0]} : sel_37115;
  assign add_37215 = array_index_37084[11:1] + 11'h247;
  assign sel_37218 = $signed({1'h0, add_37117, array_index_36982[0]}) < $signed({1'h0, sel_37120}) ? {add_37117, array_index_36982[0]} : sel_37120;
  assign add_37220 = array_index_37087[11:1] + 11'h247;
  assign sel_37223 = $signed({1'h0, add_37122, array_index_36985[0]}) < $signed({1'h0, sel_37125}) ? {add_37122, array_index_36985[0]} : sel_37125;
  assign add_37271 = array_index_36880[11:1] + 11'h79d;
  assign sel_37273 = $signed({1'h0, add_37189, array_index_36778[0]}) < $signed({1'h0, sel_37191}) ? {add_37189, array_index_36778[0]} : sel_37191;
  assign add_37275 = array_index_36883[11:1] + 11'h79d;
  assign sel_37277 = $signed({1'h0, add_37193, array_index_36781[0]}) < $signed({1'h0, sel_37195}) ? {add_37193, array_index_36781[0]} : sel_37195;
  assign add_37279 = array_index_36982[11:1] + 11'h347;
  assign sel_37281 = $signed({1'h0, add_37197, array_index_36880[0]}) < $signed({1'h0, sel_37199}) ? {add_37197, array_index_36880[0]} : sel_37199;
  assign add_37283 = array_index_36985[11:1] + 11'h347;
  assign sel_37285 = $signed({1'h0, add_37201, array_index_36883[0]}) < $signed({1'h0, sel_37203}) ? {add_37201, array_index_36883[0]} : sel_37203;
  assign add_37287 = array_index_37084[11:3] + 9'h0bd;
  assign sel_37290 = $signed({1'h0, add_37205, array_index_36982[2:0]}) < $signed({1'h0, sel_37208}) ? {add_37205, array_index_36982[2:0]} : sel_37208;
  assign add_37292 = array_index_37087[11:3] + 9'h0bd;
  assign sel_37295 = $signed({1'h0, add_37210, array_index_36985[2:0]}) < $signed({1'h0, sel_37213}) ? {add_37210, array_index_36985[2:0]} : sel_37213;
  assign concat_37298 = {1'h0, ($signed({1'h0, add_37149}) < $signed({1'h0, sel_37151}) ? add_37149 : sel_37151) == ($signed({1'h0, add_37153}) < $signed({1'h0, sel_37155}) ? add_37153 : sel_37155)};
  assign add_37313 = concat_37298 + 2'h1;
  assign add_37333 = array_index_36982[11:1] + 11'h79d;
  assign sel_37335 = $signed({1'h0, add_37271, array_index_36880[0]}) < $signed({1'h0, sel_37273}) ? {add_37271, array_index_36880[0]} : sel_37273;
  assign add_37337 = array_index_36985[11:1] + 11'h79d;
  assign sel_37339 = $signed({1'h0, add_37275, array_index_36883[0]}) < $signed({1'h0, sel_37277}) ? {add_37275, array_index_36883[0]} : sel_37277;
  assign add_37341 = array_index_37084[11:1] + 11'h347;
  assign sel_37343 = $signed({1'h0, add_37279, array_index_36982[0]}) < $signed({1'h0, sel_37281}) ? {add_37279, array_index_36982[0]} : sel_37281;
  assign add_37345 = array_index_37087[11:1] + 11'h347;
  assign sel_37347 = $signed({1'h0, add_37283, array_index_36985[0]}) < $signed({1'h0, sel_37285}) ? {add_37283, array_index_36985[0]} : sel_37285;
  assign concat_37350 = {1'h0, ($signed({1'h0, add_37215, array_index_37084[0]}) < $signed({1'h0, sel_37218}) ? {add_37215, array_index_37084[0]} : sel_37218) == ($signed({1'h0, add_37220, array_index_37087[0]}) < $signed({1'h0, sel_37223}) ? {add_37220, array_index_37087[0]} : sel_37223) ? add_37313 : concat_37298};
  assign add_37361 = concat_37350 + 3'h1;
  assign add_37375 = array_index_37084[11:1] + 11'h79d;
  assign sel_37377 = $signed({1'h0, add_37333, array_index_36982[0]}) < $signed({1'h0, sel_37335}) ? {add_37333, array_index_36982[0]} : sel_37335;
  assign add_37379 = array_index_37087[11:1] + 11'h79d;
  assign sel_37381 = $signed({1'h0, add_37337, array_index_36985[0]}) < $signed({1'h0, sel_37339}) ? {add_37337, array_index_36985[0]} : sel_37339;
  assign concat_37384 = {1'h0, ($signed({1'h0, add_37287, array_index_37084[2:0]}) < $signed({1'h0, sel_37290}) ? {add_37287, array_index_37084[2:0]} : sel_37290) == ($signed({1'h0, add_37292, array_index_37087[2:0]}) < $signed({1'h0, sel_37295}) ? {add_37292, array_index_37087[2:0]} : sel_37295) ? add_37361 : concat_37350};
  assign add_37391 = concat_37384 + 4'h1;
  assign concat_37400 = {1'h0, ($signed({1'h0, add_37341, array_index_37084[0]}) < $signed({1'h0, sel_37343}) ? {add_37341, array_index_37084[0]} : sel_37343) == ($signed({1'h0, add_37345, array_index_37087[0]}) < $signed({1'h0, sel_37347}) ? {add_37345, array_index_37087[0]} : sel_37347) ? add_37391 : concat_37384};
  assign add_37403 = concat_37400 + 5'h01;
  assign out = {{11'h000, ($signed({1'h0, add_37375, array_index_37084[0]}) < $signed({1'h0, sel_37377}) ? {add_37375, array_index_37084[0]} : sel_37377) == ($signed({1'h0, add_37379, array_index_37087[0]}) < $signed({1'h0, sel_37381}) ? {add_37379, array_index_37087[0]} : sel_37381) ? add_37403 : concat_37400}, {set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
