module min_hash(
  input wire [1599:0] set1,
  input wire [1599:0] set2,
  output wire [3207:0] out
);
  wire [15:0] set1_unflattened[100];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  assign set1_unflattened[30] = set1[495:480];
  assign set1_unflattened[31] = set1[511:496];
  assign set1_unflattened[32] = set1[527:512];
  assign set1_unflattened[33] = set1[543:528];
  assign set1_unflattened[34] = set1[559:544];
  assign set1_unflattened[35] = set1[575:560];
  assign set1_unflattened[36] = set1[591:576];
  assign set1_unflattened[37] = set1[607:592];
  assign set1_unflattened[38] = set1[623:608];
  assign set1_unflattened[39] = set1[639:624];
  assign set1_unflattened[40] = set1[655:640];
  assign set1_unflattened[41] = set1[671:656];
  assign set1_unflattened[42] = set1[687:672];
  assign set1_unflattened[43] = set1[703:688];
  assign set1_unflattened[44] = set1[719:704];
  assign set1_unflattened[45] = set1[735:720];
  assign set1_unflattened[46] = set1[751:736];
  assign set1_unflattened[47] = set1[767:752];
  assign set1_unflattened[48] = set1[783:768];
  assign set1_unflattened[49] = set1[799:784];
  assign set1_unflattened[50] = set1[815:800];
  assign set1_unflattened[51] = set1[831:816];
  assign set1_unflattened[52] = set1[847:832];
  assign set1_unflattened[53] = set1[863:848];
  assign set1_unflattened[54] = set1[879:864];
  assign set1_unflattened[55] = set1[895:880];
  assign set1_unflattened[56] = set1[911:896];
  assign set1_unflattened[57] = set1[927:912];
  assign set1_unflattened[58] = set1[943:928];
  assign set1_unflattened[59] = set1[959:944];
  assign set1_unflattened[60] = set1[975:960];
  assign set1_unflattened[61] = set1[991:976];
  assign set1_unflattened[62] = set1[1007:992];
  assign set1_unflattened[63] = set1[1023:1008];
  assign set1_unflattened[64] = set1[1039:1024];
  assign set1_unflattened[65] = set1[1055:1040];
  assign set1_unflattened[66] = set1[1071:1056];
  assign set1_unflattened[67] = set1[1087:1072];
  assign set1_unflattened[68] = set1[1103:1088];
  assign set1_unflattened[69] = set1[1119:1104];
  assign set1_unflattened[70] = set1[1135:1120];
  assign set1_unflattened[71] = set1[1151:1136];
  assign set1_unflattened[72] = set1[1167:1152];
  assign set1_unflattened[73] = set1[1183:1168];
  assign set1_unflattened[74] = set1[1199:1184];
  assign set1_unflattened[75] = set1[1215:1200];
  assign set1_unflattened[76] = set1[1231:1216];
  assign set1_unflattened[77] = set1[1247:1232];
  assign set1_unflattened[78] = set1[1263:1248];
  assign set1_unflattened[79] = set1[1279:1264];
  assign set1_unflattened[80] = set1[1295:1280];
  assign set1_unflattened[81] = set1[1311:1296];
  assign set1_unflattened[82] = set1[1327:1312];
  assign set1_unflattened[83] = set1[1343:1328];
  assign set1_unflattened[84] = set1[1359:1344];
  assign set1_unflattened[85] = set1[1375:1360];
  assign set1_unflattened[86] = set1[1391:1376];
  assign set1_unflattened[87] = set1[1407:1392];
  assign set1_unflattened[88] = set1[1423:1408];
  assign set1_unflattened[89] = set1[1439:1424];
  assign set1_unflattened[90] = set1[1455:1440];
  assign set1_unflattened[91] = set1[1471:1456];
  assign set1_unflattened[92] = set1[1487:1472];
  assign set1_unflattened[93] = set1[1503:1488];
  assign set1_unflattened[94] = set1[1519:1504];
  assign set1_unflattened[95] = set1[1535:1520];
  assign set1_unflattened[96] = set1[1551:1536];
  assign set1_unflattened[97] = set1[1567:1552];
  assign set1_unflattened[98] = set1[1583:1568];
  assign set1_unflattened[99] = set1[1599:1584];
  wire [15:0] set2_unflattened[100];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  assign set2_unflattened[30] = set2[495:480];
  assign set2_unflattened[31] = set2[511:496];
  assign set2_unflattened[32] = set2[527:512];
  assign set2_unflattened[33] = set2[543:528];
  assign set2_unflattened[34] = set2[559:544];
  assign set2_unflattened[35] = set2[575:560];
  assign set2_unflattened[36] = set2[591:576];
  assign set2_unflattened[37] = set2[607:592];
  assign set2_unflattened[38] = set2[623:608];
  assign set2_unflattened[39] = set2[639:624];
  assign set2_unflattened[40] = set2[655:640];
  assign set2_unflattened[41] = set2[671:656];
  assign set2_unflattened[42] = set2[687:672];
  assign set2_unflattened[43] = set2[703:688];
  assign set2_unflattened[44] = set2[719:704];
  assign set2_unflattened[45] = set2[735:720];
  assign set2_unflattened[46] = set2[751:736];
  assign set2_unflattened[47] = set2[767:752];
  assign set2_unflattened[48] = set2[783:768];
  assign set2_unflattened[49] = set2[799:784];
  assign set2_unflattened[50] = set2[815:800];
  assign set2_unflattened[51] = set2[831:816];
  assign set2_unflattened[52] = set2[847:832];
  assign set2_unflattened[53] = set2[863:848];
  assign set2_unflattened[54] = set2[879:864];
  assign set2_unflattened[55] = set2[895:880];
  assign set2_unflattened[56] = set2[911:896];
  assign set2_unflattened[57] = set2[927:912];
  assign set2_unflattened[58] = set2[943:928];
  assign set2_unflattened[59] = set2[959:944];
  assign set2_unflattened[60] = set2[975:960];
  assign set2_unflattened[61] = set2[991:976];
  assign set2_unflattened[62] = set2[1007:992];
  assign set2_unflattened[63] = set2[1023:1008];
  assign set2_unflattened[64] = set2[1039:1024];
  assign set2_unflattened[65] = set2[1055:1040];
  assign set2_unflattened[66] = set2[1071:1056];
  assign set2_unflattened[67] = set2[1087:1072];
  assign set2_unflattened[68] = set2[1103:1088];
  assign set2_unflattened[69] = set2[1119:1104];
  assign set2_unflattened[70] = set2[1135:1120];
  assign set2_unflattened[71] = set2[1151:1136];
  assign set2_unflattened[72] = set2[1167:1152];
  assign set2_unflattened[73] = set2[1183:1168];
  assign set2_unflattened[74] = set2[1199:1184];
  assign set2_unflattened[75] = set2[1215:1200];
  assign set2_unflattened[76] = set2[1231:1216];
  assign set2_unflattened[77] = set2[1247:1232];
  assign set2_unflattened[78] = set2[1263:1248];
  assign set2_unflattened[79] = set2[1279:1264];
  assign set2_unflattened[80] = set2[1295:1280];
  assign set2_unflattened[81] = set2[1311:1296];
  assign set2_unflattened[82] = set2[1327:1312];
  assign set2_unflattened[83] = set2[1343:1328];
  assign set2_unflattened[84] = set2[1359:1344];
  assign set2_unflattened[85] = set2[1375:1360];
  assign set2_unflattened[86] = set2[1391:1376];
  assign set2_unflattened[87] = set2[1407:1392];
  assign set2_unflattened[88] = set2[1423:1408];
  assign set2_unflattened[89] = set2[1439:1424];
  assign set2_unflattened[90] = set2[1455:1440];
  assign set2_unflattened[91] = set2[1471:1456];
  assign set2_unflattened[92] = set2[1487:1472];
  assign set2_unflattened[93] = set2[1503:1488];
  assign set2_unflattened[94] = set2[1519:1504];
  assign set2_unflattened[95] = set2[1535:1520];
  assign set2_unflattened[96] = set2[1551:1536];
  assign set2_unflattened[97] = set2[1567:1552];
  assign set2_unflattened[98] = set2[1583:1568];
  assign set2_unflattened[99] = set2[1599:1584];
  wire [15:0] array_index_948482;
  wire [15:0] array_index_948483;
  wire [15:0] array_index_948487;
  wire [1:0] concat_948488;
  wire [1:0] add_948491;
  wire [15:0] array_index_948495;
  wire [2:0] concat_948496;
  wire [2:0] add_948499;
  wire [15:0] array_index_948503;
  wire [3:0] concat_948504;
  wire [3:0] add_948507;
  wire [15:0] array_index_948511;
  wire [4:0] concat_948512;
  wire [4:0] add_948515;
  wire [15:0] array_index_948519;
  wire [5:0] concat_948520;
  wire [5:0] add_948523;
  wire [15:0] array_index_948527;
  wire [6:0] concat_948528;
  wire [6:0] add_948531;
  wire [15:0] array_index_948535;
  wire [7:0] concat_948536;
  wire [7:0] add_948540;
  wire [15:0] array_index_948541;
  wire [7:0] sel_948542;
  wire [7:0] add_948546;
  wire [15:0] array_index_948547;
  wire [7:0] sel_948548;
  wire [7:0] add_948552;
  wire [15:0] array_index_948553;
  wire [7:0] sel_948554;
  wire [7:0] add_948558;
  wire [15:0] array_index_948559;
  wire [7:0] sel_948560;
  wire [7:0] add_948564;
  wire [15:0] array_index_948565;
  wire [7:0] sel_948566;
  wire [7:0] add_948570;
  wire [15:0] array_index_948571;
  wire [7:0] sel_948572;
  wire [7:0] add_948576;
  wire [15:0] array_index_948577;
  wire [7:0] sel_948578;
  wire [7:0] add_948582;
  wire [15:0] array_index_948583;
  wire [7:0] sel_948584;
  wire [7:0] add_948588;
  wire [15:0] array_index_948589;
  wire [7:0] sel_948590;
  wire [7:0] add_948594;
  wire [15:0] array_index_948595;
  wire [7:0] sel_948596;
  wire [7:0] add_948600;
  wire [15:0] array_index_948601;
  wire [7:0] sel_948602;
  wire [7:0] add_948606;
  wire [15:0] array_index_948607;
  wire [7:0] sel_948608;
  wire [7:0] add_948612;
  wire [15:0] array_index_948613;
  wire [7:0] sel_948614;
  wire [7:0] add_948618;
  wire [15:0] array_index_948619;
  wire [7:0] sel_948620;
  wire [7:0] add_948624;
  wire [15:0] array_index_948625;
  wire [7:0] sel_948626;
  wire [7:0] add_948630;
  wire [15:0] array_index_948631;
  wire [7:0] sel_948632;
  wire [7:0] add_948636;
  wire [15:0] array_index_948637;
  wire [7:0] sel_948638;
  wire [7:0] add_948642;
  wire [15:0] array_index_948643;
  wire [7:0] sel_948644;
  wire [7:0] add_948648;
  wire [15:0] array_index_948649;
  wire [7:0] sel_948650;
  wire [7:0] add_948654;
  wire [15:0] array_index_948655;
  wire [7:0] sel_948656;
  wire [7:0] add_948660;
  wire [15:0] array_index_948661;
  wire [7:0] sel_948662;
  wire [7:0] add_948666;
  wire [15:0] array_index_948667;
  wire [7:0] sel_948668;
  wire [7:0] add_948672;
  wire [15:0] array_index_948673;
  wire [7:0] sel_948674;
  wire [7:0] add_948678;
  wire [15:0] array_index_948679;
  wire [7:0] sel_948680;
  wire [7:0] add_948684;
  wire [15:0] array_index_948685;
  wire [7:0] sel_948686;
  wire [7:0] add_948690;
  wire [15:0] array_index_948691;
  wire [7:0] sel_948692;
  wire [7:0] add_948696;
  wire [15:0] array_index_948697;
  wire [7:0] sel_948698;
  wire [7:0] add_948702;
  wire [15:0] array_index_948703;
  wire [7:0] sel_948704;
  wire [7:0] add_948708;
  wire [15:0] array_index_948709;
  wire [7:0] sel_948710;
  wire [7:0] add_948714;
  wire [15:0] array_index_948715;
  wire [7:0] sel_948716;
  wire [7:0] add_948720;
  wire [15:0] array_index_948721;
  wire [7:0] sel_948722;
  wire [7:0] add_948726;
  wire [15:0] array_index_948727;
  wire [7:0] sel_948728;
  wire [7:0] add_948732;
  wire [15:0] array_index_948733;
  wire [7:0] sel_948734;
  wire [7:0] add_948738;
  wire [15:0] array_index_948739;
  wire [7:0] sel_948740;
  wire [7:0] add_948744;
  wire [15:0] array_index_948745;
  wire [7:0] sel_948746;
  wire [7:0] add_948750;
  wire [15:0] array_index_948751;
  wire [7:0] sel_948752;
  wire [7:0] add_948756;
  wire [15:0] array_index_948757;
  wire [7:0] sel_948758;
  wire [7:0] add_948762;
  wire [15:0] array_index_948763;
  wire [7:0] sel_948764;
  wire [7:0] add_948768;
  wire [15:0] array_index_948769;
  wire [7:0] sel_948770;
  wire [7:0] add_948774;
  wire [15:0] array_index_948775;
  wire [7:0] sel_948776;
  wire [7:0] add_948780;
  wire [15:0] array_index_948781;
  wire [7:0] sel_948782;
  wire [7:0] add_948786;
  wire [15:0] array_index_948787;
  wire [7:0] sel_948788;
  wire [7:0] add_948792;
  wire [15:0] array_index_948793;
  wire [7:0] sel_948794;
  wire [7:0] add_948798;
  wire [15:0] array_index_948799;
  wire [7:0] sel_948800;
  wire [7:0] add_948804;
  wire [15:0] array_index_948805;
  wire [7:0] sel_948806;
  wire [7:0] add_948810;
  wire [15:0] array_index_948811;
  wire [7:0] sel_948812;
  wire [7:0] add_948816;
  wire [15:0] array_index_948817;
  wire [7:0] sel_948818;
  wire [7:0] add_948822;
  wire [15:0] array_index_948823;
  wire [7:0] sel_948824;
  wire [7:0] add_948828;
  wire [15:0] array_index_948829;
  wire [7:0] sel_948830;
  wire [7:0] add_948834;
  wire [15:0] array_index_948835;
  wire [7:0] sel_948836;
  wire [7:0] add_948840;
  wire [15:0] array_index_948841;
  wire [7:0] sel_948842;
  wire [7:0] add_948846;
  wire [15:0] array_index_948847;
  wire [7:0] sel_948848;
  wire [7:0] add_948852;
  wire [15:0] array_index_948853;
  wire [7:0] sel_948854;
  wire [7:0] add_948858;
  wire [15:0] array_index_948859;
  wire [7:0] sel_948860;
  wire [7:0] add_948864;
  wire [15:0] array_index_948865;
  wire [7:0] sel_948866;
  wire [7:0] add_948870;
  wire [15:0] array_index_948871;
  wire [7:0] sel_948872;
  wire [7:0] add_948876;
  wire [15:0] array_index_948877;
  wire [7:0] sel_948878;
  wire [7:0] add_948882;
  wire [15:0] array_index_948883;
  wire [7:0] sel_948884;
  wire [7:0] add_948888;
  wire [15:0] array_index_948889;
  wire [7:0] sel_948890;
  wire [7:0] add_948894;
  wire [15:0] array_index_948895;
  wire [7:0] sel_948896;
  wire [7:0] add_948900;
  wire [15:0] array_index_948901;
  wire [7:0] sel_948902;
  wire [7:0] add_948906;
  wire [15:0] array_index_948907;
  wire [7:0] sel_948908;
  wire [7:0] add_948912;
  wire [15:0] array_index_948913;
  wire [7:0] sel_948914;
  wire [7:0] add_948918;
  wire [15:0] array_index_948919;
  wire [7:0] sel_948920;
  wire [7:0] add_948924;
  wire [15:0] array_index_948925;
  wire [7:0] sel_948926;
  wire [7:0] add_948930;
  wire [15:0] array_index_948931;
  wire [7:0] sel_948932;
  wire [7:0] add_948936;
  wire [15:0] array_index_948937;
  wire [7:0] sel_948938;
  wire [7:0] add_948942;
  wire [15:0] array_index_948943;
  wire [7:0] sel_948944;
  wire [7:0] add_948948;
  wire [15:0] array_index_948949;
  wire [7:0] sel_948950;
  wire [7:0] add_948954;
  wire [15:0] array_index_948955;
  wire [7:0] sel_948956;
  wire [7:0] add_948960;
  wire [15:0] array_index_948961;
  wire [7:0] sel_948962;
  wire [7:0] add_948966;
  wire [15:0] array_index_948967;
  wire [7:0] sel_948968;
  wire [7:0] add_948972;
  wire [15:0] array_index_948973;
  wire [7:0] sel_948974;
  wire [7:0] add_948978;
  wire [15:0] array_index_948979;
  wire [7:0] sel_948980;
  wire [7:0] add_948984;
  wire [15:0] array_index_948985;
  wire [7:0] sel_948986;
  wire [7:0] add_948990;
  wire [15:0] array_index_948991;
  wire [7:0] sel_948992;
  wire [7:0] add_948996;
  wire [15:0] array_index_948997;
  wire [7:0] sel_948998;
  wire [7:0] add_949002;
  wire [15:0] array_index_949003;
  wire [7:0] sel_949004;
  wire [7:0] add_949008;
  wire [15:0] array_index_949009;
  wire [7:0] sel_949010;
  wire [7:0] add_949014;
  wire [15:0] array_index_949015;
  wire [7:0] sel_949016;
  wire [7:0] add_949020;
  wire [15:0] array_index_949021;
  wire [7:0] sel_949022;
  wire [7:0] add_949026;
  wire [15:0] array_index_949027;
  wire [7:0] sel_949028;
  wire [7:0] add_949032;
  wire [15:0] array_index_949033;
  wire [7:0] sel_949034;
  wire [7:0] add_949038;
  wire [15:0] array_index_949039;
  wire [7:0] sel_949040;
  wire [7:0] add_949044;
  wire [15:0] array_index_949045;
  wire [7:0] sel_949046;
  wire [7:0] add_949050;
  wire [15:0] array_index_949051;
  wire [7:0] sel_949052;
  wire [7:0] add_949056;
  wire [15:0] array_index_949057;
  wire [7:0] sel_949058;
  wire [7:0] add_949062;
  wire [15:0] array_index_949063;
  wire [7:0] sel_949064;
  wire [7:0] add_949068;
  wire [15:0] array_index_949069;
  wire [7:0] sel_949070;
  wire [7:0] add_949074;
  wire [15:0] array_index_949075;
  wire [7:0] sel_949076;
  wire [7:0] add_949080;
  wire [15:0] array_index_949081;
  wire [7:0] sel_949082;
  wire [7:0] add_949086;
  wire [15:0] array_index_949087;
  wire [7:0] sel_949088;
  wire [7:0] add_949092;
  wire [15:0] array_index_949093;
  wire [7:0] sel_949094;
  wire [7:0] add_949097;
  wire [7:0] sel_949098;
  wire [7:0] add_949101;
  wire [7:0] sel_949102;
  wire [7:0] add_949105;
  wire [7:0] sel_949106;
  wire [7:0] add_949109;
  wire [7:0] sel_949110;
  wire [7:0] add_949113;
  wire [7:0] sel_949114;
  wire [7:0] add_949117;
  wire [7:0] sel_949118;
  wire [7:0] add_949121;
  wire [7:0] sel_949122;
  wire [7:0] add_949125;
  wire [7:0] sel_949126;
  wire [7:0] add_949129;
  wire [7:0] sel_949130;
  wire [7:0] add_949133;
  wire [7:0] sel_949134;
  wire [7:0] add_949137;
  wire [7:0] sel_949138;
  wire [7:0] add_949141;
  wire [7:0] sel_949142;
  wire [7:0] add_949145;
  wire [7:0] sel_949146;
  wire [7:0] add_949149;
  wire [7:0] sel_949150;
  wire [7:0] add_949153;
  wire [7:0] sel_949154;
  wire [7:0] add_949157;
  wire [7:0] sel_949158;
  wire [7:0] add_949161;
  wire [7:0] sel_949162;
  wire [7:0] add_949165;
  wire [7:0] sel_949166;
  wire [7:0] add_949169;
  wire [7:0] sel_949170;
  wire [7:0] add_949173;
  wire [7:0] sel_949174;
  wire [7:0] add_949177;
  wire [7:0] sel_949178;
  wire [7:0] add_949181;
  wire [7:0] sel_949182;
  wire [7:0] add_949185;
  wire [7:0] sel_949186;
  wire [7:0] add_949189;
  wire [7:0] sel_949190;
  wire [7:0] add_949193;
  wire [7:0] sel_949194;
  wire [7:0] add_949197;
  wire [7:0] sel_949198;
  wire [7:0] add_949201;
  wire [7:0] sel_949202;
  wire [7:0] add_949205;
  wire [7:0] sel_949206;
  wire [7:0] add_949209;
  wire [7:0] sel_949210;
  wire [7:0] add_949213;
  wire [7:0] sel_949214;
  wire [7:0] add_949217;
  wire [7:0] sel_949218;
  wire [7:0] add_949221;
  wire [7:0] sel_949222;
  wire [7:0] add_949225;
  wire [7:0] sel_949226;
  wire [7:0] add_949229;
  wire [7:0] sel_949230;
  wire [7:0] add_949233;
  wire [7:0] sel_949234;
  wire [7:0] add_949237;
  wire [7:0] sel_949238;
  wire [7:0] add_949241;
  wire [7:0] sel_949242;
  wire [7:0] add_949245;
  wire [7:0] sel_949246;
  wire [7:0] add_949249;
  wire [7:0] sel_949250;
  wire [7:0] add_949253;
  wire [7:0] sel_949254;
  wire [7:0] add_949257;
  wire [7:0] sel_949258;
  wire [7:0] add_949261;
  wire [7:0] sel_949262;
  wire [7:0] add_949265;
  wire [7:0] sel_949266;
  wire [7:0] add_949269;
  wire [7:0] sel_949270;
  wire [7:0] add_949273;
  wire [7:0] sel_949274;
  wire [7:0] add_949277;
  wire [7:0] sel_949278;
  wire [7:0] add_949281;
  wire [7:0] sel_949282;
  wire [7:0] add_949285;
  wire [7:0] sel_949286;
  wire [7:0] add_949289;
  wire [7:0] sel_949290;
  wire [7:0] add_949293;
  wire [7:0] sel_949294;
  wire [7:0] add_949297;
  wire [7:0] sel_949298;
  wire [7:0] add_949301;
  wire [7:0] sel_949302;
  wire [7:0] add_949305;
  wire [7:0] sel_949306;
  wire [7:0] add_949309;
  wire [7:0] sel_949310;
  wire [7:0] add_949313;
  wire [7:0] sel_949314;
  wire [7:0] add_949317;
  wire [7:0] sel_949318;
  wire [7:0] add_949321;
  wire [7:0] sel_949322;
  wire [7:0] add_949325;
  wire [7:0] sel_949326;
  wire [7:0] add_949329;
  wire [7:0] sel_949330;
  wire [7:0] add_949333;
  wire [7:0] sel_949334;
  wire [7:0] add_949337;
  wire [7:0] sel_949338;
  wire [7:0] add_949341;
  wire [7:0] sel_949342;
  wire [7:0] add_949345;
  wire [7:0] sel_949346;
  wire [7:0] add_949349;
  wire [7:0] sel_949350;
  wire [7:0] add_949353;
  wire [7:0] sel_949354;
  wire [7:0] add_949357;
  wire [7:0] sel_949358;
  wire [7:0] add_949361;
  wire [7:0] sel_949362;
  wire [7:0] add_949365;
  wire [7:0] sel_949366;
  wire [7:0] add_949369;
  wire [7:0] sel_949370;
  wire [7:0] add_949373;
  wire [7:0] sel_949374;
  wire [7:0] add_949377;
  wire [7:0] sel_949378;
  wire [7:0] add_949381;
  wire [7:0] sel_949382;
  wire [7:0] add_949385;
  wire [7:0] sel_949386;
  wire [7:0] add_949389;
  wire [7:0] sel_949390;
  wire [7:0] add_949393;
  wire [7:0] sel_949394;
  wire [7:0] add_949397;
  wire [7:0] sel_949398;
  wire [7:0] add_949401;
  wire [7:0] sel_949402;
  wire [7:0] add_949405;
  wire [7:0] sel_949406;
  wire [7:0] add_949409;
  wire [7:0] sel_949410;
  wire [7:0] add_949413;
  wire [7:0] sel_949414;
  wire [7:0] add_949417;
  wire [7:0] sel_949418;
  wire [7:0] add_949421;
  wire [7:0] sel_949422;
  wire [7:0] add_949425;
  wire [7:0] sel_949426;
  wire [7:0] add_949429;
  wire [7:0] sel_949430;
  wire [7:0] add_949433;
  wire [7:0] sel_949434;
  wire [7:0] add_949437;
  wire [7:0] sel_949438;
  wire [7:0] add_949441;
  wire [7:0] sel_949442;
  wire [7:0] add_949445;
  wire [7:0] sel_949446;
  wire [7:0] add_949449;
  wire [7:0] sel_949450;
  wire [7:0] add_949453;
  wire [7:0] sel_949454;
  wire [7:0] add_949457;
  wire [7:0] sel_949458;
  wire [7:0] add_949461;
  wire [7:0] sel_949462;
  wire [7:0] add_949465;
  wire [7:0] sel_949466;
  wire [7:0] add_949469;
  wire [7:0] sel_949470;
  wire [7:0] add_949473;
  wire [7:0] sel_949474;
  wire [7:0] add_949477;
  wire [7:0] sel_949478;
  wire [7:0] add_949481;
  wire [7:0] sel_949482;
  wire [7:0] add_949485;
  wire [7:0] sel_949486;
  wire [7:0] add_949489;
  wire [7:0] sel_949490;
  wire [7:0] add_949494;
  wire [15:0] array_index_949495;
  wire [7:0] sel_949496;
  wire [7:0] add_949499;
  wire [7:0] sel_949500;
  wire [7:0] add_949503;
  wire [7:0] sel_949504;
  wire [7:0] add_949507;
  wire [7:0] sel_949508;
  wire [7:0] add_949511;
  wire [7:0] sel_949512;
  wire [7:0] add_949515;
  wire [7:0] sel_949516;
  wire [7:0] add_949519;
  wire [7:0] sel_949520;
  wire [7:0] add_949523;
  wire [7:0] sel_949524;
  wire [7:0] add_949527;
  wire [7:0] sel_949528;
  wire [7:0] add_949531;
  wire [7:0] sel_949532;
  wire [7:0] add_949535;
  wire [7:0] sel_949536;
  wire [7:0] add_949539;
  wire [7:0] sel_949540;
  wire [7:0] add_949543;
  wire [7:0] sel_949544;
  wire [7:0] add_949547;
  wire [7:0] sel_949548;
  wire [7:0] add_949551;
  wire [7:0] sel_949552;
  wire [7:0] add_949555;
  wire [7:0] sel_949556;
  wire [7:0] add_949559;
  wire [7:0] sel_949560;
  wire [7:0] add_949563;
  wire [7:0] sel_949564;
  wire [7:0] add_949567;
  wire [7:0] sel_949568;
  wire [7:0] add_949571;
  wire [7:0] sel_949572;
  wire [7:0] add_949575;
  wire [7:0] sel_949576;
  wire [7:0] add_949579;
  wire [7:0] sel_949580;
  wire [7:0] add_949583;
  wire [7:0] sel_949584;
  wire [7:0] add_949587;
  wire [7:0] sel_949588;
  wire [7:0] add_949591;
  wire [7:0] sel_949592;
  wire [7:0] add_949595;
  wire [7:0] sel_949596;
  wire [7:0] add_949599;
  wire [7:0] sel_949600;
  wire [7:0] add_949603;
  wire [7:0] sel_949604;
  wire [7:0] add_949607;
  wire [7:0] sel_949608;
  wire [7:0] add_949611;
  wire [7:0] sel_949612;
  wire [7:0] add_949615;
  wire [7:0] sel_949616;
  wire [7:0] add_949619;
  wire [7:0] sel_949620;
  wire [7:0] add_949623;
  wire [7:0] sel_949624;
  wire [7:0] add_949627;
  wire [7:0] sel_949628;
  wire [7:0] add_949631;
  wire [7:0] sel_949632;
  wire [7:0] add_949635;
  wire [7:0] sel_949636;
  wire [7:0] add_949639;
  wire [7:0] sel_949640;
  wire [7:0] add_949643;
  wire [7:0] sel_949644;
  wire [7:0] add_949647;
  wire [7:0] sel_949648;
  wire [7:0] add_949651;
  wire [7:0] sel_949652;
  wire [7:0] add_949655;
  wire [7:0] sel_949656;
  wire [7:0] add_949659;
  wire [7:0] sel_949660;
  wire [7:0] add_949663;
  wire [7:0] sel_949664;
  wire [7:0] add_949667;
  wire [7:0] sel_949668;
  wire [7:0] add_949671;
  wire [7:0] sel_949672;
  wire [7:0] add_949675;
  wire [7:0] sel_949676;
  wire [7:0] add_949679;
  wire [7:0] sel_949680;
  wire [7:0] add_949683;
  wire [7:0] sel_949684;
  wire [7:0] add_949687;
  wire [7:0] sel_949688;
  wire [7:0] add_949691;
  wire [7:0] sel_949692;
  wire [7:0] add_949695;
  wire [7:0] sel_949696;
  wire [7:0] add_949699;
  wire [7:0] sel_949700;
  wire [7:0] add_949703;
  wire [7:0] sel_949704;
  wire [7:0] add_949707;
  wire [7:0] sel_949708;
  wire [7:0] add_949711;
  wire [7:0] sel_949712;
  wire [7:0] add_949715;
  wire [7:0] sel_949716;
  wire [7:0] add_949719;
  wire [7:0] sel_949720;
  wire [7:0] add_949723;
  wire [7:0] sel_949724;
  wire [7:0] add_949727;
  wire [7:0] sel_949728;
  wire [7:0] add_949731;
  wire [7:0] sel_949732;
  wire [7:0] add_949735;
  wire [7:0] sel_949736;
  wire [7:0] add_949739;
  wire [7:0] sel_949740;
  wire [7:0] add_949743;
  wire [7:0] sel_949744;
  wire [7:0] add_949747;
  wire [7:0] sel_949748;
  wire [7:0] add_949751;
  wire [7:0] sel_949752;
  wire [7:0] add_949755;
  wire [7:0] sel_949756;
  wire [7:0] add_949759;
  wire [7:0] sel_949760;
  wire [7:0] add_949763;
  wire [7:0] sel_949764;
  wire [7:0] add_949767;
  wire [7:0] sel_949768;
  wire [7:0] add_949771;
  wire [7:0] sel_949772;
  wire [7:0] add_949775;
  wire [7:0] sel_949776;
  wire [7:0] add_949779;
  wire [7:0] sel_949780;
  wire [7:0] add_949783;
  wire [7:0] sel_949784;
  wire [7:0] add_949787;
  wire [7:0] sel_949788;
  wire [7:0] add_949791;
  wire [7:0] sel_949792;
  wire [7:0] add_949795;
  wire [7:0] sel_949796;
  wire [7:0] add_949799;
  wire [7:0] sel_949800;
  wire [7:0] add_949803;
  wire [7:0] sel_949804;
  wire [7:0] add_949807;
  wire [7:0] sel_949808;
  wire [7:0] add_949811;
  wire [7:0] sel_949812;
  wire [7:0] add_949815;
  wire [7:0] sel_949816;
  wire [7:0] add_949819;
  wire [7:0] sel_949820;
  wire [7:0] add_949823;
  wire [7:0] sel_949824;
  wire [7:0] add_949827;
  wire [7:0] sel_949828;
  wire [7:0] add_949831;
  wire [7:0] sel_949832;
  wire [7:0] add_949835;
  wire [7:0] sel_949836;
  wire [7:0] add_949839;
  wire [7:0] sel_949840;
  wire [7:0] add_949843;
  wire [7:0] sel_949844;
  wire [7:0] add_949847;
  wire [7:0] sel_949848;
  wire [7:0] add_949851;
  wire [7:0] sel_949852;
  wire [7:0] add_949855;
  wire [7:0] sel_949856;
  wire [7:0] add_949859;
  wire [7:0] sel_949860;
  wire [7:0] add_949863;
  wire [7:0] sel_949864;
  wire [7:0] add_949867;
  wire [7:0] sel_949868;
  wire [7:0] add_949871;
  wire [7:0] sel_949872;
  wire [7:0] add_949875;
  wire [7:0] sel_949876;
  wire [7:0] add_949879;
  wire [7:0] sel_949880;
  wire [7:0] add_949883;
  wire [7:0] sel_949884;
  wire [7:0] add_949887;
  wire [7:0] sel_949888;
  wire [7:0] add_949891;
  wire [7:0] sel_949892;
  wire [7:0] add_949896;
  wire [15:0] array_index_949897;
  wire [7:0] sel_949898;
  wire [7:0] add_949901;
  wire [7:0] sel_949902;
  wire [7:0] add_949905;
  wire [7:0] sel_949906;
  wire [7:0] add_949909;
  wire [7:0] sel_949910;
  wire [7:0] add_949913;
  wire [7:0] sel_949914;
  wire [7:0] add_949917;
  wire [7:0] sel_949918;
  wire [7:0] add_949921;
  wire [7:0] sel_949922;
  wire [7:0] add_949925;
  wire [7:0] sel_949926;
  wire [7:0] add_949929;
  wire [7:0] sel_949930;
  wire [7:0] add_949933;
  wire [7:0] sel_949934;
  wire [7:0] add_949937;
  wire [7:0] sel_949938;
  wire [7:0] add_949941;
  wire [7:0] sel_949942;
  wire [7:0] add_949945;
  wire [7:0] sel_949946;
  wire [7:0] add_949949;
  wire [7:0] sel_949950;
  wire [7:0] add_949953;
  wire [7:0] sel_949954;
  wire [7:0] add_949957;
  wire [7:0] sel_949958;
  wire [7:0] add_949961;
  wire [7:0] sel_949962;
  wire [7:0] add_949965;
  wire [7:0] sel_949966;
  wire [7:0] add_949969;
  wire [7:0] sel_949970;
  wire [7:0] add_949973;
  wire [7:0] sel_949974;
  wire [7:0] add_949977;
  wire [7:0] sel_949978;
  wire [7:0] add_949981;
  wire [7:0] sel_949982;
  wire [7:0] add_949985;
  wire [7:0] sel_949986;
  wire [7:0] add_949989;
  wire [7:0] sel_949990;
  wire [7:0] add_949993;
  wire [7:0] sel_949994;
  wire [7:0] add_949997;
  wire [7:0] sel_949998;
  wire [7:0] add_950001;
  wire [7:0] sel_950002;
  wire [7:0] add_950005;
  wire [7:0] sel_950006;
  wire [7:0] add_950009;
  wire [7:0] sel_950010;
  wire [7:0] add_950013;
  wire [7:0] sel_950014;
  wire [7:0] add_950017;
  wire [7:0] sel_950018;
  wire [7:0] add_950021;
  wire [7:0] sel_950022;
  wire [7:0] add_950025;
  wire [7:0] sel_950026;
  wire [7:0] add_950029;
  wire [7:0] sel_950030;
  wire [7:0] add_950033;
  wire [7:0] sel_950034;
  wire [7:0] add_950037;
  wire [7:0] sel_950038;
  wire [7:0] add_950041;
  wire [7:0] sel_950042;
  wire [7:0] add_950045;
  wire [7:0] sel_950046;
  wire [7:0] add_950049;
  wire [7:0] sel_950050;
  wire [7:0] add_950053;
  wire [7:0] sel_950054;
  wire [7:0] add_950057;
  wire [7:0] sel_950058;
  wire [7:0] add_950061;
  wire [7:0] sel_950062;
  wire [7:0] add_950065;
  wire [7:0] sel_950066;
  wire [7:0] add_950069;
  wire [7:0] sel_950070;
  wire [7:0] add_950073;
  wire [7:0] sel_950074;
  wire [7:0] add_950077;
  wire [7:0] sel_950078;
  wire [7:0] add_950081;
  wire [7:0] sel_950082;
  wire [7:0] add_950085;
  wire [7:0] sel_950086;
  wire [7:0] add_950089;
  wire [7:0] sel_950090;
  wire [7:0] add_950093;
  wire [7:0] sel_950094;
  wire [7:0] add_950097;
  wire [7:0] sel_950098;
  wire [7:0] add_950101;
  wire [7:0] sel_950102;
  wire [7:0] add_950105;
  wire [7:0] sel_950106;
  wire [7:0] add_950109;
  wire [7:0] sel_950110;
  wire [7:0] add_950113;
  wire [7:0] sel_950114;
  wire [7:0] add_950117;
  wire [7:0] sel_950118;
  wire [7:0] add_950121;
  wire [7:0] sel_950122;
  wire [7:0] add_950125;
  wire [7:0] sel_950126;
  wire [7:0] add_950129;
  wire [7:0] sel_950130;
  wire [7:0] add_950133;
  wire [7:0] sel_950134;
  wire [7:0] add_950137;
  wire [7:0] sel_950138;
  wire [7:0] add_950141;
  wire [7:0] sel_950142;
  wire [7:0] add_950145;
  wire [7:0] sel_950146;
  wire [7:0] add_950149;
  wire [7:0] sel_950150;
  wire [7:0] add_950153;
  wire [7:0] sel_950154;
  wire [7:0] add_950157;
  wire [7:0] sel_950158;
  wire [7:0] add_950161;
  wire [7:0] sel_950162;
  wire [7:0] add_950165;
  wire [7:0] sel_950166;
  wire [7:0] add_950169;
  wire [7:0] sel_950170;
  wire [7:0] add_950173;
  wire [7:0] sel_950174;
  wire [7:0] add_950177;
  wire [7:0] sel_950178;
  wire [7:0] add_950181;
  wire [7:0] sel_950182;
  wire [7:0] add_950185;
  wire [7:0] sel_950186;
  wire [7:0] add_950189;
  wire [7:0] sel_950190;
  wire [7:0] add_950193;
  wire [7:0] sel_950194;
  wire [7:0] add_950197;
  wire [7:0] sel_950198;
  wire [7:0] add_950201;
  wire [7:0] sel_950202;
  wire [7:0] add_950205;
  wire [7:0] sel_950206;
  wire [7:0] add_950209;
  wire [7:0] sel_950210;
  wire [7:0] add_950213;
  wire [7:0] sel_950214;
  wire [7:0] add_950217;
  wire [7:0] sel_950218;
  wire [7:0] add_950221;
  wire [7:0] sel_950222;
  wire [7:0] add_950225;
  wire [7:0] sel_950226;
  wire [7:0] add_950229;
  wire [7:0] sel_950230;
  wire [7:0] add_950233;
  wire [7:0] sel_950234;
  wire [7:0] add_950237;
  wire [7:0] sel_950238;
  wire [7:0] add_950241;
  wire [7:0] sel_950242;
  wire [7:0] add_950245;
  wire [7:0] sel_950246;
  wire [7:0] add_950249;
  wire [7:0] sel_950250;
  wire [7:0] add_950253;
  wire [7:0] sel_950254;
  wire [7:0] add_950257;
  wire [7:0] sel_950258;
  wire [7:0] add_950261;
  wire [7:0] sel_950262;
  wire [7:0] add_950265;
  wire [7:0] sel_950266;
  wire [7:0] add_950269;
  wire [7:0] sel_950270;
  wire [7:0] add_950273;
  wire [7:0] sel_950274;
  wire [7:0] add_950277;
  wire [7:0] sel_950278;
  wire [7:0] add_950281;
  wire [7:0] sel_950282;
  wire [7:0] add_950285;
  wire [7:0] sel_950286;
  wire [7:0] add_950289;
  wire [7:0] sel_950290;
  wire [7:0] add_950293;
  wire [7:0] sel_950294;
  wire [7:0] add_950298;
  wire [15:0] array_index_950299;
  wire [7:0] sel_950300;
  wire [7:0] add_950303;
  wire [7:0] sel_950304;
  wire [7:0] add_950307;
  wire [7:0] sel_950308;
  wire [7:0] add_950311;
  wire [7:0] sel_950312;
  wire [7:0] add_950315;
  wire [7:0] sel_950316;
  wire [7:0] add_950319;
  wire [7:0] sel_950320;
  wire [7:0] add_950323;
  wire [7:0] sel_950324;
  wire [7:0] add_950327;
  wire [7:0] sel_950328;
  wire [7:0] add_950331;
  wire [7:0] sel_950332;
  wire [7:0] add_950335;
  wire [7:0] sel_950336;
  wire [7:0] add_950339;
  wire [7:0] sel_950340;
  wire [7:0] add_950343;
  wire [7:0] sel_950344;
  wire [7:0] add_950347;
  wire [7:0] sel_950348;
  wire [7:0] add_950351;
  wire [7:0] sel_950352;
  wire [7:0] add_950355;
  wire [7:0] sel_950356;
  wire [7:0] add_950359;
  wire [7:0] sel_950360;
  wire [7:0] add_950363;
  wire [7:0] sel_950364;
  wire [7:0] add_950367;
  wire [7:0] sel_950368;
  wire [7:0] add_950371;
  wire [7:0] sel_950372;
  wire [7:0] add_950375;
  wire [7:0] sel_950376;
  wire [7:0] add_950379;
  wire [7:0] sel_950380;
  wire [7:0] add_950383;
  wire [7:0] sel_950384;
  wire [7:0] add_950387;
  wire [7:0] sel_950388;
  wire [7:0] add_950391;
  wire [7:0] sel_950392;
  wire [7:0] add_950395;
  wire [7:0] sel_950396;
  wire [7:0] add_950399;
  wire [7:0] sel_950400;
  wire [7:0] add_950403;
  wire [7:0] sel_950404;
  wire [7:0] add_950407;
  wire [7:0] sel_950408;
  wire [7:0] add_950411;
  wire [7:0] sel_950412;
  wire [7:0] add_950415;
  wire [7:0] sel_950416;
  wire [7:0] add_950419;
  wire [7:0] sel_950420;
  wire [7:0] add_950423;
  wire [7:0] sel_950424;
  wire [7:0] add_950427;
  wire [7:0] sel_950428;
  wire [7:0] add_950431;
  wire [7:0] sel_950432;
  wire [7:0] add_950435;
  wire [7:0] sel_950436;
  wire [7:0] add_950439;
  wire [7:0] sel_950440;
  wire [7:0] add_950443;
  wire [7:0] sel_950444;
  wire [7:0] add_950447;
  wire [7:0] sel_950448;
  wire [7:0] add_950451;
  wire [7:0] sel_950452;
  wire [7:0] add_950455;
  wire [7:0] sel_950456;
  wire [7:0] add_950459;
  wire [7:0] sel_950460;
  wire [7:0] add_950463;
  wire [7:0] sel_950464;
  wire [7:0] add_950467;
  wire [7:0] sel_950468;
  wire [7:0] add_950471;
  wire [7:0] sel_950472;
  wire [7:0] add_950475;
  wire [7:0] sel_950476;
  wire [7:0] add_950479;
  wire [7:0] sel_950480;
  wire [7:0] add_950483;
  wire [7:0] sel_950484;
  wire [7:0] add_950487;
  wire [7:0] sel_950488;
  wire [7:0] add_950491;
  wire [7:0] sel_950492;
  wire [7:0] add_950495;
  wire [7:0] sel_950496;
  wire [7:0] add_950499;
  wire [7:0] sel_950500;
  wire [7:0] add_950503;
  wire [7:0] sel_950504;
  wire [7:0] add_950507;
  wire [7:0] sel_950508;
  wire [7:0] add_950511;
  wire [7:0] sel_950512;
  wire [7:0] add_950515;
  wire [7:0] sel_950516;
  wire [7:0] add_950519;
  wire [7:0] sel_950520;
  wire [7:0] add_950523;
  wire [7:0] sel_950524;
  wire [7:0] add_950527;
  wire [7:0] sel_950528;
  wire [7:0] add_950531;
  wire [7:0] sel_950532;
  wire [7:0] add_950535;
  wire [7:0] sel_950536;
  wire [7:0] add_950539;
  wire [7:0] sel_950540;
  wire [7:0] add_950543;
  wire [7:0] sel_950544;
  wire [7:0] add_950547;
  wire [7:0] sel_950548;
  wire [7:0] add_950551;
  wire [7:0] sel_950552;
  wire [7:0] add_950555;
  wire [7:0] sel_950556;
  wire [7:0] add_950559;
  wire [7:0] sel_950560;
  wire [7:0] add_950563;
  wire [7:0] sel_950564;
  wire [7:0] add_950567;
  wire [7:0] sel_950568;
  wire [7:0] add_950571;
  wire [7:0] sel_950572;
  wire [7:0] add_950575;
  wire [7:0] sel_950576;
  wire [7:0] add_950579;
  wire [7:0] sel_950580;
  wire [7:0] add_950583;
  wire [7:0] sel_950584;
  wire [7:0] add_950587;
  wire [7:0] sel_950588;
  wire [7:0] add_950591;
  wire [7:0] sel_950592;
  wire [7:0] add_950595;
  wire [7:0] sel_950596;
  wire [7:0] add_950599;
  wire [7:0] sel_950600;
  wire [7:0] add_950603;
  wire [7:0] sel_950604;
  wire [7:0] add_950607;
  wire [7:0] sel_950608;
  wire [7:0] add_950611;
  wire [7:0] sel_950612;
  wire [7:0] add_950615;
  wire [7:0] sel_950616;
  wire [7:0] add_950619;
  wire [7:0] sel_950620;
  wire [7:0] add_950623;
  wire [7:0] sel_950624;
  wire [7:0] add_950627;
  wire [7:0] sel_950628;
  wire [7:0] add_950631;
  wire [7:0] sel_950632;
  wire [7:0] add_950635;
  wire [7:0] sel_950636;
  wire [7:0] add_950639;
  wire [7:0] sel_950640;
  wire [7:0] add_950643;
  wire [7:0] sel_950644;
  wire [7:0] add_950647;
  wire [7:0] sel_950648;
  wire [7:0] add_950651;
  wire [7:0] sel_950652;
  wire [7:0] add_950655;
  wire [7:0] sel_950656;
  wire [7:0] add_950659;
  wire [7:0] sel_950660;
  wire [7:0] add_950663;
  wire [7:0] sel_950664;
  wire [7:0] add_950667;
  wire [7:0] sel_950668;
  wire [7:0] add_950671;
  wire [7:0] sel_950672;
  wire [7:0] add_950675;
  wire [7:0] sel_950676;
  wire [7:0] add_950679;
  wire [7:0] sel_950680;
  wire [7:0] add_950683;
  wire [7:0] sel_950684;
  wire [7:0] add_950687;
  wire [7:0] sel_950688;
  wire [7:0] add_950691;
  wire [7:0] sel_950692;
  wire [7:0] add_950695;
  wire [7:0] sel_950696;
  wire [7:0] add_950700;
  wire [15:0] array_index_950701;
  wire [7:0] sel_950702;
  wire [7:0] add_950705;
  wire [7:0] sel_950706;
  wire [7:0] add_950709;
  wire [7:0] sel_950710;
  wire [7:0] add_950713;
  wire [7:0] sel_950714;
  wire [7:0] add_950717;
  wire [7:0] sel_950718;
  wire [7:0] add_950721;
  wire [7:0] sel_950722;
  wire [7:0] add_950725;
  wire [7:0] sel_950726;
  wire [7:0] add_950729;
  wire [7:0] sel_950730;
  wire [7:0] add_950733;
  wire [7:0] sel_950734;
  wire [7:0] add_950737;
  wire [7:0] sel_950738;
  wire [7:0] add_950741;
  wire [7:0] sel_950742;
  wire [7:0] add_950745;
  wire [7:0] sel_950746;
  wire [7:0] add_950749;
  wire [7:0] sel_950750;
  wire [7:0] add_950753;
  wire [7:0] sel_950754;
  wire [7:0] add_950757;
  wire [7:0] sel_950758;
  wire [7:0] add_950761;
  wire [7:0] sel_950762;
  wire [7:0] add_950765;
  wire [7:0] sel_950766;
  wire [7:0] add_950769;
  wire [7:0] sel_950770;
  wire [7:0] add_950773;
  wire [7:0] sel_950774;
  wire [7:0] add_950777;
  wire [7:0] sel_950778;
  wire [7:0] add_950781;
  wire [7:0] sel_950782;
  wire [7:0] add_950785;
  wire [7:0] sel_950786;
  wire [7:0] add_950789;
  wire [7:0] sel_950790;
  wire [7:0] add_950793;
  wire [7:0] sel_950794;
  wire [7:0] add_950797;
  wire [7:0] sel_950798;
  wire [7:0] add_950801;
  wire [7:0] sel_950802;
  wire [7:0] add_950805;
  wire [7:0] sel_950806;
  wire [7:0] add_950809;
  wire [7:0] sel_950810;
  wire [7:0] add_950813;
  wire [7:0] sel_950814;
  wire [7:0] add_950817;
  wire [7:0] sel_950818;
  wire [7:0] add_950821;
  wire [7:0] sel_950822;
  wire [7:0] add_950825;
  wire [7:0] sel_950826;
  wire [7:0] add_950829;
  wire [7:0] sel_950830;
  wire [7:0] add_950833;
  wire [7:0] sel_950834;
  wire [7:0] add_950837;
  wire [7:0] sel_950838;
  wire [7:0] add_950841;
  wire [7:0] sel_950842;
  wire [7:0] add_950845;
  wire [7:0] sel_950846;
  wire [7:0] add_950849;
  wire [7:0] sel_950850;
  wire [7:0] add_950853;
  wire [7:0] sel_950854;
  wire [7:0] add_950857;
  wire [7:0] sel_950858;
  wire [7:0] add_950861;
  wire [7:0] sel_950862;
  wire [7:0] add_950865;
  wire [7:0] sel_950866;
  wire [7:0] add_950869;
  wire [7:0] sel_950870;
  wire [7:0] add_950873;
  wire [7:0] sel_950874;
  wire [7:0] add_950877;
  wire [7:0] sel_950878;
  wire [7:0] add_950881;
  wire [7:0] sel_950882;
  wire [7:0] add_950885;
  wire [7:0] sel_950886;
  wire [7:0] add_950889;
  wire [7:0] sel_950890;
  wire [7:0] add_950893;
  wire [7:0] sel_950894;
  wire [7:0] add_950897;
  wire [7:0] sel_950898;
  wire [7:0] add_950901;
  wire [7:0] sel_950902;
  wire [7:0] add_950905;
  wire [7:0] sel_950906;
  wire [7:0] add_950909;
  wire [7:0] sel_950910;
  wire [7:0] add_950913;
  wire [7:0] sel_950914;
  wire [7:0] add_950917;
  wire [7:0] sel_950918;
  wire [7:0] add_950921;
  wire [7:0] sel_950922;
  wire [7:0] add_950925;
  wire [7:0] sel_950926;
  wire [7:0] add_950929;
  wire [7:0] sel_950930;
  wire [7:0] add_950933;
  wire [7:0] sel_950934;
  wire [7:0] add_950937;
  wire [7:0] sel_950938;
  wire [7:0] add_950941;
  wire [7:0] sel_950942;
  wire [7:0] add_950945;
  wire [7:0] sel_950946;
  wire [7:0] add_950949;
  wire [7:0] sel_950950;
  wire [7:0] add_950953;
  wire [7:0] sel_950954;
  wire [7:0] add_950957;
  wire [7:0] sel_950958;
  wire [7:0] add_950961;
  wire [7:0] sel_950962;
  wire [7:0] add_950965;
  wire [7:0] sel_950966;
  wire [7:0] add_950969;
  wire [7:0] sel_950970;
  wire [7:0] add_950973;
  wire [7:0] sel_950974;
  wire [7:0] add_950977;
  wire [7:0] sel_950978;
  wire [7:0] add_950981;
  wire [7:0] sel_950982;
  wire [7:0] add_950985;
  wire [7:0] sel_950986;
  wire [7:0] add_950989;
  wire [7:0] sel_950990;
  wire [7:0] add_950993;
  wire [7:0] sel_950994;
  wire [7:0] add_950997;
  wire [7:0] sel_950998;
  wire [7:0] add_951001;
  wire [7:0] sel_951002;
  wire [7:0] add_951005;
  wire [7:0] sel_951006;
  wire [7:0] add_951009;
  wire [7:0] sel_951010;
  wire [7:0] add_951013;
  wire [7:0] sel_951014;
  wire [7:0] add_951017;
  wire [7:0] sel_951018;
  wire [7:0] add_951021;
  wire [7:0] sel_951022;
  wire [7:0] add_951025;
  wire [7:0] sel_951026;
  wire [7:0] add_951029;
  wire [7:0] sel_951030;
  wire [7:0] add_951033;
  wire [7:0] sel_951034;
  wire [7:0] add_951037;
  wire [7:0] sel_951038;
  wire [7:0] add_951041;
  wire [7:0] sel_951042;
  wire [7:0] add_951045;
  wire [7:0] sel_951046;
  wire [7:0] add_951049;
  wire [7:0] sel_951050;
  wire [7:0] add_951053;
  wire [7:0] sel_951054;
  wire [7:0] add_951057;
  wire [7:0] sel_951058;
  wire [7:0] add_951061;
  wire [7:0] sel_951062;
  wire [7:0] add_951065;
  wire [7:0] sel_951066;
  wire [7:0] add_951069;
  wire [7:0] sel_951070;
  wire [7:0] add_951073;
  wire [7:0] sel_951074;
  wire [7:0] add_951077;
  wire [7:0] sel_951078;
  wire [7:0] add_951081;
  wire [7:0] sel_951082;
  wire [7:0] add_951085;
  wire [7:0] sel_951086;
  wire [7:0] add_951089;
  wire [7:0] sel_951090;
  wire [7:0] add_951093;
  wire [7:0] sel_951094;
  wire [7:0] add_951097;
  wire [7:0] sel_951098;
  wire [7:0] add_951102;
  wire [15:0] array_index_951103;
  wire [7:0] sel_951104;
  wire [7:0] add_951107;
  wire [7:0] sel_951108;
  wire [7:0] add_951111;
  wire [7:0] sel_951112;
  wire [7:0] add_951115;
  wire [7:0] sel_951116;
  wire [7:0] add_951119;
  wire [7:0] sel_951120;
  wire [7:0] add_951123;
  wire [7:0] sel_951124;
  wire [7:0] add_951127;
  wire [7:0] sel_951128;
  wire [7:0] add_951131;
  wire [7:0] sel_951132;
  wire [7:0] add_951135;
  wire [7:0] sel_951136;
  wire [7:0] add_951139;
  wire [7:0] sel_951140;
  wire [7:0] add_951143;
  wire [7:0] sel_951144;
  wire [7:0] add_951147;
  wire [7:0] sel_951148;
  wire [7:0] add_951151;
  wire [7:0] sel_951152;
  wire [7:0] add_951155;
  wire [7:0] sel_951156;
  wire [7:0] add_951159;
  wire [7:0] sel_951160;
  wire [7:0] add_951163;
  wire [7:0] sel_951164;
  wire [7:0] add_951167;
  wire [7:0] sel_951168;
  wire [7:0] add_951171;
  wire [7:0] sel_951172;
  wire [7:0] add_951175;
  wire [7:0] sel_951176;
  wire [7:0] add_951179;
  wire [7:0] sel_951180;
  wire [7:0] add_951183;
  wire [7:0] sel_951184;
  wire [7:0] add_951187;
  wire [7:0] sel_951188;
  wire [7:0] add_951191;
  wire [7:0] sel_951192;
  wire [7:0] add_951195;
  wire [7:0] sel_951196;
  wire [7:0] add_951199;
  wire [7:0] sel_951200;
  wire [7:0] add_951203;
  wire [7:0] sel_951204;
  wire [7:0] add_951207;
  wire [7:0] sel_951208;
  wire [7:0] add_951211;
  wire [7:0] sel_951212;
  wire [7:0] add_951215;
  wire [7:0] sel_951216;
  wire [7:0] add_951219;
  wire [7:0] sel_951220;
  wire [7:0] add_951223;
  wire [7:0] sel_951224;
  wire [7:0] add_951227;
  wire [7:0] sel_951228;
  wire [7:0] add_951231;
  wire [7:0] sel_951232;
  wire [7:0] add_951235;
  wire [7:0] sel_951236;
  wire [7:0] add_951239;
  wire [7:0] sel_951240;
  wire [7:0] add_951243;
  wire [7:0] sel_951244;
  wire [7:0] add_951247;
  wire [7:0] sel_951248;
  wire [7:0] add_951251;
  wire [7:0] sel_951252;
  wire [7:0] add_951255;
  wire [7:0] sel_951256;
  wire [7:0] add_951259;
  wire [7:0] sel_951260;
  wire [7:0] add_951263;
  wire [7:0] sel_951264;
  wire [7:0] add_951267;
  wire [7:0] sel_951268;
  wire [7:0] add_951271;
  wire [7:0] sel_951272;
  wire [7:0] add_951275;
  wire [7:0] sel_951276;
  wire [7:0] add_951279;
  wire [7:0] sel_951280;
  wire [7:0] add_951283;
  wire [7:0] sel_951284;
  wire [7:0] add_951287;
  wire [7:0] sel_951288;
  wire [7:0] add_951291;
  wire [7:0] sel_951292;
  wire [7:0] add_951295;
  wire [7:0] sel_951296;
  wire [7:0] add_951299;
  wire [7:0] sel_951300;
  wire [7:0] add_951303;
  wire [7:0] sel_951304;
  wire [7:0] add_951307;
  wire [7:0] sel_951308;
  wire [7:0] add_951311;
  wire [7:0] sel_951312;
  wire [7:0] add_951315;
  wire [7:0] sel_951316;
  wire [7:0] add_951319;
  wire [7:0] sel_951320;
  wire [7:0] add_951323;
  wire [7:0] sel_951324;
  wire [7:0] add_951327;
  wire [7:0] sel_951328;
  wire [7:0] add_951331;
  wire [7:0] sel_951332;
  wire [7:0] add_951335;
  wire [7:0] sel_951336;
  wire [7:0] add_951339;
  wire [7:0] sel_951340;
  wire [7:0] add_951343;
  wire [7:0] sel_951344;
  wire [7:0] add_951347;
  wire [7:0] sel_951348;
  wire [7:0] add_951351;
  wire [7:0] sel_951352;
  wire [7:0] add_951355;
  wire [7:0] sel_951356;
  wire [7:0] add_951359;
  wire [7:0] sel_951360;
  wire [7:0] add_951363;
  wire [7:0] sel_951364;
  wire [7:0] add_951367;
  wire [7:0] sel_951368;
  wire [7:0] add_951371;
  wire [7:0] sel_951372;
  wire [7:0] add_951375;
  wire [7:0] sel_951376;
  wire [7:0] add_951379;
  wire [7:0] sel_951380;
  wire [7:0] add_951383;
  wire [7:0] sel_951384;
  wire [7:0] add_951387;
  wire [7:0] sel_951388;
  wire [7:0] add_951391;
  wire [7:0] sel_951392;
  wire [7:0] add_951395;
  wire [7:0] sel_951396;
  wire [7:0] add_951399;
  wire [7:0] sel_951400;
  wire [7:0] add_951403;
  wire [7:0] sel_951404;
  wire [7:0] add_951407;
  wire [7:0] sel_951408;
  wire [7:0] add_951411;
  wire [7:0] sel_951412;
  wire [7:0] add_951415;
  wire [7:0] sel_951416;
  wire [7:0] add_951419;
  wire [7:0] sel_951420;
  wire [7:0] add_951423;
  wire [7:0] sel_951424;
  wire [7:0] add_951427;
  wire [7:0] sel_951428;
  wire [7:0] add_951431;
  wire [7:0] sel_951432;
  wire [7:0] add_951435;
  wire [7:0] sel_951436;
  wire [7:0] add_951439;
  wire [7:0] sel_951440;
  wire [7:0] add_951443;
  wire [7:0] sel_951444;
  wire [7:0] add_951447;
  wire [7:0] sel_951448;
  wire [7:0] add_951451;
  wire [7:0] sel_951452;
  wire [7:0] add_951455;
  wire [7:0] sel_951456;
  wire [7:0] add_951459;
  wire [7:0] sel_951460;
  wire [7:0] add_951463;
  wire [7:0] sel_951464;
  wire [7:0] add_951467;
  wire [7:0] sel_951468;
  wire [7:0] add_951471;
  wire [7:0] sel_951472;
  wire [7:0] add_951475;
  wire [7:0] sel_951476;
  wire [7:0] add_951479;
  wire [7:0] sel_951480;
  wire [7:0] add_951483;
  wire [7:0] sel_951484;
  wire [7:0] add_951487;
  wire [7:0] sel_951488;
  wire [7:0] add_951491;
  wire [7:0] sel_951492;
  wire [7:0] add_951495;
  wire [7:0] sel_951496;
  wire [7:0] add_951499;
  wire [7:0] sel_951500;
  wire [7:0] add_951504;
  wire [15:0] array_index_951505;
  wire [7:0] sel_951506;
  wire [7:0] add_951509;
  wire [7:0] sel_951510;
  wire [7:0] add_951513;
  wire [7:0] sel_951514;
  wire [7:0] add_951517;
  wire [7:0] sel_951518;
  wire [7:0] add_951521;
  wire [7:0] sel_951522;
  wire [7:0] add_951525;
  wire [7:0] sel_951526;
  wire [7:0] add_951529;
  wire [7:0] sel_951530;
  wire [7:0] add_951533;
  wire [7:0] sel_951534;
  wire [7:0] add_951537;
  wire [7:0] sel_951538;
  wire [7:0] add_951541;
  wire [7:0] sel_951542;
  wire [7:0] add_951545;
  wire [7:0] sel_951546;
  wire [7:0] add_951549;
  wire [7:0] sel_951550;
  wire [7:0] add_951553;
  wire [7:0] sel_951554;
  wire [7:0] add_951557;
  wire [7:0] sel_951558;
  wire [7:0] add_951561;
  wire [7:0] sel_951562;
  wire [7:0] add_951565;
  wire [7:0] sel_951566;
  wire [7:0] add_951569;
  wire [7:0] sel_951570;
  wire [7:0] add_951573;
  wire [7:0] sel_951574;
  wire [7:0] add_951577;
  wire [7:0] sel_951578;
  wire [7:0] add_951581;
  wire [7:0] sel_951582;
  wire [7:0] add_951585;
  wire [7:0] sel_951586;
  wire [7:0] add_951589;
  wire [7:0] sel_951590;
  wire [7:0] add_951593;
  wire [7:0] sel_951594;
  wire [7:0] add_951597;
  wire [7:0] sel_951598;
  wire [7:0] add_951601;
  wire [7:0] sel_951602;
  wire [7:0] add_951605;
  wire [7:0] sel_951606;
  wire [7:0] add_951609;
  wire [7:0] sel_951610;
  wire [7:0] add_951613;
  wire [7:0] sel_951614;
  wire [7:0] add_951617;
  wire [7:0] sel_951618;
  wire [7:0] add_951621;
  wire [7:0] sel_951622;
  wire [7:0] add_951625;
  wire [7:0] sel_951626;
  wire [7:0] add_951629;
  wire [7:0] sel_951630;
  wire [7:0] add_951633;
  wire [7:0] sel_951634;
  wire [7:0] add_951637;
  wire [7:0] sel_951638;
  wire [7:0] add_951641;
  wire [7:0] sel_951642;
  wire [7:0] add_951645;
  wire [7:0] sel_951646;
  wire [7:0] add_951649;
  wire [7:0] sel_951650;
  wire [7:0] add_951653;
  wire [7:0] sel_951654;
  wire [7:0] add_951657;
  wire [7:0] sel_951658;
  wire [7:0] add_951661;
  wire [7:0] sel_951662;
  wire [7:0] add_951665;
  wire [7:0] sel_951666;
  wire [7:0] add_951669;
  wire [7:0] sel_951670;
  wire [7:0] add_951673;
  wire [7:0] sel_951674;
  wire [7:0] add_951677;
  wire [7:0] sel_951678;
  wire [7:0] add_951681;
  wire [7:0] sel_951682;
  wire [7:0] add_951685;
  wire [7:0] sel_951686;
  wire [7:0] add_951689;
  wire [7:0] sel_951690;
  wire [7:0] add_951693;
  wire [7:0] sel_951694;
  wire [7:0] add_951697;
  wire [7:0] sel_951698;
  wire [7:0] add_951701;
  wire [7:0] sel_951702;
  wire [7:0] add_951705;
  wire [7:0] sel_951706;
  wire [7:0] add_951709;
  wire [7:0] sel_951710;
  wire [7:0] add_951713;
  wire [7:0] sel_951714;
  wire [7:0] add_951717;
  wire [7:0] sel_951718;
  wire [7:0] add_951721;
  wire [7:0] sel_951722;
  wire [7:0] add_951725;
  wire [7:0] sel_951726;
  wire [7:0] add_951729;
  wire [7:0] sel_951730;
  wire [7:0] add_951733;
  wire [7:0] sel_951734;
  wire [7:0] add_951737;
  wire [7:0] sel_951738;
  wire [7:0] add_951741;
  wire [7:0] sel_951742;
  wire [7:0] add_951745;
  wire [7:0] sel_951746;
  wire [7:0] add_951749;
  wire [7:0] sel_951750;
  wire [7:0] add_951753;
  wire [7:0] sel_951754;
  wire [7:0] add_951757;
  wire [7:0] sel_951758;
  wire [7:0] add_951761;
  wire [7:0] sel_951762;
  wire [7:0] add_951765;
  wire [7:0] sel_951766;
  wire [7:0] add_951769;
  wire [7:0] sel_951770;
  wire [7:0] add_951773;
  wire [7:0] sel_951774;
  wire [7:0] add_951777;
  wire [7:0] sel_951778;
  wire [7:0] add_951781;
  wire [7:0] sel_951782;
  wire [7:0] add_951785;
  wire [7:0] sel_951786;
  wire [7:0] add_951789;
  wire [7:0] sel_951790;
  wire [7:0] add_951793;
  wire [7:0] sel_951794;
  wire [7:0] add_951797;
  wire [7:0] sel_951798;
  wire [7:0] add_951801;
  wire [7:0] sel_951802;
  wire [7:0] add_951805;
  wire [7:0] sel_951806;
  wire [7:0] add_951809;
  wire [7:0] sel_951810;
  wire [7:0] add_951813;
  wire [7:0] sel_951814;
  wire [7:0] add_951817;
  wire [7:0] sel_951818;
  wire [7:0] add_951821;
  wire [7:0] sel_951822;
  wire [7:0] add_951825;
  wire [7:0] sel_951826;
  wire [7:0] add_951829;
  wire [7:0] sel_951830;
  wire [7:0] add_951833;
  wire [7:0] sel_951834;
  wire [7:0] add_951837;
  wire [7:0] sel_951838;
  wire [7:0] add_951841;
  wire [7:0] sel_951842;
  wire [7:0] add_951845;
  wire [7:0] sel_951846;
  wire [7:0] add_951849;
  wire [7:0] sel_951850;
  wire [7:0] add_951853;
  wire [7:0] sel_951854;
  wire [7:0] add_951857;
  wire [7:0] sel_951858;
  wire [7:0] add_951861;
  wire [7:0] sel_951862;
  wire [7:0] add_951865;
  wire [7:0] sel_951866;
  wire [7:0] add_951869;
  wire [7:0] sel_951870;
  wire [7:0] add_951873;
  wire [7:0] sel_951874;
  wire [7:0] add_951877;
  wire [7:0] sel_951878;
  wire [7:0] add_951881;
  wire [7:0] sel_951882;
  wire [7:0] add_951885;
  wire [7:0] sel_951886;
  wire [7:0] add_951889;
  wire [7:0] sel_951890;
  wire [7:0] add_951893;
  wire [7:0] sel_951894;
  wire [7:0] add_951897;
  wire [7:0] sel_951898;
  wire [7:0] add_951901;
  wire [7:0] sel_951902;
  wire [7:0] add_951906;
  wire [15:0] array_index_951907;
  wire [7:0] sel_951908;
  wire [7:0] add_951911;
  wire [7:0] sel_951912;
  wire [7:0] add_951915;
  wire [7:0] sel_951916;
  wire [7:0] add_951919;
  wire [7:0] sel_951920;
  wire [7:0] add_951923;
  wire [7:0] sel_951924;
  wire [7:0] add_951927;
  wire [7:0] sel_951928;
  wire [7:0] add_951931;
  wire [7:0] sel_951932;
  wire [7:0] add_951935;
  wire [7:0] sel_951936;
  wire [7:0] add_951939;
  wire [7:0] sel_951940;
  wire [7:0] add_951943;
  wire [7:0] sel_951944;
  wire [7:0] add_951947;
  wire [7:0] sel_951948;
  wire [7:0] add_951951;
  wire [7:0] sel_951952;
  wire [7:0] add_951955;
  wire [7:0] sel_951956;
  wire [7:0] add_951959;
  wire [7:0] sel_951960;
  wire [7:0] add_951963;
  wire [7:0] sel_951964;
  wire [7:0] add_951967;
  wire [7:0] sel_951968;
  wire [7:0] add_951971;
  wire [7:0] sel_951972;
  wire [7:0] add_951975;
  wire [7:0] sel_951976;
  wire [7:0] add_951979;
  wire [7:0] sel_951980;
  wire [7:0] add_951983;
  wire [7:0] sel_951984;
  wire [7:0] add_951987;
  wire [7:0] sel_951988;
  wire [7:0] add_951991;
  wire [7:0] sel_951992;
  wire [7:0] add_951995;
  wire [7:0] sel_951996;
  wire [7:0] add_951999;
  wire [7:0] sel_952000;
  wire [7:0] add_952003;
  wire [7:0] sel_952004;
  wire [7:0] add_952007;
  wire [7:0] sel_952008;
  wire [7:0] add_952011;
  wire [7:0] sel_952012;
  wire [7:0] add_952015;
  wire [7:0] sel_952016;
  wire [7:0] add_952019;
  wire [7:0] sel_952020;
  wire [7:0] add_952023;
  wire [7:0] sel_952024;
  wire [7:0] add_952027;
  wire [7:0] sel_952028;
  wire [7:0] add_952031;
  wire [7:0] sel_952032;
  wire [7:0] add_952035;
  wire [7:0] sel_952036;
  wire [7:0] add_952039;
  wire [7:0] sel_952040;
  wire [7:0] add_952043;
  wire [7:0] sel_952044;
  wire [7:0] add_952047;
  wire [7:0] sel_952048;
  wire [7:0] add_952051;
  wire [7:0] sel_952052;
  wire [7:0] add_952055;
  wire [7:0] sel_952056;
  wire [7:0] add_952059;
  wire [7:0] sel_952060;
  wire [7:0] add_952063;
  wire [7:0] sel_952064;
  wire [7:0] add_952067;
  wire [7:0] sel_952068;
  wire [7:0] add_952071;
  wire [7:0] sel_952072;
  wire [7:0] add_952075;
  wire [7:0] sel_952076;
  wire [7:0] add_952079;
  wire [7:0] sel_952080;
  wire [7:0] add_952083;
  wire [7:0] sel_952084;
  wire [7:0] add_952087;
  wire [7:0] sel_952088;
  wire [7:0] add_952091;
  wire [7:0] sel_952092;
  wire [7:0] add_952095;
  wire [7:0] sel_952096;
  wire [7:0] add_952099;
  wire [7:0] sel_952100;
  wire [7:0] add_952103;
  wire [7:0] sel_952104;
  wire [7:0] add_952107;
  wire [7:0] sel_952108;
  wire [7:0] add_952111;
  wire [7:0] sel_952112;
  wire [7:0] add_952115;
  wire [7:0] sel_952116;
  wire [7:0] add_952119;
  wire [7:0] sel_952120;
  wire [7:0] add_952123;
  wire [7:0] sel_952124;
  wire [7:0] add_952127;
  wire [7:0] sel_952128;
  wire [7:0] add_952131;
  wire [7:0] sel_952132;
  wire [7:0] add_952135;
  wire [7:0] sel_952136;
  wire [7:0] add_952139;
  wire [7:0] sel_952140;
  wire [7:0] add_952143;
  wire [7:0] sel_952144;
  wire [7:0] add_952147;
  wire [7:0] sel_952148;
  wire [7:0] add_952151;
  wire [7:0] sel_952152;
  wire [7:0] add_952155;
  wire [7:0] sel_952156;
  wire [7:0] add_952159;
  wire [7:0] sel_952160;
  wire [7:0] add_952163;
  wire [7:0] sel_952164;
  wire [7:0] add_952167;
  wire [7:0] sel_952168;
  wire [7:0] add_952171;
  wire [7:0] sel_952172;
  wire [7:0] add_952175;
  wire [7:0] sel_952176;
  wire [7:0] add_952179;
  wire [7:0] sel_952180;
  wire [7:0] add_952183;
  wire [7:0] sel_952184;
  wire [7:0] add_952187;
  wire [7:0] sel_952188;
  wire [7:0] add_952191;
  wire [7:0] sel_952192;
  wire [7:0] add_952195;
  wire [7:0] sel_952196;
  wire [7:0] add_952199;
  wire [7:0] sel_952200;
  wire [7:0] add_952203;
  wire [7:0] sel_952204;
  wire [7:0] add_952207;
  wire [7:0] sel_952208;
  wire [7:0] add_952211;
  wire [7:0] sel_952212;
  wire [7:0] add_952215;
  wire [7:0] sel_952216;
  wire [7:0] add_952219;
  wire [7:0] sel_952220;
  wire [7:0] add_952223;
  wire [7:0] sel_952224;
  wire [7:0] add_952227;
  wire [7:0] sel_952228;
  wire [7:0] add_952231;
  wire [7:0] sel_952232;
  wire [7:0] add_952235;
  wire [7:0] sel_952236;
  wire [7:0] add_952239;
  wire [7:0] sel_952240;
  wire [7:0] add_952243;
  wire [7:0] sel_952244;
  wire [7:0] add_952247;
  wire [7:0] sel_952248;
  wire [7:0] add_952251;
  wire [7:0] sel_952252;
  wire [7:0] add_952255;
  wire [7:0] sel_952256;
  wire [7:0] add_952259;
  wire [7:0] sel_952260;
  wire [7:0] add_952263;
  wire [7:0] sel_952264;
  wire [7:0] add_952267;
  wire [7:0] sel_952268;
  wire [7:0] add_952271;
  wire [7:0] sel_952272;
  wire [7:0] add_952275;
  wire [7:0] sel_952276;
  wire [7:0] add_952279;
  wire [7:0] sel_952280;
  wire [7:0] add_952283;
  wire [7:0] sel_952284;
  wire [7:0] add_952287;
  wire [7:0] sel_952288;
  wire [7:0] add_952291;
  wire [7:0] sel_952292;
  wire [7:0] add_952295;
  wire [7:0] sel_952296;
  wire [7:0] add_952299;
  wire [7:0] sel_952300;
  wire [7:0] add_952303;
  wire [7:0] sel_952304;
  wire [7:0] add_952308;
  wire [15:0] array_index_952309;
  wire [7:0] sel_952310;
  wire [7:0] add_952313;
  wire [7:0] sel_952314;
  wire [7:0] add_952317;
  wire [7:0] sel_952318;
  wire [7:0] add_952321;
  wire [7:0] sel_952322;
  wire [7:0] add_952325;
  wire [7:0] sel_952326;
  wire [7:0] add_952329;
  wire [7:0] sel_952330;
  wire [7:0] add_952333;
  wire [7:0] sel_952334;
  wire [7:0] add_952337;
  wire [7:0] sel_952338;
  wire [7:0] add_952341;
  wire [7:0] sel_952342;
  wire [7:0] add_952345;
  wire [7:0] sel_952346;
  wire [7:0] add_952349;
  wire [7:0] sel_952350;
  wire [7:0] add_952353;
  wire [7:0] sel_952354;
  wire [7:0] add_952357;
  wire [7:0] sel_952358;
  wire [7:0] add_952361;
  wire [7:0] sel_952362;
  wire [7:0] add_952365;
  wire [7:0] sel_952366;
  wire [7:0] add_952369;
  wire [7:0] sel_952370;
  wire [7:0] add_952373;
  wire [7:0] sel_952374;
  wire [7:0] add_952377;
  wire [7:0] sel_952378;
  wire [7:0] add_952381;
  wire [7:0] sel_952382;
  wire [7:0] add_952385;
  wire [7:0] sel_952386;
  wire [7:0] add_952389;
  wire [7:0] sel_952390;
  wire [7:0] add_952393;
  wire [7:0] sel_952394;
  wire [7:0] add_952397;
  wire [7:0] sel_952398;
  wire [7:0] add_952401;
  wire [7:0] sel_952402;
  wire [7:0] add_952405;
  wire [7:0] sel_952406;
  wire [7:0] add_952409;
  wire [7:0] sel_952410;
  wire [7:0] add_952413;
  wire [7:0] sel_952414;
  wire [7:0] add_952417;
  wire [7:0] sel_952418;
  wire [7:0] add_952421;
  wire [7:0] sel_952422;
  wire [7:0] add_952425;
  wire [7:0] sel_952426;
  wire [7:0] add_952429;
  wire [7:0] sel_952430;
  wire [7:0] add_952433;
  wire [7:0] sel_952434;
  wire [7:0] add_952437;
  wire [7:0] sel_952438;
  wire [7:0] add_952441;
  wire [7:0] sel_952442;
  wire [7:0] add_952445;
  wire [7:0] sel_952446;
  wire [7:0] add_952449;
  wire [7:0] sel_952450;
  wire [7:0] add_952453;
  wire [7:0] sel_952454;
  wire [7:0] add_952457;
  wire [7:0] sel_952458;
  wire [7:0] add_952461;
  wire [7:0] sel_952462;
  wire [7:0] add_952465;
  wire [7:0] sel_952466;
  wire [7:0] add_952469;
  wire [7:0] sel_952470;
  wire [7:0] add_952473;
  wire [7:0] sel_952474;
  wire [7:0] add_952477;
  wire [7:0] sel_952478;
  wire [7:0] add_952481;
  wire [7:0] sel_952482;
  wire [7:0] add_952485;
  wire [7:0] sel_952486;
  wire [7:0] add_952489;
  wire [7:0] sel_952490;
  wire [7:0] add_952493;
  wire [7:0] sel_952494;
  wire [7:0] add_952497;
  wire [7:0] sel_952498;
  wire [7:0] add_952501;
  wire [7:0] sel_952502;
  wire [7:0] add_952505;
  wire [7:0] sel_952506;
  wire [7:0] add_952509;
  wire [7:0] sel_952510;
  wire [7:0] add_952513;
  wire [7:0] sel_952514;
  wire [7:0] add_952517;
  wire [7:0] sel_952518;
  wire [7:0] add_952521;
  wire [7:0] sel_952522;
  wire [7:0] add_952525;
  wire [7:0] sel_952526;
  wire [7:0] add_952529;
  wire [7:0] sel_952530;
  wire [7:0] add_952533;
  wire [7:0] sel_952534;
  wire [7:0] add_952537;
  wire [7:0] sel_952538;
  wire [7:0] add_952541;
  wire [7:0] sel_952542;
  wire [7:0] add_952545;
  wire [7:0] sel_952546;
  wire [7:0] add_952549;
  wire [7:0] sel_952550;
  wire [7:0] add_952553;
  wire [7:0] sel_952554;
  wire [7:0] add_952557;
  wire [7:0] sel_952558;
  wire [7:0] add_952561;
  wire [7:0] sel_952562;
  wire [7:0] add_952565;
  wire [7:0] sel_952566;
  wire [7:0] add_952569;
  wire [7:0] sel_952570;
  wire [7:0] add_952573;
  wire [7:0] sel_952574;
  wire [7:0] add_952577;
  wire [7:0] sel_952578;
  wire [7:0] add_952581;
  wire [7:0] sel_952582;
  wire [7:0] add_952585;
  wire [7:0] sel_952586;
  wire [7:0] add_952589;
  wire [7:0] sel_952590;
  wire [7:0] add_952593;
  wire [7:0] sel_952594;
  wire [7:0] add_952597;
  wire [7:0] sel_952598;
  wire [7:0] add_952601;
  wire [7:0] sel_952602;
  wire [7:0] add_952605;
  wire [7:0] sel_952606;
  wire [7:0] add_952609;
  wire [7:0] sel_952610;
  wire [7:0] add_952613;
  wire [7:0] sel_952614;
  wire [7:0] add_952617;
  wire [7:0] sel_952618;
  wire [7:0] add_952621;
  wire [7:0] sel_952622;
  wire [7:0] add_952625;
  wire [7:0] sel_952626;
  wire [7:0] add_952629;
  wire [7:0] sel_952630;
  wire [7:0] add_952633;
  wire [7:0] sel_952634;
  wire [7:0] add_952637;
  wire [7:0] sel_952638;
  wire [7:0] add_952641;
  wire [7:0] sel_952642;
  wire [7:0] add_952645;
  wire [7:0] sel_952646;
  wire [7:0] add_952649;
  wire [7:0] sel_952650;
  wire [7:0] add_952653;
  wire [7:0] sel_952654;
  wire [7:0] add_952657;
  wire [7:0] sel_952658;
  wire [7:0] add_952661;
  wire [7:0] sel_952662;
  wire [7:0] add_952665;
  wire [7:0] sel_952666;
  wire [7:0] add_952669;
  wire [7:0] sel_952670;
  wire [7:0] add_952673;
  wire [7:0] sel_952674;
  wire [7:0] add_952677;
  wire [7:0] sel_952678;
  wire [7:0] add_952681;
  wire [7:0] sel_952682;
  wire [7:0] add_952685;
  wire [7:0] sel_952686;
  wire [7:0] add_952689;
  wire [7:0] sel_952690;
  wire [7:0] add_952693;
  wire [7:0] sel_952694;
  wire [7:0] add_952697;
  wire [7:0] sel_952698;
  wire [7:0] add_952701;
  wire [7:0] sel_952702;
  wire [7:0] add_952705;
  wire [7:0] sel_952706;
  wire [7:0] add_952710;
  wire [15:0] array_index_952711;
  wire [7:0] sel_952712;
  wire [7:0] add_952715;
  wire [7:0] sel_952716;
  wire [7:0] add_952719;
  wire [7:0] sel_952720;
  wire [7:0] add_952723;
  wire [7:0] sel_952724;
  wire [7:0] add_952727;
  wire [7:0] sel_952728;
  wire [7:0] add_952731;
  wire [7:0] sel_952732;
  wire [7:0] add_952735;
  wire [7:0] sel_952736;
  wire [7:0] add_952739;
  wire [7:0] sel_952740;
  wire [7:0] add_952743;
  wire [7:0] sel_952744;
  wire [7:0] add_952747;
  wire [7:0] sel_952748;
  wire [7:0] add_952751;
  wire [7:0] sel_952752;
  wire [7:0] add_952755;
  wire [7:0] sel_952756;
  wire [7:0] add_952759;
  wire [7:0] sel_952760;
  wire [7:0] add_952763;
  wire [7:0] sel_952764;
  wire [7:0] add_952767;
  wire [7:0] sel_952768;
  wire [7:0] add_952771;
  wire [7:0] sel_952772;
  wire [7:0] add_952775;
  wire [7:0] sel_952776;
  wire [7:0] add_952779;
  wire [7:0] sel_952780;
  wire [7:0] add_952783;
  wire [7:0] sel_952784;
  wire [7:0] add_952787;
  wire [7:0] sel_952788;
  wire [7:0] add_952791;
  wire [7:0] sel_952792;
  wire [7:0] add_952795;
  wire [7:0] sel_952796;
  wire [7:0] add_952799;
  wire [7:0] sel_952800;
  wire [7:0] add_952803;
  wire [7:0] sel_952804;
  wire [7:0] add_952807;
  wire [7:0] sel_952808;
  wire [7:0] add_952811;
  wire [7:0] sel_952812;
  wire [7:0] add_952815;
  wire [7:0] sel_952816;
  wire [7:0] add_952819;
  wire [7:0] sel_952820;
  wire [7:0] add_952823;
  wire [7:0] sel_952824;
  wire [7:0] add_952827;
  wire [7:0] sel_952828;
  wire [7:0] add_952831;
  wire [7:0] sel_952832;
  wire [7:0] add_952835;
  wire [7:0] sel_952836;
  wire [7:0] add_952839;
  wire [7:0] sel_952840;
  wire [7:0] add_952843;
  wire [7:0] sel_952844;
  wire [7:0] add_952847;
  wire [7:0] sel_952848;
  wire [7:0] add_952851;
  wire [7:0] sel_952852;
  wire [7:0] add_952855;
  wire [7:0] sel_952856;
  wire [7:0] add_952859;
  wire [7:0] sel_952860;
  wire [7:0] add_952863;
  wire [7:0] sel_952864;
  wire [7:0] add_952867;
  wire [7:0] sel_952868;
  wire [7:0] add_952871;
  wire [7:0] sel_952872;
  wire [7:0] add_952875;
  wire [7:0] sel_952876;
  wire [7:0] add_952879;
  wire [7:0] sel_952880;
  wire [7:0] add_952883;
  wire [7:0] sel_952884;
  wire [7:0] add_952887;
  wire [7:0] sel_952888;
  wire [7:0] add_952891;
  wire [7:0] sel_952892;
  wire [7:0] add_952895;
  wire [7:0] sel_952896;
  wire [7:0] add_952899;
  wire [7:0] sel_952900;
  wire [7:0] add_952903;
  wire [7:0] sel_952904;
  wire [7:0] add_952907;
  wire [7:0] sel_952908;
  wire [7:0] add_952911;
  wire [7:0] sel_952912;
  wire [7:0] add_952915;
  wire [7:0] sel_952916;
  wire [7:0] add_952919;
  wire [7:0] sel_952920;
  wire [7:0] add_952923;
  wire [7:0] sel_952924;
  wire [7:0] add_952927;
  wire [7:0] sel_952928;
  wire [7:0] add_952931;
  wire [7:0] sel_952932;
  wire [7:0] add_952935;
  wire [7:0] sel_952936;
  wire [7:0] add_952939;
  wire [7:0] sel_952940;
  wire [7:0] add_952943;
  wire [7:0] sel_952944;
  wire [7:0] add_952947;
  wire [7:0] sel_952948;
  wire [7:0] add_952951;
  wire [7:0] sel_952952;
  wire [7:0] add_952955;
  wire [7:0] sel_952956;
  wire [7:0] add_952959;
  wire [7:0] sel_952960;
  wire [7:0] add_952963;
  wire [7:0] sel_952964;
  wire [7:0] add_952967;
  wire [7:0] sel_952968;
  wire [7:0] add_952971;
  wire [7:0] sel_952972;
  wire [7:0] add_952975;
  wire [7:0] sel_952976;
  wire [7:0] add_952979;
  wire [7:0] sel_952980;
  wire [7:0] add_952983;
  wire [7:0] sel_952984;
  wire [7:0] add_952987;
  wire [7:0] sel_952988;
  wire [7:0] add_952991;
  wire [7:0] sel_952992;
  wire [7:0] add_952995;
  wire [7:0] sel_952996;
  wire [7:0] add_952999;
  wire [7:0] sel_953000;
  wire [7:0] add_953003;
  wire [7:0] sel_953004;
  wire [7:0] add_953007;
  wire [7:0] sel_953008;
  wire [7:0] add_953011;
  wire [7:0] sel_953012;
  wire [7:0] add_953015;
  wire [7:0] sel_953016;
  wire [7:0] add_953019;
  wire [7:0] sel_953020;
  wire [7:0] add_953023;
  wire [7:0] sel_953024;
  wire [7:0] add_953027;
  wire [7:0] sel_953028;
  wire [7:0] add_953031;
  wire [7:0] sel_953032;
  wire [7:0] add_953035;
  wire [7:0] sel_953036;
  wire [7:0] add_953039;
  wire [7:0] sel_953040;
  wire [7:0] add_953043;
  wire [7:0] sel_953044;
  wire [7:0] add_953047;
  wire [7:0] sel_953048;
  wire [7:0] add_953051;
  wire [7:0] sel_953052;
  wire [7:0] add_953055;
  wire [7:0] sel_953056;
  wire [7:0] add_953059;
  wire [7:0] sel_953060;
  wire [7:0] add_953063;
  wire [7:0] sel_953064;
  wire [7:0] add_953067;
  wire [7:0] sel_953068;
  wire [7:0] add_953071;
  wire [7:0] sel_953072;
  wire [7:0] add_953075;
  wire [7:0] sel_953076;
  wire [7:0] add_953079;
  wire [7:0] sel_953080;
  wire [7:0] add_953083;
  wire [7:0] sel_953084;
  wire [7:0] add_953087;
  wire [7:0] sel_953088;
  wire [7:0] add_953091;
  wire [7:0] sel_953092;
  wire [7:0] add_953095;
  wire [7:0] sel_953096;
  wire [7:0] add_953099;
  wire [7:0] sel_953100;
  wire [7:0] add_953103;
  wire [7:0] sel_953104;
  wire [7:0] add_953107;
  wire [7:0] sel_953108;
  wire [7:0] add_953112;
  wire [15:0] array_index_953113;
  wire [7:0] sel_953114;
  wire [7:0] add_953117;
  wire [7:0] sel_953118;
  wire [7:0] add_953121;
  wire [7:0] sel_953122;
  wire [7:0] add_953125;
  wire [7:0] sel_953126;
  wire [7:0] add_953129;
  wire [7:0] sel_953130;
  wire [7:0] add_953133;
  wire [7:0] sel_953134;
  wire [7:0] add_953137;
  wire [7:0] sel_953138;
  wire [7:0] add_953141;
  wire [7:0] sel_953142;
  wire [7:0] add_953145;
  wire [7:0] sel_953146;
  wire [7:0] add_953149;
  wire [7:0] sel_953150;
  wire [7:0] add_953153;
  wire [7:0] sel_953154;
  wire [7:0] add_953157;
  wire [7:0] sel_953158;
  wire [7:0] add_953161;
  wire [7:0] sel_953162;
  wire [7:0] add_953165;
  wire [7:0] sel_953166;
  wire [7:0] add_953169;
  wire [7:0] sel_953170;
  wire [7:0] add_953173;
  wire [7:0] sel_953174;
  wire [7:0] add_953177;
  wire [7:0] sel_953178;
  wire [7:0] add_953181;
  wire [7:0] sel_953182;
  wire [7:0] add_953185;
  wire [7:0] sel_953186;
  wire [7:0] add_953189;
  wire [7:0] sel_953190;
  wire [7:0] add_953193;
  wire [7:0] sel_953194;
  wire [7:0] add_953197;
  wire [7:0] sel_953198;
  wire [7:0] add_953201;
  wire [7:0] sel_953202;
  wire [7:0] add_953205;
  wire [7:0] sel_953206;
  wire [7:0] add_953209;
  wire [7:0] sel_953210;
  wire [7:0] add_953213;
  wire [7:0] sel_953214;
  wire [7:0] add_953217;
  wire [7:0] sel_953218;
  wire [7:0] add_953221;
  wire [7:0] sel_953222;
  wire [7:0] add_953225;
  wire [7:0] sel_953226;
  wire [7:0] add_953229;
  wire [7:0] sel_953230;
  wire [7:0] add_953233;
  wire [7:0] sel_953234;
  wire [7:0] add_953237;
  wire [7:0] sel_953238;
  wire [7:0] add_953241;
  wire [7:0] sel_953242;
  wire [7:0] add_953245;
  wire [7:0] sel_953246;
  wire [7:0] add_953249;
  wire [7:0] sel_953250;
  wire [7:0] add_953253;
  wire [7:0] sel_953254;
  wire [7:0] add_953257;
  wire [7:0] sel_953258;
  wire [7:0] add_953261;
  wire [7:0] sel_953262;
  wire [7:0] add_953265;
  wire [7:0] sel_953266;
  wire [7:0] add_953269;
  wire [7:0] sel_953270;
  wire [7:0] add_953273;
  wire [7:0] sel_953274;
  wire [7:0] add_953277;
  wire [7:0] sel_953278;
  wire [7:0] add_953281;
  wire [7:0] sel_953282;
  wire [7:0] add_953285;
  wire [7:0] sel_953286;
  wire [7:0] add_953289;
  wire [7:0] sel_953290;
  wire [7:0] add_953293;
  wire [7:0] sel_953294;
  wire [7:0] add_953297;
  wire [7:0] sel_953298;
  wire [7:0] add_953301;
  wire [7:0] sel_953302;
  wire [7:0] add_953305;
  wire [7:0] sel_953306;
  wire [7:0] add_953309;
  wire [7:0] sel_953310;
  wire [7:0] add_953313;
  wire [7:0] sel_953314;
  wire [7:0] add_953317;
  wire [7:0] sel_953318;
  wire [7:0] add_953321;
  wire [7:0] sel_953322;
  wire [7:0] add_953325;
  wire [7:0] sel_953326;
  wire [7:0] add_953329;
  wire [7:0] sel_953330;
  wire [7:0] add_953333;
  wire [7:0] sel_953334;
  wire [7:0] add_953337;
  wire [7:0] sel_953338;
  wire [7:0] add_953341;
  wire [7:0] sel_953342;
  wire [7:0] add_953345;
  wire [7:0] sel_953346;
  wire [7:0] add_953349;
  wire [7:0] sel_953350;
  wire [7:0] add_953353;
  wire [7:0] sel_953354;
  wire [7:0] add_953357;
  wire [7:0] sel_953358;
  wire [7:0] add_953361;
  wire [7:0] sel_953362;
  wire [7:0] add_953365;
  wire [7:0] sel_953366;
  wire [7:0] add_953369;
  wire [7:0] sel_953370;
  wire [7:0] add_953373;
  wire [7:0] sel_953374;
  wire [7:0] add_953377;
  wire [7:0] sel_953378;
  wire [7:0] add_953381;
  wire [7:0] sel_953382;
  wire [7:0] add_953385;
  wire [7:0] sel_953386;
  wire [7:0] add_953389;
  wire [7:0] sel_953390;
  wire [7:0] add_953393;
  wire [7:0] sel_953394;
  wire [7:0] add_953397;
  wire [7:0] sel_953398;
  wire [7:0] add_953401;
  wire [7:0] sel_953402;
  wire [7:0] add_953405;
  wire [7:0] sel_953406;
  wire [7:0] add_953409;
  wire [7:0] sel_953410;
  wire [7:0] add_953413;
  wire [7:0] sel_953414;
  wire [7:0] add_953417;
  wire [7:0] sel_953418;
  wire [7:0] add_953421;
  wire [7:0] sel_953422;
  wire [7:0] add_953425;
  wire [7:0] sel_953426;
  wire [7:0] add_953429;
  wire [7:0] sel_953430;
  wire [7:0] add_953433;
  wire [7:0] sel_953434;
  wire [7:0] add_953437;
  wire [7:0] sel_953438;
  wire [7:0] add_953441;
  wire [7:0] sel_953442;
  wire [7:0] add_953445;
  wire [7:0] sel_953446;
  wire [7:0] add_953449;
  wire [7:0] sel_953450;
  wire [7:0] add_953453;
  wire [7:0] sel_953454;
  wire [7:0] add_953457;
  wire [7:0] sel_953458;
  wire [7:0] add_953461;
  wire [7:0] sel_953462;
  wire [7:0] add_953465;
  wire [7:0] sel_953466;
  wire [7:0] add_953469;
  wire [7:0] sel_953470;
  wire [7:0] add_953473;
  wire [7:0] sel_953474;
  wire [7:0] add_953477;
  wire [7:0] sel_953478;
  wire [7:0] add_953481;
  wire [7:0] sel_953482;
  wire [7:0] add_953485;
  wire [7:0] sel_953486;
  wire [7:0] add_953489;
  wire [7:0] sel_953490;
  wire [7:0] add_953493;
  wire [7:0] sel_953494;
  wire [7:0] add_953497;
  wire [7:0] sel_953498;
  wire [7:0] add_953501;
  wire [7:0] sel_953502;
  wire [7:0] add_953505;
  wire [7:0] sel_953506;
  wire [7:0] add_953509;
  wire [7:0] sel_953510;
  wire [7:0] add_953514;
  wire [15:0] array_index_953515;
  wire [7:0] sel_953516;
  wire [7:0] add_953519;
  wire [7:0] sel_953520;
  wire [7:0] add_953523;
  wire [7:0] sel_953524;
  wire [7:0] add_953527;
  wire [7:0] sel_953528;
  wire [7:0] add_953531;
  wire [7:0] sel_953532;
  wire [7:0] add_953535;
  wire [7:0] sel_953536;
  wire [7:0] add_953539;
  wire [7:0] sel_953540;
  wire [7:0] add_953543;
  wire [7:0] sel_953544;
  wire [7:0] add_953547;
  wire [7:0] sel_953548;
  wire [7:0] add_953551;
  wire [7:0] sel_953552;
  wire [7:0] add_953555;
  wire [7:0] sel_953556;
  wire [7:0] add_953559;
  wire [7:0] sel_953560;
  wire [7:0] add_953563;
  wire [7:0] sel_953564;
  wire [7:0] add_953567;
  wire [7:0] sel_953568;
  wire [7:0] add_953571;
  wire [7:0] sel_953572;
  wire [7:0] add_953575;
  wire [7:0] sel_953576;
  wire [7:0] add_953579;
  wire [7:0] sel_953580;
  wire [7:0] add_953583;
  wire [7:0] sel_953584;
  wire [7:0] add_953587;
  wire [7:0] sel_953588;
  wire [7:0] add_953591;
  wire [7:0] sel_953592;
  wire [7:0] add_953595;
  wire [7:0] sel_953596;
  wire [7:0] add_953599;
  wire [7:0] sel_953600;
  wire [7:0] add_953603;
  wire [7:0] sel_953604;
  wire [7:0] add_953607;
  wire [7:0] sel_953608;
  wire [7:0] add_953611;
  wire [7:0] sel_953612;
  wire [7:0] add_953615;
  wire [7:0] sel_953616;
  wire [7:0] add_953619;
  wire [7:0] sel_953620;
  wire [7:0] add_953623;
  wire [7:0] sel_953624;
  wire [7:0] add_953627;
  wire [7:0] sel_953628;
  wire [7:0] add_953631;
  wire [7:0] sel_953632;
  wire [7:0] add_953635;
  wire [7:0] sel_953636;
  wire [7:0] add_953639;
  wire [7:0] sel_953640;
  wire [7:0] add_953643;
  wire [7:0] sel_953644;
  wire [7:0] add_953647;
  wire [7:0] sel_953648;
  wire [7:0] add_953651;
  wire [7:0] sel_953652;
  wire [7:0] add_953655;
  wire [7:0] sel_953656;
  wire [7:0] add_953659;
  wire [7:0] sel_953660;
  wire [7:0] add_953663;
  wire [7:0] sel_953664;
  wire [7:0] add_953667;
  wire [7:0] sel_953668;
  wire [7:0] add_953671;
  wire [7:0] sel_953672;
  wire [7:0] add_953675;
  wire [7:0] sel_953676;
  wire [7:0] add_953679;
  wire [7:0] sel_953680;
  wire [7:0] add_953683;
  wire [7:0] sel_953684;
  wire [7:0] add_953687;
  wire [7:0] sel_953688;
  wire [7:0] add_953691;
  wire [7:0] sel_953692;
  wire [7:0] add_953695;
  wire [7:0] sel_953696;
  wire [7:0] add_953699;
  wire [7:0] sel_953700;
  wire [7:0] add_953703;
  wire [7:0] sel_953704;
  wire [7:0] add_953707;
  wire [7:0] sel_953708;
  wire [7:0] add_953711;
  wire [7:0] sel_953712;
  wire [7:0] add_953715;
  wire [7:0] sel_953716;
  wire [7:0] add_953719;
  wire [7:0] sel_953720;
  wire [7:0] add_953723;
  wire [7:0] sel_953724;
  wire [7:0] add_953727;
  wire [7:0] sel_953728;
  wire [7:0] add_953731;
  wire [7:0] sel_953732;
  wire [7:0] add_953735;
  wire [7:0] sel_953736;
  wire [7:0] add_953739;
  wire [7:0] sel_953740;
  wire [7:0] add_953743;
  wire [7:0] sel_953744;
  wire [7:0] add_953747;
  wire [7:0] sel_953748;
  wire [7:0] add_953751;
  wire [7:0] sel_953752;
  wire [7:0] add_953755;
  wire [7:0] sel_953756;
  wire [7:0] add_953759;
  wire [7:0] sel_953760;
  wire [7:0] add_953763;
  wire [7:0] sel_953764;
  wire [7:0] add_953767;
  wire [7:0] sel_953768;
  wire [7:0] add_953771;
  wire [7:0] sel_953772;
  wire [7:0] add_953775;
  wire [7:0] sel_953776;
  wire [7:0] add_953779;
  wire [7:0] sel_953780;
  wire [7:0] add_953783;
  wire [7:0] sel_953784;
  wire [7:0] add_953787;
  wire [7:0] sel_953788;
  wire [7:0] add_953791;
  wire [7:0] sel_953792;
  wire [7:0] add_953795;
  wire [7:0] sel_953796;
  wire [7:0] add_953799;
  wire [7:0] sel_953800;
  wire [7:0] add_953803;
  wire [7:0] sel_953804;
  wire [7:0] add_953807;
  wire [7:0] sel_953808;
  wire [7:0] add_953811;
  wire [7:0] sel_953812;
  wire [7:0] add_953815;
  wire [7:0] sel_953816;
  wire [7:0] add_953819;
  wire [7:0] sel_953820;
  wire [7:0] add_953823;
  wire [7:0] sel_953824;
  wire [7:0] add_953827;
  wire [7:0] sel_953828;
  wire [7:0] add_953831;
  wire [7:0] sel_953832;
  wire [7:0] add_953835;
  wire [7:0] sel_953836;
  wire [7:0] add_953839;
  wire [7:0] sel_953840;
  wire [7:0] add_953843;
  wire [7:0] sel_953844;
  wire [7:0] add_953847;
  wire [7:0] sel_953848;
  wire [7:0] add_953851;
  wire [7:0] sel_953852;
  wire [7:0] add_953855;
  wire [7:0] sel_953856;
  wire [7:0] add_953859;
  wire [7:0] sel_953860;
  wire [7:0] add_953863;
  wire [7:0] sel_953864;
  wire [7:0] add_953867;
  wire [7:0] sel_953868;
  wire [7:0] add_953871;
  wire [7:0] sel_953872;
  wire [7:0] add_953875;
  wire [7:0] sel_953876;
  wire [7:0] add_953879;
  wire [7:0] sel_953880;
  wire [7:0] add_953883;
  wire [7:0] sel_953884;
  wire [7:0] add_953887;
  wire [7:0] sel_953888;
  wire [7:0] add_953891;
  wire [7:0] sel_953892;
  wire [7:0] add_953895;
  wire [7:0] sel_953896;
  wire [7:0] add_953899;
  wire [7:0] sel_953900;
  wire [7:0] add_953903;
  wire [7:0] sel_953904;
  wire [7:0] add_953907;
  wire [7:0] sel_953908;
  wire [7:0] add_953911;
  wire [7:0] sel_953912;
  wire [7:0] add_953916;
  wire [15:0] array_index_953917;
  wire [7:0] sel_953918;
  wire [7:0] add_953921;
  wire [7:0] sel_953922;
  wire [7:0] add_953925;
  wire [7:0] sel_953926;
  wire [7:0] add_953929;
  wire [7:0] sel_953930;
  wire [7:0] add_953933;
  wire [7:0] sel_953934;
  wire [7:0] add_953937;
  wire [7:0] sel_953938;
  wire [7:0] add_953941;
  wire [7:0] sel_953942;
  wire [7:0] add_953945;
  wire [7:0] sel_953946;
  wire [7:0] add_953949;
  wire [7:0] sel_953950;
  wire [7:0] add_953953;
  wire [7:0] sel_953954;
  wire [7:0] add_953957;
  wire [7:0] sel_953958;
  wire [7:0] add_953961;
  wire [7:0] sel_953962;
  wire [7:0] add_953965;
  wire [7:0] sel_953966;
  wire [7:0] add_953969;
  wire [7:0] sel_953970;
  wire [7:0] add_953973;
  wire [7:0] sel_953974;
  wire [7:0] add_953977;
  wire [7:0] sel_953978;
  wire [7:0] add_953981;
  wire [7:0] sel_953982;
  wire [7:0] add_953985;
  wire [7:0] sel_953986;
  wire [7:0] add_953989;
  wire [7:0] sel_953990;
  wire [7:0] add_953993;
  wire [7:0] sel_953994;
  wire [7:0] add_953997;
  wire [7:0] sel_953998;
  wire [7:0] add_954001;
  wire [7:0] sel_954002;
  wire [7:0] add_954005;
  wire [7:0] sel_954006;
  wire [7:0] add_954009;
  wire [7:0] sel_954010;
  wire [7:0] add_954013;
  wire [7:0] sel_954014;
  wire [7:0] add_954017;
  wire [7:0] sel_954018;
  wire [7:0] add_954021;
  wire [7:0] sel_954022;
  wire [7:0] add_954025;
  wire [7:0] sel_954026;
  wire [7:0] add_954029;
  wire [7:0] sel_954030;
  wire [7:0] add_954033;
  wire [7:0] sel_954034;
  wire [7:0] add_954037;
  wire [7:0] sel_954038;
  wire [7:0] add_954041;
  wire [7:0] sel_954042;
  wire [7:0] add_954045;
  wire [7:0] sel_954046;
  wire [7:0] add_954049;
  wire [7:0] sel_954050;
  wire [7:0] add_954053;
  wire [7:0] sel_954054;
  wire [7:0] add_954057;
  wire [7:0] sel_954058;
  wire [7:0] add_954061;
  wire [7:0] sel_954062;
  wire [7:0] add_954065;
  wire [7:0] sel_954066;
  wire [7:0] add_954069;
  wire [7:0] sel_954070;
  wire [7:0] add_954073;
  wire [7:0] sel_954074;
  wire [7:0] add_954077;
  wire [7:0] sel_954078;
  wire [7:0] add_954081;
  wire [7:0] sel_954082;
  wire [7:0] add_954085;
  wire [7:0] sel_954086;
  wire [7:0] add_954089;
  wire [7:0] sel_954090;
  wire [7:0] add_954093;
  wire [7:0] sel_954094;
  wire [7:0] add_954097;
  wire [7:0] sel_954098;
  wire [7:0] add_954101;
  wire [7:0] sel_954102;
  wire [7:0] add_954105;
  wire [7:0] sel_954106;
  wire [7:0] add_954109;
  wire [7:0] sel_954110;
  wire [7:0] add_954113;
  wire [7:0] sel_954114;
  wire [7:0] add_954117;
  wire [7:0] sel_954118;
  wire [7:0] add_954121;
  wire [7:0] sel_954122;
  wire [7:0] add_954125;
  wire [7:0] sel_954126;
  wire [7:0] add_954129;
  wire [7:0] sel_954130;
  wire [7:0] add_954133;
  wire [7:0] sel_954134;
  wire [7:0] add_954137;
  wire [7:0] sel_954138;
  wire [7:0] add_954141;
  wire [7:0] sel_954142;
  wire [7:0] add_954145;
  wire [7:0] sel_954146;
  wire [7:0] add_954149;
  wire [7:0] sel_954150;
  wire [7:0] add_954153;
  wire [7:0] sel_954154;
  wire [7:0] add_954157;
  wire [7:0] sel_954158;
  wire [7:0] add_954161;
  wire [7:0] sel_954162;
  wire [7:0] add_954165;
  wire [7:0] sel_954166;
  wire [7:0] add_954169;
  wire [7:0] sel_954170;
  wire [7:0] add_954173;
  wire [7:0] sel_954174;
  wire [7:0] add_954177;
  wire [7:0] sel_954178;
  wire [7:0] add_954181;
  wire [7:0] sel_954182;
  wire [7:0] add_954185;
  wire [7:0] sel_954186;
  wire [7:0] add_954189;
  wire [7:0] sel_954190;
  wire [7:0] add_954193;
  wire [7:0] sel_954194;
  wire [7:0] add_954197;
  wire [7:0] sel_954198;
  wire [7:0] add_954201;
  wire [7:0] sel_954202;
  wire [7:0] add_954205;
  wire [7:0] sel_954206;
  wire [7:0] add_954209;
  wire [7:0] sel_954210;
  wire [7:0] add_954213;
  wire [7:0] sel_954214;
  wire [7:0] add_954217;
  wire [7:0] sel_954218;
  wire [7:0] add_954221;
  wire [7:0] sel_954222;
  wire [7:0] add_954225;
  wire [7:0] sel_954226;
  wire [7:0] add_954229;
  wire [7:0] sel_954230;
  wire [7:0] add_954233;
  wire [7:0] sel_954234;
  wire [7:0] add_954237;
  wire [7:0] sel_954238;
  wire [7:0] add_954241;
  wire [7:0] sel_954242;
  wire [7:0] add_954245;
  wire [7:0] sel_954246;
  wire [7:0] add_954249;
  wire [7:0] sel_954250;
  wire [7:0] add_954253;
  wire [7:0] sel_954254;
  wire [7:0] add_954257;
  wire [7:0] sel_954258;
  wire [7:0] add_954261;
  wire [7:0] sel_954262;
  wire [7:0] add_954265;
  wire [7:0] sel_954266;
  wire [7:0] add_954269;
  wire [7:0] sel_954270;
  wire [7:0] add_954273;
  wire [7:0] sel_954274;
  wire [7:0] add_954277;
  wire [7:0] sel_954278;
  wire [7:0] add_954281;
  wire [7:0] sel_954282;
  wire [7:0] add_954285;
  wire [7:0] sel_954286;
  wire [7:0] add_954289;
  wire [7:0] sel_954290;
  wire [7:0] add_954293;
  wire [7:0] sel_954294;
  wire [7:0] add_954297;
  wire [7:0] sel_954298;
  wire [7:0] add_954301;
  wire [7:0] sel_954302;
  wire [7:0] add_954305;
  wire [7:0] sel_954306;
  wire [7:0] add_954309;
  wire [7:0] sel_954310;
  wire [7:0] add_954313;
  wire [7:0] sel_954314;
  wire [7:0] add_954318;
  wire [15:0] array_index_954319;
  wire [7:0] sel_954320;
  wire [7:0] add_954323;
  wire [7:0] sel_954324;
  wire [7:0] add_954327;
  wire [7:0] sel_954328;
  wire [7:0] add_954331;
  wire [7:0] sel_954332;
  wire [7:0] add_954335;
  wire [7:0] sel_954336;
  wire [7:0] add_954339;
  wire [7:0] sel_954340;
  wire [7:0] add_954343;
  wire [7:0] sel_954344;
  wire [7:0] add_954347;
  wire [7:0] sel_954348;
  wire [7:0] add_954351;
  wire [7:0] sel_954352;
  wire [7:0] add_954355;
  wire [7:0] sel_954356;
  wire [7:0] add_954359;
  wire [7:0] sel_954360;
  wire [7:0] add_954363;
  wire [7:0] sel_954364;
  wire [7:0] add_954367;
  wire [7:0] sel_954368;
  wire [7:0] add_954371;
  wire [7:0] sel_954372;
  wire [7:0] add_954375;
  wire [7:0] sel_954376;
  wire [7:0] add_954379;
  wire [7:0] sel_954380;
  wire [7:0] add_954383;
  wire [7:0] sel_954384;
  wire [7:0] add_954387;
  wire [7:0] sel_954388;
  wire [7:0] add_954391;
  wire [7:0] sel_954392;
  wire [7:0] add_954395;
  wire [7:0] sel_954396;
  wire [7:0] add_954399;
  wire [7:0] sel_954400;
  wire [7:0] add_954403;
  wire [7:0] sel_954404;
  wire [7:0] add_954407;
  wire [7:0] sel_954408;
  wire [7:0] add_954411;
  wire [7:0] sel_954412;
  wire [7:0] add_954415;
  wire [7:0] sel_954416;
  wire [7:0] add_954419;
  wire [7:0] sel_954420;
  wire [7:0] add_954423;
  wire [7:0] sel_954424;
  wire [7:0] add_954427;
  wire [7:0] sel_954428;
  wire [7:0] add_954431;
  wire [7:0] sel_954432;
  wire [7:0] add_954435;
  wire [7:0] sel_954436;
  wire [7:0] add_954439;
  wire [7:0] sel_954440;
  wire [7:0] add_954443;
  wire [7:0] sel_954444;
  wire [7:0] add_954447;
  wire [7:0] sel_954448;
  wire [7:0] add_954451;
  wire [7:0] sel_954452;
  wire [7:0] add_954455;
  wire [7:0] sel_954456;
  wire [7:0] add_954459;
  wire [7:0] sel_954460;
  wire [7:0] add_954463;
  wire [7:0] sel_954464;
  wire [7:0] add_954467;
  wire [7:0] sel_954468;
  wire [7:0] add_954471;
  wire [7:0] sel_954472;
  wire [7:0] add_954475;
  wire [7:0] sel_954476;
  wire [7:0] add_954479;
  wire [7:0] sel_954480;
  wire [7:0] add_954483;
  wire [7:0] sel_954484;
  wire [7:0] add_954487;
  wire [7:0] sel_954488;
  wire [7:0] add_954491;
  wire [7:0] sel_954492;
  wire [7:0] add_954495;
  wire [7:0] sel_954496;
  wire [7:0] add_954499;
  wire [7:0] sel_954500;
  wire [7:0] add_954503;
  wire [7:0] sel_954504;
  wire [7:0] add_954507;
  wire [7:0] sel_954508;
  wire [7:0] add_954511;
  wire [7:0] sel_954512;
  wire [7:0] add_954515;
  wire [7:0] sel_954516;
  wire [7:0] add_954519;
  wire [7:0] sel_954520;
  wire [7:0] add_954523;
  wire [7:0] sel_954524;
  wire [7:0] add_954527;
  wire [7:0] sel_954528;
  wire [7:0] add_954531;
  wire [7:0] sel_954532;
  wire [7:0] add_954535;
  wire [7:0] sel_954536;
  wire [7:0] add_954539;
  wire [7:0] sel_954540;
  wire [7:0] add_954543;
  wire [7:0] sel_954544;
  wire [7:0] add_954547;
  wire [7:0] sel_954548;
  wire [7:0] add_954551;
  wire [7:0] sel_954552;
  wire [7:0] add_954555;
  wire [7:0] sel_954556;
  wire [7:0] add_954559;
  wire [7:0] sel_954560;
  wire [7:0] add_954563;
  wire [7:0] sel_954564;
  wire [7:0] add_954567;
  wire [7:0] sel_954568;
  wire [7:0] add_954571;
  wire [7:0] sel_954572;
  wire [7:0] add_954575;
  wire [7:0] sel_954576;
  wire [7:0] add_954579;
  wire [7:0] sel_954580;
  wire [7:0] add_954583;
  wire [7:0] sel_954584;
  wire [7:0] add_954587;
  wire [7:0] sel_954588;
  wire [7:0] add_954591;
  wire [7:0] sel_954592;
  wire [7:0] add_954595;
  wire [7:0] sel_954596;
  wire [7:0] add_954599;
  wire [7:0] sel_954600;
  wire [7:0] add_954603;
  wire [7:0] sel_954604;
  wire [7:0] add_954607;
  wire [7:0] sel_954608;
  wire [7:0] add_954611;
  wire [7:0] sel_954612;
  wire [7:0] add_954615;
  wire [7:0] sel_954616;
  wire [7:0] add_954619;
  wire [7:0] sel_954620;
  wire [7:0] add_954623;
  wire [7:0] sel_954624;
  wire [7:0] add_954627;
  wire [7:0] sel_954628;
  wire [7:0] add_954631;
  wire [7:0] sel_954632;
  wire [7:0] add_954635;
  wire [7:0] sel_954636;
  wire [7:0] add_954639;
  wire [7:0] sel_954640;
  wire [7:0] add_954643;
  wire [7:0] sel_954644;
  wire [7:0] add_954647;
  wire [7:0] sel_954648;
  wire [7:0] add_954651;
  wire [7:0] sel_954652;
  wire [7:0] add_954655;
  wire [7:0] sel_954656;
  wire [7:0] add_954659;
  wire [7:0] sel_954660;
  wire [7:0] add_954663;
  wire [7:0] sel_954664;
  wire [7:0] add_954667;
  wire [7:0] sel_954668;
  wire [7:0] add_954671;
  wire [7:0] sel_954672;
  wire [7:0] add_954675;
  wire [7:0] sel_954676;
  wire [7:0] add_954679;
  wire [7:0] sel_954680;
  wire [7:0] add_954683;
  wire [7:0] sel_954684;
  wire [7:0] add_954687;
  wire [7:0] sel_954688;
  wire [7:0] add_954691;
  wire [7:0] sel_954692;
  wire [7:0] add_954695;
  wire [7:0] sel_954696;
  wire [7:0] add_954699;
  wire [7:0] sel_954700;
  wire [7:0] add_954703;
  wire [7:0] sel_954704;
  wire [7:0] add_954707;
  wire [7:0] sel_954708;
  wire [7:0] add_954711;
  wire [7:0] sel_954712;
  wire [7:0] add_954715;
  wire [7:0] sel_954716;
  wire [7:0] add_954720;
  wire [15:0] array_index_954721;
  wire [7:0] sel_954722;
  wire [7:0] add_954725;
  wire [7:0] sel_954726;
  wire [7:0] add_954729;
  wire [7:0] sel_954730;
  wire [7:0] add_954733;
  wire [7:0] sel_954734;
  wire [7:0] add_954737;
  wire [7:0] sel_954738;
  wire [7:0] add_954741;
  wire [7:0] sel_954742;
  wire [7:0] add_954745;
  wire [7:0] sel_954746;
  wire [7:0] add_954749;
  wire [7:0] sel_954750;
  wire [7:0] add_954753;
  wire [7:0] sel_954754;
  wire [7:0] add_954757;
  wire [7:0] sel_954758;
  wire [7:0] add_954761;
  wire [7:0] sel_954762;
  wire [7:0] add_954765;
  wire [7:0] sel_954766;
  wire [7:0] add_954769;
  wire [7:0] sel_954770;
  wire [7:0] add_954773;
  wire [7:0] sel_954774;
  wire [7:0] add_954777;
  wire [7:0] sel_954778;
  wire [7:0] add_954781;
  wire [7:0] sel_954782;
  wire [7:0] add_954785;
  wire [7:0] sel_954786;
  wire [7:0] add_954789;
  wire [7:0] sel_954790;
  wire [7:0] add_954793;
  wire [7:0] sel_954794;
  wire [7:0] add_954797;
  wire [7:0] sel_954798;
  wire [7:0] add_954801;
  wire [7:0] sel_954802;
  wire [7:0] add_954805;
  wire [7:0] sel_954806;
  wire [7:0] add_954809;
  wire [7:0] sel_954810;
  wire [7:0] add_954813;
  wire [7:0] sel_954814;
  wire [7:0] add_954817;
  wire [7:0] sel_954818;
  wire [7:0] add_954821;
  wire [7:0] sel_954822;
  wire [7:0] add_954825;
  wire [7:0] sel_954826;
  wire [7:0] add_954829;
  wire [7:0] sel_954830;
  wire [7:0] add_954833;
  wire [7:0] sel_954834;
  wire [7:0] add_954837;
  wire [7:0] sel_954838;
  wire [7:0] add_954841;
  wire [7:0] sel_954842;
  wire [7:0] add_954845;
  wire [7:0] sel_954846;
  wire [7:0] add_954849;
  wire [7:0] sel_954850;
  wire [7:0] add_954853;
  wire [7:0] sel_954854;
  wire [7:0] add_954857;
  wire [7:0] sel_954858;
  wire [7:0] add_954861;
  wire [7:0] sel_954862;
  wire [7:0] add_954865;
  wire [7:0] sel_954866;
  wire [7:0] add_954869;
  wire [7:0] sel_954870;
  wire [7:0] add_954873;
  wire [7:0] sel_954874;
  wire [7:0] add_954877;
  wire [7:0] sel_954878;
  wire [7:0] add_954881;
  wire [7:0] sel_954882;
  wire [7:0] add_954885;
  wire [7:0] sel_954886;
  wire [7:0] add_954889;
  wire [7:0] sel_954890;
  wire [7:0] add_954893;
  wire [7:0] sel_954894;
  wire [7:0] add_954897;
  wire [7:0] sel_954898;
  wire [7:0] add_954901;
  wire [7:0] sel_954902;
  wire [7:0] add_954905;
  wire [7:0] sel_954906;
  wire [7:0] add_954909;
  wire [7:0] sel_954910;
  wire [7:0] add_954913;
  wire [7:0] sel_954914;
  wire [7:0] add_954917;
  wire [7:0] sel_954918;
  wire [7:0] add_954921;
  wire [7:0] sel_954922;
  wire [7:0] add_954925;
  wire [7:0] sel_954926;
  wire [7:0] add_954929;
  wire [7:0] sel_954930;
  wire [7:0] add_954933;
  wire [7:0] sel_954934;
  wire [7:0] add_954937;
  wire [7:0] sel_954938;
  wire [7:0] add_954941;
  wire [7:0] sel_954942;
  wire [7:0] add_954945;
  wire [7:0] sel_954946;
  wire [7:0] add_954949;
  wire [7:0] sel_954950;
  wire [7:0] add_954953;
  wire [7:0] sel_954954;
  wire [7:0] add_954957;
  wire [7:0] sel_954958;
  wire [7:0] add_954961;
  wire [7:0] sel_954962;
  wire [7:0] add_954965;
  wire [7:0] sel_954966;
  wire [7:0] add_954969;
  wire [7:0] sel_954970;
  wire [7:0] add_954973;
  wire [7:0] sel_954974;
  wire [7:0] add_954977;
  wire [7:0] sel_954978;
  wire [7:0] add_954981;
  wire [7:0] sel_954982;
  wire [7:0] add_954985;
  wire [7:0] sel_954986;
  wire [7:0] add_954989;
  wire [7:0] sel_954990;
  wire [7:0] add_954993;
  wire [7:0] sel_954994;
  wire [7:0] add_954997;
  wire [7:0] sel_954998;
  wire [7:0] add_955001;
  wire [7:0] sel_955002;
  wire [7:0] add_955005;
  wire [7:0] sel_955006;
  wire [7:0] add_955009;
  wire [7:0] sel_955010;
  wire [7:0] add_955013;
  wire [7:0] sel_955014;
  wire [7:0] add_955017;
  wire [7:0] sel_955018;
  wire [7:0] add_955021;
  wire [7:0] sel_955022;
  wire [7:0] add_955025;
  wire [7:0] sel_955026;
  wire [7:0] add_955029;
  wire [7:0] sel_955030;
  wire [7:0] add_955033;
  wire [7:0] sel_955034;
  wire [7:0] add_955037;
  wire [7:0] sel_955038;
  wire [7:0] add_955041;
  wire [7:0] sel_955042;
  wire [7:0] add_955045;
  wire [7:0] sel_955046;
  wire [7:0] add_955049;
  wire [7:0] sel_955050;
  wire [7:0] add_955053;
  wire [7:0] sel_955054;
  wire [7:0] add_955057;
  wire [7:0] sel_955058;
  wire [7:0] add_955061;
  wire [7:0] sel_955062;
  wire [7:0] add_955065;
  wire [7:0] sel_955066;
  wire [7:0] add_955069;
  wire [7:0] sel_955070;
  wire [7:0] add_955073;
  wire [7:0] sel_955074;
  wire [7:0] add_955077;
  wire [7:0] sel_955078;
  wire [7:0] add_955081;
  wire [7:0] sel_955082;
  wire [7:0] add_955085;
  wire [7:0] sel_955086;
  wire [7:0] add_955089;
  wire [7:0] sel_955090;
  wire [7:0] add_955093;
  wire [7:0] sel_955094;
  wire [7:0] add_955097;
  wire [7:0] sel_955098;
  wire [7:0] add_955101;
  wire [7:0] sel_955102;
  wire [7:0] add_955105;
  wire [7:0] sel_955106;
  wire [7:0] add_955109;
  wire [7:0] sel_955110;
  wire [7:0] add_955113;
  wire [7:0] sel_955114;
  wire [7:0] add_955117;
  wire [7:0] sel_955118;
  wire [7:0] add_955122;
  wire [15:0] array_index_955123;
  wire [7:0] sel_955124;
  wire [7:0] add_955127;
  wire [7:0] sel_955128;
  wire [7:0] add_955131;
  wire [7:0] sel_955132;
  wire [7:0] add_955135;
  wire [7:0] sel_955136;
  wire [7:0] add_955139;
  wire [7:0] sel_955140;
  wire [7:0] add_955143;
  wire [7:0] sel_955144;
  wire [7:0] add_955147;
  wire [7:0] sel_955148;
  wire [7:0] add_955151;
  wire [7:0] sel_955152;
  wire [7:0] add_955155;
  wire [7:0] sel_955156;
  wire [7:0] add_955159;
  wire [7:0] sel_955160;
  wire [7:0] add_955163;
  wire [7:0] sel_955164;
  wire [7:0] add_955167;
  wire [7:0] sel_955168;
  wire [7:0] add_955171;
  wire [7:0] sel_955172;
  wire [7:0] add_955175;
  wire [7:0] sel_955176;
  wire [7:0] add_955179;
  wire [7:0] sel_955180;
  wire [7:0] add_955183;
  wire [7:0] sel_955184;
  wire [7:0] add_955187;
  wire [7:0] sel_955188;
  wire [7:0] add_955191;
  wire [7:0] sel_955192;
  wire [7:0] add_955195;
  wire [7:0] sel_955196;
  wire [7:0] add_955199;
  wire [7:0] sel_955200;
  wire [7:0] add_955203;
  wire [7:0] sel_955204;
  wire [7:0] add_955207;
  wire [7:0] sel_955208;
  wire [7:0] add_955211;
  wire [7:0] sel_955212;
  wire [7:0] add_955215;
  wire [7:0] sel_955216;
  wire [7:0] add_955219;
  wire [7:0] sel_955220;
  wire [7:0] add_955223;
  wire [7:0] sel_955224;
  wire [7:0] add_955227;
  wire [7:0] sel_955228;
  wire [7:0] add_955231;
  wire [7:0] sel_955232;
  wire [7:0] add_955235;
  wire [7:0] sel_955236;
  wire [7:0] add_955239;
  wire [7:0] sel_955240;
  wire [7:0] add_955243;
  wire [7:0] sel_955244;
  wire [7:0] add_955247;
  wire [7:0] sel_955248;
  wire [7:0] add_955251;
  wire [7:0] sel_955252;
  wire [7:0] add_955255;
  wire [7:0] sel_955256;
  wire [7:0] add_955259;
  wire [7:0] sel_955260;
  wire [7:0] add_955263;
  wire [7:0] sel_955264;
  wire [7:0] add_955267;
  wire [7:0] sel_955268;
  wire [7:0] add_955271;
  wire [7:0] sel_955272;
  wire [7:0] add_955275;
  wire [7:0] sel_955276;
  wire [7:0] add_955279;
  wire [7:0] sel_955280;
  wire [7:0] add_955283;
  wire [7:0] sel_955284;
  wire [7:0] add_955287;
  wire [7:0] sel_955288;
  wire [7:0] add_955291;
  wire [7:0] sel_955292;
  wire [7:0] add_955295;
  wire [7:0] sel_955296;
  wire [7:0] add_955299;
  wire [7:0] sel_955300;
  wire [7:0] add_955303;
  wire [7:0] sel_955304;
  wire [7:0] add_955307;
  wire [7:0] sel_955308;
  wire [7:0] add_955311;
  wire [7:0] sel_955312;
  wire [7:0] add_955315;
  wire [7:0] sel_955316;
  wire [7:0] add_955319;
  wire [7:0] sel_955320;
  wire [7:0] add_955323;
  wire [7:0] sel_955324;
  wire [7:0] add_955327;
  wire [7:0] sel_955328;
  wire [7:0] add_955331;
  wire [7:0] sel_955332;
  wire [7:0] add_955335;
  wire [7:0] sel_955336;
  wire [7:0] add_955339;
  wire [7:0] sel_955340;
  wire [7:0] add_955343;
  wire [7:0] sel_955344;
  wire [7:0] add_955347;
  wire [7:0] sel_955348;
  wire [7:0] add_955351;
  wire [7:0] sel_955352;
  wire [7:0] add_955355;
  wire [7:0] sel_955356;
  wire [7:0] add_955359;
  wire [7:0] sel_955360;
  wire [7:0] add_955363;
  wire [7:0] sel_955364;
  wire [7:0] add_955367;
  wire [7:0] sel_955368;
  wire [7:0] add_955371;
  wire [7:0] sel_955372;
  wire [7:0] add_955375;
  wire [7:0] sel_955376;
  wire [7:0] add_955379;
  wire [7:0] sel_955380;
  wire [7:0] add_955383;
  wire [7:0] sel_955384;
  wire [7:0] add_955387;
  wire [7:0] sel_955388;
  wire [7:0] add_955391;
  wire [7:0] sel_955392;
  wire [7:0] add_955395;
  wire [7:0] sel_955396;
  wire [7:0] add_955399;
  wire [7:0] sel_955400;
  wire [7:0] add_955403;
  wire [7:0] sel_955404;
  wire [7:0] add_955407;
  wire [7:0] sel_955408;
  wire [7:0] add_955411;
  wire [7:0] sel_955412;
  wire [7:0] add_955415;
  wire [7:0] sel_955416;
  wire [7:0] add_955419;
  wire [7:0] sel_955420;
  wire [7:0] add_955423;
  wire [7:0] sel_955424;
  wire [7:0] add_955427;
  wire [7:0] sel_955428;
  wire [7:0] add_955431;
  wire [7:0] sel_955432;
  wire [7:0] add_955435;
  wire [7:0] sel_955436;
  wire [7:0] add_955439;
  wire [7:0] sel_955440;
  wire [7:0] add_955443;
  wire [7:0] sel_955444;
  wire [7:0] add_955447;
  wire [7:0] sel_955448;
  wire [7:0] add_955451;
  wire [7:0] sel_955452;
  wire [7:0] add_955455;
  wire [7:0] sel_955456;
  wire [7:0] add_955459;
  wire [7:0] sel_955460;
  wire [7:0] add_955463;
  wire [7:0] sel_955464;
  wire [7:0] add_955467;
  wire [7:0] sel_955468;
  wire [7:0] add_955471;
  wire [7:0] sel_955472;
  wire [7:0] add_955475;
  wire [7:0] sel_955476;
  wire [7:0] add_955479;
  wire [7:0] sel_955480;
  wire [7:0] add_955483;
  wire [7:0] sel_955484;
  wire [7:0] add_955487;
  wire [7:0] sel_955488;
  wire [7:0] add_955491;
  wire [7:0] sel_955492;
  wire [7:0] add_955495;
  wire [7:0] sel_955496;
  wire [7:0] add_955499;
  wire [7:0] sel_955500;
  wire [7:0] add_955503;
  wire [7:0] sel_955504;
  wire [7:0] add_955507;
  wire [7:0] sel_955508;
  wire [7:0] add_955511;
  wire [7:0] sel_955512;
  wire [7:0] add_955515;
  wire [7:0] sel_955516;
  wire [7:0] add_955519;
  wire [7:0] sel_955520;
  wire [7:0] add_955524;
  wire [15:0] array_index_955525;
  wire [7:0] sel_955526;
  wire [7:0] add_955529;
  wire [7:0] sel_955530;
  wire [7:0] add_955533;
  wire [7:0] sel_955534;
  wire [7:0] add_955537;
  wire [7:0] sel_955538;
  wire [7:0] add_955541;
  wire [7:0] sel_955542;
  wire [7:0] add_955545;
  wire [7:0] sel_955546;
  wire [7:0] add_955549;
  wire [7:0] sel_955550;
  wire [7:0] add_955553;
  wire [7:0] sel_955554;
  wire [7:0] add_955557;
  wire [7:0] sel_955558;
  wire [7:0] add_955561;
  wire [7:0] sel_955562;
  wire [7:0] add_955565;
  wire [7:0] sel_955566;
  wire [7:0] add_955569;
  wire [7:0] sel_955570;
  wire [7:0] add_955573;
  wire [7:0] sel_955574;
  wire [7:0] add_955577;
  wire [7:0] sel_955578;
  wire [7:0] add_955581;
  wire [7:0] sel_955582;
  wire [7:0] add_955585;
  wire [7:0] sel_955586;
  wire [7:0] add_955589;
  wire [7:0] sel_955590;
  wire [7:0] add_955593;
  wire [7:0] sel_955594;
  wire [7:0] add_955597;
  wire [7:0] sel_955598;
  wire [7:0] add_955601;
  wire [7:0] sel_955602;
  wire [7:0] add_955605;
  wire [7:0] sel_955606;
  wire [7:0] add_955609;
  wire [7:0] sel_955610;
  wire [7:0] add_955613;
  wire [7:0] sel_955614;
  wire [7:0] add_955617;
  wire [7:0] sel_955618;
  wire [7:0] add_955621;
  wire [7:0] sel_955622;
  wire [7:0] add_955625;
  wire [7:0] sel_955626;
  wire [7:0] add_955629;
  wire [7:0] sel_955630;
  wire [7:0] add_955633;
  wire [7:0] sel_955634;
  wire [7:0] add_955637;
  wire [7:0] sel_955638;
  wire [7:0] add_955641;
  wire [7:0] sel_955642;
  wire [7:0] add_955645;
  wire [7:0] sel_955646;
  wire [7:0] add_955649;
  wire [7:0] sel_955650;
  wire [7:0] add_955653;
  wire [7:0] sel_955654;
  wire [7:0] add_955657;
  wire [7:0] sel_955658;
  wire [7:0] add_955661;
  wire [7:0] sel_955662;
  wire [7:0] add_955665;
  wire [7:0] sel_955666;
  wire [7:0] add_955669;
  wire [7:0] sel_955670;
  wire [7:0] add_955673;
  wire [7:0] sel_955674;
  wire [7:0] add_955677;
  wire [7:0] sel_955678;
  wire [7:0] add_955681;
  wire [7:0] sel_955682;
  wire [7:0] add_955685;
  wire [7:0] sel_955686;
  wire [7:0] add_955689;
  wire [7:0] sel_955690;
  wire [7:0] add_955693;
  wire [7:0] sel_955694;
  wire [7:0] add_955697;
  wire [7:0] sel_955698;
  wire [7:0] add_955701;
  wire [7:0] sel_955702;
  wire [7:0] add_955705;
  wire [7:0] sel_955706;
  wire [7:0] add_955709;
  wire [7:0] sel_955710;
  wire [7:0] add_955713;
  wire [7:0] sel_955714;
  wire [7:0] add_955717;
  wire [7:0] sel_955718;
  wire [7:0] add_955721;
  wire [7:0] sel_955722;
  wire [7:0] add_955725;
  wire [7:0] sel_955726;
  wire [7:0] add_955729;
  wire [7:0] sel_955730;
  wire [7:0] add_955733;
  wire [7:0] sel_955734;
  wire [7:0] add_955737;
  wire [7:0] sel_955738;
  wire [7:0] add_955741;
  wire [7:0] sel_955742;
  wire [7:0] add_955745;
  wire [7:0] sel_955746;
  wire [7:0] add_955749;
  wire [7:0] sel_955750;
  wire [7:0] add_955753;
  wire [7:0] sel_955754;
  wire [7:0] add_955757;
  wire [7:0] sel_955758;
  wire [7:0] add_955761;
  wire [7:0] sel_955762;
  wire [7:0] add_955765;
  wire [7:0] sel_955766;
  wire [7:0] add_955769;
  wire [7:0] sel_955770;
  wire [7:0] add_955773;
  wire [7:0] sel_955774;
  wire [7:0] add_955777;
  wire [7:0] sel_955778;
  wire [7:0] add_955781;
  wire [7:0] sel_955782;
  wire [7:0] add_955785;
  wire [7:0] sel_955786;
  wire [7:0] add_955789;
  wire [7:0] sel_955790;
  wire [7:0] add_955793;
  wire [7:0] sel_955794;
  wire [7:0] add_955797;
  wire [7:0] sel_955798;
  wire [7:0] add_955801;
  wire [7:0] sel_955802;
  wire [7:0] add_955805;
  wire [7:0] sel_955806;
  wire [7:0] add_955809;
  wire [7:0] sel_955810;
  wire [7:0] add_955813;
  wire [7:0] sel_955814;
  wire [7:0] add_955817;
  wire [7:0] sel_955818;
  wire [7:0] add_955821;
  wire [7:0] sel_955822;
  wire [7:0] add_955825;
  wire [7:0] sel_955826;
  wire [7:0] add_955829;
  wire [7:0] sel_955830;
  wire [7:0] add_955833;
  wire [7:0] sel_955834;
  wire [7:0] add_955837;
  wire [7:0] sel_955838;
  wire [7:0] add_955841;
  wire [7:0] sel_955842;
  wire [7:0] add_955845;
  wire [7:0] sel_955846;
  wire [7:0] add_955849;
  wire [7:0] sel_955850;
  wire [7:0] add_955853;
  wire [7:0] sel_955854;
  wire [7:0] add_955857;
  wire [7:0] sel_955858;
  wire [7:0] add_955861;
  wire [7:0] sel_955862;
  wire [7:0] add_955865;
  wire [7:0] sel_955866;
  wire [7:0] add_955869;
  wire [7:0] sel_955870;
  wire [7:0] add_955873;
  wire [7:0] sel_955874;
  wire [7:0] add_955877;
  wire [7:0] sel_955878;
  wire [7:0] add_955881;
  wire [7:0] sel_955882;
  wire [7:0] add_955885;
  wire [7:0] sel_955886;
  wire [7:0] add_955889;
  wire [7:0] sel_955890;
  wire [7:0] add_955893;
  wire [7:0] sel_955894;
  wire [7:0] add_955897;
  wire [7:0] sel_955898;
  wire [7:0] add_955901;
  wire [7:0] sel_955902;
  wire [7:0] add_955905;
  wire [7:0] sel_955906;
  wire [7:0] add_955909;
  wire [7:0] sel_955910;
  wire [7:0] add_955913;
  wire [7:0] sel_955914;
  wire [7:0] add_955917;
  wire [7:0] sel_955918;
  wire [7:0] add_955921;
  wire [7:0] sel_955922;
  wire [7:0] add_955926;
  wire [15:0] array_index_955927;
  wire [7:0] sel_955928;
  wire [7:0] add_955931;
  wire [7:0] sel_955932;
  wire [7:0] add_955935;
  wire [7:0] sel_955936;
  wire [7:0] add_955939;
  wire [7:0] sel_955940;
  wire [7:0] add_955943;
  wire [7:0] sel_955944;
  wire [7:0] add_955947;
  wire [7:0] sel_955948;
  wire [7:0] add_955951;
  wire [7:0] sel_955952;
  wire [7:0] add_955955;
  wire [7:0] sel_955956;
  wire [7:0] add_955959;
  wire [7:0] sel_955960;
  wire [7:0] add_955963;
  wire [7:0] sel_955964;
  wire [7:0] add_955967;
  wire [7:0] sel_955968;
  wire [7:0] add_955971;
  wire [7:0] sel_955972;
  wire [7:0] add_955975;
  wire [7:0] sel_955976;
  wire [7:0] add_955979;
  wire [7:0] sel_955980;
  wire [7:0] add_955983;
  wire [7:0] sel_955984;
  wire [7:0] add_955987;
  wire [7:0] sel_955988;
  wire [7:0] add_955991;
  wire [7:0] sel_955992;
  wire [7:0] add_955995;
  wire [7:0] sel_955996;
  wire [7:0] add_955999;
  wire [7:0] sel_956000;
  wire [7:0] add_956003;
  wire [7:0] sel_956004;
  wire [7:0] add_956007;
  wire [7:0] sel_956008;
  wire [7:0] add_956011;
  wire [7:0] sel_956012;
  wire [7:0] add_956015;
  wire [7:0] sel_956016;
  wire [7:0] add_956019;
  wire [7:0] sel_956020;
  wire [7:0] add_956023;
  wire [7:0] sel_956024;
  wire [7:0] add_956027;
  wire [7:0] sel_956028;
  wire [7:0] add_956031;
  wire [7:0] sel_956032;
  wire [7:0] add_956035;
  wire [7:0] sel_956036;
  wire [7:0] add_956039;
  wire [7:0] sel_956040;
  wire [7:0] add_956043;
  wire [7:0] sel_956044;
  wire [7:0] add_956047;
  wire [7:0] sel_956048;
  wire [7:0] add_956051;
  wire [7:0] sel_956052;
  wire [7:0] add_956055;
  wire [7:0] sel_956056;
  wire [7:0] add_956059;
  wire [7:0] sel_956060;
  wire [7:0] add_956063;
  wire [7:0] sel_956064;
  wire [7:0] add_956067;
  wire [7:0] sel_956068;
  wire [7:0] add_956071;
  wire [7:0] sel_956072;
  wire [7:0] add_956075;
  wire [7:0] sel_956076;
  wire [7:0] add_956079;
  wire [7:0] sel_956080;
  wire [7:0] add_956083;
  wire [7:0] sel_956084;
  wire [7:0] add_956087;
  wire [7:0] sel_956088;
  wire [7:0] add_956091;
  wire [7:0] sel_956092;
  wire [7:0] add_956095;
  wire [7:0] sel_956096;
  wire [7:0] add_956099;
  wire [7:0] sel_956100;
  wire [7:0] add_956103;
  wire [7:0] sel_956104;
  wire [7:0] add_956107;
  wire [7:0] sel_956108;
  wire [7:0] add_956111;
  wire [7:0] sel_956112;
  wire [7:0] add_956115;
  wire [7:0] sel_956116;
  wire [7:0] add_956119;
  wire [7:0] sel_956120;
  wire [7:0] add_956123;
  wire [7:0] sel_956124;
  wire [7:0] add_956127;
  wire [7:0] sel_956128;
  wire [7:0] add_956131;
  wire [7:0] sel_956132;
  wire [7:0] add_956135;
  wire [7:0] sel_956136;
  wire [7:0] add_956139;
  wire [7:0] sel_956140;
  wire [7:0] add_956143;
  wire [7:0] sel_956144;
  wire [7:0] add_956147;
  wire [7:0] sel_956148;
  wire [7:0] add_956151;
  wire [7:0] sel_956152;
  wire [7:0] add_956155;
  wire [7:0] sel_956156;
  wire [7:0] add_956159;
  wire [7:0] sel_956160;
  wire [7:0] add_956163;
  wire [7:0] sel_956164;
  wire [7:0] add_956167;
  wire [7:0] sel_956168;
  wire [7:0] add_956171;
  wire [7:0] sel_956172;
  wire [7:0] add_956175;
  wire [7:0] sel_956176;
  wire [7:0] add_956179;
  wire [7:0] sel_956180;
  wire [7:0] add_956183;
  wire [7:0] sel_956184;
  wire [7:0] add_956187;
  wire [7:0] sel_956188;
  wire [7:0] add_956191;
  wire [7:0] sel_956192;
  wire [7:0] add_956195;
  wire [7:0] sel_956196;
  wire [7:0] add_956199;
  wire [7:0] sel_956200;
  wire [7:0] add_956203;
  wire [7:0] sel_956204;
  wire [7:0] add_956207;
  wire [7:0] sel_956208;
  wire [7:0] add_956211;
  wire [7:0] sel_956212;
  wire [7:0] add_956215;
  wire [7:0] sel_956216;
  wire [7:0] add_956219;
  wire [7:0] sel_956220;
  wire [7:0] add_956223;
  wire [7:0] sel_956224;
  wire [7:0] add_956227;
  wire [7:0] sel_956228;
  wire [7:0] add_956231;
  wire [7:0] sel_956232;
  wire [7:0] add_956235;
  wire [7:0] sel_956236;
  wire [7:0] add_956239;
  wire [7:0] sel_956240;
  wire [7:0] add_956243;
  wire [7:0] sel_956244;
  wire [7:0] add_956247;
  wire [7:0] sel_956248;
  wire [7:0] add_956251;
  wire [7:0] sel_956252;
  wire [7:0] add_956255;
  wire [7:0] sel_956256;
  wire [7:0] add_956259;
  wire [7:0] sel_956260;
  wire [7:0] add_956263;
  wire [7:0] sel_956264;
  wire [7:0] add_956267;
  wire [7:0] sel_956268;
  wire [7:0] add_956271;
  wire [7:0] sel_956272;
  wire [7:0] add_956275;
  wire [7:0] sel_956276;
  wire [7:0] add_956279;
  wire [7:0] sel_956280;
  wire [7:0] add_956283;
  wire [7:0] sel_956284;
  wire [7:0] add_956287;
  wire [7:0] sel_956288;
  wire [7:0] add_956291;
  wire [7:0] sel_956292;
  wire [7:0] add_956295;
  wire [7:0] sel_956296;
  wire [7:0] add_956299;
  wire [7:0] sel_956300;
  wire [7:0] add_956303;
  wire [7:0] sel_956304;
  wire [7:0] add_956307;
  wire [7:0] sel_956308;
  wire [7:0] add_956311;
  wire [7:0] sel_956312;
  wire [7:0] add_956315;
  wire [7:0] sel_956316;
  wire [7:0] add_956319;
  wire [7:0] sel_956320;
  wire [7:0] add_956323;
  wire [7:0] sel_956324;
  wire [7:0] add_956328;
  wire [15:0] array_index_956329;
  wire [7:0] sel_956330;
  wire [7:0] add_956333;
  wire [7:0] sel_956334;
  wire [7:0] add_956337;
  wire [7:0] sel_956338;
  wire [7:0] add_956341;
  wire [7:0] sel_956342;
  wire [7:0] add_956345;
  wire [7:0] sel_956346;
  wire [7:0] add_956349;
  wire [7:0] sel_956350;
  wire [7:0] add_956353;
  wire [7:0] sel_956354;
  wire [7:0] add_956357;
  wire [7:0] sel_956358;
  wire [7:0] add_956361;
  wire [7:0] sel_956362;
  wire [7:0] add_956365;
  wire [7:0] sel_956366;
  wire [7:0] add_956369;
  wire [7:0] sel_956370;
  wire [7:0] add_956373;
  wire [7:0] sel_956374;
  wire [7:0] add_956377;
  wire [7:0] sel_956378;
  wire [7:0] add_956381;
  wire [7:0] sel_956382;
  wire [7:0] add_956385;
  wire [7:0] sel_956386;
  wire [7:0] add_956389;
  wire [7:0] sel_956390;
  wire [7:0] add_956393;
  wire [7:0] sel_956394;
  wire [7:0] add_956397;
  wire [7:0] sel_956398;
  wire [7:0] add_956401;
  wire [7:0] sel_956402;
  wire [7:0] add_956405;
  wire [7:0] sel_956406;
  wire [7:0] add_956409;
  wire [7:0] sel_956410;
  wire [7:0] add_956413;
  wire [7:0] sel_956414;
  wire [7:0] add_956417;
  wire [7:0] sel_956418;
  wire [7:0] add_956421;
  wire [7:0] sel_956422;
  wire [7:0] add_956425;
  wire [7:0] sel_956426;
  wire [7:0] add_956429;
  wire [7:0] sel_956430;
  wire [7:0] add_956433;
  wire [7:0] sel_956434;
  wire [7:0] add_956437;
  wire [7:0] sel_956438;
  wire [7:0] add_956441;
  wire [7:0] sel_956442;
  wire [7:0] add_956445;
  wire [7:0] sel_956446;
  wire [7:0] add_956449;
  wire [7:0] sel_956450;
  wire [7:0] add_956453;
  wire [7:0] sel_956454;
  wire [7:0] add_956457;
  wire [7:0] sel_956458;
  wire [7:0] add_956461;
  wire [7:0] sel_956462;
  wire [7:0] add_956465;
  wire [7:0] sel_956466;
  wire [7:0] add_956469;
  wire [7:0] sel_956470;
  wire [7:0] add_956473;
  wire [7:0] sel_956474;
  wire [7:0] add_956477;
  wire [7:0] sel_956478;
  wire [7:0] add_956481;
  wire [7:0] sel_956482;
  wire [7:0] add_956485;
  wire [7:0] sel_956486;
  wire [7:0] add_956489;
  wire [7:0] sel_956490;
  wire [7:0] add_956493;
  wire [7:0] sel_956494;
  wire [7:0] add_956497;
  wire [7:0] sel_956498;
  wire [7:0] add_956501;
  wire [7:0] sel_956502;
  wire [7:0] add_956505;
  wire [7:0] sel_956506;
  wire [7:0] add_956509;
  wire [7:0] sel_956510;
  wire [7:0] add_956513;
  wire [7:0] sel_956514;
  wire [7:0] add_956517;
  wire [7:0] sel_956518;
  wire [7:0] add_956521;
  wire [7:0] sel_956522;
  wire [7:0] add_956525;
  wire [7:0] sel_956526;
  wire [7:0] add_956529;
  wire [7:0] sel_956530;
  wire [7:0] add_956533;
  wire [7:0] sel_956534;
  wire [7:0] add_956537;
  wire [7:0] sel_956538;
  wire [7:0] add_956541;
  wire [7:0] sel_956542;
  wire [7:0] add_956545;
  wire [7:0] sel_956546;
  wire [7:0] add_956549;
  wire [7:0] sel_956550;
  wire [7:0] add_956553;
  wire [7:0] sel_956554;
  wire [7:0] add_956557;
  wire [7:0] sel_956558;
  wire [7:0] add_956561;
  wire [7:0] sel_956562;
  wire [7:0] add_956565;
  wire [7:0] sel_956566;
  wire [7:0] add_956569;
  wire [7:0] sel_956570;
  wire [7:0] add_956573;
  wire [7:0] sel_956574;
  wire [7:0] add_956577;
  wire [7:0] sel_956578;
  wire [7:0] add_956581;
  wire [7:0] sel_956582;
  wire [7:0] add_956585;
  wire [7:0] sel_956586;
  wire [7:0] add_956589;
  wire [7:0] sel_956590;
  wire [7:0] add_956593;
  wire [7:0] sel_956594;
  wire [7:0] add_956597;
  wire [7:0] sel_956598;
  wire [7:0] add_956601;
  wire [7:0] sel_956602;
  wire [7:0] add_956605;
  wire [7:0] sel_956606;
  wire [7:0] add_956609;
  wire [7:0] sel_956610;
  wire [7:0] add_956613;
  wire [7:0] sel_956614;
  wire [7:0] add_956617;
  wire [7:0] sel_956618;
  wire [7:0] add_956621;
  wire [7:0] sel_956622;
  wire [7:0] add_956625;
  wire [7:0] sel_956626;
  wire [7:0] add_956629;
  wire [7:0] sel_956630;
  wire [7:0] add_956633;
  wire [7:0] sel_956634;
  wire [7:0] add_956637;
  wire [7:0] sel_956638;
  wire [7:0] add_956641;
  wire [7:0] sel_956642;
  wire [7:0] add_956645;
  wire [7:0] sel_956646;
  wire [7:0] add_956649;
  wire [7:0] sel_956650;
  wire [7:0] add_956653;
  wire [7:0] sel_956654;
  wire [7:0] add_956657;
  wire [7:0] sel_956658;
  wire [7:0] add_956661;
  wire [7:0] sel_956662;
  wire [7:0] add_956665;
  wire [7:0] sel_956666;
  wire [7:0] add_956669;
  wire [7:0] sel_956670;
  wire [7:0] add_956673;
  wire [7:0] sel_956674;
  wire [7:0] add_956677;
  wire [7:0] sel_956678;
  wire [7:0] add_956681;
  wire [7:0] sel_956682;
  wire [7:0] add_956685;
  wire [7:0] sel_956686;
  wire [7:0] add_956689;
  wire [7:0] sel_956690;
  wire [7:0] add_956693;
  wire [7:0] sel_956694;
  wire [7:0] add_956697;
  wire [7:0] sel_956698;
  wire [7:0] add_956701;
  wire [7:0] sel_956702;
  wire [7:0] add_956705;
  wire [7:0] sel_956706;
  wire [7:0] add_956709;
  wire [7:0] sel_956710;
  wire [7:0] add_956713;
  wire [7:0] sel_956714;
  wire [7:0] add_956717;
  wire [7:0] sel_956718;
  wire [7:0] add_956721;
  wire [7:0] sel_956722;
  wire [7:0] add_956725;
  wire [7:0] sel_956726;
  wire [7:0] add_956730;
  wire [15:0] array_index_956731;
  wire [7:0] sel_956732;
  wire [7:0] add_956735;
  wire [7:0] sel_956736;
  wire [7:0] add_956739;
  wire [7:0] sel_956740;
  wire [7:0] add_956743;
  wire [7:0] sel_956744;
  wire [7:0] add_956747;
  wire [7:0] sel_956748;
  wire [7:0] add_956751;
  wire [7:0] sel_956752;
  wire [7:0] add_956755;
  wire [7:0] sel_956756;
  wire [7:0] add_956759;
  wire [7:0] sel_956760;
  wire [7:0] add_956763;
  wire [7:0] sel_956764;
  wire [7:0] add_956767;
  wire [7:0] sel_956768;
  wire [7:0] add_956771;
  wire [7:0] sel_956772;
  wire [7:0] add_956775;
  wire [7:0] sel_956776;
  wire [7:0] add_956779;
  wire [7:0] sel_956780;
  wire [7:0] add_956783;
  wire [7:0] sel_956784;
  wire [7:0] add_956787;
  wire [7:0] sel_956788;
  wire [7:0] add_956791;
  wire [7:0] sel_956792;
  wire [7:0] add_956795;
  wire [7:0] sel_956796;
  wire [7:0] add_956799;
  wire [7:0] sel_956800;
  wire [7:0] add_956803;
  wire [7:0] sel_956804;
  wire [7:0] add_956807;
  wire [7:0] sel_956808;
  wire [7:0] add_956811;
  wire [7:0] sel_956812;
  wire [7:0] add_956815;
  wire [7:0] sel_956816;
  wire [7:0] add_956819;
  wire [7:0] sel_956820;
  wire [7:0] add_956823;
  wire [7:0] sel_956824;
  wire [7:0] add_956827;
  wire [7:0] sel_956828;
  wire [7:0] add_956831;
  wire [7:0] sel_956832;
  wire [7:0] add_956835;
  wire [7:0] sel_956836;
  wire [7:0] add_956839;
  wire [7:0] sel_956840;
  wire [7:0] add_956843;
  wire [7:0] sel_956844;
  wire [7:0] add_956847;
  wire [7:0] sel_956848;
  wire [7:0] add_956851;
  wire [7:0] sel_956852;
  wire [7:0] add_956855;
  wire [7:0] sel_956856;
  wire [7:0] add_956859;
  wire [7:0] sel_956860;
  wire [7:0] add_956863;
  wire [7:0] sel_956864;
  wire [7:0] add_956867;
  wire [7:0] sel_956868;
  wire [7:0] add_956871;
  wire [7:0] sel_956872;
  wire [7:0] add_956875;
  wire [7:0] sel_956876;
  wire [7:0] add_956879;
  wire [7:0] sel_956880;
  wire [7:0] add_956883;
  wire [7:0] sel_956884;
  wire [7:0] add_956887;
  wire [7:0] sel_956888;
  wire [7:0] add_956891;
  wire [7:0] sel_956892;
  wire [7:0] add_956895;
  wire [7:0] sel_956896;
  wire [7:0] add_956899;
  wire [7:0] sel_956900;
  wire [7:0] add_956903;
  wire [7:0] sel_956904;
  wire [7:0] add_956907;
  wire [7:0] sel_956908;
  wire [7:0] add_956911;
  wire [7:0] sel_956912;
  wire [7:0] add_956915;
  wire [7:0] sel_956916;
  wire [7:0] add_956919;
  wire [7:0] sel_956920;
  wire [7:0] add_956923;
  wire [7:0] sel_956924;
  wire [7:0] add_956927;
  wire [7:0] sel_956928;
  wire [7:0] add_956931;
  wire [7:0] sel_956932;
  wire [7:0] add_956935;
  wire [7:0] sel_956936;
  wire [7:0] add_956939;
  wire [7:0] sel_956940;
  wire [7:0] add_956943;
  wire [7:0] sel_956944;
  wire [7:0] add_956947;
  wire [7:0] sel_956948;
  wire [7:0] add_956951;
  wire [7:0] sel_956952;
  wire [7:0] add_956955;
  wire [7:0] sel_956956;
  wire [7:0] add_956959;
  wire [7:0] sel_956960;
  wire [7:0] add_956963;
  wire [7:0] sel_956964;
  wire [7:0] add_956967;
  wire [7:0] sel_956968;
  wire [7:0] add_956971;
  wire [7:0] sel_956972;
  wire [7:0] add_956975;
  wire [7:0] sel_956976;
  wire [7:0] add_956979;
  wire [7:0] sel_956980;
  wire [7:0] add_956983;
  wire [7:0] sel_956984;
  wire [7:0] add_956987;
  wire [7:0] sel_956988;
  wire [7:0] add_956991;
  wire [7:0] sel_956992;
  wire [7:0] add_956995;
  wire [7:0] sel_956996;
  wire [7:0] add_956999;
  wire [7:0] sel_957000;
  wire [7:0] add_957003;
  wire [7:0] sel_957004;
  wire [7:0] add_957007;
  wire [7:0] sel_957008;
  wire [7:0] add_957011;
  wire [7:0] sel_957012;
  wire [7:0] add_957015;
  wire [7:0] sel_957016;
  wire [7:0] add_957019;
  wire [7:0] sel_957020;
  wire [7:0] add_957023;
  wire [7:0] sel_957024;
  wire [7:0] add_957027;
  wire [7:0] sel_957028;
  wire [7:0] add_957031;
  wire [7:0] sel_957032;
  wire [7:0] add_957035;
  wire [7:0] sel_957036;
  wire [7:0] add_957039;
  wire [7:0] sel_957040;
  wire [7:0] add_957043;
  wire [7:0] sel_957044;
  wire [7:0] add_957047;
  wire [7:0] sel_957048;
  wire [7:0] add_957051;
  wire [7:0] sel_957052;
  wire [7:0] add_957055;
  wire [7:0] sel_957056;
  wire [7:0] add_957059;
  wire [7:0] sel_957060;
  wire [7:0] add_957063;
  wire [7:0] sel_957064;
  wire [7:0] add_957067;
  wire [7:0] sel_957068;
  wire [7:0] add_957071;
  wire [7:0] sel_957072;
  wire [7:0] add_957075;
  wire [7:0] sel_957076;
  wire [7:0] add_957079;
  wire [7:0] sel_957080;
  wire [7:0] add_957083;
  wire [7:0] sel_957084;
  wire [7:0] add_957087;
  wire [7:0] sel_957088;
  wire [7:0] add_957091;
  wire [7:0] sel_957092;
  wire [7:0] add_957095;
  wire [7:0] sel_957096;
  wire [7:0] add_957099;
  wire [7:0] sel_957100;
  wire [7:0] add_957103;
  wire [7:0] sel_957104;
  wire [7:0] add_957107;
  wire [7:0] sel_957108;
  wire [7:0] add_957111;
  wire [7:0] sel_957112;
  wire [7:0] add_957115;
  wire [7:0] sel_957116;
  wire [7:0] add_957119;
  wire [7:0] sel_957120;
  wire [7:0] add_957123;
  wire [7:0] sel_957124;
  wire [7:0] add_957127;
  wire [7:0] sel_957128;
  wire [7:0] add_957132;
  wire [15:0] array_index_957133;
  wire [7:0] sel_957134;
  wire [7:0] add_957137;
  wire [7:0] sel_957138;
  wire [7:0] add_957141;
  wire [7:0] sel_957142;
  wire [7:0] add_957145;
  wire [7:0] sel_957146;
  wire [7:0] add_957149;
  wire [7:0] sel_957150;
  wire [7:0] add_957153;
  wire [7:0] sel_957154;
  wire [7:0] add_957157;
  wire [7:0] sel_957158;
  wire [7:0] add_957161;
  wire [7:0] sel_957162;
  wire [7:0] add_957165;
  wire [7:0] sel_957166;
  wire [7:0] add_957169;
  wire [7:0] sel_957170;
  wire [7:0] add_957173;
  wire [7:0] sel_957174;
  wire [7:0] add_957177;
  wire [7:0] sel_957178;
  wire [7:0] add_957181;
  wire [7:0] sel_957182;
  wire [7:0] add_957185;
  wire [7:0] sel_957186;
  wire [7:0] add_957189;
  wire [7:0] sel_957190;
  wire [7:0] add_957193;
  wire [7:0] sel_957194;
  wire [7:0] add_957197;
  wire [7:0] sel_957198;
  wire [7:0] add_957201;
  wire [7:0] sel_957202;
  wire [7:0] add_957205;
  wire [7:0] sel_957206;
  wire [7:0] add_957209;
  wire [7:0] sel_957210;
  wire [7:0] add_957213;
  wire [7:0] sel_957214;
  wire [7:0] add_957217;
  wire [7:0] sel_957218;
  wire [7:0] add_957221;
  wire [7:0] sel_957222;
  wire [7:0] add_957225;
  wire [7:0] sel_957226;
  wire [7:0] add_957229;
  wire [7:0] sel_957230;
  wire [7:0] add_957233;
  wire [7:0] sel_957234;
  wire [7:0] add_957237;
  wire [7:0] sel_957238;
  wire [7:0] add_957241;
  wire [7:0] sel_957242;
  wire [7:0] add_957245;
  wire [7:0] sel_957246;
  wire [7:0] add_957249;
  wire [7:0] sel_957250;
  wire [7:0] add_957253;
  wire [7:0] sel_957254;
  wire [7:0] add_957257;
  wire [7:0] sel_957258;
  wire [7:0] add_957261;
  wire [7:0] sel_957262;
  wire [7:0] add_957265;
  wire [7:0] sel_957266;
  wire [7:0] add_957269;
  wire [7:0] sel_957270;
  wire [7:0] add_957273;
  wire [7:0] sel_957274;
  wire [7:0] add_957277;
  wire [7:0] sel_957278;
  wire [7:0] add_957281;
  wire [7:0] sel_957282;
  wire [7:0] add_957285;
  wire [7:0] sel_957286;
  wire [7:0] add_957289;
  wire [7:0] sel_957290;
  wire [7:0] add_957293;
  wire [7:0] sel_957294;
  wire [7:0] add_957297;
  wire [7:0] sel_957298;
  wire [7:0] add_957301;
  wire [7:0] sel_957302;
  wire [7:0] add_957305;
  wire [7:0] sel_957306;
  wire [7:0] add_957309;
  wire [7:0] sel_957310;
  wire [7:0] add_957313;
  wire [7:0] sel_957314;
  wire [7:0] add_957317;
  wire [7:0] sel_957318;
  wire [7:0] add_957321;
  wire [7:0] sel_957322;
  wire [7:0] add_957325;
  wire [7:0] sel_957326;
  wire [7:0] add_957329;
  wire [7:0] sel_957330;
  wire [7:0] add_957333;
  wire [7:0] sel_957334;
  wire [7:0] add_957337;
  wire [7:0] sel_957338;
  wire [7:0] add_957341;
  wire [7:0] sel_957342;
  wire [7:0] add_957345;
  wire [7:0] sel_957346;
  wire [7:0] add_957349;
  wire [7:0] sel_957350;
  wire [7:0] add_957353;
  wire [7:0] sel_957354;
  wire [7:0] add_957357;
  wire [7:0] sel_957358;
  wire [7:0] add_957361;
  wire [7:0] sel_957362;
  wire [7:0] add_957365;
  wire [7:0] sel_957366;
  wire [7:0] add_957369;
  wire [7:0] sel_957370;
  wire [7:0] add_957373;
  wire [7:0] sel_957374;
  wire [7:0] add_957377;
  wire [7:0] sel_957378;
  wire [7:0] add_957381;
  wire [7:0] sel_957382;
  wire [7:0] add_957385;
  wire [7:0] sel_957386;
  wire [7:0] add_957389;
  wire [7:0] sel_957390;
  wire [7:0] add_957393;
  wire [7:0] sel_957394;
  wire [7:0] add_957397;
  wire [7:0] sel_957398;
  wire [7:0] add_957401;
  wire [7:0] sel_957402;
  wire [7:0] add_957405;
  wire [7:0] sel_957406;
  wire [7:0] add_957409;
  wire [7:0] sel_957410;
  wire [7:0] add_957413;
  wire [7:0] sel_957414;
  wire [7:0] add_957417;
  wire [7:0] sel_957418;
  wire [7:0] add_957421;
  wire [7:0] sel_957422;
  wire [7:0] add_957425;
  wire [7:0] sel_957426;
  wire [7:0] add_957429;
  wire [7:0] sel_957430;
  wire [7:0] add_957433;
  wire [7:0] sel_957434;
  wire [7:0] add_957437;
  wire [7:0] sel_957438;
  wire [7:0] add_957441;
  wire [7:0] sel_957442;
  wire [7:0] add_957445;
  wire [7:0] sel_957446;
  wire [7:0] add_957449;
  wire [7:0] sel_957450;
  wire [7:0] add_957453;
  wire [7:0] sel_957454;
  wire [7:0] add_957457;
  wire [7:0] sel_957458;
  wire [7:0] add_957461;
  wire [7:0] sel_957462;
  wire [7:0] add_957465;
  wire [7:0] sel_957466;
  wire [7:0] add_957469;
  wire [7:0] sel_957470;
  wire [7:0] add_957473;
  wire [7:0] sel_957474;
  wire [7:0] add_957477;
  wire [7:0] sel_957478;
  wire [7:0] add_957481;
  wire [7:0] sel_957482;
  wire [7:0] add_957485;
  wire [7:0] sel_957486;
  wire [7:0] add_957489;
  wire [7:0] sel_957490;
  wire [7:0] add_957493;
  wire [7:0] sel_957494;
  wire [7:0] add_957497;
  wire [7:0] sel_957498;
  wire [7:0] add_957501;
  wire [7:0] sel_957502;
  wire [7:0] add_957505;
  wire [7:0] sel_957506;
  wire [7:0] add_957509;
  wire [7:0] sel_957510;
  wire [7:0] add_957513;
  wire [7:0] sel_957514;
  wire [7:0] add_957517;
  wire [7:0] sel_957518;
  wire [7:0] add_957521;
  wire [7:0] sel_957522;
  wire [7:0] add_957525;
  wire [7:0] sel_957526;
  wire [7:0] add_957529;
  wire [7:0] sel_957530;
  wire [7:0] add_957534;
  wire [15:0] array_index_957535;
  wire [7:0] sel_957536;
  wire [7:0] add_957539;
  wire [7:0] sel_957540;
  wire [7:0] add_957543;
  wire [7:0] sel_957544;
  wire [7:0] add_957547;
  wire [7:0] sel_957548;
  wire [7:0] add_957551;
  wire [7:0] sel_957552;
  wire [7:0] add_957555;
  wire [7:0] sel_957556;
  wire [7:0] add_957559;
  wire [7:0] sel_957560;
  wire [7:0] add_957563;
  wire [7:0] sel_957564;
  wire [7:0] add_957567;
  wire [7:0] sel_957568;
  wire [7:0] add_957571;
  wire [7:0] sel_957572;
  wire [7:0] add_957575;
  wire [7:0] sel_957576;
  wire [7:0] add_957579;
  wire [7:0] sel_957580;
  wire [7:0] add_957583;
  wire [7:0] sel_957584;
  wire [7:0] add_957587;
  wire [7:0] sel_957588;
  wire [7:0] add_957591;
  wire [7:0] sel_957592;
  wire [7:0] add_957595;
  wire [7:0] sel_957596;
  wire [7:0] add_957599;
  wire [7:0] sel_957600;
  wire [7:0] add_957603;
  wire [7:0] sel_957604;
  wire [7:0] add_957607;
  wire [7:0] sel_957608;
  wire [7:0] add_957611;
  wire [7:0] sel_957612;
  wire [7:0] add_957615;
  wire [7:0] sel_957616;
  wire [7:0] add_957619;
  wire [7:0] sel_957620;
  wire [7:0] add_957623;
  wire [7:0] sel_957624;
  wire [7:0] add_957627;
  wire [7:0] sel_957628;
  wire [7:0] add_957631;
  wire [7:0] sel_957632;
  wire [7:0] add_957635;
  wire [7:0] sel_957636;
  wire [7:0] add_957639;
  wire [7:0] sel_957640;
  wire [7:0] add_957643;
  wire [7:0] sel_957644;
  wire [7:0] add_957647;
  wire [7:0] sel_957648;
  wire [7:0] add_957651;
  wire [7:0] sel_957652;
  wire [7:0] add_957655;
  wire [7:0] sel_957656;
  wire [7:0] add_957659;
  wire [7:0] sel_957660;
  wire [7:0] add_957663;
  wire [7:0] sel_957664;
  wire [7:0] add_957667;
  wire [7:0] sel_957668;
  wire [7:0] add_957671;
  wire [7:0] sel_957672;
  wire [7:0] add_957675;
  wire [7:0] sel_957676;
  wire [7:0] add_957679;
  wire [7:0] sel_957680;
  wire [7:0] add_957683;
  wire [7:0] sel_957684;
  wire [7:0] add_957687;
  wire [7:0] sel_957688;
  wire [7:0] add_957691;
  wire [7:0] sel_957692;
  wire [7:0] add_957695;
  wire [7:0] sel_957696;
  wire [7:0] add_957699;
  wire [7:0] sel_957700;
  wire [7:0] add_957703;
  wire [7:0] sel_957704;
  wire [7:0] add_957707;
  wire [7:0] sel_957708;
  wire [7:0] add_957711;
  wire [7:0] sel_957712;
  wire [7:0] add_957715;
  wire [7:0] sel_957716;
  wire [7:0] add_957719;
  wire [7:0] sel_957720;
  wire [7:0] add_957723;
  wire [7:0] sel_957724;
  wire [7:0] add_957727;
  wire [7:0] sel_957728;
  wire [7:0] add_957731;
  wire [7:0] sel_957732;
  wire [7:0] add_957735;
  wire [7:0] sel_957736;
  wire [7:0] add_957739;
  wire [7:0] sel_957740;
  wire [7:0] add_957743;
  wire [7:0] sel_957744;
  wire [7:0] add_957747;
  wire [7:0] sel_957748;
  wire [7:0] add_957751;
  wire [7:0] sel_957752;
  wire [7:0] add_957755;
  wire [7:0] sel_957756;
  wire [7:0] add_957759;
  wire [7:0] sel_957760;
  wire [7:0] add_957763;
  wire [7:0] sel_957764;
  wire [7:0] add_957767;
  wire [7:0] sel_957768;
  wire [7:0] add_957771;
  wire [7:0] sel_957772;
  wire [7:0] add_957775;
  wire [7:0] sel_957776;
  wire [7:0] add_957779;
  wire [7:0] sel_957780;
  wire [7:0] add_957783;
  wire [7:0] sel_957784;
  wire [7:0] add_957787;
  wire [7:0] sel_957788;
  wire [7:0] add_957791;
  wire [7:0] sel_957792;
  wire [7:0] add_957795;
  wire [7:0] sel_957796;
  wire [7:0] add_957799;
  wire [7:0] sel_957800;
  wire [7:0] add_957803;
  wire [7:0] sel_957804;
  wire [7:0] add_957807;
  wire [7:0] sel_957808;
  wire [7:0] add_957811;
  wire [7:0] sel_957812;
  wire [7:0] add_957815;
  wire [7:0] sel_957816;
  wire [7:0] add_957819;
  wire [7:0] sel_957820;
  wire [7:0] add_957823;
  wire [7:0] sel_957824;
  wire [7:0] add_957827;
  wire [7:0] sel_957828;
  wire [7:0] add_957831;
  wire [7:0] sel_957832;
  wire [7:0] add_957835;
  wire [7:0] sel_957836;
  wire [7:0] add_957839;
  wire [7:0] sel_957840;
  wire [7:0] add_957843;
  wire [7:0] sel_957844;
  wire [7:0] add_957847;
  wire [7:0] sel_957848;
  wire [7:0] add_957851;
  wire [7:0] sel_957852;
  wire [7:0] add_957855;
  wire [7:0] sel_957856;
  wire [7:0] add_957859;
  wire [7:0] sel_957860;
  wire [7:0] add_957863;
  wire [7:0] sel_957864;
  wire [7:0] add_957867;
  wire [7:0] sel_957868;
  wire [7:0] add_957871;
  wire [7:0] sel_957872;
  wire [7:0] add_957875;
  wire [7:0] sel_957876;
  wire [7:0] add_957879;
  wire [7:0] sel_957880;
  wire [7:0] add_957883;
  wire [7:0] sel_957884;
  wire [7:0] add_957887;
  wire [7:0] sel_957888;
  wire [7:0] add_957891;
  wire [7:0] sel_957892;
  wire [7:0] add_957895;
  wire [7:0] sel_957896;
  wire [7:0] add_957899;
  wire [7:0] sel_957900;
  wire [7:0] add_957903;
  wire [7:0] sel_957904;
  wire [7:0] add_957907;
  wire [7:0] sel_957908;
  wire [7:0] add_957911;
  wire [7:0] sel_957912;
  wire [7:0] add_957915;
  wire [7:0] sel_957916;
  wire [7:0] add_957919;
  wire [7:0] sel_957920;
  wire [7:0] add_957923;
  wire [7:0] sel_957924;
  wire [7:0] add_957927;
  wire [7:0] sel_957928;
  wire [7:0] add_957931;
  wire [7:0] sel_957932;
  wire [7:0] add_957936;
  wire [15:0] array_index_957937;
  wire [7:0] sel_957938;
  wire [7:0] add_957941;
  wire [7:0] sel_957942;
  wire [7:0] add_957945;
  wire [7:0] sel_957946;
  wire [7:0] add_957949;
  wire [7:0] sel_957950;
  wire [7:0] add_957953;
  wire [7:0] sel_957954;
  wire [7:0] add_957957;
  wire [7:0] sel_957958;
  wire [7:0] add_957961;
  wire [7:0] sel_957962;
  wire [7:0] add_957965;
  wire [7:0] sel_957966;
  wire [7:0] add_957969;
  wire [7:0] sel_957970;
  wire [7:0] add_957973;
  wire [7:0] sel_957974;
  wire [7:0] add_957977;
  wire [7:0] sel_957978;
  wire [7:0] add_957981;
  wire [7:0] sel_957982;
  wire [7:0] add_957985;
  wire [7:0] sel_957986;
  wire [7:0] add_957989;
  wire [7:0] sel_957990;
  wire [7:0] add_957993;
  wire [7:0] sel_957994;
  wire [7:0] add_957997;
  wire [7:0] sel_957998;
  wire [7:0] add_958001;
  wire [7:0] sel_958002;
  wire [7:0] add_958005;
  wire [7:0] sel_958006;
  wire [7:0] add_958009;
  wire [7:0] sel_958010;
  wire [7:0] add_958013;
  wire [7:0] sel_958014;
  wire [7:0] add_958017;
  wire [7:0] sel_958018;
  wire [7:0] add_958021;
  wire [7:0] sel_958022;
  wire [7:0] add_958025;
  wire [7:0] sel_958026;
  wire [7:0] add_958029;
  wire [7:0] sel_958030;
  wire [7:0] add_958033;
  wire [7:0] sel_958034;
  wire [7:0] add_958037;
  wire [7:0] sel_958038;
  wire [7:0] add_958041;
  wire [7:0] sel_958042;
  wire [7:0] add_958045;
  wire [7:0] sel_958046;
  wire [7:0] add_958049;
  wire [7:0] sel_958050;
  wire [7:0] add_958053;
  wire [7:0] sel_958054;
  wire [7:0] add_958057;
  wire [7:0] sel_958058;
  wire [7:0] add_958061;
  wire [7:0] sel_958062;
  wire [7:0] add_958065;
  wire [7:0] sel_958066;
  wire [7:0] add_958069;
  wire [7:0] sel_958070;
  wire [7:0] add_958073;
  wire [7:0] sel_958074;
  wire [7:0] add_958077;
  wire [7:0] sel_958078;
  wire [7:0] add_958081;
  wire [7:0] sel_958082;
  wire [7:0] add_958085;
  wire [7:0] sel_958086;
  wire [7:0] add_958089;
  wire [7:0] sel_958090;
  wire [7:0] add_958093;
  wire [7:0] sel_958094;
  wire [7:0] add_958097;
  wire [7:0] sel_958098;
  wire [7:0] add_958101;
  wire [7:0] sel_958102;
  wire [7:0] add_958105;
  wire [7:0] sel_958106;
  wire [7:0] add_958109;
  wire [7:0] sel_958110;
  wire [7:0] add_958113;
  wire [7:0] sel_958114;
  wire [7:0] add_958117;
  wire [7:0] sel_958118;
  wire [7:0] add_958121;
  wire [7:0] sel_958122;
  wire [7:0] add_958125;
  wire [7:0] sel_958126;
  wire [7:0] add_958129;
  wire [7:0] sel_958130;
  wire [7:0] add_958133;
  wire [7:0] sel_958134;
  wire [7:0] add_958137;
  wire [7:0] sel_958138;
  wire [7:0] add_958141;
  wire [7:0] sel_958142;
  wire [7:0] add_958145;
  wire [7:0] sel_958146;
  wire [7:0] add_958149;
  wire [7:0] sel_958150;
  wire [7:0] add_958153;
  wire [7:0] sel_958154;
  wire [7:0] add_958157;
  wire [7:0] sel_958158;
  wire [7:0] add_958161;
  wire [7:0] sel_958162;
  wire [7:0] add_958165;
  wire [7:0] sel_958166;
  wire [7:0] add_958169;
  wire [7:0] sel_958170;
  wire [7:0] add_958173;
  wire [7:0] sel_958174;
  wire [7:0] add_958177;
  wire [7:0] sel_958178;
  wire [7:0] add_958181;
  wire [7:0] sel_958182;
  wire [7:0] add_958185;
  wire [7:0] sel_958186;
  wire [7:0] add_958189;
  wire [7:0] sel_958190;
  wire [7:0] add_958193;
  wire [7:0] sel_958194;
  wire [7:0] add_958197;
  wire [7:0] sel_958198;
  wire [7:0] add_958201;
  wire [7:0] sel_958202;
  wire [7:0] add_958205;
  wire [7:0] sel_958206;
  wire [7:0] add_958209;
  wire [7:0] sel_958210;
  wire [7:0] add_958213;
  wire [7:0] sel_958214;
  wire [7:0] add_958217;
  wire [7:0] sel_958218;
  wire [7:0] add_958221;
  wire [7:0] sel_958222;
  wire [7:0] add_958225;
  wire [7:0] sel_958226;
  wire [7:0] add_958229;
  wire [7:0] sel_958230;
  wire [7:0] add_958233;
  wire [7:0] sel_958234;
  wire [7:0] add_958237;
  wire [7:0] sel_958238;
  wire [7:0] add_958241;
  wire [7:0] sel_958242;
  wire [7:0] add_958245;
  wire [7:0] sel_958246;
  wire [7:0] add_958249;
  wire [7:0] sel_958250;
  wire [7:0] add_958253;
  wire [7:0] sel_958254;
  wire [7:0] add_958257;
  wire [7:0] sel_958258;
  wire [7:0] add_958261;
  wire [7:0] sel_958262;
  wire [7:0] add_958265;
  wire [7:0] sel_958266;
  wire [7:0] add_958269;
  wire [7:0] sel_958270;
  wire [7:0] add_958273;
  wire [7:0] sel_958274;
  wire [7:0] add_958277;
  wire [7:0] sel_958278;
  wire [7:0] add_958281;
  wire [7:0] sel_958282;
  wire [7:0] add_958285;
  wire [7:0] sel_958286;
  wire [7:0] add_958289;
  wire [7:0] sel_958290;
  wire [7:0] add_958293;
  wire [7:0] sel_958294;
  wire [7:0] add_958297;
  wire [7:0] sel_958298;
  wire [7:0] add_958301;
  wire [7:0] sel_958302;
  wire [7:0] add_958305;
  wire [7:0] sel_958306;
  wire [7:0] add_958309;
  wire [7:0] sel_958310;
  wire [7:0] add_958313;
  wire [7:0] sel_958314;
  wire [7:0] add_958317;
  wire [7:0] sel_958318;
  wire [7:0] add_958321;
  wire [7:0] sel_958322;
  wire [7:0] add_958325;
  wire [7:0] sel_958326;
  wire [7:0] add_958329;
  wire [7:0] sel_958330;
  wire [7:0] add_958333;
  wire [7:0] sel_958334;
  wire [7:0] add_958338;
  wire [15:0] array_index_958339;
  wire [7:0] sel_958340;
  wire [7:0] add_958343;
  wire [7:0] sel_958344;
  wire [7:0] add_958347;
  wire [7:0] sel_958348;
  wire [7:0] add_958351;
  wire [7:0] sel_958352;
  wire [7:0] add_958355;
  wire [7:0] sel_958356;
  wire [7:0] add_958359;
  wire [7:0] sel_958360;
  wire [7:0] add_958363;
  wire [7:0] sel_958364;
  wire [7:0] add_958367;
  wire [7:0] sel_958368;
  wire [7:0] add_958371;
  wire [7:0] sel_958372;
  wire [7:0] add_958375;
  wire [7:0] sel_958376;
  wire [7:0] add_958379;
  wire [7:0] sel_958380;
  wire [7:0] add_958383;
  wire [7:0] sel_958384;
  wire [7:0] add_958387;
  wire [7:0] sel_958388;
  wire [7:0] add_958391;
  wire [7:0] sel_958392;
  wire [7:0] add_958395;
  wire [7:0] sel_958396;
  wire [7:0] add_958399;
  wire [7:0] sel_958400;
  wire [7:0] add_958403;
  wire [7:0] sel_958404;
  wire [7:0] add_958407;
  wire [7:0] sel_958408;
  wire [7:0] add_958411;
  wire [7:0] sel_958412;
  wire [7:0] add_958415;
  wire [7:0] sel_958416;
  wire [7:0] add_958419;
  wire [7:0] sel_958420;
  wire [7:0] add_958423;
  wire [7:0] sel_958424;
  wire [7:0] add_958427;
  wire [7:0] sel_958428;
  wire [7:0] add_958431;
  wire [7:0] sel_958432;
  wire [7:0] add_958435;
  wire [7:0] sel_958436;
  wire [7:0] add_958439;
  wire [7:0] sel_958440;
  wire [7:0] add_958443;
  wire [7:0] sel_958444;
  wire [7:0] add_958447;
  wire [7:0] sel_958448;
  wire [7:0] add_958451;
  wire [7:0] sel_958452;
  wire [7:0] add_958455;
  wire [7:0] sel_958456;
  wire [7:0] add_958459;
  wire [7:0] sel_958460;
  wire [7:0] add_958463;
  wire [7:0] sel_958464;
  wire [7:0] add_958467;
  wire [7:0] sel_958468;
  wire [7:0] add_958471;
  wire [7:0] sel_958472;
  wire [7:0] add_958475;
  wire [7:0] sel_958476;
  wire [7:0] add_958479;
  wire [7:0] sel_958480;
  wire [7:0] add_958483;
  wire [7:0] sel_958484;
  wire [7:0] add_958487;
  wire [7:0] sel_958488;
  wire [7:0] add_958491;
  wire [7:0] sel_958492;
  wire [7:0] add_958495;
  wire [7:0] sel_958496;
  wire [7:0] add_958499;
  wire [7:0] sel_958500;
  wire [7:0] add_958503;
  wire [7:0] sel_958504;
  wire [7:0] add_958507;
  wire [7:0] sel_958508;
  wire [7:0] add_958511;
  wire [7:0] sel_958512;
  wire [7:0] add_958515;
  wire [7:0] sel_958516;
  wire [7:0] add_958519;
  wire [7:0] sel_958520;
  wire [7:0] add_958523;
  wire [7:0] sel_958524;
  wire [7:0] add_958527;
  wire [7:0] sel_958528;
  wire [7:0] add_958531;
  wire [7:0] sel_958532;
  wire [7:0] add_958535;
  wire [7:0] sel_958536;
  wire [7:0] add_958539;
  wire [7:0] sel_958540;
  wire [7:0] add_958543;
  wire [7:0] sel_958544;
  wire [7:0] add_958547;
  wire [7:0] sel_958548;
  wire [7:0] add_958551;
  wire [7:0] sel_958552;
  wire [7:0] add_958555;
  wire [7:0] sel_958556;
  wire [7:0] add_958559;
  wire [7:0] sel_958560;
  wire [7:0] add_958563;
  wire [7:0] sel_958564;
  wire [7:0] add_958567;
  wire [7:0] sel_958568;
  wire [7:0] add_958571;
  wire [7:0] sel_958572;
  wire [7:0] add_958575;
  wire [7:0] sel_958576;
  wire [7:0] add_958579;
  wire [7:0] sel_958580;
  wire [7:0] add_958583;
  wire [7:0] sel_958584;
  wire [7:0] add_958587;
  wire [7:0] sel_958588;
  wire [7:0] add_958591;
  wire [7:0] sel_958592;
  wire [7:0] add_958595;
  wire [7:0] sel_958596;
  wire [7:0] add_958599;
  wire [7:0] sel_958600;
  wire [7:0] add_958603;
  wire [7:0] sel_958604;
  wire [7:0] add_958607;
  wire [7:0] sel_958608;
  wire [7:0] add_958611;
  wire [7:0] sel_958612;
  wire [7:0] add_958615;
  wire [7:0] sel_958616;
  wire [7:0] add_958619;
  wire [7:0] sel_958620;
  wire [7:0] add_958623;
  wire [7:0] sel_958624;
  wire [7:0] add_958627;
  wire [7:0] sel_958628;
  wire [7:0] add_958631;
  wire [7:0] sel_958632;
  wire [7:0] add_958635;
  wire [7:0] sel_958636;
  wire [7:0] add_958639;
  wire [7:0] sel_958640;
  wire [7:0] add_958643;
  wire [7:0] sel_958644;
  wire [7:0] add_958647;
  wire [7:0] sel_958648;
  wire [7:0] add_958651;
  wire [7:0] sel_958652;
  wire [7:0] add_958655;
  wire [7:0] sel_958656;
  wire [7:0] add_958659;
  wire [7:0] sel_958660;
  wire [7:0] add_958663;
  wire [7:0] sel_958664;
  wire [7:0] add_958667;
  wire [7:0] sel_958668;
  wire [7:0] add_958671;
  wire [7:0] sel_958672;
  wire [7:0] add_958675;
  wire [7:0] sel_958676;
  wire [7:0] add_958679;
  wire [7:0] sel_958680;
  wire [7:0] add_958683;
  wire [7:0] sel_958684;
  wire [7:0] add_958687;
  wire [7:0] sel_958688;
  wire [7:0] add_958691;
  wire [7:0] sel_958692;
  wire [7:0] add_958695;
  wire [7:0] sel_958696;
  wire [7:0] add_958699;
  wire [7:0] sel_958700;
  wire [7:0] add_958703;
  wire [7:0] sel_958704;
  wire [7:0] add_958707;
  wire [7:0] sel_958708;
  wire [7:0] add_958711;
  wire [7:0] sel_958712;
  wire [7:0] add_958715;
  wire [7:0] sel_958716;
  wire [7:0] add_958719;
  wire [7:0] sel_958720;
  wire [7:0] add_958723;
  wire [7:0] sel_958724;
  wire [7:0] add_958727;
  wire [7:0] sel_958728;
  wire [7:0] add_958731;
  wire [7:0] sel_958732;
  wire [7:0] add_958735;
  wire [7:0] sel_958736;
  wire [7:0] add_958740;
  wire [15:0] array_index_958741;
  wire [7:0] sel_958742;
  wire [7:0] add_958745;
  wire [7:0] sel_958746;
  wire [7:0] add_958749;
  wire [7:0] sel_958750;
  wire [7:0] add_958753;
  wire [7:0] sel_958754;
  wire [7:0] add_958757;
  wire [7:0] sel_958758;
  wire [7:0] add_958761;
  wire [7:0] sel_958762;
  wire [7:0] add_958765;
  wire [7:0] sel_958766;
  wire [7:0] add_958769;
  wire [7:0] sel_958770;
  wire [7:0] add_958773;
  wire [7:0] sel_958774;
  wire [7:0] add_958777;
  wire [7:0] sel_958778;
  wire [7:0] add_958781;
  wire [7:0] sel_958782;
  wire [7:0] add_958785;
  wire [7:0] sel_958786;
  wire [7:0] add_958789;
  wire [7:0] sel_958790;
  wire [7:0] add_958793;
  wire [7:0] sel_958794;
  wire [7:0] add_958797;
  wire [7:0] sel_958798;
  wire [7:0] add_958801;
  wire [7:0] sel_958802;
  wire [7:0] add_958805;
  wire [7:0] sel_958806;
  wire [7:0] add_958809;
  wire [7:0] sel_958810;
  wire [7:0] add_958813;
  wire [7:0] sel_958814;
  wire [7:0] add_958817;
  wire [7:0] sel_958818;
  wire [7:0] add_958821;
  wire [7:0] sel_958822;
  wire [7:0] add_958825;
  wire [7:0] sel_958826;
  wire [7:0] add_958829;
  wire [7:0] sel_958830;
  wire [7:0] add_958833;
  wire [7:0] sel_958834;
  wire [7:0] add_958837;
  wire [7:0] sel_958838;
  wire [7:0] add_958841;
  wire [7:0] sel_958842;
  wire [7:0] add_958845;
  wire [7:0] sel_958846;
  wire [7:0] add_958849;
  wire [7:0] sel_958850;
  wire [7:0] add_958853;
  wire [7:0] sel_958854;
  wire [7:0] add_958857;
  wire [7:0] sel_958858;
  wire [7:0] add_958861;
  wire [7:0] sel_958862;
  wire [7:0] add_958865;
  wire [7:0] sel_958866;
  wire [7:0] add_958869;
  wire [7:0] sel_958870;
  wire [7:0] add_958873;
  wire [7:0] sel_958874;
  wire [7:0] add_958877;
  wire [7:0] sel_958878;
  wire [7:0] add_958881;
  wire [7:0] sel_958882;
  wire [7:0] add_958885;
  wire [7:0] sel_958886;
  wire [7:0] add_958889;
  wire [7:0] sel_958890;
  wire [7:0] add_958893;
  wire [7:0] sel_958894;
  wire [7:0] add_958897;
  wire [7:0] sel_958898;
  wire [7:0] add_958901;
  wire [7:0] sel_958902;
  wire [7:0] add_958905;
  wire [7:0] sel_958906;
  wire [7:0] add_958909;
  wire [7:0] sel_958910;
  wire [7:0] add_958913;
  wire [7:0] sel_958914;
  wire [7:0] add_958917;
  wire [7:0] sel_958918;
  wire [7:0] add_958921;
  wire [7:0] sel_958922;
  wire [7:0] add_958925;
  wire [7:0] sel_958926;
  wire [7:0] add_958929;
  wire [7:0] sel_958930;
  wire [7:0] add_958933;
  wire [7:0] sel_958934;
  wire [7:0] add_958937;
  wire [7:0] sel_958938;
  wire [7:0] add_958941;
  wire [7:0] sel_958942;
  wire [7:0] add_958945;
  wire [7:0] sel_958946;
  wire [7:0] add_958949;
  wire [7:0] sel_958950;
  wire [7:0] add_958953;
  wire [7:0] sel_958954;
  wire [7:0] add_958957;
  wire [7:0] sel_958958;
  wire [7:0] add_958961;
  wire [7:0] sel_958962;
  wire [7:0] add_958965;
  wire [7:0] sel_958966;
  wire [7:0] add_958969;
  wire [7:0] sel_958970;
  wire [7:0] add_958973;
  wire [7:0] sel_958974;
  wire [7:0] add_958977;
  wire [7:0] sel_958978;
  wire [7:0] add_958981;
  wire [7:0] sel_958982;
  wire [7:0] add_958985;
  wire [7:0] sel_958986;
  wire [7:0] add_958989;
  wire [7:0] sel_958990;
  wire [7:0] add_958993;
  wire [7:0] sel_958994;
  wire [7:0] add_958997;
  wire [7:0] sel_958998;
  wire [7:0] add_959001;
  wire [7:0] sel_959002;
  wire [7:0] add_959005;
  wire [7:0] sel_959006;
  wire [7:0] add_959009;
  wire [7:0] sel_959010;
  wire [7:0] add_959013;
  wire [7:0] sel_959014;
  wire [7:0] add_959017;
  wire [7:0] sel_959018;
  wire [7:0] add_959021;
  wire [7:0] sel_959022;
  wire [7:0] add_959025;
  wire [7:0] sel_959026;
  wire [7:0] add_959029;
  wire [7:0] sel_959030;
  wire [7:0] add_959033;
  wire [7:0] sel_959034;
  wire [7:0] add_959037;
  wire [7:0] sel_959038;
  wire [7:0] add_959041;
  wire [7:0] sel_959042;
  wire [7:0] add_959045;
  wire [7:0] sel_959046;
  wire [7:0] add_959049;
  wire [7:0] sel_959050;
  wire [7:0] add_959053;
  wire [7:0] sel_959054;
  wire [7:0] add_959057;
  wire [7:0] sel_959058;
  wire [7:0] add_959061;
  wire [7:0] sel_959062;
  wire [7:0] add_959065;
  wire [7:0] sel_959066;
  wire [7:0] add_959069;
  wire [7:0] sel_959070;
  wire [7:0] add_959073;
  wire [7:0] sel_959074;
  wire [7:0] add_959077;
  wire [7:0] sel_959078;
  wire [7:0] add_959081;
  wire [7:0] sel_959082;
  wire [7:0] add_959085;
  wire [7:0] sel_959086;
  wire [7:0] add_959089;
  wire [7:0] sel_959090;
  wire [7:0] add_959093;
  wire [7:0] sel_959094;
  wire [7:0] add_959097;
  wire [7:0] sel_959098;
  wire [7:0] add_959101;
  wire [7:0] sel_959102;
  wire [7:0] add_959105;
  wire [7:0] sel_959106;
  wire [7:0] add_959109;
  wire [7:0] sel_959110;
  wire [7:0] add_959113;
  wire [7:0] sel_959114;
  wire [7:0] add_959117;
  wire [7:0] sel_959118;
  wire [7:0] add_959121;
  wire [7:0] sel_959122;
  wire [7:0] add_959125;
  wire [7:0] sel_959126;
  wire [7:0] add_959129;
  wire [7:0] sel_959130;
  wire [7:0] add_959133;
  wire [7:0] sel_959134;
  wire [7:0] add_959137;
  wire [7:0] sel_959138;
  wire [7:0] add_959142;
  wire [15:0] array_index_959143;
  wire [7:0] sel_959144;
  wire [7:0] add_959147;
  wire [7:0] sel_959148;
  wire [7:0] add_959151;
  wire [7:0] sel_959152;
  wire [7:0] add_959155;
  wire [7:0] sel_959156;
  wire [7:0] add_959159;
  wire [7:0] sel_959160;
  wire [7:0] add_959163;
  wire [7:0] sel_959164;
  wire [7:0] add_959167;
  wire [7:0] sel_959168;
  wire [7:0] add_959171;
  wire [7:0] sel_959172;
  wire [7:0] add_959175;
  wire [7:0] sel_959176;
  wire [7:0] add_959179;
  wire [7:0] sel_959180;
  wire [7:0] add_959183;
  wire [7:0] sel_959184;
  wire [7:0] add_959187;
  wire [7:0] sel_959188;
  wire [7:0] add_959191;
  wire [7:0] sel_959192;
  wire [7:0] add_959195;
  wire [7:0] sel_959196;
  wire [7:0] add_959199;
  wire [7:0] sel_959200;
  wire [7:0] add_959203;
  wire [7:0] sel_959204;
  wire [7:0] add_959207;
  wire [7:0] sel_959208;
  wire [7:0] add_959211;
  wire [7:0] sel_959212;
  wire [7:0] add_959215;
  wire [7:0] sel_959216;
  wire [7:0] add_959219;
  wire [7:0] sel_959220;
  wire [7:0] add_959223;
  wire [7:0] sel_959224;
  wire [7:0] add_959227;
  wire [7:0] sel_959228;
  wire [7:0] add_959231;
  wire [7:0] sel_959232;
  wire [7:0] add_959235;
  wire [7:0] sel_959236;
  wire [7:0] add_959239;
  wire [7:0] sel_959240;
  wire [7:0] add_959243;
  wire [7:0] sel_959244;
  wire [7:0] add_959247;
  wire [7:0] sel_959248;
  wire [7:0] add_959251;
  wire [7:0] sel_959252;
  wire [7:0] add_959255;
  wire [7:0] sel_959256;
  wire [7:0] add_959259;
  wire [7:0] sel_959260;
  wire [7:0] add_959263;
  wire [7:0] sel_959264;
  wire [7:0] add_959267;
  wire [7:0] sel_959268;
  wire [7:0] add_959271;
  wire [7:0] sel_959272;
  wire [7:0] add_959275;
  wire [7:0] sel_959276;
  wire [7:0] add_959279;
  wire [7:0] sel_959280;
  wire [7:0] add_959283;
  wire [7:0] sel_959284;
  wire [7:0] add_959287;
  wire [7:0] sel_959288;
  wire [7:0] add_959291;
  wire [7:0] sel_959292;
  wire [7:0] add_959295;
  wire [7:0] sel_959296;
  wire [7:0] add_959299;
  wire [7:0] sel_959300;
  wire [7:0] add_959303;
  wire [7:0] sel_959304;
  wire [7:0] add_959307;
  wire [7:0] sel_959308;
  wire [7:0] add_959311;
  wire [7:0] sel_959312;
  wire [7:0] add_959315;
  wire [7:0] sel_959316;
  wire [7:0] add_959319;
  wire [7:0] sel_959320;
  wire [7:0] add_959323;
  wire [7:0] sel_959324;
  wire [7:0] add_959327;
  wire [7:0] sel_959328;
  wire [7:0] add_959331;
  wire [7:0] sel_959332;
  wire [7:0] add_959335;
  wire [7:0] sel_959336;
  wire [7:0] add_959339;
  wire [7:0] sel_959340;
  wire [7:0] add_959343;
  wire [7:0] sel_959344;
  wire [7:0] add_959347;
  wire [7:0] sel_959348;
  wire [7:0] add_959351;
  wire [7:0] sel_959352;
  wire [7:0] add_959355;
  wire [7:0] sel_959356;
  wire [7:0] add_959359;
  wire [7:0] sel_959360;
  wire [7:0] add_959363;
  wire [7:0] sel_959364;
  wire [7:0] add_959367;
  wire [7:0] sel_959368;
  wire [7:0] add_959371;
  wire [7:0] sel_959372;
  wire [7:0] add_959375;
  wire [7:0] sel_959376;
  wire [7:0] add_959379;
  wire [7:0] sel_959380;
  wire [7:0] add_959383;
  wire [7:0] sel_959384;
  wire [7:0] add_959387;
  wire [7:0] sel_959388;
  wire [7:0] add_959391;
  wire [7:0] sel_959392;
  wire [7:0] add_959395;
  wire [7:0] sel_959396;
  wire [7:0] add_959399;
  wire [7:0] sel_959400;
  wire [7:0] add_959403;
  wire [7:0] sel_959404;
  wire [7:0] add_959407;
  wire [7:0] sel_959408;
  wire [7:0] add_959411;
  wire [7:0] sel_959412;
  wire [7:0] add_959415;
  wire [7:0] sel_959416;
  wire [7:0] add_959419;
  wire [7:0] sel_959420;
  wire [7:0] add_959423;
  wire [7:0] sel_959424;
  wire [7:0] add_959427;
  wire [7:0] sel_959428;
  wire [7:0] add_959431;
  wire [7:0] sel_959432;
  wire [7:0] add_959435;
  wire [7:0] sel_959436;
  wire [7:0] add_959439;
  wire [7:0] sel_959440;
  wire [7:0] add_959443;
  wire [7:0] sel_959444;
  wire [7:0] add_959447;
  wire [7:0] sel_959448;
  wire [7:0] add_959451;
  wire [7:0] sel_959452;
  wire [7:0] add_959455;
  wire [7:0] sel_959456;
  wire [7:0] add_959459;
  wire [7:0] sel_959460;
  wire [7:0] add_959463;
  wire [7:0] sel_959464;
  wire [7:0] add_959467;
  wire [7:0] sel_959468;
  wire [7:0] add_959471;
  wire [7:0] sel_959472;
  wire [7:0] add_959475;
  wire [7:0] sel_959476;
  wire [7:0] add_959479;
  wire [7:0] sel_959480;
  wire [7:0] add_959483;
  wire [7:0] sel_959484;
  wire [7:0] add_959487;
  wire [7:0] sel_959488;
  wire [7:0] add_959491;
  wire [7:0] sel_959492;
  wire [7:0] add_959495;
  wire [7:0] sel_959496;
  wire [7:0] add_959499;
  wire [7:0] sel_959500;
  wire [7:0] add_959503;
  wire [7:0] sel_959504;
  wire [7:0] add_959507;
  wire [7:0] sel_959508;
  wire [7:0] add_959511;
  wire [7:0] sel_959512;
  wire [7:0] add_959515;
  wire [7:0] sel_959516;
  wire [7:0] add_959519;
  wire [7:0] sel_959520;
  wire [7:0] add_959523;
  wire [7:0] sel_959524;
  wire [7:0] add_959527;
  wire [7:0] sel_959528;
  wire [7:0] add_959531;
  wire [7:0] sel_959532;
  wire [7:0] add_959535;
  wire [7:0] sel_959536;
  wire [7:0] add_959539;
  wire [7:0] sel_959540;
  wire [7:0] add_959544;
  wire [15:0] array_index_959545;
  wire [7:0] sel_959546;
  wire [7:0] add_959549;
  wire [7:0] sel_959550;
  wire [7:0] add_959553;
  wire [7:0] sel_959554;
  wire [7:0] add_959557;
  wire [7:0] sel_959558;
  wire [7:0] add_959561;
  wire [7:0] sel_959562;
  wire [7:0] add_959565;
  wire [7:0] sel_959566;
  wire [7:0] add_959569;
  wire [7:0] sel_959570;
  wire [7:0] add_959573;
  wire [7:0] sel_959574;
  wire [7:0] add_959577;
  wire [7:0] sel_959578;
  wire [7:0] add_959581;
  wire [7:0] sel_959582;
  wire [7:0] add_959585;
  wire [7:0] sel_959586;
  wire [7:0] add_959589;
  wire [7:0] sel_959590;
  wire [7:0] add_959593;
  wire [7:0] sel_959594;
  wire [7:0] add_959597;
  wire [7:0] sel_959598;
  wire [7:0] add_959601;
  wire [7:0] sel_959602;
  wire [7:0] add_959605;
  wire [7:0] sel_959606;
  wire [7:0] add_959609;
  wire [7:0] sel_959610;
  wire [7:0] add_959613;
  wire [7:0] sel_959614;
  wire [7:0] add_959617;
  wire [7:0] sel_959618;
  wire [7:0] add_959621;
  wire [7:0] sel_959622;
  wire [7:0] add_959625;
  wire [7:0] sel_959626;
  wire [7:0] add_959629;
  wire [7:0] sel_959630;
  wire [7:0] add_959633;
  wire [7:0] sel_959634;
  wire [7:0] add_959637;
  wire [7:0] sel_959638;
  wire [7:0] add_959641;
  wire [7:0] sel_959642;
  wire [7:0] add_959645;
  wire [7:0] sel_959646;
  wire [7:0] add_959649;
  wire [7:0] sel_959650;
  wire [7:0] add_959653;
  wire [7:0] sel_959654;
  wire [7:0] add_959657;
  wire [7:0] sel_959658;
  wire [7:0] add_959661;
  wire [7:0] sel_959662;
  wire [7:0] add_959665;
  wire [7:0] sel_959666;
  wire [7:0] add_959669;
  wire [7:0] sel_959670;
  wire [7:0] add_959673;
  wire [7:0] sel_959674;
  wire [7:0] add_959677;
  wire [7:0] sel_959678;
  wire [7:0] add_959681;
  wire [7:0] sel_959682;
  wire [7:0] add_959685;
  wire [7:0] sel_959686;
  wire [7:0] add_959689;
  wire [7:0] sel_959690;
  wire [7:0] add_959693;
  wire [7:0] sel_959694;
  wire [7:0] add_959697;
  wire [7:0] sel_959698;
  wire [7:0] add_959701;
  wire [7:0] sel_959702;
  wire [7:0] add_959705;
  wire [7:0] sel_959706;
  wire [7:0] add_959709;
  wire [7:0] sel_959710;
  wire [7:0] add_959713;
  wire [7:0] sel_959714;
  wire [7:0] add_959717;
  wire [7:0] sel_959718;
  wire [7:0] add_959721;
  wire [7:0] sel_959722;
  wire [7:0] add_959725;
  wire [7:0] sel_959726;
  wire [7:0] add_959729;
  wire [7:0] sel_959730;
  wire [7:0] add_959733;
  wire [7:0] sel_959734;
  wire [7:0] add_959737;
  wire [7:0] sel_959738;
  wire [7:0] add_959741;
  wire [7:0] sel_959742;
  wire [7:0] add_959745;
  wire [7:0] sel_959746;
  wire [7:0] add_959749;
  wire [7:0] sel_959750;
  wire [7:0] add_959753;
  wire [7:0] sel_959754;
  wire [7:0] add_959757;
  wire [7:0] sel_959758;
  wire [7:0] add_959761;
  wire [7:0] sel_959762;
  wire [7:0] add_959765;
  wire [7:0] sel_959766;
  wire [7:0] add_959769;
  wire [7:0] sel_959770;
  wire [7:0] add_959773;
  wire [7:0] sel_959774;
  wire [7:0] add_959777;
  wire [7:0] sel_959778;
  wire [7:0] add_959781;
  wire [7:0] sel_959782;
  wire [7:0] add_959785;
  wire [7:0] sel_959786;
  wire [7:0] add_959789;
  wire [7:0] sel_959790;
  wire [7:0] add_959793;
  wire [7:0] sel_959794;
  wire [7:0] add_959797;
  wire [7:0] sel_959798;
  wire [7:0] add_959801;
  wire [7:0] sel_959802;
  wire [7:0] add_959805;
  wire [7:0] sel_959806;
  wire [7:0] add_959809;
  wire [7:0] sel_959810;
  wire [7:0] add_959813;
  wire [7:0] sel_959814;
  wire [7:0] add_959817;
  wire [7:0] sel_959818;
  wire [7:0] add_959821;
  wire [7:0] sel_959822;
  wire [7:0] add_959825;
  wire [7:0] sel_959826;
  wire [7:0] add_959829;
  wire [7:0] sel_959830;
  wire [7:0] add_959833;
  wire [7:0] sel_959834;
  wire [7:0] add_959837;
  wire [7:0] sel_959838;
  wire [7:0] add_959841;
  wire [7:0] sel_959842;
  wire [7:0] add_959845;
  wire [7:0] sel_959846;
  wire [7:0] add_959849;
  wire [7:0] sel_959850;
  wire [7:0] add_959853;
  wire [7:0] sel_959854;
  wire [7:0] add_959857;
  wire [7:0] sel_959858;
  wire [7:0] add_959861;
  wire [7:0] sel_959862;
  wire [7:0] add_959865;
  wire [7:0] sel_959866;
  wire [7:0] add_959869;
  wire [7:0] sel_959870;
  wire [7:0] add_959873;
  wire [7:0] sel_959874;
  wire [7:0] add_959877;
  wire [7:0] sel_959878;
  wire [7:0] add_959881;
  wire [7:0] sel_959882;
  wire [7:0] add_959885;
  wire [7:0] sel_959886;
  wire [7:0] add_959889;
  wire [7:0] sel_959890;
  wire [7:0] add_959893;
  wire [7:0] sel_959894;
  wire [7:0] add_959897;
  wire [7:0] sel_959898;
  wire [7:0] add_959901;
  wire [7:0] sel_959902;
  wire [7:0] add_959905;
  wire [7:0] sel_959906;
  wire [7:0] add_959909;
  wire [7:0] sel_959910;
  wire [7:0] add_959913;
  wire [7:0] sel_959914;
  wire [7:0] add_959917;
  wire [7:0] sel_959918;
  wire [7:0] add_959921;
  wire [7:0] sel_959922;
  wire [7:0] add_959925;
  wire [7:0] sel_959926;
  wire [7:0] add_959929;
  wire [7:0] sel_959930;
  wire [7:0] add_959933;
  wire [7:0] sel_959934;
  wire [7:0] add_959937;
  wire [7:0] sel_959938;
  wire [7:0] add_959941;
  wire [7:0] sel_959942;
  wire [7:0] add_959946;
  wire [15:0] array_index_959947;
  wire [7:0] sel_959948;
  wire [7:0] add_959951;
  wire [7:0] sel_959952;
  wire [7:0] add_959955;
  wire [7:0] sel_959956;
  wire [7:0] add_959959;
  wire [7:0] sel_959960;
  wire [7:0] add_959963;
  wire [7:0] sel_959964;
  wire [7:0] add_959967;
  wire [7:0] sel_959968;
  wire [7:0] add_959971;
  wire [7:0] sel_959972;
  wire [7:0] add_959975;
  wire [7:0] sel_959976;
  wire [7:0] add_959979;
  wire [7:0] sel_959980;
  wire [7:0] add_959983;
  wire [7:0] sel_959984;
  wire [7:0] add_959987;
  wire [7:0] sel_959988;
  wire [7:0] add_959991;
  wire [7:0] sel_959992;
  wire [7:0] add_959995;
  wire [7:0] sel_959996;
  wire [7:0] add_959999;
  wire [7:0] sel_960000;
  wire [7:0] add_960003;
  wire [7:0] sel_960004;
  wire [7:0] add_960007;
  wire [7:0] sel_960008;
  wire [7:0] add_960011;
  wire [7:0] sel_960012;
  wire [7:0] add_960015;
  wire [7:0] sel_960016;
  wire [7:0] add_960019;
  wire [7:0] sel_960020;
  wire [7:0] add_960023;
  wire [7:0] sel_960024;
  wire [7:0] add_960027;
  wire [7:0] sel_960028;
  wire [7:0] add_960031;
  wire [7:0] sel_960032;
  wire [7:0] add_960035;
  wire [7:0] sel_960036;
  wire [7:0] add_960039;
  wire [7:0] sel_960040;
  wire [7:0] add_960043;
  wire [7:0] sel_960044;
  wire [7:0] add_960047;
  wire [7:0] sel_960048;
  wire [7:0] add_960051;
  wire [7:0] sel_960052;
  wire [7:0] add_960055;
  wire [7:0] sel_960056;
  wire [7:0] add_960059;
  wire [7:0] sel_960060;
  wire [7:0] add_960063;
  wire [7:0] sel_960064;
  wire [7:0] add_960067;
  wire [7:0] sel_960068;
  wire [7:0] add_960071;
  wire [7:0] sel_960072;
  wire [7:0] add_960075;
  wire [7:0] sel_960076;
  wire [7:0] add_960079;
  wire [7:0] sel_960080;
  wire [7:0] add_960083;
  wire [7:0] sel_960084;
  wire [7:0] add_960087;
  wire [7:0] sel_960088;
  wire [7:0] add_960091;
  wire [7:0] sel_960092;
  wire [7:0] add_960095;
  wire [7:0] sel_960096;
  wire [7:0] add_960099;
  wire [7:0] sel_960100;
  wire [7:0] add_960103;
  wire [7:0] sel_960104;
  wire [7:0] add_960107;
  wire [7:0] sel_960108;
  wire [7:0] add_960111;
  wire [7:0] sel_960112;
  wire [7:0] add_960115;
  wire [7:0] sel_960116;
  wire [7:0] add_960119;
  wire [7:0] sel_960120;
  wire [7:0] add_960123;
  wire [7:0] sel_960124;
  wire [7:0] add_960127;
  wire [7:0] sel_960128;
  wire [7:0] add_960131;
  wire [7:0] sel_960132;
  wire [7:0] add_960135;
  wire [7:0] sel_960136;
  wire [7:0] add_960139;
  wire [7:0] sel_960140;
  wire [7:0] add_960143;
  wire [7:0] sel_960144;
  wire [7:0] add_960147;
  wire [7:0] sel_960148;
  wire [7:0] add_960151;
  wire [7:0] sel_960152;
  wire [7:0] add_960155;
  wire [7:0] sel_960156;
  wire [7:0] add_960159;
  wire [7:0] sel_960160;
  wire [7:0] add_960163;
  wire [7:0] sel_960164;
  wire [7:0] add_960167;
  wire [7:0] sel_960168;
  wire [7:0] add_960171;
  wire [7:0] sel_960172;
  wire [7:0] add_960175;
  wire [7:0] sel_960176;
  wire [7:0] add_960179;
  wire [7:0] sel_960180;
  wire [7:0] add_960183;
  wire [7:0] sel_960184;
  wire [7:0] add_960187;
  wire [7:0] sel_960188;
  wire [7:0] add_960191;
  wire [7:0] sel_960192;
  wire [7:0] add_960195;
  wire [7:0] sel_960196;
  wire [7:0] add_960199;
  wire [7:0] sel_960200;
  wire [7:0] add_960203;
  wire [7:0] sel_960204;
  wire [7:0] add_960207;
  wire [7:0] sel_960208;
  wire [7:0] add_960211;
  wire [7:0] sel_960212;
  wire [7:0] add_960215;
  wire [7:0] sel_960216;
  wire [7:0] add_960219;
  wire [7:0] sel_960220;
  wire [7:0] add_960223;
  wire [7:0] sel_960224;
  wire [7:0] add_960227;
  wire [7:0] sel_960228;
  wire [7:0] add_960231;
  wire [7:0] sel_960232;
  wire [7:0] add_960235;
  wire [7:0] sel_960236;
  wire [7:0] add_960239;
  wire [7:0] sel_960240;
  wire [7:0] add_960243;
  wire [7:0] sel_960244;
  wire [7:0] add_960247;
  wire [7:0] sel_960248;
  wire [7:0] add_960251;
  wire [7:0] sel_960252;
  wire [7:0] add_960255;
  wire [7:0] sel_960256;
  wire [7:0] add_960259;
  wire [7:0] sel_960260;
  wire [7:0] add_960263;
  wire [7:0] sel_960264;
  wire [7:0] add_960267;
  wire [7:0] sel_960268;
  wire [7:0] add_960271;
  wire [7:0] sel_960272;
  wire [7:0] add_960275;
  wire [7:0] sel_960276;
  wire [7:0] add_960279;
  wire [7:0] sel_960280;
  wire [7:0] add_960283;
  wire [7:0] sel_960284;
  wire [7:0] add_960287;
  wire [7:0] sel_960288;
  wire [7:0] add_960291;
  wire [7:0] sel_960292;
  wire [7:0] add_960295;
  wire [7:0] sel_960296;
  wire [7:0] add_960299;
  wire [7:0] sel_960300;
  wire [7:0] add_960303;
  wire [7:0] sel_960304;
  wire [7:0] add_960307;
  wire [7:0] sel_960308;
  wire [7:0] add_960311;
  wire [7:0] sel_960312;
  wire [7:0] add_960315;
  wire [7:0] sel_960316;
  wire [7:0] add_960319;
  wire [7:0] sel_960320;
  wire [7:0] add_960323;
  wire [7:0] sel_960324;
  wire [7:0] add_960327;
  wire [7:0] sel_960328;
  wire [7:0] add_960331;
  wire [7:0] sel_960332;
  wire [7:0] add_960335;
  wire [7:0] sel_960336;
  wire [7:0] add_960339;
  wire [7:0] sel_960340;
  wire [7:0] add_960343;
  wire [7:0] sel_960344;
  wire [7:0] add_960348;
  wire [15:0] array_index_960349;
  wire [7:0] sel_960350;
  wire [7:0] add_960353;
  wire [7:0] sel_960354;
  wire [7:0] add_960357;
  wire [7:0] sel_960358;
  wire [7:0] add_960361;
  wire [7:0] sel_960362;
  wire [7:0] add_960365;
  wire [7:0] sel_960366;
  wire [7:0] add_960369;
  wire [7:0] sel_960370;
  wire [7:0] add_960373;
  wire [7:0] sel_960374;
  wire [7:0] add_960377;
  wire [7:0] sel_960378;
  wire [7:0] add_960381;
  wire [7:0] sel_960382;
  wire [7:0] add_960385;
  wire [7:0] sel_960386;
  wire [7:0] add_960389;
  wire [7:0] sel_960390;
  wire [7:0] add_960393;
  wire [7:0] sel_960394;
  wire [7:0] add_960397;
  wire [7:0] sel_960398;
  wire [7:0] add_960401;
  wire [7:0] sel_960402;
  wire [7:0] add_960405;
  wire [7:0] sel_960406;
  wire [7:0] add_960409;
  wire [7:0] sel_960410;
  wire [7:0] add_960413;
  wire [7:0] sel_960414;
  wire [7:0] add_960417;
  wire [7:0] sel_960418;
  wire [7:0] add_960421;
  wire [7:0] sel_960422;
  wire [7:0] add_960425;
  wire [7:0] sel_960426;
  wire [7:0] add_960429;
  wire [7:0] sel_960430;
  wire [7:0] add_960433;
  wire [7:0] sel_960434;
  wire [7:0] add_960437;
  wire [7:0] sel_960438;
  wire [7:0] add_960441;
  wire [7:0] sel_960442;
  wire [7:0] add_960445;
  wire [7:0] sel_960446;
  wire [7:0] add_960449;
  wire [7:0] sel_960450;
  wire [7:0] add_960453;
  wire [7:0] sel_960454;
  wire [7:0] add_960457;
  wire [7:0] sel_960458;
  wire [7:0] add_960461;
  wire [7:0] sel_960462;
  wire [7:0] add_960465;
  wire [7:0] sel_960466;
  wire [7:0] add_960469;
  wire [7:0] sel_960470;
  wire [7:0] add_960473;
  wire [7:0] sel_960474;
  wire [7:0] add_960477;
  wire [7:0] sel_960478;
  wire [7:0] add_960481;
  wire [7:0] sel_960482;
  wire [7:0] add_960485;
  wire [7:0] sel_960486;
  wire [7:0] add_960489;
  wire [7:0] sel_960490;
  wire [7:0] add_960493;
  wire [7:0] sel_960494;
  wire [7:0] add_960497;
  wire [7:0] sel_960498;
  wire [7:0] add_960501;
  wire [7:0] sel_960502;
  wire [7:0] add_960505;
  wire [7:0] sel_960506;
  wire [7:0] add_960509;
  wire [7:0] sel_960510;
  wire [7:0] add_960513;
  wire [7:0] sel_960514;
  wire [7:0] add_960517;
  wire [7:0] sel_960518;
  wire [7:0] add_960521;
  wire [7:0] sel_960522;
  wire [7:0] add_960525;
  wire [7:0] sel_960526;
  wire [7:0] add_960529;
  wire [7:0] sel_960530;
  wire [7:0] add_960533;
  wire [7:0] sel_960534;
  wire [7:0] add_960537;
  wire [7:0] sel_960538;
  wire [7:0] add_960541;
  wire [7:0] sel_960542;
  wire [7:0] add_960545;
  wire [7:0] sel_960546;
  wire [7:0] add_960549;
  wire [7:0] sel_960550;
  wire [7:0] add_960553;
  wire [7:0] sel_960554;
  wire [7:0] add_960557;
  wire [7:0] sel_960558;
  wire [7:0] add_960561;
  wire [7:0] sel_960562;
  wire [7:0] add_960565;
  wire [7:0] sel_960566;
  wire [7:0] add_960569;
  wire [7:0] sel_960570;
  wire [7:0] add_960573;
  wire [7:0] sel_960574;
  wire [7:0] add_960577;
  wire [7:0] sel_960578;
  wire [7:0] add_960581;
  wire [7:0] sel_960582;
  wire [7:0] add_960585;
  wire [7:0] sel_960586;
  wire [7:0] add_960589;
  wire [7:0] sel_960590;
  wire [7:0] add_960593;
  wire [7:0] sel_960594;
  wire [7:0] add_960597;
  wire [7:0] sel_960598;
  wire [7:0] add_960601;
  wire [7:0] sel_960602;
  wire [7:0] add_960605;
  wire [7:0] sel_960606;
  wire [7:0] add_960609;
  wire [7:0] sel_960610;
  wire [7:0] add_960613;
  wire [7:0] sel_960614;
  wire [7:0] add_960617;
  wire [7:0] sel_960618;
  wire [7:0] add_960621;
  wire [7:0] sel_960622;
  wire [7:0] add_960625;
  wire [7:0] sel_960626;
  wire [7:0] add_960629;
  wire [7:0] sel_960630;
  wire [7:0] add_960633;
  wire [7:0] sel_960634;
  wire [7:0] add_960637;
  wire [7:0] sel_960638;
  wire [7:0] add_960641;
  wire [7:0] sel_960642;
  wire [7:0] add_960645;
  wire [7:0] sel_960646;
  wire [7:0] add_960649;
  wire [7:0] sel_960650;
  wire [7:0] add_960653;
  wire [7:0] sel_960654;
  wire [7:0] add_960657;
  wire [7:0] sel_960658;
  wire [7:0] add_960661;
  wire [7:0] sel_960662;
  wire [7:0] add_960665;
  wire [7:0] sel_960666;
  wire [7:0] add_960669;
  wire [7:0] sel_960670;
  wire [7:0] add_960673;
  wire [7:0] sel_960674;
  wire [7:0] add_960677;
  wire [7:0] sel_960678;
  wire [7:0] add_960681;
  wire [7:0] sel_960682;
  wire [7:0] add_960685;
  wire [7:0] sel_960686;
  wire [7:0] add_960689;
  wire [7:0] sel_960690;
  wire [7:0] add_960693;
  wire [7:0] sel_960694;
  wire [7:0] add_960697;
  wire [7:0] sel_960698;
  wire [7:0] add_960701;
  wire [7:0] sel_960702;
  wire [7:0] add_960705;
  wire [7:0] sel_960706;
  wire [7:0] add_960709;
  wire [7:0] sel_960710;
  wire [7:0] add_960713;
  wire [7:0] sel_960714;
  wire [7:0] add_960717;
  wire [7:0] sel_960718;
  wire [7:0] add_960721;
  wire [7:0] sel_960722;
  wire [7:0] add_960725;
  wire [7:0] sel_960726;
  wire [7:0] add_960729;
  wire [7:0] sel_960730;
  wire [7:0] add_960733;
  wire [7:0] sel_960734;
  wire [7:0] add_960737;
  wire [7:0] sel_960738;
  wire [7:0] add_960741;
  wire [7:0] sel_960742;
  wire [7:0] add_960745;
  wire [7:0] sel_960746;
  wire [7:0] add_960750;
  wire [15:0] array_index_960751;
  wire [7:0] sel_960752;
  wire [7:0] add_960755;
  wire [7:0] sel_960756;
  wire [7:0] add_960759;
  wire [7:0] sel_960760;
  wire [7:0] add_960763;
  wire [7:0] sel_960764;
  wire [7:0] add_960767;
  wire [7:0] sel_960768;
  wire [7:0] add_960771;
  wire [7:0] sel_960772;
  wire [7:0] add_960775;
  wire [7:0] sel_960776;
  wire [7:0] add_960779;
  wire [7:0] sel_960780;
  wire [7:0] add_960783;
  wire [7:0] sel_960784;
  wire [7:0] add_960787;
  wire [7:0] sel_960788;
  wire [7:0] add_960791;
  wire [7:0] sel_960792;
  wire [7:0] add_960795;
  wire [7:0] sel_960796;
  wire [7:0] add_960799;
  wire [7:0] sel_960800;
  wire [7:0] add_960803;
  wire [7:0] sel_960804;
  wire [7:0] add_960807;
  wire [7:0] sel_960808;
  wire [7:0] add_960811;
  wire [7:0] sel_960812;
  wire [7:0] add_960815;
  wire [7:0] sel_960816;
  wire [7:0] add_960819;
  wire [7:0] sel_960820;
  wire [7:0] add_960823;
  wire [7:0] sel_960824;
  wire [7:0] add_960827;
  wire [7:0] sel_960828;
  wire [7:0] add_960831;
  wire [7:0] sel_960832;
  wire [7:0] add_960835;
  wire [7:0] sel_960836;
  wire [7:0] add_960839;
  wire [7:0] sel_960840;
  wire [7:0] add_960843;
  wire [7:0] sel_960844;
  wire [7:0] add_960847;
  wire [7:0] sel_960848;
  wire [7:0] add_960851;
  wire [7:0] sel_960852;
  wire [7:0] add_960855;
  wire [7:0] sel_960856;
  wire [7:0] add_960859;
  wire [7:0] sel_960860;
  wire [7:0] add_960863;
  wire [7:0] sel_960864;
  wire [7:0] add_960867;
  wire [7:0] sel_960868;
  wire [7:0] add_960871;
  wire [7:0] sel_960872;
  wire [7:0] add_960875;
  wire [7:0] sel_960876;
  wire [7:0] add_960879;
  wire [7:0] sel_960880;
  wire [7:0] add_960883;
  wire [7:0] sel_960884;
  wire [7:0] add_960887;
  wire [7:0] sel_960888;
  wire [7:0] add_960891;
  wire [7:0] sel_960892;
  wire [7:0] add_960895;
  wire [7:0] sel_960896;
  wire [7:0] add_960899;
  wire [7:0] sel_960900;
  wire [7:0] add_960903;
  wire [7:0] sel_960904;
  wire [7:0] add_960907;
  wire [7:0] sel_960908;
  wire [7:0] add_960911;
  wire [7:0] sel_960912;
  wire [7:0] add_960915;
  wire [7:0] sel_960916;
  wire [7:0] add_960919;
  wire [7:0] sel_960920;
  wire [7:0] add_960923;
  wire [7:0] sel_960924;
  wire [7:0] add_960927;
  wire [7:0] sel_960928;
  wire [7:0] add_960931;
  wire [7:0] sel_960932;
  wire [7:0] add_960935;
  wire [7:0] sel_960936;
  wire [7:0] add_960939;
  wire [7:0] sel_960940;
  wire [7:0] add_960943;
  wire [7:0] sel_960944;
  wire [7:0] add_960947;
  wire [7:0] sel_960948;
  wire [7:0] add_960951;
  wire [7:0] sel_960952;
  wire [7:0] add_960955;
  wire [7:0] sel_960956;
  wire [7:0] add_960959;
  wire [7:0] sel_960960;
  wire [7:0] add_960963;
  wire [7:0] sel_960964;
  wire [7:0] add_960967;
  wire [7:0] sel_960968;
  wire [7:0] add_960971;
  wire [7:0] sel_960972;
  wire [7:0] add_960975;
  wire [7:0] sel_960976;
  wire [7:0] add_960979;
  wire [7:0] sel_960980;
  wire [7:0] add_960983;
  wire [7:0] sel_960984;
  wire [7:0] add_960987;
  wire [7:0] sel_960988;
  wire [7:0] add_960991;
  wire [7:0] sel_960992;
  wire [7:0] add_960995;
  wire [7:0] sel_960996;
  wire [7:0] add_960999;
  wire [7:0] sel_961000;
  wire [7:0] add_961003;
  wire [7:0] sel_961004;
  wire [7:0] add_961007;
  wire [7:0] sel_961008;
  wire [7:0] add_961011;
  wire [7:0] sel_961012;
  wire [7:0] add_961015;
  wire [7:0] sel_961016;
  wire [7:0] add_961019;
  wire [7:0] sel_961020;
  wire [7:0] add_961023;
  wire [7:0] sel_961024;
  wire [7:0] add_961027;
  wire [7:0] sel_961028;
  wire [7:0] add_961031;
  wire [7:0] sel_961032;
  wire [7:0] add_961035;
  wire [7:0] sel_961036;
  wire [7:0] add_961039;
  wire [7:0] sel_961040;
  wire [7:0] add_961043;
  wire [7:0] sel_961044;
  wire [7:0] add_961047;
  wire [7:0] sel_961048;
  wire [7:0] add_961051;
  wire [7:0] sel_961052;
  wire [7:0] add_961055;
  wire [7:0] sel_961056;
  wire [7:0] add_961059;
  wire [7:0] sel_961060;
  wire [7:0] add_961063;
  wire [7:0] sel_961064;
  wire [7:0] add_961067;
  wire [7:0] sel_961068;
  wire [7:0] add_961071;
  wire [7:0] sel_961072;
  wire [7:0] add_961075;
  wire [7:0] sel_961076;
  wire [7:0] add_961079;
  wire [7:0] sel_961080;
  wire [7:0] add_961083;
  wire [7:0] sel_961084;
  wire [7:0] add_961087;
  wire [7:0] sel_961088;
  wire [7:0] add_961091;
  wire [7:0] sel_961092;
  wire [7:0] add_961095;
  wire [7:0] sel_961096;
  wire [7:0] add_961099;
  wire [7:0] sel_961100;
  wire [7:0] add_961103;
  wire [7:0] sel_961104;
  wire [7:0] add_961107;
  wire [7:0] sel_961108;
  wire [7:0] add_961111;
  wire [7:0] sel_961112;
  wire [7:0] add_961115;
  wire [7:0] sel_961116;
  wire [7:0] add_961119;
  wire [7:0] sel_961120;
  wire [7:0] add_961123;
  wire [7:0] sel_961124;
  wire [7:0] add_961127;
  wire [7:0] sel_961128;
  wire [7:0] add_961131;
  wire [7:0] sel_961132;
  wire [7:0] add_961135;
  wire [7:0] sel_961136;
  wire [7:0] add_961139;
  wire [7:0] sel_961140;
  wire [7:0] add_961143;
  wire [7:0] sel_961144;
  wire [7:0] add_961147;
  wire [7:0] sel_961148;
  wire [7:0] add_961152;
  wire [15:0] array_index_961153;
  wire [7:0] sel_961154;
  wire [7:0] add_961157;
  wire [7:0] sel_961158;
  wire [7:0] add_961161;
  wire [7:0] sel_961162;
  wire [7:0] add_961165;
  wire [7:0] sel_961166;
  wire [7:0] add_961169;
  wire [7:0] sel_961170;
  wire [7:0] add_961173;
  wire [7:0] sel_961174;
  wire [7:0] add_961177;
  wire [7:0] sel_961178;
  wire [7:0] add_961181;
  wire [7:0] sel_961182;
  wire [7:0] add_961185;
  wire [7:0] sel_961186;
  wire [7:0] add_961189;
  wire [7:0] sel_961190;
  wire [7:0] add_961193;
  wire [7:0] sel_961194;
  wire [7:0] add_961197;
  wire [7:0] sel_961198;
  wire [7:0] add_961201;
  wire [7:0] sel_961202;
  wire [7:0] add_961205;
  wire [7:0] sel_961206;
  wire [7:0] add_961209;
  wire [7:0] sel_961210;
  wire [7:0] add_961213;
  wire [7:0] sel_961214;
  wire [7:0] add_961217;
  wire [7:0] sel_961218;
  wire [7:0] add_961221;
  wire [7:0] sel_961222;
  wire [7:0] add_961225;
  wire [7:0] sel_961226;
  wire [7:0] add_961229;
  wire [7:0] sel_961230;
  wire [7:0] add_961233;
  wire [7:0] sel_961234;
  wire [7:0] add_961237;
  wire [7:0] sel_961238;
  wire [7:0] add_961241;
  wire [7:0] sel_961242;
  wire [7:0] add_961245;
  wire [7:0] sel_961246;
  wire [7:0] add_961249;
  wire [7:0] sel_961250;
  wire [7:0] add_961253;
  wire [7:0] sel_961254;
  wire [7:0] add_961257;
  wire [7:0] sel_961258;
  wire [7:0] add_961261;
  wire [7:0] sel_961262;
  wire [7:0] add_961265;
  wire [7:0] sel_961266;
  wire [7:0] add_961269;
  wire [7:0] sel_961270;
  wire [7:0] add_961273;
  wire [7:0] sel_961274;
  wire [7:0] add_961277;
  wire [7:0] sel_961278;
  wire [7:0] add_961281;
  wire [7:0] sel_961282;
  wire [7:0] add_961285;
  wire [7:0] sel_961286;
  wire [7:0] add_961289;
  wire [7:0] sel_961290;
  wire [7:0] add_961293;
  wire [7:0] sel_961294;
  wire [7:0] add_961297;
  wire [7:0] sel_961298;
  wire [7:0] add_961301;
  wire [7:0] sel_961302;
  wire [7:0] add_961305;
  wire [7:0] sel_961306;
  wire [7:0] add_961309;
  wire [7:0] sel_961310;
  wire [7:0] add_961313;
  wire [7:0] sel_961314;
  wire [7:0] add_961317;
  wire [7:0] sel_961318;
  wire [7:0] add_961321;
  wire [7:0] sel_961322;
  wire [7:0] add_961325;
  wire [7:0] sel_961326;
  wire [7:0] add_961329;
  wire [7:0] sel_961330;
  wire [7:0] add_961333;
  wire [7:0] sel_961334;
  wire [7:0] add_961337;
  wire [7:0] sel_961338;
  wire [7:0] add_961341;
  wire [7:0] sel_961342;
  wire [7:0] add_961345;
  wire [7:0] sel_961346;
  wire [7:0] add_961349;
  wire [7:0] sel_961350;
  wire [7:0] add_961353;
  wire [7:0] sel_961354;
  wire [7:0] add_961357;
  wire [7:0] sel_961358;
  wire [7:0] add_961361;
  wire [7:0] sel_961362;
  wire [7:0] add_961365;
  wire [7:0] sel_961366;
  wire [7:0] add_961369;
  wire [7:0] sel_961370;
  wire [7:0] add_961373;
  wire [7:0] sel_961374;
  wire [7:0] add_961377;
  wire [7:0] sel_961378;
  wire [7:0] add_961381;
  wire [7:0] sel_961382;
  wire [7:0] add_961385;
  wire [7:0] sel_961386;
  wire [7:0] add_961389;
  wire [7:0] sel_961390;
  wire [7:0] add_961393;
  wire [7:0] sel_961394;
  wire [7:0] add_961397;
  wire [7:0] sel_961398;
  wire [7:0] add_961401;
  wire [7:0] sel_961402;
  wire [7:0] add_961405;
  wire [7:0] sel_961406;
  wire [7:0] add_961409;
  wire [7:0] sel_961410;
  wire [7:0] add_961413;
  wire [7:0] sel_961414;
  wire [7:0] add_961417;
  wire [7:0] sel_961418;
  wire [7:0] add_961421;
  wire [7:0] sel_961422;
  wire [7:0] add_961425;
  wire [7:0] sel_961426;
  wire [7:0] add_961429;
  wire [7:0] sel_961430;
  wire [7:0] add_961433;
  wire [7:0] sel_961434;
  wire [7:0] add_961437;
  wire [7:0] sel_961438;
  wire [7:0] add_961441;
  wire [7:0] sel_961442;
  wire [7:0] add_961445;
  wire [7:0] sel_961446;
  wire [7:0] add_961449;
  wire [7:0] sel_961450;
  wire [7:0] add_961453;
  wire [7:0] sel_961454;
  wire [7:0] add_961457;
  wire [7:0] sel_961458;
  wire [7:0] add_961461;
  wire [7:0] sel_961462;
  wire [7:0] add_961465;
  wire [7:0] sel_961466;
  wire [7:0] add_961469;
  wire [7:0] sel_961470;
  wire [7:0] add_961473;
  wire [7:0] sel_961474;
  wire [7:0] add_961477;
  wire [7:0] sel_961478;
  wire [7:0] add_961481;
  wire [7:0] sel_961482;
  wire [7:0] add_961485;
  wire [7:0] sel_961486;
  wire [7:0] add_961489;
  wire [7:0] sel_961490;
  wire [7:0] add_961493;
  wire [7:0] sel_961494;
  wire [7:0] add_961497;
  wire [7:0] sel_961498;
  wire [7:0] add_961501;
  wire [7:0] sel_961502;
  wire [7:0] add_961505;
  wire [7:0] sel_961506;
  wire [7:0] add_961509;
  wire [7:0] sel_961510;
  wire [7:0] add_961513;
  wire [7:0] sel_961514;
  wire [7:0] add_961517;
  wire [7:0] sel_961518;
  wire [7:0] add_961521;
  wire [7:0] sel_961522;
  wire [7:0] add_961525;
  wire [7:0] sel_961526;
  wire [7:0] add_961529;
  wire [7:0] sel_961530;
  wire [7:0] add_961533;
  wire [7:0] sel_961534;
  wire [7:0] add_961537;
  wire [7:0] sel_961538;
  wire [7:0] add_961541;
  wire [7:0] sel_961542;
  wire [7:0] add_961545;
  wire [7:0] sel_961546;
  wire [7:0] add_961549;
  wire [7:0] sel_961550;
  wire [7:0] add_961554;
  wire [15:0] array_index_961555;
  wire [7:0] sel_961556;
  wire [7:0] add_961559;
  wire [7:0] sel_961560;
  wire [7:0] add_961563;
  wire [7:0] sel_961564;
  wire [7:0] add_961567;
  wire [7:0] sel_961568;
  wire [7:0] add_961571;
  wire [7:0] sel_961572;
  wire [7:0] add_961575;
  wire [7:0] sel_961576;
  wire [7:0] add_961579;
  wire [7:0] sel_961580;
  wire [7:0] add_961583;
  wire [7:0] sel_961584;
  wire [7:0] add_961587;
  wire [7:0] sel_961588;
  wire [7:0] add_961591;
  wire [7:0] sel_961592;
  wire [7:0] add_961595;
  wire [7:0] sel_961596;
  wire [7:0] add_961599;
  wire [7:0] sel_961600;
  wire [7:0] add_961603;
  wire [7:0] sel_961604;
  wire [7:0] add_961607;
  wire [7:0] sel_961608;
  wire [7:0] add_961611;
  wire [7:0] sel_961612;
  wire [7:0] add_961615;
  wire [7:0] sel_961616;
  wire [7:0] add_961619;
  wire [7:0] sel_961620;
  wire [7:0] add_961623;
  wire [7:0] sel_961624;
  wire [7:0] add_961627;
  wire [7:0] sel_961628;
  wire [7:0] add_961631;
  wire [7:0] sel_961632;
  wire [7:0] add_961635;
  wire [7:0] sel_961636;
  wire [7:0] add_961639;
  wire [7:0] sel_961640;
  wire [7:0] add_961643;
  wire [7:0] sel_961644;
  wire [7:0] add_961647;
  wire [7:0] sel_961648;
  wire [7:0] add_961651;
  wire [7:0] sel_961652;
  wire [7:0] add_961655;
  wire [7:0] sel_961656;
  wire [7:0] add_961659;
  wire [7:0] sel_961660;
  wire [7:0] add_961663;
  wire [7:0] sel_961664;
  wire [7:0] add_961667;
  wire [7:0] sel_961668;
  wire [7:0] add_961671;
  wire [7:0] sel_961672;
  wire [7:0] add_961675;
  wire [7:0] sel_961676;
  wire [7:0] add_961679;
  wire [7:0] sel_961680;
  wire [7:0] add_961683;
  wire [7:0] sel_961684;
  wire [7:0] add_961687;
  wire [7:0] sel_961688;
  wire [7:0] add_961691;
  wire [7:0] sel_961692;
  wire [7:0] add_961695;
  wire [7:0] sel_961696;
  wire [7:0] add_961699;
  wire [7:0] sel_961700;
  wire [7:0] add_961703;
  wire [7:0] sel_961704;
  wire [7:0] add_961707;
  wire [7:0] sel_961708;
  wire [7:0] add_961711;
  wire [7:0] sel_961712;
  wire [7:0] add_961715;
  wire [7:0] sel_961716;
  wire [7:0] add_961719;
  wire [7:0] sel_961720;
  wire [7:0] add_961723;
  wire [7:0] sel_961724;
  wire [7:0] add_961727;
  wire [7:0] sel_961728;
  wire [7:0] add_961731;
  wire [7:0] sel_961732;
  wire [7:0] add_961735;
  wire [7:0] sel_961736;
  wire [7:0] add_961739;
  wire [7:0] sel_961740;
  wire [7:0] add_961743;
  wire [7:0] sel_961744;
  wire [7:0] add_961747;
  wire [7:0] sel_961748;
  wire [7:0] add_961751;
  wire [7:0] sel_961752;
  wire [7:0] add_961755;
  wire [7:0] sel_961756;
  wire [7:0] add_961759;
  wire [7:0] sel_961760;
  wire [7:0] add_961763;
  wire [7:0] sel_961764;
  wire [7:0] add_961767;
  wire [7:0] sel_961768;
  wire [7:0] add_961771;
  wire [7:0] sel_961772;
  wire [7:0] add_961775;
  wire [7:0] sel_961776;
  wire [7:0] add_961779;
  wire [7:0] sel_961780;
  wire [7:0] add_961783;
  wire [7:0] sel_961784;
  wire [7:0] add_961787;
  wire [7:0] sel_961788;
  wire [7:0] add_961791;
  wire [7:0] sel_961792;
  wire [7:0] add_961795;
  wire [7:0] sel_961796;
  wire [7:0] add_961799;
  wire [7:0] sel_961800;
  wire [7:0] add_961803;
  wire [7:0] sel_961804;
  wire [7:0] add_961807;
  wire [7:0] sel_961808;
  wire [7:0] add_961811;
  wire [7:0] sel_961812;
  wire [7:0] add_961815;
  wire [7:0] sel_961816;
  wire [7:0] add_961819;
  wire [7:0] sel_961820;
  wire [7:0] add_961823;
  wire [7:0] sel_961824;
  wire [7:0] add_961827;
  wire [7:0] sel_961828;
  wire [7:0] add_961831;
  wire [7:0] sel_961832;
  wire [7:0] add_961835;
  wire [7:0] sel_961836;
  wire [7:0] add_961839;
  wire [7:0] sel_961840;
  wire [7:0] add_961843;
  wire [7:0] sel_961844;
  wire [7:0] add_961847;
  wire [7:0] sel_961848;
  wire [7:0] add_961851;
  wire [7:0] sel_961852;
  wire [7:0] add_961855;
  wire [7:0] sel_961856;
  wire [7:0] add_961859;
  wire [7:0] sel_961860;
  wire [7:0] add_961863;
  wire [7:0] sel_961864;
  wire [7:0] add_961867;
  wire [7:0] sel_961868;
  wire [7:0] add_961871;
  wire [7:0] sel_961872;
  wire [7:0] add_961875;
  wire [7:0] sel_961876;
  wire [7:0] add_961879;
  wire [7:0] sel_961880;
  wire [7:0] add_961883;
  wire [7:0] sel_961884;
  wire [7:0] add_961887;
  wire [7:0] sel_961888;
  wire [7:0] add_961891;
  wire [7:0] sel_961892;
  wire [7:0] add_961895;
  wire [7:0] sel_961896;
  wire [7:0] add_961899;
  wire [7:0] sel_961900;
  wire [7:0] add_961903;
  wire [7:0] sel_961904;
  wire [7:0] add_961907;
  wire [7:0] sel_961908;
  wire [7:0] add_961911;
  wire [7:0] sel_961912;
  wire [7:0] add_961915;
  wire [7:0] sel_961916;
  wire [7:0] add_961919;
  wire [7:0] sel_961920;
  wire [7:0] add_961923;
  wire [7:0] sel_961924;
  wire [7:0] add_961927;
  wire [7:0] sel_961928;
  wire [7:0] add_961931;
  wire [7:0] sel_961932;
  wire [7:0] add_961935;
  wire [7:0] sel_961936;
  wire [7:0] add_961939;
  wire [7:0] sel_961940;
  wire [7:0] add_961943;
  wire [7:0] sel_961944;
  wire [7:0] add_961947;
  wire [7:0] sel_961948;
  wire [7:0] add_961951;
  wire [7:0] sel_961952;
  wire [7:0] add_961956;
  wire [15:0] array_index_961957;
  wire [7:0] sel_961958;
  wire [7:0] add_961961;
  wire [7:0] sel_961962;
  wire [7:0] add_961965;
  wire [7:0] sel_961966;
  wire [7:0] add_961969;
  wire [7:0] sel_961970;
  wire [7:0] add_961973;
  wire [7:0] sel_961974;
  wire [7:0] add_961977;
  wire [7:0] sel_961978;
  wire [7:0] add_961981;
  wire [7:0] sel_961982;
  wire [7:0] add_961985;
  wire [7:0] sel_961986;
  wire [7:0] add_961989;
  wire [7:0] sel_961990;
  wire [7:0] add_961993;
  wire [7:0] sel_961994;
  wire [7:0] add_961997;
  wire [7:0] sel_961998;
  wire [7:0] add_962001;
  wire [7:0] sel_962002;
  wire [7:0] add_962005;
  wire [7:0] sel_962006;
  wire [7:0] add_962009;
  wire [7:0] sel_962010;
  wire [7:0] add_962013;
  wire [7:0] sel_962014;
  wire [7:0] add_962017;
  wire [7:0] sel_962018;
  wire [7:0] add_962021;
  wire [7:0] sel_962022;
  wire [7:0] add_962025;
  wire [7:0] sel_962026;
  wire [7:0] add_962029;
  wire [7:0] sel_962030;
  wire [7:0] add_962033;
  wire [7:0] sel_962034;
  wire [7:0] add_962037;
  wire [7:0] sel_962038;
  wire [7:0] add_962041;
  wire [7:0] sel_962042;
  wire [7:0] add_962045;
  wire [7:0] sel_962046;
  wire [7:0] add_962049;
  wire [7:0] sel_962050;
  wire [7:0] add_962053;
  wire [7:0] sel_962054;
  wire [7:0] add_962057;
  wire [7:0] sel_962058;
  wire [7:0] add_962061;
  wire [7:0] sel_962062;
  wire [7:0] add_962065;
  wire [7:0] sel_962066;
  wire [7:0] add_962069;
  wire [7:0] sel_962070;
  wire [7:0] add_962073;
  wire [7:0] sel_962074;
  wire [7:0] add_962077;
  wire [7:0] sel_962078;
  wire [7:0] add_962081;
  wire [7:0] sel_962082;
  wire [7:0] add_962085;
  wire [7:0] sel_962086;
  wire [7:0] add_962089;
  wire [7:0] sel_962090;
  wire [7:0] add_962093;
  wire [7:0] sel_962094;
  wire [7:0] add_962097;
  wire [7:0] sel_962098;
  wire [7:0] add_962101;
  wire [7:0] sel_962102;
  wire [7:0] add_962105;
  wire [7:0] sel_962106;
  wire [7:0] add_962109;
  wire [7:0] sel_962110;
  wire [7:0] add_962113;
  wire [7:0] sel_962114;
  wire [7:0] add_962117;
  wire [7:0] sel_962118;
  wire [7:0] add_962121;
  wire [7:0] sel_962122;
  wire [7:0] add_962125;
  wire [7:0] sel_962126;
  wire [7:0] add_962129;
  wire [7:0] sel_962130;
  wire [7:0] add_962133;
  wire [7:0] sel_962134;
  wire [7:0] add_962137;
  wire [7:0] sel_962138;
  wire [7:0] add_962141;
  wire [7:0] sel_962142;
  wire [7:0] add_962145;
  wire [7:0] sel_962146;
  wire [7:0] add_962149;
  wire [7:0] sel_962150;
  wire [7:0] add_962153;
  wire [7:0] sel_962154;
  wire [7:0] add_962157;
  wire [7:0] sel_962158;
  wire [7:0] add_962161;
  wire [7:0] sel_962162;
  wire [7:0] add_962165;
  wire [7:0] sel_962166;
  wire [7:0] add_962169;
  wire [7:0] sel_962170;
  wire [7:0] add_962173;
  wire [7:0] sel_962174;
  wire [7:0] add_962177;
  wire [7:0] sel_962178;
  wire [7:0] add_962181;
  wire [7:0] sel_962182;
  wire [7:0] add_962185;
  wire [7:0] sel_962186;
  wire [7:0] add_962189;
  wire [7:0] sel_962190;
  wire [7:0] add_962193;
  wire [7:0] sel_962194;
  wire [7:0] add_962197;
  wire [7:0] sel_962198;
  wire [7:0] add_962201;
  wire [7:0] sel_962202;
  wire [7:0] add_962205;
  wire [7:0] sel_962206;
  wire [7:0] add_962209;
  wire [7:0] sel_962210;
  wire [7:0] add_962213;
  wire [7:0] sel_962214;
  wire [7:0] add_962217;
  wire [7:0] sel_962218;
  wire [7:0] add_962221;
  wire [7:0] sel_962222;
  wire [7:0] add_962225;
  wire [7:0] sel_962226;
  wire [7:0] add_962229;
  wire [7:0] sel_962230;
  wire [7:0] add_962233;
  wire [7:0] sel_962234;
  wire [7:0] add_962237;
  wire [7:0] sel_962238;
  wire [7:0] add_962241;
  wire [7:0] sel_962242;
  wire [7:0] add_962245;
  wire [7:0] sel_962246;
  wire [7:0] add_962249;
  wire [7:0] sel_962250;
  wire [7:0] add_962253;
  wire [7:0] sel_962254;
  wire [7:0] add_962257;
  wire [7:0] sel_962258;
  wire [7:0] add_962261;
  wire [7:0] sel_962262;
  wire [7:0] add_962265;
  wire [7:0] sel_962266;
  wire [7:0] add_962269;
  wire [7:0] sel_962270;
  wire [7:0] add_962273;
  wire [7:0] sel_962274;
  wire [7:0] add_962277;
  wire [7:0] sel_962278;
  wire [7:0] add_962281;
  wire [7:0] sel_962282;
  wire [7:0] add_962285;
  wire [7:0] sel_962286;
  wire [7:0] add_962289;
  wire [7:0] sel_962290;
  wire [7:0] add_962293;
  wire [7:0] sel_962294;
  wire [7:0] add_962297;
  wire [7:0] sel_962298;
  wire [7:0] add_962301;
  wire [7:0] sel_962302;
  wire [7:0] add_962305;
  wire [7:0] sel_962306;
  wire [7:0] add_962309;
  wire [7:0] sel_962310;
  wire [7:0] add_962313;
  wire [7:0] sel_962314;
  wire [7:0] add_962317;
  wire [7:0] sel_962318;
  wire [7:0] add_962321;
  wire [7:0] sel_962322;
  wire [7:0] add_962325;
  wire [7:0] sel_962326;
  wire [7:0] add_962329;
  wire [7:0] sel_962330;
  wire [7:0] add_962333;
  wire [7:0] sel_962334;
  wire [7:0] add_962337;
  wire [7:0] sel_962338;
  wire [7:0] add_962341;
  wire [7:0] sel_962342;
  wire [7:0] add_962345;
  wire [7:0] sel_962346;
  wire [7:0] add_962349;
  wire [7:0] sel_962350;
  wire [7:0] add_962353;
  wire [7:0] sel_962354;
  wire [7:0] add_962358;
  wire [15:0] array_index_962359;
  wire [7:0] sel_962360;
  wire [7:0] add_962363;
  wire [7:0] sel_962364;
  wire [7:0] add_962367;
  wire [7:0] sel_962368;
  wire [7:0] add_962371;
  wire [7:0] sel_962372;
  wire [7:0] add_962375;
  wire [7:0] sel_962376;
  wire [7:0] add_962379;
  wire [7:0] sel_962380;
  wire [7:0] add_962383;
  wire [7:0] sel_962384;
  wire [7:0] add_962387;
  wire [7:0] sel_962388;
  wire [7:0] add_962391;
  wire [7:0] sel_962392;
  wire [7:0] add_962395;
  wire [7:0] sel_962396;
  wire [7:0] add_962399;
  wire [7:0] sel_962400;
  wire [7:0] add_962403;
  wire [7:0] sel_962404;
  wire [7:0] add_962407;
  wire [7:0] sel_962408;
  wire [7:0] add_962411;
  wire [7:0] sel_962412;
  wire [7:0] add_962415;
  wire [7:0] sel_962416;
  wire [7:0] add_962419;
  wire [7:0] sel_962420;
  wire [7:0] add_962423;
  wire [7:0] sel_962424;
  wire [7:0] add_962427;
  wire [7:0] sel_962428;
  wire [7:0] add_962431;
  wire [7:0] sel_962432;
  wire [7:0] add_962435;
  wire [7:0] sel_962436;
  wire [7:0] add_962439;
  wire [7:0] sel_962440;
  wire [7:0] add_962443;
  wire [7:0] sel_962444;
  wire [7:0] add_962447;
  wire [7:0] sel_962448;
  wire [7:0] add_962451;
  wire [7:0] sel_962452;
  wire [7:0] add_962455;
  wire [7:0] sel_962456;
  wire [7:0] add_962459;
  wire [7:0] sel_962460;
  wire [7:0] add_962463;
  wire [7:0] sel_962464;
  wire [7:0] add_962467;
  wire [7:0] sel_962468;
  wire [7:0] add_962471;
  wire [7:0] sel_962472;
  wire [7:0] add_962475;
  wire [7:0] sel_962476;
  wire [7:0] add_962479;
  wire [7:0] sel_962480;
  wire [7:0] add_962483;
  wire [7:0] sel_962484;
  wire [7:0] add_962487;
  wire [7:0] sel_962488;
  wire [7:0] add_962491;
  wire [7:0] sel_962492;
  wire [7:0] add_962495;
  wire [7:0] sel_962496;
  wire [7:0] add_962499;
  wire [7:0] sel_962500;
  wire [7:0] add_962503;
  wire [7:0] sel_962504;
  wire [7:0] add_962507;
  wire [7:0] sel_962508;
  wire [7:0] add_962511;
  wire [7:0] sel_962512;
  wire [7:0] add_962515;
  wire [7:0] sel_962516;
  wire [7:0] add_962519;
  wire [7:0] sel_962520;
  wire [7:0] add_962523;
  wire [7:0] sel_962524;
  wire [7:0] add_962527;
  wire [7:0] sel_962528;
  wire [7:0] add_962531;
  wire [7:0] sel_962532;
  wire [7:0] add_962535;
  wire [7:0] sel_962536;
  wire [7:0] add_962539;
  wire [7:0] sel_962540;
  wire [7:0] add_962543;
  wire [7:0] sel_962544;
  wire [7:0] add_962547;
  wire [7:0] sel_962548;
  wire [7:0] add_962551;
  wire [7:0] sel_962552;
  wire [7:0] add_962555;
  wire [7:0] sel_962556;
  wire [7:0] add_962559;
  wire [7:0] sel_962560;
  wire [7:0] add_962563;
  wire [7:0] sel_962564;
  wire [7:0] add_962567;
  wire [7:0] sel_962568;
  wire [7:0] add_962571;
  wire [7:0] sel_962572;
  wire [7:0] add_962575;
  wire [7:0] sel_962576;
  wire [7:0] add_962579;
  wire [7:0] sel_962580;
  wire [7:0] add_962583;
  wire [7:0] sel_962584;
  wire [7:0] add_962587;
  wire [7:0] sel_962588;
  wire [7:0] add_962591;
  wire [7:0] sel_962592;
  wire [7:0] add_962595;
  wire [7:0] sel_962596;
  wire [7:0] add_962599;
  wire [7:0] sel_962600;
  wire [7:0] add_962603;
  wire [7:0] sel_962604;
  wire [7:0] add_962607;
  wire [7:0] sel_962608;
  wire [7:0] add_962611;
  wire [7:0] sel_962612;
  wire [7:0] add_962615;
  wire [7:0] sel_962616;
  wire [7:0] add_962619;
  wire [7:0] sel_962620;
  wire [7:0] add_962623;
  wire [7:0] sel_962624;
  wire [7:0] add_962627;
  wire [7:0] sel_962628;
  wire [7:0] add_962631;
  wire [7:0] sel_962632;
  wire [7:0] add_962635;
  wire [7:0] sel_962636;
  wire [7:0] add_962639;
  wire [7:0] sel_962640;
  wire [7:0] add_962643;
  wire [7:0] sel_962644;
  wire [7:0] add_962647;
  wire [7:0] sel_962648;
  wire [7:0] add_962651;
  wire [7:0] sel_962652;
  wire [7:0] add_962655;
  wire [7:0] sel_962656;
  wire [7:0] add_962659;
  wire [7:0] sel_962660;
  wire [7:0] add_962663;
  wire [7:0] sel_962664;
  wire [7:0] add_962667;
  wire [7:0] sel_962668;
  wire [7:0] add_962671;
  wire [7:0] sel_962672;
  wire [7:0] add_962675;
  wire [7:0] sel_962676;
  wire [7:0] add_962679;
  wire [7:0] sel_962680;
  wire [7:0] add_962683;
  wire [7:0] sel_962684;
  wire [7:0] add_962687;
  wire [7:0] sel_962688;
  wire [7:0] add_962691;
  wire [7:0] sel_962692;
  wire [7:0] add_962695;
  wire [7:0] sel_962696;
  wire [7:0] add_962699;
  wire [7:0] sel_962700;
  wire [7:0] add_962703;
  wire [7:0] sel_962704;
  wire [7:0] add_962707;
  wire [7:0] sel_962708;
  wire [7:0] add_962711;
  wire [7:0] sel_962712;
  wire [7:0] add_962715;
  wire [7:0] sel_962716;
  wire [7:0] add_962719;
  wire [7:0] sel_962720;
  wire [7:0] add_962723;
  wire [7:0] sel_962724;
  wire [7:0] add_962727;
  wire [7:0] sel_962728;
  wire [7:0] add_962731;
  wire [7:0] sel_962732;
  wire [7:0] add_962735;
  wire [7:0] sel_962736;
  wire [7:0] add_962739;
  wire [7:0] sel_962740;
  wire [7:0] add_962743;
  wire [7:0] sel_962744;
  wire [7:0] add_962747;
  wire [7:0] sel_962748;
  wire [7:0] add_962751;
  wire [7:0] sel_962752;
  wire [7:0] add_962755;
  wire [7:0] sel_962756;
  wire [7:0] add_962760;
  wire [15:0] array_index_962761;
  wire [7:0] sel_962762;
  wire [7:0] add_962765;
  wire [7:0] sel_962766;
  wire [7:0] add_962769;
  wire [7:0] sel_962770;
  wire [7:0] add_962773;
  wire [7:0] sel_962774;
  wire [7:0] add_962777;
  wire [7:0] sel_962778;
  wire [7:0] add_962781;
  wire [7:0] sel_962782;
  wire [7:0] add_962785;
  wire [7:0] sel_962786;
  wire [7:0] add_962789;
  wire [7:0] sel_962790;
  wire [7:0] add_962793;
  wire [7:0] sel_962794;
  wire [7:0] add_962797;
  wire [7:0] sel_962798;
  wire [7:0] add_962801;
  wire [7:0] sel_962802;
  wire [7:0] add_962805;
  wire [7:0] sel_962806;
  wire [7:0] add_962809;
  wire [7:0] sel_962810;
  wire [7:0] add_962813;
  wire [7:0] sel_962814;
  wire [7:0] add_962817;
  wire [7:0] sel_962818;
  wire [7:0] add_962821;
  wire [7:0] sel_962822;
  wire [7:0] add_962825;
  wire [7:0] sel_962826;
  wire [7:0] add_962829;
  wire [7:0] sel_962830;
  wire [7:0] add_962833;
  wire [7:0] sel_962834;
  wire [7:0] add_962837;
  wire [7:0] sel_962838;
  wire [7:0] add_962841;
  wire [7:0] sel_962842;
  wire [7:0] add_962845;
  wire [7:0] sel_962846;
  wire [7:0] add_962849;
  wire [7:0] sel_962850;
  wire [7:0] add_962853;
  wire [7:0] sel_962854;
  wire [7:0] add_962857;
  wire [7:0] sel_962858;
  wire [7:0] add_962861;
  wire [7:0] sel_962862;
  wire [7:0] add_962865;
  wire [7:0] sel_962866;
  wire [7:0] add_962869;
  wire [7:0] sel_962870;
  wire [7:0] add_962873;
  wire [7:0] sel_962874;
  wire [7:0] add_962877;
  wire [7:0] sel_962878;
  wire [7:0] add_962881;
  wire [7:0] sel_962882;
  wire [7:0] add_962885;
  wire [7:0] sel_962886;
  wire [7:0] add_962889;
  wire [7:0] sel_962890;
  wire [7:0] add_962893;
  wire [7:0] sel_962894;
  wire [7:0] add_962897;
  wire [7:0] sel_962898;
  wire [7:0] add_962901;
  wire [7:0] sel_962902;
  wire [7:0] add_962905;
  wire [7:0] sel_962906;
  wire [7:0] add_962909;
  wire [7:0] sel_962910;
  wire [7:0] add_962913;
  wire [7:0] sel_962914;
  wire [7:0] add_962917;
  wire [7:0] sel_962918;
  wire [7:0] add_962921;
  wire [7:0] sel_962922;
  wire [7:0] add_962925;
  wire [7:0] sel_962926;
  wire [7:0] add_962929;
  wire [7:0] sel_962930;
  wire [7:0] add_962933;
  wire [7:0] sel_962934;
  wire [7:0] add_962937;
  wire [7:0] sel_962938;
  wire [7:0] add_962941;
  wire [7:0] sel_962942;
  wire [7:0] add_962945;
  wire [7:0] sel_962946;
  wire [7:0] add_962949;
  wire [7:0] sel_962950;
  wire [7:0] add_962953;
  wire [7:0] sel_962954;
  wire [7:0] add_962957;
  wire [7:0] sel_962958;
  wire [7:0] add_962961;
  wire [7:0] sel_962962;
  wire [7:0] add_962965;
  wire [7:0] sel_962966;
  wire [7:0] add_962969;
  wire [7:0] sel_962970;
  wire [7:0] add_962973;
  wire [7:0] sel_962974;
  wire [7:0] add_962977;
  wire [7:0] sel_962978;
  wire [7:0] add_962981;
  wire [7:0] sel_962982;
  wire [7:0] add_962985;
  wire [7:0] sel_962986;
  wire [7:0] add_962989;
  wire [7:0] sel_962990;
  wire [7:0] add_962993;
  wire [7:0] sel_962994;
  wire [7:0] add_962997;
  wire [7:0] sel_962998;
  wire [7:0] add_963001;
  wire [7:0] sel_963002;
  wire [7:0] add_963005;
  wire [7:0] sel_963006;
  wire [7:0] add_963009;
  wire [7:0] sel_963010;
  wire [7:0] add_963013;
  wire [7:0] sel_963014;
  wire [7:0] add_963017;
  wire [7:0] sel_963018;
  wire [7:0] add_963021;
  wire [7:0] sel_963022;
  wire [7:0] add_963025;
  wire [7:0] sel_963026;
  wire [7:0] add_963029;
  wire [7:0] sel_963030;
  wire [7:0] add_963033;
  wire [7:0] sel_963034;
  wire [7:0] add_963037;
  wire [7:0] sel_963038;
  wire [7:0] add_963041;
  wire [7:0] sel_963042;
  wire [7:0] add_963045;
  wire [7:0] sel_963046;
  wire [7:0] add_963049;
  wire [7:0] sel_963050;
  wire [7:0] add_963053;
  wire [7:0] sel_963054;
  wire [7:0] add_963057;
  wire [7:0] sel_963058;
  wire [7:0] add_963061;
  wire [7:0] sel_963062;
  wire [7:0] add_963065;
  wire [7:0] sel_963066;
  wire [7:0] add_963069;
  wire [7:0] sel_963070;
  wire [7:0] add_963073;
  wire [7:0] sel_963074;
  wire [7:0] add_963077;
  wire [7:0] sel_963078;
  wire [7:0] add_963081;
  wire [7:0] sel_963082;
  wire [7:0] add_963085;
  wire [7:0] sel_963086;
  wire [7:0] add_963089;
  wire [7:0] sel_963090;
  wire [7:0] add_963093;
  wire [7:0] sel_963094;
  wire [7:0] add_963097;
  wire [7:0] sel_963098;
  wire [7:0] add_963101;
  wire [7:0] sel_963102;
  wire [7:0] add_963105;
  wire [7:0] sel_963106;
  wire [7:0] add_963109;
  wire [7:0] sel_963110;
  wire [7:0] add_963113;
  wire [7:0] sel_963114;
  wire [7:0] add_963117;
  wire [7:0] sel_963118;
  wire [7:0] add_963121;
  wire [7:0] sel_963122;
  wire [7:0] add_963125;
  wire [7:0] sel_963126;
  wire [7:0] add_963129;
  wire [7:0] sel_963130;
  wire [7:0] add_963133;
  wire [7:0] sel_963134;
  wire [7:0] add_963137;
  wire [7:0] sel_963138;
  wire [7:0] add_963141;
  wire [7:0] sel_963142;
  wire [7:0] add_963145;
  wire [7:0] sel_963146;
  wire [7:0] add_963149;
  wire [7:0] sel_963150;
  wire [7:0] add_963153;
  wire [7:0] sel_963154;
  wire [7:0] add_963157;
  wire [7:0] sel_963158;
  wire [7:0] add_963162;
  wire [15:0] array_index_963163;
  wire [7:0] sel_963164;
  wire [7:0] add_963167;
  wire [7:0] sel_963168;
  wire [7:0] add_963171;
  wire [7:0] sel_963172;
  wire [7:0] add_963175;
  wire [7:0] sel_963176;
  wire [7:0] add_963179;
  wire [7:0] sel_963180;
  wire [7:0] add_963183;
  wire [7:0] sel_963184;
  wire [7:0] add_963187;
  wire [7:0] sel_963188;
  wire [7:0] add_963191;
  wire [7:0] sel_963192;
  wire [7:0] add_963195;
  wire [7:0] sel_963196;
  wire [7:0] add_963199;
  wire [7:0] sel_963200;
  wire [7:0] add_963203;
  wire [7:0] sel_963204;
  wire [7:0] add_963207;
  wire [7:0] sel_963208;
  wire [7:0] add_963211;
  wire [7:0] sel_963212;
  wire [7:0] add_963215;
  wire [7:0] sel_963216;
  wire [7:0] add_963219;
  wire [7:0] sel_963220;
  wire [7:0] add_963223;
  wire [7:0] sel_963224;
  wire [7:0] add_963227;
  wire [7:0] sel_963228;
  wire [7:0] add_963231;
  wire [7:0] sel_963232;
  wire [7:0] add_963235;
  wire [7:0] sel_963236;
  wire [7:0] add_963239;
  wire [7:0] sel_963240;
  wire [7:0] add_963243;
  wire [7:0] sel_963244;
  wire [7:0] add_963247;
  wire [7:0] sel_963248;
  wire [7:0] add_963251;
  wire [7:0] sel_963252;
  wire [7:0] add_963255;
  wire [7:0] sel_963256;
  wire [7:0] add_963259;
  wire [7:0] sel_963260;
  wire [7:0] add_963263;
  wire [7:0] sel_963264;
  wire [7:0] add_963267;
  wire [7:0] sel_963268;
  wire [7:0] add_963271;
  wire [7:0] sel_963272;
  wire [7:0] add_963275;
  wire [7:0] sel_963276;
  wire [7:0] add_963279;
  wire [7:0] sel_963280;
  wire [7:0] add_963283;
  wire [7:0] sel_963284;
  wire [7:0] add_963287;
  wire [7:0] sel_963288;
  wire [7:0] add_963291;
  wire [7:0] sel_963292;
  wire [7:0] add_963295;
  wire [7:0] sel_963296;
  wire [7:0] add_963299;
  wire [7:0] sel_963300;
  wire [7:0] add_963303;
  wire [7:0] sel_963304;
  wire [7:0] add_963307;
  wire [7:0] sel_963308;
  wire [7:0] add_963311;
  wire [7:0] sel_963312;
  wire [7:0] add_963315;
  wire [7:0] sel_963316;
  wire [7:0] add_963319;
  wire [7:0] sel_963320;
  wire [7:0] add_963323;
  wire [7:0] sel_963324;
  wire [7:0] add_963327;
  wire [7:0] sel_963328;
  wire [7:0] add_963331;
  wire [7:0] sel_963332;
  wire [7:0] add_963335;
  wire [7:0] sel_963336;
  wire [7:0] add_963339;
  wire [7:0] sel_963340;
  wire [7:0] add_963343;
  wire [7:0] sel_963344;
  wire [7:0] add_963347;
  wire [7:0] sel_963348;
  wire [7:0] add_963351;
  wire [7:0] sel_963352;
  wire [7:0] add_963355;
  wire [7:0] sel_963356;
  wire [7:0] add_963359;
  wire [7:0] sel_963360;
  wire [7:0] add_963363;
  wire [7:0] sel_963364;
  wire [7:0] add_963367;
  wire [7:0] sel_963368;
  wire [7:0] add_963371;
  wire [7:0] sel_963372;
  wire [7:0] add_963375;
  wire [7:0] sel_963376;
  wire [7:0] add_963379;
  wire [7:0] sel_963380;
  wire [7:0] add_963383;
  wire [7:0] sel_963384;
  wire [7:0] add_963387;
  wire [7:0] sel_963388;
  wire [7:0] add_963391;
  wire [7:0] sel_963392;
  wire [7:0] add_963395;
  wire [7:0] sel_963396;
  wire [7:0] add_963399;
  wire [7:0] sel_963400;
  wire [7:0] add_963403;
  wire [7:0] sel_963404;
  wire [7:0] add_963407;
  wire [7:0] sel_963408;
  wire [7:0] add_963411;
  wire [7:0] sel_963412;
  wire [7:0] add_963415;
  wire [7:0] sel_963416;
  wire [7:0] add_963419;
  wire [7:0] sel_963420;
  wire [7:0] add_963423;
  wire [7:0] sel_963424;
  wire [7:0] add_963427;
  wire [7:0] sel_963428;
  wire [7:0] add_963431;
  wire [7:0] sel_963432;
  wire [7:0] add_963435;
  wire [7:0] sel_963436;
  wire [7:0] add_963439;
  wire [7:0] sel_963440;
  wire [7:0] add_963443;
  wire [7:0] sel_963444;
  wire [7:0] add_963447;
  wire [7:0] sel_963448;
  wire [7:0] add_963451;
  wire [7:0] sel_963452;
  wire [7:0] add_963455;
  wire [7:0] sel_963456;
  wire [7:0] add_963459;
  wire [7:0] sel_963460;
  wire [7:0] add_963463;
  wire [7:0] sel_963464;
  wire [7:0] add_963467;
  wire [7:0] sel_963468;
  wire [7:0] add_963471;
  wire [7:0] sel_963472;
  wire [7:0] add_963475;
  wire [7:0] sel_963476;
  wire [7:0] add_963479;
  wire [7:0] sel_963480;
  wire [7:0] add_963483;
  wire [7:0] sel_963484;
  wire [7:0] add_963487;
  wire [7:0] sel_963488;
  wire [7:0] add_963491;
  wire [7:0] sel_963492;
  wire [7:0] add_963495;
  wire [7:0] sel_963496;
  wire [7:0] add_963499;
  wire [7:0] sel_963500;
  wire [7:0] add_963503;
  wire [7:0] sel_963504;
  wire [7:0] add_963507;
  wire [7:0] sel_963508;
  wire [7:0] add_963511;
  wire [7:0] sel_963512;
  wire [7:0] add_963515;
  wire [7:0] sel_963516;
  wire [7:0] add_963519;
  wire [7:0] sel_963520;
  wire [7:0] add_963523;
  wire [7:0] sel_963524;
  wire [7:0] add_963527;
  wire [7:0] sel_963528;
  wire [7:0] add_963531;
  wire [7:0] sel_963532;
  wire [7:0] add_963535;
  wire [7:0] sel_963536;
  wire [7:0] add_963539;
  wire [7:0] sel_963540;
  wire [7:0] add_963543;
  wire [7:0] sel_963544;
  wire [7:0] add_963547;
  wire [7:0] sel_963548;
  wire [7:0] add_963551;
  wire [7:0] sel_963552;
  wire [7:0] add_963555;
  wire [7:0] sel_963556;
  wire [7:0] add_963559;
  wire [7:0] sel_963560;
  wire [7:0] add_963564;
  wire [15:0] array_index_963565;
  wire [7:0] sel_963566;
  wire [7:0] add_963569;
  wire [7:0] sel_963570;
  wire [7:0] add_963573;
  wire [7:0] sel_963574;
  wire [7:0] add_963577;
  wire [7:0] sel_963578;
  wire [7:0] add_963581;
  wire [7:0] sel_963582;
  wire [7:0] add_963585;
  wire [7:0] sel_963586;
  wire [7:0] add_963589;
  wire [7:0] sel_963590;
  wire [7:0] add_963593;
  wire [7:0] sel_963594;
  wire [7:0] add_963597;
  wire [7:0] sel_963598;
  wire [7:0] add_963601;
  wire [7:0] sel_963602;
  wire [7:0] add_963605;
  wire [7:0] sel_963606;
  wire [7:0] add_963609;
  wire [7:0] sel_963610;
  wire [7:0] add_963613;
  wire [7:0] sel_963614;
  wire [7:0] add_963617;
  wire [7:0] sel_963618;
  wire [7:0] add_963621;
  wire [7:0] sel_963622;
  wire [7:0] add_963625;
  wire [7:0] sel_963626;
  wire [7:0] add_963629;
  wire [7:0] sel_963630;
  wire [7:0] add_963633;
  wire [7:0] sel_963634;
  wire [7:0] add_963637;
  wire [7:0] sel_963638;
  wire [7:0] add_963641;
  wire [7:0] sel_963642;
  wire [7:0] add_963645;
  wire [7:0] sel_963646;
  wire [7:0] add_963649;
  wire [7:0] sel_963650;
  wire [7:0] add_963653;
  wire [7:0] sel_963654;
  wire [7:0] add_963657;
  wire [7:0] sel_963658;
  wire [7:0] add_963661;
  wire [7:0] sel_963662;
  wire [7:0] add_963665;
  wire [7:0] sel_963666;
  wire [7:0] add_963669;
  wire [7:0] sel_963670;
  wire [7:0] add_963673;
  wire [7:0] sel_963674;
  wire [7:0] add_963677;
  wire [7:0] sel_963678;
  wire [7:0] add_963681;
  wire [7:0] sel_963682;
  wire [7:0] add_963685;
  wire [7:0] sel_963686;
  wire [7:0] add_963689;
  wire [7:0] sel_963690;
  wire [7:0] add_963693;
  wire [7:0] sel_963694;
  wire [7:0] add_963697;
  wire [7:0] sel_963698;
  wire [7:0] add_963701;
  wire [7:0] sel_963702;
  wire [7:0] add_963705;
  wire [7:0] sel_963706;
  wire [7:0] add_963709;
  wire [7:0] sel_963710;
  wire [7:0] add_963713;
  wire [7:0] sel_963714;
  wire [7:0] add_963717;
  wire [7:0] sel_963718;
  wire [7:0] add_963721;
  wire [7:0] sel_963722;
  wire [7:0] add_963725;
  wire [7:0] sel_963726;
  wire [7:0] add_963729;
  wire [7:0] sel_963730;
  wire [7:0] add_963733;
  wire [7:0] sel_963734;
  wire [7:0] add_963737;
  wire [7:0] sel_963738;
  wire [7:0] add_963741;
  wire [7:0] sel_963742;
  wire [7:0] add_963745;
  wire [7:0] sel_963746;
  wire [7:0] add_963749;
  wire [7:0] sel_963750;
  wire [7:0] add_963753;
  wire [7:0] sel_963754;
  wire [7:0] add_963757;
  wire [7:0] sel_963758;
  wire [7:0] add_963761;
  wire [7:0] sel_963762;
  wire [7:0] add_963765;
  wire [7:0] sel_963766;
  wire [7:0] add_963769;
  wire [7:0] sel_963770;
  wire [7:0] add_963773;
  wire [7:0] sel_963774;
  wire [7:0] add_963777;
  wire [7:0] sel_963778;
  wire [7:0] add_963781;
  wire [7:0] sel_963782;
  wire [7:0] add_963785;
  wire [7:0] sel_963786;
  wire [7:0] add_963789;
  wire [7:0] sel_963790;
  wire [7:0] add_963793;
  wire [7:0] sel_963794;
  wire [7:0] add_963797;
  wire [7:0] sel_963798;
  wire [7:0] add_963801;
  wire [7:0] sel_963802;
  wire [7:0] add_963805;
  wire [7:0] sel_963806;
  wire [7:0] add_963809;
  wire [7:0] sel_963810;
  wire [7:0] add_963813;
  wire [7:0] sel_963814;
  wire [7:0] add_963817;
  wire [7:0] sel_963818;
  wire [7:0] add_963821;
  wire [7:0] sel_963822;
  wire [7:0] add_963825;
  wire [7:0] sel_963826;
  wire [7:0] add_963829;
  wire [7:0] sel_963830;
  wire [7:0] add_963833;
  wire [7:0] sel_963834;
  wire [7:0] add_963837;
  wire [7:0] sel_963838;
  wire [7:0] add_963841;
  wire [7:0] sel_963842;
  wire [7:0] add_963845;
  wire [7:0] sel_963846;
  wire [7:0] add_963849;
  wire [7:0] sel_963850;
  wire [7:0] add_963853;
  wire [7:0] sel_963854;
  wire [7:0] add_963857;
  wire [7:0] sel_963858;
  wire [7:0] add_963861;
  wire [7:0] sel_963862;
  wire [7:0] add_963865;
  wire [7:0] sel_963866;
  wire [7:0] add_963869;
  wire [7:0] sel_963870;
  wire [7:0] add_963873;
  wire [7:0] sel_963874;
  wire [7:0] add_963877;
  wire [7:0] sel_963878;
  wire [7:0] add_963881;
  wire [7:0] sel_963882;
  wire [7:0] add_963885;
  wire [7:0] sel_963886;
  wire [7:0] add_963889;
  wire [7:0] sel_963890;
  wire [7:0] add_963893;
  wire [7:0] sel_963894;
  wire [7:0] add_963897;
  wire [7:0] sel_963898;
  wire [7:0] add_963901;
  wire [7:0] sel_963902;
  wire [7:0] add_963905;
  wire [7:0] sel_963906;
  wire [7:0] add_963909;
  wire [7:0] sel_963910;
  wire [7:0] add_963913;
  wire [7:0] sel_963914;
  wire [7:0] add_963917;
  wire [7:0] sel_963918;
  wire [7:0] add_963921;
  wire [7:0] sel_963922;
  wire [7:0] add_963925;
  wire [7:0] sel_963926;
  wire [7:0] add_963929;
  wire [7:0] sel_963930;
  wire [7:0] add_963933;
  wire [7:0] sel_963934;
  wire [7:0] add_963937;
  wire [7:0] sel_963938;
  wire [7:0] add_963941;
  wire [7:0] sel_963942;
  wire [7:0] add_963945;
  wire [7:0] sel_963946;
  wire [7:0] add_963949;
  wire [7:0] sel_963950;
  wire [7:0] add_963953;
  wire [7:0] sel_963954;
  wire [7:0] add_963957;
  wire [7:0] sel_963958;
  wire [7:0] add_963961;
  wire [7:0] sel_963962;
  wire [7:0] add_963966;
  wire [15:0] array_index_963967;
  wire [7:0] sel_963968;
  wire [7:0] add_963971;
  wire [7:0] sel_963972;
  wire [7:0] add_963975;
  wire [7:0] sel_963976;
  wire [7:0] add_963979;
  wire [7:0] sel_963980;
  wire [7:0] add_963983;
  wire [7:0] sel_963984;
  wire [7:0] add_963987;
  wire [7:0] sel_963988;
  wire [7:0] add_963991;
  wire [7:0] sel_963992;
  wire [7:0] add_963995;
  wire [7:0] sel_963996;
  wire [7:0] add_963999;
  wire [7:0] sel_964000;
  wire [7:0] add_964003;
  wire [7:0] sel_964004;
  wire [7:0] add_964007;
  wire [7:0] sel_964008;
  wire [7:0] add_964011;
  wire [7:0] sel_964012;
  wire [7:0] add_964015;
  wire [7:0] sel_964016;
  wire [7:0] add_964019;
  wire [7:0] sel_964020;
  wire [7:0] add_964023;
  wire [7:0] sel_964024;
  wire [7:0] add_964027;
  wire [7:0] sel_964028;
  wire [7:0] add_964031;
  wire [7:0] sel_964032;
  wire [7:0] add_964035;
  wire [7:0] sel_964036;
  wire [7:0] add_964039;
  wire [7:0] sel_964040;
  wire [7:0] add_964043;
  wire [7:0] sel_964044;
  wire [7:0] add_964047;
  wire [7:0] sel_964048;
  wire [7:0] add_964051;
  wire [7:0] sel_964052;
  wire [7:0] add_964055;
  wire [7:0] sel_964056;
  wire [7:0] add_964059;
  wire [7:0] sel_964060;
  wire [7:0] add_964063;
  wire [7:0] sel_964064;
  wire [7:0] add_964067;
  wire [7:0] sel_964068;
  wire [7:0] add_964071;
  wire [7:0] sel_964072;
  wire [7:0] add_964075;
  wire [7:0] sel_964076;
  wire [7:0] add_964079;
  wire [7:0] sel_964080;
  wire [7:0] add_964083;
  wire [7:0] sel_964084;
  wire [7:0] add_964087;
  wire [7:0] sel_964088;
  wire [7:0] add_964091;
  wire [7:0] sel_964092;
  wire [7:0] add_964095;
  wire [7:0] sel_964096;
  wire [7:0] add_964099;
  wire [7:0] sel_964100;
  wire [7:0] add_964103;
  wire [7:0] sel_964104;
  wire [7:0] add_964107;
  wire [7:0] sel_964108;
  wire [7:0] add_964111;
  wire [7:0] sel_964112;
  wire [7:0] add_964115;
  wire [7:0] sel_964116;
  wire [7:0] add_964119;
  wire [7:0] sel_964120;
  wire [7:0] add_964123;
  wire [7:0] sel_964124;
  wire [7:0] add_964127;
  wire [7:0] sel_964128;
  wire [7:0] add_964131;
  wire [7:0] sel_964132;
  wire [7:0] add_964135;
  wire [7:0] sel_964136;
  wire [7:0] add_964139;
  wire [7:0] sel_964140;
  wire [7:0] add_964143;
  wire [7:0] sel_964144;
  wire [7:0] add_964147;
  wire [7:0] sel_964148;
  wire [7:0] add_964151;
  wire [7:0] sel_964152;
  wire [7:0] add_964155;
  wire [7:0] sel_964156;
  wire [7:0] add_964159;
  wire [7:0] sel_964160;
  wire [7:0] add_964163;
  wire [7:0] sel_964164;
  wire [7:0] add_964167;
  wire [7:0] sel_964168;
  wire [7:0] add_964171;
  wire [7:0] sel_964172;
  wire [7:0] add_964175;
  wire [7:0] sel_964176;
  wire [7:0] add_964179;
  wire [7:0] sel_964180;
  wire [7:0] add_964183;
  wire [7:0] sel_964184;
  wire [7:0] add_964187;
  wire [7:0] sel_964188;
  wire [7:0] add_964191;
  wire [7:0] sel_964192;
  wire [7:0] add_964195;
  wire [7:0] sel_964196;
  wire [7:0] add_964199;
  wire [7:0] sel_964200;
  wire [7:0] add_964203;
  wire [7:0] sel_964204;
  wire [7:0] add_964207;
  wire [7:0] sel_964208;
  wire [7:0] add_964211;
  wire [7:0] sel_964212;
  wire [7:0] add_964215;
  wire [7:0] sel_964216;
  wire [7:0] add_964219;
  wire [7:0] sel_964220;
  wire [7:0] add_964223;
  wire [7:0] sel_964224;
  wire [7:0] add_964227;
  wire [7:0] sel_964228;
  wire [7:0] add_964231;
  wire [7:0] sel_964232;
  wire [7:0] add_964235;
  wire [7:0] sel_964236;
  wire [7:0] add_964239;
  wire [7:0] sel_964240;
  wire [7:0] add_964243;
  wire [7:0] sel_964244;
  wire [7:0] add_964247;
  wire [7:0] sel_964248;
  wire [7:0] add_964251;
  wire [7:0] sel_964252;
  wire [7:0] add_964255;
  wire [7:0] sel_964256;
  wire [7:0] add_964259;
  wire [7:0] sel_964260;
  wire [7:0] add_964263;
  wire [7:0] sel_964264;
  wire [7:0] add_964267;
  wire [7:0] sel_964268;
  wire [7:0] add_964271;
  wire [7:0] sel_964272;
  wire [7:0] add_964275;
  wire [7:0] sel_964276;
  wire [7:0] add_964279;
  wire [7:0] sel_964280;
  wire [7:0] add_964283;
  wire [7:0] sel_964284;
  wire [7:0] add_964287;
  wire [7:0] sel_964288;
  wire [7:0] add_964291;
  wire [7:0] sel_964292;
  wire [7:0] add_964295;
  wire [7:0] sel_964296;
  wire [7:0] add_964299;
  wire [7:0] sel_964300;
  wire [7:0] add_964303;
  wire [7:0] sel_964304;
  wire [7:0] add_964307;
  wire [7:0] sel_964308;
  wire [7:0] add_964311;
  wire [7:0] sel_964312;
  wire [7:0] add_964315;
  wire [7:0] sel_964316;
  wire [7:0] add_964319;
  wire [7:0] sel_964320;
  wire [7:0] add_964323;
  wire [7:0] sel_964324;
  wire [7:0] add_964327;
  wire [7:0] sel_964328;
  wire [7:0] add_964331;
  wire [7:0] sel_964332;
  wire [7:0] add_964335;
  wire [7:0] sel_964336;
  wire [7:0] add_964339;
  wire [7:0] sel_964340;
  wire [7:0] add_964343;
  wire [7:0] sel_964344;
  wire [7:0] add_964347;
  wire [7:0] sel_964348;
  wire [7:0] add_964351;
  wire [7:0] sel_964352;
  wire [7:0] add_964355;
  wire [7:0] sel_964356;
  wire [7:0] add_964359;
  wire [7:0] sel_964360;
  wire [7:0] add_964363;
  wire [7:0] sel_964364;
  wire [7:0] add_964368;
  wire [15:0] array_index_964369;
  wire [7:0] sel_964370;
  wire [7:0] add_964373;
  wire [7:0] sel_964374;
  wire [7:0] add_964377;
  wire [7:0] sel_964378;
  wire [7:0] add_964381;
  wire [7:0] sel_964382;
  wire [7:0] add_964385;
  wire [7:0] sel_964386;
  wire [7:0] add_964389;
  wire [7:0] sel_964390;
  wire [7:0] add_964393;
  wire [7:0] sel_964394;
  wire [7:0] add_964397;
  wire [7:0] sel_964398;
  wire [7:0] add_964401;
  wire [7:0] sel_964402;
  wire [7:0] add_964405;
  wire [7:0] sel_964406;
  wire [7:0] add_964409;
  wire [7:0] sel_964410;
  wire [7:0] add_964413;
  wire [7:0] sel_964414;
  wire [7:0] add_964417;
  wire [7:0] sel_964418;
  wire [7:0] add_964421;
  wire [7:0] sel_964422;
  wire [7:0] add_964425;
  wire [7:0] sel_964426;
  wire [7:0] add_964429;
  wire [7:0] sel_964430;
  wire [7:0] add_964433;
  wire [7:0] sel_964434;
  wire [7:0] add_964437;
  wire [7:0] sel_964438;
  wire [7:0] add_964441;
  wire [7:0] sel_964442;
  wire [7:0] add_964445;
  wire [7:0] sel_964446;
  wire [7:0] add_964449;
  wire [7:0] sel_964450;
  wire [7:0] add_964453;
  wire [7:0] sel_964454;
  wire [7:0] add_964457;
  wire [7:0] sel_964458;
  wire [7:0] add_964461;
  wire [7:0] sel_964462;
  wire [7:0] add_964465;
  wire [7:0] sel_964466;
  wire [7:0] add_964469;
  wire [7:0] sel_964470;
  wire [7:0] add_964473;
  wire [7:0] sel_964474;
  wire [7:0] add_964477;
  wire [7:0] sel_964478;
  wire [7:0] add_964481;
  wire [7:0] sel_964482;
  wire [7:0] add_964485;
  wire [7:0] sel_964486;
  wire [7:0] add_964489;
  wire [7:0] sel_964490;
  wire [7:0] add_964493;
  wire [7:0] sel_964494;
  wire [7:0] add_964497;
  wire [7:0] sel_964498;
  wire [7:0] add_964501;
  wire [7:0] sel_964502;
  wire [7:0] add_964505;
  wire [7:0] sel_964506;
  wire [7:0] add_964509;
  wire [7:0] sel_964510;
  wire [7:0] add_964513;
  wire [7:0] sel_964514;
  wire [7:0] add_964517;
  wire [7:0] sel_964518;
  wire [7:0] add_964521;
  wire [7:0] sel_964522;
  wire [7:0] add_964525;
  wire [7:0] sel_964526;
  wire [7:0] add_964529;
  wire [7:0] sel_964530;
  wire [7:0] add_964533;
  wire [7:0] sel_964534;
  wire [7:0] add_964537;
  wire [7:0] sel_964538;
  wire [7:0] add_964541;
  wire [7:0] sel_964542;
  wire [7:0] add_964545;
  wire [7:0] sel_964546;
  wire [7:0] add_964549;
  wire [7:0] sel_964550;
  wire [7:0] add_964553;
  wire [7:0] sel_964554;
  wire [7:0] add_964557;
  wire [7:0] sel_964558;
  wire [7:0] add_964561;
  wire [7:0] sel_964562;
  wire [7:0] add_964565;
  wire [7:0] sel_964566;
  wire [7:0] add_964569;
  wire [7:0] sel_964570;
  wire [7:0] add_964573;
  wire [7:0] sel_964574;
  wire [7:0] add_964577;
  wire [7:0] sel_964578;
  wire [7:0] add_964581;
  wire [7:0] sel_964582;
  wire [7:0] add_964585;
  wire [7:0] sel_964586;
  wire [7:0] add_964589;
  wire [7:0] sel_964590;
  wire [7:0] add_964593;
  wire [7:0] sel_964594;
  wire [7:0] add_964597;
  wire [7:0] sel_964598;
  wire [7:0] add_964601;
  wire [7:0] sel_964602;
  wire [7:0] add_964605;
  wire [7:0] sel_964606;
  wire [7:0] add_964609;
  wire [7:0] sel_964610;
  wire [7:0] add_964613;
  wire [7:0] sel_964614;
  wire [7:0] add_964617;
  wire [7:0] sel_964618;
  wire [7:0] add_964621;
  wire [7:0] sel_964622;
  wire [7:0] add_964625;
  wire [7:0] sel_964626;
  wire [7:0] add_964629;
  wire [7:0] sel_964630;
  wire [7:0] add_964633;
  wire [7:0] sel_964634;
  wire [7:0] add_964637;
  wire [7:0] sel_964638;
  wire [7:0] add_964641;
  wire [7:0] sel_964642;
  wire [7:0] add_964645;
  wire [7:0] sel_964646;
  wire [7:0] add_964649;
  wire [7:0] sel_964650;
  wire [7:0] add_964653;
  wire [7:0] sel_964654;
  wire [7:0] add_964657;
  wire [7:0] sel_964658;
  wire [7:0] add_964661;
  wire [7:0] sel_964662;
  wire [7:0] add_964665;
  wire [7:0] sel_964666;
  wire [7:0] add_964669;
  wire [7:0] sel_964670;
  wire [7:0] add_964673;
  wire [7:0] sel_964674;
  wire [7:0] add_964677;
  wire [7:0] sel_964678;
  wire [7:0] add_964681;
  wire [7:0] sel_964682;
  wire [7:0] add_964685;
  wire [7:0] sel_964686;
  wire [7:0] add_964689;
  wire [7:0] sel_964690;
  wire [7:0] add_964693;
  wire [7:0] sel_964694;
  wire [7:0] add_964697;
  wire [7:0] sel_964698;
  wire [7:0] add_964701;
  wire [7:0] sel_964702;
  wire [7:0] add_964705;
  wire [7:0] sel_964706;
  wire [7:0] add_964709;
  wire [7:0] sel_964710;
  wire [7:0] add_964713;
  wire [7:0] sel_964714;
  wire [7:0] add_964717;
  wire [7:0] sel_964718;
  wire [7:0] add_964721;
  wire [7:0] sel_964722;
  wire [7:0] add_964725;
  wire [7:0] sel_964726;
  wire [7:0] add_964729;
  wire [7:0] sel_964730;
  wire [7:0] add_964733;
  wire [7:0] sel_964734;
  wire [7:0] add_964737;
  wire [7:0] sel_964738;
  wire [7:0] add_964741;
  wire [7:0] sel_964742;
  wire [7:0] add_964745;
  wire [7:0] sel_964746;
  wire [7:0] add_964749;
  wire [7:0] sel_964750;
  wire [7:0] add_964753;
  wire [7:0] sel_964754;
  wire [7:0] add_964757;
  wire [7:0] sel_964758;
  wire [7:0] add_964761;
  wire [7:0] sel_964762;
  wire [7:0] add_964765;
  wire [7:0] sel_964766;
  wire [7:0] add_964770;
  wire [15:0] array_index_964771;
  wire [7:0] sel_964772;
  wire [7:0] add_964775;
  wire [7:0] sel_964776;
  wire [7:0] add_964779;
  wire [7:0] sel_964780;
  wire [7:0] add_964783;
  wire [7:0] sel_964784;
  wire [7:0] add_964787;
  wire [7:0] sel_964788;
  wire [7:0] add_964791;
  wire [7:0] sel_964792;
  wire [7:0] add_964795;
  wire [7:0] sel_964796;
  wire [7:0] add_964799;
  wire [7:0] sel_964800;
  wire [7:0] add_964803;
  wire [7:0] sel_964804;
  wire [7:0] add_964807;
  wire [7:0] sel_964808;
  wire [7:0] add_964811;
  wire [7:0] sel_964812;
  wire [7:0] add_964815;
  wire [7:0] sel_964816;
  wire [7:0] add_964819;
  wire [7:0] sel_964820;
  wire [7:0] add_964823;
  wire [7:0] sel_964824;
  wire [7:0] add_964827;
  wire [7:0] sel_964828;
  wire [7:0] add_964831;
  wire [7:0] sel_964832;
  wire [7:0] add_964835;
  wire [7:0] sel_964836;
  wire [7:0] add_964839;
  wire [7:0] sel_964840;
  wire [7:0] add_964843;
  wire [7:0] sel_964844;
  wire [7:0] add_964847;
  wire [7:0] sel_964848;
  wire [7:0] add_964851;
  wire [7:0] sel_964852;
  wire [7:0] add_964855;
  wire [7:0] sel_964856;
  wire [7:0] add_964859;
  wire [7:0] sel_964860;
  wire [7:0] add_964863;
  wire [7:0] sel_964864;
  wire [7:0] add_964867;
  wire [7:0] sel_964868;
  wire [7:0] add_964871;
  wire [7:0] sel_964872;
  wire [7:0] add_964875;
  wire [7:0] sel_964876;
  wire [7:0] add_964879;
  wire [7:0] sel_964880;
  wire [7:0] add_964883;
  wire [7:0] sel_964884;
  wire [7:0] add_964887;
  wire [7:0] sel_964888;
  wire [7:0] add_964891;
  wire [7:0] sel_964892;
  wire [7:0] add_964895;
  wire [7:0] sel_964896;
  wire [7:0] add_964899;
  wire [7:0] sel_964900;
  wire [7:0] add_964903;
  wire [7:0] sel_964904;
  wire [7:0] add_964907;
  wire [7:0] sel_964908;
  wire [7:0] add_964911;
  wire [7:0] sel_964912;
  wire [7:0] add_964915;
  wire [7:0] sel_964916;
  wire [7:0] add_964919;
  wire [7:0] sel_964920;
  wire [7:0] add_964923;
  wire [7:0] sel_964924;
  wire [7:0] add_964927;
  wire [7:0] sel_964928;
  wire [7:0] add_964931;
  wire [7:0] sel_964932;
  wire [7:0] add_964935;
  wire [7:0] sel_964936;
  wire [7:0] add_964939;
  wire [7:0] sel_964940;
  wire [7:0] add_964943;
  wire [7:0] sel_964944;
  wire [7:0] add_964947;
  wire [7:0] sel_964948;
  wire [7:0] add_964951;
  wire [7:0] sel_964952;
  wire [7:0] add_964955;
  wire [7:0] sel_964956;
  wire [7:0] add_964959;
  wire [7:0] sel_964960;
  wire [7:0] add_964963;
  wire [7:0] sel_964964;
  wire [7:0] add_964967;
  wire [7:0] sel_964968;
  wire [7:0] add_964971;
  wire [7:0] sel_964972;
  wire [7:0] add_964975;
  wire [7:0] sel_964976;
  wire [7:0] add_964979;
  wire [7:0] sel_964980;
  wire [7:0] add_964983;
  wire [7:0] sel_964984;
  wire [7:0] add_964987;
  wire [7:0] sel_964988;
  wire [7:0] add_964991;
  wire [7:0] sel_964992;
  wire [7:0] add_964995;
  wire [7:0] sel_964996;
  wire [7:0] add_964999;
  wire [7:0] sel_965000;
  wire [7:0] add_965003;
  wire [7:0] sel_965004;
  wire [7:0] add_965007;
  wire [7:0] sel_965008;
  wire [7:0] add_965011;
  wire [7:0] sel_965012;
  wire [7:0] add_965015;
  wire [7:0] sel_965016;
  wire [7:0] add_965019;
  wire [7:0] sel_965020;
  wire [7:0] add_965023;
  wire [7:0] sel_965024;
  wire [7:0] add_965027;
  wire [7:0] sel_965028;
  wire [7:0] add_965031;
  wire [7:0] sel_965032;
  wire [7:0] add_965035;
  wire [7:0] sel_965036;
  wire [7:0] add_965039;
  wire [7:0] sel_965040;
  wire [7:0] add_965043;
  wire [7:0] sel_965044;
  wire [7:0] add_965047;
  wire [7:0] sel_965048;
  wire [7:0] add_965051;
  wire [7:0] sel_965052;
  wire [7:0] add_965055;
  wire [7:0] sel_965056;
  wire [7:0] add_965059;
  wire [7:0] sel_965060;
  wire [7:0] add_965063;
  wire [7:0] sel_965064;
  wire [7:0] add_965067;
  wire [7:0] sel_965068;
  wire [7:0] add_965071;
  wire [7:0] sel_965072;
  wire [7:0] add_965075;
  wire [7:0] sel_965076;
  wire [7:0] add_965079;
  wire [7:0] sel_965080;
  wire [7:0] add_965083;
  wire [7:0] sel_965084;
  wire [7:0] add_965087;
  wire [7:0] sel_965088;
  wire [7:0] add_965091;
  wire [7:0] sel_965092;
  wire [7:0] add_965095;
  wire [7:0] sel_965096;
  wire [7:0] add_965099;
  wire [7:0] sel_965100;
  wire [7:0] add_965103;
  wire [7:0] sel_965104;
  wire [7:0] add_965107;
  wire [7:0] sel_965108;
  wire [7:0] add_965111;
  wire [7:0] sel_965112;
  wire [7:0] add_965115;
  wire [7:0] sel_965116;
  wire [7:0] add_965119;
  wire [7:0] sel_965120;
  wire [7:0] add_965123;
  wire [7:0] sel_965124;
  wire [7:0] add_965127;
  wire [7:0] sel_965128;
  wire [7:0] add_965131;
  wire [7:0] sel_965132;
  wire [7:0] add_965135;
  wire [7:0] sel_965136;
  wire [7:0] add_965139;
  wire [7:0] sel_965140;
  wire [7:0] add_965143;
  wire [7:0] sel_965144;
  wire [7:0] add_965147;
  wire [7:0] sel_965148;
  wire [7:0] add_965151;
  wire [7:0] sel_965152;
  wire [7:0] add_965155;
  wire [7:0] sel_965156;
  wire [7:0] add_965159;
  wire [7:0] sel_965160;
  wire [7:0] add_965163;
  wire [7:0] sel_965164;
  wire [7:0] add_965167;
  wire [7:0] sel_965168;
  wire [7:0] add_965172;
  wire [15:0] array_index_965173;
  wire [7:0] sel_965174;
  wire [7:0] add_965177;
  wire [7:0] sel_965178;
  wire [7:0] add_965181;
  wire [7:0] sel_965182;
  wire [7:0] add_965185;
  wire [7:0] sel_965186;
  wire [7:0] add_965189;
  wire [7:0] sel_965190;
  wire [7:0] add_965193;
  wire [7:0] sel_965194;
  wire [7:0] add_965197;
  wire [7:0] sel_965198;
  wire [7:0] add_965201;
  wire [7:0] sel_965202;
  wire [7:0] add_965205;
  wire [7:0] sel_965206;
  wire [7:0] add_965209;
  wire [7:0] sel_965210;
  wire [7:0] add_965213;
  wire [7:0] sel_965214;
  wire [7:0] add_965217;
  wire [7:0] sel_965218;
  wire [7:0] add_965221;
  wire [7:0] sel_965222;
  wire [7:0] add_965225;
  wire [7:0] sel_965226;
  wire [7:0] add_965229;
  wire [7:0] sel_965230;
  wire [7:0] add_965233;
  wire [7:0] sel_965234;
  wire [7:0] add_965237;
  wire [7:0] sel_965238;
  wire [7:0] add_965241;
  wire [7:0] sel_965242;
  wire [7:0] add_965245;
  wire [7:0] sel_965246;
  wire [7:0] add_965249;
  wire [7:0] sel_965250;
  wire [7:0] add_965253;
  wire [7:0] sel_965254;
  wire [7:0] add_965257;
  wire [7:0] sel_965258;
  wire [7:0] add_965261;
  wire [7:0] sel_965262;
  wire [7:0] add_965265;
  wire [7:0] sel_965266;
  wire [7:0] add_965269;
  wire [7:0] sel_965270;
  wire [7:0] add_965273;
  wire [7:0] sel_965274;
  wire [7:0] add_965277;
  wire [7:0] sel_965278;
  wire [7:0] add_965281;
  wire [7:0] sel_965282;
  wire [7:0] add_965285;
  wire [7:0] sel_965286;
  wire [7:0] add_965289;
  wire [7:0] sel_965290;
  wire [7:0] add_965293;
  wire [7:0] sel_965294;
  wire [7:0] add_965297;
  wire [7:0] sel_965298;
  wire [7:0] add_965301;
  wire [7:0] sel_965302;
  wire [7:0] add_965305;
  wire [7:0] sel_965306;
  wire [7:0] add_965309;
  wire [7:0] sel_965310;
  wire [7:0] add_965313;
  wire [7:0] sel_965314;
  wire [7:0] add_965317;
  wire [7:0] sel_965318;
  wire [7:0] add_965321;
  wire [7:0] sel_965322;
  wire [7:0] add_965325;
  wire [7:0] sel_965326;
  wire [7:0] add_965329;
  wire [7:0] sel_965330;
  wire [7:0] add_965333;
  wire [7:0] sel_965334;
  wire [7:0] add_965337;
  wire [7:0] sel_965338;
  wire [7:0] add_965341;
  wire [7:0] sel_965342;
  wire [7:0] add_965345;
  wire [7:0] sel_965346;
  wire [7:0] add_965349;
  wire [7:0] sel_965350;
  wire [7:0] add_965353;
  wire [7:0] sel_965354;
  wire [7:0] add_965357;
  wire [7:0] sel_965358;
  wire [7:0] add_965361;
  wire [7:0] sel_965362;
  wire [7:0] add_965365;
  wire [7:0] sel_965366;
  wire [7:0] add_965369;
  wire [7:0] sel_965370;
  wire [7:0] add_965373;
  wire [7:0] sel_965374;
  wire [7:0] add_965377;
  wire [7:0] sel_965378;
  wire [7:0] add_965381;
  wire [7:0] sel_965382;
  wire [7:0] add_965385;
  wire [7:0] sel_965386;
  wire [7:0] add_965389;
  wire [7:0] sel_965390;
  wire [7:0] add_965393;
  wire [7:0] sel_965394;
  wire [7:0] add_965397;
  wire [7:0] sel_965398;
  wire [7:0] add_965401;
  wire [7:0] sel_965402;
  wire [7:0] add_965405;
  wire [7:0] sel_965406;
  wire [7:0] add_965409;
  wire [7:0] sel_965410;
  wire [7:0] add_965413;
  wire [7:0] sel_965414;
  wire [7:0] add_965417;
  wire [7:0] sel_965418;
  wire [7:0] add_965421;
  wire [7:0] sel_965422;
  wire [7:0] add_965425;
  wire [7:0] sel_965426;
  wire [7:0] add_965429;
  wire [7:0] sel_965430;
  wire [7:0] add_965433;
  wire [7:0] sel_965434;
  wire [7:0] add_965437;
  wire [7:0] sel_965438;
  wire [7:0] add_965441;
  wire [7:0] sel_965442;
  wire [7:0] add_965445;
  wire [7:0] sel_965446;
  wire [7:0] add_965449;
  wire [7:0] sel_965450;
  wire [7:0] add_965453;
  wire [7:0] sel_965454;
  wire [7:0] add_965457;
  wire [7:0] sel_965458;
  wire [7:0] add_965461;
  wire [7:0] sel_965462;
  wire [7:0] add_965465;
  wire [7:0] sel_965466;
  wire [7:0] add_965469;
  wire [7:0] sel_965470;
  wire [7:0] add_965473;
  wire [7:0] sel_965474;
  wire [7:0] add_965477;
  wire [7:0] sel_965478;
  wire [7:0] add_965481;
  wire [7:0] sel_965482;
  wire [7:0] add_965485;
  wire [7:0] sel_965486;
  wire [7:0] add_965489;
  wire [7:0] sel_965490;
  wire [7:0] add_965493;
  wire [7:0] sel_965494;
  wire [7:0] add_965497;
  wire [7:0] sel_965498;
  wire [7:0] add_965501;
  wire [7:0] sel_965502;
  wire [7:0] add_965505;
  wire [7:0] sel_965506;
  wire [7:0] add_965509;
  wire [7:0] sel_965510;
  wire [7:0] add_965513;
  wire [7:0] sel_965514;
  wire [7:0] add_965517;
  wire [7:0] sel_965518;
  wire [7:0] add_965521;
  wire [7:0] sel_965522;
  wire [7:0] add_965525;
  wire [7:0] sel_965526;
  wire [7:0] add_965529;
  wire [7:0] sel_965530;
  wire [7:0] add_965533;
  wire [7:0] sel_965534;
  wire [7:0] add_965537;
  wire [7:0] sel_965538;
  wire [7:0] add_965541;
  wire [7:0] sel_965542;
  wire [7:0] add_965545;
  wire [7:0] sel_965546;
  wire [7:0] add_965549;
  wire [7:0] sel_965550;
  wire [7:0] add_965553;
  wire [7:0] sel_965554;
  wire [7:0] add_965557;
  wire [7:0] sel_965558;
  wire [7:0] add_965561;
  wire [7:0] sel_965562;
  wire [7:0] add_965565;
  wire [7:0] sel_965566;
  wire [7:0] add_965569;
  wire [7:0] sel_965570;
  wire [7:0] add_965574;
  wire [15:0] array_index_965575;
  wire [7:0] sel_965576;
  wire [7:0] add_965579;
  wire [7:0] sel_965580;
  wire [7:0] add_965583;
  wire [7:0] sel_965584;
  wire [7:0] add_965587;
  wire [7:0] sel_965588;
  wire [7:0] add_965591;
  wire [7:0] sel_965592;
  wire [7:0] add_965595;
  wire [7:0] sel_965596;
  wire [7:0] add_965599;
  wire [7:0] sel_965600;
  wire [7:0] add_965603;
  wire [7:0] sel_965604;
  wire [7:0] add_965607;
  wire [7:0] sel_965608;
  wire [7:0] add_965611;
  wire [7:0] sel_965612;
  wire [7:0] add_965615;
  wire [7:0] sel_965616;
  wire [7:0] add_965619;
  wire [7:0] sel_965620;
  wire [7:0] add_965623;
  wire [7:0] sel_965624;
  wire [7:0] add_965627;
  wire [7:0] sel_965628;
  wire [7:0] add_965631;
  wire [7:0] sel_965632;
  wire [7:0] add_965635;
  wire [7:0] sel_965636;
  wire [7:0] add_965639;
  wire [7:0] sel_965640;
  wire [7:0] add_965643;
  wire [7:0] sel_965644;
  wire [7:0] add_965647;
  wire [7:0] sel_965648;
  wire [7:0] add_965651;
  wire [7:0] sel_965652;
  wire [7:0] add_965655;
  wire [7:0] sel_965656;
  wire [7:0] add_965659;
  wire [7:0] sel_965660;
  wire [7:0] add_965663;
  wire [7:0] sel_965664;
  wire [7:0] add_965667;
  wire [7:0] sel_965668;
  wire [7:0] add_965671;
  wire [7:0] sel_965672;
  wire [7:0] add_965675;
  wire [7:0] sel_965676;
  wire [7:0] add_965679;
  wire [7:0] sel_965680;
  wire [7:0] add_965683;
  wire [7:0] sel_965684;
  wire [7:0] add_965687;
  wire [7:0] sel_965688;
  wire [7:0] add_965691;
  wire [7:0] sel_965692;
  wire [7:0] add_965695;
  wire [7:0] sel_965696;
  wire [7:0] add_965699;
  wire [7:0] sel_965700;
  wire [7:0] add_965703;
  wire [7:0] sel_965704;
  wire [7:0] add_965707;
  wire [7:0] sel_965708;
  wire [7:0] add_965711;
  wire [7:0] sel_965712;
  wire [7:0] add_965715;
  wire [7:0] sel_965716;
  wire [7:0] add_965719;
  wire [7:0] sel_965720;
  wire [7:0] add_965723;
  wire [7:0] sel_965724;
  wire [7:0] add_965727;
  wire [7:0] sel_965728;
  wire [7:0] add_965731;
  wire [7:0] sel_965732;
  wire [7:0] add_965735;
  wire [7:0] sel_965736;
  wire [7:0] add_965739;
  wire [7:0] sel_965740;
  wire [7:0] add_965743;
  wire [7:0] sel_965744;
  wire [7:0] add_965747;
  wire [7:0] sel_965748;
  wire [7:0] add_965751;
  wire [7:0] sel_965752;
  wire [7:0] add_965755;
  wire [7:0] sel_965756;
  wire [7:0] add_965759;
  wire [7:0] sel_965760;
  wire [7:0] add_965763;
  wire [7:0] sel_965764;
  wire [7:0] add_965767;
  wire [7:0] sel_965768;
  wire [7:0] add_965771;
  wire [7:0] sel_965772;
  wire [7:0] add_965775;
  wire [7:0] sel_965776;
  wire [7:0] add_965779;
  wire [7:0] sel_965780;
  wire [7:0] add_965783;
  wire [7:0] sel_965784;
  wire [7:0] add_965787;
  wire [7:0] sel_965788;
  wire [7:0] add_965791;
  wire [7:0] sel_965792;
  wire [7:0] add_965795;
  wire [7:0] sel_965796;
  wire [7:0] add_965799;
  wire [7:0] sel_965800;
  wire [7:0] add_965803;
  wire [7:0] sel_965804;
  wire [7:0] add_965807;
  wire [7:0] sel_965808;
  wire [7:0] add_965811;
  wire [7:0] sel_965812;
  wire [7:0] add_965815;
  wire [7:0] sel_965816;
  wire [7:0] add_965819;
  wire [7:0] sel_965820;
  wire [7:0] add_965823;
  wire [7:0] sel_965824;
  wire [7:0] add_965827;
  wire [7:0] sel_965828;
  wire [7:0] add_965831;
  wire [7:0] sel_965832;
  wire [7:0] add_965835;
  wire [7:0] sel_965836;
  wire [7:0] add_965839;
  wire [7:0] sel_965840;
  wire [7:0] add_965843;
  wire [7:0] sel_965844;
  wire [7:0] add_965847;
  wire [7:0] sel_965848;
  wire [7:0] add_965851;
  wire [7:0] sel_965852;
  wire [7:0] add_965855;
  wire [7:0] sel_965856;
  wire [7:0] add_965859;
  wire [7:0] sel_965860;
  wire [7:0] add_965863;
  wire [7:0] sel_965864;
  wire [7:0] add_965867;
  wire [7:0] sel_965868;
  wire [7:0] add_965871;
  wire [7:0] sel_965872;
  wire [7:0] add_965875;
  wire [7:0] sel_965876;
  wire [7:0] add_965879;
  wire [7:0] sel_965880;
  wire [7:0] add_965883;
  wire [7:0] sel_965884;
  wire [7:0] add_965887;
  wire [7:0] sel_965888;
  wire [7:0] add_965891;
  wire [7:0] sel_965892;
  wire [7:0] add_965895;
  wire [7:0] sel_965896;
  wire [7:0] add_965899;
  wire [7:0] sel_965900;
  wire [7:0] add_965903;
  wire [7:0] sel_965904;
  wire [7:0] add_965907;
  wire [7:0] sel_965908;
  wire [7:0] add_965911;
  wire [7:0] sel_965912;
  wire [7:0] add_965915;
  wire [7:0] sel_965916;
  wire [7:0] add_965919;
  wire [7:0] sel_965920;
  wire [7:0] add_965923;
  wire [7:0] sel_965924;
  wire [7:0] add_965927;
  wire [7:0] sel_965928;
  wire [7:0] add_965931;
  wire [7:0] sel_965932;
  wire [7:0] add_965935;
  wire [7:0] sel_965936;
  wire [7:0] add_965939;
  wire [7:0] sel_965940;
  wire [7:0] add_965943;
  wire [7:0] sel_965944;
  wire [7:0] add_965947;
  wire [7:0] sel_965948;
  wire [7:0] add_965951;
  wire [7:0] sel_965952;
  wire [7:0] add_965955;
  wire [7:0] sel_965956;
  wire [7:0] add_965959;
  wire [7:0] sel_965960;
  wire [7:0] add_965963;
  wire [7:0] sel_965964;
  wire [7:0] add_965967;
  wire [7:0] sel_965968;
  wire [7:0] add_965971;
  wire [7:0] sel_965972;
  wire [7:0] add_965976;
  wire [15:0] array_index_965977;
  wire [7:0] sel_965978;
  wire [7:0] add_965981;
  wire [7:0] sel_965982;
  wire [7:0] add_965985;
  wire [7:0] sel_965986;
  wire [7:0] add_965989;
  wire [7:0] sel_965990;
  wire [7:0] add_965993;
  wire [7:0] sel_965994;
  wire [7:0] add_965997;
  wire [7:0] sel_965998;
  wire [7:0] add_966001;
  wire [7:0] sel_966002;
  wire [7:0] add_966005;
  wire [7:0] sel_966006;
  wire [7:0] add_966009;
  wire [7:0] sel_966010;
  wire [7:0] add_966013;
  wire [7:0] sel_966014;
  wire [7:0] add_966017;
  wire [7:0] sel_966018;
  wire [7:0] add_966021;
  wire [7:0] sel_966022;
  wire [7:0] add_966025;
  wire [7:0] sel_966026;
  wire [7:0] add_966029;
  wire [7:0] sel_966030;
  wire [7:0] add_966033;
  wire [7:0] sel_966034;
  wire [7:0] add_966037;
  wire [7:0] sel_966038;
  wire [7:0] add_966041;
  wire [7:0] sel_966042;
  wire [7:0] add_966045;
  wire [7:0] sel_966046;
  wire [7:0] add_966049;
  wire [7:0] sel_966050;
  wire [7:0] add_966053;
  wire [7:0] sel_966054;
  wire [7:0] add_966057;
  wire [7:0] sel_966058;
  wire [7:0] add_966061;
  wire [7:0] sel_966062;
  wire [7:0] add_966065;
  wire [7:0] sel_966066;
  wire [7:0] add_966069;
  wire [7:0] sel_966070;
  wire [7:0] add_966073;
  wire [7:0] sel_966074;
  wire [7:0] add_966077;
  wire [7:0] sel_966078;
  wire [7:0] add_966081;
  wire [7:0] sel_966082;
  wire [7:0] add_966085;
  wire [7:0] sel_966086;
  wire [7:0] add_966089;
  wire [7:0] sel_966090;
  wire [7:0] add_966093;
  wire [7:0] sel_966094;
  wire [7:0] add_966097;
  wire [7:0] sel_966098;
  wire [7:0] add_966101;
  wire [7:0] sel_966102;
  wire [7:0] add_966105;
  wire [7:0] sel_966106;
  wire [7:0] add_966109;
  wire [7:0] sel_966110;
  wire [7:0] add_966113;
  wire [7:0] sel_966114;
  wire [7:0] add_966117;
  wire [7:0] sel_966118;
  wire [7:0] add_966121;
  wire [7:0] sel_966122;
  wire [7:0] add_966125;
  wire [7:0] sel_966126;
  wire [7:0] add_966129;
  wire [7:0] sel_966130;
  wire [7:0] add_966133;
  wire [7:0] sel_966134;
  wire [7:0] add_966137;
  wire [7:0] sel_966138;
  wire [7:0] add_966141;
  wire [7:0] sel_966142;
  wire [7:0] add_966145;
  wire [7:0] sel_966146;
  wire [7:0] add_966149;
  wire [7:0] sel_966150;
  wire [7:0] add_966153;
  wire [7:0] sel_966154;
  wire [7:0] add_966157;
  wire [7:0] sel_966158;
  wire [7:0] add_966161;
  wire [7:0] sel_966162;
  wire [7:0] add_966165;
  wire [7:0] sel_966166;
  wire [7:0] add_966169;
  wire [7:0] sel_966170;
  wire [7:0] add_966173;
  wire [7:0] sel_966174;
  wire [7:0] add_966177;
  wire [7:0] sel_966178;
  wire [7:0] add_966181;
  wire [7:0] sel_966182;
  wire [7:0] add_966185;
  wire [7:0] sel_966186;
  wire [7:0] add_966189;
  wire [7:0] sel_966190;
  wire [7:0] add_966193;
  wire [7:0] sel_966194;
  wire [7:0] add_966197;
  wire [7:0] sel_966198;
  wire [7:0] add_966201;
  wire [7:0] sel_966202;
  wire [7:0] add_966205;
  wire [7:0] sel_966206;
  wire [7:0] add_966209;
  wire [7:0] sel_966210;
  wire [7:0] add_966213;
  wire [7:0] sel_966214;
  wire [7:0] add_966217;
  wire [7:0] sel_966218;
  wire [7:0] add_966221;
  wire [7:0] sel_966222;
  wire [7:0] add_966225;
  wire [7:0] sel_966226;
  wire [7:0] add_966229;
  wire [7:0] sel_966230;
  wire [7:0] add_966233;
  wire [7:0] sel_966234;
  wire [7:0] add_966237;
  wire [7:0] sel_966238;
  wire [7:0] add_966241;
  wire [7:0] sel_966242;
  wire [7:0] add_966245;
  wire [7:0] sel_966246;
  wire [7:0] add_966249;
  wire [7:0] sel_966250;
  wire [7:0] add_966253;
  wire [7:0] sel_966254;
  wire [7:0] add_966257;
  wire [7:0] sel_966258;
  wire [7:0] add_966261;
  wire [7:0] sel_966262;
  wire [7:0] add_966265;
  wire [7:0] sel_966266;
  wire [7:0] add_966269;
  wire [7:0] sel_966270;
  wire [7:0] add_966273;
  wire [7:0] sel_966274;
  wire [7:0] add_966277;
  wire [7:0] sel_966278;
  wire [7:0] add_966281;
  wire [7:0] sel_966282;
  wire [7:0] add_966285;
  wire [7:0] sel_966286;
  wire [7:0] add_966289;
  wire [7:0] sel_966290;
  wire [7:0] add_966293;
  wire [7:0] sel_966294;
  wire [7:0] add_966297;
  wire [7:0] sel_966298;
  wire [7:0] add_966301;
  wire [7:0] sel_966302;
  wire [7:0] add_966305;
  wire [7:0] sel_966306;
  wire [7:0] add_966309;
  wire [7:0] sel_966310;
  wire [7:0] add_966313;
  wire [7:0] sel_966314;
  wire [7:0] add_966317;
  wire [7:0] sel_966318;
  wire [7:0] add_966321;
  wire [7:0] sel_966322;
  wire [7:0] add_966325;
  wire [7:0] sel_966326;
  wire [7:0] add_966329;
  wire [7:0] sel_966330;
  wire [7:0] add_966333;
  wire [7:0] sel_966334;
  wire [7:0] add_966337;
  wire [7:0] sel_966338;
  wire [7:0] add_966341;
  wire [7:0] sel_966342;
  wire [7:0] add_966345;
  wire [7:0] sel_966346;
  wire [7:0] add_966349;
  wire [7:0] sel_966350;
  wire [7:0] add_966353;
  wire [7:0] sel_966354;
  wire [7:0] add_966357;
  wire [7:0] sel_966358;
  wire [7:0] add_966361;
  wire [7:0] sel_966362;
  wire [7:0] add_966365;
  wire [7:0] sel_966366;
  wire [7:0] add_966369;
  wire [7:0] sel_966370;
  wire [7:0] add_966373;
  wire [7:0] sel_966374;
  wire [7:0] add_966378;
  wire [15:0] array_index_966379;
  wire [7:0] sel_966380;
  wire [7:0] add_966383;
  wire [7:0] sel_966384;
  wire [7:0] add_966387;
  wire [7:0] sel_966388;
  wire [7:0] add_966391;
  wire [7:0] sel_966392;
  wire [7:0] add_966395;
  wire [7:0] sel_966396;
  wire [7:0] add_966399;
  wire [7:0] sel_966400;
  wire [7:0] add_966403;
  wire [7:0] sel_966404;
  wire [7:0] add_966407;
  wire [7:0] sel_966408;
  wire [7:0] add_966411;
  wire [7:0] sel_966412;
  wire [7:0] add_966415;
  wire [7:0] sel_966416;
  wire [7:0] add_966419;
  wire [7:0] sel_966420;
  wire [7:0] add_966423;
  wire [7:0] sel_966424;
  wire [7:0] add_966427;
  wire [7:0] sel_966428;
  wire [7:0] add_966431;
  wire [7:0] sel_966432;
  wire [7:0] add_966435;
  wire [7:0] sel_966436;
  wire [7:0] add_966439;
  wire [7:0] sel_966440;
  wire [7:0] add_966443;
  wire [7:0] sel_966444;
  wire [7:0] add_966447;
  wire [7:0] sel_966448;
  wire [7:0] add_966451;
  wire [7:0] sel_966452;
  wire [7:0] add_966455;
  wire [7:0] sel_966456;
  wire [7:0] add_966459;
  wire [7:0] sel_966460;
  wire [7:0] add_966463;
  wire [7:0] sel_966464;
  wire [7:0] add_966467;
  wire [7:0] sel_966468;
  wire [7:0] add_966471;
  wire [7:0] sel_966472;
  wire [7:0] add_966475;
  wire [7:0] sel_966476;
  wire [7:0] add_966479;
  wire [7:0] sel_966480;
  wire [7:0] add_966483;
  wire [7:0] sel_966484;
  wire [7:0] add_966487;
  wire [7:0] sel_966488;
  wire [7:0] add_966491;
  wire [7:0] sel_966492;
  wire [7:0] add_966495;
  wire [7:0] sel_966496;
  wire [7:0] add_966499;
  wire [7:0] sel_966500;
  wire [7:0] add_966503;
  wire [7:0] sel_966504;
  wire [7:0] add_966507;
  wire [7:0] sel_966508;
  wire [7:0] add_966511;
  wire [7:0] sel_966512;
  wire [7:0] add_966515;
  wire [7:0] sel_966516;
  wire [7:0] add_966519;
  wire [7:0] sel_966520;
  wire [7:0] add_966523;
  wire [7:0] sel_966524;
  wire [7:0] add_966527;
  wire [7:0] sel_966528;
  wire [7:0] add_966531;
  wire [7:0] sel_966532;
  wire [7:0] add_966535;
  wire [7:0] sel_966536;
  wire [7:0] add_966539;
  wire [7:0] sel_966540;
  wire [7:0] add_966543;
  wire [7:0] sel_966544;
  wire [7:0] add_966547;
  wire [7:0] sel_966548;
  wire [7:0] add_966551;
  wire [7:0] sel_966552;
  wire [7:0] add_966555;
  wire [7:0] sel_966556;
  wire [7:0] add_966559;
  wire [7:0] sel_966560;
  wire [7:0] add_966563;
  wire [7:0] sel_966564;
  wire [7:0] add_966567;
  wire [7:0] sel_966568;
  wire [7:0] add_966571;
  wire [7:0] sel_966572;
  wire [7:0] add_966575;
  wire [7:0] sel_966576;
  wire [7:0] add_966579;
  wire [7:0] sel_966580;
  wire [7:0] add_966583;
  wire [7:0] sel_966584;
  wire [7:0] add_966587;
  wire [7:0] sel_966588;
  wire [7:0] add_966591;
  wire [7:0] sel_966592;
  wire [7:0] add_966595;
  wire [7:0] sel_966596;
  wire [7:0] add_966599;
  wire [7:0] sel_966600;
  wire [7:0] add_966603;
  wire [7:0] sel_966604;
  wire [7:0] add_966607;
  wire [7:0] sel_966608;
  wire [7:0] add_966611;
  wire [7:0] sel_966612;
  wire [7:0] add_966615;
  wire [7:0] sel_966616;
  wire [7:0] add_966619;
  wire [7:0] sel_966620;
  wire [7:0] add_966623;
  wire [7:0] sel_966624;
  wire [7:0] add_966627;
  wire [7:0] sel_966628;
  wire [7:0] add_966631;
  wire [7:0] sel_966632;
  wire [7:0] add_966635;
  wire [7:0] sel_966636;
  wire [7:0] add_966639;
  wire [7:0] sel_966640;
  wire [7:0] add_966643;
  wire [7:0] sel_966644;
  wire [7:0] add_966647;
  wire [7:0] sel_966648;
  wire [7:0] add_966651;
  wire [7:0] sel_966652;
  wire [7:0] add_966655;
  wire [7:0] sel_966656;
  wire [7:0] add_966659;
  wire [7:0] sel_966660;
  wire [7:0] add_966663;
  wire [7:0] sel_966664;
  wire [7:0] add_966667;
  wire [7:0] sel_966668;
  wire [7:0] add_966671;
  wire [7:0] sel_966672;
  wire [7:0] add_966675;
  wire [7:0] sel_966676;
  wire [7:0] add_966679;
  wire [7:0] sel_966680;
  wire [7:0] add_966683;
  wire [7:0] sel_966684;
  wire [7:0] add_966687;
  wire [7:0] sel_966688;
  wire [7:0] add_966691;
  wire [7:0] sel_966692;
  wire [7:0] add_966695;
  wire [7:0] sel_966696;
  wire [7:0] add_966699;
  wire [7:0] sel_966700;
  wire [7:0] add_966703;
  wire [7:0] sel_966704;
  wire [7:0] add_966707;
  wire [7:0] sel_966708;
  wire [7:0] add_966711;
  wire [7:0] sel_966712;
  wire [7:0] add_966715;
  wire [7:0] sel_966716;
  wire [7:0] add_966719;
  wire [7:0] sel_966720;
  wire [7:0] add_966723;
  wire [7:0] sel_966724;
  wire [7:0] add_966727;
  wire [7:0] sel_966728;
  wire [7:0] add_966731;
  wire [7:0] sel_966732;
  wire [7:0] add_966735;
  wire [7:0] sel_966736;
  wire [7:0] add_966739;
  wire [7:0] sel_966740;
  wire [7:0] add_966743;
  wire [7:0] sel_966744;
  wire [7:0] add_966747;
  wire [7:0] sel_966748;
  wire [7:0] add_966751;
  wire [7:0] sel_966752;
  wire [7:0] add_966755;
  wire [7:0] sel_966756;
  wire [7:0] add_966759;
  wire [7:0] sel_966760;
  wire [7:0] add_966763;
  wire [7:0] sel_966764;
  wire [7:0] add_966767;
  wire [7:0] sel_966768;
  wire [7:0] add_966771;
  wire [7:0] sel_966772;
  wire [7:0] add_966775;
  wire [7:0] sel_966776;
  wire [7:0] add_966780;
  wire [15:0] array_index_966781;
  wire [7:0] sel_966782;
  wire [7:0] add_966785;
  wire [7:0] sel_966786;
  wire [7:0] add_966789;
  wire [7:0] sel_966790;
  wire [7:0] add_966793;
  wire [7:0] sel_966794;
  wire [7:0] add_966797;
  wire [7:0] sel_966798;
  wire [7:0] add_966801;
  wire [7:0] sel_966802;
  wire [7:0] add_966805;
  wire [7:0] sel_966806;
  wire [7:0] add_966809;
  wire [7:0] sel_966810;
  wire [7:0] add_966813;
  wire [7:0] sel_966814;
  wire [7:0] add_966817;
  wire [7:0] sel_966818;
  wire [7:0] add_966821;
  wire [7:0] sel_966822;
  wire [7:0] add_966825;
  wire [7:0] sel_966826;
  wire [7:0] add_966829;
  wire [7:0] sel_966830;
  wire [7:0] add_966833;
  wire [7:0] sel_966834;
  wire [7:0] add_966837;
  wire [7:0] sel_966838;
  wire [7:0] add_966841;
  wire [7:0] sel_966842;
  wire [7:0] add_966845;
  wire [7:0] sel_966846;
  wire [7:0] add_966849;
  wire [7:0] sel_966850;
  wire [7:0] add_966853;
  wire [7:0] sel_966854;
  wire [7:0] add_966857;
  wire [7:0] sel_966858;
  wire [7:0] add_966861;
  wire [7:0] sel_966862;
  wire [7:0] add_966865;
  wire [7:0] sel_966866;
  wire [7:0] add_966869;
  wire [7:0] sel_966870;
  wire [7:0] add_966873;
  wire [7:0] sel_966874;
  wire [7:0] add_966877;
  wire [7:0] sel_966878;
  wire [7:0] add_966881;
  wire [7:0] sel_966882;
  wire [7:0] add_966885;
  wire [7:0] sel_966886;
  wire [7:0] add_966889;
  wire [7:0] sel_966890;
  wire [7:0] add_966893;
  wire [7:0] sel_966894;
  wire [7:0] add_966897;
  wire [7:0] sel_966898;
  wire [7:0] add_966901;
  wire [7:0] sel_966902;
  wire [7:0] add_966905;
  wire [7:0] sel_966906;
  wire [7:0] add_966909;
  wire [7:0] sel_966910;
  wire [7:0] add_966913;
  wire [7:0] sel_966914;
  wire [7:0] add_966917;
  wire [7:0] sel_966918;
  wire [7:0] add_966921;
  wire [7:0] sel_966922;
  wire [7:0] add_966925;
  wire [7:0] sel_966926;
  wire [7:0] add_966929;
  wire [7:0] sel_966930;
  wire [7:0] add_966933;
  wire [7:0] sel_966934;
  wire [7:0] add_966937;
  wire [7:0] sel_966938;
  wire [7:0] add_966941;
  wire [7:0] sel_966942;
  wire [7:0] add_966945;
  wire [7:0] sel_966946;
  wire [7:0] add_966949;
  wire [7:0] sel_966950;
  wire [7:0] add_966953;
  wire [7:0] sel_966954;
  wire [7:0] add_966957;
  wire [7:0] sel_966958;
  wire [7:0] add_966961;
  wire [7:0] sel_966962;
  wire [7:0] add_966965;
  wire [7:0] sel_966966;
  wire [7:0] add_966969;
  wire [7:0] sel_966970;
  wire [7:0] add_966973;
  wire [7:0] sel_966974;
  wire [7:0] add_966977;
  wire [7:0] sel_966978;
  wire [7:0] add_966981;
  wire [7:0] sel_966982;
  wire [7:0] add_966985;
  wire [7:0] sel_966986;
  wire [7:0] add_966989;
  wire [7:0] sel_966990;
  wire [7:0] add_966993;
  wire [7:0] sel_966994;
  wire [7:0] add_966997;
  wire [7:0] sel_966998;
  wire [7:0] add_967001;
  wire [7:0] sel_967002;
  wire [7:0] add_967005;
  wire [7:0] sel_967006;
  wire [7:0] add_967009;
  wire [7:0] sel_967010;
  wire [7:0] add_967013;
  wire [7:0] sel_967014;
  wire [7:0] add_967017;
  wire [7:0] sel_967018;
  wire [7:0] add_967021;
  wire [7:0] sel_967022;
  wire [7:0] add_967025;
  wire [7:0] sel_967026;
  wire [7:0] add_967029;
  wire [7:0] sel_967030;
  wire [7:0] add_967033;
  wire [7:0] sel_967034;
  wire [7:0] add_967037;
  wire [7:0] sel_967038;
  wire [7:0] add_967041;
  wire [7:0] sel_967042;
  wire [7:0] add_967045;
  wire [7:0] sel_967046;
  wire [7:0] add_967049;
  wire [7:0] sel_967050;
  wire [7:0] add_967053;
  wire [7:0] sel_967054;
  wire [7:0] add_967057;
  wire [7:0] sel_967058;
  wire [7:0] add_967061;
  wire [7:0] sel_967062;
  wire [7:0] add_967065;
  wire [7:0] sel_967066;
  wire [7:0] add_967069;
  wire [7:0] sel_967070;
  wire [7:0] add_967073;
  wire [7:0] sel_967074;
  wire [7:0] add_967077;
  wire [7:0] sel_967078;
  wire [7:0] add_967081;
  wire [7:0] sel_967082;
  wire [7:0] add_967085;
  wire [7:0] sel_967086;
  wire [7:0] add_967089;
  wire [7:0] sel_967090;
  wire [7:0] add_967093;
  wire [7:0] sel_967094;
  wire [7:0] add_967097;
  wire [7:0] sel_967098;
  wire [7:0] add_967101;
  wire [7:0] sel_967102;
  wire [7:0] add_967105;
  wire [7:0] sel_967106;
  wire [7:0] add_967109;
  wire [7:0] sel_967110;
  wire [7:0] add_967113;
  wire [7:0] sel_967114;
  wire [7:0] add_967117;
  wire [7:0] sel_967118;
  wire [7:0] add_967121;
  wire [7:0] sel_967122;
  wire [7:0] add_967125;
  wire [7:0] sel_967126;
  wire [7:0] add_967129;
  wire [7:0] sel_967130;
  wire [7:0] add_967133;
  wire [7:0] sel_967134;
  wire [7:0] add_967137;
  wire [7:0] sel_967138;
  wire [7:0] add_967141;
  wire [7:0] sel_967142;
  wire [7:0] add_967145;
  wire [7:0] sel_967146;
  wire [7:0] add_967149;
  wire [7:0] sel_967150;
  wire [7:0] add_967153;
  wire [7:0] sel_967154;
  wire [7:0] add_967157;
  wire [7:0] sel_967158;
  wire [7:0] add_967161;
  wire [7:0] sel_967162;
  wire [7:0] add_967165;
  wire [7:0] sel_967166;
  wire [7:0] add_967169;
  wire [7:0] sel_967170;
  wire [7:0] add_967173;
  wire [7:0] sel_967174;
  wire [7:0] add_967177;
  wire [7:0] sel_967178;
  wire [7:0] add_967182;
  wire [15:0] array_index_967183;
  wire [7:0] sel_967184;
  wire [7:0] add_967187;
  wire [7:0] sel_967188;
  wire [7:0] add_967191;
  wire [7:0] sel_967192;
  wire [7:0] add_967195;
  wire [7:0] sel_967196;
  wire [7:0] add_967199;
  wire [7:0] sel_967200;
  wire [7:0] add_967203;
  wire [7:0] sel_967204;
  wire [7:0] add_967207;
  wire [7:0] sel_967208;
  wire [7:0] add_967211;
  wire [7:0] sel_967212;
  wire [7:0] add_967215;
  wire [7:0] sel_967216;
  wire [7:0] add_967219;
  wire [7:0] sel_967220;
  wire [7:0] add_967223;
  wire [7:0] sel_967224;
  wire [7:0] add_967227;
  wire [7:0] sel_967228;
  wire [7:0] add_967231;
  wire [7:0] sel_967232;
  wire [7:0] add_967235;
  wire [7:0] sel_967236;
  wire [7:0] add_967239;
  wire [7:0] sel_967240;
  wire [7:0] add_967243;
  wire [7:0] sel_967244;
  wire [7:0] add_967247;
  wire [7:0] sel_967248;
  wire [7:0] add_967251;
  wire [7:0] sel_967252;
  wire [7:0] add_967255;
  wire [7:0] sel_967256;
  wire [7:0] add_967259;
  wire [7:0] sel_967260;
  wire [7:0] add_967263;
  wire [7:0] sel_967264;
  wire [7:0] add_967267;
  wire [7:0] sel_967268;
  wire [7:0] add_967271;
  wire [7:0] sel_967272;
  wire [7:0] add_967275;
  wire [7:0] sel_967276;
  wire [7:0] add_967279;
  wire [7:0] sel_967280;
  wire [7:0] add_967283;
  wire [7:0] sel_967284;
  wire [7:0] add_967287;
  wire [7:0] sel_967288;
  wire [7:0] add_967291;
  wire [7:0] sel_967292;
  wire [7:0] add_967295;
  wire [7:0] sel_967296;
  wire [7:0] add_967299;
  wire [7:0] sel_967300;
  wire [7:0] add_967303;
  wire [7:0] sel_967304;
  wire [7:0] add_967307;
  wire [7:0] sel_967308;
  wire [7:0] add_967311;
  wire [7:0] sel_967312;
  wire [7:0] add_967315;
  wire [7:0] sel_967316;
  wire [7:0] add_967319;
  wire [7:0] sel_967320;
  wire [7:0] add_967323;
  wire [7:0] sel_967324;
  wire [7:0] add_967327;
  wire [7:0] sel_967328;
  wire [7:0] add_967331;
  wire [7:0] sel_967332;
  wire [7:0] add_967335;
  wire [7:0] sel_967336;
  wire [7:0] add_967339;
  wire [7:0] sel_967340;
  wire [7:0] add_967343;
  wire [7:0] sel_967344;
  wire [7:0] add_967347;
  wire [7:0] sel_967348;
  wire [7:0] add_967351;
  wire [7:0] sel_967352;
  wire [7:0] add_967355;
  wire [7:0] sel_967356;
  wire [7:0] add_967359;
  wire [7:0] sel_967360;
  wire [7:0] add_967363;
  wire [7:0] sel_967364;
  wire [7:0] add_967367;
  wire [7:0] sel_967368;
  wire [7:0] add_967371;
  wire [7:0] sel_967372;
  wire [7:0] add_967375;
  wire [7:0] sel_967376;
  wire [7:0] add_967379;
  wire [7:0] sel_967380;
  wire [7:0] add_967383;
  wire [7:0] sel_967384;
  wire [7:0] add_967387;
  wire [7:0] sel_967388;
  wire [7:0] add_967391;
  wire [7:0] sel_967392;
  wire [7:0] add_967395;
  wire [7:0] sel_967396;
  wire [7:0] add_967399;
  wire [7:0] sel_967400;
  wire [7:0] add_967403;
  wire [7:0] sel_967404;
  wire [7:0] add_967407;
  wire [7:0] sel_967408;
  wire [7:0] add_967411;
  wire [7:0] sel_967412;
  wire [7:0] add_967415;
  wire [7:0] sel_967416;
  wire [7:0] add_967419;
  wire [7:0] sel_967420;
  wire [7:0] add_967423;
  wire [7:0] sel_967424;
  wire [7:0] add_967427;
  wire [7:0] sel_967428;
  wire [7:0] add_967431;
  wire [7:0] sel_967432;
  wire [7:0] add_967435;
  wire [7:0] sel_967436;
  wire [7:0] add_967439;
  wire [7:0] sel_967440;
  wire [7:0] add_967443;
  wire [7:0] sel_967444;
  wire [7:0] add_967447;
  wire [7:0] sel_967448;
  wire [7:0] add_967451;
  wire [7:0] sel_967452;
  wire [7:0] add_967455;
  wire [7:0] sel_967456;
  wire [7:0] add_967459;
  wire [7:0] sel_967460;
  wire [7:0] add_967463;
  wire [7:0] sel_967464;
  wire [7:0] add_967467;
  wire [7:0] sel_967468;
  wire [7:0] add_967471;
  wire [7:0] sel_967472;
  wire [7:0] add_967475;
  wire [7:0] sel_967476;
  wire [7:0] add_967479;
  wire [7:0] sel_967480;
  wire [7:0] add_967483;
  wire [7:0] sel_967484;
  wire [7:0] add_967487;
  wire [7:0] sel_967488;
  wire [7:0] add_967491;
  wire [7:0] sel_967492;
  wire [7:0] add_967495;
  wire [7:0] sel_967496;
  wire [7:0] add_967499;
  wire [7:0] sel_967500;
  wire [7:0] add_967503;
  wire [7:0] sel_967504;
  wire [7:0] add_967507;
  wire [7:0] sel_967508;
  wire [7:0] add_967511;
  wire [7:0] sel_967512;
  wire [7:0] add_967515;
  wire [7:0] sel_967516;
  wire [7:0] add_967519;
  wire [7:0] sel_967520;
  wire [7:0] add_967523;
  wire [7:0] sel_967524;
  wire [7:0] add_967527;
  wire [7:0] sel_967528;
  wire [7:0] add_967531;
  wire [7:0] sel_967532;
  wire [7:0] add_967535;
  wire [7:0] sel_967536;
  wire [7:0] add_967539;
  wire [7:0] sel_967540;
  wire [7:0] add_967543;
  wire [7:0] sel_967544;
  wire [7:0] add_967547;
  wire [7:0] sel_967548;
  wire [7:0] add_967551;
  wire [7:0] sel_967552;
  wire [7:0] add_967555;
  wire [7:0] sel_967556;
  wire [7:0] add_967559;
  wire [7:0] sel_967560;
  wire [7:0] add_967563;
  wire [7:0] sel_967564;
  wire [7:0] add_967567;
  wire [7:0] sel_967568;
  wire [7:0] add_967571;
  wire [7:0] sel_967572;
  wire [7:0] add_967575;
  wire [7:0] sel_967576;
  wire [7:0] add_967579;
  wire [7:0] sel_967580;
  wire [7:0] add_967584;
  wire [15:0] array_index_967585;
  wire [7:0] sel_967586;
  wire [7:0] add_967589;
  wire [7:0] sel_967590;
  wire [7:0] add_967593;
  wire [7:0] sel_967594;
  wire [7:0] add_967597;
  wire [7:0] sel_967598;
  wire [7:0] add_967601;
  wire [7:0] sel_967602;
  wire [7:0] add_967605;
  wire [7:0] sel_967606;
  wire [7:0] add_967609;
  wire [7:0] sel_967610;
  wire [7:0] add_967613;
  wire [7:0] sel_967614;
  wire [7:0] add_967617;
  wire [7:0] sel_967618;
  wire [7:0] add_967621;
  wire [7:0] sel_967622;
  wire [7:0] add_967625;
  wire [7:0] sel_967626;
  wire [7:0] add_967629;
  wire [7:0] sel_967630;
  wire [7:0] add_967633;
  wire [7:0] sel_967634;
  wire [7:0] add_967637;
  wire [7:0] sel_967638;
  wire [7:0] add_967641;
  wire [7:0] sel_967642;
  wire [7:0] add_967645;
  wire [7:0] sel_967646;
  wire [7:0] add_967649;
  wire [7:0] sel_967650;
  wire [7:0] add_967653;
  wire [7:0] sel_967654;
  wire [7:0] add_967657;
  wire [7:0] sel_967658;
  wire [7:0] add_967661;
  wire [7:0] sel_967662;
  wire [7:0] add_967665;
  wire [7:0] sel_967666;
  wire [7:0] add_967669;
  wire [7:0] sel_967670;
  wire [7:0] add_967673;
  wire [7:0] sel_967674;
  wire [7:0] add_967677;
  wire [7:0] sel_967678;
  wire [7:0] add_967681;
  wire [7:0] sel_967682;
  wire [7:0] add_967685;
  wire [7:0] sel_967686;
  wire [7:0] add_967689;
  wire [7:0] sel_967690;
  wire [7:0] add_967693;
  wire [7:0] sel_967694;
  wire [7:0] add_967697;
  wire [7:0] sel_967698;
  wire [7:0] add_967701;
  wire [7:0] sel_967702;
  wire [7:0] add_967705;
  wire [7:0] sel_967706;
  wire [7:0] add_967709;
  wire [7:0] sel_967710;
  wire [7:0] add_967713;
  wire [7:0] sel_967714;
  wire [7:0] add_967717;
  wire [7:0] sel_967718;
  wire [7:0] add_967721;
  wire [7:0] sel_967722;
  wire [7:0] add_967725;
  wire [7:0] sel_967726;
  wire [7:0] add_967729;
  wire [7:0] sel_967730;
  wire [7:0] add_967733;
  wire [7:0] sel_967734;
  wire [7:0] add_967737;
  wire [7:0] sel_967738;
  wire [7:0] add_967741;
  wire [7:0] sel_967742;
  wire [7:0] add_967745;
  wire [7:0] sel_967746;
  wire [7:0] add_967749;
  wire [7:0] sel_967750;
  wire [7:0] add_967753;
  wire [7:0] sel_967754;
  wire [7:0] add_967757;
  wire [7:0] sel_967758;
  wire [7:0] add_967761;
  wire [7:0] sel_967762;
  wire [7:0] add_967765;
  wire [7:0] sel_967766;
  wire [7:0] add_967769;
  wire [7:0] sel_967770;
  wire [7:0] add_967773;
  wire [7:0] sel_967774;
  wire [7:0] add_967777;
  wire [7:0] sel_967778;
  wire [7:0] add_967781;
  wire [7:0] sel_967782;
  wire [7:0] add_967785;
  wire [7:0] sel_967786;
  wire [7:0] add_967789;
  wire [7:0] sel_967790;
  wire [7:0] add_967793;
  wire [7:0] sel_967794;
  wire [7:0] add_967797;
  wire [7:0] sel_967798;
  wire [7:0] add_967801;
  wire [7:0] sel_967802;
  wire [7:0] add_967805;
  wire [7:0] sel_967806;
  wire [7:0] add_967809;
  wire [7:0] sel_967810;
  wire [7:0] add_967813;
  wire [7:0] sel_967814;
  wire [7:0] add_967817;
  wire [7:0] sel_967818;
  wire [7:0] add_967821;
  wire [7:0] sel_967822;
  wire [7:0] add_967825;
  wire [7:0] sel_967826;
  wire [7:0] add_967829;
  wire [7:0] sel_967830;
  wire [7:0] add_967833;
  wire [7:0] sel_967834;
  wire [7:0] add_967837;
  wire [7:0] sel_967838;
  wire [7:0] add_967841;
  wire [7:0] sel_967842;
  wire [7:0] add_967845;
  wire [7:0] sel_967846;
  wire [7:0] add_967849;
  wire [7:0] sel_967850;
  wire [7:0] add_967853;
  wire [7:0] sel_967854;
  wire [7:0] add_967857;
  wire [7:0] sel_967858;
  wire [7:0] add_967861;
  wire [7:0] sel_967862;
  wire [7:0] add_967865;
  wire [7:0] sel_967866;
  wire [7:0] add_967869;
  wire [7:0] sel_967870;
  wire [7:0] add_967873;
  wire [7:0] sel_967874;
  wire [7:0] add_967877;
  wire [7:0] sel_967878;
  wire [7:0] add_967881;
  wire [7:0] sel_967882;
  wire [7:0] add_967885;
  wire [7:0] sel_967886;
  wire [7:0] add_967889;
  wire [7:0] sel_967890;
  wire [7:0] add_967893;
  wire [7:0] sel_967894;
  wire [7:0] add_967897;
  wire [7:0] sel_967898;
  wire [7:0] add_967901;
  wire [7:0] sel_967902;
  wire [7:0] add_967905;
  wire [7:0] sel_967906;
  wire [7:0] add_967909;
  wire [7:0] sel_967910;
  wire [7:0] add_967913;
  wire [7:0] sel_967914;
  wire [7:0] add_967917;
  wire [7:0] sel_967918;
  wire [7:0] add_967921;
  wire [7:0] sel_967922;
  wire [7:0] add_967925;
  wire [7:0] sel_967926;
  wire [7:0] add_967929;
  wire [7:0] sel_967930;
  wire [7:0] add_967933;
  wire [7:0] sel_967934;
  wire [7:0] add_967937;
  wire [7:0] sel_967938;
  wire [7:0] add_967941;
  wire [7:0] sel_967942;
  wire [7:0] add_967945;
  wire [7:0] sel_967946;
  wire [7:0] add_967949;
  wire [7:0] sel_967950;
  wire [7:0] add_967953;
  wire [7:0] sel_967954;
  wire [7:0] add_967957;
  wire [7:0] sel_967958;
  wire [7:0] add_967961;
  wire [7:0] sel_967962;
  wire [7:0] add_967965;
  wire [7:0] sel_967966;
  wire [7:0] add_967969;
  wire [7:0] sel_967970;
  wire [7:0] add_967973;
  wire [7:0] sel_967974;
  wire [7:0] add_967977;
  wire [7:0] sel_967978;
  wire [7:0] add_967981;
  wire [7:0] sel_967982;
  wire [7:0] add_967986;
  wire [15:0] array_index_967987;
  wire [7:0] sel_967988;
  wire [7:0] add_967991;
  wire [7:0] sel_967992;
  wire [7:0] add_967995;
  wire [7:0] sel_967996;
  wire [7:0] add_967999;
  wire [7:0] sel_968000;
  wire [7:0] add_968003;
  wire [7:0] sel_968004;
  wire [7:0] add_968007;
  wire [7:0] sel_968008;
  wire [7:0] add_968011;
  wire [7:0] sel_968012;
  wire [7:0] add_968015;
  wire [7:0] sel_968016;
  wire [7:0] add_968019;
  wire [7:0] sel_968020;
  wire [7:0] add_968023;
  wire [7:0] sel_968024;
  wire [7:0] add_968027;
  wire [7:0] sel_968028;
  wire [7:0] add_968031;
  wire [7:0] sel_968032;
  wire [7:0] add_968035;
  wire [7:0] sel_968036;
  wire [7:0] add_968039;
  wire [7:0] sel_968040;
  wire [7:0] add_968043;
  wire [7:0] sel_968044;
  wire [7:0] add_968047;
  wire [7:0] sel_968048;
  wire [7:0] add_968051;
  wire [7:0] sel_968052;
  wire [7:0] add_968055;
  wire [7:0] sel_968056;
  wire [7:0] add_968059;
  wire [7:0] sel_968060;
  wire [7:0] add_968063;
  wire [7:0] sel_968064;
  wire [7:0] add_968067;
  wire [7:0] sel_968068;
  wire [7:0] add_968071;
  wire [7:0] sel_968072;
  wire [7:0] add_968075;
  wire [7:0] sel_968076;
  wire [7:0] add_968079;
  wire [7:0] sel_968080;
  wire [7:0] add_968083;
  wire [7:0] sel_968084;
  wire [7:0] add_968087;
  wire [7:0] sel_968088;
  wire [7:0] add_968091;
  wire [7:0] sel_968092;
  wire [7:0] add_968095;
  wire [7:0] sel_968096;
  wire [7:0] add_968099;
  wire [7:0] sel_968100;
  wire [7:0] add_968103;
  wire [7:0] sel_968104;
  wire [7:0] add_968107;
  wire [7:0] sel_968108;
  wire [7:0] add_968111;
  wire [7:0] sel_968112;
  wire [7:0] add_968115;
  wire [7:0] sel_968116;
  wire [7:0] add_968119;
  wire [7:0] sel_968120;
  wire [7:0] add_968123;
  wire [7:0] sel_968124;
  wire [7:0] add_968127;
  wire [7:0] sel_968128;
  wire [7:0] add_968131;
  wire [7:0] sel_968132;
  wire [7:0] add_968135;
  wire [7:0] sel_968136;
  wire [7:0] add_968139;
  wire [7:0] sel_968140;
  wire [7:0] add_968143;
  wire [7:0] sel_968144;
  wire [7:0] add_968147;
  wire [7:0] sel_968148;
  wire [7:0] add_968151;
  wire [7:0] sel_968152;
  wire [7:0] add_968155;
  wire [7:0] sel_968156;
  wire [7:0] add_968159;
  wire [7:0] sel_968160;
  wire [7:0] add_968163;
  wire [7:0] sel_968164;
  wire [7:0] add_968167;
  wire [7:0] sel_968168;
  wire [7:0] add_968171;
  wire [7:0] sel_968172;
  wire [7:0] add_968175;
  wire [7:0] sel_968176;
  wire [7:0] add_968179;
  wire [7:0] sel_968180;
  wire [7:0] add_968183;
  wire [7:0] sel_968184;
  wire [7:0] add_968187;
  wire [7:0] sel_968188;
  wire [7:0] add_968191;
  wire [7:0] sel_968192;
  wire [7:0] add_968195;
  wire [7:0] sel_968196;
  wire [7:0] add_968199;
  wire [7:0] sel_968200;
  wire [7:0] add_968203;
  wire [7:0] sel_968204;
  wire [7:0] add_968207;
  wire [7:0] sel_968208;
  wire [7:0] add_968211;
  wire [7:0] sel_968212;
  wire [7:0] add_968215;
  wire [7:0] sel_968216;
  wire [7:0] add_968219;
  wire [7:0] sel_968220;
  wire [7:0] add_968223;
  wire [7:0] sel_968224;
  wire [7:0] add_968227;
  wire [7:0] sel_968228;
  wire [7:0] add_968231;
  wire [7:0] sel_968232;
  wire [7:0] add_968235;
  wire [7:0] sel_968236;
  wire [7:0] add_968239;
  wire [7:0] sel_968240;
  wire [7:0] add_968243;
  wire [7:0] sel_968244;
  wire [7:0] add_968247;
  wire [7:0] sel_968248;
  wire [7:0] add_968251;
  wire [7:0] sel_968252;
  wire [7:0] add_968255;
  wire [7:0] sel_968256;
  wire [7:0] add_968259;
  wire [7:0] sel_968260;
  wire [7:0] add_968263;
  wire [7:0] sel_968264;
  wire [7:0] add_968267;
  wire [7:0] sel_968268;
  wire [7:0] add_968271;
  wire [7:0] sel_968272;
  wire [7:0] add_968275;
  wire [7:0] sel_968276;
  wire [7:0] add_968279;
  wire [7:0] sel_968280;
  wire [7:0] add_968283;
  wire [7:0] sel_968284;
  wire [7:0] add_968287;
  wire [7:0] sel_968288;
  wire [7:0] add_968291;
  wire [7:0] sel_968292;
  wire [7:0] add_968295;
  wire [7:0] sel_968296;
  wire [7:0] add_968299;
  wire [7:0] sel_968300;
  wire [7:0] add_968303;
  wire [7:0] sel_968304;
  wire [7:0] add_968307;
  wire [7:0] sel_968308;
  wire [7:0] add_968311;
  wire [7:0] sel_968312;
  wire [7:0] add_968315;
  wire [7:0] sel_968316;
  wire [7:0] add_968319;
  wire [7:0] sel_968320;
  wire [7:0] add_968323;
  wire [7:0] sel_968324;
  wire [7:0] add_968327;
  wire [7:0] sel_968328;
  wire [7:0] add_968331;
  wire [7:0] sel_968332;
  wire [7:0] add_968335;
  wire [7:0] sel_968336;
  wire [7:0] add_968339;
  wire [7:0] sel_968340;
  wire [7:0] add_968343;
  wire [7:0] sel_968344;
  wire [7:0] add_968347;
  wire [7:0] sel_968348;
  wire [7:0] add_968351;
  wire [7:0] sel_968352;
  wire [7:0] add_968355;
  wire [7:0] sel_968356;
  wire [7:0] add_968359;
  wire [7:0] sel_968360;
  wire [7:0] add_968363;
  wire [7:0] sel_968364;
  wire [7:0] add_968367;
  wire [7:0] sel_968368;
  wire [7:0] add_968371;
  wire [7:0] sel_968372;
  wire [7:0] add_968375;
  wire [7:0] sel_968376;
  wire [7:0] add_968379;
  wire [7:0] sel_968380;
  wire [7:0] add_968383;
  wire [7:0] sel_968384;
  wire [7:0] add_968388;
  wire [15:0] array_index_968389;
  wire [7:0] sel_968390;
  wire [7:0] add_968393;
  wire [7:0] sel_968394;
  wire [7:0] add_968397;
  wire [7:0] sel_968398;
  wire [7:0] add_968401;
  wire [7:0] sel_968402;
  wire [7:0] add_968405;
  wire [7:0] sel_968406;
  wire [7:0] add_968409;
  wire [7:0] sel_968410;
  wire [7:0] add_968413;
  wire [7:0] sel_968414;
  wire [7:0] add_968417;
  wire [7:0] sel_968418;
  wire [7:0] add_968421;
  wire [7:0] sel_968422;
  wire [7:0] add_968425;
  wire [7:0] sel_968426;
  wire [7:0] add_968429;
  wire [7:0] sel_968430;
  wire [7:0] add_968433;
  wire [7:0] sel_968434;
  wire [7:0] add_968437;
  wire [7:0] sel_968438;
  wire [7:0] add_968441;
  wire [7:0] sel_968442;
  wire [7:0] add_968445;
  wire [7:0] sel_968446;
  wire [7:0] add_968449;
  wire [7:0] sel_968450;
  wire [7:0] add_968453;
  wire [7:0] sel_968454;
  wire [7:0] add_968457;
  wire [7:0] sel_968458;
  wire [7:0] add_968461;
  wire [7:0] sel_968462;
  wire [7:0] add_968465;
  wire [7:0] sel_968466;
  wire [7:0] add_968469;
  wire [7:0] sel_968470;
  wire [7:0] add_968473;
  wire [7:0] sel_968474;
  wire [7:0] add_968477;
  wire [7:0] sel_968478;
  wire [7:0] add_968481;
  wire [7:0] sel_968482;
  wire [7:0] add_968485;
  wire [7:0] sel_968486;
  wire [7:0] add_968489;
  wire [7:0] sel_968490;
  wire [7:0] add_968493;
  wire [7:0] sel_968494;
  wire [7:0] add_968497;
  wire [7:0] sel_968498;
  wire [7:0] add_968501;
  wire [7:0] sel_968502;
  wire [7:0] add_968505;
  wire [7:0] sel_968506;
  wire [7:0] add_968509;
  wire [7:0] sel_968510;
  wire [7:0] add_968513;
  wire [7:0] sel_968514;
  wire [7:0] add_968517;
  wire [7:0] sel_968518;
  wire [7:0] add_968521;
  wire [7:0] sel_968522;
  wire [7:0] add_968525;
  wire [7:0] sel_968526;
  wire [7:0] add_968529;
  wire [7:0] sel_968530;
  wire [7:0] add_968533;
  wire [7:0] sel_968534;
  wire [7:0] add_968537;
  wire [7:0] sel_968538;
  wire [7:0] add_968541;
  wire [7:0] sel_968542;
  wire [7:0] add_968545;
  wire [7:0] sel_968546;
  wire [7:0] add_968549;
  wire [7:0] sel_968550;
  wire [7:0] add_968553;
  wire [7:0] sel_968554;
  wire [7:0] add_968557;
  wire [7:0] sel_968558;
  wire [7:0] add_968561;
  wire [7:0] sel_968562;
  wire [7:0] add_968565;
  wire [7:0] sel_968566;
  wire [7:0] add_968569;
  wire [7:0] sel_968570;
  wire [7:0] add_968573;
  wire [7:0] sel_968574;
  wire [7:0] add_968577;
  wire [7:0] sel_968578;
  wire [7:0] add_968581;
  wire [7:0] sel_968582;
  wire [7:0] add_968585;
  wire [7:0] sel_968586;
  wire [7:0] add_968589;
  wire [7:0] sel_968590;
  wire [7:0] add_968593;
  wire [7:0] sel_968594;
  wire [7:0] add_968597;
  wire [7:0] sel_968598;
  wire [7:0] add_968601;
  wire [7:0] sel_968602;
  wire [7:0] add_968605;
  wire [7:0] sel_968606;
  wire [7:0] add_968609;
  wire [7:0] sel_968610;
  wire [7:0] add_968613;
  wire [7:0] sel_968614;
  wire [7:0] add_968617;
  wire [7:0] sel_968618;
  wire [7:0] add_968621;
  wire [7:0] sel_968622;
  wire [7:0] add_968625;
  wire [7:0] sel_968626;
  wire [7:0] add_968629;
  wire [7:0] sel_968630;
  wire [7:0] add_968633;
  wire [7:0] sel_968634;
  wire [7:0] add_968637;
  wire [7:0] sel_968638;
  wire [7:0] add_968641;
  wire [7:0] sel_968642;
  wire [7:0] add_968645;
  wire [7:0] sel_968646;
  wire [7:0] add_968649;
  wire [7:0] sel_968650;
  wire [7:0] add_968653;
  wire [7:0] sel_968654;
  wire [7:0] add_968657;
  wire [7:0] sel_968658;
  wire [7:0] add_968661;
  wire [7:0] sel_968662;
  wire [7:0] add_968665;
  wire [7:0] sel_968666;
  wire [7:0] add_968669;
  wire [7:0] sel_968670;
  wire [7:0] add_968673;
  wire [7:0] sel_968674;
  wire [7:0] add_968677;
  wire [7:0] sel_968678;
  wire [7:0] add_968681;
  wire [7:0] sel_968682;
  wire [7:0] add_968685;
  wire [7:0] sel_968686;
  wire [7:0] add_968689;
  wire [7:0] sel_968690;
  wire [7:0] add_968693;
  wire [7:0] sel_968694;
  wire [7:0] add_968697;
  wire [7:0] sel_968698;
  wire [7:0] add_968701;
  wire [7:0] sel_968702;
  wire [7:0] add_968705;
  wire [7:0] sel_968706;
  wire [7:0] add_968709;
  wire [7:0] sel_968710;
  wire [7:0] add_968713;
  wire [7:0] sel_968714;
  wire [7:0] add_968717;
  wire [7:0] sel_968718;
  wire [7:0] add_968721;
  wire [7:0] sel_968722;
  wire [7:0] add_968725;
  wire [7:0] sel_968726;
  wire [7:0] add_968729;
  wire [7:0] sel_968730;
  wire [7:0] add_968733;
  wire [7:0] sel_968734;
  wire [7:0] add_968737;
  wire [7:0] sel_968738;
  wire [7:0] add_968741;
  wire [7:0] sel_968742;
  wire [7:0] add_968745;
  wire [7:0] sel_968746;
  wire [7:0] add_968749;
  wire [7:0] sel_968750;
  wire [7:0] add_968753;
  wire [7:0] sel_968754;
  wire [7:0] add_968757;
  wire [7:0] sel_968758;
  wire [7:0] add_968761;
  wire [7:0] sel_968762;
  wire [7:0] add_968765;
  wire [7:0] sel_968766;
  wire [7:0] add_968769;
  wire [7:0] sel_968770;
  wire [7:0] add_968773;
  wire [7:0] sel_968774;
  wire [7:0] add_968777;
  wire [7:0] sel_968778;
  wire [7:0] add_968781;
  wire [7:0] sel_968782;
  wire [7:0] add_968785;
  wire [7:0] sel_968786;
  wire [7:0] add_968790;
  wire [15:0] array_index_968791;
  wire [7:0] sel_968792;
  wire [7:0] add_968795;
  wire [7:0] sel_968796;
  wire [7:0] add_968799;
  wire [7:0] sel_968800;
  wire [7:0] add_968803;
  wire [7:0] sel_968804;
  wire [7:0] add_968807;
  wire [7:0] sel_968808;
  wire [7:0] add_968811;
  wire [7:0] sel_968812;
  wire [7:0] add_968815;
  wire [7:0] sel_968816;
  wire [7:0] add_968819;
  wire [7:0] sel_968820;
  wire [7:0] add_968823;
  wire [7:0] sel_968824;
  wire [7:0] add_968827;
  wire [7:0] sel_968828;
  wire [7:0] add_968831;
  wire [7:0] sel_968832;
  wire [7:0] add_968835;
  wire [7:0] sel_968836;
  wire [7:0] add_968839;
  wire [7:0] sel_968840;
  wire [7:0] add_968843;
  wire [7:0] sel_968844;
  wire [7:0] add_968847;
  wire [7:0] sel_968848;
  wire [7:0] add_968851;
  wire [7:0] sel_968852;
  wire [7:0] add_968855;
  wire [7:0] sel_968856;
  wire [7:0] add_968859;
  wire [7:0] sel_968860;
  wire [7:0] add_968863;
  wire [7:0] sel_968864;
  wire [7:0] add_968867;
  wire [7:0] sel_968868;
  wire [7:0] add_968871;
  wire [7:0] sel_968872;
  wire [7:0] add_968875;
  wire [7:0] sel_968876;
  wire [7:0] add_968879;
  wire [7:0] sel_968880;
  wire [7:0] add_968883;
  wire [7:0] sel_968884;
  wire [7:0] add_968887;
  wire [7:0] sel_968888;
  wire [7:0] add_968891;
  wire [7:0] sel_968892;
  wire [7:0] add_968895;
  wire [7:0] sel_968896;
  wire [7:0] add_968899;
  wire [7:0] sel_968900;
  wire [7:0] add_968903;
  wire [7:0] sel_968904;
  wire [7:0] add_968907;
  wire [7:0] sel_968908;
  wire [7:0] add_968911;
  wire [7:0] sel_968912;
  wire [7:0] add_968915;
  wire [7:0] sel_968916;
  wire [7:0] add_968919;
  wire [7:0] sel_968920;
  wire [7:0] add_968923;
  wire [7:0] sel_968924;
  wire [7:0] add_968927;
  wire [7:0] sel_968928;
  wire [7:0] add_968931;
  wire [7:0] sel_968932;
  wire [7:0] add_968935;
  wire [7:0] sel_968936;
  wire [7:0] add_968939;
  wire [7:0] sel_968940;
  wire [7:0] add_968943;
  wire [7:0] sel_968944;
  wire [7:0] add_968947;
  wire [7:0] sel_968948;
  wire [7:0] add_968951;
  wire [7:0] sel_968952;
  wire [7:0] add_968955;
  wire [7:0] sel_968956;
  wire [7:0] add_968959;
  wire [7:0] sel_968960;
  wire [7:0] add_968963;
  wire [7:0] sel_968964;
  wire [7:0] add_968967;
  wire [7:0] sel_968968;
  wire [7:0] add_968971;
  wire [7:0] sel_968972;
  wire [7:0] add_968975;
  wire [7:0] sel_968976;
  wire [7:0] add_968979;
  wire [7:0] sel_968980;
  wire [7:0] add_968983;
  wire [7:0] sel_968984;
  wire [7:0] add_968987;
  wire [7:0] sel_968988;
  wire [7:0] add_968991;
  wire [7:0] sel_968992;
  wire [7:0] add_968995;
  wire [7:0] sel_968996;
  wire [7:0] add_968999;
  wire [7:0] sel_969000;
  wire [7:0] add_969003;
  wire [7:0] sel_969004;
  wire [7:0] add_969007;
  wire [7:0] sel_969008;
  wire [7:0] add_969011;
  wire [7:0] sel_969012;
  wire [7:0] add_969015;
  wire [7:0] sel_969016;
  wire [7:0] add_969019;
  wire [7:0] sel_969020;
  wire [7:0] add_969023;
  wire [7:0] sel_969024;
  wire [7:0] add_969027;
  wire [7:0] sel_969028;
  wire [7:0] add_969031;
  wire [7:0] sel_969032;
  wire [7:0] add_969035;
  wire [7:0] sel_969036;
  wire [7:0] add_969039;
  wire [7:0] sel_969040;
  wire [7:0] add_969043;
  wire [7:0] sel_969044;
  wire [7:0] add_969047;
  wire [7:0] sel_969048;
  wire [7:0] add_969051;
  wire [7:0] sel_969052;
  wire [7:0] add_969055;
  wire [7:0] sel_969056;
  wire [7:0] add_969059;
  wire [7:0] sel_969060;
  wire [7:0] add_969063;
  wire [7:0] sel_969064;
  wire [7:0] add_969067;
  wire [7:0] sel_969068;
  wire [7:0] add_969071;
  wire [7:0] sel_969072;
  wire [7:0] add_969075;
  wire [7:0] sel_969076;
  wire [7:0] add_969079;
  wire [7:0] sel_969080;
  wire [7:0] add_969083;
  wire [7:0] sel_969084;
  wire [7:0] add_969087;
  wire [7:0] sel_969088;
  wire [7:0] add_969091;
  wire [7:0] sel_969092;
  wire [7:0] add_969095;
  wire [7:0] sel_969096;
  wire [7:0] add_969099;
  wire [7:0] sel_969100;
  wire [7:0] add_969103;
  wire [7:0] sel_969104;
  wire [7:0] add_969107;
  wire [7:0] sel_969108;
  wire [7:0] add_969111;
  wire [7:0] sel_969112;
  wire [7:0] add_969115;
  wire [7:0] sel_969116;
  wire [7:0] add_969119;
  wire [7:0] sel_969120;
  wire [7:0] add_969123;
  wire [7:0] sel_969124;
  wire [7:0] add_969127;
  wire [7:0] sel_969128;
  wire [7:0] add_969131;
  wire [7:0] sel_969132;
  wire [7:0] add_969135;
  wire [7:0] sel_969136;
  wire [7:0] add_969139;
  wire [7:0] sel_969140;
  wire [7:0] add_969143;
  wire [7:0] sel_969144;
  wire [7:0] add_969147;
  wire [7:0] sel_969148;
  wire [7:0] add_969151;
  wire [7:0] sel_969152;
  wire [7:0] add_969155;
  wire [7:0] sel_969156;
  wire [7:0] add_969159;
  wire [7:0] sel_969160;
  wire [7:0] add_969163;
  wire [7:0] sel_969164;
  wire [7:0] add_969167;
  wire [7:0] sel_969168;
  wire [7:0] add_969171;
  wire [7:0] sel_969172;
  wire [7:0] add_969175;
  wire [7:0] sel_969176;
  wire [7:0] add_969179;
  wire [7:0] sel_969180;
  wire [7:0] add_969183;
  wire [7:0] sel_969184;
  wire [7:0] add_969187;
  wire [7:0] sel_969188;
  wire [7:0] add_969192;
  wire [15:0] array_index_969193;
  wire [7:0] sel_969194;
  wire [7:0] add_969197;
  wire [7:0] sel_969198;
  wire [7:0] add_969201;
  wire [7:0] sel_969202;
  wire [7:0] add_969205;
  wire [7:0] sel_969206;
  wire [7:0] add_969209;
  wire [7:0] sel_969210;
  wire [7:0] add_969213;
  wire [7:0] sel_969214;
  wire [7:0] add_969217;
  wire [7:0] sel_969218;
  wire [7:0] add_969221;
  wire [7:0] sel_969222;
  wire [7:0] add_969225;
  wire [7:0] sel_969226;
  wire [7:0] add_969229;
  wire [7:0] sel_969230;
  wire [7:0] add_969233;
  wire [7:0] sel_969234;
  wire [7:0] add_969237;
  wire [7:0] sel_969238;
  wire [7:0] add_969241;
  wire [7:0] sel_969242;
  wire [7:0] add_969245;
  wire [7:0] sel_969246;
  wire [7:0] add_969249;
  wire [7:0] sel_969250;
  wire [7:0] add_969253;
  wire [7:0] sel_969254;
  wire [7:0] add_969257;
  wire [7:0] sel_969258;
  wire [7:0] add_969261;
  wire [7:0] sel_969262;
  wire [7:0] add_969265;
  wire [7:0] sel_969266;
  wire [7:0] add_969269;
  wire [7:0] sel_969270;
  wire [7:0] add_969273;
  wire [7:0] sel_969274;
  wire [7:0] add_969277;
  wire [7:0] sel_969278;
  wire [7:0] add_969281;
  wire [7:0] sel_969282;
  wire [7:0] add_969285;
  wire [7:0] sel_969286;
  wire [7:0] add_969289;
  wire [7:0] sel_969290;
  wire [7:0] add_969293;
  wire [7:0] sel_969294;
  wire [7:0] add_969297;
  wire [7:0] sel_969298;
  wire [7:0] add_969301;
  wire [7:0] sel_969302;
  wire [7:0] add_969305;
  wire [7:0] sel_969306;
  wire [7:0] add_969309;
  wire [7:0] sel_969310;
  wire [7:0] add_969313;
  wire [7:0] sel_969314;
  wire [7:0] add_969317;
  wire [7:0] sel_969318;
  wire [7:0] add_969321;
  wire [7:0] sel_969322;
  wire [7:0] add_969325;
  wire [7:0] sel_969326;
  wire [7:0] add_969329;
  wire [7:0] sel_969330;
  wire [7:0] add_969333;
  wire [7:0] sel_969334;
  wire [7:0] add_969337;
  wire [7:0] sel_969338;
  wire [7:0] add_969341;
  wire [7:0] sel_969342;
  wire [7:0] add_969345;
  wire [7:0] sel_969346;
  wire [7:0] add_969349;
  wire [7:0] sel_969350;
  wire [7:0] add_969353;
  wire [7:0] sel_969354;
  wire [7:0] add_969357;
  wire [7:0] sel_969358;
  wire [7:0] add_969361;
  wire [7:0] sel_969362;
  wire [7:0] add_969365;
  wire [7:0] sel_969366;
  wire [7:0] add_969369;
  wire [7:0] sel_969370;
  wire [7:0] add_969373;
  wire [7:0] sel_969374;
  wire [7:0] add_969377;
  wire [7:0] sel_969378;
  wire [7:0] add_969381;
  wire [7:0] sel_969382;
  wire [7:0] add_969385;
  wire [7:0] sel_969386;
  wire [7:0] add_969389;
  wire [7:0] sel_969390;
  wire [7:0] add_969393;
  wire [7:0] sel_969394;
  wire [7:0] add_969397;
  wire [7:0] sel_969398;
  wire [7:0] add_969401;
  wire [7:0] sel_969402;
  wire [7:0] add_969405;
  wire [7:0] sel_969406;
  wire [7:0] add_969409;
  wire [7:0] sel_969410;
  wire [7:0] add_969413;
  wire [7:0] sel_969414;
  wire [7:0] add_969417;
  wire [7:0] sel_969418;
  wire [7:0] add_969421;
  wire [7:0] sel_969422;
  wire [7:0] add_969425;
  wire [7:0] sel_969426;
  wire [7:0] add_969429;
  wire [7:0] sel_969430;
  wire [7:0] add_969433;
  wire [7:0] sel_969434;
  wire [7:0] add_969437;
  wire [7:0] sel_969438;
  wire [7:0] add_969441;
  wire [7:0] sel_969442;
  wire [7:0] add_969445;
  wire [7:0] sel_969446;
  wire [7:0] add_969449;
  wire [7:0] sel_969450;
  wire [7:0] add_969453;
  wire [7:0] sel_969454;
  wire [7:0] add_969457;
  wire [7:0] sel_969458;
  wire [7:0] add_969461;
  wire [7:0] sel_969462;
  wire [7:0] add_969465;
  wire [7:0] sel_969466;
  wire [7:0] add_969469;
  wire [7:0] sel_969470;
  wire [7:0] add_969473;
  wire [7:0] sel_969474;
  wire [7:0] add_969477;
  wire [7:0] sel_969478;
  wire [7:0] add_969481;
  wire [7:0] sel_969482;
  wire [7:0] add_969485;
  wire [7:0] sel_969486;
  wire [7:0] add_969489;
  wire [7:0] sel_969490;
  wire [7:0] add_969493;
  wire [7:0] sel_969494;
  wire [7:0] add_969497;
  wire [7:0] sel_969498;
  wire [7:0] add_969501;
  wire [7:0] sel_969502;
  wire [7:0] add_969505;
  wire [7:0] sel_969506;
  wire [7:0] add_969509;
  wire [7:0] sel_969510;
  wire [7:0] add_969513;
  wire [7:0] sel_969514;
  wire [7:0] add_969517;
  wire [7:0] sel_969518;
  wire [7:0] add_969521;
  wire [7:0] sel_969522;
  wire [7:0] add_969525;
  wire [7:0] sel_969526;
  wire [7:0] add_969529;
  wire [7:0] sel_969530;
  wire [7:0] add_969533;
  wire [7:0] sel_969534;
  wire [7:0] add_969537;
  wire [7:0] sel_969538;
  wire [7:0] add_969541;
  wire [7:0] sel_969542;
  wire [7:0] add_969545;
  wire [7:0] sel_969546;
  wire [7:0] add_969549;
  wire [7:0] sel_969550;
  wire [7:0] add_969553;
  wire [7:0] sel_969554;
  wire [7:0] add_969557;
  wire [7:0] sel_969558;
  wire [7:0] add_969561;
  wire [7:0] sel_969562;
  wire [7:0] add_969565;
  wire [7:0] sel_969566;
  wire [7:0] add_969569;
  wire [7:0] sel_969570;
  wire [7:0] add_969573;
  wire [7:0] sel_969574;
  wire [7:0] add_969577;
  wire [7:0] sel_969578;
  wire [7:0] add_969581;
  wire [7:0] sel_969582;
  wire [7:0] add_969585;
  wire [7:0] sel_969586;
  wire [7:0] add_969589;
  wire [7:0] sel_969590;
  wire [7:0] add_969594;
  wire [15:0] array_index_969595;
  wire [7:0] sel_969596;
  wire [7:0] add_969599;
  wire [7:0] sel_969600;
  wire [7:0] add_969603;
  wire [7:0] sel_969604;
  wire [7:0] add_969607;
  wire [7:0] sel_969608;
  wire [7:0] add_969611;
  wire [7:0] sel_969612;
  wire [7:0] add_969615;
  wire [7:0] sel_969616;
  wire [7:0] add_969619;
  wire [7:0] sel_969620;
  wire [7:0] add_969623;
  wire [7:0] sel_969624;
  wire [7:0] add_969627;
  wire [7:0] sel_969628;
  wire [7:0] add_969631;
  wire [7:0] sel_969632;
  wire [7:0] add_969635;
  wire [7:0] sel_969636;
  wire [7:0] add_969639;
  wire [7:0] sel_969640;
  wire [7:0] add_969643;
  wire [7:0] sel_969644;
  wire [7:0] add_969647;
  wire [7:0] sel_969648;
  wire [7:0] add_969651;
  wire [7:0] sel_969652;
  wire [7:0] add_969655;
  wire [7:0] sel_969656;
  wire [7:0] add_969659;
  wire [7:0] sel_969660;
  wire [7:0] add_969663;
  wire [7:0] sel_969664;
  wire [7:0] add_969667;
  wire [7:0] sel_969668;
  wire [7:0] add_969671;
  wire [7:0] sel_969672;
  wire [7:0] add_969675;
  wire [7:0] sel_969676;
  wire [7:0] add_969679;
  wire [7:0] sel_969680;
  wire [7:0] add_969683;
  wire [7:0] sel_969684;
  wire [7:0] add_969687;
  wire [7:0] sel_969688;
  wire [7:0] add_969691;
  wire [7:0] sel_969692;
  wire [7:0] add_969695;
  wire [7:0] sel_969696;
  wire [7:0] add_969699;
  wire [7:0] sel_969700;
  wire [7:0] add_969703;
  wire [7:0] sel_969704;
  wire [7:0] add_969707;
  wire [7:0] sel_969708;
  wire [7:0] add_969711;
  wire [7:0] sel_969712;
  wire [7:0] add_969715;
  wire [7:0] sel_969716;
  wire [7:0] add_969719;
  wire [7:0] sel_969720;
  wire [7:0] add_969723;
  wire [7:0] sel_969724;
  wire [7:0] add_969727;
  wire [7:0] sel_969728;
  wire [7:0] add_969731;
  wire [7:0] sel_969732;
  wire [7:0] add_969735;
  wire [7:0] sel_969736;
  wire [7:0] add_969739;
  wire [7:0] sel_969740;
  wire [7:0] add_969743;
  wire [7:0] sel_969744;
  wire [7:0] add_969747;
  wire [7:0] sel_969748;
  wire [7:0] add_969751;
  wire [7:0] sel_969752;
  wire [7:0] add_969755;
  wire [7:0] sel_969756;
  wire [7:0] add_969759;
  wire [7:0] sel_969760;
  wire [7:0] add_969763;
  wire [7:0] sel_969764;
  wire [7:0] add_969767;
  wire [7:0] sel_969768;
  wire [7:0] add_969771;
  wire [7:0] sel_969772;
  wire [7:0] add_969775;
  wire [7:0] sel_969776;
  wire [7:0] add_969779;
  wire [7:0] sel_969780;
  wire [7:0] add_969783;
  wire [7:0] sel_969784;
  wire [7:0] add_969787;
  wire [7:0] sel_969788;
  wire [7:0] add_969791;
  wire [7:0] sel_969792;
  wire [7:0] add_969795;
  wire [7:0] sel_969796;
  wire [7:0] add_969799;
  wire [7:0] sel_969800;
  wire [7:0] add_969803;
  wire [7:0] sel_969804;
  wire [7:0] add_969807;
  wire [7:0] sel_969808;
  wire [7:0] add_969811;
  wire [7:0] sel_969812;
  wire [7:0] add_969815;
  wire [7:0] sel_969816;
  wire [7:0] add_969819;
  wire [7:0] sel_969820;
  wire [7:0] add_969823;
  wire [7:0] sel_969824;
  wire [7:0] add_969827;
  wire [7:0] sel_969828;
  wire [7:0] add_969831;
  wire [7:0] sel_969832;
  wire [7:0] add_969835;
  wire [7:0] sel_969836;
  wire [7:0] add_969839;
  wire [7:0] sel_969840;
  wire [7:0] add_969843;
  wire [7:0] sel_969844;
  wire [7:0] add_969847;
  wire [7:0] sel_969848;
  wire [7:0] add_969851;
  wire [7:0] sel_969852;
  wire [7:0] add_969855;
  wire [7:0] sel_969856;
  wire [7:0] add_969859;
  wire [7:0] sel_969860;
  wire [7:0] add_969863;
  wire [7:0] sel_969864;
  wire [7:0] add_969867;
  wire [7:0] sel_969868;
  wire [7:0] add_969871;
  wire [7:0] sel_969872;
  wire [7:0] add_969875;
  wire [7:0] sel_969876;
  wire [7:0] add_969879;
  wire [7:0] sel_969880;
  wire [7:0] add_969883;
  wire [7:0] sel_969884;
  wire [7:0] add_969887;
  wire [7:0] sel_969888;
  wire [7:0] add_969891;
  wire [7:0] sel_969892;
  wire [7:0] add_969895;
  wire [7:0] sel_969896;
  wire [7:0] add_969899;
  wire [7:0] sel_969900;
  wire [7:0] add_969903;
  wire [7:0] sel_969904;
  wire [7:0] add_969907;
  wire [7:0] sel_969908;
  wire [7:0] add_969911;
  wire [7:0] sel_969912;
  wire [7:0] add_969915;
  wire [7:0] sel_969916;
  wire [7:0] add_969919;
  wire [7:0] sel_969920;
  wire [7:0] add_969923;
  wire [7:0] sel_969924;
  wire [7:0] add_969927;
  wire [7:0] sel_969928;
  wire [7:0] add_969931;
  wire [7:0] sel_969932;
  wire [7:0] add_969935;
  wire [7:0] sel_969936;
  wire [7:0] add_969939;
  wire [7:0] sel_969940;
  wire [7:0] add_969943;
  wire [7:0] sel_969944;
  wire [7:0] add_969947;
  wire [7:0] sel_969948;
  wire [7:0] add_969951;
  wire [7:0] sel_969952;
  wire [7:0] add_969955;
  wire [7:0] sel_969956;
  wire [7:0] add_969959;
  wire [7:0] sel_969960;
  wire [7:0] add_969963;
  wire [7:0] sel_969964;
  wire [7:0] add_969967;
  wire [7:0] sel_969968;
  wire [7:0] add_969971;
  wire [7:0] sel_969972;
  wire [7:0] add_969975;
  wire [7:0] sel_969976;
  wire [7:0] add_969979;
  wire [7:0] sel_969980;
  wire [7:0] add_969983;
  wire [7:0] sel_969984;
  wire [7:0] add_969987;
  wire [7:0] sel_969988;
  wire [7:0] add_969991;
  wire [7:0] sel_969992;
  wire [7:0] add_969996;
  wire [15:0] array_index_969997;
  wire [7:0] sel_969998;
  wire [7:0] add_970001;
  wire [7:0] sel_970002;
  wire [7:0] add_970005;
  wire [7:0] sel_970006;
  wire [7:0] add_970009;
  wire [7:0] sel_970010;
  wire [7:0] add_970013;
  wire [7:0] sel_970014;
  wire [7:0] add_970017;
  wire [7:0] sel_970018;
  wire [7:0] add_970021;
  wire [7:0] sel_970022;
  wire [7:0] add_970025;
  wire [7:0] sel_970026;
  wire [7:0] add_970029;
  wire [7:0] sel_970030;
  wire [7:0] add_970033;
  wire [7:0] sel_970034;
  wire [7:0] add_970037;
  wire [7:0] sel_970038;
  wire [7:0] add_970041;
  wire [7:0] sel_970042;
  wire [7:0] add_970045;
  wire [7:0] sel_970046;
  wire [7:0] add_970049;
  wire [7:0] sel_970050;
  wire [7:0] add_970053;
  wire [7:0] sel_970054;
  wire [7:0] add_970057;
  wire [7:0] sel_970058;
  wire [7:0] add_970061;
  wire [7:0] sel_970062;
  wire [7:0] add_970065;
  wire [7:0] sel_970066;
  wire [7:0] add_970069;
  wire [7:0] sel_970070;
  wire [7:0] add_970073;
  wire [7:0] sel_970074;
  wire [7:0] add_970077;
  wire [7:0] sel_970078;
  wire [7:0] add_970081;
  wire [7:0] sel_970082;
  wire [7:0] add_970085;
  wire [7:0] sel_970086;
  wire [7:0] add_970089;
  wire [7:0] sel_970090;
  wire [7:0] add_970093;
  wire [7:0] sel_970094;
  wire [7:0] add_970097;
  wire [7:0] sel_970098;
  wire [7:0] add_970101;
  wire [7:0] sel_970102;
  wire [7:0] add_970105;
  wire [7:0] sel_970106;
  wire [7:0] add_970109;
  wire [7:0] sel_970110;
  wire [7:0] add_970113;
  wire [7:0] sel_970114;
  wire [7:0] add_970117;
  wire [7:0] sel_970118;
  wire [7:0] add_970121;
  wire [7:0] sel_970122;
  wire [7:0] add_970125;
  wire [7:0] sel_970126;
  wire [7:0] add_970129;
  wire [7:0] sel_970130;
  wire [7:0] add_970133;
  wire [7:0] sel_970134;
  wire [7:0] add_970137;
  wire [7:0] sel_970138;
  wire [7:0] add_970141;
  wire [7:0] sel_970142;
  wire [7:0] add_970145;
  wire [7:0] sel_970146;
  wire [7:0] add_970149;
  wire [7:0] sel_970150;
  wire [7:0] add_970153;
  wire [7:0] sel_970154;
  wire [7:0] add_970157;
  wire [7:0] sel_970158;
  wire [7:0] add_970161;
  wire [7:0] sel_970162;
  wire [7:0] add_970165;
  wire [7:0] sel_970166;
  wire [7:0] add_970169;
  wire [7:0] sel_970170;
  wire [7:0] add_970173;
  wire [7:0] sel_970174;
  wire [7:0] add_970177;
  wire [7:0] sel_970178;
  wire [7:0] add_970181;
  wire [7:0] sel_970182;
  wire [7:0] add_970185;
  wire [7:0] sel_970186;
  wire [7:0] add_970189;
  wire [7:0] sel_970190;
  wire [7:0] add_970193;
  wire [7:0] sel_970194;
  wire [7:0] add_970197;
  wire [7:0] sel_970198;
  wire [7:0] add_970201;
  wire [7:0] sel_970202;
  wire [7:0] add_970205;
  wire [7:0] sel_970206;
  wire [7:0] add_970209;
  wire [7:0] sel_970210;
  wire [7:0] add_970213;
  wire [7:0] sel_970214;
  wire [7:0] add_970217;
  wire [7:0] sel_970218;
  wire [7:0] add_970221;
  wire [7:0] sel_970222;
  wire [7:0] add_970225;
  wire [7:0] sel_970226;
  wire [7:0] add_970229;
  wire [7:0] sel_970230;
  wire [7:0] add_970233;
  wire [7:0] sel_970234;
  wire [7:0] add_970237;
  wire [7:0] sel_970238;
  wire [7:0] add_970241;
  wire [7:0] sel_970242;
  wire [7:0] add_970245;
  wire [7:0] sel_970246;
  wire [7:0] add_970249;
  wire [7:0] sel_970250;
  wire [7:0] add_970253;
  wire [7:0] sel_970254;
  wire [7:0] add_970257;
  wire [7:0] sel_970258;
  wire [7:0] add_970261;
  wire [7:0] sel_970262;
  wire [7:0] add_970265;
  wire [7:0] sel_970266;
  wire [7:0] add_970269;
  wire [7:0] sel_970270;
  wire [7:0] add_970273;
  wire [7:0] sel_970274;
  wire [7:0] add_970277;
  wire [7:0] sel_970278;
  wire [7:0] add_970281;
  wire [7:0] sel_970282;
  wire [7:0] add_970285;
  wire [7:0] sel_970286;
  wire [7:0] add_970289;
  wire [7:0] sel_970290;
  wire [7:0] add_970293;
  wire [7:0] sel_970294;
  wire [7:0] add_970297;
  wire [7:0] sel_970298;
  wire [7:0] add_970301;
  wire [7:0] sel_970302;
  wire [7:0] add_970305;
  wire [7:0] sel_970306;
  wire [7:0] add_970309;
  wire [7:0] sel_970310;
  wire [7:0] add_970313;
  wire [7:0] sel_970314;
  wire [7:0] add_970317;
  wire [7:0] sel_970318;
  wire [7:0] add_970321;
  wire [7:0] sel_970322;
  wire [7:0] add_970325;
  wire [7:0] sel_970326;
  wire [7:0] add_970329;
  wire [7:0] sel_970330;
  wire [7:0] add_970333;
  wire [7:0] sel_970334;
  wire [7:0] add_970337;
  wire [7:0] sel_970338;
  wire [7:0] add_970341;
  wire [7:0] sel_970342;
  wire [7:0] add_970345;
  wire [7:0] sel_970346;
  wire [7:0] add_970349;
  wire [7:0] sel_970350;
  wire [7:0] add_970353;
  wire [7:0] sel_970354;
  wire [7:0] add_970357;
  wire [7:0] sel_970358;
  wire [7:0] add_970361;
  wire [7:0] sel_970362;
  wire [7:0] add_970365;
  wire [7:0] sel_970366;
  wire [7:0] add_970369;
  wire [7:0] sel_970370;
  wire [7:0] add_970373;
  wire [7:0] sel_970374;
  wire [7:0] add_970377;
  wire [7:0] sel_970378;
  wire [7:0] add_970381;
  wire [7:0] sel_970382;
  wire [7:0] add_970385;
  wire [7:0] sel_970386;
  wire [7:0] add_970389;
  wire [7:0] sel_970390;
  wire [7:0] add_970393;
  wire [7:0] sel_970394;
  wire [7:0] add_970398;
  wire [15:0] array_index_970399;
  wire [7:0] sel_970400;
  wire [7:0] add_970403;
  wire [7:0] sel_970404;
  wire [7:0] add_970407;
  wire [7:0] sel_970408;
  wire [7:0] add_970411;
  wire [7:0] sel_970412;
  wire [7:0] add_970415;
  wire [7:0] sel_970416;
  wire [7:0] add_970419;
  wire [7:0] sel_970420;
  wire [7:0] add_970423;
  wire [7:0] sel_970424;
  wire [7:0] add_970427;
  wire [7:0] sel_970428;
  wire [7:0] add_970431;
  wire [7:0] sel_970432;
  wire [7:0] add_970435;
  wire [7:0] sel_970436;
  wire [7:0] add_970439;
  wire [7:0] sel_970440;
  wire [7:0] add_970443;
  wire [7:0] sel_970444;
  wire [7:0] add_970447;
  wire [7:0] sel_970448;
  wire [7:0] add_970451;
  wire [7:0] sel_970452;
  wire [7:0] add_970455;
  wire [7:0] sel_970456;
  wire [7:0] add_970459;
  wire [7:0] sel_970460;
  wire [7:0] add_970463;
  wire [7:0] sel_970464;
  wire [7:0] add_970467;
  wire [7:0] sel_970468;
  wire [7:0] add_970471;
  wire [7:0] sel_970472;
  wire [7:0] add_970475;
  wire [7:0] sel_970476;
  wire [7:0] add_970479;
  wire [7:0] sel_970480;
  wire [7:0] add_970483;
  wire [7:0] sel_970484;
  wire [7:0] add_970487;
  wire [7:0] sel_970488;
  wire [7:0] add_970491;
  wire [7:0] sel_970492;
  wire [7:0] add_970495;
  wire [7:0] sel_970496;
  wire [7:0] add_970499;
  wire [7:0] sel_970500;
  wire [7:0] add_970503;
  wire [7:0] sel_970504;
  wire [7:0] add_970507;
  wire [7:0] sel_970508;
  wire [7:0] add_970511;
  wire [7:0] sel_970512;
  wire [7:0] add_970515;
  wire [7:0] sel_970516;
  wire [7:0] add_970519;
  wire [7:0] sel_970520;
  wire [7:0] add_970523;
  wire [7:0] sel_970524;
  wire [7:0] add_970527;
  wire [7:0] sel_970528;
  wire [7:0] add_970531;
  wire [7:0] sel_970532;
  wire [7:0] add_970535;
  wire [7:0] sel_970536;
  wire [7:0] add_970539;
  wire [7:0] sel_970540;
  wire [7:0] add_970543;
  wire [7:0] sel_970544;
  wire [7:0] add_970547;
  wire [7:0] sel_970548;
  wire [7:0] add_970551;
  wire [7:0] sel_970552;
  wire [7:0] add_970555;
  wire [7:0] sel_970556;
  wire [7:0] add_970559;
  wire [7:0] sel_970560;
  wire [7:0] add_970563;
  wire [7:0] sel_970564;
  wire [7:0] add_970567;
  wire [7:0] sel_970568;
  wire [7:0] add_970571;
  wire [7:0] sel_970572;
  wire [7:0] add_970575;
  wire [7:0] sel_970576;
  wire [7:0] add_970579;
  wire [7:0] sel_970580;
  wire [7:0] add_970583;
  wire [7:0] sel_970584;
  wire [7:0] add_970587;
  wire [7:0] sel_970588;
  wire [7:0] add_970591;
  wire [7:0] sel_970592;
  wire [7:0] add_970595;
  wire [7:0] sel_970596;
  wire [7:0] add_970599;
  wire [7:0] sel_970600;
  wire [7:0] add_970603;
  wire [7:0] sel_970604;
  wire [7:0] add_970607;
  wire [7:0] sel_970608;
  wire [7:0] add_970611;
  wire [7:0] sel_970612;
  wire [7:0] add_970615;
  wire [7:0] sel_970616;
  wire [7:0] add_970619;
  wire [7:0] sel_970620;
  wire [7:0] add_970623;
  wire [7:0] sel_970624;
  wire [7:0] add_970627;
  wire [7:0] sel_970628;
  wire [7:0] add_970631;
  wire [7:0] sel_970632;
  wire [7:0] add_970635;
  wire [7:0] sel_970636;
  wire [7:0] add_970639;
  wire [7:0] sel_970640;
  wire [7:0] add_970643;
  wire [7:0] sel_970644;
  wire [7:0] add_970647;
  wire [7:0] sel_970648;
  wire [7:0] add_970651;
  wire [7:0] sel_970652;
  wire [7:0] add_970655;
  wire [7:0] sel_970656;
  wire [7:0] add_970659;
  wire [7:0] sel_970660;
  wire [7:0] add_970663;
  wire [7:0] sel_970664;
  wire [7:0] add_970667;
  wire [7:0] sel_970668;
  wire [7:0] add_970671;
  wire [7:0] sel_970672;
  wire [7:0] add_970675;
  wire [7:0] sel_970676;
  wire [7:0] add_970679;
  wire [7:0] sel_970680;
  wire [7:0] add_970683;
  wire [7:0] sel_970684;
  wire [7:0] add_970687;
  wire [7:0] sel_970688;
  wire [7:0] add_970691;
  wire [7:0] sel_970692;
  wire [7:0] add_970695;
  wire [7:0] sel_970696;
  wire [7:0] add_970699;
  wire [7:0] sel_970700;
  wire [7:0] add_970703;
  wire [7:0] sel_970704;
  wire [7:0] add_970707;
  wire [7:0] sel_970708;
  wire [7:0] add_970711;
  wire [7:0] sel_970712;
  wire [7:0] add_970715;
  wire [7:0] sel_970716;
  wire [7:0] add_970719;
  wire [7:0] sel_970720;
  wire [7:0] add_970723;
  wire [7:0] sel_970724;
  wire [7:0] add_970727;
  wire [7:0] sel_970728;
  wire [7:0] add_970731;
  wire [7:0] sel_970732;
  wire [7:0] add_970735;
  wire [7:0] sel_970736;
  wire [7:0] add_970739;
  wire [7:0] sel_970740;
  wire [7:0] add_970743;
  wire [7:0] sel_970744;
  wire [7:0] add_970747;
  wire [7:0] sel_970748;
  wire [7:0] add_970751;
  wire [7:0] sel_970752;
  wire [7:0] add_970755;
  wire [7:0] sel_970756;
  wire [7:0] add_970759;
  wire [7:0] sel_970760;
  wire [7:0] add_970763;
  wire [7:0] sel_970764;
  wire [7:0] add_970767;
  wire [7:0] sel_970768;
  wire [7:0] add_970771;
  wire [7:0] sel_970772;
  wire [7:0] add_970775;
  wire [7:0] sel_970776;
  wire [7:0] add_970779;
  wire [7:0] sel_970780;
  wire [7:0] add_970783;
  wire [7:0] sel_970784;
  wire [7:0] add_970787;
  wire [7:0] sel_970788;
  wire [7:0] add_970791;
  wire [7:0] sel_970792;
  wire [7:0] add_970795;
  wire [7:0] sel_970796;
  wire [7:0] add_970800;
  wire [15:0] array_index_970801;
  wire [7:0] sel_970802;
  wire [7:0] add_970805;
  wire [7:0] sel_970806;
  wire [7:0] add_970809;
  wire [7:0] sel_970810;
  wire [7:0] add_970813;
  wire [7:0] sel_970814;
  wire [7:0] add_970817;
  wire [7:0] sel_970818;
  wire [7:0] add_970821;
  wire [7:0] sel_970822;
  wire [7:0] add_970825;
  wire [7:0] sel_970826;
  wire [7:0] add_970829;
  wire [7:0] sel_970830;
  wire [7:0] add_970833;
  wire [7:0] sel_970834;
  wire [7:0] add_970837;
  wire [7:0] sel_970838;
  wire [7:0] add_970841;
  wire [7:0] sel_970842;
  wire [7:0] add_970845;
  wire [7:0] sel_970846;
  wire [7:0] add_970849;
  wire [7:0] sel_970850;
  wire [7:0] add_970853;
  wire [7:0] sel_970854;
  wire [7:0] add_970857;
  wire [7:0] sel_970858;
  wire [7:0] add_970861;
  wire [7:0] sel_970862;
  wire [7:0] add_970865;
  wire [7:0] sel_970866;
  wire [7:0] add_970869;
  wire [7:0] sel_970870;
  wire [7:0] add_970873;
  wire [7:0] sel_970874;
  wire [7:0] add_970877;
  wire [7:0] sel_970878;
  wire [7:0] add_970881;
  wire [7:0] sel_970882;
  wire [7:0] add_970885;
  wire [7:0] sel_970886;
  wire [7:0] add_970889;
  wire [7:0] sel_970890;
  wire [7:0] add_970893;
  wire [7:0] sel_970894;
  wire [7:0] add_970897;
  wire [7:0] sel_970898;
  wire [7:0] add_970901;
  wire [7:0] sel_970902;
  wire [7:0] add_970905;
  wire [7:0] sel_970906;
  wire [7:0] add_970909;
  wire [7:0] sel_970910;
  wire [7:0] add_970913;
  wire [7:0] sel_970914;
  wire [7:0] add_970917;
  wire [7:0] sel_970918;
  wire [7:0] add_970921;
  wire [7:0] sel_970922;
  wire [7:0] add_970925;
  wire [7:0] sel_970926;
  wire [7:0] add_970929;
  wire [7:0] sel_970930;
  wire [7:0] add_970933;
  wire [7:0] sel_970934;
  wire [7:0] add_970937;
  wire [7:0] sel_970938;
  wire [7:0] add_970941;
  wire [7:0] sel_970942;
  wire [7:0] add_970945;
  wire [7:0] sel_970946;
  wire [7:0] add_970949;
  wire [7:0] sel_970950;
  wire [7:0] add_970953;
  wire [7:0] sel_970954;
  wire [7:0] add_970957;
  wire [7:0] sel_970958;
  wire [7:0] add_970961;
  wire [7:0] sel_970962;
  wire [7:0] add_970965;
  wire [7:0] sel_970966;
  wire [7:0] add_970969;
  wire [7:0] sel_970970;
  wire [7:0] add_970973;
  wire [7:0] sel_970974;
  wire [7:0] add_970977;
  wire [7:0] sel_970978;
  wire [7:0] add_970981;
  wire [7:0] sel_970982;
  wire [7:0] add_970985;
  wire [7:0] sel_970986;
  wire [7:0] add_970989;
  wire [7:0] sel_970990;
  wire [7:0] add_970993;
  wire [7:0] sel_970994;
  wire [7:0] add_970997;
  wire [7:0] sel_970998;
  wire [7:0] add_971001;
  wire [7:0] sel_971002;
  wire [7:0] add_971005;
  wire [7:0] sel_971006;
  wire [7:0] add_971009;
  wire [7:0] sel_971010;
  wire [7:0] add_971013;
  wire [7:0] sel_971014;
  wire [7:0] add_971017;
  wire [7:0] sel_971018;
  wire [7:0] add_971021;
  wire [7:0] sel_971022;
  wire [7:0] add_971025;
  wire [7:0] sel_971026;
  wire [7:0] add_971029;
  wire [7:0] sel_971030;
  wire [7:0] add_971033;
  wire [7:0] sel_971034;
  wire [7:0] add_971037;
  wire [7:0] sel_971038;
  wire [7:0] add_971041;
  wire [7:0] sel_971042;
  wire [7:0] add_971045;
  wire [7:0] sel_971046;
  wire [7:0] add_971049;
  wire [7:0] sel_971050;
  wire [7:0] add_971053;
  wire [7:0] sel_971054;
  wire [7:0] add_971057;
  wire [7:0] sel_971058;
  wire [7:0] add_971061;
  wire [7:0] sel_971062;
  wire [7:0] add_971065;
  wire [7:0] sel_971066;
  wire [7:0] add_971069;
  wire [7:0] sel_971070;
  wire [7:0] add_971073;
  wire [7:0] sel_971074;
  wire [7:0] add_971077;
  wire [7:0] sel_971078;
  wire [7:0] add_971081;
  wire [7:0] sel_971082;
  wire [7:0] add_971085;
  wire [7:0] sel_971086;
  wire [7:0] add_971089;
  wire [7:0] sel_971090;
  wire [7:0] add_971093;
  wire [7:0] sel_971094;
  wire [7:0] add_971097;
  wire [7:0] sel_971098;
  wire [7:0] add_971101;
  wire [7:0] sel_971102;
  wire [7:0] add_971105;
  wire [7:0] sel_971106;
  wire [7:0] add_971109;
  wire [7:0] sel_971110;
  wire [7:0] add_971113;
  wire [7:0] sel_971114;
  wire [7:0] add_971117;
  wire [7:0] sel_971118;
  wire [7:0] add_971121;
  wire [7:0] sel_971122;
  wire [7:0] add_971125;
  wire [7:0] sel_971126;
  wire [7:0] add_971129;
  wire [7:0] sel_971130;
  wire [7:0] add_971133;
  wire [7:0] sel_971134;
  wire [7:0] add_971137;
  wire [7:0] sel_971138;
  wire [7:0] add_971141;
  wire [7:0] sel_971142;
  wire [7:0] add_971145;
  wire [7:0] sel_971146;
  wire [7:0] add_971149;
  wire [7:0] sel_971150;
  wire [7:0] add_971153;
  wire [7:0] sel_971154;
  wire [7:0] add_971157;
  wire [7:0] sel_971158;
  wire [7:0] add_971161;
  wire [7:0] sel_971162;
  wire [7:0] add_971165;
  wire [7:0] sel_971166;
  wire [7:0] add_971169;
  wire [7:0] sel_971170;
  wire [7:0] add_971173;
  wire [7:0] sel_971174;
  wire [7:0] add_971177;
  wire [7:0] sel_971178;
  wire [7:0] add_971181;
  wire [7:0] sel_971182;
  wire [7:0] add_971185;
  wire [7:0] sel_971186;
  wire [7:0] add_971189;
  wire [7:0] sel_971190;
  wire [7:0] add_971193;
  wire [7:0] sel_971194;
  wire [7:0] add_971197;
  wire [7:0] sel_971198;
  wire [7:0] add_971202;
  wire [15:0] array_index_971203;
  wire [7:0] sel_971204;
  wire [7:0] add_971207;
  wire [7:0] sel_971208;
  wire [7:0] add_971211;
  wire [7:0] sel_971212;
  wire [7:0] add_971215;
  wire [7:0] sel_971216;
  wire [7:0] add_971219;
  wire [7:0] sel_971220;
  wire [7:0] add_971223;
  wire [7:0] sel_971224;
  wire [7:0] add_971227;
  wire [7:0] sel_971228;
  wire [7:0] add_971231;
  wire [7:0] sel_971232;
  wire [7:0] add_971235;
  wire [7:0] sel_971236;
  wire [7:0] add_971239;
  wire [7:0] sel_971240;
  wire [7:0] add_971243;
  wire [7:0] sel_971244;
  wire [7:0] add_971247;
  wire [7:0] sel_971248;
  wire [7:0] add_971251;
  wire [7:0] sel_971252;
  wire [7:0] add_971255;
  wire [7:0] sel_971256;
  wire [7:0] add_971259;
  wire [7:0] sel_971260;
  wire [7:0] add_971263;
  wire [7:0] sel_971264;
  wire [7:0] add_971267;
  wire [7:0] sel_971268;
  wire [7:0] add_971271;
  wire [7:0] sel_971272;
  wire [7:0] add_971275;
  wire [7:0] sel_971276;
  wire [7:0] add_971279;
  wire [7:0] sel_971280;
  wire [7:0] add_971283;
  wire [7:0] sel_971284;
  wire [7:0] add_971287;
  wire [7:0] sel_971288;
  wire [7:0] add_971291;
  wire [7:0] sel_971292;
  wire [7:0] add_971295;
  wire [7:0] sel_971296;
  wire [7:0] add_971299;
  wire [7:0] sel_971300;
  wire [7:0] add_971303;
  wire [7:0] sel_971304;
  wire [7:0] add_971307;
  wire [7:0] sel_971308;
  wire [7:0] add_971311;
  wire [7:0] sel_971312;
  wire [7:0] add_971315;
  wire [7:0] sel_971316;
  wire [7:0] add_971319;
  wire [7:0] sel_971320;
  wire [7:0] add_971323;
  wire [7:0] sel_971324;
  wire [7:0] add_971327;
  wire [7:0] sel_971328;
  wire [7:0] add_971331;
  wire [7:0] sel_971332;
  wire [7:0] add_971335;
  wire [7:0] sel_971336;
  wire [7:0] add_971339;
  wire [7:0] sel_971340;
  wire [7:0] add_971343;
  wire [7:0] sel_971344;
  wire [7:0] add_971347;
  wire [7:0] sel_971348;
  wire [7:0] add_971351;
  wire [7:0] sel_971352;
  wire [7:0] add_971355;
  wire [7:0] sel_971356;
  wire [7:0] add_971359;
  wire [7:0] sel_971360;
  wire [7:0] add_971363;
  wire [7:0] sel_971364;
  wire [7:0] add_971367;
  wire [7:0] sel_971368;
  wire [7:0] add_971371;
  wire [7:0] sel_971372;
  wire [7:0] add_971375;
  wire [7:0] sel_971376;
  wire [7:0] add_971379;
  wire [7:0] sel_971380;
  wire [7:0] add_971383;
  wire [7:0] sel_971384;
  wire [7:0] add_971387;
  wire [7:0] sel_971388;
  wire [7:0] add_971391;
  wire [7:0] sel_971392;
  wire [7:0] add_971395;
  wire [7:0] sel_971396;
  wire [7:0] add_971399;
  wire [7:0] sel_971400;
  wire [7:0] add_971403;
  wire [7:0] sel_971404;
  wire [7:0] add_971407;
  wire [7:0] sel_971408;
  wire [7:0] add_971411;
  wire [7:0] sel_971412;
  wire [7:0] add_971415;
  wire [7:0] sel_971416;
  wire [7:0] add_971419;
  wire [7:0] sel_971420;
  wire [7:0] add_971423;
  wire [7:0] sel_971424;
  wire [7:0] add_971427;
  wire [7:0] sel_971428;
  wire [7:0] add_971431;
  wire [7:0] sel_971432;
  wire [7:0] add_971435;
  wire [7:0] sel_971436;
  wire [7:0] add_971439;
  wire [7:0] sel_971440;
  wire [7:0] add_971443;
  wire [7:0] sel_971444;
  wire [7:0] add_971447;
  wire [7:0] sel_971448;
  wire [7:0] add_971451;
  wire [7:0] sel_971452;
  wire [7:0] add_971455;
  wire [7:0] sel_971456;
  wire [7:0] add_971459;
  wire [7:0] sel_971460;
  wire [7:0] add_971463;
  wire [7:0] sel_971464;
  wire [7:0] add_971467;
  wire [7:0] sel_971468;
  wire [7:0] add_971471;
  wire [7:0] sel_971472;
  wire [7:0] add_971475;
  wire [7:0] sel_971476;
  wire [7:0] add_971479;
  wire [7:0] sel_971480;
  wire [7:0] add_971483;
  wire [7:0] sel_971484;
  wire [7:0] add_971487;
  wire [7:0] sel_971488;
  wire [7:0] add_971491;
  wire [7:0] sel_971492;
  wire [7:0] add_971495;
  wire [7:0] sel_971496;
  wire [7:0] add_971499;
  wire [7:0] sel_971500;
  wire [7:0] add_971503;
  wire [7:0] sel_971504;
  wire [7:0] add_971507;
  wire [7:0] sel_971508;
  wire [7:0] add_971511;
  wire [7:0] sel_971512;
  wire [7:0] add_971515;
  wire [7:0] sel_971516;
  wire [7:0] add_971519;
  wire [7:0] sel_971520;
  wire [7:0] add_971523;
  wire [7:0] sel_971524;
  wire [7:0] add_971527;
  wire [7:0] sel_971528;
  wire [7:0] add_971531;
  wire [7:0] sel_971532;
  wire [7:0] add_971535;
  wire [7:0] sel_971536;
  wire [7:0] add_971539;
  wire [7:0] sel_971540;
  wire [7:0] add_971543;
  wire [7:0] sel_971544;
  wire [7:0] add_971547;
  wire [7:0] sel_971548;
  wire [7:0] add_971551;
  wire [7:0] sel_971552;
  wire [7:0] add_971555;
  wire [7:0] sel_971556;
  wire [7:0] add_971559;
  wire [7:0] sel_971560;
  wire [7:0] add_971563;
  wire [7:0] sel_971564;
  wire [7:0] add_971567;
  wire [7:0] sel_971568;
  wire [7:0] add_971571;
  wire [7:0] sel_971572;
  wire [7:0] add_971575;
  wire [7:0] sel_971576;
  wire [7:0] add_971579;
  wire [7:0] sel_971580;
  wire [7:0] add_971583;
  wire [7:0] sel_971584;
  wire [7:0] add_971587;
  wire [7:0] sel_971588;
  wire [7:0] add_971591;
  wire [7:0] sel_971592;
  wire [7:0] add_971595;
  wire [7:0] sel_971596;
  wire [7:0] add_971599;
  wire [7:0] sel_971600;
  wire [7:0] add_971604;
  wire [15:0] array_index_971605;
  wire [7:0] sel_971606;
  wire [7:0] add_971609;
  wire [7:0] sel_971610;
  wire [7:0] add_971613;
  wire [7:0] sel_971614;
  wire [7:0] add_971617;
  wire [7:0] sel_971618;
  wire [7:0] add_971621;
  wire [7:0] sel_971622;
  wire [7:0] add_971625;
  wire [7:0] sel_971626;
  wire [7:0] add_971629;
  wire [7:0] sel_971630;
  wire [7:0] add_971633;
  wire [7:0] sel_971634;
  wire [7:0] add_971637;
  wire [7:0] sel_971638;
  wire [7:0] add_971641;
  wire [7:0] sel_971642;
  wire [7:0] add_971645;
  wire [7:0] sel_971646;
  wire [7:0] add_971649;
  wire [7:0] sel_971650;
  wire [7:0] add_971653;
  wire [7:0] sel_971654;
  wire [7:0] add_971657;
  wire [7:0] sel_971658;
  wire [7:0] add_971661;
  wire [7:0] sel_971662;
  wire [7:0] add_971665;
  wire [7:0] sel_971666;
  wire [7:0] add_971669;
  wire [7:0] sel_971670;
  wire [7:0] add_971673;
  wire [7:0] sel_971674;
  wire [7:0] add_971677;
  wire [7:0] sel_971678;
  wire [7:0] add_971681;
  wire [7:0] sel_971682;
  wire [7:0] add_971685;
  wire [7:0] sel_971686;
  wire [7:0] add_971689;
  wire [7:0] sel_971690;
  wire [7:0] add_971693;
  wire [7:0] sel_971694;
  wire [7:0] add_971697;
  wire [7:0] sel_971698;
  wire [7:0] add_971701;
  wire [7:0] sel_971702;
  wire [7:0] add_971705;
  wire [7:0] sel_971706;
  wire [7:0] add_971709;
  wire [7:0] sel_971710;
  wire [7:0] add_971713;
  wire [7:0] sel_971714;
  wire [7:0] add_971717;
  wire [7:0] sel_971718;
  wire [7:0] add_971721;
  wire [7:0] sel_971722;
  wire [7:0] add_971725;
  wire [7:0] sel_971726;
  wire [7:0] add_971729;
  wire [7:0] sel_971730;
  wire [7:0] add_971733;
  wire [7:0] sel_971734;
  wire [7:0] add_971737;
  wire [7:0] sel_971738;
  wire [7:0] add_971741;
  wire [7:0] sel_971742;
  wire [7:0] add_971745;
  wire [7:0] sel_971746;
  wire [7:0] add_971749;
  wire [7:0] sel_971750;
  wire [7:0] add_971753;
  wire [7:0] sel_971754;
  wire [7:0] add_971757;
  wire [7:0] sel_971758;
  wire [7:0] add_971761;
  wire [7:0] sel_971762;
  wire [7:0] add_971765;
  wire [7:0] sel_971766;
  wire [7:0] add_971769;
  wire [7:0] sel_971770;
  wire [7:0] add_971773;
  wire [7:0] sel_971774;
  wire [7:0] add_971777;
  wire [7:0] sel_971778;
  wire [7:0] add_971781;
  wire [7:0] sel_971782;
  wire [7:0] add_971785;
  wire [7:0] sel_971786;
  wire [7:0] add_971789;
  wire [7:0] sel_971790;
  wire [7:0] add_971793;
  wire [7:0] sel_971794;
  wire [7:0] add_971797;
  wire [7:0] sel_971798;
  wire [7:0] add_971801;
  wire [7:0] sel_971802;
  wire [7:0] add_971805;
  wire [7:0] sel_971806;
  wire [7:0] add_971809;
  wire [7:0] sel_971810;
  wire [7:0] add_971813;
  wire [7:0] sel_971814;
  wire [7:0] add_971817;
  wire [7:0] sel_971818;
  wire [7:0] add_971821;
  wire [7:0] sel_971822;
  wire [7:0] add_971825;
  wire [7:0] sel_971826;
  wire [7:0] add_971829;
  wire [7:0] sel_971830;
  wire [7:0] add_971833;
  wire [7:0] sel_971834;
  wire [7:0] add_971837;
  wire [7:0] sel_971838;
  wire [7:0] add_971841;
  wire [7:0] sel_971842;
  wire [7:0] add_971845;
  wire [7:0] sel_971846;
  wire [7:0] add_971849;
  wire [7:0] sel_971850;
  wire [7:0] add_971853;
  wire [7:0] sel_971854;
  wire [7:0] add_971857;
  wire [7:0] sel_971858;
  wire [7:0] add_971861;
  wire [7:0] sel_971862;
  wire [7:0] add_971865;
  wire [7:0] sel_971866;
  wire [7:0] add_971869;
  wire [7:0] sel_971870;
  wire [7:0] add_971873;
  wire [7:0] sel_971874;
  wire [7:0] add_971877;
  wire [7:0] sel_971878;
  wire [7:0] add_971881;
  wire [7:0] sel_971882;
  wire [7:0] add_971885;
  wire [7:0] sel_971886;
  wire [7:0] add_971889;
  wire [7:0] sel_971890;
  wire [7:0] add_971893;
  wire [7:0] sel_971894;
  wire [7:0] add_971897;
  wire [7:0] sel_971898;
  wire [7:0] add_971901;
  wire [7:0] sel_971902;
  wire [7:0] add_971905;
  wire [7:0] sel_971906;
  wire [7:0] add_971909;
  wire [7:0] sel_971910;
  wire [7:0] add_971913;
  wire [7:0] sel_971914;
  wire [7:0] add_971917;
  wire [7:0] sel_971918;
  wire [7:0] add_971921;
  wire [7:0] sel_971922;
  wire [7:0] add_971925;
  wire [7:0] sel_971926;
  wire [7:0] add_971929;
  wire [7:0] sel_971930;
  wire [7:0] add_971933;
  wire [7:0] sel_971934;
  wire [7:0] add_971937;
  wire [7:0] sel_971938;
  wire [7:0] add_971941;
  wire [7:0] sel_971942;
  wire [7:0] add_971945;
  wire [7:0] sel_971946;
  wire [7:0] add_971949;
  wire [7:0] sel_971950;
  wire [7:0] add_971953;
  wire [7:0] sel_971954;
  wire [7:0] add_971957;
  wire [7:0] sel_971958;
  wire [7:0] add_971961;
  wire [7:0] sel_971962;
  wire [7:0] add_971965;
  wire [7:0] sel_971966;
  wire [7:0] add_971969;
  wire [7:0] sel_971970;
  wire [7:0] add_971973;
  wire [7:0] sel_971974;
  wire [7:0] add_971977;
  wire [7:0] sel_971978;
  wire [7:0] add_971981;
  wire [7:0] sel_971982;
  wire [7:0] add_971985;
  wire [7:0] sel_971986;
  wire [7:0] add_971989;
  wire [7:0] sel_971990;
  wire [7:0] add_971993;
  wire [7:0] sel_971994;
  wire [7:0] add_971997;
  wire [7:0] sel_971998;
  wire [7:0] add_972001;
  wire [7:0] sel_972002;
  wire [7:0] add_972006;
  wire [15:0] array_index_972007;
  wire [7:0] sel_972008;
  wire [7:0] add_972011;
  wire [7:0] sel_972012;
  wire [7:0] add_972015;
  wire [7:0] sel_972016;
  wire [7:0] add_972019;
  wire [7:0] sel_972020;
  wire [7:0] add_972023;
  wire [7:0] sel_972024;
  wire [7:0] add_972027;
  wire [7:0] sel_972028;
  wire [7:0] add_972031;
  wire [7:0] sel_972032;
  wire [7:0] add_972035;
  wire [7:0] sel_972036;
  wire [7:0] add_972039;
  wire [7:0] sel_972040;
  wire [7:0] add_972043;
  wire [7:0] sel_972044;
  wire [7:0] add_972047;
  wire [7:0] sel_972048;
  wire [7:0] add_972051;
  wire [7:0] sel_972052;
  wire [7:0] add_972055;
  wire [7:0] sel_972056;
  wire [7:0] add_972059;
  wire [7:0] sel_972060;
  wire [7:0] add_972063;
  wire [7:0] sel_972064;
  wire [7:0] add_972067;
  wire [7:0] sel_972068;
  wire [7:0] add_972071;
  wire [7:0] sel_972072;
  wire [7:0] add_972075;
  wire [7:0] sel_972076;
  wire [7:0] add_972079;
  wire [7:0] sel_972080;
  wire [7:0] add_972083;
  wire [7:0] sel_972084;
  wire [7:0] add_972087;
  wire [7:0] sel_972088;
  wire [7:0] add_972091;
  wire [7:0] sel_972092;
  wire [7:0] add_972095;
  wire [7:0] sel_972096;
  wire [7:0] add_972099;
  wire [7:0] sel_972100;
  wire [7:0] add_972103;
  wire [7:0] sel_972104;
  wire [7:0] add_972107;
  wire [7:0] sel_972108;
  wire [7:0] add_972111;
  wire [7:0] sel_972112;
  wire [7:0] add_972115;
  wire [7:0] sel_972116;
  wire [7:0] add_972119;
  wire [7:0] sel_972120;
  wire [7:0] add_972123;
  wire [7:0] sel_972124;
  wire [7:0] add_972127;
  wire [7:0] sel_972128;
  wire [7:0] add_972131;
  wire [7:0] sel_972132;
  wire [7:0] add_972135;
  wire [7:0] sel_972136;
  wire [7:0] add_972139;
  wire [7:0] sel_972140;
  wire [7:0] add_972143;
  wire [7:0] sel_972144;
  wire [7:0] add_972147;
  wire [7:0] sel_972148;
  wire [7:0] add_972151;
  wire [7:0] sel_972152;
  wire [7:0] add_972155;
  wire [7:0] sel_972156;
  wire [7:0] add_972159;
  wire [7:0] sel_972160;
  wire [7:0] add_972163;
  wire [7:0] sel_972164;
  wire [7:0] add_972167;
  wire [7:0] sel_972168;
  wire [7:0] add_972171;
  wire [7:0] sel_972172;
  wire [7:0] add_972175;
  wire [7:0] sel_972176;
  wire [7:0] add_972179;
  wire [7:0] sel_972180;
  wire [7:0] add_972183;
  wire [7:0] sel_972184;
  wire [7:0] add_972187;
  wire [7:0] sel_972188;
  wire [7:0] add_972191;
  wire [7:0] sel_972192;
  wire [7:0] add_972195;
  wire [7:0] sel_972196;
  wire [7:0] add_972199;
  wire [7:0] sel_972200;
  wire [7:0] add_972203;
  wire [7:0] sel_972204;
  wire [7:0] add_972207;
  wire [7:0] sel_972208;
  wire [7:0] add_972211;
  wire [7:0] sel_972212;
  wire [7:0] add_972215;
  wire [7:0] sel_972216;
  wire [7:0] add_972219;
  wire [7:0] sel_972220;
  wire [7:0] add_972223;
  wire [7:0] sel_972224;
  wire [7:0] add_972227;
  wire [7:0] sel_972228;
  wire [7:0] add_972231;
  wire [7:0] sel_972232;
  wire [7:0] add_972235;
  wire [7:0] sel_972236;
  wire [7:0] add_972239;
  wire [7:0] sel_972240;
  wire [7:0] add_972243;
  wire [7:0] sel_972244;
  wire [7:0] add_972247;
  wire [7:0] sel_972248;
  wire [7:0] add_972251;
  wire [7:0] sel_972252;
  wire [7:0] add_972255;
  wire [7:0] sel_972256;
  wire [7:0] add_972259;
  wire [7:0] sel_972260;
  wire [7:0] add_972263;
  wire [7:0] sel_972264;
  wire [7:0] add_972267;
  wire [7:0] sel_972268;
  wire [7:0] add_972271;
  wire [7:0] sel_972272;
  wire [7:0] add_972275;
  wire [7:0] sel_972276;
  wire [7:0] add_972279;
  wire [7:0] sel_972280;
  wire [7:0] add_972283;
  wire [7:0] sel_972284;
  wire [7:0] add_972287;
  wire [7:0] sel_972288;
  wire [7:0] add_972291;
  wire [7:0] sel_972292;
  wire [7:0] add_972295;
  wire [7:0] sel_972296;
  wire [7:0] add_972299;
  wire [7:0] sel_972300;
  wire [7:0] add_972303;
  wire [7:0] sel_972304;
  wire [7:0] add_972307;
  wire [7:0] sel_972308;
  wire [7:0] add_972311;
  wire [7:0] sel_972312;
  wire [7:0] add_972315;
  wire [7:0] sel_972316;
  wire [7:0] add_972319;
  wire [7:0] sel_972320;
  wire [7:0] add_972323;
  wire [7:0] sel_972324;
  wire [7:0] add_972327;
  wire [7:0] sel_972328;
  wire [7:0] add_972331;
  wire [7:0] sel_972332;
  wire [7:0] add_972335;
  wire [7:0] sel_972336;
  wire [7:0] add_972339;
  wire [7:0] sel_972340;
  wire [7:0] add_972343;
  wire [7:0] sel_972344;
  wire [7:0] add_972347;
  wire [7:0] sel_972348;
  wire [7:0] add_972351;
  wire [7:0] sel_972352;
  wire [7:0] add_972355;
  wire [7:0] sel_972356;
  wire [7:0] add_972359;
  wire [7:0] sel_972360;
  wire [7:0] add_972363;
  wire [7:0] sel_972364;
  wire [7:0] add_972367;
  wire [7:0] sel_972368;
  wire [7:0] add_972371;
  wire [7:0] sel_972372;
  wire [7:0] add_972375;
  wire [7:0] sel_972376;
  wire [7:0] add_972379;
  wire [7:0] sel_972380;
  wire [7:0] add_972383;
  wire [7:0] sel_972384;
  wire [7:0] add_972387;
  wire [7:0] sel_972388;
  wire [7:0] add_972391;
  wire [7:0] sel_972392;
  wire [7:0] add_972395;
  wire [7:0] sel_972396;
  wire [7:0] add_972399;
  wire [7:0] sel_972400;
  wire [7:0] add_972403;
  wire [7:0] sel_972404;
  wire [7:0] add_972408;
  wire [15:0] array_index_972409;
  wire [7:0] sel_972410;
  wire [7:0] add_972413;
  wire [7:0] sel_972414;
  wire [7:0] add_972417;
  wire [7:0] sel_972418;
  wire [7:0] add_972421;
  wire [7:0] sel_972422;
  wire [7:0] add_972425;
  wire [7:0] sel_972426;
  wire [7:0] add_972429;
  wire [7:0] sel_972430;
  wire [7:0] add_972433;
  wire [7:0] sel_972434;
  wire [7:0] add_972437;
  wire [7:0] sel_972438;
  wire [7:0] add_972441;
  wire [7:0] sel_972442;
  wire [7:0] add_972445;
  wire [7:0] sel_972446;
  wire [7:0] add_972449;
  wire [7:0] sel_972450;
  wire [7:0] add_972453;
  wire [7:0] sel_972454;
  wire [7:0] add_972457;
  wire [7:0] sel_972458;
  wire [7:0] add_972461;
  wire [7:0] sel_972462;
  wire [7:0] add_972465;
  wire [7:0] sel_972466;
  wire [7:0] add_972469;
  wire [7:0] sel_972470;
  wire [7:0] add_972473;
  wire [7:0] sel_972474;
  wire [7:0] add_972477;
  wire [7:0] sel_972478;
  wire [7:0] add_972481;
  wire [7:0] sel_972482;
  wire [7:0] add_972485;
  wire [7:0] sel_972486;
  wire [7:0] add_972489;
  wire [7:0] sel_972490;
  wire [7:0] add_972493;
  wire [7:0] sel_972494;
  wire [7:0] add_972497;
  wire [7:0] sel_972498;
  wire [7:0] add_972501;
  wire [7:0] sel_972502;
  wire [7:0] add_972505;
  wire [7:0] sel_972506;
  wire [7:0] add_972509;
  wire [7:0] sel_972510;
  wire [7:0] add_972513;
  wire [7:0] sel_972514;
  wire [7:0] add_972517;
  wire [7:0] sel_972518;
  wire [7:0] add_972521;
  wire [7:0] sel_972522;
  wire [7:0] add_972525;
  wire [7:0] sel_972526;
  wire [7:0] add_972529;
  wire [7:0] sel_972530;
  wire [7:0] add_972533;
  wire [7:0] sel_972534;
  wire [7:0] add_972537;
  wire [7:0] sel_972538;
  wire [7:0] add_972541;
  wire [7:0] sel_972542;
  wire [7:0] add_972545;
  wire [7:0] sel_972546;
  wire [7:0] add_972549;
  wire [7:0] sel_972550;
  wire [7:0] add_972553;
  wire [7:0] sel_972554;
  wire [7:0] add_972557;
  wire [7:0] sel_972558;
  wire [7:0] add_972561;
  wire [7:0] sel_972562;
  wire [7:0] add_972565;
  wire [7:0] sel_972566;
  wire [7:0] add_972569;
  wire [7:0] sel_972570;
  wire [7:0] add_972573;
  wire [7:0] sel_972574;
  wire [7:0] add_972577;
  wire [7:0] sel_972578;
  wire [7:0] add_972581;
  wire [7:0] sel_972582;
  wire [7:0] add_972585;
  wire [7:0] sel_972586;
  wire [7:0] add_972589;
  wire [7:0] sel_972590;
  wire [7:0] add_972593;
  wire [7:0] sel_972594;
  wire [7:0] add_972597;
  wire [7:0] sel_972598;
  wire [7:0] add_972601;
  wire [7:0] sel_972602;
  wire [7:0] add_972605;
  wire [7:0] sel_972606;
  wire [7:0] add_972609;
  wire [7:0] sel_972610;
  wire [7:0] add_972613;
  wire [7:0] sel_972614;
  wire [7:0] add_972617;
  wire [7:0] sel_972618;
  wire [7:0] add_972621;
  wire [7:0] sel_972622;
  wire [7:0] add_972625;
  wire [7:0] sel_972626;
  wire [7:0] add_972629;
  wire [7:0] sel_972630;
  wire [7:0] add_972633;
  wire [7:0] sel_972634;
  wire [7:0] add_972637;
  wire [7:0] sel_972638;
  wire [7:0] add_972641;
  wire [7:0] sel_972642;
  wire [7:0] add_972645;
  wire [7:0] sel_972646;
  wire [7:0] add_972649;
  wire [7:0] sel_972650;
  wire [7:0] add_972653;
  wire [7:0] sel_972654;
  wire [7:0] add_972657;
  wire [7:0] sel_972658;
  wire [7:0] add_972661;
  wire [7:0] sel_972662;
  wire [7:0] add_972665;
  wire [7:0] sel_972666;
  wire [7:0] add_972669;
  wire [7:0] sel_972670;
  wire [7:0] add_972673;
  wire [7:0] sel_972674;
  wire [7:0] add_972677;
  wire [7:0] sel_972678;
  wire [7:0] add_972681;
  wire [7:0] sel_972682;
  wire [7:0] add_972685;
  wire [7:0] sel_972686;
  wire [7:0] add_972689;
  wire [7:0] sel_972690;
  wire [7:0] add_972693;
  wire [7:0] sel_972694;
  wire [7:0] add_972697;
  wire [7:0] sel_972698;
  wire [7:0] add_972701;
  wire [7:0] sel_972702;
  wire [7:0] add_972705;
  wire [7:0] sel_972706;
  wire [7:0] add_972709;
  wire [7:0] sel_972710;
  wire [7:0] add_972713;
  wire [7:0] sel_972714;
  wire [7:0] add_972717;
  wire [7:0] sel_972718;
  wire [7:0] add_972721;
  wire [7:0] sel_972722;
  wire [7:0] add_972725;
  wire [7:0] sel_972726;
  wire [7:0] add_972729;
  wire [7:0] sel_972730;
  wire [7:0] add_972733;
  wire [7:0] sel_972734;
  wire [7:0] add_972737;
  wire [7:0] sel_972738;
  wire [7:0] add_972741;
  wire [7:0] sel_972742;
  wire [7:0] add_972745;
  wire [7:0] sel_972746;
  wire [7:0] add_972749;
  wire [7:0] sel_972750;
  wire [7:0] add_972753;
  wire [7:0] sel_972754;
  wire [7:0] add_972757;
  wire [7:0] sel_972758;
  wire [7:0] add_972761;
  wire [7:0] sel_972762;
  wire [7:0] add_972765;
  wire [7:0] sel_972766;
  wire [7:0] add_972769;
  wire [7:0] sel_972770;
  wire [7:0] add_972773;
  wire [7:0] sel_972774;
  wire [7:0] add_972777;
  wire [7:0] sel_972778;
  wire [7:0] add_972781;
  wire [7:0] sel_972782;
  wire [7:0] add_972785;
  wire [7:0] sel_972786;
  wire [7:0] add_972789;
  wire [7:0] sel_972790;
  wire [7:0] add_972793;
  wire [7:0] sel_972794;
  wire [7:0] add_972797;
  wire [7:0] sel_972798;
  wire [7:0] add_972801;
  wire [7:0] sel_972802;
  wire [7:0] add_972805;
  wire [7:0] sel_972806;
  wire [7:0] add_972810;
  wire [15:0] array_index_972811;
  wire [7:0] sel_972812;
  wire [7:0] add_972815;
  wire [7:0] sel_972816;
  wire [7:0] add_972819;
  wire [7:0] sel_972820;
  wire [7:0] add_972823;
  wire [7:0] sel_972824;
  wire [7:0] add_972827;
  wire [7:0] sel_972828;
  wire [7:0] add_972831;
  wire [7:0] sel_972832;
  wire [7:0] add_972835;
  wire [7:0] sel_972836;
  wire [7:0] add_972839;
  wire [7:0] sel_972840;
  wire [7:0] add_972843;
  wire [7:0] sel_972844;
  wire [7:0] add_972847;
  wire [7:0] sel_972848;
  wire [7:0] add_972851;
  wire [7:0] sel_972852;
  wire [7:0] add_972855;
  wire [7:0] sel_972856;
  wire [7:0] add_972859;
  wire [7:0] sel_972860;
  wire [7:0] add_972863;
  wire [7:0] sel_972864;
  wire [7:0] add_972867;
  wire [7:0] sel_972868;
  wire [7:0] add_972871;
  wire [7:0] sel_972872;
  wire [7:0] add_972875;
  wire [7:0] sel_972876;
  wire [7:0] add_972879;
  wire [7:0] sel_972880;
  wire [7:0] add_972883;
  wire [7:0] sel_972884;
  wire [7:0] add_972887;
  wire [7:0] sel_972888;
  wire [7:0] add_972891;
  wire [7:0] sel_972892;
  wire [7:0] add_972895;
  wire [7:0] sel_972896;
  wire [7:0] add_972899;
  wire [7:0] sel_972900;
  wire [7:0] add_972903;
  wire [7:0] sel_972904;
  wire [7:0] add_972907;
  wire [7:0] sel_972908;
  wire [7:0] add_972911;
  wire [7:0] sel_972912;
  wire [7:0] add_972915;
  wire [7:0] sel_972916;
  wire [7:0] add_972919;
  wire [7:0] sel_972920;
  wire [7:0] add_972923;
  wire [7:0] sel_972924;
  wire [7:0] add_972927;
  wire [7:0] sel_972928;
  wire [7:0] add_972931;
  wire [7:0] sel_972932;
  wire [7:0] add_972935;
  wire [7:0] sel_972936;
  wire [7:0] add_972939;
  wire [7:0] sel_972940;
  wire [7:0] add_972943;
  wire [7:0] sel_972944;
  wire [7:0] add_972947;
  wire [7:0] sel_972948;
  wire [7:0] add_972951;
  wire [7:0] sel_972952;
  wire [7:0] add_972955;
  wire [7:0] sel_972956;
  wire [7:0] add_972959;
  wire [7:0] sel_972960;
  wire [7:0] add_972963;
  wire [7:0] sel_972964;
  wire [7:0] add_972967;
  wire [7:0] sel_972968;
  wire [7:0] add_972971;
  wire [7:0] sel_972972;
  wire [7:0] add_972975;
  wire [7:0] sel_972976;
  wire [7:0] add_972979;
  wire [7:0] sel_972980;
  wire [7:0] add_972983;
  wire [7:0] sel_972984;
  wire [7:0] add_972987;
  wire [7:0] sel_972988;
  wire [7:0] add_972991;
  wire [7:0] sel_972992;
  wire [7:0] add_972995;
  wire [7:0] sel_972996;
  wire [7:0] add_972999;
  wire [7:0] sel_973000;
  wire [7:0] add_973003;
  wire [7:0] sel_973004;
  wire [7:0] add_973007;
  wire [7:0] sel_973008;
  wire [7:0] add_973011;
  wire [7:0] sel_973012;
  wire [7:0] add_973015;
  wire [7:0] sel_973016;
  wire [7:0] add_973019;
  wire [7:0] sel_973020;
  wire [7:0] add_973023;
  wire [7:0] sel_973024;
  wire [7:0] add_973027;
  wire [7:0] sel_973028;
  wire [7:0] add_973031;
  wire [7:0] sel_973032;
  wire [7:0] add_973035;
  wire [7:0] sel_973036;
  wire [7:0] add_973039;
  wire [7:0] sel_973040;
  wire [7:0] add_973043;
  wire [7:0] sel_973044;
  wire [7:0] add_973047;
  wire [7:0] sel_973048;
  wire [7:0] add_973051;
  wire [7:0] sel_973052;
  wire [7:0] add_973055;
  wire [7:0] sel_973056;
  wire [7:0] add_973059;
  wire [7:0] sel_973060;
  wire [7:0] add_973063;
  wire [7:0] sel_973064;
  wire [7:0] add_973067;
  wire [7:0] sel_973068;
  wire [7:0] add_973071;
  wire [7:0] sel_973072;
  wire [7:0] add_973075;
  wire [7:0] sel_973076;
  wire [7:0] add_973079;
  wire [7:0] sel_973080;
  wire [7:0] add_973083;
  wire [7:0] sel_973084;
  wire [7:0] add_973087;
  wire [7:0] sel_973088;
  wire [7:0] add_973091;
  wire [7:0] sel_973092;
  wire [7:0] add_973095;
  wire [7:0] sel_973096;
  wire [7:0] add_973099;
  wire [7:0] sel_973100;
  wire [7:0] add_973103;
  wire [7:0] sel_973104;
  wire [7:0] add_973107;
  wire [7:0] sel_973108;
  wire [7:0] add_973111;
  wire [7:0] sel_973112;
  wire [7:0] add_973115;
  wire [7:0] sel_973116;
  wire [7:0] add_973119;
  wire [7:0] sel_973120;
  wire [7:0] add_973123;
  wire [7:0] sel_973124;
  wire [7:0] add_973127;
  wire [7:0] sel_973128;
  wire [7:0] add_973131;
  wire [7:0] sel_973132;
  wire [7:0] add_973135;
  wire [7:0] sel_973136;
  wire [7:0] add_973139;
  wire [7:0] sel_973140;
  wire [7:0] add_973143;
  wire [7:0] sel_973144;
  wire [7:0] add_973147;
  wire [7:0] sel_973148;
  wire [7:0] add_973151;
  wire [7:0] sel_973152;
  wire [7:0] add_973155;
  wire [7:0] sel_973156;
  wire [7:0] add_973159;
  wire [7:0] sel_973160;
  wire [7:0] add_973163;
  wire [7:0] sel_973164;
  wire [7:0] add_973167;
  wire [7:0] sel_973168;
  wire [7:0] add_973171;
  wire [7:0] sel_973172;
  wire [7:0] add_973175;
  wire [7:0] sel_973176;
  wire [7:0] add_973179;
  wire [7:0] sel_973180;
  wire [7:0] add_973183;
  wire [7:0] sel_973184;
  wire [7:0] add_973187;
  wire [7:0] sel_973188;
  wire [7:0] add_973191;
  wire [7:0] sel_973192;
  wire [7:0] add_973195;
  wire [7:0] sel_973196;
  wire [7:0] add_973199;
  wire [7:0] sel_973200;
  wire [7:0] add_973203;
  wire [7:0] sel_973204;
  wire [7:0] add_973207;
  wire [7:0] sel_973208;
  wire [7:0] add_973212;
  wire [15:0] array_index_973213;
  wire [7:0] sel_973214;
  wire [7:0] add_973217;
  wire [7:0] sel_973218;
  wire [7:0] add_973221;
  wire [7:0] sel_973222;
  wire [7:0] add_973225;
  wire [7:0] sel_973226;
  wire [7:0] add_973229;
  wire [7:0] sel_973230;
  wire [7:0] add_973233;
  wire [7:0] sel_973234;
  wire [7:0] add_973237;
  wire [7:0] sel_973238;
  wire [7:0] add_973241;
  wire [7:0] sel_973242;
  wire [7:0] add_973245;
  wire [7:0] sel_973246;
  wire [7:0] add_973249;
  wire [7:0] sel_973250;
  wire [7:0] add_973253;
  wire [7:0] sel_973254;
  wire [7:0] add_973257;
  wire [7:0] sel_973258;
  wire [7:0] add_973261;
  wire [7:0] sel_973262;
  wire [7:0] add_973265;
  wire [7:0] sel_973266;
  wire [7:0] add_973269;
  wire [7:0] sel_973270;
  wire [7:0] add_973273;
  wire [7:0] sel_973274;
  wire [7:0] add_973277;
  wire [7:0] sel_973278;
  wire [7:0] add_973281;
  wire [7:0] sel_973282;
  wire [7:0] add_973285;
  wire [7:0] sel_973286;
  wire [7:0] add_973289;
  wire [7:0] sel_973290;
  wire [7:0] add_973293;
  wire [7:0] sel_973294;
  wire [7:0] add_973297;
  wire [7:0] sel_973298;
  wire [7:0] add_973301;
  wire [7:0] sel_973302;
  wire [7:0] add_973305;
  wire [7:0] sel_973306;
  wire [7:0] add_973309;
  wire [7:0] sel_973310;
  wire [7:0] add_973313;
  wire [7:0] sel_973314;
  wire [7:0] add_973317;
  wire [7:0] sel_973318;
  wire [7:0] add_973321;
  wire [7:0] sel_973322;
  wire [7:0] add_973325;
  wire [7:0] sel_973326;
  wire [7:0] add_973329;
  wire [7:0] sel_973330;
  wire [7:0] add_973333;
  wire [7:0] sel_973334;
  wire [7:0] add_973337;
  wire [7:0] sel_973338;
  wire [7:0] add_973341;
  wire [7:0] sel_973342;
  wire [7:0] add_973345;
  wire [7:0] sel_973346;
  wire [7:0] add_973349;
  wire [7:0] sel_973350;
  wire [7:0] add_973353;
  wire [7:0] sel_973354;
  wire [7:0] add_973357;
  wire [7:0] sel_973358;
  wire [7:0] add_973361;
  wire [7:0] sel_973362;
  wire [7:0] add_973365;
  wire [7:0] sel_973366;
  wire [7:0] add_973369;
  wire [7:0] sel_973370;
  wire [7:0] add_973373;
  wire [7:0] sel_973374;
  wire [7:0] add_973377;
  wire [7:0] sel_973378;
  wire [7:0] add_973381;
  wire [7:0] sel_973382;
  wire [7:0] add_973385;
  wire [7:0] sel_973386;
  wire [7:0] add_973389;
  wire [7:0] sel_973390;
  wire [7:0] add_973393;
  wire [7:0] sel_973394;
  wire [7:0] add_973397;
  wire [7:0] sel_973398;
  wire [7:0] add_973401;
  wire [7:0] sel_973402;
  wire [7:0] add_973405;
  wire [7:0] sel_973406;
  wire [7:0] add_973409;
  wire [7:0] sel_973410;
  wire [7:0] add_973413;
  wire [7:0] sel_973414;
  wire [7:0] add_973417;
  wire [7:0] sel_973418;
  wire [7:0] add_973421;
  wire [7:0] sel_973422;
  wire [7:0] add_973425;
  wire [7:0] sel_973426;
  wire [7:0] add_973429;
  wire [7:0] sel_973430;
  wire [7:0] add_973433;
  wire [7:0] sel_973434;
  wire [7:0] add_973437;
  wire [7:0] sel_973438;
  wire [7:0] add_973441;
  wire [7:0] sel_973442;
  wire [7:0] add_973445;
  wire [7:0] sel_973446;
  wire [7:0] add_973449;
  wire [7:0] sel_973450;
  wire [7:0] add_973453;
  wire [7:0] sel_973454;
  wire [7:0] add_973457;
  wire [7:0] sel_973458;
  wire [7:0] add_973461;
  wire [7:0] sel_973462;
  wire [7:0] add_973465;
  wire [7:0] sel_973466;
  wire [7:0] add_973469;
  wire [7:0] sel_973470;
  wire [7:0] add_973473;
  wire [7:0] sel_973474;
  wire [7:0] add_973477;
  wire [7:0] sel_973478;
  wire [7:0] add_973481;
  wire [7:0] sel_973482;
  wire [7:0] add_973485;
  wire [7:0] sel_973486;
  wire [7:0] add_973489;
  wire [7:0] sel_973490;
  wire [7:0] add_973493;
  wire [7:0] sel_973494;
  wire [7:0] add_973497;
  wire [7:0] sel_973498;
  wire [7:0] add_973501;
  wire [7:0] sel_973502;
  wire [7:0] add_973505;
  wire [7:0] sel_973506;
  wire [7:0] add_973509;
  wire [7:0] sel_973510;
  wire [7:0] add_973513;
  wire [7:0] sel_973514;
  wire [7:0] add_973517;
  wire [7:0] sel_973518;
  wire [7:0] add_973521;
  wire [7:0] sel_973522;
  wire [7:0] add_973525;
  wire [7:0] sel_973526;
  wire [7:0] add_973529;
  wire [7:0] sel_973530;
  wire [7:0] add_973533;
  wire [7:0] sel_973534;
  wire [7:0] add_973537;
  wire [7:0] sel_973538;
  wire [7:0] add_973541;
  wire [7:0] sel_973542;
  wire [7:0] add_973545;
  wire [7:0] sel_973546;
  wire [7:0] add_973549;
  wire [7:0] sel_973550;
  wire [7:0] add_973553;
  wire [7:0] sel_973554;
  wire [7:0] add_973557;
  wire [7:0] sel_973558;
  wire [7:0] add_973561;
  wire [7:0] sel_973562;
  wire [7:0] add_973565;
  wire [7:0] sel_973566;
  wire [7:0] add_973569;
  wire [7:0] sel_973570;
  wire [7:0] add_973573;
  wire [7:0] sel_973574;
  wire [7:0] add_973577;
  wire [7:0] sel_973578;
  wire [7:0] add_973581;
  wire [7:0] sel_973582;
  wire [7:0] add_973585;
  wire [7:0] sel_973586;
  wire [7:0] add_973589;
  wire [7:0] sel_973590;
  wire [7:0] add_973593;
  wire [7:0] sel_973594;
  wire [7:0] add_973597;
  wire [7:0] sel_973598;
  wire [7:0] add_973601;
  wire [7:0] sel_973602;
  wire [7:0] add_973605;
  wire [7:0] sel_973606;
  wire [7:0] add_973609;
  wire [7:0] sel_973610;
  wire [7:0] add_973614;
  wire [15:0] array_index_973615;
  wire [7:0] sel_973616;
  wire [7:0] add_973619;
  wire [7:0] sel_973620;
  wire [7:0] add_973623;
  wire [7:0] sel_973624;
  wire [7:0] add_973627;
  wire [7:0] sel_973628;
  wire [7:0] add_973631;
  wire [7:0] sel_973632;
  wire [7:0] add_973635;
  wire [7:0] sel_973636;
  wire [7:0] add_973639;
  wire [7:0] sel_973640;
  wire [7:0] add_973643;
  wire [7:0] sel_973644;
  wire [7:0] add_973647;
  wire [7:0] sel_973648;
  wire [7:0] add_973651;
  wire [7:0] sel_973652;
  wire [7:0] add_973655;
  wire [7:0] sel_973656;
  wire [7:0] add_973659;
  wire [7:0] sel_973660;
  wire [7:0] add_973663;
  wire [7:0] sel_973664;
  wire [7:0] add_973667;
  wire [7:0] sel_973668;
  wire [7:0] add_973671;
  wire [7:0] sel_973672;
  wire [7:0] add_973675;
  wire [7:0] sel_973676;
  wire [7:0] add_973679;
  wire [7:0] sel_973680;
  wire [7:0] add_973683;
  wire [7:0] sel_973684;
  wire [7:0] add_973687;
  wire [7:0] sel_973688;
  wire [7:0] add_973691;
  wire [7:0] sel_973692;
  wire [7:0] add_973695;
  wire [7:0] sel_973696;
  wire [7:0] add_973699;
  wire [7:0] sel_973700;
  wire [7:0] add_973703;
  wire [7:0] sel_973704;
  wire [7:0] add_973707;
  wire [7:0] sel_973708;
  wire [7:0] add_973711;
  wire [7:0] sel_973712;
  wire [7:0] add_973715;
  wire [7:0] sel_973716;
  wire [7:0] add_973719;
  wire [7:0] sel_973720;
  wire [7:0] add_973723;
  wire [7:0] sel_973724;
  wire [7:0] add_973727;
  wire [7:0] sel_973728;
  wire [7:0] add_973731;
  wire [7:0] sel_973732;
  wire [7:0] add_973735;
  wire [7:0] sel_973736;
  wire [7:0] add_973739;
  wire [7:0] sel_973740;
  wire [7:0] add_973743;
  wire [7:0] sel_973744;
  wire [7:0] add_973747;
  wire [7:0] sel_973748;
  wire [7:0] add_973751;
  wire [7:0] sel_973752;
  wire [7:0] add_973755;
  wire [7:0] sel_973756;
  wire [7:0] add_973759;
  wire [7:0] sel_973760;
  wire [7:0] add_973763;
  wire [7:0] sel_973764;
  wire [7:0] add_973767;
  wire [7:0] sel_973768;
  wire [7:0] add_973771;
  wire [7:0] sel_973772;
  wire [7:0] add_973775;
  wire [7:0] sel_973776;
  wire [7:0] add_973779;
  wire [7:0] sel_973780;
  wire [7:0] add_973783;
  wire [7:0] sel_973784;
  wire [7:0] add_973787;
  wire [7:0] sel_973788;
  wire [7:0] add_973791;
  wire [7:0] sel_973792;
  wire [7:0] add_973795;
  wire [7:0] sel_973796;
  wire [7:0] add_973799;
  wire [7:0] sel_973800;
  wire [7:0] add_973803;
  wire [7:0] sel_973804;
  wire [7:0] add_973807;
  wire [7:0] sel_973808;
  wire [7:0] add_973811;
  wire [7:0] sel_973812;
  wire [7:0] add_973815;
  wire [7:0] sel_973816;
  wire [7:0] add_973819;
  wire [7:0] sel_973820;
  wire [7:0] add_973823;
  wire [7:0] sel_973824;
  wire [7:0] add_973827;
  wire [7:0] sel_973828;
  wire [7:0] add_973831;
  wire [7:0] sel_973832;
  wire [7:0] add_973835;
  wire [7:0] sel_973836;
  wire [7:0] add_973839;
  wire [7:0] sel_973840;
  wire [7:0] add_973843;
  wire [7:0] sel_973844;
  wire [7:0] add_973847;
  wire [7:0] sel_973848;
  wire [7:0] add_973851;
  wire [7:0] sel_973852;
  wire [7:0] add_973855;
  wire [7:0] sel_973856;
  wire [7:0] add_973859;
  wire [7:0] sel_973860;
  wire [7:0] add_973863;
  wire [7:0] sel_973864;
  wire [7:0] add_973867;
  wire [7:0] sel_973868;
  wire [7:0] add_973871;
  wire [7:0] sel_973872;
  wire [7:0] add_973875;
  wire [7:0] sel_973876;
  wire [7:0] add_973879;
  wire [7:0] sel_973880;
  wire [7:0] add_973883;
  wire [7:0] sel_973884;
  wire [7:0] add_973887;
  wire [7:0] sel_973888;
  wire [7:0] add_973891;
  wire [7:0] sel_973892;
  wire [7:0] add_973895;
  wire [7:0] sel_973896;
  wire [7:0] add_973899;
  wire [7:0] sel_973900;
  wire [7:0] add_973903;
  wire [7:0] sel_973904;
  wire [7:0] add_973907;
  wire [7:0] sel_973908;
  wire [7:0] add_973911;
  wire [7:0] sel_973912;
  wire [7:0] add_973915;
  wire [7:0] sel_973916;
  wire [7:0] add_973919;
  wire [7:0] sel_973920;
  wire [7:0] add_973923;
  wire [7:0] sel_973924;
  wire [7:0] add_973927;
  wire [7:0] sel_973928;
  wire [7:0] add_973931;
  wire [7:0] sel_973932;
  wire [7:0] add_973935;
  wire [7:0] sel_973936;
  wire [7:0] add_973939;
  wire [7:0] sel_973940;
  wire [7:0] add_973943;
  wire [7:0] sel_973944;
  wire [7:0] add_973947;
  wire [7:0] sel_973948;
  wire [7:0] add_973951;
  wire [7:0] sel_973952;
  wire [7:0] add_973955;
  wire [7:0] sel_973956;
  wire [7:0] add_973959;
  wire [7:0] sel_973960;
  wire [7:0] add_973963;
  wire [7:0] sel_973964;
  wire [7:0] add_973967;
  wire [7:0] sel_973968;
  wire [7:0] add_973971;
  wire [7:0] sel_973972;
  wire [7:0] add_973975;
  wire [7:0] sel_973976;
  wire [7:0] add_973979;
  wire [7:0] sel_973980;
  wire [7:0] add_973983;
  wire [7:0] sel_973984;
  wire [7:0] add_973987;
  wire [7:0] sel_973988;
  wire [7:0] add_973991;
  wire [7:0] sel_973992;
  wire [7:0] add_973995;
  wire [7:0] sel_973996;
  wire [7:0] add_973999;
  wire [7:0] sel_974000;
  wire [7:0] add_974003;
  wire [7:0] sel_974004;
  wire [7:0] add_974007;
  wire [7:0] sel_974008;
  wire [7:0] add_974011;
  wire [7:0] sel_974012;
  wire [7:0] add_974016;
  wire [15:0] array_index_974017;
  wire [7:0] sel_974018;
  wire [7:0] add_974021;
  wire [7:0] sel_974022;
  wire [7:0] add_974025;
  wire [7:0] sel_974026;
  wire [7:0] add_974029;
  wire [7:0] sel_974030;
  wire [7:0] add_974033;
  wire [7:0] sel_974034;
  wire [7:0] add_974037;
  wire [7:0] sel_974038;
  wire [7:0] add_974041;
  wire [7:0] sel_974042;
  wire [7:0] add_974045;
  wire [7:0] sel_974046;
  wire [7:0] add_974049;
  wire [7:0] sel_974050;
  wire [7:0] add_974053;
  wire [7:0] sel_974054;
  wire [7:0] add_974057;
  wire [7:0] sel_974058;
  wire [7:0] add_974061;
  wire [7:0] sel_974062;
  wire [7:0] add_974065;
  wire [7:0] sel_974066;
  wire [7:0] add_974069;
  wire [7:0] sel_974070;
  wire [7:0] add_974073;
  wire [7:0] sel_974074;
  wire [7:0] add_974077;
  wire [7:0] sel_974078;
  wire [7:0] add_974081;
  wire [7:0] sel_974082;
  wire [7:0] add_974085;
  wire [7:0] sel_974086;
  wire [7:0] add_974089;
  wire [7:0] sel_974090;
  wire [7:0] add_974093;
  wire [7:0] sel_974094;
  wire [7:0] add_974097;
  wire [7:0] sel_974098;
  wire [7:0] add_974101;
  wire [7:0] sel_974102;
  wire [7:0] add_974105;
  wire [7:0] sel_974106;
  wire [7:0] add_974109;
  wire [7:0] sel_974110;
  wire [7:0] add_974113;
  wire [7:0] sel_974114;
  wire [7:0] add_974117;
  wire [7:0] sel_974118;
  wire [7:0] add_974121;
  wire [7:0] sel_974122;
  wire [7:0] add_974125;
  wire [7:0] sel_974126;
  wire [7:0] add_974129;
  wire [7:0] sel_974130;
  wire [7:0] add_974133;
  wire [7:0] sel_974134;
  wire [7:0] add_974137;
  wire [7:0] sel_974138;
  wire [7:0] add_974141;
  wire [7:0] sel_974142;
  wire [7:0] add_974145;
  wire [7:0] sel_974146;
  wire [7:0] add_974149;
  wire [7:0] sel_974150;
  wire [7:0] add_974153;
  wire [7:0] sel_974154;
  wire [7:0] add_974157;
  wire [7:0] sel_974158;
  wire [7:0] add_974161;
  wire [7:0] sel_974162;
  wire [7:0] add_974165;
  wire [7:0] sel_974166;
  wire [7:0] add_974169;
  wire [7:0] sel_974170;
  wire [7:0] add_974173;
  wire [7:0] sel_974174;
  wire [7:0] add_974177;
  wire [7:0] sel_974178;
  wire [7:0] add_974181;
  wire [7:0] sel_974182;
  wire [7:0] add_974185;
  wire [7:0] sel_974186;
  wire [7:0] add_974189;
  wire [7:0] sel_974190;
  wire [7:0] add_974193;
  wire [7:0] sel_974194;
  wire [7:0] add_974197;
  wire [7:0] sel_974198;
  wire [7:0] add_974201;
  wire [7:0] sel_974202;
  wire [7:0] add_974205;
  wire [7:0] sel_974206;
  wire [7:0] add_974209;
  wire [7:0] sel_974210;
  wire [7:0] add_974213;
  wire [7:0] sel_974214;
  wire [7:0] add_974217;
  wire [7:0] sel_974218;
  wire [7:0] add_974221;
  wire [7:0] sel_974222;
  wire [7:0] add_974225;
  wire [7:0] sel_974226;
  wire [7:0] add_974229;
  wire [7:0] sel_974230;
  wire [7:0] add_974233;
  wire [7:0] sel_974234;
  wire [7:0] add_974237;
  wire [7:0] sel_974238;
  wire [7:0] add_974241;
  wire [7:0] sel_974242;
  wire [7:0] add_974245;
  wire [7:0] sel_974246;
  wire [7:0] add_974249;
  wire [7:0] sel_974250;
  wire [7:0] add_974253;
  wire [7:0] sel_974254;
  wire [7:0] add_974257;
  wire [7:0] sel_974258;
  wire [7:0] add_974261;
  wire [7:0] sel_974262;
  wire [7:0] add_974265;
  wire [7:0] sel_974266;
  wire [7:0] add_974269;
  wire [7:0] sel_974270;
  wire [7:0] add_974273;
  wire [7:0] sel_974274;
  wire [7:0] add_974277;
  wire [7:0] sel_974278;
  wire [7:0] add_974281;
  wire [7:0] sel_974282;
  wire [7:0] add_974285;
  wire [7:0] sel_974286;
  wire [7:0] add_974289;
  wire [7:0] sel_974290;
  wire [7:0] add_974293;
  wire [7:0] sel_974294;
  wire [7:0] add_974297;
  wire [7:0] sel_974298;
  wire [7:0] add_974301;
  wire [7:0] sel_974302;
  wire [7:0] add_974305;
  wire [7:0] sel_974306;
  wire [7:0] add_974309;
  wire [7:0] sel_974310;
  wire [7:0] add_974313;
  wire [7:0] sel_974314;
  wire [7:0] add_974317;
  wire [7:0] sel_974318;
  wire [7:0] add_974321;
  wire [7:0] sel_974322;
  wire [7:0] add_974325;
  wire [7:0] sel_974326;
  wire [7:0] add_974329;
  wire [7:0] sel_974330;
  wire [7:0] add_974333;
  wire [7:0] sel_974334;
  wire [7:0] add_974337;
  wire [7:0] sel_974338;
  wire [7:0] add_974341;
  wire [7:0] sel_974342;
  wire [7:0] add_974345;
  wire [7:0] sel_974346;
  wire [7:0] add_974349;
  wire [7:0] sel_974350;
  wire [7:0] add_974353;
  wire [7:0] sel_974354;
  wire [7:0] add_974357;
  wire [7:0] sel_974358;
  wire [7:0] add_974361;
  wire [7:0] sel_974362;
  wire [7:0] add_974365;
  wire [7:0] sel_974366;
  wire [7:0] add_974369;
  wire [7:0] sel_974370;
  wire [7:0] add_974373;
  wire [7:0] sel_974374;
  wire [7:0] add_974377;
  wire [7:0] sel_974378;
  wire [7:0] add_974381;
  wire [7:0] sel_974382;
  wire [7:0] add_974385;
  wire [7:0] sel_974386;
  wire [7:0] add_974389;
  wire [7:0] sel_974390;
  wire [7:0] add_974393;
  wire [7:0] sel_974394;
  wire [7:0] add_974397;
  wire [7:0] sel_974398;
  wire [7:0] add_974401;
  wire [7:0] sel_974402;
  wire [7:0] add_974405;
  wire [7:0] sel_974406;
  wire [7:0] add_974409;
  wire [7:0] sel_974410;
  wire [7:0] add_974413;
  wire [7:0] sel_974414;
  wire [7:0] add_974418;
  wire [15:0] array_index_974419;
  wire [7:0] sel_974420;
  wire [7:0] add_974423;
  wire [7:0] sel_974424;
  wire [7:0] add_974427;
  wire [7:0] sel_974428;
  wire [7:0] add_974431;
  wire [7:0] sel_974432;
  wire [7:0] add_974435;
  wire [7:0] sel_974436;
  wire [7:0] add_974439;
  wire [7:0] sel_974440;
  wire [7:0] add_974443;
  wire [7:0] sel_974444;
  wire [7:0] add_974447;
  wire [7:0] sel_974448;
  wire [7:0] add_974451;
  wire [7:0] sel_974452;
  wire [7:0] add_974455;
  wire [7:0] sel_974456;
  wire [7:0] add_974459;
  wire [7:0] sel_974460;
  wire [7:0] add_974463;
  wire [7:0] sel_974464;
  wire [7:0] add_974467;
  wire [7:0] sel_974468;
  wire [7:0] add_974471;
  wire [7:0] sel_974472;
  wire [7:0] add_974475;
  wire [7:0] sel_974476;
  wire [7:0] add_974479;
  wire [7:0] sel_974480;
  wire [7:0] add_974483;
  wire [7:0] sel_974484;
  wire [7:0] add_974487;
  wire [7:0] sel_974488;
  wire [7:0] add_974491;
  wire [7:0] sel_974492;
  wire [7:0] add_974495;
  wire [7:0] sel_974496;
  wire [7:0] add_974499;
  wire [7:0] sel_974500;
  wire [7:0] add_974503;
  wire [7:0] sel_974504;
  wire [7:0] add_974507;
  wire [7:0] sel_974508;
  wire [7:0] add_974511;
  wire [7:0] sel_974512;
  wire [7:0] add_974515;
  wire [7:0] sel_974516;
  wire [7:0] add_974519;
  wire [7:0] sel_974520;
  wire [7:0] add_974523;
  wire [7:0] sel_974524;
  wire [7:0] add_974527;
  wire [7:0] sel_974528;
  wire [7:0] add_974531;
  wire [7:0] sel_974532;
  wire [7:0] add_974535;
  wire [7:0] sel_974536;
  wire [7:0] add_974539;
  wire [7:0] sel_974540;
  wire [7:0] add_974543;
  wire [7:0] sel_974544;
  wire [7:0] add_974547;
  wire [7:0] sel_974548;
  wire [7:0] add_974551;
  wire [7:0] sel_974552;
  wire [7:0] add_974555;
  wire [7:0] sel_974556;
  wire [7:0] add_974559;
  wire [7:0] sel_974560;
  wire [7:0] add_974563;
  wire [7:0] sel_974564;
  wire [7:0] add_974567;
  wire [7:0] sel_974568;
  wire [7:0] add_974571;
  wire [7:0] sel_974572;
  wire [7:0] add_974575;
  wire [7:0] sel_974576;
  wire [7:0] add_974579;
  wire [7:0] sel_974580;
  wire [7:0] add_974583;
  wire [7:0] sel_974584;
  wire [7:0] add_974587;
  wire [7:0] sel_974588;
  wire [7:0] add_974591;
  wire [7:0] sel_974592;
  wire [7:0] add_974595;
  wire [7:0] sel_974596;
  wire [7:0] add_974599;
  wire [7:0] sel_974600;
  wire [7:0] add_974603;
  wire [7:0] sel_974604;
  wire [7:0] add_974607;
  wire [7:0] sel_974608;
  wire [7:0] add_974611;
  wire [7:0] sel_974612;
  wire [7:0] add_974615;
  wire [7:0] sel_974616;
  wire [7:0] add_974619;
  wire [7:0] sel_974620;
  wire [7:0] add_974623;
  wire [7:0] sel_974624;
  wire [7:0] add_974627;
  wire [7:0] sel_974628;
  wire [7:0] add_974631;
  wire [7:0] sel_974632;
  wire [7:0] add_974635;
  wire [7:0] sel_974636;
  wire [7:0] add_974639;
  wire [7:0] sel_974640;
  wire [7:0] add_974643;
  wire [7:0] sel_974644;
  wire [7:0] add_974647;
  wire [7:0] sel_974648;
  wire [7:0] add_974651;
  wire [7:0] sel_974652;
  wire [7:0] add_974655;
  wire [7:0] sel_974656;
  wire [7:0] add_974659;
  wire [7:0] sel_974660;
  wire [7:0] add_974663;
  wire [7:0] sel_974664;
  wire [7:0] add_974667;
  wire [7:0] sel_974668;
  wire [7:0] add_974671;
  wire [7:0] sel_974672;
  wire [7:0] add_974675;
  wire [7:0] sel_974676;
  wire [7:0] add_974679;
  wire [7:0] sel_974680;
  wire [7:0] add_974683;
  wire [7:0] sel_974684;
  wire [7:0] add_974687;
  wire [7:0] sel_974688;
  wire [7:0] add_974691;
  wire [7:0] sel_974692;
  wire [7:0] add_974695;
  wire [7:0] sel_974696;
  wire [7:0] add_974699;
  wire [7:0] sel_974700;
  wire [7:0] add_974703;
  wire [7:0] sel_974704;
  wire [7:0] add_974707;
  wire [7:0] sel_974708;
  wire [7:0] add_974711;
  wire [7:0] sel_974712;
  wire [7:0] add_974715;
  wire [7:0] sel_974716;
  wire [7:0] add_974719;
  wire [7:0] sel_974720;
  wire [7:0] add_974723;
  wire [7:0] sel_974724;
  wire [7:0] add_974727;
  wire [7:0] sel_974728;
  wire [7:0] add_974731;
  wire [7:0] sel_974732;
  wire [7:0] add_974735;
  wire [7:0] sel_974736;
  wire [7:0] add_974739;
  wire [7:0] sel_974740;
  wire [7:0] add_974743;
  wire [7:0] sel_974744;
  wire [7:0] add_974747;
  wire [7:0] sel_974748;
  wire [7:0] add_974751;
  wire [7:0] sel_974752;
  wire [7:0] add_974755;
  wire [7:0] sel_974756;
  wire [7:0] add_974759;
  wire [7:0] sel_974760;
  wire [7:0] add_974763;
  wire [7:0] sel_974764;
  wire [7:0] add_974767;
  wire [7:0] sel_974768;
  wire [7:0] add_974771;
  wire [7:0] sel_974772;
  wire [7:0] add_974775;
  wire [7:0] sel_974776;
  wire [7:0] add_974779;
  wire [7:0] sel_974780;
  wire [7:0] add_974783;
  wire [7:0] sel_974784;
  wire [7:0] add_974787;
  wire [7:0] sel_974788;
  wire [7:0] add_974791;
  wire [7:0] sel_974792;
  wire [7:0] add_974795;
  wire [7:0] sel_974796;
  wire [7:0] add_974799;
  wire [7:0] sel_974800;
  wire [7:0] add_974803;
  wire [7:0] sel_974804;
  wire [7:0] add_974807;
  wire [7:0] sel_974808;
  wire [7:0] add_974811;
  wire [7:0] sel_974812;
  wire [7:0] add_974815;
  wire [7:0] sel_974816;
  wire [7:0] add_974820;
  wire [15:0] array_index_974821;
  wire [7:0] sel_974822;
  wire [7:0] add_974825;
  wire [7:0] sel_974826;
  wire [7:0] add_974829;
  wire [7:0] sel_974830;
  wire [7:0] add_974833;
  wire [7:0] sel_974834;
  wire [7:0] add_974837;
  wire [7:0] sel_974838;
  wire [7:0] add_974841;
  wire [7:0] sel_974842;
  wire [7:0] add_974845;
  wire [7:0] sel_974846;
  wire [7:0] add_974849;
  wire [7:0] sel_974850;
  wire [7:0] add_974853;
  wire [7:0] sel_974854;
  wire [7:0] add_974857;
  wire [7:0] sel_974858;
  wire [7:0] add_974861;
  wire [7:0] sel_974862;
  wire [7:0] add_974865;
  wire [7:0] sel_974866;
  wire [7:0] add_974869;
  wire [7:0] sel_974870;
  wire [7:0] add_974873;
  wire [7:0] sel_974874;
  wire [7:0] add_974877;
  wire [7:0] sel_974878;
  wire [7:0] add_974881;
  wire [7:0] sel_974882;
  wire [7:0] add_974885;
  wire [7:0] sel_974886;
  wire [7:0] add_974889;
  wire [7:0] sel_974890;
  wire [7:0] add_974893;
  wire [7:0] sel_974894;
  wire [7:0] add_974897;
  wire [7:0] sel_974898;
  wire [7:0] add_974901;
  wire [7:0] sel_974902;
  wire [7:0] add_974905;
  wire [7:0] sel_974906;
  wire [7:0] add_974909;
  wire [7:0] sel_974910;
  wire [7:0] add_974913;
  wire [7:0] sel_974914;
  wire [7:0] add_974917;
  wire [7:0] sel_974918;
  wire [7:0] add_974921;
  wire [7:0] sel_974922;
  wire [7:0] add_974925;
  wire [7:0] sel_974926;
  wire [7:0] add_974929;
  wire [7:0] sel_974930;
  wire [7:0] add_974933;
  wire [7:0] sel_974934;
  wire [7:0] add_974937;
  wire [7:0] sel_974938;
  wire [7:0] add_974941;
  wire [7:0] sel_974942;
  wire [7:0] add_974945;
  wire [7:0] sel_974946;
  wire [7:0] add_974949;
  wire [7:0] sel_974950;
  wire [7:0] add_974953;
  wire [7:0] sel_974954;
  wire [7:0] add_974957;
  wire [7:0] sel_974958;
  wire [7:0] add_974961;
  wire [7:0] sel_974962;
  wire [7:0] add_974965;
  wire [7:0] sel_974966;
  wire [7:0] add_974969;
  wire [7:0] sel_974970;
  wire [7:0] add_974973;
  wire [7:0] sel_974974;
  wire [7:0] add_974977;
  wire [7:0] sel_974978;
  wire [7:0] add_974981;
  wire [7:0] sel_974982;
  wire [7:0] add_974985;
  wire [7:0] sel_974986;
  wire [7:0] add_974989;
  wire [7:0] sel_974990;
  wire [7:0] add_974993;
  wire [7:0] sel_974994;
  wire [7:0] add_974997;
  wire [7:0] sel_974998;
  wire [7:0] add_975001;
  wire [7:0] sel_975002;
  wire [7:0] add_975005;
  wire [7:0] sel_975006;
  wire [7:0] add_975009;
  wire [7:0] sel_975010;
  wire [7:0] add_975013;
  wire [7:0] sel_975014;
  wire [7:0] add_975017;
  wire [7:0] sel_975018;
  wire [7:0] add_975021;
  wire [7:0] sel_975022;
  wire [7:0] add_975025;
  wire [7:0] sel_975026;
  wire [7:0] add_975029;
  wire [7:0] sel_975030;
  wire [7:0] add_975033;
  wire [7:0] sel_975034;
  wire [7:0] add_975037;
  wire [7:0] sel_975038;
  wire [7:0] add_975041;
  wire [7:0] sel_975042;
  wire [7:0] add_975045;
  wire [7:0] sel_975046;
  wire [7:0] add_975049;
  wire [7:0] sel_975050;
  wire [7:0] add_975053;
  wire [7:0] sel_975054;
  wire [7:0] add_975057;
  wire [7:0] sel_975058;
  wire [7:0] add_975061;
  wire [7:0] sel_975062;
  wire [7:0] add_975065;
  wire [7:0] sel_975066;
  wire [7:0] add_975069;
  wire [7:0] sel_975070;
  wire [7:0] add_975073;
  wire [7:0] sel_975074;
  wire [7:0] add_975077;
  wire [7:0] sel_975078;
  wire [7:0] add_975081;
  wire [7:0] sel_975082;
  wire [7:0] add_975085;
  wire [7:0] sel_975086;
  wire [7:0] add_975089;
  wire [7:0] sel_975090;
  wire [7:0] add_975093;
  wire [7:0] sel_975094;
  wire [7:0] add_975097;
  wire [7:0] sel_975098;
  wire [7:0] add_975101;
  wire [7:0] sel_975102;
  wire [7:0] add_975105;
  wire [7:0] sel_975106;
  wire [7:0] add_975109;
  wire [7:0] sel_975110;
  wire [7:0] add_975113;
  wire [7:0] sel_975114;
  wire [7:0] add_975117;
  wire [7:0] sel_975118;
  wire [7:0] add_975121;
  wire [7:0] sel_975122;
  wire [7:0] add_975125;
  wire [7:0] sel_975126;
  wire [7:0] add_975129;
  wire [7:0] sel_975130;
  wire [7:0] add_975133;
  wire [7:0] sel_975134;
  wire [7:0] add_975137;
  wire [7:0] sel_975138;
  wire [7:0] add_975141;
  wire [7:0] sel_975142;
  wire [7:0] add_975145;
  wire [7:0] sel_975146;
  wire [7:0] add_975149;
  wire [7:0] sel_975150;
  wire [7:0] add_975153;
  wire [7:0] sel_975154;
  wire [7:0] add_975157;
  wire [7:0] sel_975158;
  wire [7:0] add_975161;
  wire [7:0] sel_975162;
  wire [7:0] add_975165;
  wire [7:0] sel_975166;
  wire [7:0] add_975169;
  wire [7:0] sel_975170;
  wire [7:0] add_975173;
  wire [7:0] sel_975174;
  wire [7:0] add_975177;
  wire [7:0] sel_975178;
  wire [7:0] add_975181;
  wire [7:0] sel_975182;
  wire [7:0] add_975185;
  wire [7:0] sel_975186;
  wire [7:0] add_975189;
  wire [7:0] sel_975190;
  wire [7:0] add_975193;
  wire [7:0] sel_975194;
  wire [7:0] add_975197;
  wire [7:0] sel_975198;
  wire [7:0] add_975201;
  wire [7:0] sel_975202;
  wire [7:0] add_975205;
  wire [7:0] sel_975206;
  wire [7:0] add_975209;
  wire [7:0] sel_975210;
  wire [7:0] add_975213;
  wire [7:0] sel_975214;
  wire [7:0] add_975217;
  wire [7:0] sel_975218;
  wire [7:0] add_975222;
  wire [15:0] array_index_975223;
  wire [7:0] sel_975224;
  wire [7:0] add_975227;
  wire [7:0] sel_975228;
  wire [7:0] add_975231;
  wire [7:0] sel_975232;
  wire [7:0] add_975235;
  wire [7:0] sel_975236;
  wire [7:0] add_975239;
  wire [7:0] sel_975240;
  wire [7:0] add_975243;
  wire [7:0] sel_975244;
  wire [7:0] add_975247;
  wire [7:0] sel_975248;
  wire [7:0] add_975251;
  wire [7:0] sel_975252;
  wire [7:0] add_975255;
  wire [7:0] sel_975256;
  wire [7:0] add_975259;
  wire [7:0] sel_975260;
  wire [7:0] add_975263;
  wire [7:0] sel_975264;
  wire [7:0] add_975267;
  wire [7:0] sel_975268;
  wire [7:0] add_975271;
  wire [7:0] sel_975272;
  wire [7:0] add_975275;
  wire [7:0] sel_975276;
  wire [7:0] add_975279;
  wire [7:0] sel_975280;
  wire [7:0] add_975283;
  wire [7:0] sel_975284;
  wire [7:0] add_975287;
  wire [7:0] sel_975288;
  wire [7:0] add_975291;
  wire [7:0] sel_975292;
  wire [7:0] add_975295;
  wire [7:0] sel_975296;
  wire [7:0] add_975299;
  wire [7:0] sel_975300;
  wire [7:0] add_975303;
  wire [7:0] sel_975304;
  wire [7:0] add_975307;
  wire [7:0] sel_975308;
  wire [7:0] add_975311;
  wire [7:0] sel_975312;
  wire [7:0] add_975315;
  wire [7:0] sel_975316;
  wire [7:0] add_975319;
  wire [7:0] sel_975320;
  wire [7:0] add_975323;
  wire [7:0] sel_975324;
  wire [7:0] add_975327;
  wire [7:0] sel_975328;
  wire [7:0] add_975331;
  wire [7:0] sel_975332;
  wire [7:0] add_975335;
  wire [7:0] sel_975336;
  wire [7:0] add_975339;
  wire [7:0] sel_975340;
  wire [7:0] add_975343;
  wire [7:0] sel_975344;
  wire [7:0] add_975347;
  wire [7:0] sel_975348;
  wire [7:0] add_975351;
  wire [7:0] sel_975352;
  wire [7:0] add_975355;
  wire [7:0] sel_975356;
  wire [7:0] add_975359;
  wire [7:0] sel_975360;
  wire [7:0] add_975363;
  wire [7:0] sel_975364;
  wire [7:0] add_975367;
  wire [7:0] sel_975368;
  wire [7:0] add_975371;
  wire [7:0] sel_975372;
  wire [7:0] add_975375;
  wire [7:0] sel_975376;
  wire [7:0] add_975379;
  wire [7:0] sel_975380;
  wire [7:0] add_975383;
  wire [7:0] sel_975384;
  wire [7:0] add_975387;
  wire [7:0] sel_975388;
  wire [7:0] add_975391;
  wire [7:0] sel_975392;
  wire [7:0] add_975395;
  wire [7:0] sel_975396;
  wire [7:0] add_975399;
  wire [7:0] sel_975400;
  wire [7:0] add_975403;
  wire [7:0] sel_975404;
  wire [7:0] add_975407;
  wire [7:0] sel_975408;
  wire [7:0] add_975411;
  wire [7:0] sel_975412;
  wire [7:0] add_975415;
  wire [7:0] sel_975416;
  wire [7:0] add_975419;
  wire [7:0] sel_975420;
  wire [7:0] add_975423;
  wire [7:0] sel_975424;
  wire [7:0] add_975427;
  wire [7:0] sel_975428;
  wire [7:0] add_975431;
  wire [7:0] sel_975432;
  wire [7:0] add_975435;
  wire [7:0] sel_975436;
  wire [7:0] add_975439;
  wire [7:0] sel_975440;
  wire [7:0] add_975443;
  wire [7:0] sel_975444;
  wire [7:0] add_975447;
  wire [7:0] sel_975448;
  wire [7:0] add_975451;
  wire [7:0] sel_975452;
  wire [7:0] add_975455;
  wire [7:0] sel_975456;
  wire [7:0] add_975459;
  wire [7:0] sel_975460;
  wire [7:0] add_975463;
  wire [7:0] sel_975464;
  wire [7:0] add_975467;
  wire [7:0] sel_975468;
  wire [7:0] add_975471;
  wire [7:0] sel_975472;
  wire [7:0] add_975475;
  wire [7:0] sel_975476;
  wire [7:0] add_975479;
  wire [7:0] sel_975480;
  wire [7:0] add_975483;
  wire [7:0] sel_975484;
  wire [7:0] add_975487;
  wire [7:0] sel_975488;
  wire [7:0] add_975491;
  wire [7:0] sel_975492;
  wire [7:0] add_975495;
  wire [7:0] sel_975496;
  wire [7:0] add_975499;
  wire [7:0] sel_975500;
  wire [7:0] add_975503;
  wire [7:0] sel_975504;
  wire [7:0] add_975507;
  wire [7:0] sel_975508;
  wire [7:0] add_975511;
  wire [7:0] sel_975512;
  wire [7:0] add_975515;
  wire [7:0] sel_975516;
  wire [7:0] add_975519;
  wire [7:0] sel_975520;
  wire [7:0] add_975523;
  wire [7:0] sel_975524;
  wire [7:0] add_975527;
  wire [7:0] sel_975528;
  wire [7:0] add_975531;
  wire [7:0] sel_975532;
  wire [7:0] add_975535;
  wire [7:0] sel_975536;
  wire [7:0] add_975539;
  wire [7:0] sel_975540;
  wire [7:0] add_975543;
  wire [7:0] sel_975544;
  wire [7:0] add_975547;
  wire [7:0] sel_975548;
  wire [7:0] add_975551;
  wire [7:0] sel_975552;
  wire [7:0] add_975555;
  wire [7:0] sel_975556;
  wire [7:0] add_975559;
  wire [7:0] sel_975560;
  wire [7:0] add_975563;
  wire [7:0] sel_975564;
  wire [7:0] add_975567;
  wire [7:0] sel_975568;
  wire [7:0] add_975571;
  wire [7:0] sel_975572;
  wire [7:0] add_975575;
  wire [7:0] sel_975576;
  wire [7:0] add_975579;
  wire [7:0] sel_975580;
  wire [7:0] add_975583;
  wire [7:0] sel_975584;
  wire [7:0] add_975587;
  wire [7:0] sel_975588;
  wire [7:0] add_975591;
  wire [7:0] sel_975592;
  wire [7:0] add_975595;
  wire [7:0] sel_975596;
  wire [7:0] add_975599;
  wire [7:0] sel_975600;
  wire [7:0] add_975603;
  wire [7:0] sel_975604;
  wire [7:0] add_975607;
  wire [7:0] sel_975608;
  wire [7:0] add_975611;
  wire [7:0] sel_975612;
  wire [7:0] add_975615;
  wire [7:0] sel_975616;
  wire [7:0] add_975619;
  wire [7:0] sel_975620;
  wire [7:0] add_975624;
  wire [15:0] array_index_975625;
  wire [7:0] sel_975626;
  wire [7:0] add_975629;
  wire [7:0] sel_975630;
  wire [7:0] add_975633;
  wire [7:0] sel_975634;
  wire [7:0] add_975637;
  wire [7:0] sel_975638;
  wire [7:0] add_975641;
  wire [7:0] sel_975642;
  wire [7:0] add_975645;
  wire [7:0] sel_975646;
  wire [7:0] add_975649;
  wire [7:0] sel_975650;
  wire [7:0] add_975653;
  wire [7:0] sel_975654;
  wire [7:0] add_975657;
  wire [7:0] sel_975658;
  wire [7:0] add_975661;
  wire [7:0] sel_975662;
  wire [7:0] add_975665;
  wire [7:0] sel_975666;
  wire [7:0] add_975669;
  wire [7:0] sel_975670;
  wire [7:0] add_975673;
  wire [7:0] sel_975674;
  wire [7:0] add_975677;
  wire [7:0] sel_975678;
  wire [7:0] add_975681;
  wire [7:0] sel_975682;
  wire [7:0] add_975685;
  wire [7:0] sel_975686;
  wire [7:0] add_975689;
  wire [7:0] sel_975690;
  wire [7:0] add_975693;
  wire [7:0] sel_975694;
  wire [7:0] add_975697;
  wire [7:0] sel_975698;
  wire [7:0] add_975701;
  wire [7:0] sel_975702;
  wire [7:0] add_975705;
  wire [7:0] sel_975706;
  wire [7:0] add_975709;
  wire [7:0] sel_975710;
  wire [7:0] add_975713;
  wire [7:0] sel_975714;
  wire [7:0] add_975717;
  wire [7:0] sel_975718;
  wire [7:0] add_975721;
  wire [7:0] sel_975722;
  wire [7:0] add_975725;
  wire [7:0] sel_975726;
  wire [7:0] add_975729;
  wire [7:0] sel_975730;
  wire [7:0] add_975733;
  wire [7:0] sel_975734;
  wire [7:0] add_975737;
  wire [7:0] sel_975738;
  wire [7:0] add_975741;
  wire [7:0] sel_975742;
  wire [7:0] add_975745;
  wire [7:0] sel_975746;
  wire [7:0] add_975749;
  wire [7:0] sel_975750;
  wire [7:0] add_975753;
  wire [7:0] sel_975754;
  wire [7:0] add_975757;
  wire [7:0] sel_975758;
  wire [7:0] add_975761;
  wire [7:0] sel_975762;
  wire [7:0] add_975765;
  wire [7:0] sel_975766;
  wire [7:0] add_975769;
  wire [7:0] sel_975770;
  wire [7:0] add_975773;
  wire [7:0] sel_975774;
  wire [7:0] add_975777;
  wire [7:0] sel_975778;
  wire [7:0] add_975781;
  wire [7:0] sel_975782;
  wire [7:0] add_975785;
  wire [7:0] sel_975786;
  wire [7:0] add_975789;
  wire [7:0] sel_975790;
  wire [7:0] add_975793;
  wire [7:0] sel_975794;
  wire [7:0] add_975797;
  wire [7:0] sel_975798;
  wire [7:0] add_975801;
  wire [7:0] sel_975802;
  wire [7:0] add_975805;
  wire [7:0] sel_975806;
  wire [7:0] add_975809;
  wire [7:0] sel_975810;
  wire [7:0] add_975813;
  wire [7:0] sel_975814;
  wire [7:0] add_975817;
  wire [7:0] sel_975818;
  wire [7:0] add_975821;
  wire [7:0] sel_975822;
  wire [7:0] add_975825;
  wire [7:0] sel_975826;
  wire [7:0] add_975829;
  wire [7:0] sel_975830;
  wire [7:0] add_975833;
  wire [7:0] sel_975834;
  wire [7:0] add_975837;
  wire [7:0] sel_975838;
  wire [7:0] add_975841;
  wire [7:0] sel_975842;
  wire [7:0] add_975845;
  wire [7:0] sel_975846;
  wire [7:0] add_975849;
  wire [7:0] sel_975850;
  wire [7:0] add_975853;
  wire [7:0] sel_975854;
  wire [7:0] add_975857;
  wire [7:0] sel_975858;
  wire [7:0] add_975861;
  wire [7:0] sel_975862;
  wire [7:0] add_975865;
  wire [7:0] sel_975866;
  wire [7:0] add_975869;
  wire [7:0] sel_975870;
  wire [7:0] add_975873;
  wire [7:0] sel_975874;
  wire [7:0] add_975877;
  wire [7:0] sel_975878;
  wire [7:0] add_975881;
  wire [7:0] sel_975882;
  wire [7:0] add_975885;
  wire [7:0] sel_975886;
  wire [7:0] add_975889;
  wire [7:0] sel_975890;
  wire [7:0] add_975893;
  wire [7:0] sel_975894;
  wire [7:0] add_975897;
  wire [7:0] sel_975898;
  wire [7:0] add_975901;
  wire [7:0] sel_975902;
  wire [7:0] add_975905;
  wire [7:0] sel_975906;
  wire [7:0] add_975909;
  wire [7:0] sel_975910;
  wire [7:0] add_975913;
  wire [7:0] sel_975914;
  wire [7:0] add_975917;
  wire [7:0] sel_975918;
  wire [7:0] add_975921;
  wire [7:0] sel_975922;
  wire [7:0] add_975925;
  wire [7:0] sel_975926;
  wire [7:0] add_975929;
  wire [7:0] sel_975930;
  wire [7:0] add_975933;
  wire [7:0] sel_975934;
  wire [7:0] add_975937;
  wire [7:0] sel_975938;
  wire [7:0] add_975941;
  wire [7:0] sel_975942;
  wire [7:0] add_975945;
  wire [7:0] sel_975946;
  wire [7:0] add_975949;
  wire [7:0] sel_975950;
  wire [7:0] add_975953;
  wire [7:0] sel_975954;
  wire [7:0] add_975957;
  wire [7:0] sel_975958;
  wire [7:0] add_975961;
  wire [7:0] sel_975962;
  wire [7:0] add_975965;
  wire [7:0] sel_975966;
  wire [7:0] add_975969;
  wire [7:0] sel_975970;
  wire [7:0] add_975973;
  wire [7:0] sel_975974;
  wire [7:0] add_975977;
  wire [7:0] sel_975978;
  wire [7:0] add_975981;
  wire [7:0] sel_975982;
  wire [7:0] add_975985;
  wire [7:0] sel_975986;
  wire [7:0] add_975989;
  wire [7:0] sel_975990;
  wire [7:0] add_975993;
  wire [7:0] sel_975994;
  wire [7:0] add_975997;
  wire [7:0] sel_975998;
  wire [7:0] add_976001;
  wire [7:0] sel_976002;
  wire [7:0] add_976005;
  wire [7:0] sel_976006;
  wire [7:0] add_976009;
  wire [7:0] sel_976010;
  wire [7:0] add_976013;
  wire [7:0] sel_976014;
  wire [7:0] add_976017;
  wire [7:0] sel_976018;
  wire [7:0] add_976021;
  wire [7:0] sel_976022;
  wire [7:0] add_976026;
  wire [15:0] array_index_976027;
  wire [7:0] sel_976028;
  wire [7:0] add_976031;
  wire [7:0] sel_976032;
  wire [7:0] add_976035;
  wire [7:0] sel_976036;
  wire [7:0] add_976039;
  wire [7:0] sel_976040;
  wire [7:0] add_976043;
  wire [7:0] sel_976044;
  wire [7:0] add_976047;
  wire [7:0] sel_976048;
  wire [7:0] add_976051;
  wire [7:0] sel_976052;
  wire [7:0] add_976055;
  wire [7:0] sel_976056;
  wire [7:0] add_976059;
  wire [7:0] sel_976060;
  wire [7:0] add_976063;
  wire [7:0] sel_976064;
  wire [7:0] add_976067;
  wire [7:0] sel_976068;
  wire [7:0] add_976071;
  wire [7:0] sel_976072;
  wire [7:0] add_976075;
  wire [7:0] sel_976076;
  wire [7:0] add_976079;
  wire [7:0] sel_976080;
  wire [7:0] add_976083;
  wire [7:0] sel_976084;
  wire [7:0] add_976087;
  wire [7:0] sel_976088;
  wire [7:0] add_976091;
  wire [7:0] sel_976092;
  wire [7:0] add_976095;
  wire [7:0] sel_976096;
  wire [7:0] add_976099;
  wire [7:0] sel_976100;
  wire [7:0] add_976103;
  wire [7:0] sel_976104;
  wire [7:0] add_976107;
  wire [7:0] sel_976108;
  wire [7:0] add_976111;
  wire [7:0] sel_976112;
  wire [7:0] add_976115;
  wire [7:0] sel_976116;
  wire [7:0] add_976119;
  wire [7:0] sel_976120;
  wire [7:0] add_976123;
  wire [7:0] sel_976124;
  wire [7:0] add_976127;
  wire [7:0] sel_976128;
  wire [7:0] add_976131;
  wire [7:0] sel_976132;
  wire [7:0] add_976135;
  wire [7:0] sel_976136;
  wire [7:0] add_976139;
  wire [7:0] sel_976140;
  wire [7:0] add_976143;
  wire [7:0] sel_976144;
  wire [7:0] add_976147;
  wire [7:0] sel_976148;
  wire [7:0] add_976151;
  wire [7:0] sel_976152;
  wire [7:0] add_976155;
  wire [7:0] sel_976156;
  wire [7:0] add_976159;
  wire [7:0] sel_976160;
  wire [7:0] add_976163;
  wire [7:0] sel_976164;
  wire [7:0] add_976167;
  wire [7:0] sel_976168;
  wire [7:0] add_976171;
  wire [7:0] sel_976172;
  wire [7:0] add_976175;
  wire [7:0] sel_976176;
  wire [7:0] add_976179;
  wire [7:0] sel_976180;
  wire [7:0] add_976183;
  wire [7:0] sel_976184;
  wire [7:0] add_976187;
  wire [7:0] sel_976188;
  wire [7:0] add_976191;
  wire [7:0] sel_976192;
  wire [7:0] add_976195;
  wire [7:0] sel_976196;
  wire [7:0] add_976199;
  wire [7:0] sel_976200;
  wire [7:0] add_976203;
  wire [7:0] sel_976204;
  wire [7:0] add_976207;
  wire [7:0] sel_976208;
  wire [7:0] add_976211;
  wire [7:0] sel_976212;
  wire [7:0] add_976215;
  wire [7:0] sel_976216;
  wire [7:0] add_976219;
  wire [7:0] sel_976220;
  wire [7:0] add_976223;
  wire [7:0] sel_976224;
  wire [7:0] add_976227;
  wire [7:0] sel_976228;
  wire [7:0] add_976231;
  wire [7:0] sel_976232;
  wire [7:0] add_976235;
  wire [7:0] sel_976236;
  wire [7:0] add_976239;
  wire [7:0] sel_976240;
  wire [7:0] add_976243;
  wire [7:0] sel_976244;
  wire [7:0] add_976247;
  wire [7:0] sel_976248;
  wire [7:0] add_976251;
  wire [7:0] sel_976252;
  wire [7:0] add_976255;
  wire [7:0] sel_976256;
  wire [7:0] add_976259;
  wire [7:0] sel_976260;
  wire [7:0] add_976263;
  wire [7:0] sel_976264;
  wire [7:0] add_976267;
  wire [7:0] sel_976268;
  wire [7:0] add_976271;
  wire [7:0] sel_976272;
  wire [7:0] add_976275;
  wire [7:0] sel_976276;
  wire [7:0] add_976279;
  wire [7:0] sel_976280;
  wire [7:0] add_976283;
  wire [7:0] sel_976284;
  wire [7:0] add_976287;
  wire [7:0] sel_976288;
  wire [7:0] add_976291;
  wire [7:0] sel_976292;
  wire [7:0] add_976295;
  wire [7:0] sel_976296;
  wire [7:0] add_976299;
  wire [7:0] sel_976300;
  wire [7:0] add_976303;
  wire [7:0] sel_976304;
  wire [7:0] add_976307;
  wire [7:0] sel_976308;
  wire [7:0] add_976311;
  wire [7:0] sel_976312;
  wire [7:0] add_976315;
  wire [7:0] sel_976316;
  wire [7:0] add_976319;
  wire [7:0] sel_976320;
  wire [7:0] add_976323;
  wire [7:0] sel_976324;
  wire [7:0] add_976327;
  wire [7:0] sel_976328;
  wire [7:0] add_976331;
  wire [7:0] sel_976332;
  wire [7:0] add_976335;
  wire [7:0] sel_976336;
  wire [7:0] add_976339;
  wire [7:0] sel_976340;
  wire [7:0] add_976343;
  wire [7:0] sel_976344;
  wire [7:0] add_976347;
  wire [7:0] sel_976348;
  wire [7:0] add_976351;
  wire [7:0] sel_976352;
  wire [7:0] add_976355;
  wire [7:0] sel_976356;
  wire [7:0] add_976359;
  wire [7:0] sel_976360;
  wire [7:0] add_976363;
  wire [7:0] sel_976364;
  wire [7:0] add_976367;
  wire [7:0] sel_976368;
  wire [7:0] add_976371;
  wire [7:0] sel_976372;
  wire [7:0] add_976375;
  wire [7:0] sel_976376;
  wire [7:0] add_976379;
  wire [7:0] sel_976380;
  wire [7:0] add_976383;
  wire [7:0] sel_976384;
  wire [7:0] add_976387;
  wire [7:0] sel_976388;
  wire [7:0] add_976391;
  wire [7:0] sel_976392;
  wire [7:0] add_976395;
  wire [7:0] sel_976396;
  wire [7:0] add_976399;
  wire [7:0] sel_976400;
  wire [7:0] add_976403;
  wire [7:0] sel_976404;
  wire [7:0] add_976407;
  wire [7:0] sel_976408;
  wire [7:0] add_976411;
  wire [7:0] sel_976412;
  wire [7:0] add_976415;
  wire [7:0] sel_976416;
  wire [7:0] add_976419;
  wire [7:0] sel_976420;
  wire [7:0] add_976423;
  wire [7:0] sel_976424;
  wire [7:0] add_976428;
  wire [15:0] array_index_976429;
  wire [7:0] sel_976430;
  wire [7:0] add_976433;
  wire [7:0] sel_976434;
  wire [7:0] add_976437;
  wire [7:0] sel_976438;
  wire [7:0] add_976441;
  wire [7:0] sel_976442;
  wire [7:0] add_976445;
  wire [7:0] sel_976446;
  wire [7:0] add_976449;
  wire [7:0] sel_976450;
  wire [7:0] add_976453;
  wire [7:0] sel_976454;
  wire [7:0] add_976457;
  wire [7:0] sel_976458;
  wire [7:0] add_976461;
  wire [7:0] sel_976462;
  wire [7:0] add_976465;
  wire [7:0] sel_976466;
  wire [7:0] add_976469;
  wire [7:0] sel_976470;
  wire [7:0] add_976473;
  wire [7:0] sel_976474;
  wire [7:0] add_976477;
  wire [7:0] sel_976478;
  wire [7:0] add_976481;
  wire [7:0] sel_976482;
  wire [7:0] add_976485;
  wire [7:0] sel_976486;
  wire [7:0] add_976489;
  wire [7:0] sel_976490;
  wire [7:0] add_976493;
  wire [7:0] sel_976494;
  wire [7:0] add_976497;
  wire [7:0] sel_976498;
  wire [7:0] add_976501;
  wire [7:0] sel_976502;
  wire [7:0] add_976505;
  wire [7:0] sel_976506;
  wire [7:0] add_976509;
  wire [7:0] sel_976510;
  wire [7:0] add_976513;
  wire [7:0] sel_976514;
  wire [7:0] add_976517;
  wire [7:0] sel_976518;
  wire [7:0] add_976521;
  wire [7:0] sel_976522;
  wire [7:0] add_976525;
  wire [7:0] sel_976526;
  wire [7:0] add_976529;
  wire [7:0] sel_976530;
  wire [7:0] add_976533;
  wire [7:0] sel_976534;
  wire [7:0] add_976537;
  wire [7:0] sel_976538;
  wire [7:0] add_976541;
  wire [7:0] sel_976542;
  wire [7:0] add_976545;
  wire [7:0] sel_976546;
  wire [7:0] add_976549;
  wire [7:0] sel_976550;
  wire [7:0] add_976553;
  wire [7:0] sel_976554;
  wire [7:0] add_976557;
  wire [7:0] sel_976558;
  wire [7:0] add_976561;
  wire [7:0] sel_976562;
  wire [7:0] add_976565;
  wire [7:0] sel_976566;
  wire [7:0] add_976569;
  wire [7:0] sel_976570;
  wire [7:0] add_976573;
  wire [7:0] sel_976574;
  wire [7:0] add_976577;
  wire [7:0] sel_976578;
  wire [7:0] add_976581;
  wire [7:0] sel_976582;
  wire [7:0] add_976585;
  wire [7:0] sel_976586;
  wire [7:0] add_976589;
  wire [7:0] sel_976590;
  wire [7:0] add_976593;
  wire [7:0] sel_976594;
  wire [7:0] add_976597;
  wire [7:0] sel_976598;
  wire [7:0] add_976601;
  wire [7:0] sel_976602;
  wire [7:0] add_976605;
  wire [7:0] sel_976606;
  wire [7:0] add_976609;
  wire [7:0] sel_976610;
  wire [7:0] add_976613;
  wire [7:0] sel_976614;
  wire [7:0] add_976617;
  wire [7:0] sel_976618;
  wire [7:0] add_976621;
  wire [7:0] sel_976622;
  wire [7:0] add_976625;
  wire [7:0] sel_976626;
  wire [7:0] add_976629;
  wire [7:0] sel_976630;
  wire [7:0] add_976633;
  wire [7:0] sel_976634;
  wire [7:0] add_976637;
  wire [7:0] sel_976638;
  wire [7:0] add_976641;
  wire [7:0] sel_976642;
  wire [7:0] add_976645;
  wire [7:0] sel_976646;
  wire [7:0] add_976649;
  wire [7:0] sel_976650;
  wire [7:0] add_976653;
  wire [7:0] sel_976654;
  wire [7:0] add_976657;
  wire [7:0] sel_976658;
  wire [7:0] add_976661;
  wire [7:0] sel_976662;
  wire [7:0] add_976665;
  wire [7:0] sel_976666;
  wire [7:0] add_976669;
  wire [7:0] sel_976670;
  wire [7:0] add_976673;
  wire [7:0] sel_976674;
  wire [7:0] add_976677;
  wire [7:0] sel_976678;
  wire [7:0] add_976681;
  wire [7:0] sel_976682;
  wire [7:0] add_976685;
  wire [7:0] sel_976686;
  wire [7:0] add_976689;
  wire [7:0] sel_976690;
  wire [7:0] add_976693;
  wire [7:0] sel_976694;
  wire [7:0] add_976697;
  wire [7:0] sel_976698;
  wire [7:0] add_976701;
  wire [7:0] sel_976702;
  wire [7:0] add_976705;
  wire [7:0] sel_976706;
  wire [7:0] add_976709;
  wire [7:0] sel_976710;
  wire [7:0] add_976713;
  wire [7:0] sel_976714;
  wire [7:0] add_976717;
  wire [7:0] sel_976718;
  wire [7:0] add_976721;
  wire [7:0] sel_976722;
  wire [7:0] add_976725;
  wire [7:0] sel_976726;
  wire [7:0] add_976729;
  wire [7:0] sel_976730;
  wire [7:0] add_976733;
  wire [7:0] sel_976734;
  wire [7:0] add_976737;
  wire [7:0] sel_976738;
  wire [7:0] add_976741;
  wire [7:0] sel_976742;
  wire [7:0] add_976745;
  wire [7:0] sel_976746;
  wire [7:0] add_976749;
  wire [7:0] sel_976750;
  wire [7:0] add_976753;
  wire [7:0] sel_976754;
  wire [7:0] add_976757;
  wire [7:0] sel_976758;
  wire [7:0] add_976761;
  wire [7:0] sel_976762;
  wire [7:0] add_976765;
  wire [7:0] sel_976766;
  wire [7:0] add_976769;
  wire [7:0] sel_976770;
  wire [7:0] add_976773;
  wire [7:0] sel_976774;
  wire [7:0] add_976777;
  wire [7:0] sel_976778;
  wire [7:0] add_976781;
  wire [7:0] sel_976782;
  wire [7:0] add_976785;
  wire [7:0] sel_976786;
  wire [7:0] add_976789;
  wire [7:0] sel_976790;
  wire [7:0] add_976793;
  wire [7:0] sel_976794;
  wire [7:0] add_976797;
  wire [7:0] sel_976798;
  wire [7:0] add_976801;
  wire [7:0] sel_976802;
  wire [7:0] add_976805;
  wire [7:0] sel_976806;
  wire [7:0] add_976809;
  wire [7:0] sel_976810;
  wire [7:0] add_976813;
  wire [7:0] sel_976814;
  wire [7:0] add_976817;
  wire [7:0] sel_976818;
  wire [7:0] add_976821;
  wire [7:0] sel_976822;
  wire [7:0] add_976825;
  wire [7:0] sel_976826;
  wire [7:0] add_976830;
  wire [15:0] array_index_976831;
  wire [7:0] sel_976832;
  wire [7:0] add_976835;
  wire [7:0] sel_976836;
  wire [7:0] add_976839;
  wire [7:0] sel_976840;
  wire [7:0] add_976843;
  wire [7:0] sel_976844;
  wire [7:0] add_976847;
  wire [7:0] sel_976848;
  wire [7:0] add_976851;
  wire [7:0] sel_976852;
  wire [7:0] add_976855;
  wire [7:0] sel_976856;
  wire [7:0] add_976859;
  wire [7:0] sel_976860;
  wire [7:0] add_976863;
  wire [7:0] sel_976864;
  wire [7:0] add_976867;
  wire [7:0] sel_976868;
  wire [7:0] add_976871;
  wire [7:0] sel_976872;
  wire [7:0] add_976875;
  wire [7:0] sel_976876;
  wire [7:0] add_976879;
  wire [7:0] sel_976880;
  wire [7:0] add_976883;
  wire [7:0] sel_976884;
  wire [7:0] add_976887;
  wire [7:0] sel_976888;
  wire [7:0] add_976891;
  wire [7:0] sel_976892;
  wire [7:0] add_976895;
  wire [7:0] sel_976896;
  wire [7:0] add_976899;
  wire [7:0] sel_976900;
  wire [7:0] add_976903;
  wire [7:0] sel_976904;
  wire [7:0] add_976907;
  wire [7:0] sel_976908;
  wire [7:0] add_976911;
  wire [7:0] sel_976912;
  wire [7:0] add_976915;
  wire [7:0] sel_976916;
  wire [7:0] add_976919;
  wire [7:0] sel_976920;
  wire [7:0] add_976923;
  wire [7:0] sel_976924;
  wire [7:0] add_976927;
  wire [7:0] sel_976928;
  wire [7:0] add_976931;
  wire [7:0] sel_976932;
  wire [7:0] add_976935;
  wire [7:0] sel_976936;
  wire [7:0] add_976939;
  wire [7:0] sel_976940;
  wire [7:0] add_976943;
  wire [7:0] sel_976944;
  wire [7:0] add_976947;
  wire [7:0] sel_976948;
  wire [7:0] add_976951;
  wire [7:0] sel_976952;
  wire [7:0] add_976955;
  wire [7:0] sel_976956;
  wire [7:0] add_976959;
  wire [7:0] sel_976960;
  wire [7:0] add_976963;
  wire [7:0] sel_976964;
  wire [7:0] add_976967;
  wire [7:0] sel_976968;
  wire [7:0] add_976971;
  wire [7:0] sel_976972;
  wire [7:0] add_976975;
  wire [7:0] sel_976976;
  wire [7:0] add_976979;
  wire [7:0] sel_976980;
  wire [7:0] add_976983;
  wire [7:0] sel_976984;
  wire [7:0] add_976987;
  wire [7:0] sel_976988;
  wire [7:0] add_976991;
  wire [7:0] sel_976992;
  wire [7:0] add_976995;
  wire [7:0] sel_976996;
  wire [7:0] add_976999;
  wire [7:0] sel_977000;
  wire [7:0] add_977003;
  wire [7:0] sel_977004;
  wire [7:0] add_977007;
  wire [7:0] sel_977008;
  wire [7:0] add_977011;
  wire [7:0] sel_977012;
  wire [7:0] add_977015;
  wire [7:0] sel_977016;
  wire [7:0] add_977019;
  wire [7:0] sel_977020;
  wire [7:0] add_977023;
  wire [7:0] sel_977024;
  wire [7:0] add_977027;
  wire [7:0] sel_977028;
  wire [7:0] add_977031;
  wire [7:0] sel_977032;
  wire [7:0] add_977035;
  wire [7:0] sel_977036;
  wire [7:0] add_977039;
  wire [7:0] sel_977040;
  wire [7:0] add_977043;
  wire [7:0] sel_977044;
  wire [7:0] add_977047;
  wire [7:0] sel_977048;
  wire [7:0] add_977051;
  wire [7:0] sel_977052;
  wire [7:0] add_977055;
  wire [7:0] sel_977056;
  wire [7:0] add_977059;
  wire [7:0] sel_977060;
  wire [7:0] add_977063;
  wire [7:0] sel_977064;
  wire [7:0] add_977067;
  wire [7:0] sel_977068;
  wire [7:0] add_977071;
  wire [7:0] sel_977072;
  wire [7:0] add_977075;
  wire [7:0] sel_977076;
  wire [7:0] add_977079;
  wire [7:0] sel_977080;
  wire [7:0] add_977083;
  wire [7:0] sel_977084;
  wire [7:0] add_977087;
  wire [7:0] sel_977088;
  wire [7:0] add_977091;
  wire [7:0] sel_977092;
  wire [7:0] add_977095;
  wire [7:0] sel_977096;
  wire [7:0] add_977099;
  wire [7:0] sel_977100;
  wire [7:0] add_977103;
  wire [7:0] sel_977104;
  wire [7:0] add_977107;
  wire [7:0] sel_977108;
  wire [7:0] add_977111;
  wire [7:0] sel_977112;
  wire [7:0] add_977115;
  wire [7:0] sel_977116;
  wire [7:0] add_977119;
  wire [7:0] sel_977120;
  wire [7:0] add_977123;
  wire [7:0] sel_977124;
  wire [7:0] add_977127;
  wire [7:0] sel_977128;
  wire [7:0] add_977131;
  wire [7:0] sel_977132;
  wire [7:0] add_977135;
  wire [7:0] sel_977136;
  wire [7:0] add_977139;
  wire [7:0] sel_977140;
  wire [7:0] add_977143;
  wire [7:0] sel_977144;
  wire [7:0] add_977147;
  wire [7:0] sel_977148;
  wire [7:0] add_977151;
  wire [7:0] sel_977152;
  wire [7:0] add_977155;
  wire [7:0] sel_977156;
  wire [7:0] add_977159;
  wire [7:0] sel_977160;
  wire [7:0] add_977163;
  wire [7:0] sel_977164;
  wire [7:0] add_977167;
  wire [7:0] sel_977168;
  wire [7:0] add_977171;
  wire [7:0] sel_977172;
  wire [7:0] add_977175;
  wire [7:0] sel_977176;
  wire [7:0] add_977179;
  wire [7:0] sel_977180;
  wire [7:0] add_977183;
  wire [7:0] sel_977184;
  wire [7:0] add_977187;
  wire [7:0] sel_977188;
  wire [7:0] add_977191;
  wire [7:0] sel_977192;
  wire [7:0] add_977195;
  wire [7:0] sel_977196;
  wire [7:0] add_977199;
  wire [7:0] sel_977200;
  wire [7:0] add_977203;
  wire [7:0] sel_977204;
  wire [7:0] add_977207;
  wire [7:0] sel_977208;
  wire [7:0] add_977211;
  wire [7:0] sel_977212;
  wire [7:0] add_977215;
  wire [7:0] sel_977216;
  wire [7:0] add_977219;
  wire [7:0] sel_977220;
  wire [7:0] add_977223;
  wire [7:0] sel_977224;
  wire [7:0] add_977227;
  wire [7:0] sel_977228;
  wire [7:0] add_977232;
  wire [15:0] array_index_977233;
  wire [7:0] sel_977234;
  wire [7:0] add_977237;
  wire [7:0] sel_977238;
  wire [7:0] add_977241;
  wire [7:0] sel_977242;
  wire [7:0] add_977245;
  wire [7:0] sel_977246;
  wire [7:0] add_977249;
  wire [7:0] sel_977250;
  wire [7:0] add_977253;
  wire [7:0] sel_977254;
  wire [7:0] add_977257;
  wire [7:0] sel_977258;
  wire [7:0] add_977261;
  wire [7:0] sel_977262;
  wire [7:0] add_977265;
  wire [7:0] sel_977266;
  wire [7:0] add_977269;
  wire [7:0] sel_977270;
  wire [7:0] add_977273;
  wire [7:0] sel_977274;
  wire [7:0] add_977277;
  wire [7:0] sel_977278;
  wire [7:0] add_977281;
  wire [7:0] sel_977282;
  wire [7:0] add_977285;
  wire [7:0] sel_977286;
  wire [7:0] add_977289;
  wire [7:0] sel_977290;
  wire [7:0] add_977293;
  wire [7:0] sel_977294;
  wire [7:0] add_977297;
  wire [7:0] sel_977298;
  wire [7:0] add_977301;
  wire [7:0] sel_977302;
  wire [7:0] add_977305;
  wire [7:0] sel_977306;
  wire [7:0] add_977309;
  wire [7:0] sel_977310;
  wire [7:0] add_977313;
  wire [7:0] sel_977314;
  wire [7:0] add_977317;
  wire [7:0] sel_977318;
  wire [7:0] add_977321;
  wire [7:0] sel_977322;
  wire [7:0] add_977325;
  wire [7:0] sel_977326;
  wire [7:0] add_977329;
  wire [7:0] sel_977330;
  wire [7:0] add_977333;
  wire [7:0] sel_977334;
  wire [7:0] add_977337;
  wire [7:0] sel_977338;
  wire [7:0] add_977341;
  wire [7:0] sel_977342;
  wire [7:0] add_977345;
  wire [7:0] sel_977346;
  wire [7:0] add_977349;
  wire [7:0] sel_977350;
  wire [7:0] add_977353;
  wire [7:0] sel_977354;
  wire [7:0] add_977357;
  wire [7:0] sel_977358;
  wire [7:0] add_977361;
  wire [7:0] sel_977362;
  wire [7:0] add_977365;
  wire [7:0] sel_977366;
  wire [7:0] add_977369;
  wire [7:0] sel_977370;
  wire [7:0] add_977373;
  wire [7:0] sel_977374;
  wire [7:0] add_977377;
  wire [7:0] sel_977378;
  wire [7:0] add_977381;
  wire [7:0] sel_977382;
  wire [7:0] add_977385;
  wire [7:0] sel_977386;
  wire [7:0] add_977389;
  wire [7:0] sel_977390;
  wire [7:0] add_977393;
  wire [7:0] sel_977394;
  wire [7:0] add_977397;
  wire [7:0] sel_977398;
  wire [7:0] add_977401;
  wire [7:0] sel_977402;
  wire [7:0] add_977405;
  wire [7:0] sel_977406;
  wire [7:0] add_977409;
  wire [7:0] sel_977410;
  wire [7:0] add_977413;
  wire [7:0] sel_977414;
  wire [7:0] add_977417;
  wire [7:0] sel_977418;
  wire [7:0] add_977421;
  wire [7:0] sel_977422;
  wire [7:0] add_977425;
  wire [7:0] sel_977426;
  wire [7:0] add_977429;
  wire [7:0] sel_977430;
  wire [7:0] add_977433;
  wire [7:0] sel_977434;
  wire [7:0] add_977437;
  wire [7:0] sel_977438;
  wire [7:0] add_977441;
  wire [7:0] sel_977442;
  wire [7:0] add_977445;
  wire [7:0] sel_977446;
  wire [7:0] add_977449;
  wire [7:0] sel_977450;
  wire [7:0] add_977453;
  wire [7:0] sel_977454;
  wire [7:0] add_977457;
  wire [7:0] sel_977458;
  wire [7:0] add_977461;
  wire [7:0] sel_977462;
  wire [7:0] add_977465;
  wire [7:0] sel_977466;
  wire [7:0] add_977469;
  wire [7:0] sel_977470;
  wire [7:0] add_977473;
  wire [7:0] sel_977474;
  wire [7:0] add_977477;
  wire [7:0] sel_977478;
  wire [7:0] add_977481;
  wire [7:0] sel_977482;
  wire [7:0] add_977485;
  wire [7:0] sel_977486;
  wire [7:0] add_977489;
  wire [7:0] sel_977490;
  wire [7:0] add_977493;
  wire [7:0] sel_977494;
  wire [7:0] add_977497;
  wire [7:0] sel_977498;
  wire [7:0] add_977501;
  wire [7:0] sel_977502;
  wire [7:0] add_977505;
  wire [7:0] sel_977506;
  wire [7:0] add_977509;
  wire [7:0] sel_977510;
  wire [7:0] add_977513;
  wire [7:0] sel_977514;
  wire [7:0] add_977517;
  wire [7:0] sel_977518;
  wire [7:0] add_977521;
  wire [7:0] sel_977522;
  wire [7:0] add_977525;
  wire [7:0] sel_977526;
  wire [7:0] add_977529;
  wire [7:0] sel_977530;
  wire [7:0] add_977533;
  wire [7:0] sel_977534;
  wire [7:0] add_977537;
  wire [7:0] sel_977538;
  wire [7:0] add_977541;
  wire [7:0] sel_977542;
  wire [7:0] add_977545;
  wire [7:0] sel_977546;
  wire [7:0] add_977549;
  wire [7:0] sel_977550;
  wire [7:0] add_977553;
  wire [7:0] sel_977554;
  wire [7:0] add_977557;
  wire [7:0] sel_977558;
  wire [7:0] add_977561;
  wire [7:0] sel_977562;
  wire [7:0] add_977565;
  wire [7:0] sel_977566;
  wire [7:0] add_977569;
  wire [7:0] sel_977570;
  wire [7:0] add_977573;
  wire [7:0] sel_977574;
  wire [7:0] add_977577;
  wire [7:0] sel_977578;
  wire [7:0] add_977581;
  wire [7:0] sel_977582;
  wire [7:0] add_977585;
  wire [7:0] sel_977586;
  wire [7:0] add_977589;
  wire [7:0] sel_977590;
  wire [7:0] add_977593;
  wire [7:0] sel_977594;
  wire [7:0] add_977597;
  wire [7:0] sel_977598;
  wire [7:0] add_977601;
  wire [7:0] sel_977602;
  wire [7:0] add_977605;
  wire [7:0] sel_977606;
  wire [7:0] add_977609;
  wire [7:0] sel_977610;
  wire [7:0] add_977613;
  wire [7:0] sel_977614;
  wire [7:0] add_977617;
  wire [7:0] sel_977618;
  wire [7:0] add_977621;
  wire [7:0] sel_977622;
  wire [7:0] add_977625;
  wire [7:0] sel_977626;
  wire [7:0] add_977629;
  wire [7:0] sel_977630;
  wire [7:0] add_977634;
  wire [15:0] array_index_977635;
  wire [7:0] sel_977636;
  wire [7:0] add_977639;
  wire [7:0] sel_977640;
  wire [7:0] add_977643;
  wire [7:0] sel_977644;
  wire [7:0] add_977647;
  wire [7:0] sel_977648;
  wire [7:0] add_977651;
  wire [7:0] sel_977652;
  wire [7:0] add_977655;
  wire [7:0] sel_977656;
  wire [7:0] add_977659;
  wire [7:0] sel_977660;
  wire [7:0] add_977663;
  wire [7:0] sel_977664;
  wire [7:0] add_977667;
  wire [7:0] sel_977668;
  wire [7:0] add_977671;
  wire [7:0] sel_977672;
  wire [7:0] add_977675;
  wire [7:0] sel_977676;
  wire [7:0] add_977679;
  wire [7:0] sel_977680;
  wire [7:0] add_977683;
  wire [7:0] sel_977684;
  wire [7:0] add_977687;
  wire [7:0] sel_977688;
  wire [7:0] add_977691;
  wire [7:0] sel_977692;
  wire [7:0] add_977695;
  wire [7:0] sel_977696;
  wire [7:0] add_977699;
  wire [7:0] sel_977700;
  wire [7:0] add_977703;
  wire [7:0] sel_977704;
  wire [7:0] add_977707;
  wire [7:0] sel_977708;
  wire [7:0] add_977711;
  wire [7:0] sel_977712;
  wire [7:0] add_977715;
  wire [7:0] sel_977716;
  wire [7:0] add_977719;
  wire [7:0] sel_977720;
  wire [7:0] add_977723;
  wire [7:0] sel_977724;
  wire [7:0] add_977727;
  wire [7:0] sel_977728;
  wire [7:0] add_977731;
  wire [7:0] sel_977732;
  wire [7:0] add_977735;
  wire [7:0] sel_977736;
  wire [7:0] add_977739;
  wire [7:0] sel_977740;
  wire [7:0] add_977743;
  wire [7:0] sel_977744;
  wire [7:0] add_977747;
  wire [7:0] sel_977748;
  wire [7:0] add_977751;
  wire [7:0] sel_977752;
  wire [7:0] add_977755;
  wire [7:0] sel_977756;
  wire [7:0] add_977759;
  wire [7:0] sel_977760;
  wire [7:0] add_977763;
  wire [7:0] sel_977764;
  wire [7:0] add_977767;
  wire [7:0] sel_977768;
  wire [7:0] add_977771;
  wire [7:0] sel_977772;
  wire [7:0] add_977775;
  wire [7:0] sel_977776;
  wire [7:0] add_977779;
  wire [7:0] sel_977780;
  wire [7:0] add_977783;
  wire [7:0] sel_977784;
  wire [7:0] add_977787;
  wire [7:0] sel_977788;
  wire [7:0] add_977791;
  wire [7:0] sel_977792;
  wire [7:0] add_977795;
  wire [7:0] sel_977796;
  wire [7:0] add_977799;
  wire [7:0] sel_977800;
  wire [7:0] add_977803;
  wire [7:0] sel_977804;
  wire [7:0] add_977807;
  wire [7:0] sel_977808;
  wire [7:0] add_977811;
  wire [7:0] sel_977812;
  wire [7:0] add_977815;
  wire [7:0] sel_977816;
  wire [7:0] add_977819;
  wire [7:0] sel_977820;
  wire [7:0] add_977823;
  wire [7:0] sel_977824;
  wire [7:0] add_977827;
  wire [7:0] sel_977828;
  wire [7:0] add_977831;
  wire [7:0] sel_977832;
  wire [7:0] add_977835;
  wire [7:0] sel_977836;
  wire [7:0] add_977839;
  wire [7:0] sel_977840;
  wire [7:0] add_977843;
  wire [7:0] sel_977844;
  wire [7:0] add_977847;
  wire [7:0] sel_977848;
  wire [7:0] add_977851;
  wire [7:0] sel_977852;
  wire [7:0] add_977855;
  wire [7:0] sel_977856;
  wire [7:0] add_977859;
  wire [7:0] sel_977860;
  wire [7:0] add_977863;
  wire [7:0] sel_977864;
  wire [7:0] add_977867;
  wire [7:0] sel_977868;
  wire [7:0] add_977871;
  wire [7:0] sel_977872;
  wire [7:0] add_977875;
  wire [7:0] sel_977876;
  wire [7:0] add_977879;
  wire [7:0] sel_977880;
  wire [7:0] add_977883;
  wire [7:0] sel_977884;
  wire [7:0] add_977887;
  wire [7:0] sel_977888;
  wire [7:0] add_977891;
  wire [7:0] sel_977892;
  wire [7:0] add_977895;
  wire [7:0] sel_977896;
  wire [7:0] add_977899;
  wire [7:0] sel_977900;
  wire [7:0] add_977903;
  wire [7:0] sel_977904;
  wire [7:0] add_977907;
  wire [7:0] sel_977908;
  wire [7:0] add_977911;
  wire [7:0] sel_977912;
  wire [7:0] add_977915;
  wire [7:0] sel_977916;
  wire [7:0] add_977919;
  wire [7:0] sel_977920;
  wire [7:0] add_977923;
  wire [7:0] sel_977924;
  wire [7:0] add_977927;
  wire [7:0] sel_977928;
  wire [7:0] add_977931;
  wire [7:0] sel_977932;
  wire [7:0] add_977935;
  wire [7:0] sel_977936;
  wire [7:0] add_977939;
  wire [7:0] sel_977940;
  wire [7:0] add_977943;
  wire [7:0] sel_977944;
  wire [7:0] add_977947;
  wire [7:0] sel_977948;
  wire [7:0] add_977951;
  wire [7:0] sel_977952;
  wire [7:0] add_977955;
  wire [7:0] sel_977956;
  wire [7:0] add_977959;
  wire [7:0] sel_977960;
  wire [7:0] add_977963;
  wire [7:0] sel_977964;
  wire [7:0] add_977967;
  wire [7:0] sel_977968;
  wire [7:0] add_977971;
  wire [7:0] sel_977972;
  wire [7:0] add_977975;
  wire [7:0] sel_977976;
  wire [7:0] add_977979;
  wire [7:0] sel_977980;
  wire [7:0] add_977983;
  wire [7:0] sel_977984;
  wire [7:0] add_977987;
  wire [7:0] sel_977988;
  wire [7:0] add_977991;
  wire [7:0] sel_977992;
  wire [7:0] add_977995;
  wire [7:0] sel_977996;
  wire [7:0] add_977999;
  wire [7:0] sel_978000;
  wire [7:0] add_978003;
  wire [7:0] sel_978004;
  wire [7:0] add_978007;
  wire [7:0] sel_978008;
  wire [7:0] add_978011;
  wire [7:0] sel_978012;
  wire [7:0] add_978015;
  wire [7:0] sel_978016;
  wire [7:0] add_978019;
  wire [7:0] sel_978020;
  wire [7:0] add_978023;
  wire [7:0] sel_978024;
  wire [7:0] add_978027;
  wire [7:0] sel_978028;
  wire [7:0] add_978031;
  wire [7:0] sel_978032;
  wire [7:0] add_978036;
  wire [15:0] array_index_978037;
  wire [7:0] sel_978038;
  wire [7:0] add_978041;
  wire [7:0] sel_978042;
  wire [7:0] add_978045;
  wire [7:0] sel_978046;
  wire [7:0] add_978049;
  wire [7:0] sel_978050;
  wire [7:0] add_978053;
  wire [7:0] sel_978054;
  wire [7:0] add_978057;
  wire [7:0] sel_978058;
  wire [7:0] add_978061;
  wire [7:0] sel_978062;
  wire [7:0] add_978065;
  wire [7:0] sel_978066;
  wire [7:0] add_978069;
  wire [7:0] sel_978070;
  wire [7:0] add_978073;
  wire [7:0] sel_978074;
  wire [7:0] add_978077;
  wire [7:0] sel_978078;
  wire [7:0] add_978081;
  wire [7:0] sel_978082;
  wire [7:0] add_978085;
  wire [7:0] sel_978086;
  wire [7:0] add_978089;
  wire [7:0] sel_978090;
  wire [7:0] add_978093;
  wire [7:0] sel_978094;
  wire [7:0] add_978097;
  wire [7:0] sel_978098;
  wire [7:0] add_978101;
  wire [7:0] sel_978102;
  wire [7:0] add_978105;
  wire [7:0] sel_978106;
  wire [7:0] add_978109;
  wire [7:0] sel_978110;
  wire [7:0] add_978113;
  wire [7:0] sel_978114;
  wire [7:0] add_978117;
  wire [7:0] sel_978118;
  wire [7:0] add_978121;
  wire [7:0] sel_978122;
  wire [7:0] add_978125;
  wire [7:0] sel_978126;
  wire [7:0] add_978129;
  wire [7:0] sel_978130;
  wire [7:0] add_978133;
  wire [7:0] sel_978134;
  wire [7:0] add_978137;
  wire [7:0] sel_978138;
  wire [7:0] add_978141;
  wire [7:0] sel_978142;
  wire [7:0] add_978145;
  wire [7:0] sel_978146;
  wire [7:0] add_978149;
  wire [7:0] sel_978150;
  wire [7:0] add_978153;
  wire [7:0] sel_978154;
  wire [7:0] add_978157;
  wire [7:0] sel_978158;
  wire [7:0] add_978161;
  wire [7:0] sel_978162;
  wire [7:0] add_978165;
  wire [7:0] sel_978166;
  wire [7:0] add_978169;
  wire [7:0] sel_978170;
  wire [7:0] add_978173;
  wire [7:0] sel_978174;
  wire [7:0] add_978177;
  wire [7:0] sel_978178;
  wire [7:0] add_978181;
  wire [7:0] sel_978182;
  wire [7:0] add_978185;
  wire [7:0] sel_978186;
  wire [7:0] add_978189;
  wire [7:0] sel_978190;
  wire [7:0] add_978193;
  wire [7:0] sel_978194;
  wire [7:0] add_978197;
  wire [7:0] sel_978198;
  wire [7:0] add_978201;
  wire [7:0] sel_978202;
  wire [7:0] add_978205;
  wire [7:0] sel_978206;
  wire [7:0] add_978209;
  wire [7:0] sel_978210;
  wire [7:0] add_978213;
  wire [7:0] sel_978214;
  wire [7:0] add_978217;
  wire [7:0] sel_978218;
  wire [7:0] add_978221;
  wire [7:0] sel_978222;
  wire [7:0] add_978225;
  wire [7:0] sel_978226;
  wire [7:0] add_978229;
  wire [7:0] sel_978230;
  wire [7:0] add_978233;
  wire [7:0] sel_978234;
  wire [7:0] add_978237;
  wire [7:0] sel_978238;
  wire [7:0] add_978241;
  wire [7:0] sel_978242;
  wire [7:0] add_978245;
  wire [7:0] sel_978246;
  wire [7:0] add_978249;
  wire [7:0] sel_978250;
  wire [7:0] add_978253;
  wire [7:0] sel_978254;
  wire [7:0] add_978257;
  wire [7:0] sel_978258;
  wire [7:0] add_978261;
  wire [7:0] sel_978262;
  wire [7:0] add_978265;
  wire [7:0] sel_978266;
  wire [7:0] add_978269;
  wire [7:0] sel_978270;
  wire [7:0] add_978273;
  wire [7:0] sel_978274;
  wire [7:0] add_978277;
  wire [7:0] sel_978278;
  wire [7:0] add_978281;
  wire [7:0] sel_978282;
  wire [7:0] add_978285;
  wire [7:0] sel_978286;
  wire [7:0] add_978289;
  wire [7:0] sel_978290;
  wire [7:0] add_978293;
  wire [7:0] sel_978294;
  wire [7:0] add_978297;
  wire [7:0] sel_978298;
  wire [7:0] add_978301;
  wire [7:0] sel_978302;
  wire [7:0] add_978305;
  wire [7:0] sel_978306;
  wire [7:0] add_978309;
  wire [7:0] sel_978310;
  wire [7:0] add_978313;
  wire [7:0] sel_978314;
  wire [7:0] add_978317;
  wire [7:0] sel_978318;
  wire [7:0] add_978321;
  wire [7:0] sel_978322;
  wire [7:0] add_978325;
  wire [7:0] sel_978326;
  wire [7:0] add_978329;
  wire [7:0] sel_978330;
  wire [7:0] add_978333;
  wire [7:0] sel_978334;
  wire [7:0] add_978337;
  wire [7:0] sel_978338;
  wire [7:0] add_978341;
  wire [7:0] sel_978342;
  wire [7:0] add_978345;
  wire [7:0] sel_978346;
  wire [7:0] add_978349;
  wire [7:0] sel_978350;
  wire [7:0] add_978353;
  wire [7:0] sel_978354;
  wire [7:0] add_978357;
  wire [7:0] sel_978358;
  wire [7:0] add_978361;
  wire [7:0] sel_978362;
  wire [7:0] add_978365;
  wire [7:0] sel_978366;
  wire [7:0] add_978369;
  wire [7:0] sel_978370;
  wire [7:0] add_978373;
  wire [7:0] sel_978374;
  wire [7:0] add_978377;
  wire [7:0] sel_978378;
  wire [7:0] add_978381;
  wire [7:0] sel_978382;
  wire [7:0] add_978385;
  wire [7:0] sel_978386;
  wire [7:0] add_978389;
  wire [7:0] sel_978390;
  wire [7:0] add_978393;
  wire [7:0] sel_978394;
  wire [7:0] add_978397;
  wire [7:0] sel_978398;
  wire [7:0] add_978401;
  wire [7:0] sel_978402;
  wire [7:0] add_978405;
  wire [7:0] sel_978406;
  wire [7:0] add_978409;
  wire [7:0] sel_978410;
  wire [7:0] add_978413;
  wire [7:0] sel_978414;
  wire [7:0] add_978417;
  wire [7:0] sel_978418;
  wire [7:0] add_978421;
  wire [7:0] sel_978422;
  wire [7:0] add_978425;
  wire [7:0] sel_978426;
  wire [7:0] add_978429;
  wire [7:0] sel_978430;
  wire [7:0] add_978433;
  wire [7:0] sel_978434;
  wire [7:0] add_978438;
  wire [15:0] array_index_978439;
  wire [7:0] sel_978440;
  wire [7:0] add_978443;
  wire [7:0] sel_978444;
  wire [7:0] add_978447;
  wire [7:0] sel_978448;
  wire [7:0] add_978451;
  wire [7:0] sel_978452;
  wire [7:0] add_978455;
  wire [7:0] sel_978456;
  wire [7:0] add_978459;
  wire [7:0] sel_978460;
  wire [7:0] add_978463;
  wire [7:0] sel_978464;
  wire [7:0] add_978467;
  wire [7:0] sel_978468;
  wire [7:0] add_978471;
  wire [7:0] sel_978472;
  wire [7:0] add_978475;
  wire [7:0] sel_978476;
  wire [7:0] add_978479;
  wire [7:0] sel_978480;
  wire [7:0] add_978483;
  wire [7:0] sel_978484;
  wire [7:0] add_978487;
  wire [7:0] sel_978488;
  wire [7:0] add_978491;
  wire [7:0] sel_978492;
  wire [7:0] add_978495;
  wire [7:0] sel_978496;
  wire [7:0] add_978499;
  wire [7:0] sel_978500;
  wire [7:0] add_978503;
  wire [7:0] sel_978504;
  wire [7:0] add_978507;
  wire [7:0] sel_978508;
  wire [7:0] add_978511;
  wire [7:0] sel_978512;
  wire [7:0] add_978515;
  wire [7:0] sel_978516;
  wire [7:0] add_978519;
  wire [7:0] sel_978520;
  wire [7:0] add_978523;
  wire [7:0] sel_978524;
  wire [7:0] add_978527;
  wire [7:0] sel_978528;
  wire [7:0] add_978531;
  wire [7:0] sel_978532;
  wire [7:0] add_978535;
  wire [7:0] sel_978536;
  wire [7:0] add_978539;
  wire [7:0] sel_978540;
  wire [7:0] add_978543;
  wire [7:0] sel_978544;
  wire [7:0] add_978547;
  wire [7:0] sel_978548;
  wire [7:0] add_978551;
  wire [7:0] sel_978552;
  wire [7:0] add_978555;
  wire [7:0] sel_978556;
  wire [7:0] add_978559;
  wire [7:0] sel_978560;
  wire [7:0] add_978563;
  wire [7:0] sel_978564;
  wire [7:0] add_978567;
  wire [7:0] sel_978568;
  wire [7:0] add_978571;
  wire [7:0] sel_978572;
  wire [7:0] add_978575;
  wire [7:0] sel_978576;
  wire [7:0] add_978579;
  wire [7:0] sel_978580;
  wire [7:0] add_978583;
  wire [7:0] sel_978584;
  wire [7:0] add_978587;
  wire [7:0] sel_978588;
  wire [7:0] add_978591;
  wire [7:0] sel_978592;
  wire [7:0] add_978595;
  wire [7:0] sel_978596;
  wire [7:0] add_978599;
  wire [7:0] sel_978600;
  wire [7:0] add_978603;
  wire [7:0] sel_978604;
  wire [7:0] add_978607;
  wire [7:0] sel_978608;
  wire [7:0] add_978611;
  wire [7:0] sel_978612;
  wire [7:0] add_978615;
  wire [7:0] sel_978616;
  wire [7:0] add_978619;
  wire [7:0] sel_978620;
  wire [7:0] add_978623;
  wire [7:0] sel_978624;
  wire [7:0] add_978627;
  wire [7:0] sel_978628;
  wire [7:0] add_978631;
  wire [7:0] sel_978632;
  wire [7:0] add_978635;
  wire [7:0] sel_978636;
  wire [7:0] add_978639;
  wire [7:0] sel_978640;
  wire [7:0] add_978643;
  wire [7:0] sel_978644;
  wire [7:0] add_978647;
  wire [7:0] sel_978648;
  wire [7:0] add_978651;
  wire [7:0] sel_978652;
  wire [7:0] add_978655;
  wire [7:0] sel_978656;
  wire [7:0] add_978659;
  wire [7:0] sel_978660;
  wire [7:0] add_978663;
  wire [7:0] sel_978664;
  wire [7:0] add_978667;
  wire [7:0] sel_978668;
  wire [7:0] add_978671;
  wire [7:0] sel_978672;
  wire [7:0] add_978675;
  wire [7:0] sel_978676;
  wire [7:0] add_978679;
  wire [7:0] sel_978680;
  wire [7:0] add_978683;
  wire [7:0] sel_978684;
  wire [7:0] add_978687;
  wire [7:0] sel_978688;
  wire [7:0] add_978691;
  wire [7:0] sel_978692;
  wire [7:0] add_978695;
  wire [7:0] sel_978696;
  wire [7:0] add_978699;
  wire [7:0] sel_978700;
  wire [7:0] add_978703;
  wire [7:0] sel_978704;
  wire [7:0] add_978707;
  wire [7:0] sel_978708;
  wire [7:0] add_978711;
  wire [7:0] sel_978712;
  wire [7:0] add_978715;
  wire [7:0] sel_978716;
  wire [7:0] add_978719;
  wire [7:0] sel_978720;
  wire [7:0] add_978723;
  wire [7:0] sel_978724;
  wire [7:0] add_978727;
  wire [7:0] sel_978728;
  wire [7:0] add_978731;
  wire [7:0] sel_978732;
  wire [7:0] add_978735;
  wire [7:0] sel_978736;
  wire [7:0] add_978739;
  wire [7:0] sel_978740;
  wire [7:0] add_978743;
  wire [7:0] sel_978744;
  wire [7:0] add_978747;
  wire [7:0] sel_978748;
  wire [7:0] add_978751;
  wire [7:0] sel_978752;
  wire [7:0] add_978755;
  wire [7:0] sel_978756;
  wire [7:0] add_978759;
  wire [7:0] sel_978760;
  wire [7:0] add_978763;
  wire [7:0] sel_978764;
  wire [7:0] add_978767;
  wire [7:0] sel_978768;
  wire [7:0] add_978771;
  wire [7:0] sel_978772;
  wire [7:0] add_978775;
  wire [7:0] sel_978776;
  wire [7:0] add_978779;
  wire [7:0] sel_978780;
  wire [7:0] add_978783;
  wire [7:0] sel_978784;
  wire [7:0] add_978787;
  wire [7:0] sel_978788;
  wire [7:0] add_978791;
  wire [7:0] sel_978792;
  wire [7:0] add_978795;
  wire [7:0] sel_978796;
  wire [7:0] add_978799;
  wire [7:0] sel_978800;
  wire [7:0] add_978803;
  wire [7:0] sel_978804;
  wire [7:0] add_978807;
  wire [7:0] sel_978808;
  wire [7:0] add_978811;
  wire [7:0] sel_978812;
  wire [7:0] add_978815;
  wire [7:0] sel_978816;
  wire [7:0] add_978819;
  wire [7:0] sel_978820;
  wire [7:0] add_978823;
  wire [7:0] sel_978824;
  wire [7:0] add_978827;
  wire [7:0] sel_978828;
  wire [7:0] add_978831;
  wire [7:0] sel_978832;
  wire [7:0] add_978835;
  wire [7:0] sel_978836;
  wire [7:0] add_978840;
  wire [15:0] array_index_978841;
  wire [7:0] sel_978842;
  wire [7:0] add_978845;
  wire [7:0] sel_978846;
  wire [7:0] add_978849;
  wire [7:0] sel_978850;
  wire [7:0] add_978853;
  wire [7:0] sel_978854;
  wire [7:0] add_978857;
  wire [7:0] sel_978858;
  wire [7:0] add_978861;
  wire [7:0] sel_978862;
  wire [7:0] add_978865;
  wire [7:0] sel_978866;
  wire [7:0] add_978869;
  wire [7:0] sel_978870;
  wire [7:0] add_978873;
  wire [7:0] sel_978874;
  wire [7:0] add_978877;
  wire [7:0] sel_978878;
  wire [7:0] add_978881;
  wire [7:0] sel_978882;
  wire [7:0] add_978885;
  wire [7:0] sel_978886;
  wire [7:0] add_978889;
  wire [7:0] sel_978890;
  wire [7:0] add_978893;
  wire [7:0] sel_978894;
  wire [7:0] add_978897;
  wire [7:0] sel_978898;
  wire [7:0] add_978901;
  wire [7:0] sel_978902;
  wire [7:0] add_978905;
  wire [7:0] sel_978906;
  wire [7:0] add_978909;
  wire [7:0] sel_978910;
  wire [7:0] add_978913;
  wire [7:0] sel_978914;
  wire [7:0] add_978917;
  wire [7:0] sel_978918;
  wire [7:0] add_978921;
  wire [7:0] sel_978922;
  wire [7:0] add_978925;
  wire [7:0] sel_978926;
  wire [7:0] add_978929;
  wire [7:0] sel_978930;
  wire [7:0] add_978933;
  wire [7:0] sel_978934;
  wire [7:0] add_978937;
  wire [7:0] sel_978938;
  wire [7:0] add_978941;
  wire [7:0] sel_978942;
  wire [7:0] add_978945;
  wire [7:0] sel_978946;
  wire [7:0] add_978949;
  wire [7:0] sel_978950;
  wire [7:0] add_978953;
  wire [7:0] sel_978954;
  wire [7:0] add_978957;
  wire [7:0] sel_978958;
  wire [7:0] add_978961;
  wire [7:0] sel_978962;
  wire [7:0] add_978965;
  wire [7:0] sel_978966;
  wire [7:0] add_978969;
  wire [7:0] sel_978970;
  wire [7:0] add_978973;
  wire [7:0] sel_978974;
  wire [7:0] add_978977;
  wire [7:0] sel_978978;
  wire [7:0] add_978981;
  wire [7:0] sel_978982;
  wire [7:0] add_978985;
  wire [7:0] sel_978986;
  wire [7:0] add_978989;
  wire [7:0] sel_978990;
  wire [7:0] add_978993;
  wire [7:0] sel_978994;
  wire [7:0] add_978997;
  wire [7:0] sel_978998;
  wire [7:0] add_979001;
  wire [7:0] sel_979002;
  wire [7:0] add_979005;
  wire [7:0] sel_979006;
  wire [7:0] add_979009;
  wire [7:0] sel_979010;
  wire [7:0] add_979013;
  wire [7:0] sel_979014;
  wire [7:0] add_979017;
  wire [7:0] sel_979018;
  wire [7:0] add_979021;
  wire [7:0] sel_979022;
  wire [7:0] add_979025;
  wire [7:0] sel_979026;
  wire [7:0] add_979029;
  wire [7:0] sel_979030;
  wire [7:0] add_979033;
  wire [7:0] sel_979034;
  wire [7:0] add_979037;
  wire [7:0] sel_979038;
  wire [7:0] add_979041;
  wire [7:0] sel_979042;
  wire [7:0] add_979045;
  wire [7:0] sel_979046;
  wire [7:0] add_979049;
  wire [7:0] sel_979050;
  wire [7:0] add_979053;
  wire [7:0] sel_979054;
  wire [7:0] add_979057;
  wire [7:0] sel_979058;
  wire [7:0] add_979061;
  wire [7:0] sel_979062;
  wire [7:0] add_979065;
  wire [7:0] sel_979066;
  wire [7:0] add_979069;
  wire [7:0] sel_979070;
  wire [7:0] add_979073;
  wire [7:0] sel_979074;
  wire [7:0] add_979077;
  wire [7:0] sel_979078;
  wire [7:0] add_979081;
  wire [7:0] sel_979082;
  wire [7:0] add_979085;
  wire [7:0] sel_979086;
  wire [7:0] add_979089;
  wire [7:0] sel_979090;
  wire [7:0] add_979093;
  wire [7:0] sel_979094;
  wire [7:0] add_979097;
  wire [7:0] sel_979098;
  wire [7:0] add_979101;
  wire [7:0] sel_979102;
  wire [7:0] add_979105;
  wire [7:0] sel_979106;
  wire [7:0] add_979109;
  wire [7:0] sel_979110;
  wire [7:0] add_979113;
  wire [7:0] sel_979114;
  wire [7:0] add_979117;
  wire [7:0] sel_979118;
  wire [7:0] add_979121;
  wire [7:0] sel_979122;
  wire [7:0] add_979125;
  wire [7:0] sel_979126;
  wire [7:0] add_979129;
  wire [7:0] sel_979130;
  wire [7:0] add_979133;
  wire [7:0] sel_979134;
  wire [7:0] add_979137;
  wire [7:0] sel_979138;
  wire [7:0] add_979141;
  wire [7:0] sel_979142;
  wire [7:0] add_979145;
  wire [7:0] sel_979146;
  wire [7:0] add_979149;
  wire [7:0] sel_979150;
  wire [7:0] add_979153;
  wire [7:0] sel_979154;
  wire [7:0] add_979157;
  wire [7:0] sel_979158;
  wire [7:0] add_979161;
  wire [7:0] sel_979162;
  wire [7:0] add_979165;
  wire [7:0] sel_979166;
  wire [7:0] add_979169;
  wire [7:0] sel_979170;
  wire [7:0] add_979173;
  wire [7:0] sel_979174;
  wire [7:0] add_979177;
  wire [7:0] sel_979178;
  wire [7:0] add_979181;
  wire [7:0] sel_979182;
  wire [7:0] add_979185;
  wire [7:0] sel_979186;
  wire [7:0] add_979189;
  wire [7:0] sel_979190;
  wire [7:0] add_979193;
  wire [7:0] sel_979194;
  wire [7:0] add_979197;
  wire [7:0] sel_979198;
  wire [7:0] add_979201;
  wire [7:0] sel_979202;
  wire [7:0] add_979205;
  wire [7:0] sel_979206;
  wire [7:0] add_979209;
  wire [7:0] sel_979210;
  wire [7:0] add_979213;
  wire [7:0] sel_979214;
  wire [7:0] add_979217;
  wire [7:0] sel_979218;
  wire [7:0] add_979221;
  wire [7:0] sel_979222;
  wire [7:0] add_979225;
  wire [7:0] sel_979226;
  wire [7:0] add_979229;
  wire [7:0] sel_979230;
  wire [7:0] add_979233;
  wire [7:0] sel_979234;
  wire [7:0] add_979237;
  wire [7:0] sel_979238;
  wire [7:0] add_979242;
  wire [15:0] array_index_979243;
  wire [7:0] sel_979244;
  wire [7:0] add_979247;
  wire [7:0] sel_979248;
  wire [7:0] add_979251;
  wire [7:0] sel_979252;
  wire [7:0] add_979255;
  wire [7:0] sel_979256;
  wire [7:0] add_979259;
  wire [7:0] sel_979260;
  wire [7:0] add_979263;
  wire [7:0] sel_979264;
  wire [7:0] add_979267;
  wire [7:0] sel_979268;
  wire [7:0] add_979271;
  wire [7:0] sel_979272;
  wire [7:0] add_979275;
  wire [7:0] sel_979276;
  wire [7:0] add_979279;
  wire [7:0] sel_979280;
  wire [7:0] add_979283;
  wire [7:0] sel_979284;
  wire [7:0] add_979287;
  wire [7:0] sel_979288;
  wire [7:0] add_979291;
  wire [7:0] sel_979292;
  wire [7:0] add_979295;
  wire [7:0] sel_979296;
  wire [7:0] add_979299;
  wire [7:0] sel_979300;
  wire [7:0] add_979303;
  wire [7:0] sel_979304;
  wire [7:0] add_979307;
  wire [7:0] sel_979308;
  wire [7:0] add_979311;
  wire [7:0] sel_979312;
  wire [7:0] add_979315;
  wire [7:0] sel_979316;
  wire [7:0] add_979319;
  wire [7:0] sel_979320;
  wire [7:0] add_979323;
  wire [7:0] sel_979324;
  wire [7:0] add_979327;
  wire [7:0] sel_979328;
  wire [7:0] add_979331;
  wire [7:0] sel_979332;
  wire [7:0] add_979335;
  wire [7:0] sel_979336;
  wire [7:0] add_979339;
  wire [7:0] sel_979340;
  wire [7:0] add_979343;
  wire [7:0] sel_979344;
  wire [7:0] add_979347;
  wire [7:0] sel_979348;
  wire [7:0] add_979351;
  wire [7:0] sel_979352;
  wire [7:0] add_979355;
  wire [7:0] sel_979356;
  wire [7:0] add_979359;
  wire [7:0] sel_979360;
  wire [7:0] add_979363;
  wire [7:0] sel_979364;
  wire [7:0] add_979367;
  wire [7:0] sel_979368;
  wire [7:0] add_979371;
  wire [7:0] sel_979372;
  wire [7:0] add_979375;
  wire [7:0] sel_979376;
  wire [7:0] add_979379;
  wire [7:0] sel_979380;
  wire [7:0] add_979383;
  wire [7:0] sel_979384;
  wire [7:0] add_979387;
  wire [7:0] sel_979388;
  wire [7:0] add_979391;
  wire [7:0] sel_979392;
  wire [7:0] add_979395;
  wire [7:0] sel_979396;
  wire [7:0] add_979399;
  wire [7:0] sel_979400;
  wire [7:0] add_979403;
  wire [7:0] sel_979404;
  wire [7:0] add_979407;
  wire [7:0] sel_979408;
  wire [7:0] add_979411;
  wire [7:0] sel_979412;
  wire [7:0] add_979415;
  wire [7:0] sel_979416;
  wire [7:0] add_979419;
  wire [7:0] sel_979420;
  wire [7:0] add_979423;
  wire [7:0] sel_979424;
  wire [7:0] add_979427;
  wire [7:0] sel_979428;
  wire [7:0] add_979431;
  wire [7:0] sel_979432;
  wire [7:0] add_979435;
  wire [7:0] sel_979436;
  wire [7:0] add_979439;
  wire [7:0] sel_979440;
  wire [7:0] add_979443;
  wire [7:0] sel_979444;
  wire [7:0] add_979447;
  wire [7:0] sel_979448;
  wire [7:0] add_979451;
  wire [7:0] sel_979452;
  wire [7:0] add_979455;
  wire [7:0] sel_979456;
  wire [7:0] add_979459;
  wire [7:0] sel_979460;
  wire [7:0] add_979463;
  wire [7:0] sel_979464;
  wire [7:0] add_979467;
  wire [7:0] sel_979468;
  wire [7:0] add_979471;
  wire [7:0] sel_979472;
  wire [7:0] add_979475;
  wire [7:0] sel_979476;
  wire [7:0] add_979479;
  wire [7:0] sel_979480;
  wire [7:0] add_979483;
  wire [7:0] sel_979484;
  wire [7:0] add_979487;
  wire [7:0] sel_979488;
  wire [7:0] add_979491;
  wire [7:0] sel_979492;
  wire [7:0] add_979495;
  wire [7:0] sel_979496;
  wire [7:0] add_979499;
  wire [7:0] sel_979500;
  wire [7:0] add_979503;
  wire [7:0] sel_979504;
  wire [7:0] add_979507;
  wire [7:0] sel_979508;
  wire [7:0] add_979511;
  wire [7:0] sel_979512;
  wire [7:0] add_979515;
  wire [7:0] sel_979516;
  wire [7:0] add_979519;
  wire [7:0] sel_979520;
  wire [7:0] add_979523;
  wire [7:0] sel_979524;
  wire [7:0] add_979527;
  wire [7:0] sel_979528;
  wire [7:0] add_979531;
  wire [7:0] sel_979532;
  wire [7:0] add_979535;
  wire [7:0] sel_979536;
  wire [7:0] add_979539;
  wire [7:0] sel_979540;
  wire [7:0] add_979543;
  wire [7:0] sel_979544;
  wire [7:0] add_979547;
  wire [7:0] sel_979548;
  wire [7:0] add_979551;
  wire [7:0] sel_979552;
  wire [7:0] add_979555;
  wire [7:0] sel_979556;
  wire [7:0] add_979559;
  wire [7:0] sel_979560;
  wire [7:0] add_979563;
  wire [7:0] sel_979564;
  wire [7:0] add_979567;
  wire [7:0] sel_979568;
  wire [7:0] add_979571;
  wire [7:0] sel_979572;
  wire [7:0] add_979575;
  wire [7:0] sel_979576;
  wire [7:0] add_979579;
  wire [7:0] sel_979580;
  wire [7:0] add_979583;
  wire [7:0] sel_979584;
  wire [7:0] add_979587;
  wire [7:0] sel_979588;
  wire [7:0] add_979591;
  wire [7:0] sel_979592;
  wire [7:0] add_979595;
  wire [7:0] sel_979596;
  wire [7:0] add_979599;
  wire [7:0] sel_979600;
  wire [7:0] add_979603;
  wire [7:0] sel_979604;
  wire [7:0] add_979607;
  wire [7:0] sel_979608;
  wire [7:0] add_979611;
  wire [7:0] sel_979612;
  wire [7:0] add_979615;
  wire [7:0] sel_979616;
  wire [7:0] add_979619;
  wire [7:0] sel_979620;
  wire [7:0] add_979623;
  wire [7:0] sel_979624;
  wire [7:0] add_979627;
  wire [7:0] sel_979628;
  wire [7:0] add_979631;
  wire [7:0] sel_979632;
  wire [7:0] add_979635;
  wire [7:0] sel_979636;
  wire [7:0] add_979639;
  wire [7:0] sel_979640;
  wire [7:0] add_979644;
  wire [15:0] array_index_979645;
  wire [7:0] sel_979646;
  wire [7:0] add_979649;
  wire [7:0] sel_979650;
  wire [7:0] add_979653;
  wire [7:0] sel_979654;
  wire [7:0] add_979657;
  wire [7:0] sel_979658;
  wire [7:0] add_979661;
  wire [7:0] sel_979662;
  wire [7:0] add_979665;
  wire [7:0] sel_979666;
  wire [7:0] add_979669;
  wire [7:0] sel_979670;
  wire [7:0] add_979673;
  wire [7:0] sel_979674;
  wire [7:0] add_979677;
  wire [7:0] sel_979678;
  wire [7:0] add_979681;
  wire [7:0] sel_979682;
  wire [7:0] add_979685;
  wire [7:0] sel_979686;
  wire [7:0] add_979689;
  wire [7:0] sel_979690;
  wire [7:0] add_979693;
  wire [7:0] sel_979694;
  wire [7:0] add_979697;
  wire [7:0] sel_979698;
  wire [7:0] add_979701;
  wire [7:0] sel_979702;
  wire [7:0] add_979705;
  wire [7:0] sel_979706;
  wire [7:0] add_979709;
  wire [7:0] sel_979710;
  wire [7:0] add_979713;
  wire [7:0] sel_979714;
  wire [7:0] add_979717;
  wire [7:0] sel_979718;
  wire [7:0] add_979721;
  wire [7:0] sel_979722;
  wire [7:0] add_979725;
  wire [7:0] sel_979726;
  wire [7:0] add_979729;
  wire [7:0] sel_979730;
  wire [7:0] add_979733;
  wire [7:0] sel_979734;
  wire [7:0] add_979737;
  wire [7:0] sel_979738;
  wire [7:0] add_979741;
  wire [7:0] sel_979742;
  wire [7:0] add_979745;
  wire [7:0] sel_979746;
  wire [7:0] add_979749;
  wire [7:0] sel_979750;
  wire [7:0] add_979753;
  wire [7:0] sel_979754;
  wire [7:0] add_979757;
  wire [7:0] sel_979758;
  wire [7:0] add_979761;
  wire [7:0] sel_979762;
  wire [7:0] add_979765;
  wire [7:0] sel_979766;
  wire [7:0] add_979769;
  wire [7:0] sel_979770;
  wire [7:0] add_979773;
  wire [7:0] sel_979774;
  wire [7:0] add_979777;
  wire [7:0] sel_979778;
  wire [7:0] add_979781;
  wire [7:0] sel_979782;
  wire [7:0] add_979785;
  wire [7:0] sel_979786;
  wire [7:0] add_979789;
  wire [7:0] sel_979790;
  wire [7:0] add_979793;
  wire [7:0] sel_979794;
  wire [7:0] add_979797;
  wire [7:0] sel_979798;
  wire [7:0] add_979801;
  wire [7:0] sel_979802;
  wire [7:0] add_979805;
  wire [7:0] sel_979806;
  wire [7:0] add_979809;
  wire [7:0] sel_979810;
  wire [7:0] add_979813;
  wire [7:0] sel_979814;
  wire [7:0] add_979817;
  wire [7:0] sel_979818;
  wire [7:0] add_979821;
  wire [7:0] sel_979822;
  wire [7:0] add_979825;
  wire [7:0] sel_979826;
  wire [7:0] add_979829;
  wire [7:0] sel_979830;
  wire [7:0] add_979833;
  wire [7:0] sel_979834;
  wire [7:0] add_979837;
  wire [7:0] sel_979838;
  wire [7:0] add_979841;
  wire [7:0] sel_979842;
  wire [7:0] add_979845;
  wire [7:0] sel_979846;
  wire [7:0] add_979849;
  wire [7:0] sel_979850;
  wire [7:0] add_979853;
  wire [7:0] sel_979854;
  wire [7:0] add_979857;
  wire [7:0] sel_979858;
  wire [7:0] add_979861;
  wire [7:0] sel_979862;
  wire [7:0] add_979865;
  wire [7:0] sel_979866;
  wire [7:0] add_979869;
  wire [7:0] sel_979870;
  wire [7:0] add_979873;
  wire [7:0] sel_979874;
  wire [7:0] add_979877;
  wire [7:0] sel_979878;
  wire [7:0] add_979881;
  wire [7:0] sel_979882;
  wire [7:0] add_979885;
  wire [7:0] sel_979886;
  wire [7:0] add_979889;
  wire [7:0] sel_979890;
  wire [7:0] add_979893;
  wire [7:0] sel_979894;
  wire [7:0] add_979897;
  wire [7:0] sel_979898;
  wire [7:0] add_979901;
  wire [7:0] sel_979902;
  wire [7:0] add_979905;
  wire [7:0] sel_979906;
  wire [7:0] add_979909;
  wire [7:0] sel_979910;
  wire [7:0] add_979913;
  wire [7:0] sel_979914;
  wire [7:0] add_979917;
  wire [7:0] sel_979918;
  wire [7:0] add_979921;
  wire [7:0] sel_979922;
  wire [7:0] add_979925;
  wire [7:0] sel_979926;
  wire [7:0] add_979929;
  wire [7:0] sel_979930;
  wire [7:0] add_979933;
  wire [7:0] sel_979934;
  wire [7:0] add_979937;
  wire [7:0] sel_979938;
  wire [7:0] add_979941;
  wire [7:0] sel_979942;
  wire [7:0] add_979945;
  wire [7:0] sel_979946;
  wire [7:0] add_979949;
  wire [7:0] sel_979950;
  wire [7:0] add_979953;
  wire [7:0] sel_979954;
  wire [7:0] add_979957;
  wire [7:0] sel_979958;
  wire [7:0] add_979961;
  wire [7:0] sel_979962;
  wire [7:0] add_979965;
  wire [7:0] sel_979966;
  wire [7:0] add_979969;
  wire [7:0] sel_979970;
  wire [7:0] add_979973;
  wire [7:0] sel_979974;
  wire [7:0] add_979977;
  wire [7:0] sel_979978;
  wire [7:0] add_979981;
  wire [7:0] sel_979982;
  wire [7:0] add_979985;
  wire [7:0] sel_979986;
  wire [7:0] add_979989;
  wire [7:0] sel_979990;
  wire [7:0] add_979993;
  wire [7:0] sel_979994;
  wire [7:0] add_979997;
  wire [7:0] sel_979998;
  wire [7:0] add_980001;
  wire [7:0] sel_980002;
  wire [7:0] add_980005;
  wire [7:0] sel_980006;
  wire [7:0] add_980009;
  wire [7:0] sel_980010;
  wire [7:0] add_980013;
  wire [7:0] sel_980014;
  wire [7:0] add_980017;
  wire [7:0] sel_980018;
  wire [7:0] add_980021;
  wire [7:0] sel_980022;
  wire [7:0] add_980025;
  wire [7:0] sel_980026;
  wire [7:0] add_980029;
  wire [7:0] sel_980030;
  wire [7:0] add_980033;
  wire [7:0] sel_980034;
  wire [7:0] add_980037;
  wire [7:0] sel_980038;
  wire [7:0] add_980041;
  wire [7:0] sel_980042;
  wire [7:0] add_980046;
  wire [15:0] array_index_980047;
  wire [7:0] sel_980048;
  wire [7:0] add_980051;
  wire [7:0] sel_980052;
  wire [7:0] add_980055;
  wire [7:0] sel_980056;
  wire [7:0] add_980059;
  wire [7:0] sel_980060;
  wire [7:0] add_980063;
  wire [7:0] sel_980064;
  wire [7:0] add_980067;
  wire [7:0] sel_980068;
  wire [7:0] add_980071;
  wire [7:0] sel_980072;
  wire [7:0] add_980075;
  wire [7:0] sel_980076;
  wire [7:0] add_980079;
  wire [7:0] sel_980080;
  wire [7:0] add_980083;
  wire [7:0] sel_980084;
  wire [7:0] add_980087;
  wire [7:0] sel_980088;
  wire [7:0] add_980091;
  wire [7:0] sel_980092;
  wire [7:0] add_980095;
  wire [7:0] sel_980096;
  wire [7:0] add_980099;
  wire [7:0] sel_980100;
  wire [7:0] add_980103;
  wire [7:0] sel_980104;
  wire [7:0] add_980107;
  wire [7:0] sel_980108;
  wire [7:0] add_980111;
  wire [7:0] sel_980112;
  wire [7:0] add_980115;
  wire [7:0] sel_980116;
  wire [7:0] add_980119;
  wire [7:0] sel_980120;
  wire [7:0] add_980123;
  wire [7:0] sel_980124;
  wire [7:0] add_980127;
  wire [7:0] sel_980128;
  wire [7:0] add_980131;
  wire [7:0] sel_980132;
  wire [7:0] add_980135;
  wire [7:0] sel_980136;
  wire [7:0] add_980139;
  wire [7:0] sel_980140;
  wire [7:0] add_980143;
  wire [7:0] sel_980144;
  wire [7:0] add_980147;
  wire [7:0] sel_980148;
  wire [7:0] add_980151;
  wire [7:0] sel_980152;
  wire [7:0] add_980155;
  wire [7:0] sel_980156;
  wire [7:0] add_980159;
  wire [7:0] sel_980160;
  wire [7:0] add_980163;
  wire [7:0] sel_980164;
  wire [7:0] add_980167;
  wire [7:0] sel_980168;
  wire [7:0] add_980171;
  wire [7:0] sel_980172;
  wire [7:0] add_980175;
  wire [7:0] sel_980176;
  wire [7:0] add_980179;
  wire [7:0] sel_980180;
  wire [7:0] add_980183;
  wire [7:0] sel_980184;
  wire [7:0] add_980187;
  wire [7:0] sel_980188;
  wire [7:0] add_980191;
  wire [7:0] sel_980192;
  wire [7:0] add_980195;
  wire [7:0] sel_980196;
  wire [7:0] add_980199;
  wire [7:0] sel_980200;
  wire [7:0] add_980203;
  wire [7:0] sel_980204;
  wire [7:0] add_980207;
  wire [7:0] sel_980208;
  wire [7:0] add_980211;
  wire [7:0] sel_980212;
  wire [7:0] add_980215;
  wire [7:0] sel_980216;
  wire [7:0] add_980219;
  wire [7:0] sel_980220;
  wire [7:0] add_980223;
  wire [7:0] sel_980224;
  wire [7:0] add_980227;
  wire [7:0] sel_980228;
  wire [7:0] add_980231;
  wire [7:0] sel_980232;
  wire [7:0] add_980235;
  wire [7:0] sel_980236;
  wire [7:0] add_980239;
  wire [7:0] sel_980240;
  wire [7:0] add_980243;
  wire [7:0] sel_980244;
  wire [7:0] add_980247;
  wire [7:0] sel_980248;
  wire [7:0] add_980251;
  wire [7:0] sel_980252;
  wire [7:0] add_980255;
  wire [7:0] sel_980256;
  wire [7:0] add_980259;
  wire [7:0] sel_980260;
  wire [7:0] add_980263;
  wire [7:0] sel_980264;
  wire [7:0] add_980267;
  wire [7:0] sel_980268;
  wire [7:0] add_980271;
  wire [7:0] sel_980272;
  wire [7:0] add_980275;
  wire [7:0] sel_980276;
  wire [7:0] add_980279;
  wire [7:0] sel_980280;
  wire [7:0] add_980283;
  wire [7:0] sel_980284;
  wire [7:0] add_980287;
  wire [7:0] sel_980288;
  wire [7:0] add_980291;
  wire [7:0] sel_980292;
  wire [7:0] add_980295;
  wire [7:0] sel_980296;
  wire [7:0] add_980299;
  wire [7:0] sel_980300;
  wire [7:0] add_980303;
  wire [7:0] sel_980304;
  wire [7:0] add_980307;
  wire [7:0] sel_980308;
  wire [7:0] add_980311;
  wire [7:0] sel_980312;
  wire [7:0] add_980315;
  wire [7:0] sel_980316;
  wire [7:0] add_980319;
  wire [7:0] sel_980320;
  wire [7:0] add_980323;
  wire [7:0] sel_980324;
  wire [7:0] add_980327;
  wire [7:0] sel_980328;
  wire [7:0] add_980331;
  wire [7:0] sel_980332;
  wire [7:0] add_980335;
  wire [7:0] sel_980336;
  wire [7:0] add_980339;
  wire [7:0] sel_980340;
  wire [7:0] add_980343;
  wire [7:0] sel_980344;
  wire [7:0] add_980347;
  wire [7:0] sel_980348;
  wire [7:0] add_980351;
  wire [7:0] sel_980352;
  wire [7:0] add_980355;
  wire [7:0] sel_980356;
  wire [7:0] add_980359;
  wire [7:0] sel_980360;
  wire [7:0] add_980363;
  wire [7:0] sel_980364;
  wire [7:0] add_980367;
  wire [7:0] sel_980368;
  wire [7:0] add_980371;
  wire [7:0] sel_980372;
  wire [7:0] add_980375;
  wire [7:0] sel_980376;
  wire [7:0] add_980379;
  wire [7:0] sel_980380;
  wire [7:0] add_980383;
  wire [7:0] sel_980384;
  wire [7:0] add_980387;
  wire [7:0] sel_980388;
  wire [7:0] add_980391;
  wire [7:0] sel_980392;
  wire [7:0] add_980395;
  wire [7:0] sel_980396;
  wire [7:0] add_980399;
  wire [7:0] sel_980400;
  wire [7:0] add_980403;
  wire [7:0] sel_980404;
  wire [7:0] add_980407;
  wire [7:0] sel_980408;
  wire [7:0] add_980411;
  wire [7:0] sel_980412;
  wire [7:0] add_980415;
  wire [7:0] sel_980416;
  wire [7:0] add_980419;
  wire [7:0] sel_980420;
  wire [7:0] add_980423;
  wire [7:0] sel_980424;
  wire [7:0] add_980427;
  wire [7:0] sel_980428;
  wire [7:0] add_980431;
  wire [7:0] sel_980432;
  wire [7:0] add_980435;
  wire [7:0] sel_980436;
  wire [7:0] add_980439;
  wire [7:0] sel_980440;
  wire [7:0] add_980443;
  wire [7:0] sel_980444;
  wire [7:0] add_980448;
  wire [15:0] array_index_980449;
  wire [7:0] sel_980450;
  wire [7:0] add_980453;
  wire [7:0] sel_980454;
  wire [7:0] add_980457;
  wire [7:0] sel_980458;
  wire [7:0] add_980461;
  wire [7:0] sel_980462;
  wire [7:0] add_980465;
  wire [7:0] sel_980466;
  wire [7:0] add_980469;
  wire [7:0] sel_980470;
  wire [7:0] add_980473;
  wire [7:0] sel_980474;
  wire [7:0] add_980477;
  wire [7:0] sel_980478;
  wire [7:0] add_980481;
  wire [7:0] sel_980482;
  wire [7:0] add_980485;
  wire [7:0] sel_980486;
  wire [7:0] add_980489;
  wire [7:0] sel_980490;
  wire [7:0] add_980493;
  wire [7:0] sel_980494;
  wire [7:0] add_980497;
  wire [7:0] sel_980498;
  wire [7:0] add_980501;
  wire [7:0] sel_980502;
  wire [7:0] add_980505;
  wire [7:0] sel_980506;
  wire [7:0] add_980509;
  wire [7:0] sel_980510;
  wire [7:0] add_980513;
  wire [7:0] sel_980514;
  wire [7:0] add_980517;
  wire [7:0] sel_980518;
  wire [7:0] add_980521;
  wire [7:0] sel_980522;
  wire [7:0] add_980525;
  wire [7:0] sel_980526;
  wire [7:0] add_980529;
  wire [7:0] sel_980530;
  wire [7:0] add_980533;
  wire [7:0] sel_980534;
  wire [7:0] add_980537;
  wire [7:0] sel_980538;
  wire [7:0] add_980541;
  wire [7:0] sel_980542;
  wire [7:0] add_980545;
  wire [7:0] sel_980546;
  wire [7:0] add_980549;
  wire [7:0] sel_980550;
  wire [7:0] add_980553;
  wire [7:0] sel_980554;
  wire [7:0] add_980557;
  wire [7:0] sel_980558;
  wire [7:0] add_980561;
  wire [7:0] sel_980562;
  wire [7:0] add_980565;
  wire [7:0] sel_980566;
  wire [7:0] add_980569;
  wire [7:0] sel_980570;
  wire [7:0] add_980573;
  wire [7:0] sel_980574;
  wire [7:0] add_980577;
  wire [7:0] sel_980578;
  wire [7:0] add_980581;
  wire [7:0] sel_980582;
  wire [7:0] add_980585;
  wire [7:0] sel_980586;
  wire [7:0] add_980589;
  wire [7:0] sel_980590;
  wire [7:0] add_980593;
  wire [7:0] sel_980594;
  wire [7:0] add_980597;
  wire [7:0] sel_980598;
  wire [7:0] add_980601;
  wire [7:0] sel_980602;
  wire [7:0] add_980605;
  wire [7:0] sel_980606;
  wire [7:0] add_980609;
  wire [7:0] sel_980610;
  wire [7:0] add_980613;
  wire [7:0] sel_980614;
  wire [7:0] add_980617;
  wire [7:0] sel_980618;
  wire [7:0] add_980621;
  wire [7:0] sel_980622;
  wire [7:0] add_980625;
  wire [7:0] sel_980626;
  wire [7:0] add_980629;
  wire [7:0] sel_980630;
  wire [7:0] add_980633;
  wire [7:0] sel_980634;
  wire [7:0] add_980637;
  wire [7:0] sel_980638;
  wire [7:0] add_980641;
  wire [7:0] sel_980642;
  wire [7:0] add_980645;
  wire [7:0] sel_980646;
  wire [7:0] add_980649;
  wire [7:0] sel_980650;
  wire [7:0] add_980653;
  wire [7:0] sel_980654;
  wire [7:0] add_980657;
  wire [7:0] sel_980658;
  wire [7:0] add_980661;
  wire [7:0] sel_980662;
  wire [7:0] add_980665;
  wire [7:0] sel_980666;
  wire [7:0] add_980669;
  wire [7:0] sel_980670;
  wire [7:0] add_980673;
  wire [7:0] sel_980674;
  wire [7:0] add_980677;
  wire [7:0] sel_980678;
  wire [7:0] add_980681;
  wire [7:0] sel_980682;
  wire [7:0] add_980685;
  wire [7:0] sel_980686;
  wire [7:0] add_980689;
  wire [7:0] sel_980690;
  wire [7:0] add_980693;
  wire [7:0] sel_980694;
  wire [7:0] add_980697;
  wire [7:0] sel_980698;
  wire [7:0] add_980701;
  wire [7:0] sel_980702;
  wire [7:0] add_980705;
  wire [7:0] sel_980706;
  wire [7:0] add_980709;
  wire [7:0] sel_980710;
  wire [7:0] add_980713;
  wire [7:0] sel_980714;
  wire [7:0] add_980717;
  wire [7:0] sel_980718;
  wire [7:0] add_980721;
  wire [7:0] sel_980722;
  wire [7:0] add_980725;
  wire [7:0] sel_980726;
  wire [7:0] add_980729;
  wire [7:0] sel_980730;
  wire [7:0] add_980733;
  wire [7:0] sel_980734;
  wire [7:0] add_980737;
  wire [7:0] sel_980738;
  wire [7:0] add_980741;
  wire [7:0] sel_980742;
  wire [7:0] add_980745;
  wire [7:0] sel_980746;
  wire [7:0] add_980749;
  wire [7:0] sel_980750;
  wire [7:0] add_980753;
  wire [7:0] sel_980754;
  wire [7:0] add_980757;
  wire [7:0] sel_980758;
  wire [7:0] add_980761;
  wire [7:0] sel_980762;
  wire [7:0] add_980765;
  wire [7:0] sel_980766;
  wire [7:0] add_980769;
  wire [7:0] sel_980770;
  wire [7:0] add_980773;
  wire [7:0] sel_980774;
  wire [7:0] add_980777;
  wire [7:0] sel_980778;
  wire [7:0] add_980781;
  wire [7:0] sel_980782;
  wire [7:0] add_980785;
  wire [7:0] sel_980786;
  wire [7:0] add_980789;
  wire [7:0] sel_980790;
  wire [7:0] add_980793;
  wire [7:0] sel_980794;
  wire [7:0] add_980797;
  wire [7:0] sel_980798;
  wire [7:0] add_980801;
  wire [7:0] sel_980802;
  wire [7:0] add_980805;
  wire [7:0] sel_980806;
  wire [7:0] add_980809;
  wire [7:0] sel_980810;
  wire [7:0] add_980813;
  wire [7:0] sel_980814;
  wire [7:0] add_980817;
  wire [7:0] sel_980818;
  wire [7:0] add_980821;
  wire [7:0] sel_980822;
  wire [7:0] add_980825;
  wire [7:0] sel_980826;
  wire [7:0] add_980829;
  wire [7:0] sel_980830;
  wire [7:0] add_980833;
  wire [7:0] sel_980834;
  wire [7:0] add_980837;
  wire [7:0] sel_980838;
  wire [7:0] add_980841;
  wire [7:0] sel_980842;
  wire [7:0] add_980845;
  wire [7:0] sel_980846;
  wire [7:0] add_980850;
  wire [15:0] array_index_980851;
  wire [7:0] sel_980852;
  wire [7:0] add_980855;
  wire [7:0] sel_980856;
  wire [7:0] add_980859;
  wire [7:0] sel_980860;
  wire [7:0] add_980863;
  wire [7:0] sel_980864;
  wire [7:0] add_980867;
  wire [7:0] sel_980868;
  wire [7:0] add_980871;
  wire [7:0] sel_980872;
  wire [7:0] add_980875;
  wire [7:0] sel_980876;
  wire [7:0] add_980879;
  wire [7:0] sel_980880;
  wire [7:0] add_980883;
  wire [7:0] sel_980884;
  wire [7:0] add_980887;
  wire [7:0] sel_980888;
  wire [7:0] add_980891;
  wire [7:0] sel_980892;
  wire [7:0] add_980895;
  wire [7:0] sel_980896;
  wire [7:0] add_980899;
  wire [7:0] sel_980900;
  wire [7:0] add_980903;
  wire [7:0] sel_980904;
  wire [7:0] add_980907;
  wire [7:0] sel_980908;
  wire [7:0] add_980911;
  wire [7:0] sel_980912;
  wire [7:0] add_980915;
  wire [7:0] sel_980916;
  wire [7:0] add_980919;
  wire [7:0] sel_980920;
  wire [7:0] add_980923;
  wire [7:0] sel_980924;
  wire [7:0] add_980927;
  wire [7:0] sel_980928;
  wire [7:0] add_980931;
  wire [7:0] sel_980932;
  wire [7:0] add_980935;
  wire [7:0] sel_980936;
  wire [7:0] add_980939;
  wire [7:0] sel_980940;
  wire [7:0] add_980943;
  wire [7:0] sel_980944;
  wire [7:0] add_980947;
  wire [7:0] sel_980948;
  wire [7:0] add_980951;
  wire [7:0] sel_980952;
  wire [7:0] add_980955;
  wire [7:0] sel_980956;
  wire [7:0] add_980959;
  wire [7:0] sel_980960;
  wire [7:0] add_980963;
  wire [7:0] sel_980964;
  wire [7:0] add_980967;
  wire [7:0] sel_980968;
  wire [7:0] add_980971;
  wire [7:0] sel_980972;
  wire [7:0] add_980975;
  wire [7:0] sel_980976;
  wire [7:0] add_980979;
  wire [7:0] sel_980980;
  wire [7:0] add_980983;
  wire [7:0] sel_980984;
  wire [7:0] add_980987;
  wire [7:0] sel_980988;
  wire [7:0] add_980991;
  wire [7:0] sel_980992;
  wire [7:0] add_980995;
  wire [7:0] sel_980996;
  wire [7:0] add_980999;
  wire [7:0] sel_981000;
  wire [7:0] add_981003;
  wire [7:0] sel_981004;
  wire [7:0] add_981007;
  wire [7:0] sel_981008;
  wire [7:0] add_981011;
  wire [7:0] sel_981012;
  wire [7:0] add_981015;
  wire [7:0] sel_981016;
  wire [7:0] add_981019;
  wire [7:0] sel_981020;
  wire [7:0] add_981023;
  wire [7:0] sel_981024;
  wire [7:0] add_981027;
  wire [7:0] sel_981028;
  wire [7:0] add_981031;
  wire [7:0] sel_981032;
  wire [7:0] add_981035;
  wire [7:0] sel_981036;
  wire [7:0] add_981039;
  wire [7:0] sel_981040;
  wire [7:0] add_981043;
  wire [7:0] sel_981044;
  wire [7:0] add_981047;
  wire [7:0] sel_981048;
  wire [7:0] add_981051;
  wire [7:0] sel_981052;
  wire [7:0] add_981055;
  wire [7:0] sel_981056;
  wire [7:0] add_981059;
  wire [7:0] sel_981060;
  wire [7:0] add_981063;
  wire [7:0] sel_981064;
  wire [7:0] add_981067;
  wire [7:0] sel_981068;
  wire [7:0] add_981071;
  wire [7:0] sel_981072;
  wire [7:0] add_981075;
  wire [7:0] sel_981076;
  wire [7:0] add_981079;
  wire [7:0] sel_981080;
  wire [7:0] add_981083;
  wire [7:0] sel_981084;
  wire [7:0] add_981087;
  wire [7:0] sel_981088;
  wire [7:0] add_981091;
  wire [7:0] sel_981092;
  wire [7:0] add_981095;
  wire [7:0] sel_981096;
  wire [7:0] add_981099;
  wire [7:0] sel_981100;
  wire [7:0] add_981103;
  wire [7:0] sel_981104;
  wire [7:0] add_981107;
  wire [7:0] sel_981108;
  wire [7:0] add_981111;
  wire [7:0] sel_981112;
  wire [7:0] add_981115;
  wire [7:0] sel_981116;
  wire [7:0] add_981119;
  wire [7:0] sel_981120;
  wire [7:0] add_981123;
  wire [7:0] sel_981124;
  wire [7:0] add_981127;
  wire [7:0] sel_981128;
  wire [7:0] add_981131;
  wire [7:0] sel_981132;
  wire [7:0] add_981135;
  wire [7:0] sel_981136;
  wire [7:0] add_981139;
  wire [7:0] sel_981140;
  wire [7:0] add_981143;
  wire [7:0] sel_981144;
  wire [7:0] add_981147;
  wire [7:0] sel_981148;
  wire [7:0] add_981151;
  wire [7:0] sel_981152;
  wire [7:0] add_981155;
  wire [7:0] sel_981156;
  wire [7:0] add_981159;
  wire [7:0] sel_981160;
  wire [7:0] add_981163;
  wire [7:0] sel_981164;
  wire [7:0] add_981167;
  wire [7:0] sel_981168;
  wire [7:0] add_981171;
  wire [7:0] sel_981172;
  wire [7:0] add_981175;
  wire [7:0] sel_981176;
  wire [7:0] add_981179;
  wire [7:0] sel_981180;
  wire [7:0] add_981183;
  wire [7:0] sel_981184;
  wire [7:0] add_981187;
  wire [7:0] sel_981188;
  wire [7:0] add_981191;
  wire [7:0] sel_981192;
  wire [7:0] add_981195;
  wire [7:0] sel_981196;
  wire [7:0] add_981199;
  wire [7:0] sel_981200;
  wire [7:0] add_981203;
  wire [7:0] sel_981204;
  wire [7:0] add_981207;
  wire [7:0] sel_981208;
  wire [7:0] add_981211;
  wire [7:0] sel_981212;
  wire [7:0] add_981215;
  wire [7:0] sel_981216;
  wire [7:0] add_981219;
  wire [7:0] sel_981220;
  wire [7:0] add_981223;
  wire [7:0] sel_981224;
  wire [7:0] add_981227;
  wire [7:0] sel_981228;
  wire [7:0] add_981231;
  wire [7:0] sel_981232;
  wire [7:0] add_981235;
  wire [7:0] sel_981236;
  wire [7:0] add_981239;
  wire [7:0] sel_981240;
  wire [7:0] add_981243;
  wire [7:0] sel_981244;
  wire [7:0] add_981247;
  wire [7:0] sel_981248;
  wire [7:0] add_981252;
  wire [15:0] array_index_981253;
  wire [7:0] sel_981254;
  wire [7:0] add_981257;
  wire [7:0] sel_981258;
  wire [7:0] add_981261;
  wire [7:0] sel_981262;
  wire [7:0] add_981265;
  wire [7:0] sel_981266;
  wire [7:0] add_981269;
  wire [7:0] sel_981270;
  wire [7:0] add_981273;
  wire [7:0] sel_981274;
  wire [7:0] add_981277;
  wire [7:0] sel_981278;
  wire [7:0] add_981281;
  wire [7:0] sel_981282;
  wire [7:0] add_981285;
  wire [7:0] sel_981286;
  wire [7:0] add_981289;
  wire [7:0] sel_981290;
  wire [7:0] add_981293;
  wire [7:0] sel_981294;
  wire [7:0] add_981297;
  wire [7:0] sel_981298;
  wire [7:0] add_981301;
  wire [7:0] sel_981302;
  wire [7:0] add_981305;
  wire [7:0] sel_981306;
  wire [7:0] add_981309;
  wire [7:0] sel_981310;
  wire [7:0] add_981313;
  wire [7:0] sel_981314;
  wire [7:0] add_981317;
  wire [7:0] sel_981318;
  wire [7:0] add_981321;
  wire [7:0] sel_981322;
  wire [7:0] add_981325;
  wire [7:0] sel_981326;
  wire [7:0] add_981329;
  wire [7:0] sel_981330;
  wire [7:0] add_981333;
  wire [7:0] sel_981334;
  wire [7:0] add_981337;
  wire [7:0] sel_981338;
  wire [7:0] add_981341;
  wire [7:0] sel_981342;
  wire [7:0] add_981345;
  wire [7:0] sel_981346;
  wire [7:0] add_981349;
  wire [7:0] sel_981350;
  wire [7:0] add_981353;
  wire [7:0] sel_981354;
  wire [7:0] add_981357;
  wire [7:0] sel_981358;
  wire [7:0] add_981361;
  wire [7:0] sel_981362;
  wire [7:0] add_981365;
  wire [7:0] sel_981366;
  wire [7:0] add_981369;
  wire [7:0] sel_981370;
  wire [7:0] add_981373;
  wire [7:0] sel_981374;
  wire [7:0] add_981377;
  wire [7:0] sel_981378;
  wire [7:0] add_981381;
  wire [7:0] sel_981382;
  wire [7:0] add_981385;
  wire [7:0] sel_981386;
  wire [7:0] add_981389;
  wire [7:0] sel_981390;
  wire [7:0] add_981393;
  wire [7:0] sel_981394;
  wire [7:0] add_981397;
  wire [7:0] sel_981398;
  wire [7:0] add_981401;
  wire [7:0] sel_981402;
  wire [7:0] add_981405;
  wire [7:0] sel_981406;
  wire [7:0] add_981409;
  wire [7:0] sel_981410;
  wire [7:0] add_981413;
  wire [7:0] sel_981414;
  wire [7:0] add_981417;
  wire [7:0] sel_981418;
  wire [7:0] add_981421;
  wire [7:0] sel_981422;
  wire [7:0] add_981425;
  wire [7:0] sel_981426;
  wire [7:0] add_981429;
  wire [7:0] sel_981430;
  wire [7:0] add_981433;
  wire [7:0] sel_981434;
  wire [7:0] add_981437;
  wire [7:0] sel_981438;
  wire [7:0] add_981441;
  wire [7:0] sel_981442;
  wire [7:0] add_981445;
  wire [7:0] sel_981446;
  wire [7:0] add_981449;
  wire [7:0] sel_981450;
  wire [7:0] add_981453;
  wire [7:0] sel_981454;
  wire [7:0] add_981457;
  wire [7:0] sel_981458;
  wire [7:0] add_981461;
  wire [7:0] sel_981462;
  wire [7:0] add_981465;
  wire [7:0] sel_981466;
  wire [7:0] add_981469;
  wire [7:0] sel_981470;
  wire [7:0] add_981473;
  wire [7:0] sel_981474;
  wire [7:0] add_981477;
  wire [7:0] sel_981478;
  wire [7:0] add_981481;
  wire [7:0] sel_981482;
  wire [7:0] add_981485;
  wire [7:0] sel_981486;
  wire [7:0] add_981489;
  wire [7:0] sel_981490;
  wire [7:0] add_981493;
  wire [7:0] sel_981494;
  wire [7:0] add_981497;
  wire [7:0] sel_981498;
  wire [7:0] add_981501;
  wire [7:0] sel_981502;
  wire [7:0] add_981505;
  wire [7:0] sel_981506;
  wire [7:0] add_981509;
  wire [7:0] sel_981510;
  wire [7:0] add_981513;
  wire [7:0] sel_981514;
  wire [7:0] add_981517;
  wire [7:0] sel_981518;
  wire [7:0] add_981521;
  wire [7:0] sel_981522;
  wire [7:0] add_981525;
  wire [7:0] sel_981526;
  wire [7:0] add_981529;
  wire [7:0] sel_981530;
  wire [7:0] add_981533;
  wire [7:0] sel_981534;
  wire [7:0] add_981537;
  wire [7:0] sel_981538;
  wire [7:0] add_981541;
  wire [7:0] sel_981542;
  wire [7:0] add_981545;
  wire [7:0] sel_981546;
  wire [7:0] add_981549;
  wire [7:0] sel_981550;
  wire [7:0] add_981553;
  wire [7:0] sel_981554;
  wire [7:0] add_981557;
  wire [7:0] sel_981558;
  wire [7:0] add_981561;
  wire [7:0] sel_981562;
  wire [7:0] add_981565;
  wire [7:0] sel_981566;
  wire [7:0] add_981569;
  wire [7:0] sel_981570;
  wire [7:0] add_981573;
  wire [7:0] sel_981574;
  wire [7:0] add_981577;
  wire [7:0] sel_981578;
  wire [7:0] add_981581;
  wire [7:0] sel_981582;
  wire [7:0] add_981585;
  wire [7:0] sel_981586;
  wire [7:0] add_981589;
  wire [7:0] sel_981590;
  wire [7:0] add_981593;
  wire [7:0] sel_981594;
  wire [7:0] add_981597;
  wire [7:0] sel_981598;
  wire [7:0] add_981601;
  wire [7:0] sel_981602;
  wire [7:0] add_981605;
  wire [7:0] sel_981606;
  wire [7:0] add_981609;
  wire [7:0] sel_981610;
  wire [7:0] add_981613;
  wire [7:0] sel_981614;
  wire [7:0] add_981617;
  wire [7:0] sel_981618;
  wire [7:0] add_981621;
  wire [7:0] sel_981622;
  wire [7:0] add_981625;
  wire [7:0] sel_981626;
  wire [7:0] add_981629;
  wire [7:0] sel_981630;
  wire [7:0] add_981633;
  wire [7:0] sel_981634;
  wire [7:0] add_981637;
  wire [7:0] sel_981638;
  wire [7:0] add_981641;
  wire [7:0] sel_981642;
  wire [7:0] add_981645;
  wire [7:0] sel_981646;
  wire [7:0] add_981649;
  wire [7:0] sel_981650;
  wire [7:0] add_981654;
  wire [15:0] array_index_981655;
  wire [7:0] sel_981656;
  wire [7:0] add_981659;
  wire [7:0] sel_981660;
  wire [7:0] add_981663;
  wire [7:0] sel_981664;
  wire [7:0] add_981667;
  wire [7:0] sel_981668;
  wire [7:0] add_981671;
  wire [7:0] sel_981672;
  wire [7:0] add_981675;
  wire [7:0] sel_981676;
  wire [7:0] add_981679;
  wire [7:0] sel_981680;
  wire [7:0] add_981683;
  wire [7:0] sel_981684;
  wire [7:0] add_981687;
  wire [7:0] sel_981688;
  wire [7:0] add_981691;
  wire [7:0] sel_981692;
  wire [7:0] add_981695;
  wire [7:0] sel_981696;
  wire [7:0] add_981699;
  wire [7:0] sel_981700;
  wire [7:0] add_981703;
  wire [7:0] sel_981704;
  wire [7:0] add_981707;
  wire [7:0] sel_981708;
  wire [7:0] add_981711;
  wire [7:0] sel_981712;
  wire [7:0] add_981715;
  wire [7:0] sel_981716;
  wire [7:0] add_981719;
  wire [7:0] sel_981720;
  wire [7:0] add_981723;
  wire [7:0] sel_981724;
  wire [7:0] add_981727;
  wire [7:0] sel_981728;
  wire [7:0] add_981731;
  wire [7:0] sel_981732;
  wire [7:0] add_981735;
  wire [7:0] sel_981736;
  wire [7:0] add_981739;
  wire [7:0] sel_981740;
  wire [7:0] add_981743;
  wire [7:0] sel_981744;
  wire [7:0] add_981747;
  wire [7:0] sel_981748;
  wire [7:0] add_981751;
  wire [7:0] sel_981752;
  wire [7:0] add_981755;
  wire [7:0] sel_981756;
  wire [7:0] add_981759;
  wire [7:0] sel_981760;
  wire [7:0] add_981763;
  wire [7:0] sel_981764;
  wire [7:0] add_981767;
  wire [7:0] sel_981768;
  wire [7:0] add_981771;
  wire [7:0] sel_981772;
  wire [7:0] add_981775;
  wire [7:0] sel_981776;
  wire [7:0] add_981779;
  wire [7:0] sel_981780;
  wire [7:0] add_981783;
  wire [7:0] sel_981784;
  wire [7:0] add_981787;
  wire [7:0] sel_981788;
  wire [7:0] add_981791;
  wire [7:0] sel_981792;
  wire [7:0] add_981795;
  wire [7:0] sel_981796;
  wire [7:0] add_981799;
  wire [7:0] sel_981800;
  wire [7:0] add_981803;
  wire [7:0] sel_981804;
  wire [7:0] add_981807;
  wire [7:0] sel_981808;
  wire [7:0] add_981811;
  wire [7:0] sel_981812;
  wire [7:0] add_981815;
  wire [7:0] sel_981816;
  wire [7:0] add_981819;
  wire [7:0] sel_981820;
  wire [7:0] add_981823;
  wire [7:0] sel_981824;
  wire [7:0] add_981827;
  wire [7:0] sel_981828;
  wire [7:0] add_981831;
  wire [7:0] sel_981832;
  wire [7:0] add_981835;
  wire [7:0] sel_981836;
  wire [7:0] add_981839;
  wire [7:0] sel_981840;
  wire [7:0] add_981843;
  wire [7:0] sel_981844;
  wire [7:0] add_981847;
  wire [7:0] sel_981848;
  wire [7:0] add_981851;
  wire [7:0] sel_981852;
  wire [7:0] add_981855;
  wire [7:0] sel_981856;
  wire [7:0] add_981859;
  wire [7:0] sel_981860;
  wire [7:0] add_981863;
  wire [7:0] sel_981864;
  wire [7:0] add_981867;
  wire [7:0] sel_981868;
  wire [7:0] add_981871;
  wire [7:0] sel_981872;
  wire [7:0] add_981875;
  wire [7:0] sel_981876;
  wire [7:0] add_981879;
  wire [7:0] sel_981880;
  wire [7:0] add_981883;
  wire [7:0] sel_981884;
  wire [7:0] add_981887;
  wire [7:0] sel_981888;
  wire [7:0] add_981891;
  wire [7:0] sel_981892;
  wire [7:0] add_981895;
  wire [7:0] sel_981896;
  wire [7:0] add_981899;
  wire [7:0] sel_981900;
  wire [7:0] add_981903;
  wire [7:0] sel_981904;
  wire [7:0] add_981907;
  wire [7:0] sel_981908;
  wire [7:0] add_981911;
  wire [7:0] sel_981912;
  wire [7:0] add_981915;
  wire [7:0] sel_981916;
  wire [7:0] add_981919;
  wire [7:0] sel_981920;
  wire [7:0] add_981923;
  wire [7:0] sel_981924;
  wire [7:0] add_981927;
  wire [7:0] sel_981928;
  wire [7:0] add_981931;
  wire [7:0] sel_981932;
  wire [7:0] add_981935;
  wire [7:0] sel_981936;
  wire [7:0] add_981939;
  wire [7:0] sel_981940;
  wire [7:0] add_981943;
  wire [7:0] sel_981944;
  wire [7:0] add_981947;
  wire [7:0] sel_981948;
  wire [7:0] add_981951;
  wire [7:0] sel_981952;
  wire [7:0] add_981955;
  wire [7:0] sel_981956;
  wire [7:0] add_981959;
  wire [7:0] sel_981960;
  wire [7:0] add_981963;
  wire [7:0] sel_981964;
  wire [7:0] add_981967;
  wire [7:0] sel_981968;
  wire [7:0] add_981971;
  wire [7:0] sel_981972;
  wire [7:0] add_981975;
  wire [7:0] sel_981976;
  wire [7:0] add_981979;
  wire [7:0] sel_981980;
  wire [7:0] add_981983;
  wire [7:0] sel_981984;
  wire [7:0] add_981987;
  wire [7:0] sel_981988;
  wire [7:0] add_981991;
  wire [7:0] sel_981992;
  wire [7:0] add_981995;
  wire [7:0] sel_981996;
  wire [7:0] add_981999;
  wire [7:0] sel_982000;
  wire [7:0] add_982003;
  wire [7:0] sel_982004;
  wire [7:0] add_982007;
  wire [7:0] sel_982008;
  wire [7:0] add_982011;
  wire [7:0] sel_982012;
  wire [7:0] add_982015;
  wire [7:0] sel_982016;
  wire [7:0] add_982019;
  wire [7:0] sel_982020;
  wire [7:0] add_982023;
  wire [7:0] sel_982024;
  wire [7:0] add_982027;
  wire [7:0] sel_982028;
  wire [7:0] add_982031;
  wire [7:0] sel_982032;
  wire [7:0] add_982035;
  wire [7:0] sel_982036;
  wire [7:0] add_982039;
  wire [7:0] sel_982040;
  wire [7:0] add_982043;
  wire [7:0] sel_982044;
  wire [7:0] add_982047;
  wire [7:0] sel_982048;
  wire [7:0] add_982051;
  wire [7:0] sel_982052;
  wire [7:0] add_982056;
  wire [15:0] array_index_982057;
  wire [7:0] sel_982058;
  wire [7:0] add_982061;
  wire [7:0] sel_982062;
  wire [7:0] add_982065;
  wire [7:0] sel_982066;
  wire [7:0] add_982069;
  wire [7:0] sel_982070;
  wire [7:0] add_982073;
  wire [7:0] sel_982074;
  wire [7:0] add_982077;
  wire [7:0] sel_982078;
  wire [7:0] add_982081;
  wire [7:0] sel_982082;
  wire [7:0] add_982085;
  wire [7:0] sel_982086;
  wire [7:0] add_982089;
  wire [7:0] sel_982090;
  wire [7:0] add_982093;
  wire [7:0] sel_982094;
  wire [7:0] add_982097;
  wire [7:0] sel_982098;
  wire [7:0] add_982101;
  wire [7:0] sel_982102;
  wire [7:0] add_982105;
  wire [7:0] sel_982106;
  wire [7:0] add_982109;
  wire [7:0] sel_982110;
  wire [7:0] add_982113;
  wire [7:0] sel_982114;
  wire [7:0] add_982117;
  wire [7:0] sel_982118;
  wire [7:0] add_982121;
  wire [7:0] sel_982122;
  wire [7:0] add_982125;
  wire [7:0] sel_982126;
  wire [7:0] add_982129;
  wire [7:0] sel_982130;
  wire [7:0] add_982133;
  wire [7:0] sel_982134;
  wire [7:0] add_982137;
  wire [7:0] sel_982138;
  wire [7:0] add_982141;
  wire [7:0] sel_982142;
  wire [7:0] add_982145;
  wire [7:0] sel_982146;
  wire [7:0] add_982149;
  wire [7:0] sel_982150;
  wire [7:0] add_982153;
  wire [7:0] sel_982154;
  wire [7:0] add_982157;
  wire [7:0] sel_982158;
  wire [7:0] add_982161;
  wire [7:0] sel_982162;
  wire [7:0] add_982165;
  wire [7:0] sel_982166;
  wire [7:0] add_982169;
  wire [7:0] sel_982170;
  wire [7:0] add_982173;
  wire [7:0] sel_982174;
  wire [7:0] add_982177;
  wire [7:0] sel_982178;
  wire [7:0] add_982181;
  wire [7:0] sel_982182;
  wire [7:0] add_982185;
  wire [7:0] sel_982186;
  wire [7:0] add_982189;
  wire [7:0] sel_982190;
  wire [7:0] add_982193;
  wire [7:0] sel_982194;
  wire [7:0] add_982197;
  wire [7:0] sel_982198;
  wire [7:0] add_982201;
  wire [7:0] sel_982202;
  wire [7:0] add_982205;
  wire [7:0] sel_982206;
  wire [7:0] add_982209;
  wire [7:0] sel_982210;
  wire [7:0] add_982213;
  wire [7:0] sel_982214;
  wire [7:0] add_982217;
  wire [7:0] sel_982218;
  wire [7:0] add_982221;
  wire [7:0] sel_982222;
  wire [7:0] add_982225;
  wire [7:0] sel_982226;
  wire [7:0] add_982229;
  wire [7:0] sel_982230;
  wire [7:0] add_982233;
  wire [7:0] sel_982234;
  wire [7:0] add_982237;
  wire [7:0] sel_982238;
  wire [7:0] add_982241;
  wire [7:0] sel_982242;
  wire [7:0] add_982245;
  wire [7:0] sel_982246;
  wire [7:0] add_982249;
  wire [7:0] sel_982250;
  wire [7:0] add_982253;
  wire [7:0] sel_982254;
  wire [7:0] add_982257;
  wire [7:0] sel_982258;
  wire [7:0] add_982261;
  wire [7:0] sel_982262;
  wire [7:0] add_982265;
  wire [7:0] sel_982266;
  wire [7:0] add_982269;
  wire [7:0] sel_982270;
  wire [7:0] add_982273;
  wire [7:0] sel_982274;
  wire [7:0] add_982277;
  wire [7:0] sel_982278;
  wire [7:0] add_982281;
  wire [7:0] sel_982282;
  wire [7:0] add_982285;
  wire [7:0] sel_982286;
  wire [7:0] add_982289;
  wire [7:0] sel_982290;
  wire [7:0] add_982293;
  wire [7:0] sel_982294;
  wire [7:0] add_982297;
  wire [7:0] sel_982298;
  wire [7:0] add_982301;
  wire [7:0] sel_982302;
  wire [7:0] add_982305;
  wire [7:0] sel_982306;
  wire [7:0] add_982309;
  wire [7:0] sel_982310;
  wire [7:0] add_982313;
  wire [7:0] sel_982314;
  wire [7:0] add_982317;
  wire [7:0] sel_982318;
  wire [7:0] add_982321;
  wire [7:0] sel_982322;
  wire [7:0] add_982325;
  wire [7:0] sel_982326;
  wire [7:0] add_982329;
  wire [7:0] sel_982330;
  wire [7:0] add_982333;
  wire [7:0] sel_982334;
  wire [7:0] add_982337;
  wire [7:0] sel_982338;
  wire [7:0] add_982341;
  wire [7:0] sel_982342;
  wire [7:0] add_982345;
  wire [7:0] sel_982346;
  wire [7:0] add_982349;
  wire [7:0] sel_982350;
  wire [7:0] add_982353;
  wire [7:0] sel_982354;
  wire [7:0] add_982357;
  wire [7:0] sel_982358;
  wire [7:0] add_982361;
  wire [7:0] sel_982362;
  wire [7:0] add_982365;
  wire [7:0] sel_982366;
  wire [7:0] add_982369;
  wire [7:0] sel_982370;
  wire [7:0] add_982373;
  wire [7:0] sel_982374;
  wire [7:0] add_982377;
  wire [7:0] sel_982378;
  wire [7:0] add_982381;
  wire [7:0] sel_982382;
  wire [7:0] add_982385;
  wire [7:0] sel_982386;
  wire [7:0] add_982389;
  wire [7:0] sel_982390;
  wire [7:0] add_982393;
  wire [7:0] sel_982394;
  wire [7:0] add_982397;
  wire [7:0] sel_982398;
  wire [7:0] add_982401;
  wire [7:0] sel_982402;
  wire [7:0] add_982405;
  wire [7:0] sel_982406;
  wire [7:0] add_982409;
  wire [7:0] sel_982410;
  wire [7:0] add_982413;
  wire [7:0] sel_982414;
  wire [7:0] add_982417;
  wire [7:0] sel_982418;
  wire [7:0] add_982421;
  wire [7:0] sel_982422;
  wire [7:0] add_982425;
  wire [7:0] sel_982426;
  wire [7:0] add_982429;
  wire [7:0] sel_982430;
  wire [7:0] add_982433;
  wire [7:0] sel_982434;
  wire [7:0] add_982437;
  wire [7:0] sel_982438;
  wire [7:0] add_982441;
  wire [7:0] sel_982442;
  wire [7:0] add_982445;
  wire [7:0] sel_982446;
  wire [7:0] add_982449;
  wire [7:0] sel_982450;
  wire [7:0] add_982453;
  wire [7:0] sel_982454;
  wire [7:0] add_982458;
  wire [15:0] array_index_982459;
  wire [7:0] sel_982460;
  wire [7:0] add_982463;
  wire [7:0] sel_982464;
  wire [7:0] add_982467;
  wire [7:0] sel_982468;
  wire [7:0] add_982471;
  wire [7:0] sel_982472;
  wire [7:0] add_982475;
  wire [7:0] sel_982476;
  wire [7:0] add_982479;
  wire [7:0] sel_982480;
  wire [7:0] add_982483;
  wire [7:0] sel_982484;
  wire [7:0] add_982487;
  wire [7:0] sel_982488;
  wire [7:0] add_982491;
  wire [7:0] sel_982492;
  wire [7:0] add_982495;
  wire [7:0] sel_982496;
  wire [7:0] add_982499;
  wire [7:0] sel_982500;
  wire [7:0] add_982503;
  wire [7:0] sel_982504;
  wire [7:0] add_982507;
  wire [7:0] sel_982508;
  wire [7:0] add_982511;
  wire [7:0] sel_982512;
  wire [7:0] add_982515;
  wire [7:0] sel_982516;
  wire [7:0] add_982519;
  wire [7:0] sel_982520;
  wire [7:0] add_982523;
  wire [7:0] sel_982524;
  wire [7:0] add_982527;
  wire [7:0] sel_982528;
  wire [7:0] add_982531;
  wire [7:0] sel_982532;
  wire [7:0] add_982535;
  wire [7:0] sel_982536;
  wire [7:0] add_982539;
  wire [7:0] sel_982540;
  wire [7:0] add_982543;
  wire [7:0] sel_982544;
  wire [7:0] add_982547;
  wire [7:0] sel_982548;
  wire [7:0] add_982551;
  wire [7:0] sel_982552;
  wire [7:0] add_982555;
  wire [7:0] sel_982556;
  wire [7:0] add_982559;
  wire [7:0] sel_982560;
  wire [7:0] add_982563;
  wire [7:0] sel_982564;
  wire [7:0] add_982567;
  wire [7:0] sel_982568;
  wire [7:0] add_982571;
  wire [7:0] sel_982572;
  wire [7:0] add_982575;
  wire [7:0] sel_982576;
  wire [7:0] add_982579;
  wire [7:0] sel_982580;
  wire [7:0] add_982583;
  wire [7:0] sel_982584;
  wire [7:0] add_982587;
  wire [7:0] sel_982588;
  wire [7:0] add_982591;
  wire [7:0] sel_982592;
  wire [7:0] add_982595;
  wire [7:0] sel_982596;
  wire [7:0] add_982599;
  wire [7:0] sel_982600;
  wire [7:0] add_982603;
  wire [7:0] sel_982604;
  wire [7:0] add_982607;
  wire [7:0] sel_982608;
  wire [7:0] add_982611;
  wire [7:0] sel_982612;
  wire [7:0] add_982615;
  wire [7:0] sel_982616;
  wire [7:0] add_982619;
  wire [7:0] sel_982620;
  wire [7:0] add_982623;
  wire [7:0] sel_982624;
  wire [7:0] add_982627;
  wire [7:0] sel_982628;
  wire [7:0] add_982631;
  wire [7:0] sel_982632;
  wire [7:0] add_982635;
  wire [7:0] sel_982636;
  wire [7:0] add_982639;
  wire [7:0] sel_982640;
  wire [7:0] add_982643;
  wire [7:0] sel_982644;
  wire [7:0] add_982647;
  wire [7:0] sel_982648;
  wire [7:0] add_982651;
  wire [7:0] sel_982652;
  wire [7:0] add_982655;
  wire [7:0] sel_982656;
  wire [7:0] add_982659;
  wire [7:0] sel_982660;
  wire [7:0] add_982663;
  wire [7:0] sel_982664;
  wire [7:0] add_982667;
  wire [7:0] sel_982668;
  wire [7:0] add_982671;
  wire [7:0] sel_982672;
  wire [7:0] add_982675;
  wire [7:0] sel_982676;
  wire [7:0] add_982679;
  wire [7:0] sel_982680;
  wire [7:0] add_982683;
  wire [7:0] sel_982684;
  wire [7:0] add_982687;
  wire [7:0] sel_982688;
  wire [7:0] add_982691;
  wire [7:0] sel_982692;
  wire [7:0] add_982695;
  wire [7:0] sel_982696;
  wire [7:0] add_982699;
  wire [7:0] sel_982700;
  wire [7:0] add_982703;
  wire [7:0] sel_982704;
  wire [7:0] add_982707;
  wire [7:0] sel_982708;
  wire [7:0] add_982711;
  wire [7:0] sel_982712;
  wire [7:0] add_982715;
  wire [7:0] sel_982716;
  wire [7:0] add_982719;
  wire [7:0] sel_982720;
  wire [7:0] add_982723;
  wire [7:0] sel_982724;
  wire [7:0] add_982727;
  wire [7:0] sel_982728;
  wire [7:0] add_982731;
  wire [7:0] sel_982732;
  wire [7:0] add_982735;
  wire [7:0] sel_982736;
  wire [7:0] add_982739;
  wire [7:0] sel_982740;
  wire [7:0] add_982743;
  wire [7:0] sel_982744;
  wire [7:0] add_982747;
  wire [7:0] sel_982748;
  wire [7:0] add_982751;
  wire [7:0] sel_982752;
  wire [7:0] add_982755;
  wire [7:0] sel_982756;
  wire [7:0] add_982759;
  wire [7:0] sel_982760;
  wire [7:0] add_982763;
  wire [7:0] sel_982764;
  wire [7:0] add_982767;
  wire [7:0] sel_982768;
  wire [7:0] add_982771;
  wire [7:0] sel_982772;
  wire [7:0] add_982775;
  wire [7:0] sel_982776;
  wire [7:0] add_982779;
  wire [7:0] sel_982780;
  wire [7:0] add_982783;
  wire [7:0] sel_982784;
  wire [7:0] add_982787;
  wire [7:0] sel_982788;
  wire [7:0] add_982791;
  wire [7:0] sel_982792;
  wire [7:0] add_982795;
  wire [7:0] sel_982796;
  wire [7:0] add_982799;
  wire [7:0] sel_982800;
  wire [7:0] add_982803;
  wire [7:0] sel_982804;
  wire [7:0] add_982807;
  wire [7:0] sel_982808;
  wire [7:0] add_982811;
  wire [7:0] sel_982812;
  wire [7:0] add_982815;
  wire [7:0] sel_982816;
  wire [7:0] add_982819;
  wire [7:0] sel_982820;
  wire [7:0] add_982823;
  wire [7:0] sel_982824;
  wire [7:0] add_982827;
  wire [7:0] sel_982828;
  wire [7:0] add_982831;
  wire [7:0] sel_982832;
  wire [7:0] add_982835;
  wire [7:0] sel_982836;
  wire [7:0] add_982839;
  wire [7:0] sel_982840;
  wire [7:0] add_982843;
  wire [7:0] sel_982844;
  wire [7:0] add_982847;
  wire [7:0] sel_982848;
  wire [7:0] add_982851;
  wire [7:0] sel_982852;
  wire [7:0] add_982855;
  wire [7:0] sel_982856;
  wire [7:0] add_982860;
  wire [15:0] array_index_982861;
  wire [7:0] sel_982862;
  wire [7:0] add_982865;
  wire [7:0] sel_982866;
  wire [7:0] add_982869;
  wire [7:0] sel_982870;
  wire [7:0] add_982873;
  wire [7:0] sel_982874;
  wire [7:0] add_982877;
  wire [7:0] sel_982878;
  wire [7:0] add_982881;
  wire [7:0] sel_982882;
  wire [7:0] add_982885;
  wire [7:0] sel_982886;
  wire [7:0] add_982889;
  wire [7:0] sel_982890;
  wire [7:0] add_982893;
  wire [7:0] sel_982894;
  wire [7:0] add_982897;
  wire [7:0] sel_982898;
  wire [7:0] add_982901;
  wire [7:0] sel_982902;
  wire [7:0] add_982905;
  wire [7:0] sel_982906;
  wire [7:0] add_982909;
  wire [7:0] sel_982910;
  wire [7:0] add_982913;
  wire [7:0] sel_982914;
  wire [7:0] add_982917;
  wire [7:0] sel_982918;
  wire [7:0] add_982921;
  wire [7:0] sel_982922;
  wire [7:0] add_982925;
  wire [7:0] sel_982926;
  wire [7:0] add_982929;
  wire [7:0] sel_982930;
  wire [7:0] add_982933;
  wire [7:0] sel_982934;
  wire [7:0] add_982937;
  wire [7:0] sel_982938;
  wire [7:0] add_982941;
  wire [7:0] sel_982942;
  wire [7:0] add_982945;
  wire [7:0] sel_982946;
  wire [7:0] add_982949;
  wire [7:0] sel_982950;
  wire [7:0] add_982953;
  wire [7:0] sel_982954;
  wire [7:0] add_982957;
  wire [7:0] sel_982958;
  wire [7:0] add_982961;
  wire [7:0] sel_982962;
  wire [7:0] add_982965;
  wire [7:0] sel_982966;
  wire [7:0] add_982969;
  wire [7:0] sel_982970;
  wire [7:0] add_982973;
  wire [7:0] sel_982974;
  wire [7:0] add_982977;
  wire [7:0] sel_982978;
  wire [7:0] add_982981;
  wire [7:0] sel_982982;
  wire [7:0] add_982985;
  wire [7:0] sel_982986;
  wire [7:0] add_982989;
  wire [7:0] sel_982990;
  wire [7:0] add_982993;
  wire [7:0] sel_982994;
  wire [7:0] add_982997;
  wire [7:0] sel_982998;
  wire [7:0] add_983001;
  wire [7:0] sel_983002;
  wire [7:0] add_983005;
  wire [7:0] sel_983006;
  wire [7:0] add_983009;
  wire [7:0] sel_983010;
  wire [7:0] add_983013;
  wire [7:0] sel_983014;
  wire [7:0] add_983017;
  wire [7:0] sel_983018;
  wire [7:0] add_983021;
  wire [7:0] sel_983022;
  wire [7:0] add_983025;
  wire [7:0] sel_983026;
  wire [7:0] add_983029;
  wire [7:0] sel_983030;
  wire [7:0] add_983033;
  wire [7:0] sel_983034;
  wire [7:0] add_983037;
  wire [7:0] sel_983038;
  wire [7:0] add_983041;
  wire [7:0] sel_983042;
  wire [7:0] add_983045;
  wire [7:0] sel_983046;
  wire [7:0] add_983049;
  wire [7:0] sel_983050;
  wire [7:0] add_983053;
  wire [7:0] sel_983054;
  wire [7:0] add_983057;
  wire [7:0] sel_983058;
  wire [7:0] add_983061;
  wire [7:0] sel_983062;
  wire [7:0] add_983065;
  wire [7:0] sel_983066;
  wire [7:0] add_983069;
  wire [7:0] sel_983070;
  wire [7:0] add_983073;
  wire [7:0] sel_983074;
  wire [7:0] add_983077;
  wire [7:0] sel_983078;
  wire [7:0] add_983081;
  wire [7:0] sel_983082;
  wire [7:0] add_983085;
  wire [7:0] sel_983086;
  wire [7:0] add_983089;
  wire [7:0] sel_983090;
  wire [7:0] add_983093;
  wire [7:0] sel_983094;
  wire [7:0] add_983097;
  wire [7:0] sel_983098;
  wire [7:0] add_983101;
  wire [7:0] sel_983102;
  wire [7:0] add_983105;
  wire [7:0] sel_983106;
  wire [7:0] add_983109;
  wire [7:0] sel_983110;
  wire [7:0] add_983113;
  wire [7:0] sel_983114;
  wire [7:0] add_983117;
  wire [7:0] sel_983118;
  wire [7:0] add_983121;
  wire [7:0] sel_983122;
  wire [7:0] add_983125;
  wire [7:0] sel_983126;
  wire [7:0] add_983129;
  wire [7:0] sel_983130;
  wire [7:0] add_983133;
  wire [7:0] sel_983134;
  wire [7:0] add_983137;
  wire [7:0] sel_983138;
  wire [7:0] add_983141;
  wire [7:0] sel_983142;
  wire [7:0] add_983145;
  wire [7:0] sel_983146;
  wire [7:0] add_983149;
  wire [7:0] sel_983150;
  wire [7:0] add_983153;
  wire [7:0] sel_983154;
  wire [7:0] add_983157;
  wire [7:0] sel_983158;
  wire [7:0] add_983161;
  wire [7:0] sel_983162;
  wire [7:0] add_983165;
  wire [7:0] sel_983166;
  wire [7:0] add_983169;
  wire [7:0] sel_983170;
  wire [7:0] add_983173;
  wire [7:0] sel_983174;
  wire [7:0] add_983177;
  wire [7:0] sel_983178;
  wire [7:0] add_983181;
  wire [7:0] sel_983182;
  wire [7:0] add_983185;
  wire [7:0] sel_983186;
  wire [7:0] add_983189;
  wire [7:0] sel_983190;
  wire [7:0] add_983193;
  wire [7:0] sel_983194;
  wire [7:0] add_983197;
  wire [7:0] sel_983198;
  wire [7:0] add_983201;
  wire [7:0] sel_983202;
  wire [7:0] add_983205;
  wire [7:0] sel_983206;
  wire [7:0] add_983209;
  wire [7:0] sel_983210;
  wire [7:0] add_983213;
  wire [7:0] sel_983214;
  wire [7:0] add_983217;
  wire [7:0] sel_983218;
  wire [7:0] add_983221;
  wire [7:0] sel_983222;
  wire [7:0] add_983225;
  wire [7:0] sel_983226;
  wire [7:0] add_983229;
  wire [7:0] sel_983230;
  wire [7:0] add_983233;
  wire [7:0] sel_983234;
  wire [7:0] add_983237;
  wire [7:0] sel_983238;
  wire [7:0] add_983241;
  wire [7:0] sel_983242;
  wire [7:0] add_983245;
  wire [7:0] sel_983246;
  wire [7:0] add_983249;
  wire [7:0] sel_983250;
  wire [7:0] add_983253;
  wire [7:0] sel_983254;
  wire [7:0] add_983257;
  wire [7:0] sel_983258;
  wire [7:0] add_983262;
  wire [15:0] array_index_983263;
  wire [7:0] sel_983264;
  wire [7:0] add_983267;
  wire [7:0] sel_983268;
  wire [7:0] add_983271;
  wire [7:0] sel_983272;
  wire [7:0] add_983275;
  wire [7:0] sel_983276;
  wire [7:0] add_983279;
  wire [7:0] sel_983280;
  wire [7:0] add_983283;
  wire [7:0] sel_983284;
  wire [7:0] add_983287;
  wire [7:0] sel_983288;
  wire [7:0] add_983291;
  wire [7:0] sel_983292;
  wire [7:0] add_983295;
  wire [7:0] sel_983296;
  wire [7:0] add_983299;
  wire [7:0] sel_983300;
  wire [7:0] add_983303;
  wire [7:0] sel_983304;
  wire [7:0] add_983307;
  wire [7:0] sel_983308;
  wire [7:0] add_983311;
  wire [7:0] sel_983312;
  wire [7:0] add_983315;
  wire [7:0] sel_983316;
  wire [7:0] add_983319;
  wire [7:0] sel_983320;
  wire [7:0] add_983323;
  wire [7:0] sel_983324;
  wire [7:0] add_983327;
  wire [7:0] sel_983328;
  wire [7:0] add_983331;
  wire [7:0] sel_983332;
  wire [7:0] add_983335;
  wire [7:0] sel_983336;
  wire [7:0] add_983339;
  wire [7:0] sel_983340;
  wire [7:0] add_983343;
  wire [7:0] sel_983344;
  wire [7:0] add_983347;
  wire [7:0] sel_983348;
  wire [7:0] add_983351;
  wire [7:0] sel_983352;
  wire [7:0] add_983355;
  wire [7:0] sel_983356;
  wire [7:0] add_983359;
  wire [7:0] sel_983360;
  wire [7:0] add_983363;
  wire [7:0] sel_983364;
  wire [7:0] add_983367;
  wire [7:0] sel_983368;
  wire [7:0] add_983371;
  wire [7:0] sel_983372;
  wire [7:0] add_983375;
  wire [7:0] sel_983376;
  wire [7:0] add_983379;
  wire [7:0] sel_983380;
  wire [7:0] add_983383;
  wire [7:0] sel_983384;
  wire [7:0] add_983387;
  wire [7:0] sel_983388;
  wire [7:0] add_983391;
  wire [7:0] sel_983392;
  wire [7:0] add_983395;
  wire [7:0] sel_983396;
  wire [7:0] add_983399;
  wire [7:0] sel_983400;
  wire [7:0] add_983403;
  wire [7:0] sel_983404;
  wire [7:0] add_983407;
  wire [7:0] sel_983408;
  wire [7:0] add_983411;
  wire [7:0] sel_983412;
  wire [7:0] add_983415;
  wire [7:0] sel_983416;
  wire [7:0] add_983419;
  wire [7:0] sel_983420;
  wire [7:0] add_983423;
  wire [7:0] sel_983424;
  wire [7:0] add_983427;
  wire [7:0] sel_983428;
  wire [7:0] add_983431;
  wire [7:0] sel_983432;
  wire [7:0] add_983435;
  wire [7:0] sel_983436;
  wire [7:0] add_983439;
  wire [7:0] sel_983440;
  wire [7:0] add_983443;
  wire [7:0] sel_983444;
  wire [7:0] add_983447;
  wire [7:0] sel_983448;
  wire [7:0] add_983451;
  wire [7:0] sel_983452;
  wire [7:0] add_983455;
  wire [7:0] sel_983456;
  wire [7:0] add_983459;
  wire [7:0] sel_983460;
  wire [7:0] add_983463;
  wire [7:0] sel_983464;
  wire [7:0] add_983467;
  wire [7:0] sel_983468;
  wire [7:0] add_983471;
  wire [7:0] sel_983472;
  wire [7:0] add_983475;
  wire [7:0] sel_983476;
  wire [7:0] add_983479;
  wire [7:0] sel_983480;
  wire [7:0] add_983483;
  wire [7:0] sel_983484;
  wire [7:0] add_983487;
  wire [7:0] sel_983488;
  wire [7:0] add_983491;
  wire [7:0] sel_983492;
  wire [7:0] add_983495;
  wire [7:0] sel_983496;
  wire [7:0] add_983499;
  wire [7:0] sel_983500;
  wire [7:0] add_983503;
  wire [7:0] sel_983504;
  wire [7:0] add_983507;
  wire [7:0] sel_983508;
  wire [7:0] add_983511;
  wire [7:0] sel_983512;
  wire [7:0] add_983515;
  wire [7:0] sel_983516;
  wire [7:0] add_983519;
  wire [7:0] sel_983520;
  wire [7:0] add_983523;
  wire [7:0] sel_983524;
  wire [7:0] add_983527;
  wire [7:0] sel_983528;
  wire [7:0] add_983531;
  wire [7:0] sel_983532;
  wire [7:0] add_983535;
  wire [7:0] sel_983536;
  wire [7:0] add_983539;
  wire [7:0] sel_983540;
  wire [7:0] add_983543;
  wire [7:0] sel_983544;
  wire [7:0] add_983547;
  wire [7:0] sel_983548;
  wire [7:0] add_983551;
  wire [7:0] sel_983552;
  wire [7:0] add_983555;
  wire [7:0] sel_983556;
  wire [7:0] add_983559;
  wire [7:0] sel_983560;
  wire [7:0] add_983563;
  wire [7:0] sel_983564;
  wire [7:0] add_983567;
  wire [7:0] sel_983568;
  wire [7:0] add_983571;
  wire [7:0] sel_983572;
  wire [7:0] add_983575;
  wire [7:0] sel_983576;
  wire [7:0] add_983579;
  wire [7:0] sel_983580;
  wire [7:0] add_983583;
  wire [7:0] sel_983584;
  wire [7:0] add_983587;
  wire [7:0] sel_983588;
  wire [7:0] add_983591;
  wire [7:0] sel_983592;
  wire [7:0] add_983595;
  wire [7:0] sel_983596;
  wire [7:0] add_983599;
  wire [7:0] sel_983600;
  wire [7:0] add_983603;
  wire [7:0] sel_983604;
  wire [7:0] add_983607;
  wire [7:0] sel_983608;
  wire [7:0] add_983611;
  wire [7:0] sel_983612;
  wire [7:0] add_983615;
  wire [7:0] sel_983616;
  wire [7:0] add_983619;
  wire [7:0] sel_983620;
  wire [7:0] add_983623;
  wire [7:0] sel_983624;
  wire [7:0] add_983627;
  wire [7:0] sel_983628;
  wire [7:0] add_983631;
  wire [7:0] sel_983632;
  wire [7:0] add_983635;
  wire [7:0] sel_983636;
  wire [7:0] add_983639;
  wire [7:0] sel_983640;
  wire [7:0] add_983643;
  wire [7:0] sel_983644;
  wire [7:0] add_983647;
  wire [7:0] sel_983648;
  wire [7:0] add_983651;
  wire [7:0] sel_983652;
  wire [7:0] add_983655;
  wire [7:0] sel_983656;
  wire [7:0] add_983659;
  wire [7:0] sel_983660;
  wire [7:0] add_983664;
  wire [15:0] array_index_983665;
  wire [7:0] sel_983666;
  wire [7:0] add_983669;
  wire [7:0] sel_983670;
  wire [7:0] add_983673;
  wire [7:0] sel_983674;
  wire [7:0] add_983677;
  wire [7:0] sel_983678;
  wire [7:0] add_983681;
  wire [7:0] sel_983682;
  wire [7:0] add_983685;
  wire [7:0] sel_983686;
  wire [7:0] add_983689;
  wire [7:0] sel_983690;
  wire [7:0] add_983693;
  wire [7:0] sel_983694;
  wire [7:0] add_983697;
  wire [7:0] sel_983698;
  wire [7:0] add_983701;
  wire [7:0] sel_983702;
  wire [7:0] add_983705;
  wire [7:0] sel_983706;
  wire [7:0] add_983709;
  wire [7:0] sel_983710;
  wire [7:0] add_983713;
  wire [7:0] sel_983714;
  wire [7:0] add_983717;
  wire [7:0] sel_983718;
  wire [7:0] add_983721;
  wire [7:0] sel_983722;
  wire [7:0] add_983725;
  wire [7:0] sel_983726;
  wire [7:0] add_983729;
  wire [7:0] sel_983730;
  wire [7:0] add_983733;
  wire [7:0] sel_983734;
  wire [7:0] add_983737;
  wire [7:0] sel_983738;
  wire [7:0] add_983741;
  wire [7:0] sel_983742;
  wire [7:0] add_983745;
  wire [7:0] sel_983746;
  wire [7:0] add_983749;
  wire [7:0] sel_983750;
  wire [7:0] add_983753;
  wire [7:0] sel_983754;
  wire [7:0] add_983757;
  wire [7:0] sel_983758;
  wire [7:0] add_983761;
  wire [7:0] sel_983762;
  wire [7:0] add_983765;
  wire [7:0] sel_983766;
  wire [7:0] add_983769;
  wire [7:0] sel_983770;
  wire [7:0] add_983773;
  wire [7:0] sel_983774;
  wire [7:0] add_983777;
  wire [7:0] sel_983778;
  wire [7:0] add_983781;
  wire [7:0] sel_983782;
  wire [7:0] add_983785;
  wire [7:0] sel_983786;
  wire [7:0] add_983789;
  wire [7:0] sel_983790;
  wire [7:0] add_983793;
  wire [7:0] sel_983794;
  wire [7:0] add_983797;
  wire [7:0] sel_983798;
  wire [7:0] add_983801;
  wire [7:0] sel_983802;
  wire [7:0] add_983805;
  wire [7:0] sel_983806;
  wire [7:0] add_983809;
  wire [7:0] sel_983810;
  wire [7:0] add_983813;
  wire [7:0] sel_983814;
  wire [7:0] add_983817;
  wire [7:0] sel_983818;
  wire [7:0] add_983821;
  wire [7:0] sel_983822;
  wire [7:0] add_983825;
  wire [7:0] sel_983826;
  wire [7:0] add_983829;
  wire [7:0] sel_983830;
  wire [7:0] add_983833;
  wire [7:0] sel_983834;
  wire [7:0] add_983837;
  wire [7:0] sel_983838;
  wire [7:0] add_983841;
  wire [7:0] sel_983842;
  wire [7:0] add_983845;
  wire [7:0] sel_983846;
  wire [7:0] add_983849;
  wire [7:0] sel_983850;
  wire [7:0] add_983853;
  wire [7:0] sel_983854;
  wire [7:0] add_983857;
  wire [7:0] sel_983858;
  wire [7:0] add_983861;
  wire [7:0] sel_983862;
  wire [7:0] add_983865;
  wire [7:0] sel_983866;
  wire [7:0] add_983869;
  wire [7:0] sel_983870;
  wire [7:0] add_983873;
  wire [7:0] sel_983874;
  wire [7:0] add_983877;
  wire [7:0] sel_983878;
  wire [7:0] add_983881;
  wire [7:0] sel_983882;
  wire [7:0] add_983885;
  wire [7:0] sel_983886;
  wire [7:0] add_983889;
  wire [7:0] sel_983890;
  wire [7:0] add_983893;
  wire [7:0] sel_983894;
  wire [7:0] add_983897;
  wire [7:0] sel_983898;
  wire [7:0] add_983901;
  wire [7:0] sel_983902;
  wire [7:0] add_983905;
  wire [7:0] sel_983906;
  wire [7:0] add_983909;
  wire [7:0] sel_983910;
  wire [7:0] add_983913;
  wire [7:0] sel_983914;
  wire [7:0] add_983917;
  wire [7:0] sel_983918;
  wire [7:0] add_983921;
  wire [7:0] sel_983922;
  wire [7:0] add_983925;
  wire [7:0] sel_983926;
  wire [7:0] add_983929;
  wire [7:0] sel_983930;
  wire [7:0] add_983933;
  wire [7:0] sel_983934;
  wire [7:0] add_983937;
  wire [7:0] sel_983938;
  wire [7:0] add_983941;
  wire [7:0] sel_983942;
  wire [7:0] add_983945;
  wire [7:0] sel_983946;
  wire [7:0] add_983949;
  wire [7:0] sel_983950;
  wire [7:0] add_983953;
  wire [7:0] sel_983954;
  wire [7:0] add_983957;
  wire [7:0] sel_983958;
  wire [7:0] add_983961;
  wire [7:0] sel_983962;
  wire [7:0] add_983965;
  wire [7:0] sel_983966;
  wire [7:0] add_983969;
  wire [7:0] sel_983970;
  wire [7:0] add_983973;
  wire [7:0] sel_983974;
  wire [7:0] add_983977;
  wire [7:0] sel_983978;
  wire [7:0] add_983981;
  wire [7:0] sel_983982;
  wire [7:0] add_983985;
  wire [7:0] sel_983986;
  wire [7:0] add_983989;
  wire [7:0] sel_983990;
  wire [7:0] add_983993;
  wire [7:0] sel_983994;
  wire [7:0] add_983997;
  wire [7:0] sel_983998;
  wire [7:0] add_984001;
  wire [7:0] sel_984002;
  wire [7:0] add_984005;
  wire [7:0] sel_984006;
  wire [7:0] add_984009;
  wire [7:0] sel_984010;
  wire [7:0] add_984013;
  wire [7:0] sel_984014;
  wire [7:0] add_984017;
  wire [7:0] sel_984018;
  wire [7:0] add_984021;
  wire [7:0] sel_984022;
  wire [7:0] add_984025;
  wire [7:0] sel_984026;
  wire [7:0] add_984029;
  wire [7:0] sel_984030;
  wire [7:0] add_984033;
  wire [7:0] sel_984034;
  wire [7:0] add_984037;
  wire [7:0] sel_984038;
  wire [7:0] add_984041;
  wire [7:0] sel_984042;
  wire [7:0] add_984045;
  wire [7:0] sel_984046;
  wire [7:0] add_984049;
  wire [7:0] sel_984050;
  wire [7:0] add_984053;
  wire [7:0] sel_984054;
  wire [7:0] add_984057;
  wire [7:0] sel_984058;
  wire [7:0] add_984061;
  wire [7:0] sel_984062;
  wire [7:0] add_984066;
  wire [15:0] array_index_984067;
  wire [7:0] sel_984068;
  wire [7:0] add_984071;
  wire [7:0] sel_984072;
  wire [7:0] add_984075;
  wire [7:0] sel_984076;
  wire [7:0] add_984079;
  wire [7:0] sel_984080;
  wire [7:0] add_984083;
  wire [7:0] sel_984084;
  wire [7:0] add_984087;
  wire [7:0] sel_984088;
  wire [7:0] add_984091;
  wire [7:0] sel_984092;
  wire [7:0] add_984095;
  wire [7:0] sel_984096;
  wire [7:0] add_984099;
  wire [7:0] sel_984100;
  wire [7:0] add_984103;
  wire [7:0] sel_984104;
  wire [7:0] add_984107;
  wire [7:0] sel_984108;
  wire [7:0] add_984111;
  wire [7:0] sel_984112;
  wire [7:0] add_984115;
  wire [7:0] sel_984116;
  wire [7:0] add_984119;
  wire [7:0] sel_984120;
  wire [7:0] add_984123;
  wire [7:0] sel_984124;
  wire [7:0] add_984127;
  wire [7:0] sel_984128;
  wire [7:0] add_984131;
  wire [7:0] sel_984132;
  wire [7:0] add_984135;
  wire [7:0] sel_984136;
  wire [7:0] add_984139;
  wire [7:0] sel_984140;
  wire [7:0] add_984143;
  wire [7:0] sel_984144;
  wire [7:0] add_984147;
  wire [7:0] sel_984148;
  wire [7:0] add_984151;
  wire [7:0] sel_984152;
  wire [7:0] add_984155;
  wire [7:0] sel_984156;
  wire [7:0] add_984159;
  wire [7:0] sel_984160;
  wire [7:0] add_984163;
  wire [7:0] sel_984164;
  wire [7:0] add_984167;
  wire [7:0] sel_984168;
  wire [7:0] add_984171;
  wire [7:0] sel_984172;
  wire [7:0] add_984175;
  wire [7:0] sel_984176;
  wire [7:0] add_984179;
  wire [7:0] sel_984180;
  wire [7:0] add_984183;
  wire [7:0] sel_984184;
  wire [7:0] add_984187;
  wire [7:0] sel_984188;
  wire [7:0] add_984191;
  wire [7:0] sel_984192;
  wire [7:0] add_984195;
  wire [7:0] sel_984196;
  wire [7:0] add_984199;
  wire [7:0] sel_984200;
  wire [7:0] add_984203;
  wire [7:0] sel_984204;
  wire [7:0] add_984207;
  wire [7:0] sel_984208;
  wire [7:0] add_984211;
  wire [7:0] sel_984212;
  wire [7:0] add_984215;
  wire [7:0] sel_984216;
  wire [7:0] add_984219;
  wire [7:0] sel_984220;
  wire [7:0] add_984223;
  wire [7:0] sel_984224;
  wire [7:0] add_984227;
  wire [7:0] sel_984228;
  wire [7:0] add_984231;
  wire [7:0] sel_984232;
  wire [7:0] add_984235;
  wire [7:0] sel_984236;
  wire [7:0] add_984239;
  wire [7:0] sel_984240;
  wire [7:0] add_984243;
  wire [7:0] sel_984244;
  wire [7:0] add_984247;
  wire [7:0] sel_984248;
  wire [7:0] add_984251;
  wire [7:0] sel_984252;
  wire [7:0] add_984255;
  wire [7:0] sel_984256;
  wire [7:0] add_984259;
  wire [7:0] sel_984260;
  wire [7:0] add_984263;
  wire [7:0] sel_984264;
  wire [7:0] add_984267;
  wire [7:0] sel_984268;
  wire [7:0] add_984271;
  wire [7:0] sel_984272;
  wire [7:0] add_984275;
  wire [7:0] sel_984276;
  wire [7:0] add_984279;
  wire [7:0] sel_984280;
  wire [7:0] add_984283;
  wire [7:0] sel_984284;
  wire [7:0] add_984287;
  wire [7:0] sel_984288;
  wire [7:0] add_984291;
  wire [7:0] sel_984292;
  wire [7:0] add_984295;
  wire [7:0] sel_984296;
  wire [7:0] add_984299;
  wire [7:0] sel_984300;
  wire [7:0] add_984303;
  wire [7:0] sel_984304;
  wire [7:0] add_984307;
  wire [7:0] sel_984308;
  wire [7:0] add_984311;
  wire [7:0] sel_984312;
  wire [7:0] add_984315;
  wire [7:0] sel_984316;
  wire [7:0] add_984319;
  wire [7:0] sel_984320;
  wire [7:0] add_984323;
  wire [7:0] sel_984324;
  wire [7:0] add_984327;
  wire [7:0] sel_984328;
  wire [7:0] add_984331;
  wire [7:0] sel_984332;
  wire [7:0] add_984335;
  wire [7:0] sel_984336;
  wire [7:0] add_984339;
  wire [7:0] sel_984340;
  wire [7:0] add_984343;
  wire [7:0] sel_984344;
  wire [7:0] add_984347;
  wire [7:0] sel_984348;
  wire [7:0] add_984351;
  wire [7:0] sel_984352;
  wire [7:0] add_984355;
  wire [7:0] sel_984356;
  wire [7:0] add_984359;
  wire [7:0] sel_984360;
  wire [7:0] add_984363;
  wire [7:0] sel_984364;
  wire [7:0] add_984367;
  wire [7:0] sel_984368;
  wire [7:0] add_984371;
  wire [7:0] sel_984372;
  wire [7:0] add_984375;
  wire [7:0] sel_984376;
  wire [7:0] add_984379;
  wire [7:0] sel_984380;
  wire [7:0] add_984383;
  wire [7:0] sel_984384;
  wire [7:0] add_984387;
  wire [7:0] sel_984388;
  wire [7:0] add_984391;
  wire [7:0] sel_984392;
  wire [7:0] add_984395;
  wire [7:0] sel_984396;
  wire [7:0] add_984399;
  wire [7:0] sel_984400;
  wire [7:0] add_984403;
  wire [7:0] sel_984404;
  wire [7:0] add_984407;
  wire [7:0] sel_984408;
  wire [7:0] add_984411;
  wire [7:0] sel_984412;
  wire [7:0] add_984415;
  wire [7:0] sel_984416;
  wire [7:0] add_984419;
  wire [7:0] sel_984420;
  wire [7:0] add_984423;
  wire [7:0] sel_984424;
  wire [7:0] add_984427;
  wire [7:0] sel_984428;
  wire [7:0] add_984431;
  wire [7:0] sel_984432;
  wire [7:0] add_984435;
  wire [7:0] sel_984436;
  wire [7:0] add_984439;
  wire [7:0] sel_984440;
  wire [7:0] add_984443;
  wire [7:0] sel_984444;
  wire [7:0] add_984447;
  wire [7:0] sel_984448;
  wire [7:0] add_984451;
  wire [7:0] sel_984452;
  wire [7:0] add_984455;
  wire [7:0] sel_984456;
  wire [7:0] add_984459;
  wire [7:0] sel_984460;
  wire [7:0] add_984463;
  wire [7:0] sel_984464;
  wire [7:0] add_984468;
  wire [15:0] array_index_984469;
  wire [7:0] sel_984470;
  wire [7:0] add_984473;
  wire [7:0] sel_984474;
  wire [7:0] add_984477;
  wire [7:0] sel_984478;
  wire [7:0] add_984481;
  wire [7:0] sel_984482;
  wire [7:0] add_984485;
  wire [7:0] sel_984486;
  wire [7:0] add_984489;
  wire [7:0] sel_984490;
  wire [7:0] add_984493;
  wire [7:0] sel_984494;
  wire [7:0] add_984497;
  wire [7:0] sel_984498;
  wire [7:0] add_984501;
  wire [7:0] sel_984502;
  wire [7:0] add_984505;
  wire [7:0] sel_984506;
  wire [7:0] add_984509;
  wire [7:0] sel_984510;
  wire [7:0] add_984513;
  wire [7:0] sel_984514;
  wire [7:0] add_984517;
  wire [7:0] sel_984518;
  wire [7:0] add_984521;
  wire [7:0] sel_984522;
  wire [7:0] add_984525;
  wire [7:0] sel_984526;
  wire [7:0] add_984529;
  wire [7:0] sel_984530;
  wire [7:0] add_984533;
  wire [7:0] sel_984534;
  wire [7:0] add_984537;
  wire [7:0] sel_984538;
  wire [7:0] add_984541;
  wire [7:0] sel_984542;
  wire [7:0] add_984545;
  wire [7:0] sel_984546;
  wire [7:0] add_984549;
  wire [7:0] sel_984550;
  wire [7:0] add_984553;
  wire [7:0] sel_984554;
  wire [7:0] add_984557;
  wire [7:0] sel_984558;
  wire [7:0] add_984561;
  wire [7:0] sel_984562;
  wire [7:0] add_984565;
  wire [7:0] sel_984566;
  wire [7:0] add_984569;
  wire [7:0] sel_984570;
  wire [7:0] add_984573;
  wire [7:0] sel_984574;
  wire [7:0] add_984577;
  wire [7:0] sel_984578;
  wire [7:0] add_984581;
  wire [7:0] sel_984582;
  wire [7:0] add_984585;
  wire [7:0] sel_984586;
  wire [7:0] add_984589;
  wire [7:0] sel_984590;
  wire [7:0] add_984593;
  wire [7:0] sel_984594;
  wire [7:0] add_984597;
  wire [7:0] sel_984598;
  wire [7:0] add_984601;
  wire [7:0] sel_984602;
  wire [7:0] add_984605;
  wire [7:0] sel_984606;
  wire [7:0] add_984609;
  wire [7:0] sel_984610;
  wire [7:0] add_984613;
  wire [7:0] sel_984614;
  wire [7:0] add_984617;
  wire [7:0] sel_984618;
  wire [7:0] add_984621;
  wire [7:0] sel_984622;
  wire [7:0] add_984625;
  wire [7:0] sel_984626;
  wire [7:0] add_984629;
  wire [7:0] sel_984630;
  wire [7:0] add_984633;
  wire [7:0] sel_984634;
  wire [7:0] add_984637;
  wire [7:0] sel_984638;
  wire [7:0] add_984641;
  wire [7:0] sel_984642;
  wire [7:0] add_984645;
  wire [7:0] sel_984646;
  wire [7:0] add_984649;
  wire [7:0] sel_984650;
  wire [7:0] add_984653;
  wire [7:0] sel_984654;
  wire [7:0] add_984657;
  wire [7:0] sel_984658;
  wire [7:0] add_984661;
  wire [7:0] sel_984662;
  wire [7:0] add_984665;
  wire [7:0] sel_984666;
  wire [7:0] add_984669;
  wire [7:0] sel_984670;
  wire [7:0] add_984673;
  wire [7:0] sel_984674;
  wire [7:0] add_984677;
  wire [7:0] sel_984678;
  wire [7:0] add_984681;
  wire [7:0] sel_984682;
  wire [7:0] add_984685;
  wire [7:0] sel_984686;
  wire [7:0] add_984689;
  wire [7:0] sel_984690;
  wire [7:0] add_984693;
  wire [7:0] sel_984694;
  wire [7:0] add_984697;
  wire [7:0] sel_984698;
  wire [7:0] add_984701;
  wire [7:0] sel_984702;
  wire [7:0] add_984705;
  wire [7:0] sel_984706;
  wire [7:0] add_984709;
  wire [7:0] sel_984710;
  wire [7:0] add_984713;
  wire [7:0] sel_984714;
  wire [7:0] add_984717;
  wire [7:0] sel_984718;
  wire [7:0] add_984721;
  wire [7:0] sel_984722;
  wire [7:0] add_984725;
  wire [7:0] sel_984726;
  wire [7:0] add_984729;
  wire [7:0] sel_984730;
  wire [7:0] add_984733;
  wire [7:0] sel_984734;
  wire [7:0] add_984737;
  wire [7:0] sel_984738;
  wire [7:0] add_984741;
  wire [7:0] sel_984742;
  wire [7:0] add_984745;
  wire [7:0] sel_984746;
  wire [7:0] add_984749;
  wire [7:0] sel_984750;
  wire [7:0] add_984753;
  wire [7:0] sel_984754;
  wire [7:0] add_984757;
  wire [7:0] sel_984758;
  wire [7:0] add_984761;
  wire [7:0] sel_984762;
  wire [7:0] add_984765;
  wire [7:0] sel_984766;
  wire [7:0] add_984769;
  wire [7:0] sel_984770;
  wire [7:0] add_984773;
  wire [7:0] sel_984774;
  wire [7:0] add_984777;
  wire [7:0] sel_984778;
  wire [7:0] add_984781;
  wire [7:0] sel_984782;
  wire [7:0] add_984785;
  wire [7:0] sel_984786;
  wire [7:0] add_984789;
  wire [7:0] sel_984790;
  wire [7:0] add_984793;
  wire [7:0] sel_984794;
  wire [7:0] add_984797;
  wire [7:0] sel_984798;
  wire [7:0] add_984801;
  wire [7:0] sel_984802;
  wire [7:0] add_984805;
  wire [7:0] sel_984806;
  wire [7:0] add_984809;
  wire [7:0] sel_984810;
  wire [7:0] add_984813;
  wire [7:0] sel_984814;
  wire [7:0] add_984817;
  wire [7:0] sel_984818;
  wire [7:0] add_984821;
  wire [7:0] sel_984822;
  wire [7:0] add_984825;
  wire [7:0] sel_984826;
  wire [7:0] add_984829;
  wire [7:0] sel_984830;
  wire [7:0] add_984833;
  wire [7:0] sel_984834;
  wire [7:0] add_984837;
  wire [7:0] sel_984838;
  wire [7:0] add_984841;
  wire [7:0] sel_984842;
  wire [7:0] add_984845;
  wire [7:0] sel_984846;
  wire [7:0] add_984849;
  wire [7:0] sel_984850;
  wire [7:0] add_984853;
  wire [7:0] sel_984854;
  wire [7:0] add_984857;
  wire [7:0] sel_984858;
  wire [7:0] add_984861;
  wire [7:0] sel_984862;
  wire [7:0] add_984865;
  wire [7:0] sel_984866;
  wire [7:0] add_984870;
  wire [15:0] array_index_984871;
  wire [7:0] sel_984872;
  wire [7:0] add_984875;
  wire [7:0] sel_984876;
  wire [7:0] add_984879;
  wire [7:0] sel_984880;
  wire [7:0] add_984883;
  wire [7:0] sel_984884;
  wire [7:0] add_984887;
  wire [7:0] sel_984888;
  wire [7:0] add_984891;
  wire [7:0] sel_984892;
  wire [7:0] add_984895;
  wire [7:0] sel_984896;
  wire [7:0] add_984899;
  wire [7:0] sel_984900;
  wire [7:0] add_984903;
  wire [7:0] sel_984904;
  wire [7:0] add_984907;
  wire [7:0] sel_984908;
  wire [7:0] add_984911;
  wire [7:0] sel_984912;
  wire [7:0] add_984915;
  wire [7:0] sel_984916;
  wire [7:0] add_984919;
  wire [7:0] sel_984920;
  wire [7:0] add_984923;
  wire [7:0] sel_984924;
  wire [7:0] add_984927;
  wire [7:0] sel_984928;
  wire [7:0] add_984931;
  wire [7:0] sel_984932;
  wire [7:0] add_984935;
  wire [7:0] sel_984936;
  wire [7:0] add_984939;
  wire [7:0] sel_984940;
  wire [7:0] add_984943;
  wire [7:0] sel_984944;
  wire [7:0] add_984947;
  wire [7:0] sel_984948;
  wire [7:0] add_984951;
  wire [7:0] sel_984952;
  wire [7:0] add_984955;
  wire [7:0] sel_984956;
  wire [7:0] add_984959;
  wire [7:0] sel_984960;
  wire [7:0] add_984963;
  wire [7:0] sel_984964;
  wire [7:0] add_984967;
  wire [7:0] sel_984968;
  wire [7:0] add_984971;
  wire [7:0] sel_984972;
  wire [7:0] add_984975;
  wire [7:0] sel_984976;
  wire [7:0] add_984979;
  wire [7:0] sel_984980;
  wire [7:0] add_984983;
  wire [7:0] sel_984984;
  wire [7:0] add_984987;
  wire [7:0] sel_984988;
  wire [7:0] add_984991;
  wire [7:0] sel_984992;
  wire [7:0] add_984995;
  wire [7:0] sel_984996;
  wire [7:0] add_984999;
  wire [7:0] sel_985000;
  wire [7:0] add_985003;
  wire [7:0] sel_985004;
  wire [7:0] add_985007;
  wire [7:0] sel_985008;
  wire [7:0] add_985011;
  wire [7:0] sel_985012;
  wire [7:0] add_985015;
  wire [7:0] sel_985016;
  wire [7:0] add_985019;
  wire [7:0] sel_985020;
  wire [7:0] add_985023;
  wire [7:0] sel_985024;
  wire [7:0] add_985027;
  wire [7:0] sel_985028;
  wire [7:0] add_985031;
  wire [7:0] sel_985032;
  wire [7:0] add_985035;
  wire [7:0] sel_985036;
  wire [7:0] add_985039;
  wire [7:0] sel_985040;
  wire [7:0] add_985043;
  wire [7:0] sel_985044;
  wire [7:0] add_985047;
  wire [7:0] sel_985048;
  wire [7:0] add_985051;
  wire [7:0] sel_985052;
  wire [7:0] add_985055;
  wire [7:0] sel_985056;
  wire [7:0] add_985059;
  wire [7:0] sel_985060;
  wire [7:0] add_985063;
  wire [7:0] sel_985064;
  wire [7:0] add_985067;
  wire [7:0] sel_985068;
  wire [7:0] add_985071;
  wire [7:0] sel_985072;
  wire [7:0] add_985075;
  wire [7:0] sel_985076;
  wire [7:0] add_985079;
  wire [7:0] sel_985080;
  wire [7:0] add_985083;
  wire [7:0] sel_985084;
  wire [7:0] add_985087;
  wire [7:0] sel_985088;
  wire [7:0] add_985091;
  wire [7:0] sel_985092;
  wire [7:0] add_985095;
  wire [7:0] sel_985096;
  wire [7:0] add_985099;
  wire [7:0] sel_985100;
  wire [7:0] add_985103;
  wire [7:0] sel_985104;
  wire [7:0] add_985107;
  wire [7:0] sel_985108;
  wire [7:0] add_985111;
  wire [7:0] sel_985112;
  wire [7:0] add_985115;
  wire [7:0] sel_985116;
  wire [7:0] add_985119;
  wire [7:0] sel_985120;
  wire [7:0] add_985123;
  wire [7:0] sel_985124;
  wire [7:0] add_985127;
  wire [7:0] sel_985128;
  wire [7:0] add_985131;
  wire [7:0] sel_985132;
  wire [7:0] add_985135;
  wire [7:0] sel_985136;
  wire [7:0] add_985139;
  wire [7:0] sel_985140;
  wire [7:0] add_985143;
  wire [7:0] sel_985144;
  wire [7:0] add_985147;
  wire [7:0] sel_985148;
  wire [7:0] add_985151;
  wire [7:0] sel_985152;
  wire [7:0] add_985155;
  wire [7:0] sel_985156;
  wire [7:0] add_985159;
  wire [7:0] sel_985160;
  wire [7:0] add_985163;
  wire [7:0] sel_985164;
  wire [7:0] add_985167;
  wire [7:0] sel_985168;
  wire [7:0] add_985171;
  wire [7:0] sel_985172;
  wire [7:0] add_985175;
  wire [7:0] sel_985176;
  wire [7:0] add_985179;
  wire [7:0] sel_985180;
  wire [7:0] add_985183;
  wire [7:0] sel_985184;
  wire [7:0] add_985187;
  wire [7:0] sel_985188;
  wire [7:0] add_985191;
  wire [7:0] sel_985192;
  wire [7:0] add_985195;
  wire [7:0] sel_985196;
  wire [7:0] add_985199;
  wire [7:0] sel_985200;
  wire [7:0] add_985203;
  wire [7:0] sel_985204;
  wire [7:0] add_985207;
  wire [7:0] sel_985208;
  wire [7:0] add_985211;
  wire [7:0] sel_985212;
  wire [7:0] add_985215;
  wire [7:0] sel_985216;
  wire [7:0] add_985219;
  wire [7:0] sel_985220;
  wire [7:0] add_985223;
  wire [7:0] sel_985224;
  wire [7:0] add_985227;
  wire [7:0] sel_985228;
  wire [7:0] add_985231;
  wire [7:0] sel_985232;
  wire [7:0] add_985235;
  wire [7:0] sel_985236;
  wire [7:0] add_985239;
  wire [7:0] sel_985240;
  wire [7:0] add_985243;
  wire [7:0] sel_985244;
  wire [7:0] add_985247;
  wire [7:0] sel_985248;
  wire [7:0] add_985251;
  wire [7:0] sel_985252;
  wire [7:0] add_985255;
  wire [7:0] sel_985256;
  wire [7:0] add_985259;
  wire [7:0] sel_985260;
  wire [7:0] add_985263;
  wire [7:0] sel_985264;
  wire [7:0] add_985267;
  wire [7:0] sel_985268;
  wire [7:0] add_985272;
  wire [15:0] array_index_985273;
  wire [7:0] sel_985274;
  wire [7:0] add_985277;
  wire [7:0] sel_985278;
  wire [7:0] add_985281;
  wire [7:0] sel_985282;
  wire [7:0] add_985285;
  wire [7:0] sel_985286;
  wire [7:0] add_985289;
  wire [7:0] sel_985290;
  wire [7:0] add_985293;
  wire [7:0] sel_985294;
  wire [7:0] add_985297;
  wire [7:0] sel_985298;
  wire [7:0] add_985301;
  wire [7:0] sel_985302;
  wire [7:0] add_985305;
  wire [7:0] sel_985306;
  wire [7:0] add_985309;
  wire [7:0] sel_985310;
  wire [7:0] add_985313;
  wire [7:0] sel_985314;
  wire [7:0] add_985317;
  wire [7:0] sel_985318;
  wire [7:0] add_985321;
  wire [7:0] sel_985322;
  wire [7:0] add_985325;
  wire [7:0] sel_985326;
  wire [7:0] add_985329;
  wire [7:0] sel_985330;
  wire [7:0] add_985333;
  wire [7:0] sel_985334;
  wire [7:0] add_985337;
  wire [7:0] sel_985338;
  wire [7:0] add_985341;
  wire [7:0] sel_985342;
  wire [7:0] add_985345;
  wire [7:0] sel_985346;
  wire [7:0] add_985349;
  wire [7:0] sel_985350;
  wire [7:0] add_985353;
  wire [7:0] sel_985354;
  wire [7:0] add_985357;
  wire [7:0] sel_985358;
  wire [7:0] add_985361;
  wire [7:0] sel_985362;
  wire [7:0] add_985365;
  wire [7:0] sel_985366;
  wire [7:0] add_985369;
  wire [7:0] sel_985370;
  wire [7:0] add_985373;
  wire [7:0] sel_985374;
  wire [7:0] add_985377;
  wire [7:0] sel_985378;
  wire [7:0] add_985381;
  wire [7:0] sel_985382;
  wire [7:0] add_985385;
  wire [7:0] sel_985386;
  wire [7:0] add_985389;
  wire [7:0] sel_985390;
  wire [7:0] add_985393;
  wire [7:0] sel_985394;
  wire [7:0] add_985397;
  wire [7:0] sel_985398;
  wire [7:0] add_985401;
  wire [7:0] sel_985402;
  wire [7:0] add_985405;
  wire [7:0] sel_985406;
  wire [7:0] add_985409;
  wire [7:0] sel_985410;
  wire [7:0] add_985413;
  wire [7:0] sel_985414;
  wire [7:0] add_985417;
  wire [7:0] sel_985418;
  wire [7:0] add_985421;
  wire [7:0] sel_985422;
  wire [7:0] add_985425;
  wire [7:0] sel_985426;
  wire [7:0] add_985429;
  wire [7:0] sel_985430;
  wire [7:0] add_985433;
  wire [7:0] sel_985434;
  wire [7:0] add_985437;
  wire [7:0] sel_985438;
  wire [7:0] add_985441;
  wire [7:0] sel_985442;
  wire [7:0] add_985445;
  wire [7:0] sel_985446;
  wire [7:0] add_985449;
  wire [7:0] sel_985450;
  wire [7:0] add_985453;
  wire [7:0] sel_985454;
  wire [7:0] add_985457;
  wire [7:0] sel_985458;
  wire [7:0] add_985461;
  wire [7:0] sel_985462;
  wire [7:0] add_985465;
  wire [7:0] sel_985466;
  wire [7:0] add_985469;
  wire [7:0] sel_985470;
  wire [7:0] add_985473;
  wire [7:0] sel_985474;
  wire [7:0] add_985477;
  wire [7:0] sel_985478;
  wire [7:0] add_985481;
  wire [7:0] sel_985482;
  wire [7:0] add_985485;
  wire [7:0] sel_985486;
  wire [7:0] add_985489;
  wire [7:0] sel_985490;
  wire [7:0] add_985493;
  wire [7:0] sel_985494;
  wire [7:0] add_985497;
  wire [7:0] sel_985498;
  wire [7:0] add_985501;
  wire [7:0] sel_985502;
  wire [7:0] add_985505;
  wire [7:0] sel_985506;
  wire [7:0] add_985509;
  wire [7:0] sel_985510;
  wire [7:0] add_985513;
  wire [7:0] sel_985514;
  wire [7:0] add_985517;
  wire [7:0] sel_985518;
  wire [7:0] add_985521;
  wire [7:0] sel_985522;
  wire [7:0] add_985525;
  wire [7:0] sel_985526;
  wire [7:0] add_985529;
  wire [7:0] sel_985530;
  wire [7:0] add_985533;
  wire [7:0] sel_985534;
  wire [7:0] add_985537;
  wire [7:0] sel_985538;
  wire [7:0] add_985541;
  wire [7:0] sel_985542;
  wire [7:0] add_985545;
  wire [7:0] sel_985546;
  wire [7:0] add_985549;
  wire [7:0] sel_985550;
  wire [7:0] add_985553;
  wire [7:0] sel_985554;
  wire [7:0] add_985557;
  wire [7:0] sel_985558;
  wire [7:0] add_985561;
  wire [7:0] sel_985562;
  wire [7:0] add_985565;
  wire [7:0] sel_985566;
  wire [7:0] add_985569;
  wire [7:0] sel_985570;
  wire [7:0] add_985573;
  wire [7:0] sel_985574;
  wire [7:0] add_985577;
  wire [7:0] sel_985578;
  wire [7:0] add_985581;
  wire [7:0] sel_985582;
  wire [7:0] add_985585;
  wire [7:0] sel_985586;
  wire [7:0] add_985589;
  wire [7:0] sel_985590;
  wire [7:0] add_985593;
  wire [7:0] sel_985594;
  wire [7:0] add_985597;
  wire [7:0] sel_985598;
  wire [7:0] add_985601;
  wire [7:0] sel_985602;
  wire [7:0] add_985605;
  wire [7:0] sel_985606;
  wire [7:0] add_985609;
  wire [7:0] sel_985610;
  wire [7:0] add_985613;
  wire [7:0] sel_985614;
  wire [7:0] add_985617;
  wire [7:0] sel_985618;
  wire [7:0] add_985621;
  wire [7:0] sel_985622;
  wire [7:0] add_985625;
  wire [7:0] sel_985626;
  wire [7:0] add_985629;
  wire [7:0] sel_985630;
  wire [7:0] add_985633;
  wire [7:0] sel_985634;
  wire [7:0] add_985637;
  wire [7:0] sel_985638;
  wire [7:0] add_985641;
  wire [7:0] sel_985642;
  wire [7:0] add_985645;
  wire [7:0] sel_985646;
  wire [7:0] add_985649;
  wire [7:0] sel_985650;
  wire [7:0] add_985653;
  wire [7:0] sel_985654;
  wire [7:0] add_985657;
  wire [7:0] sel_985658;
  wire [7:0] add_985661;
  wire [7:0] sel_985662;
  wire [7:0] add_985665;
  wire [7:0] sel_985666;
  wire [7:0] add_985669;
  wire [7:0] sel_985670;
  wire [7:0] add_985674;
  wire [15:0] array_index_985675;
  wire [7:0] sel_985676;
  wire [7:0] add_985679;
  wire [7:0] sel_985680;
  wire [7:0] add_985683;
  wire [7:0] sel_985684;
  wire [7:0] add_985687;
  wire [7:0] sel_985688;
  wire [7:0] add_985691;
  wire [7:0] sel_985692;
  wire [7:0] add_985695;
  wire [7:0] sel_985696;
  wire [7:0] add_985699;
  wire [7:0] sel_985700;
  wire [7:0] add_985703;
  wire [7:0] sel_985704;
  wire [7:0] add_985707;
  wire [7:0] sel_985708;
  wire [7:0] add_985711;
  wire [7:0] sel_985712;
  wire [7:0] add_985715;
  wire [7:0] sel_985716;
  wire [7:0] add_985719;
  wire [7:0] sel_985720;
  wire [7:0] add_985723;
  wire [7:0] sel_985724;
  wire [7:0] add_985727;
  wire [7:0] sel_985728;
  wire [7:0] add_985731;
  wire [7:0] sel_985732;
  wire [7:0] add_985735;
  wire [7:0] sel_985736;
  wire [7:0] add_985739;
  wire [7:0] sel_985740;
  wire [7:0] add_985743;
  wire [7:0] sel_985744;
  wire [7:0] add_985747;
  wire [7:0] sel_985748;
  wire [7:0] add_985751;
  wire [7:0] sel_985752;
  wire [7:0] add_985755;
  wire [7:0] sel_985756;
  wire [7:0] add_985759;
  wire [7:0] sel_985760;
  wire [7:0] add_985763;
  wire [7:0] sel_985764;
  wire [7:0] add_985767;
  wire [7:0] sel_985768;
  wire [7:0] add_985771;
  wire [7:0] sel_985772;
  wire [7:0] add_985775;
  wire [7:0] sel_985776;
  wire [7:0] add_985779;
  wire [7:0] sel_985780;
  wire [7:0] add_985783;
  wire [7:0] sel_985784;
  wire [7:0] add_985787;
  wire [7:0] sel_985788;
  wire [7:0] add_985791;
  wire [7:0] sel_985792;
  wire [7:0] add_985795;
  wire [7:0] sel_985796;
  wire [7:0] add_985799;
  wire [7:0] sel_985800;
  wire [7:0] add_985803;
  wire [7:0] sel_985804;
  wire [7:0] add_985807;
  wire [7:0] sel_985808;
  wire [7:0] add_985811;
  wire [7:0] sel_985812;
  wire [7:0] add_985815;
  wire [7:0] sel_985816;
  wire [7:0] add_985819;
  wire [7:0] sel_985820;
  wire [7:0] add_985823;
  wire [7:0] sel_985824;
  wire [7:0] add_985827;
  wire [7:0] sel_985828;
  wire [7:0] add_985831;
  wire [7:0] sel_985832;
  wire [7:0] add_985835;
  wire [7:0] sel_985836;
  wire [7:0] add_985839;
  wire [7:0] sel_985840;
  wire [7:0] add_985843;
  wire [7:0] sel_985844;
  wire [7:0] add_985847;
  wire [7:0] sel_985848;
  wire [7:0] add_985851;
  wire [7:0] sel_985852;
  wire [7:0] add_985855;
  wire [7:0] sel_985856;
  wire [7:0] add_985859;
  wire [7:0] sel_985860;
  wire [7:0] add_985863;
  wire [7:0] sel_985864;
  wire [7:0] add_985867;
  wire [7:0] sel_985868;
  wire [7:0] add_985871;
  wire [7:0] sel_985872;
  wire [7:0] add_985875;
  wire [7:0] sel_985876;
  wire [7:0] add_985879;
  wire [7:0] sel_985880;
  wire [7:0] add_985883;
  wire [7:0] sel_985884;
  wire [7:0] add_985887;
  wire [7:0] sel_985888;
  wire [7:0] add_985891;
  wire [7:0] sel_985892;
  wire [7:0] add_985895;
  wire [7:0] sel_985896;
  wire [7:0] add_985899;
  wire [7:0] sel_985900;
  wire [7:0] add_985903;
  wire [7:0] sel_985904;
  wire [7:0] add_985907;
  wire [7:0] sel_985908;
  wire [7:0] add_985911;
  wire [7:0] sel_985912;
  wire [7:0] add_985915;
  wire [7:0] sel_985916;
  wire [7:0] add_985919;
  wire [7:0] sel_985920;
  wire [7:0] add_985923;
  wire [7:0] sel_985924;
  wire [7:0] add_985927;
  wire [7:0] sel_985928;
  wire [7:0] add_985931;
  wire [7:0] sel_985932;
  wire [7:0] add_985935;
  wire [7:0] sel_985936;
  wire [7:0] add_985939;
  wire [7:0] sel_985940;
  wire [7:0] add_985943;
  wire [7:0] sel_985944;
  wire [7:0] add_985947;
  wire [7:0] sel_985948;
  wire [7:0] add_985951;
  wire [7:0] sel_985952;
  wire [7:0] add_985955;
  wire [7:0] sel_985956;
  wire [7:0] add_985959;
  wire [7:0] sel_985960;
  wire [7:0] add_985963;
  wire [7:0] sel_985964;
  wire [7:0] add_985967;
  wire [7:0] sel_985968;
  wire [7:0] add_985971;
  wire [7:0] sel_985972;
  wire [7:0] add_985975;
  wire [7:0] sel_985976;
  wire [7:0] add_985979;
  wire [7:0] sel_985980;
  wire [7:0] add_985983;
  wire [7:0] sel_985984;
  wire [7:0] add_985987;
  wire [7:0] sel_985988;
  wire [7:0] add_985991;
  wire [7:0] sel_985992;
  wire [7:0] add_985995;
  wire [7:0] sel_985996;
  wire [7:0] add_985999;
  wire [7:0] sel_986000;
  wire [7:0] add_986003;
  wire [7:0] sel_986004;
  wire [7:0] add_986007;
  wire [7:0] sel_986008;
  wire [7:0] add_986011;
  wire [7:0] sel_986012;
  wire [7:0] add_986015;
  wire [7:0] sel_986016;
  wire [7:0] add_986019;
  wire [7:0] sel_986020;
  wire [7:0] add_986023;
  wire [7:0] sel_986024;
  wire [7:0] add_986027;
  wire [7:0] sel_986028;
  wire [7:0] add_986031;
  wire [7:0] sel_986032;
  wire [7:0] add_986035;
  wire [7:0] sel_986036;
  wire [7:0] add_986039;
  wire [7:0] sel_986040;
  wire [7:0] add_986043;
  wire [7:0] sel_986044;
  wire [7:0] add_986047;
  wire [7:0] sel_986048;
  wire [7:0] add_986051;
  wire [7:0] sel_986052;
  wire [7:0] add_986055;
  wire [7:0] sel_986056;
  wire [7:0] add_986059;
  wire [7:0] sel_986060;
  wire [7:0] add_986063;
  wire [7:0] sel_986064;
  wire [7:0] add_986067;
  wire [7:0] sel_986068;
  wire [7:0] add_986071;
  wire [7:0] sel_986072;
  wire [7:0] add_986076;
  wire [15:0] array_index_986077;
  wire [7:0] sel_986078;
  wire [7:0] add_986081;
  wire [7:0] sel_986082;
  wire [7:0] add_986085;
  wire [7:0] sel_986086;
  wire [7:0] add_986089;
  wire [7:0] sel_986090;
  wire [7:0] add_986093;
  wire [7:0] sel_986094;
  wire [7:0] add_986097;
  wire [7:0] sel_986098;
  wire [7:0] add_986101;
  wire [7:0] sel_986102;
  wire [7:0] add_986105;
  wire [7:0] sel_986106;
  wire [7:0] add_986109;
  wire [7:0] sel_986110;
  wire [7:0] add_986113;
  wire [7:0] sel_986114;
  wire [7:0] add_986117;
  wire [7:0] sel_986118;
  wire [7:0] add_986121;
  wire [7:0] sel_986122;
  wire [7:0] add_986125;
  wire [7:0] sel_986126;
  wire [7:0] add_986129;
  wire [7:0] sel_986130;
  wire [7:0] add_986133;
  wire [7:0] sel_986134;
  wire [7:0] add_986137;
  wire [7:0] sel_986138;
  wire [7:0] add_986141;
  wire [7:0] sel_986142;
  wire [7:0] add_986145;
  wire [7:0] sel_986146;
  wire [7:0] add_986149;
  wire [7:0] sel_986150;
  wire [7:0] add_986153;
  wire [7:0] sel_986154;
  wire [7:0] add_986157;
  wire [7:0] sel_986158;
  wire [7:0] add_986161;
  wire [7:0] sel_986162;
  wire [7:0] add_986165;
  wire [7:0] sel_986166;
  wire [7:0] add_986169;
  wire [7:0] sel_986170;
  wire [7:0] add_986173;
  wire [7:0] sel_986174;
  wire [7:0] add_986177;
  wire [7:0] sel_986178;
  wire [7:0] add_986181;
  wire [7:0] sel_986182;
  wire [7:0] add_986185;
  wire [7:0] sel_986186;
  wire [7:0] add_986189;
  wire [7:0] sel_986190;
  wire [7:0] add_986193;
  wire [7:0] sel_986194;
  wire [7:0] add_986197;
  wire [7:0] sel_986198;
  wire [7:0] add_986201;
  wire [7:0] sel_986202;
  wire [7:0] add_986205;
  wire [7:0] sel_986206;
  wire [7:0] add_986209;
  wire [7:0] sel_986210;
  wire [7:0] add_986213;
  wire [7:0] sel_986214;
  wire [7:0] add_986217;
  wire [7:0] sel_986218;
  wire [7:0] add_986221;
  wire [7:0] sel_986222;
  wire [7:0] add_986225;
  wire [7:0] sel_986226;
  wire [7:0] add_986229;
  wire [7:0] sel_986230;
  wire [7:0] add_986233;
  wire [7:0] sel_986234;
  wire [7:0] add_986237;
  wire [7:0] sel_986238;
  wire [7:0] add_986241;
  wire [7:0] sel_986242;
  wire [7:0] add_986245;
  wire [7:0] sel_986246;
  wire [7:0] add_986249;
  wire [7:0] sel_986250;
  wire [7:0] add_986253;
  wire [7:0] sel_986254;
  wire [7:0] add_986257;
  wire [7:0] sel_986258;
  wire [7:0] add_986261;
  wire [7:0] sel_986262;
  wire [7:0] add_986265;
  wire [7:0] sel_986266;
  wire [7:0] add_986269;
  wire [7:0] sel_986270;
  wire [7:0] add_986273;
  wire [7:0] sel_986274;
  wire [7:0] add_986277;
  wire [7:0] sel_986278;
  wire [7:0] add_986281;
  wire [7:0] sel_986282;
  wire [7:0] add_986285;
  wire [7:0] sel_986286;
  wire [7:0] add_986289;
  wire [7:0] sel_986290;
  wire [7:0] add_986293;
  wire [7:0] sel_986294;
  wire [7:0] add_986297;
  wire [7:0] sel_986298;
  wire [7:0] add_986301;
  wire [7:0] sel_986302;
  wire [7:0] add_986305;
  wire [7:0] sel_986306;
  wire [7:0] add_986309;
  wire [7:0] sel_986310;
  wire [7:0] add_986313;
  wire [7:0] sel_986314;
  wire [7:0] add_986317;
  wire [7:0] sel_986318;
  wire [7:0] add_986321;
  wire [7:0] sel_986322;
  wire [7:0] add_986325;
  wire [7:0] sel_986326;
  wire [7:0] add_986329;
  wire [7:0] sel_986330;
  wire [7:0] add_986333;
  wire [7:0] sel_986334;
  wire [7:0] add_986337;
  wire [7:0] sel_986338;
  wire [7:0] add_986341;
  wire [7:0] sel_986342;
  wire [7:0] add_986345;
  wire [7:0] sel_986346;
  wire [7:0] add_986349;
  wire [7:0] sel_986350;
  wire [7:0] add_986353;
  wire [7:0] sel_986354;
  wire [7:0] add_986357;
  wire [7:0] sel_986358;
  wire [7:0] add_986361;
  wire [7:0] sel_986362;
  wire [7:0] add_986365;
  wire [7:0] sel_986366;
  wire [7:0] add_986369;
  wire [7:0] sel_986370;
  wire [7:0] add_986373;
  wire [7:0] sel_986374;
  wire [7:0] add_986377;
  wire [7:0] sel_986378;
  wire [7:0] add_986381;
  wire [7:0] sel_986382;
  wire [7:0] add_986385;
  wire [7:0] sel_986386;
  wire [7:0] add_986389;
  wire [7:0] sel_986390;
  wire [7:0] add_986393;
  wire [7:0] sel_986394;
  wire [7:0] add_986397;
  wire [7:0] sel_986398;
  wire [7:0] add_986401;
  wire [7:0] sel_986402;
  wire [7:0] add_986405;
  wire [7:0] sel_986406;
  wire [7:0] add_986409;
  wire [7:0] sel_986410;
  wire [7:0] add_986413;
  wire [7:0] sel_986414;
  wire [7:0] add_986417;
  wire [7:0] sel_986418;
  wire [7:0] add_986421;
  wire [7:0] sel_986422;
  wire [7:0] add_986425;
  wire [7:0] sel_986426;
  wire [7:0] add_986429;
  wire [7:0] sel_986430;
  wire [7:0] add_986433;
  wire [7:0] sel_986434;
  wire [7:0] add_986437;
  wire [7:0] sel_986438;
  wire [7:0] add_986441;
  wire [7:0] sel_986442;
  wire [7:0] add_986445;
  wire [7:0] sel_986446;
  wire [7:0] add_986449;
  wire [7:0] sel_986450;
  wire [7:0] add_986453;
  wire [7:0] sel_986454;
  wire [7:0] add_986457;
  wire [7:0] sel_986458;
  wire [7:0] add_986461;
  wire [7:0] sel_986462;
  wire [7:0] add_986465;
  wire [7:0] sel_986466;
  wire [7:0] add_986469;
  wire [7:0] sel_986470;
  wire [7:0] add_986473;
  wire [7:0] sel_986474;
  wire [7:0] add_986478;
  wire [15:0] array_index_986479;
  wire [7:0] sel_986480;
  wire [7:0] add_986483;
  wire [7:0] sel_986484;
  wire [7:0] add_986487;
  wire [7:0] sel_986488;
  wire [7:0] add_986491;
  wire [7:0] sel_986492;
  wire [7:0] add_986495;
  wire [7:0] sel_986496;
  wire [7:0] add_986499;
  wire [7:0] sel_986500;
  wire [7:0] add_986503;
  wire [7:0] sel_986504;
  wire [7:0] add_986507;
  wire [7:0] sel_986508;
  wire [7:0] add_986511;
  wire [7:0] sel_986512;
  wire [7:0] add_986515;
  wire [7:0] sel_986516;
  wire [7:0] add_986519;
  wire [7:0] sel_986520;
  wire [7:0] add_986523;
  wire [7:0] sel_986524;
  wire [7:0] add_986527;
  wire [7:0] sel_986528;
  wire [7:0] add_986531;
  wire [7:0] sel_986532;
  wire [7:0] add_986535;
  wire [7:0] sel_986536;
  wire [7:0] add_986539;
  wire [7:0] sel_986540;
  wire [7:0] add_986543;
  wire [7:0] sel_986544;
  wire [7:0] add_986547;
  wire [7:0] sel_986548;
  wire [7:0] add_986551;
  wire [7:0] sel_986552;
  wire [7:0] add_986555;
  wire [7:0] sel_986556;
  wire [7:0] add_986559;
  wire [7:0] sel_986560;
  wire [7:0] add_986563;
  wire [7:0] sel_986564;
  wire [7:0] add_986567;
  wire [7:0] sel_986568;
  wire [7:0] add_986571;
  wire [7:0] sel_986572;
  wire [7:0] add_986575;
  wire [7:0] sel_986576;
  wire [7:0] add_986579;
  wire [7:0] sel_986580;
  wire [7:0] add_986583;
  wire [7:0] sel_986584;
  wire [7:0] add_986587;
  wire [7:0] sel_986588;
  wire [7:0] add_986591;
  wire [7:0] sel_986592;
  wire [7:0] add_986595;
  wire [7:0] sel_986596;
  wire [7:0] add_986599;
  wire [7:0] sel_986600;
  wire [7:0] add_986603;
  wire [7:0] sel_986604;
  wire [7:0] add_986607;
  wire [7:0] sel_986608;
  wire [7:0] add_986611;
  wire [7:0] sel_986612;
  wire [7:0] add_986615;
  wire [7:0] sel_986616;
  wire [7:0] add_986619;
  wire [7:0] sel_986620;
  wire [7:0] add_986623;
  wire [7:0] sel_986624;
  wire [7:0] add_986627;
  wire [7:0] sel_986628;
  wire [7:0] add_986631;
  wire [7:0] sel_986632;
  wire [7:0] add_986635;
  wire [7:0] sel_986636;
  wire [7:0] add_986639;
  wire [7:0] sel_986640;
  wire [7:0] add_986643;
  wire [7:0] sel_986644;
  wire [7:0] add_986647;
  wire [7:0] sel_986648;
  wire [7:0] add_986651;
  wire [7:0] sel_986652;
  wire [7:0] add_986655;
  wire [7:0] sel_986656;
  wire [7:0] add_986659;
  wire [7:0] sel_986660;
  wire [7:0] add_986663;
  wire [7:0] sel_986664;
  wire [7:0] add_986667;
  wire [7:0] sel_986668;
  wire [7:0] add_986671;
  wire [7:0] sel_986672;
  wire [7:0] add_986675;
  wire [7:0] sel_986676;
  wire [7:0] add_986679;
  wire [7:0] sel_986680;
  wire [7:0] add_986683;
  wire [7:0] sel_986684;
  wire [7:0] add_986687;
  wire [7:0] sel_986688;
  wire [7:0] add_986691;
  wire [7:0] sel_986692;
  wire [7:0] add_986695;
  wire [7:0] sel_986696;
  wire [7:0] add_986699;
  wire [7:0] sel_986700;
  wire [7:0] add_986703;
  wire [7:0] sel_986704;
  wire [7:0] add_986707;
  wire [7:0] sel_986708;
  wire [7:0] add_986711;
  wire [7:0] sel_986712;
  wire [7:0] add_986715;
  wire [7:0] sel_986716;
  wire [7:0] add_986719;
  wire [7:0] sel_986720;
  wire [7:0] add_986723;
  wire [7:0] sel_986724;
  wire [7:0] add_986727;
  wire [7:0] sel_986728;
  wire [7:0] add_986731;
  wire [7:0] sel_986732;
  wire [7:0] add_986735;
  wire [7:0] sel_986736;
  wire [7:0] add_986739;
  wire [7:0] sel_986740;
  wire [7:0] add_986743;
  wire [7:0] sel_986744;
  wire [7:0] add_986747;
  wire [7:0] sel_986748;
  wire [7:0] add_986751;
  wire [7:0] sel_986752;
  wire [7:0] add_986755;
  wire [7:0] sel_986756;
  wire [7:0] add_986759;
  wire [7:0] sel_986760;
  wire [7:0] add_986763;
  wire [7:0] sel_986764;
  wire [7:0] add_986767;
  wire [7:0] sel_986768;
  wire [7:0] add_986771;
  wire [7:0] sel_986772;
  wire [7:0] add_986775;
  wire [7:0] sel_986776;
  wire [7:0] add_986779;
  wire [7:0] sel_986780;
  wire [7:0] add_986783;
  wire [7:0] sel_986784;
  wire [7:0] add_986787;
  wire [7:0] sel_986788;
  wire [7:0] add_986791;
  wire [7:0] sel_986792;
  wire [7:0] add_986795;
  wire [7:0] sel_986796;
  wire [7:0] add_986799;
  wire [7:0] sel_986800;
  wire [7:0] add_986803;
  wire [7:0] sel_986804;
  wire [7:0] add_986807;
  wire [7:0] sel_986808;
  wire [7:0] add_986811;
  wire [7:0] sel_986812;
  wire [7:0] add_986815;
  wire [7:0] sel_986816;
  wire [7:0] add_986819;
  wire [7:0] sel_986820;
  wire [7:0] add_986823;
  wire [7:0] sel_986824;
  wire [7:0] add_986827;
  wire [7:0] sel_986828;
  wire [7:0] add_986831;
  wire [7:0] sel_986832;
  wire [7:0] add_986835;
  wire [7:0] sel_986836;
  wire [7:0] add_986839;
  wire [7:0] sel_986840;
  wire [7:0] add_986843;
  wire [7:0] sel_986844;
  wire [7:0] add_986847;
  wire [7:0] sel_986848;
  wire [7:0] add_986851;
  wire [7:0] sel_986852;
  wire [7:0] add_986855;
  wire [7:0] sel_986856;
  wire [7:0] add_986859;
  wire [7:0] sel_986860;
  wire [7:0] add_986863;
  wire [7:0] sel_986864;
  wire [7:0] add_986867;
  wire [7:0] sel_986868;
  wire [7:0] add_986871;
  wire [7:0] sel_986872;
  wire [7:0] add_986875;
  wire [7:0] sel_986876;
  wire [7:0] add_986880;
  wire [15:0] array_index_986881;
  wire [7:0] sel_986882;
  wire [7:0] add_986885;
  wire [7:0] sel_986886;
  wire [7:0] add_986889;
  wire [7:0] sel_986890;
  wire [7:0] add_986893;
  wire [7:0] sel_986894;
  wire [7:0] add_986897;
  wire [7:0] sel_986898;
  wire [7:0] add_986901;
  wire [7:0] sel_986902;
  wire [7:0] add_986905;
  wire [7:0] sel_986906;
  wire [7:0] add_986909;
  wire [7:0] sel_986910;
  wire [7:0] add_986913;
  wire [7:0] sel_986914;
  wire [7:0] add_986917;
  wire [7:0] sel_986918;
  wire [7:0] add_986921;
  wire [7:0] sel_986922;
  wire [7:0] add_986925;
  wire [7:0] sel_986926;
  wire [7:0] add_986929;
  wire [7:0] sel_986930;
  wire [7:0] add_986933;
  wire [7:0] sel_986934;
  wire [7:0] add_986937;
  wire [7:0] sel_986938;
  wire [7:0] add_986941;
  wire [7:0] sel_986942;
  wire [7:0] add_986945;
  wire [7:0] sel_986946;
  wire [7:0] add_986949;
  wire [7:0] sel_986950;
  wire [7:0] add_986953;
  wire [7:0] sel_986954;
  wire [7:0] add_986957;
  wire [7:0] sel_986958;
  wire [7:0] add_986961;
  wire [7:0] sel_986962;
  wire [7:0] add_986965;
  wire [7:0] sel_986966;
  wire [7:0] add_986969;
  wire [7:0] sel_986970;
  wire [7:0] add_986973;
  wire [7:0] sel_986974;
  wire [7:0] add_986977;
  wire [7:0] sel_986978;
  wire [7:0] add_986981;
  wire [7:0] sel_986982;
  wire [7:0] add_986985;
  wire [7:0] sel_986986;
  wire [7:0] add_986989;
  wire [7:0] sel_986990;
  wire [7:0] add_986993;
  wire [7:0] sel_986994;
  wire [7:0] add_986997;
  wire [7:0] sel_986998;
  wire [7:0] add_987001;
  wire [7:0] sel_987002;
  wire [7:0] add_987005;
  wire [7:0] sel_987006;
  wire [7:0] add_987009;
  wire [7:0] sel_987010;
  wire [7:0] add_987013;
  wire [7:0] sel_987014;
  wire [7:0] add_987017;
  wire [7:0] sel_987018;
  wire [7:0] add_987021;
  wire [7:0] sel_987022;
  wire [7:0] add_987025;
  wire [7:0] sel_987026;
  wire [7:0] add_987029;
  wire [7:0] sel_987030;
  wire [7:0] add_987033;
  wire [7:0] sel_987034;
  wire [7:0] add_987037;
  wire [7:0] sel_987038;
  wire [7:0] add_987041;
  wire [7:0] sel_987042;
  wire [7:0] add_987045;
  wire [7:0] sel_987046;
  wire [7:0] add_987049;
  wire [7:0] sel_987050;
  wire [7:0] add_987053;
  wire [7:0] sel_987054;
  wire [7:0] add_987057;
  wire [7:0] sel_987058;
  wire [7:0] add_987061;
  wire [7:0] sel_987062;
  wire [7:0] add_987065;
  wire [7:0] sel_987066;
  wire [7:0] add_987069;
  wire [7:0] sel_987070;
  wire [7:0] add_987073;
  wire [7:0] sel_987074;
  wire [7:0] add_987077;
  wire [7:0] sel_987078;
  wire [7:0] add_987081;
  wire [7:0] sel_987082;
  wire [7:0] add_987085;
  wire [7:0] sel_987086;
  wire [7:0] add_987089;
  wire [7:0] sel_987090;
  wire [7:0] add_987093;
  wire [7:0] sel_987094;
  wire [7:0] add_987097;
  wire [7:0] sel_987098;
  wire [7:0] add_987101;
  wire [7:0] sel_987102;
  wire [7:0] add_987105;
  wire [7:0] sel_987106;
  wire [7:0] add_987109;
  wire [7:0] sel_987110;
  wire [7:0] add_987113;
  wire [7:0] sel_987114;
  wire [7:0] add_987117;
  wire [7:0] sel_987118;
  wire [7:0] add_987121;
  wire [7:0] sel_987122;
  wire [7:0] add_987125;
  wire [7:0] sel_987126;
  wire [7:0] add_987129;
  wire [7:0] sel_987130;
  wire [7:0] add_987133;
  wire [7:0] sel_987134;
  wire [7:0] add_987137;
  wire [7:0] sel_987138;
  wire [7:0] add_987141;
  wire [7:0] sel_987142;
  wire [7:0] add_987145;
  wire [7:0] sel_987146;
  wire [7:0] add_987149;
  wire [7:0] sel_987150;
  wire [7:0] add_987153;
  wire [7:0] sel_987154;
  wire [7:0] add_987157;
  wire [7:0] sel_987158;
  wire [7:0] add_987161;
  wire [7:0] sel_987162;
  wire [7:0] add_987165;
  wire [7:0] sel_987166;
  wire [7:0] add_987169;
  wire [7:0] sel_987170;
  wire [7:0] add_987173;
  wire [7:0] sel_987174;
  wire [7:0] add_987177;
  wire [7:0] sel_987178;
  wire [7:0] add_987181;
  wire [7:0] sel_987182;
  wire [7:0] add_987185;
  wire [7:0] sel_987186;
  wire [7:0] add_987189;
  wire [7:0] sel_987190;
  wire [7:0] add_987193;
  wire [7:0] sel_987194;
  wire [7:0] add_987197;
  wire [7:0] sel_987198;
  wire [7:0] add_987201;
  wire [7:0] sel_987202;
  wire [7:0] add_987205;
  wire [7:0] sel_987206;
  wire [7:0] add_987209;
  wire [7:0] sel_987210;
  wire [7:0] add_987213;
  wire [7:0] sel_987214;
  wire [7:0] add_987217;
  wire [7:0] sel_987218;
  wire [7:0] add_987221;
  wire [7:0] sel_987222;
  wire [7:0] add_987225;
  wire [7:0] sel_987226;
  wire [7:0] add_987229;
  wire [7:0] sel_987230;
  wire [7:0] add_987233;
  wire [7:0] sel_987234;
  wire [7:0] add_987237;
  wire [7:0] sel_987238;
  wire [7:0] add_987241;
  wire [7:0] sel_987242;
  wire [7:0] add_987245;
  wire [7:0] sel_987246;
  wire [7:0] add_987249;
  wire [7:0] sel_987250;
  wire [7:0] add_987253;
  wire [7:0] sel_987254;
  wire [7:0] add_987257;
  wire [7:0] sel_987258;
  wire [7:0] add_987261;
  wire [7:0] sel_987262;
  wire [7:0] add_987265;
  wire [7:0] sel_987266;
  wire [7:0] add_987269;
  wire [7:0] sel_987270;
  wire [7:0] add_987273;
  wire [7:0] sel_987274;
  wire [7:0] add_987277;
  wire [7:0] sel_987278;
  wire [7:0] add_987282;
  wire [15:0] array_index_987283;
  wire [7:0] sel_987284;
  wire [7:0] add_987287;
  wire [7:0] sel_987288;
  wire [7:0] add_987291;
  wire [7:0] sel_987292;
  wire [7:0] add_987295;
  wire [7:0] sel_987296;
  wire [7:0] add_987299;
  wire [7:0] sel_987300;
  wire [7:0] add_987303;
  wire [7:0] sel_987304;
  wire [7:0] add_987307;
  wire [7:0] sel_987308;
  wire [7:0] add_987311;
  wire [7:0] sel_987312;
  wire [7:0] add_987315;
  wire [7:0] sel_987316;
  wire [7:0] add_987319;
  wire [7:0] sel_987320;
  wire [7:0] add_987323;
  wire [7:0] sel_987324;
  wire [7:0] add_987327;
  wire [7:0] sel_987328;
  wire [7:0] add_987331;
  wire [7:0] sel_987332;
  wire [7:0] add_987335;
  wire [7:0] sel_987336;
  wire [7:0] add_987339;
  wire [7:0] sel_987340;
  wire [7:0] add_987343;
  wire [7:0] sel_987344;
  wire [7:0] add_987347;
  wire [7:0] sel_987348;
  wire [7:0] add_987351;
  wire [7:0] sel_987352;
  wire [7:0] add_987355;
  wire [7:0] sel_987356;
  wire [7:0] add_987359;
  wire [7:0] sel_987360;
  wire [7:0] add_987363;
  wire [7:0] sel_987364;
  wire [7:0] add_987367;
  wire [7:0] sel_987368;
  wire [7:0] add_987371;
  wire [7:0] sel_987372;
  wire [7:0] add_987375;
  wire [7:0] sel_987376;
  wire [7:0] add_987379;
  wire [7:0] sel_987380;
  wire [7:0] add_987383;
  wire [7:0] sel_987384;
  wire [7:0] add_987387;
  wire [7:0] sel_987388;
  wire [7:0] add_987391;
  wire [7:0] sel_987392;
  wire [7:0] add_987395;
  wire [7:0] sel_987396;
  wire [7:0] add_987399;
  wire [7:0] sel_987400;
  wire [7:0] add_987403;
  wire [7:0] sel_987404;
  wire [7:0] add_987407;
  wire [7:0] sel_987408;
  wire [7:0] add_987411;
  wire [7:0] sel_987412;
  wire [7:0] add_987415;
  wire [7:0] sel_987416;
  wire [7:0] add_987419;
  wire [7:0] sel_987420;
  wire [7:0] add_987423;
  wire [7:0] sel_987424;
  wire [7:0] add_987427;
  wire [7:0] sel_987428;
  wire [7:0] add_987431;
  wire [7:0] sel_987432;
  wire [7:0] add_987435;
  wire [7:0] sel_987436;
  wire [7:0] add_987439;
  wire [7:0] sel_987440;
  wire [7:0] add_987443;
  wire [7:0] sel_987444;
  wire [7:0] add_987447;
  wire [7:0] sel_987448;
  wire [7:0] add_987451;
  wire [7:0] sel_987452;
  wire [7:0] add_987455;
  wire [7:0] sel_987456;
  wire [7:0] add_987459;
  wire [7:0] sel_987460;
  wire [7:0] add_987463;
  wire [7:0] sel_987464;
  wire [7:0] add_987467;
  wire [7:0] sel_987468;
  wire [7:0] add_987471;
  wire [7:0] sel_987472;
  wire [7:0] add_987475;
  wire [7:0] sel_987476;
  wire [7:0] add_987479;
  wire [7:0] sel_987480;
  wire [7:0] add_987483;
  wire [7:0] sel_987484;
  wire [7:0] add_987487;
  wire [7:0] sel_987488;
  wire [7:0] add_987491;
  wire [7:0] sel_987492;
  wire [7:0] add_987495;
  wire [7:0] sel_987496;
  wire [7:0] add_987499;
  wire [7:0] sel_987500;
  wire [7:0] add_987503;
  wire [7:0] sel_987504;
  wire [7:0] add_987507;
  wire [7:0] sel_987508;
  wire [7:0] add_987511;
  wire [7:0] sel_987512;
  wire [7:0] add_987515;
  wire [7:0] sel_987516;
  wire [7:0] add_987519;
  wire [7:0] sel_987520;
  wire [7:0] add_987523;
  wire [7:0] sel_987524;
  wire [7:0] add_987527;
  wire [7:0] sel_987528;
  wire [7:0] add_987531;
  wire [7:0] sel_987532;
  wire [7:0] add_987535;
  wire [7:0] sel_987536;
  wire [7:0] add_987539;
  wire [7:0] sel_987540;
  wire [7:0] add_987543;
  wire [7:0] sel_987544;
  wire [7:0] add_987547;
  wire [7:0] sel_987548;
  wire [7:0] add_987551;
  wire [7:0] sel_987552;
  wire [7:0] add_987555;
  wire [7:0] sel_987556;
  wire [7:0] add_987559;
  wire [7:0] sel_987560;
  wire [7:0] add_987563;
  wire [7:0] sel_987564;
  wire [7:0] add_987567;
  wire [7:0] sel_987568;
  wire [7:0] add_987571;
  wire [7:0] sel_987572;
  wire [7:0] add_987575;
  wire [7:0] sel_987576;
  wire [7:0] add_987579;
  wire [7:0] sel_987580;
  wire [7:0] add_987583;
  wire [7:0] sel_987584;
  wire [7:0] add_987587;
  wire [7:0] sel_987588;
  wire [7:0] add_987591;
  wire [7:0] sel_987592;
  wire [7:0] add_987595;
  wire [7:0] sel_987596;
  wire [7:0] add_987599;
  wire [7:0] sel_987600;
  wire [7:0] add_987603;
  wire [7:0] sel_987604;
  wire [7:0] add_987607;
  wire [7:0] sel_987608;
  wire [7:0] add_987611;
  wire [7:0] sel_987612;
  wire [7:0] add_987615;
  wire [7:0] sel_987616;
  wire [7:0] add_987619;
  wire [7:0] sel_987620;
  wire [7:0] add_987623;
  wire [7:0] sel_987624;
  wire [7:0] add_987627;
  wire [7:0] sel_987628;
  wire [7:0] add_987631;
  wire [7:0] sel_987632;
  wire [7:0] add_987635;
  wire [7:0] sel_987636;
  wire [7:0] add_987639;
  wire [7:0] sel_987640;
  wire [7:0] add_987643;
  wire [7:0] sel_987644;
  wire [7:0] add_987647;
  wire [7:0] sel_987648;
  wire [7:0] add_987651;
  wire [7:0] sel_987652;
  wire [7:0] add_987655;
  wire [7:0] sel_987656;
  wire [7:0] add_987659;
  wire [7:0] sel_987660;
  wire [7:0] add_987663;
  wire [7:0] sel_987664;
  wire [7:0] add_987667;
  wire [7:0] sel_987668;
  wire [7:0] add_987671;
  wire [7:0] sel_987672;
  wire [7:0] add_987675;
  wire [7:0] sel_987676;
  wire [7:0] add_987679;
  wire [7:0] sel_987680;
  wire [7:0] add_987684;
  wire [15:0] array_index_987685;
  wire [7:0] sel_987686;
  wire [7:0] add_987689;
  wire [7:0] sel_987690;
  wire [7:0] add_987693;
  wire [7:0] sel_987694;
  wire [7:0] add_987697;
  wire [7:0] sel_987698;
  wire [7:0] add_987701;
  wire [7:0] sel_987702;
  wire [7:0] add_987705;
  wire [7:0] sel_987706;
  wire [7:0] add_987709;
  wire [7:0] sel_987710;
  wire [7:0] add_987713;
  wire [7:0] sel_987714;
  wire [7:0] add_987717;
  wire [7:0] sel_987718;
  wire [7:0] add_987721;
  wire [7:0] sel_987722;
  wire [7:0] add_987725;
  wire [7:0] sel_987726;
  wire [7:0] add_987729;
  wire [7:0] sel_987730;
  wire [7:0] add_987733;
  wire [7:0] sel_987734;
  wire [7:0] add_987737;
  wire [7:0] sel_987738;
  wire [7:0] add_987741;
  wire [7:0] sel_987742;
  wire [7:0] add_987745;
  wire [7:0] sel_987746;
  wire [7:0] add_987749;
  wire [7:0] sel_987750;
  wire [7:0] add_987753;
  wire [7:0] sel_987754;
  wire [7:0] add_987757;
  wire [7:0] sel_987758;
  wire [7:0] add_987761;
  wire [7:0] sel_987762;
  wire [7:0] add_987765;
  wire [7:0] sel_987766;
  wire [7:0] add_987769;
  wire [7:0] sel_987770;
  wire [7:0] add_987773;
  wire [7:0] sel_987774;
  wire [7:0] add_987777;
  wire [7:0] sel_987778;
  wire [7:0] add_987781;
  wire [7:0] sel_987782;
  wire [7:0] add_987785;
  wire [7:0] sel_987786;
  wire [7:0] add_987789;
  wire [7:0] sel_987790;
  wire [7:0] add_987793;
  wire [7:0] sel_987794;
  wire [7:0] add_987797;
  wire [7:0] sel_987798;
  wire [7:0] add_987801;
  wire [7:0] sel_987802;
  wire [7:0] add_987805;
  wire [7:0] sel_987806;
  wire [7:0] add_987809;
  wire [7:0] sel_987810;
  wire [7:0] add_987813;
  wire [7:0] sel_987814;
  wire [7:0] add_987817;
  wire [7:0] sel_987818;
  wire [7:0] add_987821;
  wire [7:0] sel_987822;
  wire [7:0] add_987825;
  wire [7:0] sel_987826;
  wire [7:0] add_987829;
  wire [7:0] sel_987830;
  wire [7:0] add_987833;
  wire [7:0] sel_987834;
  wire [7:0] add_987837;
  wire [7:0] sel_987838;
  wire [7:0] add_987841;
  wire [7:0] sel_987842;
  wire [7:0] add_987845;
  wire [7:0] sel_987846;
  wire [7:0] add_987849;
  wire [7:0] sel_987850;
  wire [7:0] add_987853;
  wire [7:0] sel_987854;
  wire [7:0] add_987857;
  wire [7:0] sel_987858;
  wire [7:0] add_987861;
  wire [7:0] sel_987862;
  wire [7:0] add_987865;
  wire [7:0] sel_987866;
  wire [7:0] add_987869;
  wire [7:0] sel_987870;
  wire [7:0] add_987873;
  wire [7:0] sel_987874;
  wire [7:0] add_987877;
  wire [7:0] sel_987878;
  wire [7:0] add_987881;
  wire [7:0] sel_987882;
  wire [7:0] add_987885;
  wire [7:0] sel_987886;
  wire [7:0] add_987889;
  wire [7:0] sel_987890;
  wire [7:0] add_987893;
  wire [7:0] sel_987894;
  wire [7:0] add_987897;
  wire [7:0] sel_987898;
  wire [7:0] add_987901;
  wire [7:0] sel_987902;
  wire [7:0] add_987905;
  wire [7:0] sel_987906;
  wire [7:0] add_987909;
  wire [7:0] sel_987910;
  wire [7:0] add_987913;
  wire [7:0] sel_987914;
  wire [7:0] add_987917;
  wire [7:0] sel_987918;
  wire [7:0] add_987921;
  wire [7:0] sel_987922;
  wire [7:0] add_987925;
  wire [7:0] sel_987926;
  wire [7:0] add_987929;
  wire [7:0] sel_987930;
  wire [7:0] add_987933;
  wire [7:0] sel_987934;
  wire [7:0] add_987937;
  wire [7:0] sel_987938;
  wire [7:0] add_987941;
  wire [7:0] sel_987942;
  wire [7:0] add_987945;
  wire [7:0] sel_987946;
  wire [7:0] add_987949;
  wire [7:0] sel_987950;
  wire [7:0] add_987953;
  wire [7:0] sel_987954;
  wire [7:0] add_987957;
  wire [7:0] sel_987958;
  wire [7:0] add_987961;
  wire [7:0] sel_987962;
  wire [7:0] add_987965;
  wire [7:0] sel_987966;
  wire [7:0] add_987969;
  wire [7:0] sel_987970;
  wire [7:0] add_987973;
  wire [7:0] sel_987974;
  wire [7:0] add_987977;
  wire [7:0] sel_987978;
  wire [7:0] add_987981;
  wire [7:0] sel_987982;
  wire [7:0] add_987985;
  wire [7:0] sel_987986;
  wire [7:0] add_987989;
  wire [7:0] sel_987990;
  wire [7:0] add_987993;
  wire [7:0] sel_987994;
  wire [7:0] add_987997;
  wire [7:0] sel_987998;
  wire [7:0] add_988001;
  wire [7:0] sel_988002;
  wire [7:0] add_988005;
  wire [7:0] sel_988006;
  wire [7:0] add_988009;
  wire [7:0] sel_988010;
  wire [7:0] add_988013;
  wire [7:0] sel_988014;
  wire [7:0] add_988017;
  wire [7:0] sel_988018;
  wire [7:0] add_988021;
  wire [7:0] sel_988022;
  wire [7:0] add_988025;
  wire [7:0] sel_988026;
  wire [7:0] add_988029;
  wire [7:0] sel_988030;
  wire [7:0] add_988033;
  wire [7:0] sel_988034;
  wire [7:0] add_988037;
  wire [7:0] sel_988038;
  wire [7:0] add_988041;
  wire [7:0] sel_988042;
  wire [7:0] add_988045;
  wire [7:0] sel_988046;
  wire [7:0] add_988049;
  wire [7:0] sel_988050;
  wire [7:0] add_988053;
  wire [7:0] sel_988054;
  wire [7:0] add_988057;
  wire [7:0] sel_988058;
  wire [7:0] add_988061;
  wire [7:0] sel_988062;
  wire [7:0] add_988065;
  wire [7:0] sel_988066;
  wire [7:0] add_988069;
  wire [7:0] sel_988070;
  wire [7:0] add_988073;
  wire [7:0] sel_988074;
  wire [7:0] add_988077;
  wire [7:0] sel_988078;
  wire [7:0] add_988081;
  wire [7:0] sel_988082;
  wire [7:0] add_988086;
  wire [15:0] array_index_988087;
  wire [7:0] sel_988088;
  wire [7:0] add_988091;
  wire [7:0] sel_988092;
  wire [7:0] add_988095;
  wire [7:0] sel_988096;
  wire [7:0] add_988099;
  wire [7:0] sel_988100;
  wire [7:0] add_988103;
  wire [7:0] sel_988104;
  wire [7:0] add_988107;
  wire [7:0] sel_988108;
  wire [7:0] add_988111;
  wire [7:0] sel_988112;
  wire [7:0] add_988115;
  wire [7:0] sel_988116;
  wire [7:0] add_988119;
  wire [7:0] sel_988120;
  wire [7:0] add_988123;
  wire [7:0] sel_988124;
  wire [7:0] add_988127;
  wire [7:0] sel_988128;
  wire [7:0] add_988131;
  wire [7:0] sel_988132;
  wire [7:0] add_988135;
  wire [7:0] sel_988136;
  wire [7:0] add_988139;
  wire [7:0] sel_988140;
  wire [7:0] add_988143;
  wire [7:0] sel_988144;
  wire [7:0] add_988147;
  wire [7:0] sel_988148;
  wire [7:0] add_988151;
  wire [7:0] sel_988152;
  wire [7:0] add_988155;
  wire [7:0] sel_988156;
  wire [7:0] add_988159;
  wire [7:0] sel_988160;
  wire [7:0] add_988163;
  wire [7:0] sel_988164;
  wire [7:0] add_988167;
  wire [7:0] sel_988168;
  wire [7:0] add_988171;
  wire [7:0] sel_988172;
  wire [7:0] add_988175;
  wire [7:0] sel_988176;
  wire [7:0] add_988179;
  wire [7:0] sel_988180;
  wire [7:0] add_988183;
  wire [7:0] sel_988184;
  wire [7:0] add_988187;
  wire [7:0] sel_988188;
  wire [7:0] add_988191;
  wire [7:0] sel_988192;
  wire [7:0] add_988195;
  wire [7:0] sel_988196;
  wire [7:0] add_988199;
  wire [7:0] sel_988200;
  wire [7:0] add_988203;
  wire [7:0] sel_988204;
  wire [7:0] add_988207;
  wire [7:0] sel_988208;
  wire [7:0] add_988211;
  wire [7:0] sel_988212;
  wire [7:0] add_988215;
  wire [7:0] sel_988216;
  wire [7:0] add_988219;
  wire [7:0] sel_988220;
  wire [7:0] add_988223;
  wire [7:0] sel_988224;
  wire [7:0] add_988227;
  wire [7:0] sel_988228;
  wire [7:0] add_988231;
  wire [7:0] sel_988232;
  wire [7:0] add_988235;
  wire [7:0] sel_988236;
  wire [7:0] add_988239;
  wire [7:0] sel_988240;
  wire [7:0] add_988243;
  wire [7:0] sel_988244;
  wire [7:0] add_988247;
  wire [7:0] sel_988248;
  wire [7:0] add_988251;
  wire [7:0] sel_988252;
  wire [7:0] add_988255;
  wire [7:0] sel_988256;
  wire [7:0] add_988259;
  wire [7:0] sel_988260;
  wire [7:0] add_988263;
  wire [7:0] sel_988264;
  wire [7:0] add_988267;
  wire [7:0] sel_988268;
  wire [7:0] add_988271;
  wire [7:0] sel_988272;
  wire [7:0] add_988275;
  wire [7:0] sel_988276;
  wire [7:0] add_988279;
  wire [7:0] sel_988280;
  wire [7:0] add_988283;
  wire [7:0] sel_988284;
  wire [7:0] add_988287;
  wire [7:0] sel_988288;
  wire [7:0] add_988291;
  wire [7:0] sel_988292;
  wire [7:0] add_988295;
  wire [7:0] sel_988296;
  wire [7:0] add_988299;
  wire [7:0] sel_988300;
  wire [7:0] add_988303;
  wire [7:0] sel_988304;
  wire [7:0] add_988307;
  wire [7:0] sel_988308;
  wire [7:0] add_988311;
  wire [7:0] sel_988312;
  wire [7:0] add_988315;
  wire [7:0] sel_988316;
  wire [7:0] add_988319;
  wire [7:0] sel_988320;
  wire [7:0] add_988323;
  wire [7:0] sel_988324;
  wire [7:0] add_988327;
  wire [7:0] sel_988328;
  wire [7:0] add_988331;
  wire [7:0] sel_988332;
  wire [7:0] add_988335;
  wire [7:0] sel_988336;
  wire [7:0] add_988339;
  wire [7:0] sel_988340;
  wire [7:0] add_988343;
  wire [7:0] sel_988344;
  wire [7:0] add_988347;
  wire [7:0] sel_988348;
  wire [7:0] add_988351;
  wire [7:0] sel_988352;
  wire [7:0] add_988355;
  wire [7:0] sel_988356;
  wire [7:0] add_988359;
  wire [7:0] sel_988360;
  wire [7:0] add_988363;
  wire [7:0] sel_988364;
  wire [7:0] add_988367;
  wire [7:0] sel_988368;
  wire [7:0] add_988371;
  wire [7:0] sel_988372;
  wire [7:0] add_988375;
  wire [7:0] sel_988376;
  wire [7:0] add_988379;
  wire [7:0] sel_988380;
  wire [7:0] add_988383;
  wire [7:0] sel_988384;
  wire [7:0] add_988387;
  wire [7:0] sel_988388;
  wire [7:0] add_988391;
  wire [7:0] sel_988392;
  wire [7:0] add_988395;
  wire [7:0] sel_988396;
  wire [7:0] add_988399;
  wire [7:0] sel_988400;
  wire [7:0] add_988403;
  wire [7:0] sel_988404;
  wire [7:0] add_988407;
  wire [7:0] sel_988408;
  wire [7:0] add_988411;
  wire [7:0] sel_988412;
  wire [7:0] add_988415;
  wire [7:0] sel_988416;
  wire [7:0] add_988419;
  wire [7:0] sel_988420;
  wire [7:0] add_988423;
  wire [7:0] sel_988424;
  wire [7:0] add_988427;
  wire [7:0] sel_988428;
  wire [7:0] add_988431;
  wire [7:0] sel_988432;
  wire [7:0] add_988435;
  wire [7:0] sel_988436;
  wire [7:0] add_988439;
  wire [7:0] sel_988440;
  wire [7:0] add_988443;
  wire [7:0] sel_988444;
  wire [7:0] add_988447;
  wire [7:0] sel_988448;
  wire [7:0] add_988451;
  wire [7:0] sel_988452;
  wire [7:0] add_988455;
  wire [7:0] sel_988456;
  wire [7:0] add_988459;
  wire [7:0] sel_988460;
  wire [7:0] add_988463;
  wire [7:0] sel_988464;
  wire [7:0] add_988467;
  wire [7:0] sel_988468;
  wire [7:0] add_988471;
  wire [7:0] sel_988472;
  wire [7:0] add_988475;
  wire [7:0] sel_988476;
  wire [7:0] add_988479;
  wire [7:0] sel_988480;
  wire [7:0] add_988483;
  wire [7:0] sel_988484;
  wire [7:0] add_988488;
  wire [15:0] array_index_988489;
  wire [7:0] sel_988490;
  wire [7:0] add_988493;
  wire [7:0] sel_988494;
  wire [7:0] add_988497;
  wire [7:0] sel_988498;
  wire [7:0] add_988501;
  wire [7:0] sel_988502;
  wire [7:0] add_988505;
  wire [7:0] sel_988506;
  wire [7:0] add_988509;
  wire [7:0] sel_988510;
  wire [7:0] add_988513;
  wire [7:0] sel_988514;
  wire [7:0] add_988517;
  wire [7:0] sel_988518;
  wire [7:0] add_988521;
  wire [7:0] sel_988522;
  wire [7:0] add_988525;
  wire [7:0] sel_988526;
  wire [7:0] add_988529;
  wire [7:0] sel_988530;
  wire [7:0] add_988533;
  wire [7:0] sel_988534;
  wire [7:0] add_988537;
  wire [7:0] sel_988538;
  wire [7:0] add_988541;
  wire [7:0] sel_988542;
  wire [7:0] add_988545;
  wire [7:0] sel_988546;
  wire [7:0] add_988549;
  wire [7:0] sel_988550;
  wire [7:0] add_988553;
  wire [7:0] sel_988554;
  wire [7:0] add_988557;
  wire [7:0] sel_988558;
  wire [7:0] add_988561;
  wire [7:0] sel_988562;
  wire [7:0] add_988565;
  wire [7:0] sel_988566;
  wire [7:0] add_988569;
  wire [7:0] sel_988570;
  wire [7:0] add_988573;
  wire [7:0] sel_988574;
  wire [7:0] add_988577;
  wire [7:0] sel_988578;
  wire [7:0] add_988581;
  wire [7:0] sel_988582;
  wire [7:0] add_988585;
  wire [7:0] sel_988586;
  wire [7:0] add_988589;
  wire [7:0] sel_988590;
  wire [7:0] add_988593;
  wire [7:0] sel_988594;
  wire [7:0] add_988597;
  wire [7:0] sel_988598;
  wire [7:0] add_988601;
  wire [7:0] sel_988602;
  wire [7:0] add_988605;
  wire [7:0] sel_988606;
  wire [7:0] add_988609;
  wire [7:0] sel_988610;
  wire [7:0] add_988613;
  wire [7:0] sel_988614;
  wire [7:0] add_988617;
  wire [7:0] sel_988618;
  wire [7:0] add_988621;
  wire [7:0] sel_988622;
  wire [7:0] add_988625;
  wire [7:0] sel_988626;
  wire [7:0] add_988629;
  wire [7:0] sel_988630;
  wire [7:0] add_988633;
  wire [7:0] sel_988634;
  wire [7:0] add_988637;
  wire [7:0] sel_988638;
  wire [7:0] add_988641;
  wire [7:0] sel_988642;
  wire [7:0] add_988645;
  wire [7:0] sel_988646;
  wire [7:0] add_988649;
  wire [7:0] sel_988650;
  wire [7:0] add_988653;
  wire [7:0] sel_988654;
  wire [7:0] add_988657;
  wire [7:0] sel_988658;
  wire [7:0] add_988661;
  wire [7:0] sel_988662;
  wire [7:0] add_988665;
  wire [7:0] sel_988666;
  wire [7:0] add_988669;
  wire [7:0] sel_988670;
  wire [7:0] add_988673;
  wire [7:0] sel_988674;
  wire [7:0] add_988677;
  wire [7:0] sel_988678;
  wire [7:0] add_988681;
  wire [7:0] sel_988682;
  wire [7:0] add_988685;
  wire [7:0] sel_988686;
  wire [7:0] add_988689;
  wire [7:0] sel_988690;
  wire [7:0] add_988693;
  wire [7:0] sel_988694;
  wire [7:0] add_988697;
  wire [7:0] sel_988698;
  wire [7:0] add_988701;
  wire [7:0] sel_988702;
  wire [7:0] add_988705;
  wire [7:0] sel_988706;
  wire [7:0] add_988709;
  wire [7:0] sel_988710;
  wire [7:0] add_988713;
  wire [7:0] sel_988714;
  wire [7:0] add_988717;
  wire [7:0] sel_988718;
  wire [7:0] add_988721;
  wire [7:0] sel_988722;
  wire [7:0] add_988725;
  wire [7:0] sel_988726;
  wire [7:0] add_988729;
  wire [7:0] sel_988730;
  wire [7:0] add_988733;
  wire [7:0] sel_988734;
  wire [7:0] add_988737;
  wire [7:0] sel_988738;
  wire [7:0] add_988741;
  wire [7:0] sel_988742;
  wire [7:0] add_988745;
  wire [7:0] sel_988746;
  wire [7:0] add_988749;
  wire [7:0] sel_988750;
  wire [7:0] add_988753;
  wire [7:0] sel_988754;
  wire [7:0] add_988757;
  wire [7:0] sel_988758;
  wire [7:0] add_988761;
  wire [7:0] sel_988762;
  wire [7:0] add_988765;
  wire [7:0] sel_988766;
  wire [7:0] add_988769;
  wire [7:0] sel_988770;
  wire [7:0] add_988773;
  wire [7:0] sel_988774;
  wire [7:0] add_988777;
  wire [7:0] sel_988778;
  wire [7:0] add_988781;
  wire [7:0] sel_988782;
  wire [7:0] add_988785;
  wire [7:0] sel_988786;
  wire [7:0] add_988789;
  wire [7:0] sel_988790;
  wire [7:0] add_988793;
  wire [7:0] sel_988794;
  wire [7:0] add_988797;
  wire [7:0] sel_988798;
  wire [7:0] add_988801;
  wire [7:0] sel_988802;
  wire [7:0] add_988805;
  wire [7:0] sel_988806;
  wire [7:0] add_988809;
  wire [7:0] sel_988810;
  wire [7:0] add_988813;
  wire [7:0] sel_988814;
  wire [7:0] add_988817;
  wire [7:0] sel_988818;
  wire [7:0] add_988821;
  wire [7:0] sel_988822;
  wire [7:0] add_988825;
  wire [7:0] sel_988826;
  wire [7:0] add_988829;
  wire [7:0] sel_988830;
  wire [7:0] add_988833;
  wire [7:0] sel_988834;
  wire [7:0] add_988837;
  wire [7:0] sel_988838;
  wire [7:0] add_988841;
  wire [7:0] sel_988842;
  wire [7:0] add_988845;
  wire [7:0] sel_988846;
  wire [7:0] add_988849;
  wire [7:0] sel_988850;
  wire [7:0] add_988853;
  wire [7:0] sel_988854;
  wire [7:0] add_988857;
  wire [7:0] sel_988858;
  wire [7:0] add_988861;
  wire [7:0] sel_988862;
  wire [7:0] add_988865;
  wire [7:0] sel_988866;
  wire [7:0] add_988869;
  wire [7:0] sel_988870;
  wire [7:0] add_988873;
  wire [7:0] sel_988874;
  wire [7:0] add_988877;
  wire [7:0] sel_988878;
  wire [7:0] add_988881;
  wire [7:0] sel_988882;
  wire [7:0] add_988885;
  wire [7:0] sel_988886;
  wire [7:0] add_988889;
  assign array_index_948482 = set1_unflattened[7'h00];
  assign array_index_948483 = set2_unflattened[7'h00];
  assign array_index_948487 = set2_unflattened[7'h01];
  assign concat_948488 = {1'h0, array_index_948482 == array_index_948483};
  assign add_948491 = concat_948488 + 2'h1;
  assign array_index_948495 = set2_unflattened[7'h02];
  assign concat_948496 = {1'h0, array_index_948482 == array_index_948487 ? add_948491 : concat_948488};
  assign add_948499 = concat_948496 + 3'h1;
  assign array_index_948503 = set2_unflattened[7'h03];
  assign concat_948504 = {1'h0, array_index_948482 == array_index_948495 ? add_948499 : concat_948496};
  assign add_948507 = concat_948504 + 4'h1;
  assign array_index_948511 = set2_unflattened[7'h04];
  assign concat_948512 = {1'h0, array_index_948482 == array_index_948503 ? add_948507 : concat_948504};
  assign add_948515 = concat_948512 + 5'h01;
  assign array_index_948519 = set2_unflattened[7'h05];
  assign concat_948520 = {1'h0, array_index_948482 == array_index_948511 ? add_948515 : concat_948512};
  assign add_948523 = concat_948520 + 6'h01;
  assign array_index_948527 = set2_unflattened[7'h06];
  assign concat_948528 = {1'h0, array_index_948482 == array_index_948519 ? add_948523 : concat_948520};
  assign add_948531 = concat_948528 + 7'h01;
  assign array_index_948535 = set2_unflattened[7'h07];
  assign concat_948536 = {1'h0, array_index_948482 == array_index_948527 ? add_948531 : concat_948528};
  assign add_948540 = concat_948536 + 8'h01;
  assign array_index_948541 = set2_unflattened[7'h08];
  assign sel_948542 = array_index_948482 == array_index_948535 ? add_948540 : concat_948536;
  assign add_948546 = sel_948542 + 8'h01;
  assign array_index_948547 = set2_unflattened[7'h09];
  assign sel_948548 = array_index_948482 == array_index_948541 ? add_948546 : sel_948542;
  assign add_948552 = sel_948548 + 8'h01;
  assign array_index_948553 = set2_unflattened[7'h0a];
  assign sel_948554 = array_index_948482 == array_index_948547 ? add_948552 : sel_948548;
  assign add_948558 = sel_948554 + 8'h01;
  assign array_index_948559 = set2_unflattened[7'h0b];
  assign sel_948560 = array_index_948482 == array_index_948553 ? add_948558 : sel_948554;
  assign add_948564 = sel_948560 + 8'h01;
  assign array_index_948565 = set2_unflattened[7'h0c];
  assign sel_948566 = array_index_948482 == array_index_948559 ? add_948564 : sel_948560;
  assign add_948570 = sel_948566 + 8'h01;
  assign array_index_948571 = set2_unflattened[7'h0d];
  assign sel_948572 = array_index_948482 == array_index_948565 ? add_948570 : sel_948566;
  assign add_948576 = sel_948572 + 8'h01;
  assign array_index_948577 = set2_unflattened[7'h0e];
  assign sel_948578 = array_index_948482 == array_index_948571 ? add_948576 : sel_948572;
  assign add_948582 = sel_948578 + 8'h01;
  assign array_index_948583 = set2_unflattened[7'h0f];
  assign sel_948584 = array_index_948482 == array_index_948577 ? add_948582 : sel_948578;
  assign add_948588 = sel_948584 + 8'h01;
  assign array_index_948589 = set2_unflattened[7'h10];
  assign sel_948590 = array_index_948482 == array_index_948583 ? add_948588 : sel_948584;
  assign add_948594 = sel_948590 + 8'h01;
  assign array_index_948595 = set2_unflattened[7'h11];
  assign sel_948596 = array_index_948482 == array_index_948589 ? add_948594 : sel_948590;
  assign add_948600 = sel_948596 + 8'h01;
  assign array_index_948601 = set2_unflattened[7'h12];
  assign sel_948602 = array_index_948482 == array_index_948595 ? add_948600 : sel_948596;
  assign add_948606 = sel_948602 + 8'h01;
  assign array_index_948607 = set2_unflattened[7'h13];
  assign sel_948608 = array_index_948482 == array_index_948601 ? add_948606 : sel_948602;
  assign add_948612 = sel_948608 + 8'h01;
  assign array_index_948613 = set2_unflattened[7'h14];
  assign sel_948614 = array_index_948482 == array_index_948607 ? add_948612 : sel_948608;
  assign add_948618 = sel_948614 + 8'h01;
  assign array_index_948619 = set2_unflattened[7'h15];
  assign sel_948620 = array_index_948482 == array_index_948613 ? add_948618 : sel_948614;
  assign add_948624 = sel_948620 + 8'h01;
  assign array_index_948625 = set2_unflattened[7'h16];
  assign sel_948626 = array_index_948482 == array_index_948619 ? add_948624 : sel_948620;
  assign add_948630 = sel_948626 + 8'h01;
  assign array_index_948631 = set2_unflattened[7'h17];
  assign sel_948632 = array_index_948482 == array_index_948625 ? add_948630 : sel_948626;
  assign add_948636 = sel_948632 + 8'h01;
  assign array_index_948637 = set2_unflattened[7'h18];
  assign sel_948638 = array_index_948482 == array_index_948631 ? add_948636 : sel_948632;
  assign add_948642 = sel_948638 + 8'h01;
  assign array_index_948643 = set2_unflattened[7'h19];
  assign sel_948644 = array_index_948482 == array_index_948637 ? add_948642 : sel_948638;
  assign add_948648 = sel_948644 + 8'h01;
  assign array_index_948649 = set2_unflattened[7'h1a];
  assign sel_948650 = array_index_948482 == array_index_948643 ? add_948648 : sel_948644;
  assign add_948654 = sel_948650 + 8'h01;
  assign array_index_948655 = set2_unflattened[7'h1b];
  assign sel_948656 = array_index_948482 == array_index_948649 ? add_948654 : sel_948650;
  assign add_948660 = sel_948656 + 8'h01;
  assign array_index_948661 = set2_unflattened[7'h1c];
  assign sel_948662 = array_index_948482 == array_index_948655 ? add_948660 : sel_948656;
  assign add_948666 = sel_948662 + 8'h01;
  assign array_index_948667 = set2_unflattened[7'h1d];
  assign sel_948668 = array_index_948482 == array_index_948661 ? add_948666 : sel_948662;
  assign add_948672 = sel_948668 + 8'h01;
  assign array_index_948673 = set2_unflattened[7'h1e];
  assign sel_948674 = array_index_948482 == array_index_948667 ? add_948672 : sel_948668;
  assign add_948678 = sel_948674 + 8'h01;
  assign array_index_948679 = set2_unflattened[7'h1f];
  assign sel_948680 = array_index_948482 == array_index_948673 ? add_948678 : sel_948674;
  assign add_948684 = sel_948680 + 8'h01;
  assign array_index_948685 = set2_unflattened[7'h20];
  assign sel_948686 = array_index_948482 == array_index_948679 ? add_948684 : sel_948680;
  assign add_948690 = sel_948686 + 8'h01;
  assign array_index_948691 = set2_unflattened[7'h21];
  assign sel_948692 = array_index_948482 == array_index_948685 ? add_948690 : sel_948686;
  assign add_948696 = sel_948692 + 8'h01;
  assign array_index_948697 = set2_unflattened[7'h22];
  assign sel_948698 = array_index_948482 == array_index_948691 ? add_948696 : sel_948692;
  assign add_948702 = sel_948698 + 8'h01;
  assign array_index_948703 = set2_unflattened[7'h23];
  assign sel_948704 = array_index_948482 == array_index_948697 ? add_948702 : sel_948698;
  assign add_948708 = sel_948704 + 8'h01;
  assign array_index_948709 = set2_unflattened[7'h24];
  assign sel_948710 = array_index_948482 == array_index_948703 ? add_948708 : sel_948704;
  assign add_948714 = sel_948710 + 8'h01;
  assign array_index_948715 = set2_unflattened[7'h25];
  assign sel_948716 = array_index_948482 == array_index_948709 ? add_948714 : sel_948710;
  assign add_948720 = sel_948716 + 8'h01;
  assign array_index_948721 = set2_unflattened[7'h26];
  assign sel_948722 = array_index_948482 == array_index_948715 ? add_948720 : sel_948716;
  assign add_948726 = sel_948722 + 8'h01;
  assign array_index_948727 = set2_unflattened[7'h27];
  assign sel_948728 = array_index_948482 == array_index_948721 ? add_948726 : sel_948722;
  assign add_948732 = sel_948728 + 8'h01;
  assign array_index_948733 = set2_unflattened[7'h28];
  assign sel_948734 = array_index_948482 == array_index_948727 ? add_948732 : sel_948728;
  assign add_948738 = sel_948734 + 8'h01;
  assign array_index_948739 = set2_unflattened[7'h29];
  assign sel_948740 = array_index_948482 == array_index_948733 ? add_948738 : sel_948734;
  assign add_948744 = sel_948740 + 8'h01;
  assign array_index_948745 = set2_unflattened[7'h2a];
  assign sel_948746 = array_index_948482 == array_index_948739 ? add_948744 : sel_948740;
  assign add_948750 = sel_948746 + 8'h01;
  assign array_index_948751 = set2_unflattened[7'h2b];
  assign sel_948752 = array_index_948482 == array_index_948745 ? add_948750 : sel_948746;
  assign add_948756 = sel_948752 + 8'h01;
  assign array_index_948757 = set2_unflattened[7'h2c];
  assign sel_948758 = array_index_948482 == array_index_948751 ? add_948756 : sel_948752;
  assign add_948762 = sel_948758 + 8'h01;
  assign array_index_948763 = set2_unflattened[7'h2d];
  assign sel_948764 = array_index_948482 == array_index_948757 ? add_948762 : sel_948758;
  assign add_948768 = sel_948764 + 8'h01;
  assign array_index_948769 = set2_unflattened[7'h2e];
  assign sel_948770 = array_index_948482 == array_index_948763 ? add_948768 : sel_948764;
  assign add_948774 = sel_948770 + 8'h01;
  assign array_index_948775 = set2_unflattened[7'h2f];
  assign sel_948776 = array_index_948482 == array_index_948769 ? add_948774 : sel_948770;
  assign add_948780 = sel_948776 + 8'h01;
  assign array_index_948781 = set2_unflattened[7'h30];
  assign sel_948782 = array_index_948482 == array_index_948775 ? add_948780 : sel_948776;
  assign add_948786 = sel_948782 + 8'h01;
  assign array_index_948787 = set2_unflattened[7'h31];
  assign sel_948788 = array_index_948482 == array_index_948781 ? add_948786 : sel_948782;
  assign add_948792 = sel_948788 + 8'h01;
  assign array_index_948793 = set2_unflattened[7'h32];
  assign sel_948794 = array_index_948482 == array_index_948787 ? add_948792 : sel_948788;
  assign add_948798 = sel_948794 + 8'h01;
  assign array_index_948799 = set2_unflattened[7'h33];
  assign sel_948800 = array_index_948482 == array_index_948793 ? add_948798 : sel_948794;
  assign add_948804 = sel_948800 + 8'h01;
  assign array_index_948805 = set2_unflattened[7'h34];
  assign sel_948806 = array_index_948482 == array_index_948799 ? add_948804 : sel_948800;
  assign add_948810 = sel_948806 + 8'h01;
  assign array_index_948811 = set2_unflattened[7'h35];
  assign sel_948812 = array_index_948482 == array_index_948805 ? add_948810 : sel_948806;
  assign add_948816 = sel_948812 + 8'h01;
  assign array_index_948817 = set2_unflattened[7'h36];
  assign sel_948818 = array_index_948482 == array_index_948811 ? add_948816 : sel_948812;
  assign add_948822 = sel_948818 + 8'h01;
  assign array_index_948823 = set2_unflattened[7'h37];
  assign sel_948824 = array_index_948482 == array_index_948817 ? add_948822 : sel_948818;
  assign add_948828 = sel_948824 + 8'h01;
  assign array_index_948829 = set2_unflattened[7'h38];
  assign sel_948830 = array_index_948482 == array_index_948823 ? add_948828 : sel_948824;
  assign add_948834 = sel_948830 + 8'h01;
  assign array_index_948835 = set2_unflattened[7'h39];
  assign sel_948836 = array_index_948482 == array_index_948829 ? add_948834 : sel_948830;
  assign add_948840 = sel_948836 + 8'h01;
  assign array_index_948841 = set2_unflattened[7'h3a];
  assign sel_948842 = array_index_948482 == array_index_948835 ? add_948840 : sel_948836;
  assign add_948846 = sel_948842 + 8'h01;
  assign array_index_948847 = set2_unflattened[7'h3b];
  assign sel_948848 = array_index_948482 == array_index_948841 ? add_948846 : sel_948842;
  assign add_948852 = sel_948848 + 8'h01;
  assign array_index_948853 = set2_unflattened[7'h3c];
  assign sel_948854 = array_index_948482 == array_index_948847 ? add_948852 : sel_948848;
  assign add_948858 = sel_948854 + 8'h01;
  assign array_index_948859 = set2_unflattened[7'h3d];
  assign sel_948860 = array_index_948482 == array_index_948853 ? add_948858 : sel_948854;
  assign add_948864 = sel_948860 + 8'h01;
  assign array_index_948865 = set2_unflattened[7'h3e];
  assign sel_948866 = array_index_948482 == array_index_948859 ? add_948864 : sel_948860;
  assign add_948870 = sel_948866 + 8'h01;
  assign array_index_948871 = set2_unflattened[7'h3f];
  assign sel_948872 = array_index_948482 == array_index_948865 ? add_948870 : sel_948866;
  assign add_948876 = sel_948872 + 8'h01;
  assign array_index_948877 = set2_unflattened[7'h40];
  assign sel_948878 = array_index_948482 == array_index_948871 ? add_948876 : sel_948872;
  assign add_948882 = sel_948878 + 8'h01;
  assign array_index_948883 = set2_unflattened[7'h41];
  assign sel_948884 = array_index_948482 == array_index_948877 ? add_948882 : sel_948878;
  assign add_948888 = sel_948884 + 8'h01;
  assign array_index_948889 = set2_unflattened[7'h42];
  assign sel_948890 = array_index_948482 == array_index_948883 ? add_948888 : sel_948884;
  assign add_948894 = sel_948890 + 8'h01;
  assign array_index_948895 = set2_unflattened[7'h43];
  assign sel_948896 = array_index_948482 == array_index_948889 ? add_948894 : sel_948890;
  assign add_948900 = sel_948896 + 8'h01;
  assign array_index_948901 = set2_unflattened[7'h44];
  assign sel_948902 = array_index_948482 == array_index_948895 ? add_948900 : sel_948896;
  assign add_948906 = sel_948902 + 8'h01;
  assign array_index_948907 = set2_unflattened[7'h45];
  assign sel_948908 = array_index_948482 == array_index_948901 ? add_948906 : sel_948902;
  assign add_948912 = sel_948908 + 8'h01;
  assign array_index_948913 = set2_unflattened[7'h46];
  assign sel_948914 = array_index_948482 == array_index_948907 ? add_948912 : sel_948908;
  assign add_948918 = sel_948914 + 8'h01;
  assign array_index_948919 = set2_unflattened[7'h47];
  assign sel_948920 = array_index_948482 == array_index_948913 ? add_948918 : sel_948914;
  assign add_948924 = sel_948920 + 8'h01;
  assign array_index_948925 = set2_unflattened[7'h48];
  assign sel_948926 = array_index_948482 == array_index_948919 ? add_948924 : sel_948920;
  assign add_948930 = sel_948926 + 8'h01;
  assign array_index_948931 = set2_unflattened[7'h49];
  assign sel_948932 = array_index_948482 == array_index_948925 ? add_948930 : sel_948926;
  assign add_948936 = sel_948932 + 8'h01;
  assign array_index_948937 = set2_unflattened[7'h4a];
  assign sel_948938 = array_index_948482 == array_index_948931 ? add_948936 : sel_948932;
  assign add_948942 = sel_948938 + 8'h01;
  assign array_index_948943 = set2_unflattened[7'h4b];
  assign sel_948944 = array_index_948482 == array_index_948937 ? add_948942 : sel_948938;
  assign add_948948 = sel_948944 + 8'h01;
  assign array_index_948949 = set2_unflattened[7'h4c];
  assign sel_948950 = array_index_948482 == array_index_948943 ? add_948948 : sel_948944;
  assign add_948954 = sel_948950 + 8'h01;
  assign array_index_948955 = set2_unflattened[7'h4d];
  assign sel_948956 = array_index_948482 == array_index_948949 ? add_948954 : sel_948950;
  assign add_948960 = sel_948956 + 8'h01;
  assign array_index_948961 = set2_unflattened[7'h4e];
  assign sel_948962 = array_index_948482 == array_index_948955 ? add_948960 : sel_948956;
  assign add_948966 = sel_948962 + 8'h01;
  assign array_index_948967 = set2_unflattened[7'h4f];
  assign sel_948968 = array_index_948482 == array_index_948961 ? add_948966 : sel_948962;
  assign add_948972 = sel_948968 + 8'h01;
  assign array_index_948973 = set2_unflattened[7'h50];
  assign sel_948974 = array_index_948482 == array_index_948967 ? add_948972 : sel_948968;
  assign add_948978 = sel_948974 + 8'h01;
  assign array_index_948979 = set2_unflattened[7'h51];
  assign sel_948980 = array_index_948482 == array_index_948973 ? add_948978 : sel_948974;
  assign add_948984 = sel_948980 + 8'h01;
  assign array_index_948985 = set2_unflattened[7'h52];
  assign sel_948986 = array_index_948482 == array_index_948979 ? add_948984 : sel_948980;
  assign add_948990 = sel_948986 + 8'h01;
  assign array_index_948991 = set2_unflattened[7'h53];
  assign sel_948992 = array_index_948482 == array_index_948985 ? add_948990 : sel_948986;
  assign add_948996 = sel_948992 + 8'h01;
  assign array_index_948997 = set2_unflattened[7'h54];
  assign sel_948998 = array_index_948482 == array_index_948991 ? add_948996 : sel_948992;
  assign add_949002 = sel_948998 + 8'h01;
  assign array_index_949003 = set2_unflattened[7'h55];
  assign sel_949004 = array_index_948482 == array_index_948997 ? add_949002 : sel_948998;
  assign add_949008 = sel_949004 + 8'h01;
  assign array_index_949009 = set2_unflattened[7'h56];
  assign sel_949010 = array_index_948482 == array_index_949003 ? add_949008 : sel_949004;
  assign add_949014 = sel_949010 + 8'h01;
  assign array_index_949015 = set2_unflattened[7'h57];
  assign sel_949016 = array_index_948482 == array_index_949009 ? add_949014 : sel_949010;
  assign add_949020 = sel_949016 + 8'h01;
  assign array_index_949021 = set2_unflattened[7'h58];
  assign sel_949022 = array_index_948482 == array_index_949015 ? add_949020 : sel_949016;
  assign add_949026 = sel_949022 + 8'h01;
  assign array_index_949027 = set2_unflattened[7'h59];
  assign sel_949028 = array_index_948482 == array_index_949021 ? add_949026 : sel_949022;
  assign add_949032 = sel_949028 + 8'h01;
  assign array_index_949033 = set2_unflattened[7'h5a];
  assign sel_949034 = array_index_948482 == array_index_949027 ? add_949032 : sel_949028;
  assign add_949038 = sel_949034 + 8'h01;
  assign array_index_949039 = set2_unflattened[7'h5b];
  assign sel_949040 = array_index_948482 == array_index_949033 ? add_949038 : sel_949034;
  assign add_949044 = sel_949040 + 8'h01;
  assign array_index_949045 = set2_unflattened[7'h5c];
  assign sel_949046 = array_index_948482 == array_index_949039 ? add_949044 : sel_949040;
  assign add_949050 = sel_949046 + 8'h01;
  assign array_index_949051 = set2_unflattened[7'h5d];
  assign sel_949052 = array_index_948482 == array_index_949045 ? add_949050 : sel_949046;
  assign add_949056 = sel_949052 + 8'h01;
  assign array_index_949057 = set2_unflattened[7'h5e];
  assign sel_949058 = array_index_948482 == array_index_949051 ? add_949056 : sel_949052;
  assign add_949062 = sel_949058 + 8'h01;
  assign array_index_949063 = set2_unflattened[7'h5f];
  assign sel_949064 = array_index_948482 == array_index_949057 ? add_949062 : sel_949058;
  assign add_949068 = sel_949064 + 8'h01;
  assign array_index_949069 = set2_unflattened[7'h60];
  assign sel_949070 = array_index_948482 == array_index_949063 ? add_949068 : sel_949064;
  assign add_949074 = sel_949070 + 8'h01;
  assign array_index_949075 = set2_unflattened[7'h61];
  assign sel_949076 = array_index_948482 == array_index_949069 ? add_949074 : sel_949070;
  assign add_949080 = sel_949076 + 8'h01;
  assign array_index_949081 = set2_unflattened[7'h62];
  assign sel_949082 = array_index_948482 == array_index_949075 ? add_949080 : sel_949076;
  assign add_949086 = sel_949082 + 8'h01;
  assign array_index_949087 = set2_unflattened[7'h63];
  assign sel_949088 = array_index_948482 == array_index_949081 ? add_949086 : sel_949082;
  assign add_949092 = sel_949088 + 8'h01;
  assign array_index_949093 = set1_unflattened[7'h01];
  assign sel_949094 = array_index_948482 == array_index_949087 ? add_949092 : sel_949088;
  assign add_949097 = sel_949094 + 8'h01;
  assign sel_949098 = array_index_949093 == array_index_948483 ? add_949097 : sel_949094;
  assign add_949101 = sel_949098 + 8'h01;
  assign sel_949102 = array_index_949093 == array_index_948487 ? add_949101 : sel_949098;
  assign add_949105 = sel_949102 + 8'h01;
  assign sel_949106 = array_index_949093 == array_index_948495 ? add_949105 : sel_949102;
  assign add_949109 = sel_949106 + 8'h01;
  assign sel_949110 = array_index_949093 == array_index_948503 ? add_949109 : sel_949106;
  assign add_949113 = sel_949110 + 8'h01;
  assign sel_949114 = array_index_949093 == array_index_948511 ? add_949113 : sel_949110;
  assign add_949117 = sel_949114 + 8'h01;
  assign sel_949118 = array_index_949093 == array_index_948519 ? add_949117 : sel_949114;
  assign add_949121 = sel_949118 + 8'h01;
  assign sel_949122 = array_index_949093 == array_index_948527 ? add_949121 : sel_949118;
  assign add_949125 = sel_949122 + 8'h01;
  assign sel_949126 = array_index_949093 == array_index_948535 ? add_949125 : sel_949122;
  assign add_949129 = sel_949126 + 8'h01;
  assign sel_949130 = array_index_949093 == array_index_948541 ? add_949129 : sel_949126;
  assign add_949133 = sel_949130 + 8'h01;
  assign sel_949134 = array_index_949093 == array_index_948547 ? add_949133 : sel_949130;
  assign add_949137 = sel_949134 + 8'h01;
  assign sel_949138 = array_index_949093 == array_index_948553 ? add_949137 : sel_949134;
  assign add_949141 = sel_949138 + 8'h01;
  assign sel_949142 = array_index_949093 == array_index_948559 ? add_949141 : sel_949138;
  assign add_949145 = sel_949142 + 8'h01;
  assign sel_949146 = array_index_949093 == array_index_948565 ? add_949145 : sel_949142;
  assign add_949149 = sel_949146 + 8'h01;
  assign sel_949150 = array_index_949093 == array_index_948571 ? add_949149 : sel_949146;
  assign add_949153 = sel_949150 + 8'h01;
  assign sel_949154 = array_index_949093 == array_index_948577 ? add_949153 : sel_949150;
  assign add_949157 = sel_949154 + 8'h01;
  assign sel_949158 = array_index_949093 == array_index_948583 ? add_949157 : sel_949154;
  assign add_949161 = sel_949158 + 8'h01;
  assign sel_949162 = array_index_949093 == array_index_948589 ? add_949161 : sel_949158;
  assign add_949165 = sel_949162 + 8'h01;
  assign sel_949166 = array_index_949093 == array_index_948595 ? add_949165 : sel_949162;
  assign add_949169 = sel_949166 + 8'h01;
  assign sel_949170 = array_index_949093 == array_index_948601 ? add_949169 : sel_949166;
  assign add_949173 = sel_949170 + 8'h01;
  assign sel_949174 = array_index_949093 == array_index_948607 ? add_949173 : sel_949170;
  assign add_949177 = sel_949174 + 8'h01;
  assign sel_949178 = array_index_949093 == array_index_948613 ? add_949177 : sel_949174;
  assign add_949181 = sel_949178 + 8'h01;
  assign sel_949182 = array_index_949093 == array_index_948619 ? add_949181 : sel_949178;
  assign add_949185 = sel_949182 + 8'h01;
  assign sel_949186 = array_index_949093 == array_index_948625 ? add_949185 : sel_949182;
  assign add_949189 = sel_949186 + 8'h01;
  assign sel_949190 = array_index_949093 == array_index_948631 ? add_949189 : sel_949186;
  assign add_949193 = sel_949190 + 8'h01;
  assign sel_949194 = array_index_949093 == array_index_948637 ? add_949193 : sel_949190;
  assign add_949197 = sel_949194 + 8'h01;
  assign sel_949198 = array_index_949093 == array_index_948643 ? add_949197 : sel_949194;
  assign add_949201 = sel_949198 + 8'h01;
  assign sel_949202 = array_index_949093 == array_index_948649 ? add_949201 : sel_949198;
  assign add_949205 = sel_949202 + 8'h01;
  assign sel_949206 = array_index_949093 == array_index_948655 ? add_949205 : sel_949202;
  assign add_949209 = sel_949206 + 8'h01;
  assign sel_949210 = array_index_949093 == array_index_948661 ? add_949209 : sel_949206;
  assign add_949213 = sel_949210 + 8'h01;
  assign sel_949214 = array_index_949093 == array_index_948667 ? add_949213 : sel_949210;
  assign add_949217 = sel_949214 + 8'h01;
  assign sel_949218 = array_index_949093 == array_index_948673 ? add_949217 : sel_949214;
  assign add_949221 = sel_949218 + 8'h01;
  assign sel_949222 = array_index_949093 == array_index_948679 ? add_949221 : sel_949218;
  assign add_949225 = sel_949222 + 8'h01;
  assign sel_949226 = array_index_949093 == array_index_948685 ? add_949225 : sel_949222;
  assign add_949229 = sel_949226 + 8'h01;
  assign sel_949230 = array_index_949093 == array_index_948691 ? add_949229 : sel_949226;
  assign add_949233 = sel_949230 + 8'h01;
  assign sel_949234 = array_index_949093 == array_index_948697 ? add_949233 : sel_949230;
  assign add_949237 = sel_949234 + 8'h01;
  assign sel_949238 = array_index_949093 == array_index_948703 ? add_949237 : sel_949234;
  assign add_949241 = sel_949238 + 8'h01;
  assign sel_949242 = array_index_949093 == array_index_948709 ? add_949241 : sel_949238;
  assign add_949245 = sel_949242 + 8'h01;
  assign sel_949246 = array_index_949093 == array_index_948715 ? add_949245 : sel_949242;
  assign add_949249 = sel_949246 + 8'h01;
  assign sel_949250 = array_index_949093 == array_index_948721 ? add_949249 : sel_949246;
  assign add_949253 = sel_949250 + 8'h01;
  assign sel_949254 = array_index_949093 == array_index_948727 ? add_949253 : sel_949250;
  assign add_949257 = sel_949254 + 8'h01;
  assign sel_949258 = array_index_949093 == array_index_948733 ? add_949257 : sel_949254;
  assign add_949261 = sel_949258 + 8'h01;
  assign sel_949262 = array_index_949093 == array_index_948739 ? add_949261 : sel_949258;
  assign add_949265 = sel_949262 + 8'h01;
  assign sel_949266 = array_index_949093 == array_index_948745 ? add_949265 : sel_949262;
  assign add_949269 = sel_949266 + 8'h01;
  assign sel_949270 = array_index_949093 == array_index_948751 ? add_949269 : sel_949266;
  assign add_949273 = sel_949270 + 8'h01;
  assign sel_949274 = array_index_949093 == array_index_948757 ? add_949273 : sel_949270;
  assign add_949277 = sel_949274 + 8'h01;
  assign sel_949278 = array_index_949093 == array_index_948763 ? add_949277 : sel_949274;
  assign add_949281 = sel_949278 + 8'h01;
  assign sel_949282 = array_index_949093 == array_index_948769 ? add_949281 : sel_949278;
  assign add_949285 = sel_949282 + 8'h01;
  assign sel_949286 = array_index_949093 == array_index_948775 ? add_949285 : sel_949282;
  assign add_949289 = sel_949286 + 8'h01;
  assign sel_949290 = array_index_949093 == array_index_948781 ? add_949289 : sel_949286;
  assign add_949293 = sel_949290 + 8'h01;
  assign sel_949294 = array_index_949093 == array_index_948787 ? add_949293 : sel_949290;
  assign add_949297 = sel_949294 + 8'h01;
  assign sel_949298 = array_index_949093 == array_index_948793 ? add_949297 : sel_949294;
  assign add_949301 = sel_949298 + 8'h01;
  assign sel_949302 = array_index_949093 == array_index_948799 ? add_949301 : sel_949298;
  assign add_949305 = sel_949302 + 8'h01;
  assign sel_949306 = array_index_949093 == array_index_948805 ? add_949305 : sel_949302;
  assign add_949309 = sel_949306 + 8'h01;
  assign sel_949310 = array_index_949093 == array_index_948811 ? add_949309 : sel_949306;
  assign add_949313 = sel_949310 + 8'h01;
  assign sel_949314 = array_index_949093 == array_index_948817 ? add_949313 : sel_949310;
  assign add_949317 = sel_949314 + 8'h01;
  assign sel_949318 = array_index_949093 == array_index_948823 ? add_949317 : sel_949314;
  assign add_949321 = sel_949318 + 8'h01;
  assign sel_949322 = array_index_949093 == array_index_948829 ? add_949321 : sel_949318;
  assign add_949325 = sel_949322 + 8'h01;
  assign sel_949326 = array_index_949093 == array_index_948835 ? add_949325 : sel_949322;
  assign add_949329 = sel_949326 + 8'h01;
  assign sel_949330 = array_index_949093 == array_index_948841 ? add_949329 : sel_949326;
  assign add_949333 = sel_949330 + 8'h01;
  assign sel_949334 = array_index_949093 == array_index_948847 ? add_949333 : sel_949330;
  assign add_949337 = sel_949334 + 8'h01;
  assign sel_949338 = array_index_949093 == array_index_948853 ? add_949337 : sel_949334;
  assign add_949341 = sel_949338 + 8'h01;
  assign sel_949342 = array_index_949093 == array_index_948859 ? add_949341 : sel_949338;
  assign add_949345 = sel_949342 + 8'h01;
  assign sel_949346 = array_index_949093 == array_index_948865 ? add_949345 : sel_949342;
  assign add_949349 = sel_949346 + 8'h01;
  assign sel_949350 = array_index_949093 == array_index_948871 ? add_949349 : sel_949346;
  assign add_949353 = sel_949350 + 8'h01;
  assign sel_949354 = array_index_949093 == array_index_948877 ? add_949353 : sel_949350;
  assign add_949357 = sel_949354 + 8'h01;
  assign sel_949358 = array_index_949093 == array_index_948883 ? add_949357 : sel_949354;
  assign add_949361 = sel_949358 + 8'h01;
  assign sel_949362 = array_index_949093 == array_index_948889 ? add_949361 : sel_949358;
  assign add_949365 = sel_949362 + 8'h01;
  assign sel_949366 = array_index_949093 == array_index_948895 ? add_949365 : sel_949362;
  assign add_949369 = sel_949366 + 8'h01;
  assign sel_949370 = array_index_949093 == array_index_948901 ? add_949369 : sel_949366;
  assign add_949373 = sel_949370 + 8'h01;
  assign sel_949374 = array_index_949093 == array_index_948907 ? add_949373 : sel_949370;
  assign add_949377 = sel_949374 + 8'h01;
  assign sel_949378 = array_index_949093 == array_index_948913 ? add_949377 : sel_949374;
  assign add_949381 = sel_949378 + 8'h01;
  assign sel_949382 = array_index_949093 == array_index_948919 ? add_949381 : sel_949378;
  assign add_949385 = sel_949382 + 8'h01;
  assign sel_949386 = array_index_949093 == array_index_948925 ? add_949385 : sel_949382;
  assign add_949389 = sel_949386 + 8'h01;
  assign sel_949390 = array_index_949093 == array_index_948931 ? add_949389 : sel_949386;
  assign add_949393 = sel_949390 + 8'h01;
  assign sel_949394 = array_index_949093 == array_index_948937 ? add_949393 : sel_949390;
  assign add_949397 = sel_949394 + 8'h01;
  assign sel_949398 = array_index_949093 == array_index_948943 ? add_949397 : sel_949394;
  assign add_949401 = sel_949398 + 8'h01;
  assign sel_949402 = array_index_949093 == array_index_948949 ? add_949401 : sel_949398;
  assign add_949405 = sel_949402 + 8'h01;
  assign sel_949406 = array_index_949093 == array_index_948955 ? add_949405 : sel_949402;
  assign add_949409 = sel_949406 + 8'h01;
  assign sel_949410 = array_index_949093 == array_index_948961 ? add_949409 : sel_949406;
  assign add_949413 = sel_949410 + 8'h01;
  assign sel_949414 = array_index_949093 == array_index_948967 ? add_949413 : sel_949410;
  assign add_949417 = sel_949414 + 8'h01;
  assign sel_949418 = array_index_949093 == array_index_948973 ? add_949417 : sel_949414;
  assign add_949421 = sel_949418 + 8'h01;
  assign sel_949422 = array_index_949093 == array_index_948979 ? add_949421 : sel_949418;
  assign add_949425 = sel_949422 + 8'h01;
  assign sel_949426 = array_index_949093 == array_index_948985 ? add_949425 : sel_949422;
  assign add_949429 = sel_949426 + 8'h01;
  assign sel_949430 = array_index_949093 == array_index_948991 ? add_949429 : sel_949426;
  assign add_949433 = sel_949430 + 8'h01;
  assign sel_949434 = array_index_949093 == array_index_948997 ? add_949433 : sel_949430;
  assign add_949437 = sel_949434 + 8'h01;
  assign sel_949438 = array_index_949093 == array_index_949003 ? add_949437 : sel_949434;
  assign add_949441 = sel_949438 + 8'h01;
  assign sel_949442 = array_index_949093 == array_index_949009 ? add_949441 : sel_949438;
  assign add_949445 = sel_949442 + 8'h01;
  assign sel_949446 = array_index_949093 == array_index_949015 ? add_949445 : sel_949442;
  assign add_949449 = sel_949446 + 8'h01;
  assign sel_949450 = array_index_949093 == array_index_949021 ? add_949449 : sel_949446;
  assign add_949453 = sel_949450 + 8'h01;
  assign sel_949454 = array_index_949093 == array_index_949027 ? add_949453 : sel_949450;
  assign add_949457 = sel_949454 + 8'h01;
  assign sel_949458 = array_index_949093 == array_index_949033 ? add_949457 : sel_949454;
  assign add_949461 = sel_949458 + 8'h01;
  assign sel_949462 = array_index_949093 == array_index_949039 ? add_949461 : sel_949458;
  assign add_949465 = sel_949462 + 8'h01;
  assign sel_949466 = array_index_949093 == array_index_949045 ? add_949465 : sel_949462;
  assign add_949469 = sel_949466 + 8'h01;
  assign sel_949470 = array_index_949093 == array_index_949051 ? add_949469 : sel_949466;
  assign add_949473 = sel_949470 + 8'h01;
  assign sel_949474 = array_index_949093 == array_index_949057 ? add_949473 : sel_949470;
  assign add_949477 = sel_949474 + 8'h01;
  assign sel_949478 = array_index_949093 == array_index_949063 ? add_949477 : sel_949474;
  assign add_949481 = sel_949478 + 8'h01;
  assign sel_949482 = array_index_949093 == array_index_949069 ? add_949481 : sel_949478;
  assign add_949485 = sel_949482 + 8'h01;
  assign sel_949486 = array_index_949093 == array_index_949075 ? add_949485 : sel_949482;
  assign add_949489 = sel_949486 + 8'h01;
  assign sel_949490 = array_index_949093 == array_index_949081 ? add_949489 : sel_949486;
  assign add_949494 = sel_949490 + 8'h01;
  assign array_index_949495 = set1_unflattened[7'h02];
  assign sel_949496 = array_index_949093 == array_index_949087 ? add_949494 : sel_949490;
  assign add_949499 = sel_949496 + 8'h01;
  assign sel_949500 = array_index_949495 == array_index_948483 ? add_949499 : sel_949496;
  assign add_949503 = sel_949500 + 8'h01;
  assign sel_949504 = array_index_949495 == array_index_948487 ? add_949503 : sel_949500;
  assign add_949507 = sel_949504 + 8'h01;
  assign sel_949508 = array_index_949495 == array_index_948495 ? add_949507 : sel_949504;
  assign add_949511 = sel_949508 + 8'h01;
  assign sel_949512 = array_index_949495 == array_index_948503 ? add_949511 : sel_949508;
  assign add_949515 = sel_949512 + 8'h01;
  assign sel_949516 = array_index_949495 == array_index_948511 ? add_949515 : sel_949512;
  assign add_949519 = sel_949516 + 8'h01;
  assign sel_949520 = array_index_949495 == array_index_948519 ? add_949519 : sel_949516;
  assign add_949523 = sel_949520 + 8'h01;
  assign sel_949524 = array_index_949495 == array_index_948527 ? add_949523 : sel_949520;
  assign add_949527 = sel_949524 + 8'h01;
  assign sel_949528 = array_index_949495 == array_index_948535 ? add_949527 : sel_949524;
  assign add_949531 = sel_949528 + 8'h01;
  assign sel_949532 = array_index_949495 == array_index_948541 ? add_949531 : sel_949528;
  assign add_949535 = sel_949532 + 8'h01;
  assign sel_949536 = array_index_949495 == array_index_948547 ? add_949535 : sel_949532;
  assign add_949539 = sel_949536 + 8'h01;
  assign sel_949540 = array_index_949495 == array_index_948553 ? add_949539 : sel_949536;
  assign add_949543 = sel_949540 + 8'h01;
  assign sel_949544 = array_index_949495 == array_index_948559 ? add_949543 : sel_949540;
  assign add_949547 = sel_949544 + 8'h01;
  assign sel_949548 = array_index_949495 == array_index_948565 ? add_949547 : sel_949544;
  assign add_949551 = sel_949548 + 8'h01;
  assign sel_949552 = array_index_949495 == array_index_948571 ? add_949551 : sel_949548;
  assign add_949555 = sel_949552 + 8'h01;
  assign sel_949556 = array_index_949495 == array_index_948577 ? add_949555 : sel_949552;
  assign add_949559 = sel_949556 + 8'h01;
  assign sel_949560 = array_index_949495 == array_index_948583 ? add_949559 : sel_949556;
  assign add_949563 = sel_949560 + 8'h01;
  assign sel_949564 = array_index_949495 == array_index_948589 ? add_949563 : sel_949560;
  assign add_949567 = sel_949564 + 8'h01;
  assign sel_949568 = array_index_949495 == array_index_948595 ? add_949567 : sel_949564;
  assign add_949571 = sel_949568 + 8'h01;
  assign sel_949572 = array_index_949495 == array_index_948601 ? add_949571 : sel_949568;
  assign add_949575 = sel_949572 + 8'h01;
  assign sel_949576 = array_index_949495 == array_index_948607 ? add_949575 : sel_949572;
  assign add_949579 = sel_949576 + 8'h01;
  assign sel_949580 = array_index_949495 == array_index_948613 ? add_949579 : sel_949576;
  assign add_949583 = sel_949580 + 8'h01;
  assign sel_949584 = array_index_949495 == array_index_948619 ? add_949583 : sel_949580;
  assign add_949587 = sel_949584 + 8'h01;
  assign sel_949588 = array_index_949495 == array_index_948625 ? add_949587 : sel_949584;
  assign add_949591 = sel_949588 + 8'h01;
  assign sel_949592 = array_index_949495 == array_index_948631 ? add_949591 : sel_949588;
  assign add_949595 = sel_949592 + 8'h01;
  assign sel_949596 = array_index_949495 == array_index_948637 ? add_949595 : sel_949592;
  assign add_949599 = sel_949596 + 8'h01;
  assign sel_949600 = array_index_949495 == array_index_948643 ? add_949599 : sel_949596;
  assign add_949603 = sel_949600 + 8'h01;
  assign sel_949604 = array_index_949495 == array_index_948649 ? add_949603 : sel_949600;
  assign add_949607 = sel_949604 + 8'h01;
  assign sel_949608 = array_index_949495 == array_index_948655 ? add_949607 : sel_949604;
  assign add_949611 = sel_949608 + 8'h01;
  assign sel_949612 = array_index_949495 == array_index_948661 ? add_949611 : sel_949608;
  assign add_949615 = sel_949612 + 8'h01;
  assign sel_949616 = array_index_949495 == array_index_948667 ? add_949615 : sel_949612;
  assign add_949619 = sel_949616 + 8'h01;
  assign sel_949620 = array_index_949495 == array_index_948673 ? add_949619 : sel_949616;
  assign add_949623 = sel_949620 + 8'h01;
  assign sel_949624 = array_index_949495 == array_index_948679 ? add_949623 : sel_949620;
  assign add_949627 = sel_949624 + 8'h01;
  assign sel_949628 = array_index_949495 == array_index_948685 ? add_949627 : sel_949624;
  assign add_949631 = sel_949628 + 8'h01;
  assign sel_949632 = array_index_949495 == array_index_948691 ? add_949631 : sel_949628;
  assign add_949635 = sel_949632 + 8'h01;
  assign sel_949636 = array_index_949495 == array_index_948697 ? add_949635 : sel_949632;
  assign add_949639 = sel_949636 + 8'h01;
  assign sel_949640 = array_index_949495 == array_index_948703 ? add_949639 : sel_949636;
  assign add_949643 = sel_949640 + 8'h01;
  assign sel_949644 = array_index_949495 == array_index_948709 ? add_949643 : sel_949640;
  assign add_949647 = sel_949644 + 8'h01;
  assign sel_949648 = array_index_949495 == array_index_948715 ? add_949647 : sel_949644;
  assign add_949651 = sel_949648 + 8'h01;
  assign sel_949652 = array_index_949495 == array_index_948721 ? add_949651 : sel_949648;
  assign add_949655 = sel_949652 + 8'h01;
  assign sel_949656 = array_index_949495 == array_index_948727 ? add_949655 : sel_949652;
  assign add_949659 = sel_949656 + 8'h01;
  assign sel_949660 = array_index_949495 == array_index_948733 ? add_949659 : sel_949656;
  assign add_949663 = sel_949660 + 8'h01;
  assign sel_949664 = array_index_949495 == array_index_948739 ? add_949663 : sel_949660;
  assign add_949667 = sel_949664 + 8'h01;
  assign sel_949668 = array_index_949495 == array_index_948745 ? add_949667 : sel_949664;
  assign add_949671 = sel_949668 + 8'h01;
  assign sel_949672 = array_index_949495 == array_index_948751 ? add_949671 : sel_949668;
  assign add_949675 = sel_949672 + 8'h01;
  assign sel_949676 = array_index_949495 == array_index_948757 ? add_949675 : sel_949672;
  assign add_949679 = sel_949676 + 8'h01;
  assign sel_949680 = array_index_949495 == array_index_948763 ? add_949679 : sel_949676;
  assign add_949683 = sel_949680 + 8'h01;
  assign sel_949684 = array_index_949495 == array_index_948769 ? add_949683 : sel_949680;
  assign add_949687 = sel_949684 + 8'h01;
  assign sel_949688 = array_index_949495 == array_index_948775 ? add_949687 : sel_949684;
  assign add_949691 = sel_949688 + 8'h01;
  assign sel_949692 = array_index_949495 == array_index_948781 ? add_949691 : sel_949688;
  assign add_949695 = sel_949692 + 8'h01;
  assign sel_949696 = array_index_949495 == array_index_948787 ? add_949695 : sel_949692;
  assign add_949699 = sel_949696 + 8'h01;
  assign sel_949700 = array_index_949495 == array_index_948793 ? add_949699 : sel_949696;
  assign add_949703 = sel_949700 + 8'h01;
  assign sel_949704 = array_index_949495 == array_index_948799 ? add_949703 : sel_949700;
  assign add_949707 = sel_949704 + 8'h01;
  assign sel_949708 = array_index_949495 == array_index_948805 ? add_949707 : sel_949704;
  assign add_949711 = sel_949708 + 8'h01;
  assign sel_949712 = array_index_949495 == array_index_948811 ? add_949711 : sel_949708;
  assign add_949715 = sel_949712 + 8'h01;
  assign sel_949716 = array_index_949495 == array_index_948817 ? add_949715 : sel_949712;
  assign add_949719 = sel_949716 + 8'h01;
  assign sel_949720 = array_index_949495 == array_index_948823 ? add_949719 : sel_949716;
  assign add_949723 = sel_949720 + 8'h01;
  assign sel_949724 = array_index_949495 == array_index_948829 ? add_949723 : sel_949720;
  assign add_949727 = sel_949724 + 8'h01;
  assign sel_949728 = array_index_949495 == array_index_948835 ? add_949727 : sel_949724;
  assign add_949731 = sel_949728 + 8'h01;
  assign sel_949732 = array_index_949495 == array_index_948841 ? add_949731 : sel_949728;
  assign add_949735 = sel_949732 + 8'h01;
  assign sel_949736 = array_index_949495 == array_index_948847 ? add_949735 : sel_949732;
  assign add_949739 = sel_949736 + 8'h01;
  assign sel_949740 = array_index_949495 == array_index_948853 ? add_949739 : sel_949736;
  assign add_949743 = sel_949740 + 8'h01;
  assign sel_949744 = array_index_949495 == array_index_948859 ? add_949743 : sel_949740;
  assign add_949747 = sel_949744 + 8'h01;
  assign sel_949748 = array_index_949495 == array_index_948865 ? add_949747 : sel_949744;
  assign add_949751 = sel_949748 + 8'h01;
  assign sel_949752 = array_index_949495 == array_index_948871 ? add_949751 : sel_949748;
  assign add_949755 = sel_949752 + 8'h01;
  assign sel_949756 = array_index_949495 == array_index_948877 ? add_949755 : sel_949752;
  assign add_949759 = sel_949756 + 8'h01;
  assign sel_949760 = array_index_949495 == array_index_948883 ? add_949759 : sel_949756;
  assign add_949763 = sel_949760 + 8'h01;
  assign sel_949764 = array_index_949495 == array_index_948889 ? add_949763 : sel_949760;
  assign add_949767 = sel_949764 + 8'h01;
  assign sel_949768 = array_index_949495 == array_index_948895 ? add_949767 : sel_949764;
  assign add_949771 = sel_949768 + 8'h01;
  assign sel_949772 = array_index_949495 == array_index_948901 ? add_949771 : sel_949768;
  assign add_949775 = sel_949772 + 8'h01;
  assign sel_949776 = array_index_949495 == array_index_948907 ? add_949775 : sel_949772;
  assign add_949779 = sel_949776 + 8'h01;
  assign sel_949780 = array_index_949495 == array_index_948913 ? add_949779 : sel_949776;
  assign add_949783 = sel_949780 + 8'h01;
  assign sel_949784 = array_index_949495 == array_index_948919 ? add_949783 : sel_949780;
  assign add_949787 = sel_949784 + 8'h01;
  assign sel_949788 = array_index_949495 == array_index_948925 ? add_949787 : sel_949784;
  assign add_949791 = sel_949788 + 8'h01;
  assign sel_949792 = array_index_949495 == array_index_948931 ? add_949791 : sel_949788;
  assign add_949795 = sel_949792 + 8'h01;
  assign sel_949796 = array_index_949495 == array_index_948937 ? add_949795 : sel_949792;
  assign add_949799 = sel_949796 + 8'h01;
  assign sel_949800 = array_index_949495 == array_index_948943 ? add_949799 : sel_949796;
  assign add_949803 = sel_949800 + 8'h01;
  assign sel_949804 = array_index_949495 == array_index_948949 ? add_949803 : sel_949800;
  assign add_949807 = sel_949804 + 8'h01;
  assign sel_949808 = array_index_949495 == array_index_948955 ? add_949807 : sel_949804;
  assign add_949811 = sel_949808 + 8'h01;
  assign sel_949812 = array_index_949495 == array_index_948961 ? add_949811 : sel_949808;
  assign add_949815 = sel_949812 + 8'h01;
  assign sel_949816 = array_index_949495 == array_index_948967 ? add_949815 : sel_949812;
  assign add_949819 = sel_949816 + 8'h01;
  assign sel_949820 = array_index_949495 == array_index_948973 ? add_949819 : sel_949816;
  assign add_949823 = sel_949820 + 8'h01;
  assign sel_949824 = array_index_949495 == array_index_948979 ? add_949823 : sel_949820;
  assign add_949827 = sel_949824 + 8'h01;
  assign sel_949828 = array_index_949495 == array_index_948985 ? add_949827 : sel_949824;
  assign add_949831 = sel_949828 + 8'h01;
  assign sel_949832 = array_index_949495 == array_index_948991 ? add_949831 : sel_949828;
  assign add_949835 = sel_949832 + 8'h01;
  assign sel_949836 = array_index_949495 == array_index_948997 ? add_949835 : sel_949832;
  assign add_949839 = sel_949836 + 8'h01;
  assign sel_949840 = array_index_949495 == array_index_949003 ? add_949839 : sel_949836;
  assign add_949843 = sel_949840 + 8'h01;
  assign sel_949844 = array_index_949495 == array_index_949009 ? add_949843 : sel_949840;
  assign add_949847 = sel_949844 + 8'h01;
  assign sel_949848 = array_index_949495 == array_index_949015 ? add_949847 : sel_949844;
  assign add_949851 = sel_949848 + 8'h01;
  assign sel_949852 = array_index_949495 == array_index_949021 ? add_949851 : sel_949848;
  assign add_949855 = sel_949852 + 8'h01;
  assign sel_949856 = array_index_949495 == array_index_949027 ? add_949855 : sel_949852;
  assign add_949859 = sel_949856 + 8'h01;
  assign sel_949860 = array_index_949495 == array_index_949033 ? add_949859 : sel_949856;
  assign add_949863 = sel_949860 + 8'h01;
  assign sel_949864 = array_index_949495 == array_index_949039 ? add_949863 : sel_949860;
  assign add_949867 = sel_949864 + 8'h01;
  assign sel_949868 = array_index_949495 == array_index_949045 ? add_949867 : sel_949864;
  assign add_949871 = sel_949868 + 8'h01;
  assign sel_949872 = array_index_949495 == array_index_949051 ? add_949871 : sel_949868;
  assign add_949875 = sel_949872 + 8'h01;
  assign sel_949876 = array_index_949495 == array_index_949057 ? add_949875 : sel_949872;
  assign add_949879 = sel_949876 + 8'h01;
  assign sel_949880 = array_index_949495 == array_index_949063 ? add_949879 : sel_949876;
  assign add_949883 = sel_949880 + 8'h01;
  assign sel_949884 = array_index_949495 == array_index_949069 ? add_949883 : sel_949880;
  assign add_949887 = sel_949884 + 8'h01;
  assign sel_949888 = array_index_949495 == array_index_949075 ? add_949887 : sel_949884;
  assign add_949891 = sel_949888 + 8'h01;
  assign sel_949892 = array_index_949495 == array_index_949081 ? add_949891 : sel_949888;
  assign add_949896 = sel_949892 + 8'h01;
  assign array_index_949897 = set1_unflattened[7'h03];
  assign sel_949898 = array_index_949495 == array_index_949087 ? add_949896 : sel_949892;
  assign add_949901 = sel_949898 + 8'h01;
  assign sel_949902 = array_index_949897 == array_index_948483 ? add_949901 : sel_949898;
  assign add_949905 = sel_949902 + 8'h01;
  assign sel_949906 = array_index_949897 == array_index_948487 ? add_949905 : sel_949902;
  assign add_949909 = sel_949906 + 8'h01;
  assign sel_949910 = array_index_949897 == array_index_948495 ? add_949909 : sel_949906;
  assign add_949913 = sel_949910 + 8'h01;
  assign sel_949914 = array_index_949897 == array_index_948503 ? add_949913 : sel_949910;
  assign add_949917 = sel_949914 + 8'h01;
  assign sel_949918 = array_index_949897 == array_index_948511 ? add_949917 : sel_949914;
  assign add_949921 = sel_949918 + 8'h01;
  assign sel_949922 = array_index_949897 == array_index_948519 ? add_949921 : sel_949918;
  assign add_949925 = sel_949922 + 8'h01;
  assign sel_949926 = array_index_949897 == array_index_948527 ? add_949925 : sel_949922;
  assign add_949929 = sel_949926 + 8'h01;
  assign sel_949930 = array_index_949897 == array_index_948535 ? add_949929 : sel_949926;
  assign add_949933 = sel_949930 + 8'h01;
  assign sel_949934 = array_index_949897 == array_index_948541 ? add_949933 : sel_949930;
  assign add_949937 = sel_949934 + 8'h01;
  assign sel_949938 = array_index_949897 == array_index_948547 ? add_949937 : sel_949934;
  assign add_949941 = sel_949938 + 8'h01;
  assign sel_949942 = array_index_949897 == array_index_948553 ? add_949941 : sel_949938;
  assign add_949945 = sel_949942 + 8'h01;
  assign sel_949946 = array_index_949897 == array_index_948559 ? add_949945 : sel_949942;
  assign add_949949 = sel_949946 + 8'h01;
  assign sel_949950 = array_index_949897 == array_index_948565 ? add_949949 : sel_949946;
  assign add_949953 = sel_949950 + 8'h01;
  assign sel_949954 = array_index_949897 == array_index_948571 ? add_949953 : sel_949950;
  assign add_949957 = sel_949954 + 8'h01;
  assign sel_949958 = array_index_949897 == array_index_948577 ? add_949957 : sel_949954;
  assign add_949961 = sel_949958 + 8'h01;
  assign sel_949962 = array_index_949897 == array_index_948583 ? add_949961 : sel_949958;
  assign add_949965 = sel_949962 + 8'h01;
  assign sel_949966 = array_index_949897 == array_index_948589 ? add_949965 : sel_949962;
  assign add_949969 = sel_949966 + 8'h01;
  assign sel_949970 = array_index_949897 == array_index_948595 ? add_949969 : sel_949966;
  assign add_949973 = sel_949970 + 8'h01;
  assign sel_949974 = array_index_949897 == array_index_948601 ? add_949973 : sel_949970;
  assign add_949977 = sel_949974 + 8'h01;
  assign sel_949978 = array_index_949897 == array_index_948607 ? add_949977 : sel_949974;
  assign add_949981 = sel_949978 + 8'h01;
  assign sel_949982 = array_index_949897 == array_index_948613 ? add_949981 : sel_949978;
  assign add_949985 = sel_949982 + 8'h01;
  assign sel_949986 = array_index_949897 == array_index_948619 ? add_949985 : sel_949982;
  assign add_949989 = sel_949986 + 8'h01;
  assign sel_949990 = array_index_949897 == array_index_948625 ? add_949989 : sel_949986;
  assign add_949993 = sel_949990 + 8'h01;
  assign sel_949994 = array_index_949897 == array_index_948631 ? add_949993 : sel_949990;
  assign add_949997 = sel_949994 + 8'h01;
  assign sel_949998 = array_index_949897 == array_index_948637 ? add_949997 : sel_949994;
  assign add_950001 = sel_949998 + 8'h01;
  assign sel_950002 = array_index_949897 == array_index_948643 ? add_950001 : sel_949998;
  assign add_950005 = sel_950002 + 8'h01;
  assign sel_950006 = array_index_949897 == array_index_948649 ? add_950005 : sel_950002;
  assign add_950009 = sel_950006 + 8'h01;
  assign sel_950010 = array_index_949897 == array_index_948655 ? add_950009 : sel_950006;
  assign add_950013 = sel_950010 + 8'h01;
  assign sel_950014 = array_index_949897 == array_index_948661 ? add_950013 : sel_950010;
  assign add_950017 = sel_950014 + 8'h01;
  assign sel_950018 = array_index_949897 == array_index_948667 ? add_950017 : sel_950014;
  assign add_950021 = sel_950018 + 8'h01;
  assign sel_950022 = array_index_949897 == array_index_948673 ? add_950021 : sel_950018;
  assign add_950025 = sel_950022 + 8'h01;
  assign sel_950026 = array_index_949897 == array_index_948679 ? add_950025 : sel_950022;
  assign add_950029 = sel_950026 + 8'h01;
  assign sel_950030 = array_index_949897 == array_index_948685 ? add_950029 : sel_950026;
  assign add_950033 = sel_950030 + 8'h01;
  assign sel_950034 = array_index_949897 == array_index_948691 ? add_950033 : sel_950030;
  assign add_950037 = sel_950034 + 8'h01;
  assign sel_950038 = array_index_949897 == array_index_948697 ? add_950037 : sel_950034;
  assign add_950041 = sel_950038 + 8'h01;
  assign sel_950042 = array_index_949897 == array_index_948703 ? add_950041 : sel_950038;
  assign add_950045 = sel_950042 + 8'h01;
  assign sel_950046 = array_index_949897 == array_index_948709 ? add_950045 : sel_950042;
  assign add_950049 = sel_950046 + 8'h01;
  assign sel_950050 = array_index_949897 == array_index_948715 ? add_950049 : sel_950046;
  assign add_950053 = sel_950050 + 8'h01;
  assign sel_950054 = array_index_949897 == array_index_948721 ? add_950053 : sel_950050;
  assign add_950057 = sel_950054 + 8'h01;
  assign sel_950058 = array_index_949897 == array_index_948727 ? add_950057 : sel_950054;
  assign add_950061 = sel_950058 + 8'h01;
  assign sel_950062 = array_index_949897 == array_index_948733 ? add_950061 : sel_950058;
  assign add_950065 = sel_950062 + 8'h01;
  assign sel_950066 = array_index_949897 == array_index_948739 ? add_950065 : sel_950062;
  assign add_950069 = sel_950066 + 8'h01;
  assign sel_950070 = array_index_949897 == array_index_948745 ? add_950069 : sel_950066;
  assign add_950073 = sel_950070 + 8'h01;
  assign sel_950074 = array_index_949897 == array_index_948751 ? add_950073 : sel_950070;
  assign add_950077 = sel_950074 + 8'h01;
  assign sel_950078 = array_index_949897 == array_index_948757 ? add_950077 : sel_950074;
  assign add_950081 = sel_950078 + 8'h01;
  assign sel_950082 = array_index_949897 == array_index_948763 ? add_950081 : sel_950078;
  assign add_950085 = sel_950082 + 8'h01;
  assign sel_950086 = array_index_949897 == array_index_948769 ? add_950085 : sel_950082;
  assign add_950089 = sel_950086 + 8'h01;
  assign sel_950090 = array_index_949897 == array_index_948775 ? add_950089 : sel_950086;
  assign add_950093 = sel_950090 + 8'h01;
  assign sel_950094 = array_index_949897 == array_index_948781 ? add_950093 : sel_950090;
  assign add_950097 = sel_950094 + 8'h01;
  assign sel_950098 = array_index_949897 == array_index_948787 ? add_950097 : sel_950094;
  assign add_950101 = sel_950098 + 8'h01;
  assign sel_950102 = array_index_949897 == array_index_948793 ? add_950101 : sel_950098;
  assign add_950105 = sel_950102 + 8'h01;
  assign sel_950106 = array_index_949897 == array_index_948799 ? add_950105 : sel_950102;
  assign add_950109 = sel_950106 + 8'h01;
  assign sel_950110 = array_index_949897 == array_index_948805 ? add_950109 : sel_950106;
  assign add_950113 = sel_950110 + 8'h01;
  assign sel_950114 = array_index_949897 == array_index_948811 ? add_950113 : sel_950110;
  assign add_950117 = sel_950114 + 8'h01;
  assign sel_950118 = array_index_949897 == array_index_948817 ? add_950117 : sel_950114;
  assign add_950121 = sel_950118 + 8'h01;
  assign sel_950122 = array_index_949897 == array_index_948823 ? add_950121 : sel_950118;
  assign add_950125 = sel_950122 + 8'h01;
  assign sel_950126 = array_index_949897 == array_index_948829 ? add_950125 : sel_950122;
  assign add_950129 = sel_950126 + 8'h01;
  assign sel_950130 = array_index_949897 == array_index_948835 ? add_950129 : sel_950126;
  assign add_950133 = sel_950130 + 8'h01;
  assign sel_950134 = array_index_949897 == array_index_948841 ? add_950133 : sel_950130;
  assign add_950137 = sel_950134 + 8'h01;
  assign sel_950138 = array_index_949897 == array_index_948847 ? add_950137 : sel_950134;
  assign add_950141 = sel_950138 + 8'h01;
  assign sel_950142 = array_index_949897 == array_index_948853 ? add_950141 : sel_950138;
  assign add_950145 = sel_950142 + 8'h01;
  assign sel_950146 = array_index_949897 == array_index_948859 ? add_950145 : sel_950142;
  assign add_950149 = sel_950146 + 8'h01;
  assign sel_950150 = array_index_949897 == array_index_948865 ? add_950149 : sel_950146;
  assign add_950153 = sel_950150 + 8'h01;
  assign sel_950154 = array_index_949897 == array_index_948871 ? add_950153 : sel_950150;
  assign add_950157 = sel_950154 + 8'h01;
  assign sel_950158 = array_index_949897 == array_index_948877 ? add_950157 : sel_950154;
  assign add_950161 = sel_950158 + 8'h01;
  assign sel_950162 = array_index_949897 == array_index_948883 ? add_950161 : sel_950158;
  assign add_950165 = sel_950162 + 8'h01;
  assign sel_950166 = array_index_949897 == array_index_948889 ? add_950165 : sel_950162;
  assign add_950169 = sel_950166 + 8'h01;
  assign sel_950170 = array_index_949897 == array_index_948895 ? add_950169 : sel_950166;
  assign add_950173 = sel_950170 + 8'h01;
  assign sel_950174 = array_index_949897 == array_index_948901 ? add_950173 : sel_950170;
  assign add_950177 = sel_950174 + 8'h01;
  assign sel_950178 = array_index_949897 == array_index_948907 ? add_950177 : sel_950174;
  assign add_950181 = sel_950178 + 8'h01;
  assign sel_950182 = array_index_949897 == array_index_948913 ? add_950181 : sel_950178;
  assign add_950185 = sel_950182 + 8'h01;
  assign sel_950186 = array_index_949897 == array_index_948919 ? add_950185 : sel_950182;
  assign add_950189 = sel_950186 + 8'h01;
  assign sel_950190 = array_index_949897 == array_index_948925 ? add_950189 : sel_950186;
  assign add_950193 = sel_950190 + 8'h01;
  assign sel_950194 = array_index_949897 == array_index_948931 ? add_950193 : sel_950190;
  assign add_950197 = sel_950194 + 8'h01;
  assign sel_950198 = array_index_949897 == array_index_948937 ? add_950197 : sel_950194;
  assign add_950201 = sel_950198 + 8'h01;
  assign sel_950202 = array_index_949897 == array_index_948943 ? add_950201 : sel_950198;
  assign add_950205 = sel_950202 + 8'h01;
  assign sel_950206 = array_index_949897 == array_index_948949 ? add_950205 : sel_950202;
  assign add_950209 = sel_950206 + 8'h01;
  assign sel_950210 = array_index_949897 == array_index_948955 ? add_950209 : sel_950206;
  assign add_950213 = sel_950210 + 8'h01;
  assign sel_950214 = array_index_949897 == array_index_948961 ? add_950213 : sel_950210;
  assign add_950217 = sel_950214 + 8'h01;
  assign sel_950218 = array_index_949897 == array_index_948967 ? add_950217 : sel_950214;
  assign add_950221 = sel_950218 + 8'h01;
  assign sel_950222 = array_index_949897 == array_index_948973 ? add_950221 : sel_950218;
  assign add_950225 = sel_950222 + 8'h01;
  assign sel_950226 = array_index_949897 == array_index_948979 ? add_950225 : sel_950222;
  assign add_950229 = sel_950226 + 8'h01;
  assign sel_950230 = array_index_949897 == array_index_948985 ? add_950229 : sel_950226;
  assign add_950233 = sel_950230 + 8'h01;
  assign sel_950234 = array_index_949897 == array_index_948991 ? add_950233 : sel_950230;
  assign add_950237 = sel_950234 + 8'h01;
  assign sel_950238 = array_index_949897 == array_index_948997 ? add_950237 : sel_950234;
  assign add_950241 = sel_950238 + 8'h01;
  assign sel_950242 = array_index_949897 == array_index_949003 ? add_950241 : sel_950238;
  assign add_950245 = sel_950242 + 8'h01;
  assign sel_950246 = array_index_949897 == array_index_949009 ? add_950245 : sel_950242;
  assign add_950249 = sel_950246 + 8'h01;
  assign sel_950250 = array_index_949897 == array_index_949015 ? add_950249 : sel_950246;
  assign add_950253 = sel_950250 + 8'h01;
  assign sel_950254 = array_index_949897 == array_index_949021 ? add_950253 : sel_950250;
  assign add_950257 = sel_950254 + 8'h01;
  assign sel_950258 = array_index_949897 == array_index_949027 ? add_950257 : sel_950254;
  assign add_950261 = sel_950258 + 8'h01;
  assign sel_950262 = array_index_949897 == array_index_949033 ? add_950261 : sel_950258;
  assign add_950265 = sel_950262 + 8'h01;
  assign sel_950266 = array_index_949897 == array_index_949039 ? add_950265 : sel_950262;
  assign add_950269 = sel_950266 + 8'h01;
  assign sel_950270 = array_index_949897 == array_index_949045 ? add_950269 : sel_950266;
  assign add_950273 = sel_950270 + 8'h01;
  assign sel_950274 = array_index_949897 == array_index_949051 ? add_950273 : sel_950270;
  assign add_950277 = sel_950274 + 8'h01;
  assign sel_950278 = array_index_949897 == array_index_949057 ? add_950277 : sel_950274;
  assign add_950281 = sel_950278 + 8'h01;
  assign sel_950282 = array_index_949897 == array_index_949063 ? add_950281 : sel_950278;
  assign add_950285 = sel_950282 + 8'h01;
  assign sel_950286 = array_index_949897 == array_index_949069 ? add_950285 : sel_950282;
  assign add_950289 = sel_950286 + 8'h01;
  assign sel_950290 = array_index_949897 == array_index_949075 ? add_950289 : sel_950286;
  assign add_950293 = sel_950290 + 8'h01;
  assign sel_950294 = array_index_949897 == array_index_949081 ? add_950293 : sel_950290;
  assign add_950298 = sel_950294 + 8'h01;
  assign array_index_950299 = set1_unflattened[7'h04];
  assign sel_950300 = array_index_949897 == array_index_949087 ? add_950298 : sel_950294;
  assign add_950303 = sel_950300 + 8'h01;
  assign sel_950304 = array_index_950299 == array_index_948483 ? add_950303 : sel_950300;
  assign add_950307 = sel_950304 + 8'h01;
  assign sel_950308 = array_index_950299 == array_index_948487 ? add_950307 : sel_950304;
  assign add_950311 = sel_950308 + 8'h01;
  assign sel_950312 = array_index_950299 == array_index_948495 ? add_950311 : sel_950308;
  assign add_950315 = sel_950312 + 8'h01;
  assign sel_950316 = array_index_950299 == array_index_948503 ? add_950315 : sel_950312;
  assign add_950319 = sel_950316 + 8'h01;
  assign sel_950320 = array_index_950299 == array_index_948511 ? add_950319 : sel_950316;
  assign add_950323 = sel_950320 + 8'h01;
  assign sel_950324 = array_index_950299 == array_index_948519 ? add_950323 : sel_950320;
  assign add_950327 = sel_950324 + 8'h01;
  assign sel_950328 = array_index_950299 == array_index_948527 ? add_950327 : sel_950324;
  assign add_950331 = sel_950328 + 8'h01;
  assign sel_950332 = array_index_950299 == array_index_948535 ? add_950331 : sel_950328;
  assign add_950335 = sel_950332 + 8'h01;
  assign sel_950336 = array_index_950299 == array_index_948541 ? add_950335 : sel_950332;
  assign add_950339 = sel_950336 + 8'h01;
  assign sel_950340 = array_index_950299 == array_index_948547 ? add_950339 : sel_950336;
  assign add_950343 = sel_950340 + 8'h01;
  assign sel_950344 = array_index_950299 == array_index_948553 ? add_950343 : sel_950340;
  assign add_950347 = sel_950344 + 8'h01;
  assign sel_950348 = array_index_950299 == array_index_948559 ? add_950347 : sel_950344;
  assign add_950351 = sel_950348 + 8'h01;
  assign sel_950352 = array_index_950299 == array_index_948565 ? add_950351 : sel_950348;
  assign add_950355 = sel_950352 + 8'h01;
  assign sel_950356 = array_index_950299 == array_index_948571 ? add_950355 : sel_950352;
  assign add_950359 = sel_950356 + 8'h01;
  assign sel_950360 = array_index_950299 == array_index_948577 ? add_950359 : sel_950356;
  assign add_950363 = sel_950360 + 8'h01;
  assign sel_950364 = array_index_950299 == array_index_948583 ? add_950363 : sel_950360;
  assign add_950367 = sel_950364 + 8'h01;
  assign sel_950368 = array_index_950299 == array_index_948589 ? add_950367 : sel_950364;
  assign add_950371 = sel_950368 + 8'h01;
  assign sel_950372 = array_index_950299 == array_index_948595 ? add_950371 : sel_950368;
  assign add_950375 = sel_950372 + 8'h01;
  assign sel_950376 = array_index_950299 == array_index_948601 ? add_950375 : sel_950372;
  assign add_950379 = sel_950376 + 8'h01;
  assign sel_950380 = array_index_950299 == array_index_948607 ? add_950379 : sel_950376;
  assign add_950383 = sel_950380 + 8'h01;
  assign sel_950384 = array_index_950299 == array_index_948613 ? add_950383 : sel_950380;
  assign add_950387 = sel_950384 + 8'h01;
  assign sel_950388 = array_index_950299 == array_index_948619 ? add_950387 : sel_950384;
  assign add_950391 = sel_950388 + 8'h01;
  assign sel_950392 = array_index_950299 == array_index_948625 ? add_950391 : sel_950388;
  assign add_950395 = sel_950392 + 8'h01;
  assign sel_950396 = array_index_950299 == array_index_948631 ? add_950395 : sel_950392;
  assign add_950399 = sel_950396 + 8'h01;
  assign sel_950400 = array_index_950299 == array_index_948637 ? add_950399 : sel_950396;
  assign add_950403 = sel_950400 + 8'h01;
  assign sel_950404 = array_index_950299 == array_index_948643 ? add_950403 : sel_950400;
  assign add_950407 = sel_950404 + 8'h01;
  assign sel_950408 = array_index_950299 == array_index_948649 ? add_950407 : sel_950404;
  assign add_950411 = sel_950408 + 8'h01;
  assign sel_950412 = array_index_950299 == array_index_948655 ? add_950411 : sel_950408;
  assign add_950415 = sel_950412 + 8'h01;
  assign sel_950416 = array_index_950299 == array_index_948661 ? add_950415 : sel_950412;
  assign add_950419 = sel_950416 + 8'h01;
  assign sel_950420 = array_index_950299 == array_index_948667 ? add_950419 : sel_950416;
  assign add_950423 = sel_950420 + 8'h01;
  assign sel_950424 = array_index_950299 == array_index_948673 ? add_950423 : sel_950420;
  assign add_950427 = sel_950424 + 8'h01;
  assign sel_950428 = array_index_950299 == array_index_948679 ? add_950427 : sel_950424;
  assign add_950431 = sel_950428 + 8'h01;
  assign sel_950432 = array_index_950299 == array_index_948685 ? add_950431 : sel_950428;
  assign add_950435 = sel_950432 + 8'h01;
  assign sel_950436 = array_index_950299 == array_index_948691 ? add_950435 : sel_950432;
  assign add_950439 = sel_950436 + 8'h01;
  assign sel_950440 = array_index_950299 == array_index_948697 ? add_950439 : sel_950436;
  assign add_950443 = sel_950440 + 8'h01;
  assign sel_950444 = array_index_950299 == array_index_948703 ? add_950443 : sel_950440;
  assign add_950447 = sel_950444 + 8'h01;
  assign sel_950448 = array_index_950299 == array_index_948709 ? add_950447 : sel_950444;
  assign add_950451 = sel_950448 + 8'h01;
  assign sel_950452 = array_index_950299 == array_index_948715 ? add_950451 : sel_950448;
  assign add_950455 = sel_950452 + 8'h01;
  assign sel_950456 = array_index_950299 == array_index_948721 ? add_950455 : sel_950452;
  assign add_950459 = sel_950456 + 8'h01;
  assign sel_950460 = array_index_950299 == array_index_948727 ? add_950459 : sel_950456;
  assign add_950463 = sel_950460 + 8'h01;
  assign sel_950464 = array_index_950299 == array_index_948733 ? add_950463 : sel_950460;
  assign add_950467 = sel_950464 + 8'h01;
  assign sel_950468 = array_index_950299 == array_index_948739 ? add_950467 : sel_950464;
  assign add_950471 = sel_950468 + 8'h01;
  assign sel_950472 = array_index_950299 == array_index_948745 ? add_950471 : sel_950468;
  assign add_950475 = sel_950472 + 8'h01;
  assign sel_950476 = array_index_950299 == array_index_948751 ? add_950475 : sel_950472;
  assign add_950479 = sel_950476 + 8'h01;
  assign sel_950480 = array_index_950299 == array_index_948757 ? add_950479 : sel_950476;
  assign add_950483 = sel_950480 + 8'h01;
  assign sel_950484 = array_index_950299 == array_index_948763 ? add_950483 : sel_950480;
  assign add_950487 = sel_950484 + 8'h01;
  assign sel_950488 = array_index_950299 == array_index_948769 ? add_950487 : sel_950484;
  assign add_950491 = sel_950488 + 8'h01;
  assign sel_950492 = array_index_950299 == array_index_948775 ? add_950491 : sel_950488;
  assign add_950495 = sel_950492 + 8'h01;
  assign sel_950496 = array_index_950299 == array_index_948781 ? add_950495 : sel_950492;
  assign add_950499 = sel_950496 + 8'h01;
  assign sel_950500 = array_index_950299 == array_index_948787 ? add_950499 : sel_950496;
  assign add_950503 = sel_950500 + 8'h01;
  assign sel_950504 = array_index_950299 == array_index_948793 ? add_950503 : sel_950500;
  assign add_950507 = sel_950504 + 8'h01;
  assign sel_950508 = array_index_950299 == array_index_948799 ? add_950507 : sel_950504;
  assign add_950511 = sel_950508 + 8'h01;
  assign sel_950512 = array_index_950299 == array_index_948805 ? add_950511 : sel_950508;
  assign add_950515 = sel_950512 + 8'h01;
  assign sel_950516 = array_index_950299 == array_index_948811 ? add_950515 : sel_950512;
  assign add_950519 = sel_950516 + 8'h01;
  assign sel_950520 = array_index_950299 == array_index_948817 ? add_950519 : sel_950516;
  assign add_950523 = sel_950520 + 8'h01;
  assign sel_950524 = array_index_950299 == array_index_948823 ? add_950523 : sel_950520;
  assign add_950527 = sel_950524 + 8'h01;
  assign sel_950528 = array_index_950299 == array_index_948829 ? add_950527 : sel_950524;
  assign add_950531 = sel_950528 + 8'h01;
  assign sel_950532 = array_index_950299 == array_index_948835 ? add_950531 : sel_950528;
  assign add_950535 = sel_950532 + 8'h01;
  assign sel_950536 = array_index_950299 == array_index_948841 ? add_950535 : sel_950532;
  assign add_950539 = sel_950536 + 8'h01;
  assign sel_950540 = array_index_950299 == array_index_948847 ? add_950539 : sel_950536;
  assign add_950543 = sel_950540 + 8'h01;
  assign sel_950544 = array_index_950299 == array_index_948853 ? add_950543 : sel_950540;
  assign add_950547 = sel_950544 + 8'h01;
  assign sel_950548 = array_index_950299 == array_index_948859 ? add_950547 : sel_950544;
  assign add_950551 = sel_950548 + 8'h01;
  assign sel_950552 = array_index_950299 == array_index_948865 ? add_950551 : sel_950548;
  assign add_950555 = sel_950552 + 8'h01;
  assign sel_950556 = array_index_950299 == array_index_948871 ? add_950555 : sel_950552;
  assign add_950559 = sel_950556 + 8'h01;
  assign sel_950560 = array_index_950299 == array_index_948877 ? add_950559 : sel_950556;
  assign add_950563 = sel_950560 + 8'h01;
  assign sel_950564 = array_index_950299 == array_index_948883 ? add_950563 : sel_950560;
  assign add_950567 = sel_950564 + 8'h01;
  assign sel_950568 = array_index_950299 == array_index_948889 ? add_950567 : sel_950564;
  assign add_950571 = sel_950568 + 8'h01;
  assign sel_950572 = array_index_950299 == array_index_948895 ? add_950571 : sel_950568;
  assign add_950575 = sel_950572 + 8'h01;
  assign sel_950576 = array_index_950299 == array_index_948901 ? add_950575 : sel_950572;
  assign add_950579 = sel_950576 + 8'h01;
  assign sel_950580 = array_index_950299 == array_index_948907 ? add_950579 : sel_950576;
  assign add_950583 = sel_950580 + 8'h01;
  assign sel_950584 = array_index_950299 == array_index_948913 ? add_950583 : sel_950580;
  assign add_950587 = sel_950584 + 8'h01;
  assign sel_950588 = array_index_950299 == array_index_948919 ? add_950587 : sel_950584;
  assign add_950591 = sel_950588 + 8'h01;
  assign sel_950592 = array_index_950299 == array_index_948925 ? add_950591 : sel_950588;
  assign add_950595 = sel_950592 + 8'h01;
  assign sel_950596 = array_index_950299 == array_index_948931 ? add_950595 : sel_950592;
  assign add_950599 = sel_950596 + 8'h01;
  assign sel_950600 = array_index_950299 == array_index_948937 ? add_950599 : sel_950596;
  assign add_950603 = sel_950600 + 8'h01;
  assign sel_950604 = array_index_950299 == array_index_948943 ? add_950603 : sel_950600;
  assign add_950607 = sel_950604 + 8'h01;
  assign sel_950608 = array_index_950299 == array_index_948949 ? add_950607 : sel_950604;
  assign add_950611 = sel_950608 + 8'h01;
  assign sel_950612 = array_index_950299 == array_index_948955 ? add_950611 : sel_950608;
  assign add_950615 = sel_950612 + 8'h01;
  assign sel_950616 = array_index_950299 == array_index_948961 ? add_950615 : sel_950612;
  assign add_950619 = sel_950616 + 8'h01;
  assign sel_950620 = array_index_950299 == array_index_948967 ? add_950619 : sel_950616;
  assign add_950623 = sel_950620 + 8'h01;
  assign sel_950624 = array_index_950299 == array_index_948973 ? add_950623 : sel_950620;
  assign add_950627 = sel_950624 + 8'h01;
  assign sel_950628 = array_index_950299 == array_index_948979 ? add_950627 : sel_950624;
  assign add_950631 = sel_950628 + 8'h01;
  assign sel_950632 = array_index_950299 == array_index_948985 ? add_950631 : sel_950628;
  assign add_950635 = sel_950632 + 8'h01;
  assign sel_950636 = array_index_950299 == array_index_948991 ? add_950635 : sel_950632;
  assign add_950639 = sel_950636 + 8'h01;
  assign sel_950640 = array_index_950299 == array_index_948997 ? add_950639 : sel_950636;
  assign add_950643 = sel_950640 + 8'h01;
  assign sel_950644 = array_index_950299 == array_index_949003 ? add_950643 : sel_950640;
  assign add_950647 = sel_950644 + 8'h01;
  assign sel_950648 = array_index_950299 == array_index_949009 ? add_950647 : sel_950644;
  assign add_950651 = sel_950648 + 8'h01;
  assign sel_950652 = array_index_950299 == array_index_949015 ? add_950651 : sel_950648;
  assign add_950655 = sel_950652 + 8'h01;
  assign sel_950656 = array_index_950299 == array_index_949021 ? add_950655 : sel_950652;
  assign add_950659 = sel_950656 + 8'h01;
  assign sel_950660 = array_index_950299 == array_index_949027 ? add_950659 : sel_950656;
  assign add_950663 = sel_950660 + 8'h01;
  assign sel_950664 = array_index_950299 == array_index_949033 ? add_950663 : sel_950660;
  assign add_950667 = sel_950664 + 8'h01;
  assign sel_950668 = array_index_950299 == array_index_949039 ? add_950667 : sel_950664;
  assign add_950671 = sel_950668 + 8'h01;
  assign sel_950672 = array_index_950299 == array_index_949045 ? add_950671 : sel_950668;
  assign add_950675 = sel_950672 + 8'h01;
  assign sel_950676 = array_index_950299 == array_index_949051 ? add_950675 : sel_950672;
  assign add_950679 = sel_950676 + 8'h01;
  assign sel_950680 = array_index_950299 == array_index_949057 ? add_950679 : sel_950676;
  assign add_950683 = sel_950680 + 8'h01;
  assign sel_950684 = array_index_950299 == array_index_949063 ? add_950683 : sel_950680;
  assign add_950687 = sel_950684 + 8'h01;
  assign sel_950688 = array_index_950299 == array_index_949069 ? add_950687 : sel_950684;
  assign add_950691 = sel_950688 + 8'h01;
  assign sel_950692 = array_index_950299 == array_index_949075 ? add_950691 : sel_950688;
  assign add_950695 = sel_950692 + 8'h01;
  assign sel_950696 = array_index_950299 == array_index_949081 ? add_950695 : sel_950692;
  assign add_950700 = sel_950696 + 8'h01;
  assign array_index_950701 = set1_unflattened[7'h05];
  assign sel_950702 = array_index_950299 == array_index_949087 ? add_950700 : sel_950696;
  assign add_950705 = sel_950702 + 8'h01;
  assign sel_950706 = array_index_950701 == array_index_948483 ? add_950705 : sel_950702;
  assign add_950709 = sel_950706 + 8'h01;
  assign sel_950710 = array_index_950701 == array_index_948487 ? add_950709 : sel_950706;
  assign add_950713 = sel_950710 + 8'h01;
  assign sel_950714 = array_index_950701 == array_index_948495 ? add_950713 : sel_950710;
  assign add_950717 = sel_950714 + 8'h01;
  assign sel_950718 = array_index_950701 == array_index_948503 ? add_950717 : sel_950714;
  assign add_950721 = sel_950718 + 8'h01;
  assign sel_950722 = array_index_950701 == array_index_948511 ? add_950721 : sel_950718;
  assign add_950725 = sel_950722 + 8'h01;
  assign sel_950726 = array_index_950701 == array_index_948519 ? add_950725 : sel_950722;
  assign add_950729 = sel_950726 + 8'h01;
  assign sel_950730 = array_index_950701 == array_index_948527 ? add_950729 : sel_950726;
  assign add_950733 = sel_950730 + 8'h01;
  assign sel_950734 = array_index_950701 == array_index_948535 ? add_950733 : sel_950730;
  assign add_950737 = sel_950734 + 8'h01;
  assign sel_950738 = array_index_950701 == array_index_948541 ? add_950737 : sel_950734;
  assign add_950741 = sel_950738 + 8'h01;
  assign sel_950742 = array_index_950701 == array_index_948547 ? add_950741 : sel_950738;
  assign add_950745 = sel_950742 + 8'h01;
  assign sel_950746 = array_index_950701 == array_index_948553 ? add_950745 : sel_950742;
  assign add_950749 = sel_950746 + 8'h01;
  assign sel_950750 = array_index_950701 == array_index_948559 ? add_950749 : sel_950746;
  assign add_950753 = sel_950750 + 8'h01;
  assign sel_950754 = array_index_950701 == array_index_948565 ? add_950753 : sel_950750;
  assign add_950757 = sel_950754 + 8'h01;
  assign sel_950758 = array_index_950701 == array_index_948571 ? add_950757 : sel_950754;
  assign add_950761 = sel_950758 + 8'h01;
  assign sel_950762 = array_index_950701 == array_index_948577 ? add_950761 : sel_950758;
  assign add_950765 = sel_950762 + 8'h01;
  assign sel_950766 = array_index_950701 == array_index_948583 ? add_950765 : sel_950762;
  assign add_950769 = sel_950766 + 8'h01;
  assign sel_950770 = array_index_950701 == array_index_948589 ? add_950769 : sel_950766;
  assign add_950773 = sel_950770 + 8'h01;
  assign sel_950774 = array_index_950701 == array_index_948595 ? add_950773 : sel_950770;
  assign add_950777 = sel_950774 + 8'h01;
  assign sel_950778 = array_index_950701 == array_index_948601 ? add_950777 : sel_950774;
  assign add_950781 = sel_950778 + 8'h01;
  assign sel_950782 = array_index_950701 == array_index_948607 ? add_950781 : sel_950778;
  assign add_950785 = sel_950782 + 8'h01;
  assign sel_950786 = array_index_950701 == array_index_948613 ? add_950785 : sel_950782;
  assign add_950789 = sel_950786 + 8'h01;
  assign sel_950790 = array_index_950701 == array_index_948619 ? add_950789 : sel_950786;
  assign add_950793 = sel_950790 + 8'h01;
  assign sel_950794 = array_index_950701 == array_index_948625 ? add_950793 : sel_950790;
  assign add_950797 = sel_950794 + 8'h01;
  assign sel_950798 = array_index_950701 == array_index_948631 ? add_950797 : sel_950794;
  assign add_950801 = sel_950798 + 8'h01;
  assign sel_950802 = array_index_950701 == array_index_948637 ? add_950801 : sel_950798;
  assign add_950805 = sel_950802 + 8'h01;
  assign sel_950806 = array_index_950701 == array_index_948643 ? add_950805 : sel_950802;
  assign add_950809 = sel_950806 + 8'h01;
  assign sel_950810 = array_index_950701 == array_index_948649 ? add_950809 : sel_950806;
  assign add_950813 = sel_950810 + 8'h01;
  assign sel_950814 = array_index_950701 == array_index_948655 ? add_950813 : sel_950810;
  assign add_950817 = sel_950814 + 8'h01;
  assign sel_950818 = array_index_950701 == array_index_948661 ? add_950817 : sel_950814;
  assign add_950821 = sel_950818 + 8'h01;
  assign sel_950822 = array_index_950701 == array_index_948667 ? add_950821 : sel_950818;
  assign add_950825 = sel_950822 + 8'h01;
  assign sel_950826 = array_index_950701 == array_index_948673 ? add_950825 : sel_950822;
  assign add_950829 = sel_950826 + 8'h01;
  assign sel_950830 = array_index_950701 == array_index_948679 ? add_950829 : sel_950826;
  assign add_950833 = sel_950830 + 8'h01;
  assign sel_950834 = array_index_950701 == array_index_948685 ? add_950833 : sel_950830;
  assign add_950837 = sel_950834 + 8'h01;
  assign sel_950838 = array_index_950701 == array_index_948691 ? add_950837 : sel_950834;
  assign add_950841 = sel_950838 + 8'h01;
  assign sel_950842 = array_index_950701 == array_index_948697 ? add_950841 : sel_950838;
  assign add_950845 = sel_950842 + 8'h01;
  assign sel_950846 = array_index_950701 == array_index_948703 ? add_950845 : sel_950842;
  assign add_950849 = sel_950846 + 8'h01;
  assign sel_950850 = array_index_950701 == array_index_948709 ? add_950849 : sel_950846;
  assign add_950853 = sel_950850 + 8'h01;
  assign sel_950854 = array_index_950701 == array_index_948715 ? add_950853 : sel_950850;
  assign add_950857 = sel_950854 + 8'h01;
  assign sel_950858 = array_index_950701 == array_index_948721 ? add_950857 : sel_950854;
  assign add_950861 = sel_950858 + 8'h01;
  assign sel_950862 = array_index_950701 == array_index_948727 ? add_950861 : sel_950858;
  assign add_950865 = sel_950862 + 8'h01;
  assign sel_950866 = array_index_950701 == array_index_948733 ? add_950865 : sel_950862;
  assign add_950869 = sel_950866 + 8'h01;
  assign sel_950870 = array_index_950701 == array_index_948739 ? add_950869 : sel_950866;
  assign add_950873 = sel_950870 + 8'h01;
  assign sel_950874 = array_index_950701 == array_index_948745 ? add_950873 : sel_950870;
  assign add_950877 = sel_950874 + 8'h01;
  assign sel_950878 = array_index_950701 == array_index_948751 ? add_950877 : sel_950874;
  assign add_950881 = sel_950878 + 8'h01;
  assign sel_950882 = array_index_950701 == array_index_948757 ? add_950881 : sel_950878;
  assign add_950885 = sel_950882 + 8'h01;
  assign sel_950886 = array_index_950701 == array_index_948763 ? add_950885 : sel_950882;
  assign add_950889 = sel_950886 + 8'h01;
  assign sel_950890 = array_index_950701 == array_index_948769 ? add_950889 : sel_950886;
  assign add_950893 = sel_950890 + 8'h01;
  assign sel_950894 = array_index_950701 == array_index_948775 ? add_950893 : sel_950890;
  assign add_950897 = sel_950894 + 8'h01;
  assign sel_950898 = array_index_950701 == array_index_948781 ? add_950897 : sel_950894;
  assign add_950901 = sel_950898 + 8'h01;
  assign sel_950902 = array_index_950701 == array_index_948787 ? add_950901 : sel_950898;
  assign add_950905 = sel_950902 + 8'h01;
  assign sel_950906 = array_index_950701 == array_index_948793 ? add_950905 : sel_950902;
  assign add_950909 = sel_950906 + 8'h01;
  assign sel_950910 = array_index_950701 == array_index_948799 ? add_950909 : sel_950906;
  assign add_950913 = sel_950910 + 8'h01;
  assign sel_950914 = array_index_950701 == array_index_948805 ? add_950913 : sel_950910;
  assign add_950917 = sel_950914 + 8'h01;
  assign sel_950918 = array_index_950701 == array_index_948811 ? add_950917 : sel_950914;
  assign add_950921 = sel_950918 + 8'h01;
  assign sel_950922 = array_index_950701 == array_index_948817 ? add_950921 : sel_950918;
  assign add_950925 = sel_950922 + 8'h01;
  assign sel_950926 = array_index_950701 == array_index_948823 ? add_950925 : sel_950922;
  assign add_950929 = sel_950926 + 8'h01;
  assign sel_950930 = array_index_950701 == array_index_948829 ? add_950929 : sel_950926;
  assign add_950933 = sel_950930 + 8'h01;
  assign sel_950934 = array_index_950701 == array_index_948835 ? add_950933 : sel_950930;
  assign add_950937 = sel_950934 + 8'h01;
  assign sel_950938 = array_index_950701 == array_index_948841 ? add_950937 : sel_950934;
  assign add_950941 = sel_950938 + 8'h01;
  assign sel_950942 = array_index_950701 == array_index_948847 ? add_950941 : sel_950938;
  assign add_950945 = sel_950942 + 8'h01;
  assign sel_950946 = array_index_950701 == array_index_948853 ? add_950945 : sel_950942;
  assign add_950949 = sel_950946 + 8'h01;
  assign sel_950950 = array_index_950701 == array_index_948859 ? add_950949 : sel_950946;
  assign add_950953 = sel_950950 + 8'h01;
  assign sel_950954 = array_index_950701 == array_index_948865 ? add_950953 : sel_950950;
  assign add_950957 = sel_950954 + 8'h01;
  assign sel_950958 = array_index_950701 == array_index_948871 ? add_950957 : sel_950954;
  assign add_950961 = sel_950958 + 8'h01;
  assign sel_950962 = array_index_950701 == array_index_948877 ? add_950961 : sel_950958;
  assign add_950965 = sel_950962 + 8'h01;
  assign sel_950966 = array_index_950701 == array_index_948883 ? add_950965 : sel_950962;
  assign add_950969 = sel_950966 + 8'h01;
  assign sel_950970 = array_index_950701 == array_index_948889 ? add_950969 : sel_950966;
  assign add_950973 = sel_950970 + 8'h01;
  assign sel_950974 = array_index_950701 == array_index_948895 ? add_950973 : sel_950970;
  assign add_950977 = sel_950974 + 8'h01;
  assign sel_950978 = array_index_950701 == array_index_948901 ? add_950977 : sel_950974;
  assign add_950981 = sel_950978 + 8'h01;
  assign sel_950982 = array_index_950701 == array_index_948907 ? add_950981 : sel_950978;
  assign add_950985 = sel_950982 + 8'h01;
  assign sel_950986 = array_index_950701 == array_index_948913 ? add_950985 : sel_950982;
  assign add_950989 = sel_950986 + 8'h01;
  assign sel_950990 = array_index_950701 == array_index_948919 ? add_950989 : sel_950986;
  assign add_950993 = sel_950990 + 8'h01;
  assign sel_950994 = array_index_950701 == array_index_948925 ? add_950993 : sel_950990;
  assign add_950997 = sel_950994 + 8'h01;
  assign sel_950998 = array_index_950701 == array_index_948931 ? add_950997 : sel_950994;
  assign add_951001 = sel_950998 + 8'h01;
  assign sel_951002 = array_index_950701 == array_index_948937 ? add_951001 : sel_950998;
  assign add_951005 = sel_951002 + 8'h01;
  assign sel_951006 = array_index_950701 == array_index_948943 ? add_951005 : sel_951002;
  assign add_951009 = sel_951006 + 8'h01;
  assign sel_951010 = array_index_950701 == array_index_948949 ? add_951009 : sel_951006;
  assign add_951013 = sel_951010 + 8'h01;
  assign sel_951014 = array_index_950701 == array_index_948955 ? add_951013 : sel_951010;
  assign add_951017 = sel_951014 + 8'h01;
  assign sel_951018 = array_index_950701 == array_index_948961 ? add_951017 : sel_951014;
  assign add_951021 = sel_951018 + 8'h01;
  assign sel_951022 = array_index_950701 == array_index_948967 ? add_951021 : sel_951018;
  assign add_951025 = sel_951022 + 8'h01;
  assign sel_951026 = array_index_950701 == array_index_948973 ? add_951025 : sel_951022;
  assign add_951029 = sel_951026 + 8'h01;
  assign sel_951030 = array_index_950701 == array_index_948979 ? add_951029 : sel_951026;
  assign add_951033 = sel_951030 + 8'h01;
  assign sel_951034 = array_index_950701 == array_index_948985 ? add_951033 : sel_951030;
  assign add_951037 = sel_951034 + 8'h01;
  assign sel_951038 = array_index_950701 == array_index_948991 ? add_951037 : sel_951034;
  assign add_951041 = sel_951038 + 8'h01;
  assign sel_951042 = array_index_950701 == array_index_948997 ? add_951041 : sel_951038;
  assign add_951045 = sel_951042 + 8'h01;
  assign sel_951046 = array_index_950701 == array_index_949003 ? add_951045 : sel_951042;
  assign add_951049 = sel_951046 + 8'h01;
  assign sel_951050 = array_index_950701 == array_index_949009 ? add_951049 : sel_951046;
  assign add_951053 = sel_951050 + 8'h01;
  assign sel_951054 = array_index_950701 == array_index_949015 ? add_951053 : sel_951050;
  assign add_951057 = sel_951054 + 8'h01;
  assign sel_951058 = array_index_950701 == array_index_949021 ? add_951057 : sel_951054;
  assign add_951061 = sel_951058 + 8'h01;
  assign sel_951062 = array_index_950701 == array_index_949027 ? add_951061 : sel_951058;
  assign add_951065 = sel_951062 + 8'h01;
  assign sel_951066 = array_index_950701 == array_index_949033 ? add_951065 : sel_951062;
  assign add_951069 = sel_951066 + 8'h01;
  assign sel_951070 = array_index_950701 == array_index_949039 ? add_951069 : sel_951066;
  assign add_951073 = sel_951070 + 8'h01;
  assign sel_951074 = array_index_950701 == array_index_949045 ? add_951073 : sel_951070;
  assign add_951077 = sel_951074 + 8'h01;
  assign sel_951078 = array_index_950701 == array_index_949051 ? add_951077 : sel_951074;
  assign add_951081 = sel_951078 + 8'h01;
  assign sel_951082 = array_index_950701 == array_index_949057 ? add_951081 : sel_951078;
  assign add_951085 = sel_951082 + 8'h01;
  assign sel_951086 = array_index_950701 == array_index_949063 ? add_951085 : sel_951082;
  assign add_951089 = sel_951086 + 8'h01;
  assign sel_951090 = array_index_950701 == array_index_949069 ? add_951089 : sel_951086;
  assign add_951093 = sel_951090 + 8'h01;
  assign sel_951094 = array_index_950701 == array_index_949075 ? add_951093 : sel_951090;
  assign add_951097 = sel_951094 + 8'h01;
  assign sel_951098 = array_index_950701 == array_index_949081 ? add_951097 : sel_951094;
  assign add_951102 = sel_951098 + 8'h01;
  assign array_index_951103 = set1_unflattened[7'h06];
  assign sel_951104 = array_index_950701 == array_index_949087 ? add_951102 : sel_951098;
  assign add_951107 = sel_951104 + 8'h01;
  assign sel_951108 = array_index_951103 == array_index_948483 ? add_951107 : sel_951104;
  assign add_951111 = sel_951108 + 8'h01;
  assign sel_951112 = array_index_951103 == array_index_948487 ? add_951111 : sel_951108;
  assign add_951115 = sel_951112 + 8'h01;
  assign sel_951116 = array_index_951103 == array_index_948495 ? add_951115 : sel_951112;
  assign add_951119 = sel_951116 + 8'h01;
  assign sel_951120 = array_index_951103 == array_index_948503 ? add_951119 : sel_951116;
  assign add_951123 = sel_951120 + 8'h01;
  assign sel_951124 = array_index_951103 == array_index_948511 ? add_951123 : sel_951120;
  assign add_951127 = sel_951124 + 8'h01;
  assign sel_951128 = array_index_951103 == array_index_948519 ? add_951127 : sel_951124;
  assign add_951131 = sel_951128 + 8'h01;
  assign sel_951132 = array_index_951103 == array_index_948527 ? add_951131 : sel_951128;
  assign add_951135 = sel_951132 + 8'h01;
  assign sel_951136 = array_index_951103 == array_index_948535 ? add_951135 : sel_951132;
  assign add_951139 = sel_951136 + 8'h01;
  assign sel_951140 = array_index_951103 == array_index_948541 ? add_951139 : sel_951136;
  assign add_951143 = sel_951140 + 8'h01;
  assign sel_951144 = array_index_951103 == array_index_948547 ? add_951143 : sel_951140;
  assign add_951147 = sel_951144 + 8'h01;
  assign sel_951148 = array_index_951103 == array_index_948553 ? add_951147 : sel_951144;
  assign add_951151 = sel_951148 + 8'h01;
  assign sel_951152 = array_index_951103 == array_index_948559 ? add_951151 : sel_951148;
  assign add_951155 = sel_951152 + 8'h01;
  assign sel_951156 = array_index_951103 == array_index_948565 ? add_951155 : sel_951152;
  assign add_951159 = sel_951156 + 8'h01;
  assign sel_951160 = array_index_951103 == array_index_948571 ? add_951159 : sel_951156;
  assign add_951163 = sel_951160 + 8'h01;
  assign sel_951164 = array_index_951103 == array_index_948577 ? add_951163 : sel_951160;
  assign add_951167 = sel_951164 + 8'h01;
  assign sel_951168 = array_index_951103 == array_index_948583 ? add_951167 : sel_951164;
  assign add_951171 = sel_951168 + 8'h01;
  assign sel_951172 = array_index_951103 == array_index_948589 ? add_951171 : sel_951168;
  assign add_951175 = sel_951172 + 8'h01;
  assign sel_951176 = array_index_951103 == array_index_948595 ? add_951175 : sel_951172;
  assign add_951179 = sel_951176 + 8'h01;
  assign sel_951180 = array_index_951103 == array_index_948601 ? add_951179 : sel_951176;
  assign add_951183 = sel_951180 + 8'h01;
  assign sel_951184 = array_index_951103 == array_index_948607 ? add_951183 : sel_951180;
  assign add_951187 = sel_951184 + 8'h01;
  assign sel_951188 = array_index_951103 == array_index_948613 ? add_951187 : sel_951184;
  assign add_951191 = sel_951188 + 8'h01;
  assign sel_951192 = array_index_951103 == array_index_948619 ? add_951191 : sel_951188;
  assign add_951195 = sel_951192 + 8'h01;
  assign sel_951196 = array_index_951103 == array_index_948625 ? add_951195 : sel_951192;
  assign add_951199 = sel_951196 + 8'h01;
  assign sel_951200 = array_index_951103 == array_index_948631 ? add_951199 : sel_951196;
  assign add_951203 = sel_951200 + 8'h01;
  assign sel_951204 = array_index_951103 == array_index_948637 ? add_951203 : sel_951200;
  assign add_951207 = sel_951204 + 8'h01;
  assign sel_951208 = array_index_951103 == array_index_948643 ? add_951207 : sel_951204;
  assign add_951211 = sel_951208 + 8'h01;
  assign sel_951212 = array_index_951103 == array_index_948649 ? add_951211 : sel_951208;
  assign add_951215 = sel_951212 + 8'h01;
  assign sel_951216 = array_index_951103 == array_index_948655 ? add_951215 : sel_951212;
  assign add_951219 = sel_951216 + 8'h01;
  assign sel_951220 = array_index_951103 == array_index_948661 ? add_951219 : sel_951216;
  assign add_951223 = sel_951220 + 8'h01;
  assign sel_951224 = array_index_951103 == array_index_948667 ? add_951223 : sel_951220;
  assign add_951227 = sel_951224 + 8'h01;
  assign sel_951228 = array_index_951103 == array_index_948673 ? add_951227 : sel_951224;
  assign add_951231 = sel_951228 + 8'h01;
  assign sel_951232 = array_index_951103 == array_index_948679 ? add_951231 : sel_951228;
  assign add_951235 = sel_951232 + 8'h01;
  assign sel_951236 = array_index_951103 == array_index_948685 ? add_951235 : sel_951232;
  assign add_951239 = sel_951236 + 8'h01;
  assign sel_951240 = array_index_951103 == array_index_948691 ? add_951239 : sel_951236;
  assign add_951243 = sel_951240 + 8'h01;
  assign sel_951244 = array_index_951103 == array_index_948697 ? add_951243 : sel_951240;
  assign add_951247 = sel_951244 + 8'h01;
  assign sel_951248 = array_index_951103 == array_index_948703 ? add_951247 : sel_951244;
  assign add_951251 = sel_951248 + 8'h01;
  assign sel_951252 = array_index_951103 == array_index_948709 ? add_951251 : sel_951248;
  assign add_951255 = sel_951252 + 8'h01;
  assign sel_951256 = array_index_951103 == array_index_948715 ? add_951255 : sel_951252;
  assign add_951259 = sel_951256 + 8'h01;
  assign sel_951260 = array_index_951103 == array_index_948721 ? add_951259 : sel_951256;
  assign add_951263 = sel_951260 + 8'h01;
  assign sel_951264 = array_index_951103 == array_index_948727 ? add_951263 : sel_951260;
  assign add_951267 = sel_951264 + 8'h01;
  assign sel_951268 = array_index_951103 == array_index_948733 ? add_951267 : sel_951264;
  assign add_951271 = sel_951268 + 8'h01;
  assign sel_951272 = array_index_951103 == array_index_948739 ? add_951271 : sel_951268;
  assign add_951275 = sel_951272 + 8'h01;
  assign sel_951276 = array_index_951103 == array_index_948745 ? add_951275 : sel_951272;
  assign add_951279 = sel_951276 + 8'h01;
  assign sel_951280 = array_index_951103 == array_index_948751 ? add_951279 : sel_951276;
  assign add_951283 = sel_951280 + 8'h01;
  assign sel_951284 = array_index_951103 == array_index_948757 ? add_951283 : sel_951280;
  assign add_951287 = sel_951284 + 8'h01;
  assign sel_951288 = array_index_951103 == array_index_948763 ? add_951287 : sel_951284;
  assign add_951291 = sel_951288 + 8'h01;
  assign sel_951292 = array_index_951103 == array_index_948769 ? add_951291 : sel_951288;
  assign add_951295 = sel_951292 + 8'h01;
  assign sel_951296 = array_index_951103 == array_index_948775 ? add_951295 : sel_951292;
  assign add_951299 = sel_951296 + 8'h01;
  assign sel_951300 = array_index_951103 == array_index_948781 ? add_951299 : sel_951296;
  assign add_951303 = sel_951300 + 8'h01;
  assign sel_951304 = array_index_951103 == array_index_948787 ? add_951303 : sel_951300;
  assign add_951307 = sel_951304 + 8'h01;
  assign sel_951308 = array_index_951103 == array_index_948793 ? add_951307 : sel_951304;
  assign add_951311 = sel_951308 + 8'h01;
  assign sel_951312 = array_index_951103 == array_index_948799 ? add_951311 : sel_951308;
  assign add_951315 = sel_951312 + 8'h01;
  assign sel_951316 = array_index_951103 == array_index_948805 ? add_951315 : sel_951312;
  assign add_951319 = sel_951316 + 8'h01;
  assign sel_951320 = array_index_951103 == array_index_948811 ? add_951319 : sel_951316;
  assign add_951323 = sel_951320 + 8'h01;
  assign sel_951324 = array_index_951103 == array_index_948817 ? add_951323 : sel_951320;
  assign add_951327 = sel_951324 + 8'h01;
  assign sel_951328 = array_index_951103 == array_index_948823 ? add_951327 : sel_951324;
  assign add_951331 = sel_951328 + 8'h01;
  assign sel_951332 = array_index_951103 == array_index_948829 ? add_951331 : sel_951328;
  assign add_951335 = sel_951332 + 8'h01;
  assign sel_951336 = array_index_951103 == array_index_948835 ? add_951335 : sel_951332;
  assign add_951339 = sel_951336 + 8'h01;
  assign sel_951340 = array_index_951103 == array_index_948841 ? add_951339 : sel_951336;
  assign add_951343 = sel_951340 + 8'h01;
  assign sel_951344 = array_index_951103 == array_index_948847 ? add_951343 : sel_951340;
  assign add_951347 = sel_951344 + 8'h01;
  assign sel_951348 = array_index_951103 == array_index_948853 ? add_951347 : sel_951344;
  assign add_951351 = sel_951348 + 8'h01;
  assign sel_951352 = array_index_951103 == array_index_948859 ? add_951351 : sel_951348;
  assign add_951355 = sel_951352 + 8'h01;
  assign sel_951356 = array_index_951103 == array_index_948865 ? add_951355 : sel_951352;
  assign add_951359 = sel_951356 + 8'h01;
  assign sel_951360 = array_index_951103 == array_index_948871 ? add_951359 : sel_951356;
  assign add_951363 = sel_951360 + 8'h01;
  assign sel_951364 = array_index_951103 == array_index_948877 ? add_951363 : sel_951360;
  assign add_951367 = sel_951364 + 8'h01;
  assign sel_951368 = array_index_951103 == array_index_948883 ? add_951367 : sel_951364;
  assign add_951371 = sel_951368 + 8'h01;
  assign sel_951372 = array_index_951103 == array_index_948889 ? add_951371 : sel_951368;
  assign add_951375 = sel_951372 + 8'h01;
  assign sel_951376 = array_index_951103 == array_index_948895 ? add_951375 : sel_951372;
  assign add_951379 = sel_951376 + 8'h01;
  assign sel_951380 = array_index_951103 == array_index_948901 ? add_951379 : sel_951376;
  assign add_951383 = sel_951380 + 8'h01;
  assign sel_951384 = array_index_951103 == array_index_948907 ? add_951383 : sel_951380;
  assign add_951387 = sel_951384 + 8'h01;
  assign sel_951388 = array_index_951103 == array_index_948913 ? add_951387 : sel_951384;
  assign add_951391 = sel_951388 + 8'h01;
  assign sel_951392 = array_index_951103 == array_index_948919 ? add_951391 : sel_951388;
  assign add_951395 = sel_951392 + 8'h01;
  assign sel_951396 = array_index_951103 == array_index_948925 ? add_951395 : sel_951392;
  assign add_951399 = sel_951396 + 8'h01;
  assign sel_951400 = array_index_951103 == array_index_948931 ? add_951399 : sel_951396;
  assign add_951403 = sel_951400 + 8'h01;
  assign sel_951404 = array_index_951103 == array_index_948937 ? add_951403 : sel_951400;
  assign add_951407 = sel_951404 + 8'h01;
  assign sel_951408 = array_index_951103 == array_index_948943 ? add_951407 : sel_951404;
  assign add_951411 = sel_951408 + 8'h01;
  assign sel_951412 = array_index_951103 == array_index_948949 ? add_951411 : sel_951408;
  assign add_951415 = sel_951412 + 8'h01;
  assign sel_951416 = array_index_951103 == array_index_948955 ? add_951415 : sel_951412;
  assign add_951419 = sel_951416 + 8'h01;
  assign sel_951420 = array_index_951103 == array_index_948961 ? add_951419 : sel_951416;
  assign add_951423 = sel_951420 + 8'h01;
  assign sel_951424 = array_index_951103 == array_index_948967 ? add_951423 : sel_951420;
  assign add_951427 = sel_951424 + 8'h01;
  assign sel_951428 = array_index_951103 == array_index_948973 ? add_951427 : sel_951424;
  assign add_951431 = sel_951428 + 8'h01;
  assign sel_951432 = array_index_951103 == array_index_948979 ? add_951431 : sel_951428;
  assign add_951435 = sel_951432 + 8'h01;
  assign sel_951436 = array_index_951103 == array_index_948985 ? add_951435 : sel_951432;
  assign add_951439 = sel_951436 + 8'h01;
  assign sel_951440 = array_index_951103 == array_index_948991 ? add_951439 : sel_951436;
  assign add_951443 = sel_951440 + 8'h01;
  assign sel_951444 = array_index_951103 == array_index_948997 ? add_951443 : sel_951440;
  assign add_951447 = sel_951444 + 8'h01;
  assign sel_951448 = array_index_951103 == array_index_949003 ? add_951447 : sel_951444;
  assign add_951451 = sel_951448 + 8'h01;
  assign sel_951452 = array_index_951103 == array_index_949009 ? add_951451 : sel_951448;
  assign add_951455 = sel_951452 + 8'h01;
  assign sel_951456 = array_index_951103 == array_index_949015 ? add_951455 : sel_951452;
  assign add_951459 = sel_951456 + 8'h01;
  assign sel_951460 = array_index_951103 == array_index_949021 ? add_951459 : sel_951456;
  assign add_951463 = sel_951460 + 8'h01;
  assign sel_951464 = array_index_951103 == array_index_949027 ? add_951463 : sel_951460;
  assign add_951467 = sel_951464 + 8'h01;
  assign sel_951468 = array_index_951103 == array_index_949033 ? add_951467 : sel_951464;
  assign add_951471 = sel_951468 + 8'h01;
  assign sel_951472 = array_index_951103 == array_index_949039 ? add_951471 : sel_951468;
  assign add_951475 = sel_951472 + 8'h01;
  assign sel_951476 = array_index_951103 == array_index_949045 ? add_951475 : sel_951472;
  assign add_951479 = sel_951476 + 8'h01;
  assign sel_951480 = array_index_951103 == array_index_949051 ? add_951479 : sel_951476;
  assign add_951483 = sel_951480 + 8'h01;
  assign sel_951484 = array_index_951103 == array_index_949057 ? add_951483 : sel_951480;
  assign add_951487 = sel_951484 + 8'h01;
  assign sel_951488 = array_index_951103 == array_index_949063 ? add_951487 : sel_951484;
  assign add_951491 = sel_951488 + 8'h01;
  assign sel_951492 = array_index_951103 == array_index_949069 ? add_951491 : sel_951488;
  assign add_951495 = sel_951492 + 8'h01;
  assign sel_951496 = array_index_951103 == array_index_949075 ? add_951495 : sel_951492;
  assign add_951499 = sel_951496 + 8'h01;
  assign sel_951500 = array_index_951103 == array_index_949081 ? add_951499 : sel_951496;
  assign add_951504 = sel_951500 + 8'h01;
  assign array_index_951505 = set1_unflattened[7'h07];
  assign sel_951506 = array_index_951103 == array_index_949087 ? add_951504 : sel_951500;
  assign add_951509 = sel_951506 + 8'h01;
  assign sel_951510 = array_index_951505 == array_index_948483 ? add_951509 : sel_951506;
  assign add_951513 = sel_951510 + 8'h01;
  assign sel_951514 = array_index_951505 == array_index_948487 ? add_951513 : sel_951510;
  assign add_951517 = sel_951514 + 8'h01;
  assign sel_951518 = array_index_951505 == array_index_948495 ? add_951517 : sel_951514;
  assign add_951521 = sel_951518 + 8'h01;
  assign sel_951522 = array_index_951505 == array_index_948503 ? add_951521 : sel_951518;
  assign add_951525 = sel_951522 + 8'h01;
  assign sel_951526 = array_index_951505 == array_index_948511 ? add_951525 : sel_951522;
  assign add_951529 = sel_951526 + 8'h01;
  assign sel_951530 = array_index_951505 == array_index_948519 ? add_951529 : sel_951526;
  assign add_951533 = sel_951530 + 8'h01;
  assign sel_951534 = array_index_951505 == array_index_948527 ? add_951533 : sel_951530;
  assign add_951537 = sel_951534 + 8'h01;
  assign sel_951538 = array_index_951505 == array_index_948535 ? add_951537 : sel_951534;
  assign add_951541 = sel_951538 + 8'h01;
  assign sel_951542 = array_index_951505 == array_index_948541 ? add_951541 : sel_951538;
  assign add_951545 = sel_951542 + 8'h01;
  assign sel_951546 = array_index_951505 == array_index_948547 ? add_951545 : sel_951542;
  assign add_951549 = sel_951546 + 8'h01;
  assign sel_951550 = array_index_951505 == array_index_948553 ? add_951549 : sel_951546;
  assign add_951553 = sel_951550 + 8'h01;
  assign sel_951554 = array_index_951505 == array_index_948559 ? add_951553 : sel_951550;
  assign add_951557 = sel_951554 + 8'h01;
  assign sel_951558 = array_index_951505 == array_index_948565 ? add_951557 : sel_951554;
  assign add_951561 = sel_951558 + 8'h01;
  assign sel_951562 = array_index_951505 == array_index_948571 ? add_951561 : sel_951558;
  assign add_951565 = sel_951562 + 8'h01;
  assign sel_951566 = array_index_951505 == array_index_948577 ? add_951565 : sel_951562;
  assign add_951569 = sel_951566 + 8'h01;
  assign sel_951570 = array_index_951505 == array_index_948583 ? add_951569 : sel_951566;
  assign add_951573 = sel_951570 + 8'h01;
  assign sel_951574 = array_index_951505 == array_index_948589 ? add_951573 : sel_951570;
  assign add_951577 = sel_951574 + 8'h01;
  assign sel_951578 = array_index_951505 == array_index_948595 ? add_951577 : sel_951574;
  assign add_951581 = sel_951578 + 8'h01;
  assign sel_951582 = array_index_951505 == array_index_948601 ? add_951581 : sel_951578;
  assign add_951585 = sel_951582 + 8'h01;
  assign sel_951586 = array_index_951505 == array_index_948607 ? add_951585 : sel_951582;
  assign add_951589 = sel_951586 + 8'h01;
  assign sel_951590 = array_index_951505 == array_index_948613 ? add_951589 : sel_951586;
  assign add_951593 = sel_951590 + 8'h01;
  assign sel_951594 = array_index_951505 == array_index_948619 ? add_951593 : sel_951590;
  assign add_951597 = sel_951594 + 8'h01;
  assign sel_951598 = array_index_951505 == array_index_948625 ? add_951597 : sel_951594;
  assign add_951601 = sel_951598 + 8'h01;
  assign sel_951602 = array_index_951505 == array_index_948631 ? add_951601 : sel_951598;
  assign add_951605 = sel_951602 + 8'h01;
  assign sel_951606 = array_index_951505 == array_index_948637 ? add_951605 : sel_951602;
  assign add_951609 = sel_951606 + 8'h01;
  assign sel_951610 = array_index_951505 == array_index_948643 ? add_951609 : sel_951606;
  assign add_951613 = sel_951610 + 8'h01;
  assign sel_951614 = array_index_951505 == array_index_948649 ? add_951613 : sel_951610;
  assign add_951617 = sel_951614 + 8'h01;
  assign sel_951618 = array_index_951505 == array_index_948655 ? add_951617 : sel_951614;
  assign add_951621 = sel_951618 + 8'h01;
  assign sel_951622 = array_index_951505 == array_index_948661 ? add_951621 : sel_951618;
  assign add_951625 = sel_951622 + 8'h01;
  assign sel_951626 = array_index_951505 == array_index_948667 ? add_951625 : sel_951622;
  assign add_951629 = sel_951626 + 8'h01;
  assign sel_951630 = array_index_951505 == array_index_948673 ? add_951629 : sel_951626;
  assign add_951633 = sel_951630 + 8'h01;
  assign sel_951634 = array_index_951505 == array_index_948679 ? add_951633 : sel_951630;
  assign add_951637 = sel_951634 + 8'h01;
  assign sel_951638 = array_index_951505 == array_index_948685 ? add_951637 : sel_951634;
  assign add_951641 = sel_951638 + 8'h01;
  assign sel_951642 = array_index_951505 == array_index_948691 ? add_951641 : sel_951638;
  assign add_951645 = sel_951642 + 8'h01;
  assign sel_951646 = array_index_951505 == array_index_948697 ? add_951645 : sel_951642;
  assign add_951649 = sel_951646 + 8'h01;
  assign sel_951650 = array_index_951505 == array_index_948703 ? add_951649 : sel_951646;
  assign add_951653 = sel_951650 + 8'h01;
  assign sel_951654 = array_index_951505 == array_index_948709 ? add_951653 : sel_951650;
  assign add_951657 = sel_951654 + 8'h01;
  assign sel_951658 = array_index_951505 == array_index_948715 ? add_951657 : sel_951654;
  assign add_951661 = sel_951658 + 8'h01;
  assign sel_951662 = array_index_951505 == array_index_948721 ? add_951661 : sel_951658;
  assign add_951665 = sel_951662 + 8'h01;
  assign sel_951666 = array_index_951505 == array_index_948727 ? add_951665 : sel_951662;
  assign add_951669 = sel_951666 + 8'h01;
  assign sel_951670 = array_index_951505 == array_index_948733 ? add_951669 : sel_951666;
  assign add_951673 = sel_951670 + 8'h01;
  assign sel_951674 = array_index_951505 == array_index_948739 ? add_951673 : sel_951670;
  assign add_951677 = sel_951674 + 8'h01;
  assign sel_951678 = array_index_951505 == array_index_948745 ? add_951677 : sel_951674;
  assign add_951681 = sel_951678 + 8'h01;
  assign sel_951682 = array_index_951505 == array_index_948751 ? add_951681 : sel_951678;
  assign add_951685 = sel_951682 + 8'h01;
  assign sel_951686 = array_index_951505 == array_index_948757 ? add_951685 : sel_951682;
  assign add_951689 = sel_951686 + 8'h01;
  assign sel_951690 = array_index_951505 == array_index_948763 ? add_951689 : sel_951686;
  assign add_951693 = sel_951690 + 8'h01;
  assign sel_951694 = array_index_951505 == array_index_948769 ? add_951693 : sel_951690;
  assign add_951697 = sel_951694 + 8'h01;
  assign sel_951698 = array_index_951505 == array_index_948775 ? add_951697 : sel_951694;
  assign add_951701 = sel_951698 + 8'h01;
  assign sel_951702 = array_index_951505 == array_index_948781 ? add_951701 : sel_951698;
  assign add_951705 = sel_951702 + 8'h01;
  assign sel_951706 = array_index_951505 == array_index_948787 ? add_951705 : sel_951702;
  assign add_951709 = sel_951706 + 8'h01;
  assign sel_951710 = array_index_951505 == array_index_948793 ? add_951709 : sel_951706;
  assign add_951713 = sel_951710 + 8'h01;
  assign sel_951714 = array_index_951505 == array_index_948799 ? add_951713 : sel_951710;
  assign add_951717 = sel_951714 + 8'h01;
  assign sel_951718 = array_index_951505 == array_index_948805 ? add_951717 : sel_951714;
  assign add_951721 = sel_951718 + 8'h01;
  assign sel_951722 = array_index_951505 == array_index_948811 ? add_951721 : sel_951718;
  assign add_951725 = sel_951722 + 8'h01;
  assign sel_951726 = array_index_951505 == array_index_948817 ? add_951725 : sel_951722;
  assign add_951729 = sel_951726 + 8'h01;
  assign sel_951730 = array_index_951505 == array_index_948823 ? add_951729 : sel_951726;
  assign add_951733 = sel_951730 + 8'h01;
  assign sel_951734 = array_index_951505 == array_index_948829 ? add_951733 : sel_951730;
  assign add_951737 = sel_951734 + 8'h01;
  assign sel_951738 = array_index_951505 == array_index_948835 ? add_951737 : sel_951734;
  assign add_951741 = sel_951738 + 8'h01;
  assign sel_951742 = array_index_951505 == array_index_948841 ? add_951741 : sel_951738;
  assign add_951745 = sel_951742 + 8'h01;
  assign sel_951746 = array_index_951505 == array_index_948847 ? add_951745 : sel_951742;
  assign add_951749 = sel_951746 + 8'h01;
  assign sel_951750 = array_index_951505 == array_index_948853 ? add_951749 : sel_951746;
  assign add_951753 = sel_951750 + 8'h01;
  assign sel_951754 = array_index_951505 == array_index_948859 ? add_951753 : sel_951750;
  assign add_951757 = sel_951754 + 8'h01;
  assign sel_951758 = array_index_951505 == array_index_948865 ? add_951757 : sel_951754;
  assign add_951761 = sel_951758 + 8'h01;
  assign sel_951762 = array_index_951505 == array_index_948871 ? add_951761 : sel_951758;
  assign add_951765 = sel_951762 + 8'h01;
  assign sel_951766 = array_index_951505 == array_index_948877 ? add_951765 : sel_951762;
  assign add_951769 = sel_951766 + 8'h01;
  assign sel_951770 = array_index_951505 == array_index_948883 ? add_951769 : sel_951766;
  assign add_951773 = sel_951770 + 8'h01;
  assign sel_951774 = array_index_951505 == array_index_948889 ? add_951773 : sel_951770;
  assign add_951777 = sel_951774 + 8'h01;
  assign sel_951778 = array_index_951505 == array_index_948895 ? add_951777 : sel_951774;
  assign add_951781 = sel_951778 + 8'h01;
  assign sel_951782 = array_index_951505 == array_index_948901 ? add_951781 : sel_951778;
  assign add_951785 = sel_951782 + 8'h01;
  assign sel_951786 = array_index_951505 == array_index_948907 ? add_951785 : sel_951782;
  assign add_951789 = sel_951786 + 8'h01;
  assign sel_951790 = array_index_951505 == array_index_948913 ? add_951789 : sel_951786;
  assign add_951793 = sel_951790 + 8'h01;
  assign sel_951794 = array_index_951505 == array_index_948919 ? add_951793 : sel_951790;
  assign add_951797 = sel_951794 + 8'h01;
  assign sel_951798 = array_index_951505 == array_index_948925 ? add_951797 : sel_951794;
  assign add_951801 = sel_951798 + 8'h01;
  assign sel_951802 = array_index_951505 == array_index_948931 ? add_951801 : sel_951798;
  assign add_951805 = sel_951802 + 8'h01;
  assign sel_951806 = array_index_951505 == array_index_948937 ? add_951805 : sel_951802;
  assign add_951809 = sel_951806 + 8'h01;
  assign sel_951810 = array_index_951505 == array_index_948943 ? add_951809 : sel_951806;
  assign add_951813 = sel_951810 + 8'h01;
  assign sel_951814 = array_index_951505 == array_index_948949 ? add_951813 : sel_951810;
  assign add_951817 = sel_951814 + 8'h01;
  assign sel_951818 = array_index_951505 == array_index_948955 ? add_951817 : sel_951814;
  assign add_951821 = sel_951818 + 8'h01;
  assign sel_951822 = array_index_951505 == array_index_948961 ? add_951821 : sel_951818;
  assign add_951825 = sel_951822 + 8'h01;
  assign sel_951826 = array_index_951505 == array_index_948967 ? add_951825 : sel_951822;
  assign add_951829 = sel_951826 + 8'h01;
  assign sel_951830 = array_index_951505 == array_index_948973 ? add_951829 : sel_951826;
  assign add_951833 = sel_951830 + 8'h01;
  assign sel_951834 = array_index_951505 == array_index_948979 ? add_951833 : sel_951830;
  assign add_951837 = sel_951834 + 8'h01;
  assign sel_951838 = array_index_951505 == array_index_948985 ? add_951837 : sel_951834;
  assign add_951841 = sel_951838 + 8'h01;
  assign sel_951842 = array_index_951505 == array_index_948991 ? add_951841 : sel_951838;
  assign add_951845 = sel_951842 + 8'h01;
  assign sel_951846 = array_index_951505 == array_index_948997 ? add_951845 : sel_951842;
  assign add_951849 = sel_951846 + 8'h01;
  assign sel_951850 = array_index_951505 == array_index_949003 ? add_951849 : sel_951846;
  assign add_951853 = sel_951850 + 8'h01;
  assign sel_951854 = array_index_951505 == array_index_949009 ? add_951853 : sel_951850;
  assign add_951857 = sel_951854 + 8'h01;
  assign sel_951858 = array_index_951505 == array_index_949015 ? add_951857 : sel_951854;
  assign add_951861 = sel_951858 + 8'h01;
  assign sel_951862 = array_index_951505 == array_index_949021 ? add_951861 : sel_951858;
  assign add_951865 = sel_951862 + 8'h01;
  assign sel_951866 = array_index_951505 == array_index_949027 ? add_951865 : sel_951862;
  assign add_951869 = sel_951866 + 8'h01;
  assign sel_951870 = array_index_951505 == array_index_949033 ? add_951869 : sel_951866;
  assign add_951873 = sel_951870 + 8'h01;
  assign sel_951874 = array_index_951505 == array_index_949039 ? add_951873 : sel_951870;
  assign add_951877 = sel_951874 + 8'h01;
  assign sel_951878 = array_index_951505 == array_index_949045 ? add_951877 : sel_951874;
  assign add_951881 = sel_951878 + 8'h01;
  assign sel_951882 = array_index_951505 == array_index_949051 ? add_951881 : sel_951878;
  assign add_951885 = sel_951882 + 8'h01;
  assign sel_951886 = array_index_951505 == array_index_949057 ? add_951885 : sel_951882;
  assign add_951889 = sel_951886 + 8'h01;
  assign sel_951890 = array_index_951505 == array_index_949063 ? add_951889 : sel_951886;
  assign add_951893 = sel_951890 + 8'h01;
  assign sel_951894 = array_index_951505 == array_index_949069 ? add_951893 : sel_951890;
  assign add_951897 = sel_951894 + 8'h01;
  assign sel_951898 = array_index_951505 == array_index_949075 ? add_951897 : sel_951894;
  assign add_951901 = sel_951898 + 8'h01;
  assign sel_951902 = array_index_951505 == array_index_949081 ? add_951901 : sel_951898;
  assign add_951906 = sel_951902 + 8'h01;
  assign array_index_951907 = set1_unflattened[7'h08];
  assign sel_951908 = array_index_951505 == array_index_949087 ? add_951906 : sel_951902;
  assign add_951911 = sel_951908 + 8'h01;
  assign sel_951912 = array_index_951907 == array_index_948483 ? add_951911 : sel_951908;
  assign add_951915 = sel_951912 + 8'h01;
  assign sel_951916 = array_index_951907 == array_index_948487 ? add_951915 : sel_951912;
  assign add_951919 = sel_951916 + 8'h01;
  assign sel_951920 = array_index_951907 == array_index_948495 ? add_951919 : sel_951916;
  assign add_951923 = sel_951920 + 8'h01;
  assign sel_951924 = array_index_951907 == array_index_948503 ? add_951923 : sel_951920;
  assign add_951927 = sel_951924 + 8'h01;
  assign sel_951928 = array_index_951907 == array_index_948511 ? add_951927 : sel_951924;
  assign add_951931 = sel_951928 + 8'h01;
  assign sel_951932 = array_index_951907 == array_index_948519 ? add_951931 : sel_951928;
  assign add_951935 = sel_951932 + 8'h01;
  assign sel_951936 = array_index_951907 == array_index_948527 ? add_951935 : sel_951932;
  assign add_951939 = sel_951936 + 8'h01;
  assign sel_951940 = array_index_951907 == array_index_948535 ? add_951939 : sel_951936;
  assign add_951943 = sel_951940 + 8'h01;
  assign sel_951944 = array_index_951907 == array_index_948541 ? add_951943 : sel_951940;
  assign add_951947 = sel_951944 + 8'h01;
  assign sel_951948 = array_index_951907 == array_index_948547 ? add_951947 : sel_951944;
  assign add_951951 = sel_951948 + 8'h01;
  assign sel_951952 = array_index_951907 == array_index_948553 ? add_951951 : sel_951948;
  assign add_951955 = sel_951952 + 8'h01;
  assign sel_951956 = array_index_951907 == array_index_948559 ? add_951955 : sel_951952;
  assign add_951959 = sel_951956 + 8'h01;
  assign sel_951960 = array_index_951907 == array_index_948565 ? add_951959 : sel_951956;
  assign add_951963 = sel_951960 + 8'h01;
  assign sel_951964 = array_index_951907 == array_index_948571 ? add_951963 : sel_951960;
  assign add_951967 = sel_951964 + 8'h01;
  assign sel_951968 = array_index_951907 == array_index_948577 ? add_951967 : sel_951964;
  assign add_951971 = sel_951968 + 8'h01;
  assign sel_951972 = array_index_951907 == array_index_948583 ? add_951971 : sel_951968;
  assign add_951975 = sel_951972 + 8'h01;
  assign sel_951976 = array_index_951907 == array_index_948589 ? add_951975 : sel_951972;
  assign add_951979 = sel_951976 + 8'h01;
  assign sel_951980 = array_index_951907 == array_index_948595 ? add_951979 : sel_951976;
  assign add_951983 = sel_951980 + 8'h01;
  assign sel_951984 = array_index_951907 == array_index_948601 ? add_951983 : sel_951980;
  assign add_951987 = sel_951984 + 8'h01;
  assign sel_951988 = array_index_951907 == array_index_948607 ? add_951987 : sel_951984;
  assign add_951991 = sel_951988 + 8'h01;
  assign sel_951992 = array_index_951907 == array_index_948613 ? add_951991 : sel_951988;
  assign add_951995 = sel_951992 + 8'h01;
  assign sel_951996 = array_index_951907 == array_index_948619 ? add_951995 : sel_951992;
  assign add_951999 = sel_951996 + 8'h01;
  assign sel_952000 = array_index_951907 == array_index_948625 ? add_951999 : sel_951996;
  assign add_952003 = sel_952000 + 8'h01;
  assign sel_952004 = array_index_951907 == array_index_948631 ? add_952003 : sel_952000;
  assign add_952007 = sel_952004 + 8'h01;
  assign sel_952008 = array_index_951907 == array_index_948637 ? add_952007 : sel_952004;
  assign add_952011 = sel_952008 + 8'h01;
  assign sel_952012 = array_index_951907 == array_index_948643 ? add_952011 : sel_952008;
  assign add_952015 = sel_952012 + 8'h01;
  assign sel_952016 = array_index_951907 == array_index_948649 ? add_952015 : sel_952012;
  assign add_952019 = sel_952016 + 8'h01;
  assign sel_952020 = array_index_951907 == array_index_948655 ? add_952019 : sel_952016;
  assign add_952023 = sel_952020 + 8'h01;
  assign sel_952024 = array_index_951907 == array_index_948661 ? add_952023 : sel_952020;
  assign add_952027 = sel_952024 + 8'h01;
  assign sel_952028 = array_index_951907 == array_index_948667 ? add_952027 : sel_952024;
  assign add_952031 = sel_952028 + 8'h01;
  assign sel_952032 = array_index_951907 == array_index_948673 ? add_952031 : sel_952028;
  assign add_952035 = sel_952032 + 8'h01;
  assign sel_952036 = array_index_951907 == array_index_948679 ? add_952035 : sel_952032;
  assign add_952039 = sel_952036 + 8'h01;
  assign sel_952040 = array_index_951907 == array_index_948685 ? add_952039 : sel_952036;
  assign add_952043 = sel_952040 + 8'h01;
  assign sel_952044 = array_index_951907 == array_index_948691 ? add_952043 : sel_952040;
  assign add_952047 = sel_952044 + 8'h01;
  assign sel_952048 = array_index_951907 == array_index_948697 ? add_952047 : sel_952044;
  assign add_952051 = sel_952048 + 8'h01;
  assign sel_952052 = array_index_951907 == array_index_948703 ? add_952051 : sel_952048;
  assign add_952055 = sel_952052 + 8'h01;
  assign sel_952056 = array_index_951907 == array_index_948709 ? add_952055 : sel_952052;
  assign add_952059 = sel_952056 + 8'h01;
  assign sel_952060 = array_index_951907 == array_index_948715 ? add_952059 : sel_952056;
  assign add_952063 = sel_952060 + 8'h01;
  assign sel_952064 = array_index_951907 == array_index_948721 ? add_952063 : sel_952060;
  assign add_952067 = sel_952064 + 8'h01;
  assign sel_952068 = array_index_951907 == array_index_948727 ? add_952067 : sel_952064;
  assign add_952071 = sel_952068 + 8'h01;
  assign sel_952072 = array_index_951907 == array_index_948733 ? add_952071 : sel_952068;
  assign add_952075 = sel_952072 + 8'h01;
  assign sel_952076 = array_index_951907 == array_index_948739 ? add_952075 : sel_952072;
  assign add_952079 = sel_952076 + 8'h01;
  assign sel_952080 = array_index_951907 == array_index_948745 ? add_952079 : sel_952076;
  assign add_952083 = sel_952080 + 8'h01;
  assign sel_952084 = array_index_951907 == array_index_948751 ? add_952083 : sel_952080;
  assign add_952087 = sel_952084 + 8'h01;
  assign sel_952088 = array_index_951907 == array_index_948757 ? add_952087 : sel_952084;
  assign add_952091 = sel_952088 + 8'h01;
  assign sel_952092 = array_index_951907 == array_index_948763 ? add_952091 : sel_952088;
  assign add_952095 = sel_952092 + 8'h01;
  assign sel_952096 = array_index_951907 == array_index_948769 ? add_952095 : sel_952092;
  assign add_952099 = sel_952096 + 8'h01;
  assign sel_952100 = array_index_951907 == array_index_948775 ? add_952099 : sel_952096;
  assign add_952103 = sel_952100 + 8'h01;
  assign sel_952104 = array_index_951907 == array_index_948781 ? add_952103 : sel_952100;
  assign add_952107 = sel_952104 + 8'h01;
  assign sel_952108 = array_index_951907 == array_index_948787 ? add_952107 : sel_952104;
  assign add_952111 = sel_952108 + 8'h01;
  assign sel_952112 = array_index_951907 == array_index_948793 ? add_952111 : sel_952108;
  assign add_952115 = sel_952112 + 8'h01;
  assign sel_952116 = array_index_951907 == array_index_948799 ? add_952115 : sel_952112;
  assign add_952119 = sel_952116 + 8'h01;
  assign sel_952120 = array_index_951907 == array_index_948805 ? add_952119 : sel_952116;
  assign add_952123 = sel_952120 + 8'h01;
  assign sel_952124 = array_index_951907 == array_index_948811 ? add_952123 : sel_952120;
  assign add_952127 = sel_952124 + 8'h01;
  assign sel_952128 = array_index_951907 == array_index_948817 ? add_952127 : sel_952124;
  assign add_952131 = sel_952128 + 8'h01;
  assign sel_952132 = array_index_951907 == array_index_948823 ? add_952131 : sel_952128;
  assign add_952135 = sel_952132 + 8'h01;
  assign sel_952136 = array_index_951907 == array_index_948829 ? add_952135 : sel_952132;
  assign add_952139 = sel_952136 + 8'h01;
  assign sel_952140 = array_index_951907 == array_index_948835 ? add_952139 : sel_952136;
  assign add_952143 = sel_952140 + 8'h01;
  assign sel_952144 = array_index_951907 == array_index_948841 ? add_952143 : sel_952140;
  assign add_952147 = sel_952144 + 8'h01;
  assign sel_952148 = array_index_951907 == array_index_948847 ? add_952147 : sel_952144;
  assign add_952151 = sel_952148 + 8'h01;
  assign sel_952152 = array_index_951907 == array_index_948853 ? add_952151 : sel_952148;
  assign add_952155 = sel_952152 + 8'h01;
  assign sel_952156 = array_index_951907 == array_index_948859 ? add_952155 : sel_952152;
  assign add_952159 = sel_952156 + 8'h01;
  assign sel_952160 = array_index_951907 == array_index_948865 ? add_952159 : sel_952156;
  assign add_952163 = sel_952160 + 8'h01;
  assign sel_952164 = array_index_951907 == array_index_948871 ? add_952163 : sel_952160;
  assign add_952167 = sel_952164 + 8'h01;
  assign sel_952168 = array_index_951907 == array_index_948877 ? add_952167 : sel_952164;
  assign add_952171 = sel_952168 + 8'h01;
  assign sel_952172 = array_index_951907 == array_index_948883 ? add_952171 : sel_952168;
  assign add_952175 = sel_952172 + 8'h01;
  assign sel_952176 = array_index_951907 == array_index_948889 ? add_952175 : sel_952172;
  assign add_952179 = sel_952176 + 8'h01;
  assign sel_952180 = array_index_951907 == array_index_948895 ? add_952179 : sel_952176;
  assign add_952183 = sel_952180 + 8'h01;
  assign sel_952184 = array_index_951907 == array_index_948901 ? add_952183 : sel_952180;
  assign add_952187 = sel_952184 + 8'h01;
  assign sel_952188 = array_index_951907 == array_index_948907 ? add_952187 : sel_952184;
  assign add_952191 = sel_952188 + 8'h01;
  assign sel_952192 = array_index_951907 == array_index_948913 ? add_952191 : sel_952188;
  assign add_952195 = sel_952192 + 8'h01;
  assign sel_952196 = array_index_951907 == array_index_948919 ? add_952195 : sel_952192;
  assign add_952199 = sel_952196 + 8'h01;
  assign sel_952200 = array_index_951907 == array_index_948925 ? add_952199 : sel_952196;
  assign add_952203 = sel_952200 + 8'h01;
  assign sel_952204 = array_index_951907 == array_index_948931 ? add_952203 : sel_952200;
  assign add_952207 = sel_952204 + 8'h01;
  assign sel_952208 = array_index_951907 == array_index_948937 ? add_952207 : sel_952204;
  assign add_952211 = sel_952208 + 8'h01;
  assign sel_952212 = array_index_951907 == array_index_948943 ? add_952211 : sel_952208;
  assign add_952215 = sel_952212 + 8'h01;
  assign sel_952216 = array_index_951907 == array_index_948949 ? add_952215 : sel_952212;
  assign add_952219 = sel_952216 + 8'h01;
  assign sel_952220 = array_index_951907 == array_index_948955 ? add_952219 : sel_952216;
  assign add_952223 = sel_952220 + 8'h01;
  assign sel_952224 = array_index_951907 == array_index_948961 ? add_952223 : sel_952220;
  assign add_952227 = sel_952224 + 8'h01;
  assign sel_952228 = array_index_951907 == array_index_948967 ? add_952227 : sel_952224;
  assign add_952231 = sel_952228 + 8'h01;
  assign sel_952232 = array_index_951907 == array_index_948973 ? add_952231 : sel_952228;
  assign add_952235 = sel_952232 + 8'h01;
  assign sel_952236 = array_index_951907 == array_index_948979 ? add_952235 : sel_952232;
  assign add_952239 = sel_952236 + 8'h01;
  assign sel_952240 = array_index_951907 == array_index_948985 ? add_952239 : sel_952236;
  assign add_952243 = sel_952240 + 8'h01;
  assign sel_952244 = array_index_951907 == array_index_948991 ? add_952243 : sel_952240;
  assign add_952247 = sel_952244 + 8'h01;
  assign sel_952248 = array_index_951907 == array_index_948997 ? add_952247 : sel_952244;
  assign add_952251 = sel_952248 + 8'h01;
  assign sel_952252 = array_index_951907 == array_index_949003 ? add_952251 : sel_952248;
  assign add_952255 = sel_952252 + 8'h01;
  assign sel_952256 = array_index_951907 == array_index_949009 ? add_952255 : sel_952252;
  assign add_952259 = sel_952256 + 8'h01;
  assign sel_952260 = array_index_951907 == array_index_949015 ? add_952259 : sel_952256;
  assign add_952263 = sel_952260 + 8'h01;
  assign sel_952264 = array_index_951907 == array_index_949021 ? add_952263 : sel_952260;
  assign add_952267 = sel_952264 + 8'h01;
  assign sel_952268 = array_index_951907 == array_index_949027 ? add_952267 : sel_952264;
  assign add_952271 = sel_952268 + 8'h01;
  assign sel_952272 = array_index_951907 == array_index_949033 ? add_952271 : sel_952268;
  assign add_952275 = sel_952272 + 8'h01;
  assign sel_952276 = array_index_951907 == array_index_949039 ? add_952275 : sel_952272;
  assign add_952279 = sel_952276 + 8'h01;
  assign sel_952280 = array_index_951907 == array_index_949045 ? add_952279 : sel_952276;
  assign add_952283 = sel_952280 + 8'h01;
  assign sel_952284 = array_index_951907 == array_index_949051 ? add_952283 : sel_952280;
  assign add_952287 = sel_952284 + 8'h01;
  assign sel_952288 = array_index_951907 == array_index_949057 ? add_952287 : sel_952284;
  assign add_952291 = sel_952288 + 8'h01;
  assign sel_952292 = array_index_951907 == array_index_949063 ? add_952291 : sel_952288;
  assign add_952295 = sel_952292 + 8'h01;
  assign sel_952296 = array_index_951907 == array_index_949069 ? add_952295 : sel_952292;
  assign add_952299 = sel_952296 + 8'h01;
  assign sel_952300 = array_index_951907 == array_index_949075 ? add_952299 : sel_952296;
  assign add_952303 = sel_952300 + 8'h01;
  assign sel_952304 = array_index_951907 == array_index_949081 ? add_952303 : sel_952300;
  assign add_952308 = sel_952304 + 8'h01;
  assign array_index_952309 = set1_unflattened[7'h09];
  assign sel_952310 = array_index_951907 == array_index_949087 ? add_952308 : sel_952304;
  assign add_952313 = sel_952310 + 8'h01;
  assign sel_952314 = array_index_952309 == array_index_948483 ? add_952313 : sel_952310;
  assign add_952317 = sel_952314 + 8'h01;
  assign sel_952318 = array_index_952309 == array_index_948487 ? add_952317 : sel_952314;
  assign add_952321 = sel_952318 + 8'h01;
  assign sel_952322 = array_index_952309 == array_index_948495 ? add_952321 : sel_952318;
  assign add_952325 = sel_952322 + 8'h01;
  assign sel_952326 = array_index_952309 == array_index_948503 ? add_952325 : sel_952322;
  assign add_952329 = sel_952326 + 8'h01;
  assign sel_952330 = array_index_952309 == array_index_948511 ? add_952329 : sel_952326;
  assign add_952333 = sel_952330 + 8'h01;
  assign sel_952334 = array_index_952309 == array_index_948519 ? add_952333 : sel_952330;
  assign add_952337 = sel_952334 + 8'h01;
  assign sel_952338 = array_index_952309 == array_index_948527 ? add_952337 : sel_952334;
  assign add_952341 = sel_952338 + 8'h01;
  assign sel_952342 = array_index_952309 == array_index_948535 ? add_952341 : sel_952338;
  assign add_952345 = sel_952342 + 8'h01;
  assign sel_952346 = array_index_952309 == array_index_948541 ? add_952345 : sel_952342;
  assign add_952349 = sel_952346 + 8'h01;
  assign sel_952350 = array_index_952309 == array_index_948547 ? add_952349 : sel_952346;
  assign add_952353 = sel_952350 + 8'h01;
  assign sel_952354 = array_index_952309 == array_index_948553 ? add_952353 : sel_952350;
  assign add_952357 = sel_952354 + 8'h01;
  assign sel_952358 = array_index_952309 == array_index_948559 ? add_952357 : sel_952354;
  assign add_952361 = sel_952358 + 8'h01;
  assign sel_952362 = array_index_952309 == array_index_948565 ? add_952361 : sel_952358;
  assign add_952365 = sel_952362 + 8'h01;
  assign sel_952366 = array_index_952309 == array_index_948571 ? add_952365 : sel_952362;
  assign add_952369 = sel_952366 + 8'h01;
  assign sel_952370 = array_index_952309 == array_index_948577 ? add_952369 : sel_952366;
  assign add_952373 = sel_952370 + 8'h01;
  assign sel_952374 = array_index_952309 == array_index_948583 ? add_952373 : sel_952370;
  assign add_952377 = sel_952374 + 8'h01;
  assign sel_952378 = array_index_952309 == array_index_948589 ? add_952377 : sel_952374;
  assign add_952381 = sel_952378 + 8'h01;
  assign sel_952382 = array_index_952309 == array_index_948595 ? add_952381 : sel_952378;
  assign add_952385 = sel_952382 + 8'h01;
  assign sel_952386 = array_index_952309 == array_index_948601 ? add_952385 : sel_952382;
  assign add_952389 = sel_952386 + 8'h01;
  assign sel_952390 = array_index_952309 == array_index_948607 ? add_952389 : sel_952386;
  assign add_952393 = sel_952390 + 8'h01;
  assign sel_952394 = array_index_952309 == array_index_948613 ? add_952393 : sel_952390;
  assign add_952397 = sel_952394 + 8'h01;
  assign sel_952398 = array_index_952309 == array_index_948619 ? add_952397 : sel_952394;
  assign add_952401 = sel_952398 + 8'h01;
  assign sel_952402 = array_index_952309 == array_index_948625 ? add_952401 : sel_952398;
  assign add_952405 = sel_952402 + 8'h01;
  assign sel_952406 = array_index_952309 == array_index_948631 ? add_952405 : sel_952402;
  assign add_952409 = sel_952406 + 8'h01;
  assign sel_952410 = array_index_952309 == array_index_948637 ? add_952409 : sel_952406;
  assign add_952413 = sel_952410 + 8'h01;
  assign sel_952414 = array_index_952309 == array_index_948643 ? add_952413 : sel_952410;
  assign add_952417 = sel_952414 + 8'h01;
  assign sel_952418 = array_index_952309 == array_index_948649 ? add_952417 : sel_952414;
  assign add_952421 = sel_952418 + 8'h01;
  assign sel_952422 = array_index_952309 == array_index_948655 ? add_952421 : sel_952418;
  assign add_952425 = sel_952422 + 8'h01;
  assign sel_952426 = array_index_952309 == array_index_948661 ? add_952425 : sel_952422;
  assign add_952429 = sel_952426 + 8'h01;
  assign sel_952430 = array_index_952309 == array_index_948667 ? add_952429 : sel_952426;
  assign add_952433 = sel_952430 + 8'h01;
  assign sel_952434 = array_index_952309 == array_index_948673 ? add_952433 : sel_952430;
  assign add_952437 = sel_952434 + 8'h01;
  assign sel_952438 = array_index_952309 == array_index_948679 ? add_952437 : sel_952434;
  assign add_952441 = sel_952438 + 8'h01;
  assign sel_952442 = array_index_952309 == array_index_948685 ? add_952441 : sel_952438;
  assign add_952445 = sel_952442 + 8'h01;
  assign sel_952446 = array_index_952309 == array_index_948691 ? add_952445 : sel_952442;
  assign add_952449 = sel_952446 + 8'h01;
  assign sel_952450 = array_index_952309 == array_index_948697 ? add_952449 : sel_952446;
  assign add_952453 = sel_952450 + 8'h01;
  assign sel_952454 = array_index_952309 == array_index_948703 ? add_952453 : sel_952450;
  assign add_952457 = sel_952454 + 8'h01;
  assign sel_952458 = array_index_952309 == array_index_948709 ? add_952457 : sel_952454;
  assign add_952461 = sel_952458 + 8'h01;
  assign sel_952462 = array_index_952309 == array_index_948715 ? add_952461 : sel_952458;
  assign add_952465 = sel_952462 + 8'h01;
  assign sel_952466 = array_index_952309 == array_index_948721 ? add_952465 : sel_952462;
  assign add_952469 = sel_952466 + 8'h01;
  assign sel_952470 = array_index_952309 == array_index_948727 ? add_952469 : sel_952466;
  assign add_952473 = sel_952470 + 8'h01;
  assign sel_952474 = array_index_952309 == array_index_948733 ? add_952473 : sel_952470;
  assign add_952477 = sel_952474 + 8'h01;
  assign sel_952478 = array_index_952309 == array_index_948739 ? add_952477 : sel_952474;
  assign add_952481 = sel_952478 + 8'h01;
  assign sel_952482 = array_index_952309 == array_index_948745 ? add_952481 : sel_952478;
  assign add_952485 = sel_952482 + 8'h01;
  assign sel_952486 = array_index_952309 == array_index_948751 ? add_952485 : sel_952482;
  assign add_952489 = sel_952486 + 8'h01;
  assign sel_952490 = array_index_952309 == array_index_948757 ? add_952489 : sel_952486;
  assign add_952493 = sel_952490 + 8'h01;
  assign sel_952494 = array_index_952309 == array_index_948763 ? add_952493 : sel_952490;
  assign add_952497 = sel_952494 + 8'h01;
  assign sel_952498 = array_index_952309 == array_index_948769 ? add_952497 : sel_952494;
  assign add_952501 = sel_952498 + 8'h01;
  assign sel_952502 = array_index_952309 == array_index_948775 ? add_952501 : sel_952498;
  assign add_952505 = sel_952502 + 8'h01;
  assign sel_952506 = array_index_952309 == array_index_948781 ? add_952505 : sel_952502;
  assign add_952509 = sel_952506 + 8'h01;
  assign sel_952510 = array_index_952309 == array_index_948787 ? add_952509 : sel_952506;
  assign add_952513 = sel_952510 + 8'h01;
  assign sel_952514 = array_index_952309 == array_index_948793 ? add_952513 : sel_952510;
  assign add_952517 = sel_952514 + 8'h01;
  assign sel_952518 = array_index_952309 == array_index_948799 ? add_952517 : sel_952514;
  assign add_952521 = sel_952518 + 8'h01;
  assign sel_952522 = array_index_952309 == array_index_948805 ? add_952521 : sel_952518;
  assign add_952525 = sel_952522 + 8'h01;
  assign sel_952526 = array_index_952309 == array_index_948811 ? add_952525 : sel_952522;
  assign add_952529 = sel_952526 + 8'h01;
  assign sel_952530 = array_index_952309 == array_index_948817 ? add_952529 : sel_952526;
  assign add_952533 = sel_952530 + 8'h01;
  assign sel_952534 = array_index_952309 == array_index_948823 ? add_952533 : sel_952530;
  assign add_952537 = sel_952534 + 8'h01;
  assign sel_952538 = array_index_952309 == array_index_948829 ? add_952537 : sel_952534;
  assign add_952541 = sel_952538 + 8'h01;
  assign sel_952542 = array_index_952309 == array_index_948835 ? add_952541 : sel_952538;
  assign add_952545 = sel_952542 + 8'h01;
  assign sel_952546 = array_index_952309 == array_index_948841 ? add_952545 : sel_952542;
  assign add_952549 = sel_952546 + 8'h01;
  assign sel_952550 = array_index_952309 == array_index_948847 ? add_952549 : sel_952546;
  assign add_952553 = sel_952550 + 8'h01;
  assign sel_952554 = array_index_952309 == array_index_948853 ? add_952553 : sel_952550;
  assign add_952557 = sel_952554 + 8'h01;
  assign sel_952558 = array_index_952309 == array_index_948859 ? add_952557 : sel_952554;
  assign add_952561 = sel_952558 + 8'h01;
  assign sel_952562 = array_index_952309 == array_index_948865 ? add_952561 : sel_952558;
  assign add_952565 = sel_952562 + 8'h01;
  assign sel_952566 = array_index_952309 == array_index_948871 ? add_952565 : sel_952562;
  assign add_952569 = sel_952566 + 8'h01;
  assign sel_952570 = array_index_952309 == array_index_948877 ? add_952569 : sel_952566;
  assign add_952573 = sel_952570 + 8'h01;
  assign sel_952574 = array_index_952309 == array_index_948883 ? add_952573 : sel_952570;
  assign add_952577 = sel_952574 + 8'h01;
  assign sel_952578 = array_index_952309 == array_index_948889 ? add_952577 : sel_952574;
  assign add_952581 = sel_952578 + 8'h01;
  assign sel_952582 = array_index_952309 == array_index_948895 ? add_952581 : sel_952578;
  assign add_952585 = sel_952582 + 8'h01;
  assign sel_952586 = array_index_952309 == array_index_948901 ? add_952585 : sel_952582;
  assign add_952589 = sel_952586 + 8'h01;
  assign sel_952590 = array_index_952309 == array_index_948907 ? add_952589 : sel_952586;
  assign add_952593 = sel_952590 + 8'h01;
  assign sel_952594 = array_index_952309 == array_index_948913 ? add_952593 : sel_952590;
  assign add_952597 = sel_952594 + 8'h01;
  assign sel_952598 = array_index_952309 == array_index_948919 ? add_952597 : sel_952594;
  assign add_952601 = sel_952598 + 8'h01;
  assign sel_952602 = array_index_952309 == array_index_948925 ? add_952601 : sel_952598;
  assign add_952605 = sel_952602 + 8'h01;
  assign sel_952606 = array_index_952309 == array_index_948931 ? add_952605 : sel_952602;
  assign add_952609 = sel_952606 + 8'h01;
  assign sel_952610 = array_index_952309 == array_index_948937 ? add_952609 : sel_952606;
  assign add_952613 = sel_952610 + 8'h01;
  assign sel_952614 = array_index_952309 == array_index_948943 ? add_952613 : sel_952610;
  assign add_952617 = sel_952614 + 8'h01;
  assign sel_952618 = array_index_952309 == array_index_948949 ? add_952617 : sel_952614;
  assign add_952621 = sel_952618 + 8'h01;
  assign sel_952622 = array_index_952309 == array_index_948955 ? add_952621 : sel_952618;
  assign add_952625 = sel_952622 + 8'h01;
  assign sel_952626 = array_index_952309 == array_index_948961 ? add_952625 : sel_952622;
  assign add_952629 = sel_952626 + 8'h01;
  assign sel_952630 = array_index_952309 == array_index_948967 ? add_952629 : sel_952626;
  assign add_952633 = sel_952630 + 8'h01;
  assign sel_952634 = array_index_952309 == array_index_948973 ? add_952633 : sel_952630;
  assign add_952637 = sel_952634 + 8'h01;
  assign sel_952638 = array_index_952309 == array_index_948979 ? add_952637 : sel_952634;
  assign add_952641 = sel_952638 + 8'h01;
  assign sel_952642 = array_index_952309 == array_index_948985 ? add_952641 : sel_952638;
  assign add_952645 = sel_952642 + 8'h01;
  assign sel_952646 = array_index_952309 == array_index_948991 ? add_952645 : sel_952642;
  assign add_952649 = sel_952646 + 8'h01;
  assign sel_952650 = array_index_952309 == array_index_948997 ? add_952649 : sel_952646;
  assign add_952653 = sel_952650 + 8'h01;
  assign sel_952654 = array_index_952309 == array_index_949003 ? add_952653 : sel_952650;
  assign add_952657 = sel_952654 + 8'h01;
  assign sel_952658 = array_index_952309 == array_index_949009 ? add_952657 : sel_952654;
  assign add_952661 = sel_952658 + 8'h01;
  assign sel_952662 = array_index_952309 == array_index_949015 ? add_952661 : sel_952658;
  assign add_952665 = sel_952662 + 8'h01;
  assign sel_952666 = array_index_952309 == array_index_949021 ? add_952665 : sel_952662;
  assign add_952669 = sel_952666 + 8'h01;
  assign sel_952670 = array_index_952309 == array_index_949027 ? add_952669 : sel_952666;
  assign add_952673 = sel_952670 + 8'h01;
  assign sel_952674 = array_index_952309 == array_index_949033 ? add_952673 : sel_952670;
  assign add_952677 = sel_952674 + 8'h01;
  assign sel_952678 = array_index_952309 == array_index_949039 ? add_952677 : sel_952674;
  assign add_952681 = sel_952678 + 8'h01;
  assign sel_952682 = array_index_952309 == array_index_949045 ? add_952681 : sel_952678;
  assign add_952685 = sel_952682 + 8'h01;
  assign sel_952686 = array_index_952309 == array_index_949051 ? add_952685 : sel_952682;
  assign add_952689 = sel_952686 + 8'h01;
  assign sel_952690 = array_index_952309 == array_index_949057 ? add_952689 : sel_952686;
  assign add_952693 = sel_952690 + 8'h01;
  assign sel_952694 = array_index_952309 == array_index_949063 ? add_952693 : sel_952690;
  assign add_952697 = sel_952694 + 8'h01;
  assign sel_952698 = array_index_952309 == array_index_949069 ? add_952697 : sel_952694;
  assign add_952701 = sel_952698 + 8'h01;
  assign sel_952702 = array_index_952309 == array_index_949075 ? add_952701 : sel_952698;
  assign add_952705 = sel_952702 + 8'h01;
  assign sel_952706 = array_index_952309 == array_index_949081 ? add_952705 : sel_952702;
  assign add_952710 = sel_952706 + 8'h01;
  assign array_index_952711 = set1_unflattened[7'h0a];
  assign sel_952712 = array_index_952309 == array_index_949087 ? add_952710 : sel_952706;
  assign add_952715 = sel_952712 + 8'h01;
  assign sel_952716 = array_index_952711 == array_index_948483 ? add_952715 : sel_952712;
  assign add_952719 = sel_952716 + 8'h01;
  assign sel_952720 = array_index_952711 == array_index_948487 ? add_952719 : sel_952716;
  assign add_952723 = sel_952720 + 8'h01;
  assign sel_952724 = array_index_952711 == array_index_948495 ? add_952723 : sel_952720;
  assign add_952727 = sel_952724 + 8'h01;
  assign sel_952728 = array_index_952711 == array_index_948503 ? add_952727 : sel_952724;
  assign add_952731 = sel_952728 + 8'h01;
  assign sel_952732 = array_index_952711 == array_index_948511 ? add_952731 : sel_952728;
  assign add_952735 = sel_952732 + 8'h01;
  assign sel_952736 = array_index_952711 == array_index_948519 ? add_952735 : sel_952732;
  assign add_952739 = sel_952736 + 8'h01;
  assign sel_952740 = array_index_952711 == array_index_948527 ? add_952739 : sel_952736;
  assign add_952743 = sel_952740 + 8'h01;
  assign sel_952744 = array_index_952711 == array_index_948535 ? add_952743 : sel_952740;
  assign add_952747 = sel_952744 + 8'h01;
  assign sel_952748 = array_index_952711 == array_index_948541 ? add_952747 : sel_952744;
  assign add_952751 = sel_952748 + 8'h01;
  assign sel_952752 = array_index_952711 == array_index_948547 ? add_952751 : sel_952748;
  assign add_952755 = sel_952752 + 8'h01;
  assign sel_952756 = array_index_952711 == array_index_948553 ? add_952755 : sel_952752;
  assign add_952759 = sel_952756 + 8'h01;
  assign sel_952760 = array_index_952711 == array_index_948559 ? add_952759 : sel_952756;
  assign add_952763 = sel_952760 + 8'h01;
  assign sel_952764 = array_index_952711 == array_index_948565 ? add_952763 : sel_952760;
  assign add_952767 = sel_952764 + 8'h01;
  assign sel_952768 = array_index_952711 == array_index_948571 ? add_952767 : sel_952764;
  assign add_952771 = sel_952768 + 8'h01;
  assign sel_952772 = array_index_952711 == array_index_948577 ? add_952771 : sel_952768;
  assign add_952775 = sel_952772 + 8'h01;
  assign sel_952776 = array_index_952711 == array_index_948583 ? add_952775 : sel_952772;
  assign add_952779 = sel_952776 + 8'h01;
  assign sel_952780 = array_index_952711 == array_index_948589 ? add_952779 : sel_952776;
  assign add_952783 = sel_952780 + 8'h01;
  assign sel_952784 = array_index_952711 == array_index_948595 ? add_952783 : sel_952780;
  assign add_952787 = sel_952784 + 8'h01;
  assign sel_952788 = array_index_952711 == array_index_948601 ? add_952787 : sel_952784;
  assign add_952791 = sel_952788 + 8'h01;
  assign sel_952792 = array_index_952711 == array_index_948607 ? add_952791 : sel_952788;
  assign add_952795 = sel_952792 + 8'h01;
  assign sel_952796 = array_index_952711 == array_index_948613 ? add_952795 : sel_952792;
  assign add_952799 = sel_952796 + 8'h01;
  assign sel_952800 = array_index_952711 == array_index_948619 ? add_952799 : sel_952796;
  assign add_952803 = sel_952800 + 8'h01;
  assign sel_952804 = array_index_952711 == array_index_948625 ? add_952803 : sel_952800;
  assign add_952807 = sel_952804 + 8'h01;
  assign sel_952808 = array_index_952711 == array_index_948631 ? add_952807 : sel_952804;
  assign add_952811 = sel_952808 + 8'h01;
  assign sel_952812 = array_index_952711 == array_index_948637 ? add_952811 : sel_952808;
  assign add_952815 = sel_952812 + 8'h01;
  assign sel_952816 = array_index_952711 == array_index_948643 ? add_952815 : sel_952812;
  assign add_952819 = sel_952816 + 8'h01;
  assign sel_952820 = array_index_952711 == array_index_948649 ? add_952819 : sel_952816;
  assign add_952823 = sel_952820 + 8'h01;
  assign sel_952824 = array_index_952711 == array_index_948655 ? add_952823 : sel_952820;
  assign add_952827 = sel_952824 + 8'h01;
  assign sel_952828 = array_index_952711 == array_index_948661 ? add_952827 : sel_952824;
  assign add_952831 = sel_952828 + 8'h01;
  assign sel_952832 = array_index_952711 == array_index_948667 ? add_952831 : sel_952828;
  assign add_952835 = sel_952832 + 8'h01;
  assign sel_952836 = array_index_952711 == array_index_948673 ? add_952835 : sel_952832;
  assign add_952839 = sel_952836 + 8'h01;
  assign sel_952840 = array_index_952711 == array_index_948679 ? add_952839 : sel_952836;
  assign add_952843 = sel_952840 + 8'h01;
  assign sel_952844 = array_index_952711 == array_index_948685 ? add_952843 : sel_952840;
  assign add_952847 = sel_952844 + 8'h01;
  assign sel_952848 = array_index_952711 == array_index_948691 ? add_952847 : sel_952844;
  assign add_952851 = sel_952848 + 8'h01;
  assign sel_952852 = array_index_952711 == array_index_948697 ? add_952851 : sel_952848;
  assign add_952855 = sel_952852 + 8'h01;
  assign sel_952856 = array_index_952711 == array_index_948703 ? add_952855 : sel_952852;
  assign add_952859 = sel_952856 + 8'h01;
  assign sel_952860 = array_index_952711 == array_index_948709 ? add_952859 : sel_952856;
  assign add_952863 = sel_952860 + 8'h01;
  assign sel_952864 = array_index_952711 == array_index_948715 ? add_952863 : sel_952860;
  assign add_952867 = sel_952864 + 8'h01;
  assign sel_952868 = array_index_952711 == array_index_948721 ? add_952867 : sel_952864;
  assign add_952871 = sel_952868 + 8'h01;
  assign sel_952872 = array_index_952711 == array_index_948727 ? add_952871 : sel_952868;
  assign add_952875 = sel_952872 + 8'h01;
  assign sel_952876 = array_index_952711 == array_index_948733 ? add_952875 : sel_952872;
  assign add_952879 = sel_952876 + 8'h01;
  assign sel_952880 = array_index_952711 == array_index_948739 ? add_952879 : sel_952876;
  assign add_952883 = sel_952880 + 8'h01;
  assign sel_952884 = array_index_952711 == array_index_948745 ? add_952883 : sel_952880;
  assign add_952887 = sel_952884 + 8'h01;
  assign sel_952888 = array_index_952711 == array_index_948751 ? add_952887 : sel_952884;
  assign add_952891 = sel_952888 + 8'h01;
  assign sel_952892 = array_index_952711 == array_index_948757 ? add_952891 : sel_952888;
  assign add_952895 = sel_952892 + 8'h01;
  assign sel_952896 = array_index_952711 == array_index_948763 ? add_952895 : sel_952892;
  assign add_952899 = sel_952896 + 8'h01;
  assign sel_952900 = array_index_952711 == array_index_948769 ? add_952899 : sel_952896;
  assign add_952903 = sel_952900 + 8'h01;
  assign sel_952904 = array_index_952711 == array_index_948775 ? add_952903 : sel_952900;
  assign add_952907 = sel_952904 + 8'h01;
  assign sel_952908 = array_index_952711 == array_index_948781 ? add_952907 : sel_952904;
  assign add_952911 = sel_952908 + 8'h01;
  assign sel_952912 = array_index_952711 == array_index_948787 ? add_952911 : sel_952908;
  assign add_952915 = sel_952912 + 8'h01;
  assign sel_952916 = array_index_952711 == array_index_948793 ? add_952915 : sel_952912;
  assign add_952919 = sel_952916 + 8'h01;
  assign sel_952920 = array_index_952711 == array_index_948799 ? add_952919 : sel_952916;
  assign add_952923 = sel_952920 + 8'h01;
  assign sel_952924 = array_index_952711 == array_index_948805 ? add_952923 : sel_952920;
  assign add_952927 = sel_952924 + 8'h01;
  assign sel_952928 = array_index_952711 == array_index_948811 ? add_952927 : sel_952924;
  assign add_952931 = sel_952928 + 8'h01;
  assign sel_952932 = array_index_952711 == array_index_948817 ? add_952931 : sel_952928;
  assign add_952935 = sel_952932 + 8'h01;
  assign sel_952936 = array_index_952711 == array_index_948823 ? add_952935 : sel_952932;
  assign add_952939 = sel_952936 + 8'h01;
  assign sel_952940 = array_index_952711 == array_index_948829 ? add_952939 : sel_952936;
  assign add_952943 = sel_952940 + 8'h01;
  assign sel_952944 = array_index_952711 == array_index_948835 ? add_952943 : sel_952940;
  assign add_952947 = sel_952944 + 8'h01;
  assign sel_952948 = array_index_952711 == array_index_948841 ? add_952947 : sel_952944;
  assign add_952951 = sel_952948 + 8'h01;
  assign sel_952952 = array_index_952711 == array_index_948847 ? add_952951 : sel_952948;
  assign add_952955 = sel_952952 + 8'h01;
  assign sel_952956 = array_index_952711 == array_index_948853 ? add_952955 : sel_952952;
  assign add_952959 = sel_952956 + 8'h01;
  assign sel_952960 = array_index_952711 == array_index_948859 ? add_952959 : sel_952956;
  assign add_952963 = sel_952960 + 8'h01;
  assign sel_952964 = array_index_952711 == array_index_948865 ? add_952963 : sel_952960;
  assign add_952967 = sel_952964 + 8'h01;
  assign sel_952968 = array_index_952711 == array_index_948871 ? add_952967 : sel_952964;
  assign add_952971 = sel_952968 + 8'h01;
  assign sel_952972 = array_index_952711 == array_index_948877 ? add_952971 : sel_952968;
  assign add_952975 = sel_952972 + 8'h01;
  assign sel_952976 = array_index_952711 == array_index_948883 ? add_952975 : sel_952972;
  assign add_952979 = sel_952976 + 8'h01;
  assign sel_952980 = array_index_952711 == array_index_948889 ? add_952979 : sel_952976;
  assign add_952983 = sel_952980 + 8'h01;
  assign sel_952984 = array_index_952711 == array_index_948895 ? add_952983 : sel_952980;
  assign add_952987 = sel_952984 + 8'h01;
  assign sel_952988 = array_index_952711 == array_index_948901 ? add_952987 : sel_952984;
  assign add_952991 = sel_952988 + 8'h01;
  assign sel_952992 = array_index_952711 == array_index_948907 ? add_952991 : sel_952988;
  assign add_952995 = sel_952992 + 8'h01;
  assign sel_952996 = array_index_952711 == array_index_948913 ? add_952995 : sel_952992;
  assign add_952999 = sel_952996 + 8'h01;
  assign sel_953000 = array_index_952711 == array_index_948919 ? add_952999 : sel_952996;
  assign add_953003 = sel_953000 + 8'h01;
  assign sel_953004 = array_index_952711 == array_index_948925 ? add_953003 : sel_953000;
  assign add_953007 = sel_953004 + 8'h01;
  assign sel_953008 = array_index_952711 == array_index_948931 ? add_953007 : sel_953004;
  assign add_953011 = sel_953008 + 8'h01;
  assign sel_953012 = array_index_952711 == array_index_948937 ? add_953011 : sel_953008;
  assign add_953015 = sel_953012 + 8'h01;
  assign sel_953016 = array_index_952711 == array_index_948943 ? add_953015 : sel_953012;
  assign add_953019 = sel_953016 + 8'h01;
  assign sel_953020 = array_index_952711 == array_index_948949 ? add_953019 : sel_953016;
  assign add_953023 = sel_953020 + 8'h01;
  assign sel_953024 = array_index_952711 == array_index_948955 ? add_953023 : sel_953020;
  assign add_953027 = sel_953024 + 8'h01;
  assign sel_953028 = array_index_952711 == array_index_948961 ? add_953027 : sel_953024;
  assign add_953031 = sel_953028 + 8'h01;
  assign sel_953032 = array_index_952711 == array_index_948967 ? add_953031 : sel_953028;
  assign add_953035 = sel_953032 + 8'h01;
  assign sel_953036 = array_index_952711 == array_index_948973 ? add_953035 : sel_953032;
  assign add_953039 = sel_953036 + 8'h01;
  assign sel_953040 = array_index_952711 == array_index_948979 ? add_953039 : sel_953036;
  assign add_953043 = sel_953040 + 8'h01;
  assign sel_953044 = array_index_952711 == array_index_948985 ? add_953043 : sel_953040;
  assign add_953047 = sel_953044 + 8'h01;
  assign sel_953048 = array_index_952711 == array_index_948991 ? add_953047 : sel_953044;
  assign add_953051 = sel_953048 + 8'h01;
  assign sel_953052 = array_index_952711 == array_index_948997 ? add_953051 : sel_953048;
  assign add_953055 = sel_953052 + 8'h01;
  assign sel_953056 = array_index_952711 == array_index_949003 ? add_953055 : sel_953052;
  assign add_953059 = sel_953056 + 8'h01;
  assign sel_953060 = array_index_952711 == array_index_949009 ? add_953059 : sel_953056;
  assign add_953063 = sel_953060 + 8'h01;
  assign sel_953064 = array_index_952711 == array_index_949015 ? add_953063 : sel_953060;
  assign add_953067 = sel_953064 + 8'h01;
  assign sel_953068 = array_index_952711 == array_index_949021 ? add_953067 : sel_953064;
  assign add_953071 = sel_953068 + 8'h01;
  assign sel_953072 = array_index_952711 == array_index_949027 ? add_953071 : sel_953068;
  assign add_953075 = sel_953072 + 8'h01;
  assign sel_953076 = array_index_952711 == array_index_949033 ? add_953075 : sel_953072;
  assign add_953079 = sel_953076 + 8'h01;
  assign sel_953080 = array_index_952711 == array_index_949039 ? add_953079 : sel_953076;
  assign add_953083 = sel_953080 + 8'h01;
  assign sel_953084 = array_index_952711 == array_index_949045 ? add_953083 : sel_953080;
  assign add_953087 = sel_953084 + 8'h01;
  assign sel_953088 = array_index_952711 == array_index_949051 ? add_953087 : sel_953084;
  assign add_953091 = sel_953088 + 8'h01;
  assign sel_953092 = array_index_952711 == array_index_949057 ? add_953091 : sel_953088;
  assign add_953095 = sel_953092 + 8'h01;
  assign sel_953096 = array_index_952711 == array_index_949063 ? add_953095 : sel_953092;
  assign add_953099 = sel_953096 + 8'h01;
  assign sel_953100 = array_index_952711 == array_index_949069 ? add_953099 : sel_953096;
  assign add_953103 = sel_953100 + 8'h01;
  assign sel_953104 = array_index_952711 == array_index_949075 ? add_953103 : sel_953100;
  assign add_953107 = sel_953104 + 8'h01;
  assign sel_953108 = array_index_952711 == array_index_949081 ? add_953107 : sel_953104;
  assign add_953112 = sel_953108 + 8'h01;
  assign array_index_953113 = set1_unflattened[7'h0b];
  assign sel_953114 = array_index_952711 == array_index_949087 ? add_953112 : sel_953108;
  assign add_953117 = sel_953114 + 8'h01;
  assign sel_953118 = array_index_953113 == array_index_948483 ? add_953117 : sel_953114;
  assign add_953121 = sel_953118 + 8'h01;
  assign sel_953122 = array_index_953113 == array_index_948487 ? add_953121 : sel_953118;
  assign add_953125 = sel_953122 + 8'h01;
  assign sel_953126 = array_index_953113 == array_index_948495 ? add_953125 : sel_953122;
  assign add_953129 = sel_953126 + 8'h01;
  assign sel_953130 = array_index_953113 == array_index_948503 ? add_953129 : sel_953126;
  assign add_953133 = sel_953130 + 8'h01;
  assign sel_953134 = array_index_953113 == array_index_948511 ? add_953133 : sel_953130;
  assign add_953137 = sel_953134 + 8'h01;
  assign sel_953138 = array_index_953113 == array_index_948519 ? add_953137 : sel_953134;
  assign add_953141 = sel_953138 + 8'h01;
  assign sel_953142 = array_index_953113 == array_index_948527 ? add_953141 : sel_953138;
  assign add_953145 = sel_953142 + 8'h01;
  assign sel_953146 = array_index_953113 == array_index_948535 ? add_953145 : sel_953142;
  assign add_953149 = sel_953146 + 8'h01;
  assign sel_953150 = array_index_953113 == array_index_948541 ? add_953149 : sel_953146;
  assign add_953153 = sel_953150 + 8'h01;
  assign sel_953154 = array_index_953113 == array_index_948547 ? add_953153 : sel_953150;
  assign add_953157 = sel_953154 + 8'h01;
  assign sel_953158 = array_index_953113 == array_index_948553 ? add_953157 : sel_953154;
  assign add_953161 = sel_953158 + 8'h01;
  assign sel_953162 = array_index_953113 == array_index_948559 ? add_953161 : sel_953158;
  assign add_953165 = sel_953162 + 8'h01;
  assign sel_953166 = array_index_953113 == array_index_948565 ? add_953165 : sel_953162;
  assign add_953169 = sel_953166 + 8'h01;
  assign sel_953170 = array_index_953113 == array_index_948571 ? add_953169 : sel_953166;
  assign add_953173 = sel_953170 + 8'h01;
  assign sel_953174 = array_index_953113 == array_index_948577 ? add_953173 : sel_953170;
  assign add_953177 = sel_953174 + 8'h01;
  assign sel_953178 = array_index_953113 == array_index_948583 ? add_953177 : sel_953174;
  assign add_953181 = sel_953178 + 8'h01;
  assign sel_953182 = array_index_953113 == array_index_948589 ? add_953181 : sel_953178;
  assign add_953185 = sel_953182 + 8'h01;
  assign sel_953186 = array_index_953113 == array_index_948595 ? add_953185 : sel_953182;
  assign add_953189 = sel_953186 + 8'h01;
  assign sel_953190 = array_index_953113 == array_index_948601 ? add_953189 : sel_953186;
  assign add_953193 = sel_953190 + 8'h01;
  assign sel_953194 = array_index_953113 == array_index_948607 ? add_953193 : sel_953190;
  assign add_953197 = sel_953194 + 8'h01;
  assign sel_953198 = array_index_953113 == array_index_948613 ? add_953197 : sel_953194;
  assign add_953201 = sel_953198 + 8'h01;
  assign sel_953202 = array_index_953113 == array_index_948619 ? add_953201 : sel_953198;
  assign add_953205 = sel_953202 + 8'h01;
  assign sel_953206 = array_index_953113 == array_index_948625 ? add_953205 : sel_953202;
  assign add_953209 = sel_953206 + 8'h01;
  assign sel_953210 = array_index_953113 == array_index_948631 ? add_953209 : sel_953206;
  assign add_953213 = sel_953210 + 8'h01;
  assign sel_953214 = array_index_953113 == array_index_948637 ? add_953213 : sel_953210;
  assign add_953217 = sel_953214 + 8'h01;
  assign sel_953218 = array_index_953113 == array_index_948643 ? add_953217 : sel_953214;
  assign add_953221 = sel_953218 + 8'h01;
  assign sel_953222 = array_index_953113 == array_index_948649 ? add_953221 : sel_953218;
  assign add_953225 = sel_953222 + 8'h01;
  assign sel_953226 = array_index_953113 == array_index_948655 ? add_953225 : sel_953222;
  assign add_953229 = sel_953226 + 8'h01;
  assign sel_953230 = array_index_953113 == array_index_948661 ? add_953229 : sel_953226;
  assign add_953233 = sel_953230 + 8'h01;
  assign sel_953234 = array_index_953113 == array_index_948667 ? add_953233 : sel_953230;
  assign add_953237 = sel_953234 + 8'h01;
  assign sel_953238 = array_index_953113 == array_index_948673 ? add_953237 : sel_953234;
  assign add_953241 = sel_953238 + 8'h01;
  assign sel_953242 = array_index_953113 == array_index_948679 ? add_953241 : sel_953238;
  assign add_953245 = sel_953242 + 8'h01;
  assign sel_953246 = array_index_953113 == array_index_948685 ? add_953245 : sel_953242;
  assign add_953249 = sel_953246 + 8'h01;
  assign sel_953250 = array_index_953113 == array_index_948691 ? add_953249 : sel_953246;
  assign add_953253 = sel_953250 + 8'h01;
  assign sel_953254 = array_index_953113 == array_index_948697 ? add_953253 : sel_953250;
  assign add_953257 = sel_953254 + 8'h01;
  assign sel_953258 = array_index_953113 == array_index_948703 ? add_953257 : sel_953254;
  assign add_953261 = sel_953258 + 8'h01;
  assign sel_953262 = array_index_953113 == array_index_948709 ? add_953261 : sel_953258;
  assign add_953265 = sel_953262 + 8'h01;
  assign sel_953266 = array_index_953113 == array_index_948715 ? add_953265 : sel_953262;
  assign add_953269 = sel_953266 + 8'h01;
  assign sel_953270 = array_index_953113 == array_index_948721 ? add_953269 : sel_953266;
  assign add_953273 = sel_953270 + 8'h01;
  assign sel_953274 = array_index_953113 == array_index_948727 ? add_953273 : sel_953270;
  assign add_953277 = sel_953274 + 8'h01;
  assign sel_953278 = array_index_953113 == array_index_948733 ? add_953277 : sel_953274;
  assign add_953281 = sel_953278 + 8'h01;
  assign sel_953282 = array_index_953113 == array_index_948739 ? add_953281 : sel_953278;
  assign add_953285 = sel_953282 + 8'h01;
  assign sel_953286 = array_index_953113 == array_index_948745 ? add_953285 : sel_953282;
  assign add_953289 = sel_953286 + 8'h01;
  assign sel_953290 = array_index_953113 == array_index_948751 ? add_953289 : sel_953286;
  assign add_953293 = sel_953290 + 8'h01;
  assign sel_953294 = array_index_953113 == array_index_948757 ? add_953293 : sel_953290;
  assign add_953297 = sel_953294 + 8'h01;
  assign sel_953298 = array_index_953113 == array_index_948763 ? add_953297 : sel_953294;
  assign add_953301 = sel_953298 + 8'h01;
  assign sel_953302 = array_index_953113 == array_index_948769 ? add_953301 : sel_953298;
  assign add_953305 = sel_953302 + 8'h01;
  assign sel_953306 = array_index_953113 == array_index_948775 ? add_953305 : sel_953302;
  assign add_953309 = sel_953306 + 8'h01;
  assign sel_953310 = array_index_953113 == array_index_948781 ? add_953309 : sel_953306;
  assign add_953313 = sel_953310 + 8'h01;
  assign sel_953314 = array_index_953113 == array_index_948787 ? add_953313 : sel_953310;
  assign add_953317 = sel_953314 + 8'h01;
  assign sel_953318 = array_index_953113 == array_index_948793 ? add_953317 : sel_953314;
  assign add_953321 = sel_953318 + 8'h01;
  assign sel_953322 = array_index_953113 == array_index_948799 ? add_953321 : sel_953318;
  assign add_953325 = sel_953322 + 8'h01;
  assign sel_953326 = array_index_953113 == array_index_948805 ? add_953325 : sel_953322;
  assign add_953329 = sel_953326 + 8'h01;
  assign sel_953330 = array_index_953113 == array_index_948811 ? add_953329 : sel_953326;
  assign add_953333 = sel_953330 + 8'h01;
  assign sel_953334 = array_index_953113 == array_index_948817 ? add_953333 : sel_953330;
  assign add_953337 = sel_953334 + 8'h01;
  assign sel_953338 = array_index_953113 == array_index_948823 ? add_953337 : sel_953334;
  assign add_953341 = sel_953338 + 8'h01;
  assign sel_953342 = array_index_953113 == array_index_948829 ? add_953341 : sel_953338;
  assign add_953345 = sel_953342 + 8'h01;
  assign sel_953346 = array_index_953113 == array_index_948835 ? add_953345 : sel_953342;
  assign add_953349 = sel_953346 + 8'h01;
  assign sel_953350 = array_index_953113 == array_index_948841 ? add_953349 : sel_953346;
  assign add_953353 = sel_953350 + 8'h01;
  assign sel_953354 = array_index_953113 == array_index_948847 ? add_953353 : sel_953350;
  assign add_953357 = sel_953354 + 8'h01;
  assign sel_953358 = array_index_953113 == array_index_948853 ? add_953357 : sel_953354;
  assign add_953361 = sel_953358 + 8'h01;
  assign sel_953362 = array_index_953113 == array_index_948859 ? add_953361 : sel_953358;
  assign add_953365 = sel_953362 + 8'h01;
  assign sel_953366 = array_index_953113 == array_index_948865 ? add_953365 : sel_953362;
  assign add_953369 = sel_953366 + 8'h01;
  assign sel_953370 = array_index_953113 == array_index_948871 ? add_953369 : sel_953366;
  assign add_953373 = sel_953370 + 8'h01;
  assign sel_953374 = array_index_953113 == array_index_948877 ? add_953373 : sel_953370;
  assign add_953377 = sel_953374 + 8'h01;
  assign sel_953378 = array_index_953113 == array_index_948883 ? add_953377 : sel_953374;
  assign add_953381 = sel_953378 + 8'h01;
  assign sel_953382 = array_index_953113 == array_index_948889 ? add_953381 : sel_953378;
  assign add_953385 = sel_953382 + 8'h01;
  assign sel_953386 = array_index_953113 == array_index_948895 ? add_953385 : sel_953382;
  assign add_953389 = sel_953386 + 8'h01;
  assign sel_953390 = array_index_953113 == array_index_948901 ? add_953389 : sel_953386;
  assign add_953393 = sel_953390 + 8'h01;
  assign sel_953394 = array_index_953113 == array_index_948907 ? add_953393 : sel_953390;
  assign add_953397 = sel_953394 + 8'h01;
  assign sel_953398 = array_index_953113 == array_index_948913 ? add_953397 : sel_953394;
  assign add_953401 = sel_953398 + 8'h01;
  assign sel_953402 = array_index_953113 == array_index_948919 ? add_953401 : sel_953398;
  assign add_953405 = sel_953402 + 8'h01;
  assign sel_953406 = array_index_953113 == array_index_948925 ? add_953405 : sel_953402;
  assign add_953409 = sel_953406 + 8'h01;
  assign sel_953410 = array_index_953113 == array_index_948931 ? add_953409 : sel_953406;
  assign add_953413 = sel_953410 + 8'h01;
  assign sel_953414 = array_index_953113 == array_index_948937 ? add_953413 : sel_953410;
  assign add_953417 = sel_953414 + 8'h01;
  assign sel_953418 = array_index_953113 == array_index_948943 ? add_953417 : sel_953414;
  assign add_953421 = sel_953418 + 8'h01;
  assign sel_953422 = array_index_953113 == array_index_948949 ? add_953421 : sel_953418;
  assign add_953425 = sel_953422 + 8'h01;
  assign sel_953426 = array_index_953113 == array_index_948955 ? add_953425 : sel_953422;
  assign add_953429 = sel_953426 + 8'h01;
  assign sel_953430 = array_index_953113 == array_index_948961 ? add_953429 : sel_953426;
  assign add_953433 = sel_953430 + 8'h01;
  assign sel_953434 = array_index_953113 == array_index_948967 ? add_953433 : sel_953430;
  assign add_953437 = sel_953434 + 8'h01;
  assign sel_953438 = array_index_953113 == array_index_948973 ? add_953437 : sel_953434;
  assign add_953441 = sel_953438 + 8'h01;
  assign sel_953442 = array_index_953113 == array_index_948979 ? add_953441 : sel_953438;
  assign add_953445 = sel_953442 + 8'h01;
  assign sel_953446 = array_index_953113 == array_index_948985 ? add_953445 : sel_953442;
  assign add_953449 = sel_953446 + 8'h01;
  assign sel_953450 = array_index_953113 == array_index_948991 ? add_953449 : sel_953446;
  assign add_953453 = sel_953450 + 8'h01;
  assign sel_953454 = array_index_953113 == array_index_948997 ? add_953453 : sel_953450;
  assign add_953457 = sel_953454 + 8'h01;
  assign sel_953458 = array_index_953113 == array_index_949003 ? add_953457 : sel_953454;
  assign add_953461 = sel_953458 + 8'h01;
  assign sel_953462 = array_index_953113 == array_index_949009 ? add_953461 : sel_953458;
  assign add_953465 = sel_953462 + 8'h01;
  assign sel_953466 = array_index_953113 == array_index_949015 ? add_953465 : sel_953462;
  assign add_953469 = sel_953466 + 8'h01;
  assign sel_953470 = array_index_953113 == array_index_949021 ? add_953469 : sel_953466;
  assign add_953473 = sel_953470 + 8'h01;
  assign sel_953474 = array_index_953113 == array_index_949027 ? add_953473 : sel_953470;
  assign add_953477 = sel_953474 + 8'h01;
  assign sel_953478 = array_index_953113 == array_index_949033 ? add_953477 : sel_953474;
  assign add_953481 = sel_953478 + 8'h01;
  assign sel_953482 = array_index_953113 == array_index_949039 ? add_953481 : sel_953478;
  assign add_953485 = sel_953482 + 8'h01;
  assign sel_953486 = array_index_953113 == array_index_949045 ? add_953485 : sel_953482;
  assign add_953489 = sel_953486 + 8'h01;
  assign sel_953490 = array_index_953113 == array_index_949051 ? add_953489 : sel_953486;
  assign add_953493 = sel_953490 + 8'h01;
  assign sel_953494 = array_index_953113 == array_index_949057 ? add_953493 : sel_953490;
  assign add_953497 = sel_953494 + 8'h01;
  assign sel_953498 = array_index_953113 == array_index_949063 ? add_953497 : sel_953494;
  assign add_953501 = sel_953498 + 8'h01;
  assign sel_953502 = array_index_953113 == array_index_949069 ? add_953501 : sel_953498;
  assign add_953505 = sel_953502 + 8'h01;
  assign sel_953506 = array_index_953113 == array_index_949075 ? add_953505 : sel_953502;
  assign add_953509 = sel_953506 + 8'h01;
  assign sel_953510 = array_index_953113 == array_index_949081 ? add_953509 : sel_953506;
  assign add_953514 = sel_953510 + 8'h01;
  assign array_index_953515 = set1_unflattened[7'h0c];
  assign sel_953516 = array_index_953113 == array_index_949087 ? add_953514 : sel_953510;
  assign add_953519 = sel_953516 + 8'h01;
  assign sel_953520 = array_index_953515 == array_index_948483 ? add_953519 : sel_953516;
  assign add_953523 = sel_953520 + 8'h01;
  assign sel_953524 = array_index_953515 == array_index_948487 ? add_953523 : sel_953520;
  assign add_953527 = sel_953524 + 8'h01;
  assign sel_953528 = array_index_953515 == array_index_948495 ? add_953527 : sel_953524;
  assign add_953531 = sel_953528 + 8'h01;
  assign sel_953532 = array_index_953515 == array_index_948503 ? add_953531 : sel_953528;
  assign add_953535 = sel_953532 + 8'h01;
  assign sel_953536 = array_index_953515 == array_index_948511 ? add_953535 : sel_953532;
  assign add_953539 = sel_953536 + 8'h01;
  assign sel_953540 = array_index_953515 == array_index_948519 ? add_953539 : sel_953536;
  assign add_953543 = sel_953540 + 8'h01;
  assign sel_953544 = array_index_953515 == array_index_948527 ? add_953543 : sel_953540;
  assign add_953547 = sel_953544 + 8'h01;
  assign sel_953548 = array_index_953515 == array_index_948535 ? add_953547 : sel_953544;
  assign add_953551 = sel_953548 + 8'h01;
  assign sel_953552 = array_index_953515 == array_index_948541 ? add_953551 : sel_953548;
  assign add_953555 = sel_953552 + 8'h01;
  assign sel_953556 = array_index_953515 == array_index_948547 ? add_953555 : sel_953552;
  assign add_953559 = sel_953556 + 8'h01;
  assign sel_953560 = array_index_953515 == array_index_948553 ? add_953559 : sel_953556;
  assign add_953563 = sel_953560 + 8'h01;
  assign sel_953564 = array_index_953515 == array_index_948559 ? add_953563 : sel_953560;
  assign add_953567 = sel_953564 + 8'h01;
  assign sel_953568 = array_index_953515 == array_index_948565 ? add_953567 : sel_953564;
  assign add_953571 = sel_953568 + 8'h01;
  assign sel_953572 = array_index_953515 == array_index_948571 ? add_953571 : sel_953568;
  assign add_953575 = sel_953572 + 8'h01;
  assign sel_953576 = array_index_953515 == array_index_948577 ? add_953575 : sel_953572;
  assign add_953579 = sel_953576 + 8'h01;
  assign sel_953580 = array_index_953515 == array_index_948583 ? add_953579 : sel_953576;
  assign add_953583 = sel_953580 + 8'h01;
  assign sel_953584 = array_index_953515 == array_index_948589 ? add_953583 : sel_953580;
  assign add_953587 = sel_953584 + 8'h01;
  assign sel_953588 = array_index_953515 == array_index_948595 ? add_953587 : sel_953584;
  assign add_953591 = sel_953588 + 8'h01;
  assign sel_953592 = array_index_953515 == array_index_948601 ? add_953591 : sel_953588;
  assign add_953595 = sel_953592 + 8'h01;
  assign sel_953596 = array_index_953515 == array_index_948607 ? add_953595 : sel_953592;
  assign add_953599 = sel_953596 + 8'h01;
  assign sel_953600 = array_index_953515 == array_index_948613 ? add_953599 : sel_953596;
  assign add_953603 = sel_953600 + 8'h01;
  assign sel_953604 = array_index_953515 == array_index_948619 ? add_953603 : sel_953600;
  assign add_953607 = sel_953604 + 8'h01;
  assign sel_953608 = array_index_953515 == array_index_948625 ? add_953607 : sel_953604;
  assign add_953611 = sel_953608 + 8'h01;
  assign sel_953612 = array_index_953515 == array_index_948631 ? add_953611 : sel_953608;
  assign add_953615 = sel_953612 + 8'h01;
  assign sel_953616 = array_index_953515 == array_index_948637 ? add_953615 : sel_953612;
  assign add_953619 = sel_953616 + 8'h01;
  assign sel_953620 = array_index_953515 == array_index_948643 ? add_953619 : sel_953616;
  assign add_953623 = sel_953620 + 8'h01;
  assign sel_953624 = array_index_953515 == array_index_948649 ? add_953623 : sel_953620;
  assign add_953627 = sel_953624 + 8'h01;
  assign sel_953628 = array_index_953515 == array_index_948655 ? add_953627 : sel_953624;
  assign add_953631 = sel_953628 + 8'h01;
  assign sel_953632 = array_index_953515 == array_index_948661 ? add_953631 : sel_953628;
  assign add_953635 = sel_953632 + 8'h01;
  assign sel_953636 = array_index_953515 == array_index_948667 ? add_953635 : sel_953632;
  assign add_953639 = sel_953636 + 8'h01;
  assign sel_953640 = array_index_953515 == array_index_948673 ? add_953639 : sel_953636;
  assign add_953643 = sel_953640 + 8'h01;
  assign sel_953644 = array_index_953515 == array_index_948679 ? add_953643 : sel_953640;
  assign add_953647 = sel_953644 + 8'h01;
  assign sel_953648 = array_index_953515 == array_index_948685 ? add_953647 : sel_953644;
  assign add_953651 = sel_953648 + 8'h01;
  assign sel_953652 = array_index_953515 == array_index_948691 ? add_953651 : sel_953648;
  assign add_953655 = sel_953652 + 8'h01;
  assign sel_953656 = array_index_953515 == array_index_948697 ? add_953655 : sel_953652;
  assign add_953659 = sel_953656 + 8'h01;
  assign sel_953660 = array_index_953515 == array_index_948703 ? add_953659 : sel_953656;
  assign add_953663 = sel_953660 + 8'h01;
  assign sel_953664 = array_index_953515 == array_index_948709 ? add_953663 : sel_953660;
  assign add_953667 = sel_953664 + 8'h01;
  assign sel_953668 = array_index_953515 == array_index_948715 ? add_953667 : sel_953664;
  assign add_953671 = sel_953668 + 8'h01;
  assign sel_953672 = array_index_953515 == array_index_948721 ? add_953671 : sel_953668;
  assign add_953675 = sel_953672 + 8'h01;
  assign sel_953676 = array_index_953515 == array_index_948727 ? add_953675 : sel_953672;
  assign add_953679 = sel_953676 + 8'h01;
  assign sel_953680 = array_index_953515 == array_index_948733 ? add_953679 : sel_953676;
  assign add_953683 = sel_953680 + 8'h01;
  assign sel_953684 = array_index_953515 == array_index_948739 ? add_953683 : sel_953680;
  assign add_953687 = sel_953684 + 8'h01;
  assign sel_953688 = array_index_953515 == array_index_948745 ? add_953687 : sel_953684;
  assign add_953691 = sel_953688 + 8'h01;
  assign sel_953692 = array_index_953515 == array_index_948751 ? add_953691 : sel_953688;
  assign add_953695 = sel_953692 + 8'h01;
  assign sel_953696 = array_index_953515 == array_index_948757 ? add_953695 : sel_953692;
  assign add_953699 = sel_953696 + 8'h01;
  assign sel_953700 = array_index_953515 == array_index_948763 ? add_953699 : sel_953696;
  assign add_953703 = sel_953700 + 8'h01;
  assign sel_953704 = array_index_953515 == array_index_948769 ? add_953703 : sel_953700;
  assign add_953707 = sel_953704 + 8'h01;
  assign sel_953708 = array_index_953515 == array_index_948775 ? add_953707 : sel_953704;
  assign add_953711 = sel_953708 + 8'h01;
  assign sel_953712 = array_index_953515 == array_index_948781 ? add_953711 : sel_953708;
  assign add_953715 = sel_953712 + 8'h01;
  assign sel_953716 = array_index_953515 == array_index_948787 ? add_953715 : sel_953712;
  assign add_953719 = sel_953716 + 8'h01;
  assign sel_953720 = array_index_953515 == array_index_948793 ? add_953719 : sel_953716;
  assign add_953723 = sel_953720 + 8'h01;
  assign sel_953724 = array_index_953515 == array_index_948799 ? add_953723 : sel_953720;
  assign add_953727 = sel_953724 + 8'h01;
  assign sel_953728 = array_index_953515 == array_index_948805 ? add_953727 : sel_953724;
  assign add_953731 = sel_953728 + 8'h01;
  assign sel_953732 = array_index_953515 == array_index_948811 ? add_953731 : sel_953728;
  assign add_953735 = sel_953732 + 8'h01;
  assign sel_953736 = array_index_953515 == array_index_948817 ? add_953735 : sel_953732;
  assign add_953739 = sel_953736 + 8'h01;
  assign sel_953740 = array_index_953515 == array_index_948823 ? add_953739 : sel_953736;
  assign add_953743 = sel_953740 + 8'h01;
  assign sel_953744 = array_index_953515 == array_index_948829 ? add_953743 : sel_953740;
  assign add_953747 = sel_953744 + 8'h01;
  assign sel_953748 = array_index_953515 == array_index_948835 ? add_953747 : sel_953744;
  assign add_953751 = sel_953748 + 8'h01;
  assign sel_953752 = array_index_953515 == array_index_948841 ? add_953751 : sel_953748;
  assign add_953755 = sel_953752 + 8'h01;
  assign sel_953756 = array_index_953515 == array_index_948847 ? add_953755 : sel_953752;
  assign add_953759 = sel_953756 + 8'h01;
  assign sel_953760 = array_index_953515 == array_index_948853 ? add_953759 : sel_953756;
  assign add_953763 = sel_953760 + 8'h01;
  assign sel_953764 = array_index_953515 == array_index_948859 ? add_953763 : sel_953760;
  assign add_953767 = sel_953764 + 8'h01;
  assign sel_953768 = array_index_953515 == array_index_948865 ? add_953767 : sel_953764;
  assign add_953771 = sel_953768 + 8'h01;
  assign sel_953772 = array_index_953515 == array_index_948871 ? add_953771 : sel_953768;
  assign add_953775 = sel_953772 + 8'h01;
  assign sel_953776 = array_index_953515 == array_index_948877 ? add_953775 : sel_953772;
  assign add_953779 = sel_953776 + 8'h01;
  assign sel_953780 = array_index_953515 == array_index_948883 ? add_953779 : sel_953776;
  assign add_953783 = sel_953780 + 8'h01;
  assign sel_953784 = array_index_953515 == array_index_948889 ? add_953783 : sel_953780;
  assign add_953787 = sel_953784 + 8'h01;
  assign sel_953788 = array_index_953515 == array_index_948895 ? add_953787 : sel_953784;
  assign add_953791 = sel_953788 + 8'h01;
  assign sel_953792 = array_index_953515 == array_index_948901 ? add_953791 : sel_953788;
  assign add_953795 = sel_953792 + 8'h01;
  assign sel_953796 = array_index_953515 == array_index_948907 ? add_953795 : sel_953792;
  assign add_953799 = sel_953796 + 8'h01;
  assign sel_953800 = array_index_953515 == array_index_948913 ? add_953799 : sel_953796;
  assign add_953803 = sel_953800 + 8'h01;
  assign sel_953804 = array_index_953515 == array_index_948919 ? add_953803 : sel_953800;
  assign add_953807 = sel_953804 + 8'h01;
  assign sel_953808 = array_index_953515 == array_index_948925 ? add_953807 : sel_953804;
  assign add_953811 = sel_953808 + 8'h01;
  assign sel_953812 = array_index_953515 == array_index_948931 ? add_953811 : sel_953808;
  assign add_953815 = sel_953812 + 8'h01;
  assign sel_953816 = array_index_953515 == array_index_948937 ? add_953815 : sel_953812;
  assign add_953819 = sel_953816 + 8'h01;
  assign sel_953820 = array_index_953515 == array_index_948943 ? add_953819 : sel_953816;
  assign add_953823 = sel_953820 + 8'h01;
  assign sel_953824 = array_index_953515 == array_index_948949 ? add_953823 : sel_953820;
  assign add_953827 = sel_953824 + 8'h01;
  assign sel_953828 = array_index_953515 == array_index_948955 ? add_953827 : sel_953824;
  assign add_953831 = sel_953828 + 8'h01;
  assign sel_953832 = array_index_953515 == array_index_948961 ? add_953831 : sel_953828;
  assign add_953835 = sel_953832 + 8'h01;
  assign sel_953836 = array_index_953515 == array_index_948967 ? add_953835 : sel_953832;
  assign add_953839 = sel_953836 + 8'h01;
  assign sel_953840 = array_index_953515 == array_index_948973 ? add_953839 : sel_953836;
  assign add_953843 = sel_953840 + 8'h01;
  assign sel_953844 = array_index_953515 == array_index_948979 ? add_953843 : sel_953840;
  assign add_953847 = sel_953844 + 8'h01;
  assign sel_953848 = array_index_953515 == array_index_948985 ? add_953847 : sel_953844;
  assign add_953851 = sel_953848 + 8'h01;
  assign sel_953852 = array_index_953515 == array_index_948991 ? add_953851 : sel_953848;
  assign add_953855 = sel_953852 + 8'h01;
  assign sel_953856 = array_index_953515 == array_index_948997 ? add_953855 : sel_953852;
  assign add_953859 = sel_953856 + 8'h01;
  assign sel_953860 = array_index_953515 == array_index_949003 ? add_953859 : sel_953856;
  assign add_953863 = sel_953860 + 8'h01;
  assign sel_953864 = array_index_953515 == array_index_949009 ? add_953863 : sel_953860;
  assign add_953867 = sel_953864 + 8'h01;
  assign sel_953868 = array_index_953515 == array_index_949015 ? add_953867 : sel_953864;
  assign add_953871 = sel_953868 + 8'h01;
  assign sel_953872 = array_index_953515 == array_index_949021 ? add_953871 : sel_953868;
  assign add_953875 = sel_953872 + 8'h01;
  assign sel_953876 = array_index_953515 == array_index_949027 ? add_953875 : sel_953872;
  assign add_953879 = sel_953876 + 8'h01;
  assign sel_953880 = array_index_953515 == array_index_949033 ? add_953879 : sel_953876;
  assign add_953883 = sel_953880 + 8'h01;
  assign sel_953884 = array_index_953515 == array_index_949039 ? add_953883 : sel_953880;
  assign add_953887 = sel_953884 + 8'h01;
  assign sel_953888 = array_index_953515 == array_index_949045 ? add_953887 : sel_953884;
  assign add_953891 = sel_953888 + 8'h01;
  assign sel_953892 = array_index_953515 == array_index_949051 ? add_953891 : sel_953888;
  assign add_953895 = sel_953892 + 8'h01;
  assign sel_953896 = array_index_953515 == array_index_949057 ? add_953895 : sel_953892;
  assign add_953899 = sel_953896 + 8'h01;
  assign sel_953900 = array_index_953515 == array_index_949063 ? add_953899 : sel_953896;
  assign add_953903 = sel_953900 + 8'h01;
  assign sel_953904 = array_index_953515 == array_index_949069 ? add_953903 : sel_953900;
  assign add_953907 = sel_953904 + 8'h01;
  assign sel_953908 = array_index_953515 == array_index_949075 ? add_953907 : sel_953904;
  assign add_953911 = sel_953908 + 8'h01;
  assign sel_953912 = array_index_953515 == array_index_949081 ? add_953911 : sel_953908;
  assign add_953916 = sel_953912 + 8'h01;
  assign array_index_953917 = set1_unflattened[7'h0d];
  assign sel_953918 = array_index_953515 == array_index_949087 ? add_953916 : sel_953912;
  assign add_953921 = sel_953918 + 8'h01;
  assign sel_953922 = array_index_953917 == array_index_948483 ? add_953921 : sel_953918;
  assign add_953925 = sel_953922 + 8'h01;
  assign sel_953926 = array_index_953917 == array_index_948487 ? add_953925 : sel_953922;
  assign add_953929 = sel_953926 + 8'h01;
  assign sel_953930 = array_index_953917 == array_index_948495 ? add_953929 : sel_953926;
  assign add_953933 = sel_953930 + 8'h01;
  assign sel_953934 = array_index_953917 == array_index_948503 ? add_953933 : sel_953930;
  assign add_953937 = sel_953934 + 8'h01;
  assign sel_953938 = array_index_953917 == array_index_948511 ? add_953937 : sel_953934;
  assign add_953941 = sel_953938 + 8'h01;
  assign sel_953942 = array_index_953917 == array_index_948519 ? add_953941 : sel_953938;
  assign add_953945 = sel_953942 + 8'h01;
  assign sel_953946 = array_index_953917 == array_index_948527 ? add_953945 : sel_953942;
  assign add_953949 = sel_953946 + 8'h01;
  assign sel_953950 = array_index_953917 == array_index_948535 ? add_953949 : sel_953946;
  assign add_953953 = sel_953950 + 8'h01;
  assign sel_953954 = array_index_953917 == array_index_948541 ? add_953953 : sel_953950;
  assign add_953957 = sel_953954 + 8'h01;
  assign sel_953958 = array_index_953917 == array_index_948547 ? add_953957 : sel_953954;
  assign add_953961 = sel_953958 + 8'h01;
  assign sel_953962 = array_index_953917 == array_index_948553 ? add_953961 : sel_953958;
  assign add_953965 = sel_953962 + 8'h01;
  assign sel_953966 = array_index_953917 == array_index_948559 ? add_953965 : sel_953962;
  assign add_953969 = sel_953966 + 8'h01;
  assign sel_953970 = array_index_953917 == array_index_948565 ? add_953969 : sel_953966;
  assign add_953973 = sel_953970 + 8'h01;
  assign sel_953974 = array_index_953917 == array_index_948571 ? add_953973 : sel_953970;
  assign add_953977 = sel_953974 + 8'h01;
  assign sel_953978 = array_index_953917 == array_index_948577 ? add_953977 : sel_953974;
  assign add_953981 = sel_953978 + 8'h01;
  assign sel_953982 = array_index_953917 == array_index_948583 ? add_953981 : sel_953978;
  assign add_953985 = sel_953982 + 8'h01;
  assign sel_953986 = array_index_953917 == array_index_948589 ? add_953985 : sel_953982;
  assign add_953989 = sel_953986 + 8'h01;
  assign sel_953990 = array_index_953917 == array_index_948595 ? add_953989 : sel_953986;
  assign add_953993 = sel_953990 + 8'h01;
  assign sel_953994 = array_index_953917 == array_index_948601 ? add_953993 : sel_953990;
  assign add_953997 = sel_953994 + 8'h01;
  assign sel_953998 = array_index_953917 == array_index_948607 ? add_953997 : sel_953994;
  assign add_954001 = sel_953998 + 8'h01;
  assign sel_954002 = array_index_953917 == array_index_948613 ? add_954001 : sel_953998;
  assign add_954005 = sel_954002 + 8'h01;
  assign sel_954006 = array_index_953917 == array_index_948619 ? add_954005 : sel_954002;
  assign add_954009 = sel_954006 + 8'h01;
  assign sel_954010 = array_index_953917 == array_index_948625 ? add_954009 : sel_954006;
  assign add_954013 = sel_954010 + 8'h01;
  assign sel_954014 = array_index_953917 == array_index_948631 ? add_954013 : sel_954010;
  assign add_954017 = sel_954014 + 8'h01;
  assign sel_954018 = array_index_953917 == array_index_948637 ? add_954017 : sel_954014;
  assign add_954021 = sel_954018 + 8'h01;
  assign sel_954022 = array_index_953917 == array_index_948643 ? add_954021 : sel_954018;
  assign add_954025 = sel_954022 + 8'h01;
  assign sel_954026 = array_index_953917 == array_index_948649 ? add_954025 : sel_954022;
  assign add_954029 = sel_954026 + 8'h01;
  assign sel_954030 = array_index_953917 == array_index_948655 ? add_954029 : sel_954026;
  assign add_954033 = sel_954030 + 8'h01;
  assign sel_954034 = array_index_953917 == array_index_948661 ? add_954033 : sel_954030;
  assign add_954037 = sel_954034 + 8'h01;
  assign sel_954038 = array_index_953917 == array_index_948667 ? add_954037 : sel_954034;
  assign add_954041 = sel_954038 + 8'h01;
  assign sel_954042 = array_index_953917 == array_index_948673 ? add_954041 : sel_954038;
  assign add_954045 = sel_954042 + 8'h01;
  assign sel_954046 = array_index_953917 == array_index_948679 ? add_954045 : sel_954042;
  assign add_954049 = sel_954046 + 8'h01;
  assign sel_954050 = array_index_953917 == array_index_948685 ? add_954049 : sel_954046;
  assign add_954053 = sel_954050 + 8'h01;
  assign sel_954054 = array_index_953917 == array_index_948691 ? add_954053 : sel_954050;
  assign add_954057 = sel_954054 + 8'h01;
  assign sel_954058 = array_index_953917 == array_index_948697 ? add_954057 : sel_954054;
  assign add_954061 = sel_954058 + 8'h01;
  assign sel_954062 = array_index_953917 == array_index_948703 ? add_954061 : sel_954058;
  assign add_954065 = sel_954062 + 8'h01;
  assign sel_954066 = array_index_953917 == array_index_948709 ? add_954065 : sel_954062;
  assign add_954069 = sel_954066 + 8'h01;
  assign sel_954070 = array_index_953917 == array_index_948715 ? add_954069 : sel_954066;
  assign add_954073 = sel_954070 + 8'h01;
  assign sel_954074 = array_index_953917 == array_index_948721 ? add_954073 : sel_954070;
  assign add_954077 = sel_954074 + 8'h01;
  assign sel_954078 = array_index_953917 == array_index_948727 ? add_954077 : sel_954074;
  assign add_954081 = sel_954078 + 8'h01;
  assign sel_954082 = array_index_953917 == array_index_948733 ? add_954081 : sel_954078;
  assign add_954085 = sel_954082 + 8'h01;
  assign sel_954086 = array_index_953917 == array_index_948739 ? add_954085 : sel_954082;
  assign add_954089 = sel_954086 + 8'h01;
  assign sel_954090 = array_index_953917 == array_index_948745 ? add_954089 : sel_954086;
  assign add_954093 = sel_954090 + 8'h01;
  assign sel_954094 = array_index_953917 == array_index_948751 ? add_954093 : sel_954090;
  assign add_954097 = sel_954094 + 8'h01;
  assign sel_954098 = array_index_953917 == array_index_948757 ? add_954097 : sel_954094;
  assign add_954101 = sel_954098 + 8'h01;
  assign sel_954102 = array_index_953917 == array_index_948763 ? add_954101 : sel_954098;
  assign add_954105 = sel_954102 + 8'h01;
  assign sel_954106 = array_index_953917 == array_index_948769 ? add_954105 : sel_954102;
  assign add_954109 = sel_954106 + 8'h01;
  assign sel_954110 = array_index_953917 == array_index_948775 ? add_954109 : sel_954106;
  assign add_954113 = sel_954110 + 8'h01;
  assign sel_954114 = array_index_953917 == array_index_948781 ? add_954113 : sel_954110;
  assign add_954117 = sel_954114 + 8'h01;
  assign sel_954118 = array_index_953917 == array_index_948787 ? add_954117 : sel_954114;
  assign add_954121 = sel_954118 + 8'h01;
  assign sel_954122 = array_index_953917 == array_index_948793 ? add_954121 : sel_954118;
  assign add_954125 = sel_954122 + 8'h01;
  assign sel_954126 = array_index_953917 == array_index_948799 ? add_954125 : sel_954122;
  assign add_954129 = sel_954126 + 8'h01;
  assign sel_954130 = array_index_953917 == array_index_948805 ? add_954129 : sel_954126;
  assign add_954133 = sel_954130 + 8'h01;
  assign sel_954134 = array_index_953917 == array_index_948811 ? add_954133 : sel_954130;
  assign add_954137 = sel_954134 + 8'h01;
  assign sel_954138 = array_index_953917 == array_index_948817 ? add_954137 : sel_954134;
  assign add_954141 = sel_954138 + 8'h01;
  assign sel_954142 = array_index_953917 == array_index_948823 ? add_954141 : sel_954138;
  assign add_954145 = sel_954142 + 8'h01;
  assign sel_954146 = array_index_953917 == array_index_948829 ? add_954145 : sel_954142;
  assign add_954149 = sel_954146 + 8'h01;
  assign sel_954150 = array_index_953917 == array_index_948835 ? add_954149 : sel_954146;
  assign add_954153 = sel_954150 + 8'h01;
  assign sel_954154 = array_index_953917 == array_index_948841 ? add_954153 : sel_954150;
  assign add_954157 = sel_954154 + 8'h01;
  assign sel_954158 = array_index_953917 == array_index_948847 ? add_954157 : sel_954154;
  assign add_954161 = sel_954158 + 8'h01;
  assign sel_954162 = array_index_953917 == array_index_948853 ? add_954161 : sel_954158;
  assign add_954165 = sel_954162 + 8'h01;
  assign sel_954166 = array_index_953917 == array_index_948859 ? add_954165 : sel_954162;
  assign add_954169 = sel_954166 + 8'h01;
  assign sel_954170 = array_index_953917 == array_index_948865 ? add_954169 : sel_954166;
  assign add_954173 = sel_954170 + 8'h01;
  assign sel_954174 = array_index_953917 == array_index_948871 ? add_954173 : sel_954170;
  assign add_954177 = sel_954174 + 8'h01;
  assign sel_954178 = array_index_953917 == array_index_948877 ? add_954177 : sel_954174;
  assign add_954181 = sel_954178 + 8'h01;
  assign sel_954182 = array_index_953917 == array_index_948883 ? add_954181 : sel_954178;
  assign add_954185 = sel_954182 + 8'h01;
  assign sel_954186 = array_index_953917 == array_index_948889 ? add_954185 : sel_954182;
  assign add_954189 = sel_954186 + 8'h01;
  assign sel_954190 = array_index_953917 == array_index_948895 ? add_954189 : sel_954186;
  assign add_954193 = sel_954190 + 8'h01;
  assign sel_954194 = array_index_953917 == array_index_948901 ? add_954193 : sel_954190;
  assign add_954197 = sel_954194 + 8'h01;
  assign sel_954198 = array_index_953917 == array_index_948907 ? add_954197 : sel_954194;
  assign add_954201 = sel_954198 + 8'h01;
  assign sel_954202 = array_index_953917 == array_index_948913 ? add_954201 : sel_954198;
  assign add_954205 = sel_954202 + 8'h01;
  assign sel_954206 = array_index_953917 == array_index_948919 ? add_954205 : sel_954202;
  assign add_954209 = sel_954206 + 8'h01;
  assign sel_954210 = array_index_953917 == array_index_948925 ? add_954209 : sel_954206;
  assign add_954213 = sel_954210 + 8'h01;
  assign sel_954214 = array_index_953917 == array_index_948931 ? add_954213 : sel_954210;
  assign add_954217 = sel_954214 + 8'h01;
  assign sel_954218 = array_index_953917 == array_index_948937 ? add_954217 : sel_954214;
  assign add_954221 = sel_954218 + 8'h01;
  assign sel_954222 = array_index_953917 == array_index_948943 ? add_954221 : sel_954218;
  assign add_954225 = sel_954222 + 8'h01;
  assign sel_954226 = array_index_953917 == array_index_948949 ? add_954225 : sel_954222;
  assign add_954229 = sel_954226 + 8'h01;
  assign sel_954230 = array_index_953917 == array_index_948955 ? add_954229 : sel_954226;
  assign add_954233 = sel_954230 + 8'h01;
  assign sel_954234 = array_index_953917 == array_index_948961 ? add_954233 : sel_954230;
  assign add_954237 = sel_954234 + 8'h01;
  assign sel_954238 = array_index_953917 == array_index_948967 ? add_954237 : sel_954234;
  assign add_954241 = sel_954238 + 8'h01;
  assign sel_954242 = array_index_953917 == array_index_948973 ? add_954241 : sel_954238;
  assign add_954245 = sel_954242 + 8'h01;
  assign sel_954246 = array_index_953917 == array_index_948979 ? add_954245 : sel_954242;
  assign add_954249 = sel_954246 + 8'h01;
  assign sel_954250 = array_index_953917 == array_index_948985 ? add_954249 : sel_954246;
  assign add_954253 = sel_954250 + 8'h01;
  assign sel_954254 = array_index_953917 == array_index_948991 ? add_954253 : sel_954250;
  assign add_954257 = sel_954254 + 8'h01;
  assign sel_954258 = array_index_953917 == array_index_948997 ? add_954257 : sel_954254;
  assign add_954261 = sel_954258 + 8'h01;
  assign sel_954262 = array_index_953917 == array_index_949003 ? add_954261 : sel_954258;
  assign add_954265 = sel_954262 + 8'h01;
  assign sel_954266 = array_index_953917 == array_index_949009 ? add_954265 : sel_954262;
  assign add_954269 = sel_954266 + 8'h01;
  assign sel_954270 = array_index_953917 == array_index_949015 ? add_954269 : sel_954266;
  assign add_954273 = sel_954270 + 8'h01;
  assign sel_954274 = array_index_953917 == array_index_949021 ? add_954273 : sel_954270;
  assign add_954277 = sel_954274 + 8'h01;
  assign sel_954278 = array_index_953917 == array_index_949027 ? add_954277 : sel_954274;
  assign add_954281 = sel_954278 + 8'h01;
  assign sel_954282 = array_index_953917 == array_index_949033 ? add_954281 : sel_954278;
  assign add_954285 = sel_954282 + 8'h01;
  assign sel_954286 = array_index_953917 == array_index_949039 ? add_954285 : sel_954282;
  assign add_954289 = sel_954286 + 8'h01;
  assign sel_954290 = array_index_953917 == array_index_949045 ? add_954289 : sel_954286;
  assign add_954293 = sel_954290 + 8'h01;
  assign sel_954294 = array_index_953917 == array_index_949051 ? add_954293 : sel_954290;
  assign add_954297 = sel_954294 + 8'h01;
  assign sel_954298 = array_index_953917 == array_index_949057 ? add_954297 : sel_954294;
  assign add_954301 = sel_954298 + 8'h01;
  assign sel_954302 = array_index_953917 == array_index_949063 ? add_954301 : sel_954298;
  assign add_954305 = sel_954302 + 8'h01;
  assign sel_954306 = array_index_953917 == array_index_949069 ? add_954305 : sel_954302;
  assign add_954309 = sel_954306 + 8'h01;
  assign sel_954310 = array_index_953917 == array_index_949075 ? add_954309 : sel_954306;
  assign add_954313 = sel_954310 + 8'h01;
  assign sel_954314 = array_index_953917 == array_index_949081 ? add_954313 : sel_954310;
  assign add_954318 = sel_954314 + 8'h01;
  assign array_index_954319 = set1_unflattened[7'h0e];
  assign sel_954320 = array_index_953917 == array_index_949087 ? add_954318 : sel_954314;
  assign add_954323 = sel_954320 + 8'h01;
  assign sel_954324 = array_index_954319 == array_index_948483 ? add_954323 : sel_954320;
  assign add_954327 = sel_954324 + 8'h01;
  assign sel_954328 = array_index_954319 == array_index_948487 ? add_954327 : sel_954324;
  assign add_954331 = sel_954328 + 8'h01;
  assign sel_954332 = array_index_954319 == array_index_948495 ? add_954331 : sel_954328;
  assign add_954335 = sel_954332 + 8'h01;
  assign sel_954336 = array_index_954319 == array_index_948503 ? add_954335 : sel_954332;
  assign add_954339 = sel_954336 + 8'h01;
  assign sel_954340 = array_index_954319 == array_index_948511 ? add_954339 : sel_954336;
  assign add_954343 = sel_954340 + 8'h01;
  assign sel_954344 = array_index_954319 == array_index_948519 ? add_954343 : sel_954340;
  assign add_954347 = sel_954344 + 8'h01;
  assign sel_954348 = array_index_954319 == array_index_948527 ? add_954347 : sel_954344;
  assign add_954351 = sel_954348 + 8'h01;
  assign sel_954352 = array_index_954319 == array_index_948535 ? add_954351 : sel_954348;
  assign add_954355 = sel_954352 + 8'h01;
  assign sel_954356 = array_index_954319 == array_index_948541 ? add_954355 : sel_954352;
  assign add_954359 = sel_954356 + 8'h01;
  assign sel_954360 = array_index_954319 == array_index_948547 ? add_954359 : sel_954356;
  assign add_954363 = sel_954360 + 8'h01;
  assign sel_954364 = array_index_954319 == array_index_948553 ? add_954363 : sel_954360;
  assign add_954367 = sel_954364 + 8'h01;
  assign sel_954368 = array_index_954319 == array_index_948559 ? add_954367 : sel_954364;
  assign add_954371 = sel_954368 + 8'h01;
  assign sel_954372 = array_index_954319 == array_index_948565 ? add_954371 : sel_954368;
  assign add_954375 = sel_954372 + 8'h01;
  assign sel_954376 = array_index_954319 == array_index_948571 ? add_954375 : sel_954372;
  assign add_954379 = sel_954376 + 8'h01;
  assign sel_954380 = array_index_954319 == array_index_948577 ? add_954379 : sel_954376;
  assign add_954383 = sel_954380 + 8'h01;
  assign sel_954384 = array_index_954319 == array_index_948583 ? add_954383 : sel_954380;
  assign add_954387 = sel_954384 + 8'h01;
  assign sel_954388 = array_index_954319 == array_index_948589 ? add_954387 : sel_954384;
  assign add_954391 = sel_954388 + 8'h01;
  assign sel_954392 = array_index_954319 == array_index_948595 ? add_954391 : sel_954388;
  assign add_954395 = sel_954392 + 8'h01;
  assign sel_954396 = array_index_954319 == array_index_948601 ? add_954395 : sel_954392;
  assign add_954399 = sel_954396 + 8'h01;
  assign sel_954400 = array_index_954319 == array_index_948607 ? add_954399 : sel_954396;
  assign add_954403 = sel_954400 + 8'h01;
  assign sel_954404 = array_index_954319 == array_index_948613 ? add_954403 : sel_954400;
  assign add_954407 = sel_954404 + 8'h01;
  assign sel_954408 = array_index_954319 == array_index_948619 ? add_954407 : sel_954404;
  assign add_954411 = sel_954408 + 8'h01;
  assign sel_954412 = array_index_954319 == array_index_948625 ? add_954411 : sel_954408;
  assign add_954415 = sel_954412 + 8'h01;
  assign sel_954416 = array_index_954319 == array_index_948631 ? add_954415 : sel_954412;
  assign add_954419 = sel_954416 + 8'h01;
  assign sel_954420 = array_index_954319 == array_index_948637 ? add_954419 : sel_954416;
  assign add_954423 = sel_954420 + 8'h01;
  assign sel_954424 = array_index_954319 == array_index_948643 ? add_954423 : sel_954420;
  assign add_954427 = sel_954424 + 8'h01;
  assign sel_954428 = array_index_954319 == array_index_948649 ? add_954427 : sel_954424;
  assign add_954431 = sel_954428 + 8'h01;
  assign sel_954432 = array_index_954319 == array_index_948655 ? add_954431 : sel_954428;
  assign add_954435 = sel_954432 + 8'h01;
  assign sel_954436 = array_index_954319 == array_index_948661 ? add_954435 : sel_954432;
  assign add_954439 = sel_954436 + 8'h01;
  assign sel_954440 = array_index_954319 == array_index_948667 ? add_954439 : sel_954436;
  assign add_954443 = sel_954440 + 8'h01;
  assign sel_954444 = array_index_954319 == array_index_948673 ? add_954443 : sel_954440;
  assign add_954447 = sel_954444 + 8'h01;
  assign sel_954448 = array_index_954319 == array_index_948679 ? add_954447 : sel_954444;
  assign add_954451 = sel_954448 + 8'h01;
  assign sel_954452 = array_index_954319 == array_index_948685 ? add_954451 : sel_954448;
  assign add_954455 = sel_954452 + 8'h01;
  assign sel_954456 = array_index_954319 == array_index_948691 ? add_954455 : sel_954452;
  assign add_954459 = sel_954456 + 8'h01;
  assign sel_954460 = array_index_954319 == array_index_948697 ? add_954459 : sel_954456;
  assign add_954463 = sel_954460 + 8'h01;
  assign sel_954464 = array_index_954319 == array_index_948703 ? add_954463 : sel_954460;
  assign add_954467 = sel_954464 + 8'h01;
  assign sel_954468 = array_index_954319 == array_index_948709 ? add_954467 : sel_954464;
  assign add_954471 = sel_954468 + 8'h01;
  assign sel_954472 = array_index_954319 == array_index_948715 ? add_954471 : sel_954468;
  assign add_954475 = sel_954472 + 8'h01;
  assign sel_954476 = array_index_954319 == array_index_948721 ? add_954475 : sel_954472;
  assign add_954479 = sel_954476 + 8'h01;
  assign sel_954480 = array_index_954319 == array_index_948727 ? add_954479 : sel_954476;
  assign add_954483 = sel_954480 + 8'h01;
  assign sel_954484 = array_index_954319 == array_index_948733 ? add_954483 : sel_954480;
  assign add_954487 = sel_954484 + 8'h01;
  assign sel_954488 = array_index_954319 == array_index_948739 ? add_954487 : sel_954484;
  assign add_954491 = sel_954488 + 8'h01;
  assign sel_954492 = array_index_954319 == array_index_948745 ? add_954491 : sel_954488;
  assign add_954495 = sel_954492 + 8'h01;
  assign sel_954496 = array_index_954319 == array_index_948751 ? add_954495 : sel_954492;
  assign add_954499 = sel_954496 + 8'h01;
  assign sel_954500 = array_index_954319 == array_index_948757 ? add_954499 : sel_954496;
  assign add_954503 = sel_954500 + 8'h01;
  assign sel_954504 = array_index_954319 == array_index_948763 ? add_954503 : sel_954500;
  assign add_954507 = sel_954504 + 8'h01;
  assign sel_954508 = array_index_954319 == array_index_948769 ? add_954507 : sel_954504;
  assign add_954511 = sel_954508 + 8'h01;
  assign sel_954512 = array_index_954319 == array_index_948775 ? add_954511 : sel_954508;
  assign add_954515 = sel_954512 + 8'h01;
  assign sel_954516 = array_index_954319 == array_index_948781 ? add_954515 : sel_954512;
  assign add_954519 = sel_954516 + 8'h01;
  assign sel_954520 = array_index_954319 == array_index_948787 ? add_954519 : sel_954516;
  assign add_954523 = sel_954520 + 8'h01;
  assign sel_954524 = array_index_954319 == array_index_948793 ? add_954523 : sel_954520;
  assign add_954527 = sel_954524 + 8'h01;
  assign sel_954528 = array_index_954319 == array_index_948799 ? add_954527 : sel_954524;
  assign add_954531 = sel_954528 + 8'h01;
  assign sel_954532 = array_index_954319 == array_index_948805 ? add_954531 : sel_954528;
  assign add_954535 = sel_954532 + 8'h01;
  assign sel_954536 = array_index_954319 == array_index_948811 ? add_954535 : sel_954532;
  assign add_954539 = sel_954536 + 8'h01;
  assign sel_954540 = array_index_954319 == array_index_948817 ? add_954539 : sel_954536;
  assign add_954543 = sel_954540 + 8'h01;
  assign sel_954544 = array_index_954319 == array_index_948823 ? add_954543 : sel_954540;
  assign add_954547 = sel_954544 + 8'h01;
  assign sel_954548 = array_index_954319 == array_index_948829 ? add_954547 : sel_954544;
  assign add_954551 = sel_954548 + 8'h01;
  assign sel_954552 = array_index_954319 == array_index_948835 ? add_954551 : sel_954548;
  assign add_954555 = sel_954552 + 8'h01;
  assign sel_954556 = array_index_954319 == array_index_948841 ? add_954555 : sel_954552;
  assign add_954559 = sel_954556 + 8'h01;
  assign sel_954560 = array_index_954319 == array_index_948847 ? add_954559 : sel_954556;
  assign add_954563 = sel_954560 + 8'h01;
  assign sel_954564 = array_index_954319 == array_index_948853 ? add_954563 : sel_954560;
  assign add_954567 = sel_954564 + 8'h01;
  assign sel_954568 = array_index_954319 == array_index_948859 ? add_954567 : sel_954564;
  assign add_954571 = sel_954568 + 8'h01;
  assign sel_954572 = array_index_954319 == array_index_948865 ? add_954571 : sel_954568;
  assign add_954575 = sel_954572 + 8'h01;
  assign sel_954576 = array_index_954319 == array_index_948871 ? add_954575 : sel_954572;
  assign add_954579 = sel_954576 + 8'h01;
  assign sel_954580 = array_index_954319 == array_index_948877 ? add_954579 : sel_954576;
  assign add_954583 = sel_954580 + 8'h01;
  assign sel_954584 = array_index_954319 == array_index_948883 ? add_954583 : sel_954580;
  assign add_954587 = sel_954584 + 8'h01;
  assign sel_954588 = array_index_954319 == array_index_948889 ? add_954587 : sel_954584;
  assign add_954591 = sel_954588 + 8'h01;
  assign sel_954592 = array_index_954319 == array_index_948895 ? add_954591 : sel_954588;
  assign add_954595 = sel_954592 + 8'h01;
  assign sel_954596 = array_index_954319 == array_index_948901 ? add_954595 : sel_954592;
  assign add_954599 = sel_954596 + 8'h01;
  assign sel_954600 = array_index_954319 == array_index_948907 ? add_954599 : sel_954596;
  assign add_954603 = sel_954600 + 8'h01;
  assign sel_954604 = array_index_954319 == array_index_948913 ? add_954603 : sel_954600;
  assign add_954607 = sel_954604 + 8'h01;
  assign sel_954608 = array_index_954319 == array_index_948919 ? add_954607 : sel_954604;
  assign add_954611 = sel_954608 + 8'h01;
  assign sel_954612 = array_index_954319 == array_index_948925 ? add_954611 : sel_954608;
  assign add_954615 = sel_954612 + 8'h01;
  assign sel_954616 = array_index_954319 == array_index_948931 ? add_954615 : sel_954612;
  assign add_954619 = sel_954616 + 8'h01;
  assign sel_954620 = array_index_954319 == array_index_948937 ? add_954619 : sel_954616;
  assign add_954623 = sel_954620 + 8'h01;
  assign sel_954624 = array_index_954319 == array_index_948943 ? add_954623 : sel_954620;
  assign add_954627 = sel_954624 + 8'h01;
  assign sel_954628 = array_index_954319 == array_index_948949 ? add_954627 : sel_954624;
  assign add_954631 = sel_954628 + 8'h01;
  assign sel_954632 = array_index_954319 == array_index_948955 ? add_954631 : sel_954628;
  assign add_954635 = sel_954632 + 8'h01;
  assign sel_954636 = array_index_954319 == array_index_948961 ? add_954635 : sel_954632;
  assign add_954639 = sel_954636 + 8'h01;
  assign sel_954640 = array_index_954319 == array_index_948967 ? add_954639 : sel_954636;
  assign add_954643 = sel_954640 + 8'h01;
  assign sel_954644 = array_index_954319 == array_index_948973 ? add_954643 : sel_954640;
  assign add_954647 = sel_954644 + 8'h01;
  assign sel_954648 = array_index_954319 == array_index_948979 ? add_954647 : sel_954644;
  assign add_954651 = sel_954648 + 8'h01;
  assign sel_954652 = array_index_954319 == array_index_948985 ? add_954651 : sel_954648;
  assign add_954655 = sel_954652 + 8'h01;
  assign sel_954656 = array_index_954319 == array_index_948991 ? add_954655 : sel_954652;
  assign add_954659 = sel_954656 + 8'h01;
  assign sel_954660 = array_index_954319 == array_index_948997 ? add_954659 : sel_954656;
  assign add_954663 = sel_954660 + 8'h01;
  assign sel_954664 = array_index_954319 == array_index_949003 ? add_954663 : sel_954660;
  assign add_954667 = sel_954664 + 8'h01;
  assign sel_954668 = array_index_954319 == array_index_949009 ? add_954667 : sel_954664;
  assign add_954671 = sel_954668 + 8'h01;
  assign sel_954672 = array_index_954319 == array_index_949015 ? add_954671 : sel_954668;
  assign add_954675 = sel_954672 + 8'h01;
  assign sel_954676 = array_index_954319 == array_index_949021 ? add_954675 : sel_954672;
  assign add_954679 = sel_954676 + 8'h01;
  assign sel_954680 = array_index_954319 == array_index_949027 ? add_954679 : sel_954676;
  assign add_954683 = sel_954680 + 8'h01;
  assign sel_954684 = array_index_954319 == array_index_949033 ? add_954683 : sel_954680;
  assign add_954687 = sel_954684 + 8'h01;
  assign sel_954688 = array_index_954319 == array_index_949039 ? add_954687 : sel_954684;
  assign add_954691 = sel_954688 + 8'h01;
  assign sel_954692 = array_index_954319 == array_index_949045 ? add_954691 : sel_954688;
  assign add_954695 = sel_954692 + 8'h01;
  assign sel_954696 = array_index_954319 == array_index_949051 ? add_954695 : sel_954692;
  assign add_954699 = sel_954696 + 8'h01;
  assign sel_954700 = array_index_954319 == array_index_949057 ? add_954699 : sel_954696;
  assign add_954703 = sel_954700 + 8'h01;
  assign sel_954704 = array_index_954319 == array_index_949063 ? add_954703 : sel_954700;
  assign add_954707 = sel_954704 + 8'h01;
  assign sel_954708 = array_index_954319 == array_index_949069 ? add_954707 : sel_954704;
  assign add_954711 = sel_954708 + 8'h01;
  assign sel_954712 = array_index_954319 == array_index_949075 ? add_954711 : sel_954708;
  assign add_954715 = sel_954712 + 8'h01;
  assign sel_954716 = array_index_954319 == array_index_949081 ? add_954715 : sel_954712;
  assign add_954720 = sel_954716 + 8'h01;
  assign array_index_954721 = set1_unflattened[7'h0f];
  assign sel_954722 = array_index_954319 == array_index_949087 ? add_954720 : sel_954716;
  assign add_954725 = sel_954722 + 8'h01;
  assign sel_954726 = array_index_954721 == array_index_948483 ? add_954725 : sel_954722;
  assign add_954729 = sel_954726 + 8'h01;
  assign sel_954730 = array_index_954721 == array_index_948487 ? add_954729 : sel_954726;
  assign add_954733 = sel_954730 + 8'h01;
  assign sel_954734 = array_index_954721 == array_index_948495 ? add_954733 : sel_954730;
  assign add_954737 = sel_954734 + 8'h01;
  assign sel_954738 = array_index_954721 == array_index_948503 ? add_954737 : sel_954734;
  assign add_954741 = sel_954738 + 8'h01;
  assign sel_954742 = array_index_954721 == array_index_948511 ? add_954741 : sel_954738;
  assign add_954745 = sel_954742 + 8'h01;
  assign sel_954746 = array_index_954721 == array_index_948519 ? add_954745 : sel_954742;
  assign add_954749 = sel_954746 + 8'h01;
  assign sel_954750 = array_index_954721 == array_index_948527 ? add_954749 : sel_954746;
  assign add_954753 = sel_954750 + 8'h01;
  assign sel_954754 = array_index_954721 == array_index_948535 ? add_954753 : sel_954750;
  assign add_954757 = sel_954754 + 8'h01;
  assign sel_954758 = array_index_954721 == array_index_948541 ? add_954757 : sel_954754;
  assign add_954761 = sel_954758 + 8'h01;
  assign sel_954762 = array_index_954721 == array_index_948547 ? add_954761 : sel_954758;
  assign add_954765 = sel_954762 + 8'h01;
  assign sel_954766 = array_index_954721 == array_index_948553 ? add_954765 : sel_954762;
  assign add_954769 = sel_954766 + 8'h01;
  assign sel_954770 = array_index_954721 == array_index_948559 ? add_954769 : sel_954766;
  assign add_954773 = sel_954770 + 8'h01;
  assign sel_954774 = array_index_954721 == array_index_948565 ? add_954773 : sel_954770;
  assign add_954777 = sel_954774 + 8'h01;
  assign sel_954778 = array_index_954721 == array_index_948571 ? add_954777 : sel_954774;
  assign add_954781 = sel_954778 + 8'h01;
  assign sel_954782 = array_index_954721 == array_index_948577 ? add_954781 : sel_954778;
  assign add_954785 = sel_954782 + 8'h01;
  assign sel_954786 = array_index_954721 == array_index_948583 ? add_954785 : sel_954782;
  assign add_954789 = sel_954786 + 8'h01;
  assign sel_954790 = array_index_954721 == array_index_948589 ? add_954789 : sel_954786;
  assign add_954793 = sel_954790 + 8'h01;
  assign sel_954794 = array_index_954721 == array_index_948595 ? add_954793 : sel_954790;
  assign add_954797 = sel_954794 + 8'h01;
  assign sel_954798 = array_index_954721 == array_index_948601 ? add_954797 : sel_954794;
  assign add_954801 = sel_954798 + 8'h01;
  assign sel_954802 = array_index_954721 == array_index_948607 ? add_954801 : sel_954798;
  assign add_954805 = sel_954802 + 8'h01;
  assign sel_954806 = array_index_954721 == array_index_948613 ? add_954805 : sel_954802;
  assign add_954809 = sel_954806 + 8'h01;
  assign sel_954810 = array_index_954721 == array_index_948619 ? add_954809 : sel_954806;
  assign add_954813 = sel_954810 + 8'h01;
  assign sel_954814 = array_index_954721 == array_index_948625 ? add_954813 : sel_954810;
  assign add_954817 = sel_954814 + 8'h01;
  assign sel_954818 = array_index_954721 == array_index_948631 ? add_954817 : sel_954814;
  assign add_954821 = sel_954818 + 8'h01;
  assign sel_954822 = array_index_954721 == array_index_948637 ? add_954821 : sel_954818;
  assign add_954825 = sel_954822 + 8'h01;
  assign sel_954826 = array_index_954721 == array_index_948643 ? add_954825 : sel_954822;
  assign add_954829 = sel_954826 + 8'h01;
  assign sel_954830 = array_index_954721 == array_index_948649 ? add_954829 : sel_954826;
  assign add_954833 = sel_954830 + 8'h01;
  assign sel_954834 = array_index_954721 == array_index_948655 ? add_954833 : sel_954830;
  assign add_954837 = sel_954834 + 8'h01;
  assign sel_954838 = array_index_954721 == array_index_948661 ? add_954837 : sel_954834;
  assign add_954841 = sel_954838 + 8'h01;
  assign sel_954842 = array_index_954721 == array_index_948667 ? add_954841 : sel_954838;
  assign add_954845 = sel_954842 + 8'h01;
  assign sel_954846 = array_index_954721 == array_index_948673 ? add_954845 : sel_954842;
  assign add_954849 = sel_954846 + 8'h01;
  assign sel_954850 = array_index_954721 == array_index_948679 ? add_954849 : sel_954846;
  assign add_954853 = sel_954850 + 8'h01;
  assign sel_954854 = array_index_954721 == array_index_948685 ? add_954853 : sel_954850;
  assign add_954857 = sel_954854 + 8'h01;
  assign sel_954858 = array_index_954721 == array_index_948691 ? add_954857 : sel_954854;
  assign add_954861 = sel_954858 + 8'h01;
  assign sel_954862 = array_index_954721 == array_index_948697 ? add_954861 : sel_954858;
  assign add_954865 = sel_954862 + 8'h01;
  assign sel_954866 = array_index_954721 == array_index_948703 ? add_954865 : sel_954862;
  assign add_954869 = sel_954866 + 8'h01;
  assign sel_954870 = array_index_954721 == array_index_948709 ? add_954869 : sel_954866;
  assign add_954873 = sel_954870 + 8'h01;
  assign sel_954874 = array_index_954721 == array_index_948715 ? add_954873 : sel_954870;
  assign add_954877 = sel_954874 + 8'h01;
  assign sel_954878 = array_index_954721 == array_index_948721 ? add_954877 : sel_954874;
  assign add_954881 = sel_954878 + 8'h01;
  assign sel_954882 = array_index_954721 == array_index_948727 ? add_954881 : sel_954878;
  assign add_954885 = sel_954882 + 8'h01;
  assign sel_954886 = array_index_954721 == array_index_948733 ? add_954885 : sel_954882;
  assign add_954889 = sel_954886 + 8'h01;
  assign sel_954890 = array_index_954721 == array_index_948739 ? add_954889 : sel_954886;
  assign add_954893 = sel_954890 + 8'h01;
  assign sel_954894 = array_index_954721 == array_index_948745 ? add_954893 : sel_954890;
  assign add_954897 = sel_954894 + 8'h01;
  assign sel_954898 = array_index_954721 == array_index_948751 ? add_954897 : sel_954894;
  assign add_954901 = sel_954898 + 8'h01;
  assign sel_954902 = array_index_954721 == array_index_948757 ? add_954901 : sel_954898;
  assign add_954905 = sel_954902 + 8'h01;
  assign sel_954906 = array_index_954721 == array_index_948763 ? add_954905 : sel_954902;
  assign add_954909 = sel_954906 + 8'h01;
  assign sel_954910 = array_index_954721 == array_index_948769 ? add_954909 : sel_954906;
  assign add_954913 = sel_954910 + 8'h01;
  assign sel_954914 = array_index_954721 == array_index_948775 ? add_954913 : sel_954910;
  assign add_954917 = sel_954914 + 8'h01;
  assign sel_954918 = array_index_954721 == array_index_948781 ? add_954917 : sel_954914;
  assign add_954921 = sel_954918 + 8'h01;
  assign sel_954922 = array_index_954721 == array_index_948787 ? add_954921 : sel_954918;
  assign add_954925 = sel_954922 + 8'h01;
  assign sel_954926 = array_index_954721 == array_index_948793 ? add_954925 : sel_954922;
  assign add_954929 = sel_954926 + 8'h01;
  assign sel_954930 = array_index_954721 == array_index_948799 ? add_954929 : sel_954926;
  assign add_954933 = sel_954930 + 8'h01;
  assign sel_954934 = array_index_954721 == array_index_948805 ? add_954933 : sel_954930;
  assign add_954937 = sel_954934 + 8'h01;
  assign sel_954938 = array_index_954721 == array_index_948811 ? add_954937 : sel_954934;
  assign add_954941 = sel_954938 + 8'h01;
  assign sel_954942 = array_index_954721 == array_index_948817 ? add_954941 : sel_954938;
  assign add_954945 = sel_954942 + 8'h01;
  assign sel_954946 = array_index_954721 == array_index_948823 ? add_954945 : sel_954942;
  assign add_954949 = sel_954946 + 8'h01;
  assign sel_954950 = array_index_954721 == array_index_948829 ? add_954949 : sel_954946;
  assign add_954953 = sel_954950 + 8'h01;
  assign sel_954954 = array_index_954721 == array_index_948835 ? add_954953 : sel_954950;
  assign add_954957 = sel_954954 + 8'h01;
  assign sel_954958 = array_index_954721 == array_index_948841 ? add_954957 : sel_954954;
  assign add_954961 = sel_954958 + 8'h01;
  assign sel_954962 = array_index_954721 == array_index_948847 ? add_954961 : sel_954958;
  assign add_954965 = sel_954962 + 8'h01;
  assign sel_954966 = array_index_954721 == array_index_948853 ? add_954965 : sel_954962;
  assign add_954969 = sel_954966 + 8'h01;
  assign sel_954970 = array_index_954721 == array_index_948859 ? add_954969 : sel_954966;
  assign add_954973 = sel_954970 + 8'h01;
  assign sel_954974 = array_index_954721 == array_index_948865 ? add_954973 : sel_954970;
  assign add_954977 = sel_954974 + 8'h01;
  assign sel_954978 = array_index_954721 == array_index_948871 ? add_954977 : sel_954974;
  assign add_954981 = sel_954978 + 8'h01;
  assign sel_954982 = array_index_954721 == array_index_948877 ? add_954981 : sel_954978;
  assign add_954985 = sel_954982 + 8'h01;
  assign sel_954986 = array_index_954721 == array_index_948883 ? add_954985 : sel_954982;
  assign add_954989 = sel_954986 + 8'h01;
  assign sel_954990 = array_index_954721 == array_index_948889 ? add_954989 : sel_954986;
  assign add_954993 = sel_954990 + 8'h01;
  assign sel_954994 = array_index_954721 == array_index_948895 ? add_954993 : sel_954990;
  assign add_954997 = sel_954994 + 8'h01;
  assign sel_954998 = array_index_954721 == array_index_948901 ? add_954997 : sel_954994;
  assign add_955001 = sel_954998 + 8'h01;
  assign sel_955002 = array_index_954721 == array_index_948907 ? add_955001 : sel_954998;
  assign add_955005 = sel_955002 + 8'h01;
  assign sel_955006 = array_index_954721 == array_index_948913 ? add_955005 : sel_955002;
  assign add_955009 = sel_955006 + 8'h01;
  assign sel_955010 = array_index_954721 == array_index_948919 ? add_955009 : sel_955006;
  assign add_955013 = sel_955010 + 8'h01;
  assign sel_955014 = array_index_954721 == array_index_948925 ? add_955013 : sel_955010;
  assign add_955017 = sel_955014 + 8'h01;
  assign sel_955018 = array_index_954721 == array_index_948931 ? add_955017 : sel_955014;
  assign add_955021 = sel_955018 + 8'h01;
  assign sel_955022 = array_index_954721 == array_index_948937 ? add_955021 : sel_955018;
  assign add_955025 = sel_955022 + 8'h01;
  assign sel_955026 = array_index_954721 == array_index_948943 ? add_955025 : sel_955022;
  assign add_955029 = sel_955026 + 8'h01;
  assign sel_955030 = array_index_954721 == array_index_948949 ? add_955029 : sel_955026;
  assign add_955033 = sel_955030 + 8'h01;
  assign sel_955034 = array_index_954721 == array_index_948955 ? add_955033 : sel_955030;
  assign add_955037 = sel_955034 + 8'h01;
  assign sel_955038 = array_index_954721 == array_index_948961 ? add_955037 : sel_955034;
  assign add_955041 = sel_955038 + 8'h01;
  assign sel_955042 = array_index_954721 == array_index_948967 ? add_955041 : sel_955038;
  assign add_955045 = sel_955042 + 8'h01;
  assign sel_955046 = array_index_954721 == array_index_948973 ? add_955045 : sel_955042;
  assign add_955049 = sel_955046 + 8'h01;
  assign sel_955050 = array_index_954721 == array_index_948979 ? add_955049 : sel_955046;
  assign add_955053 = sel_955050 + 8'h01;
  assign sel_955054 = array_index_954721 == array_index_948985 ? add_955053 : sel_955050;
  assign add_955057 = sel_955054 + 8'h01;
  assign sel_955058 = array_index_954721 == array_index_948991 ? add_955057 : sel_955054;
  assign add_955061 = sel_955058 + 8'h01;
  assign sel_955062 = array_index_954721 == array_index_948997 ? add_955061 : sel_955058;
  assign add_955065 = sel_955062 + 8'h01;
  assign sel_955066 = array_index_954721 == array_index_949003 ? add_955065 : sel_955062;
  assign add_955069 = sel_955066 + 8'h01;
  assign sel_955070 = array_index_954721 == array_index_949009 ? add_955069 : sel_955066;
  assign add_955073 = sel_955070 + 8'h01;
  assign sel_955074 = array_index_954721 == array_index_949015 ? add_955073 : sel_955070;
  assign add_955077 = sel_955074 + 8'h01;
  assign sel_955078 = array_index_954721 == array_index_949021 ? add_955077 : sel_955074;
  assign add_955081 = sel_955078 + 8'h01;
  assign sel_955082 = array_index_954721 == array_index_949027 ? add_955081 : sel_955078;
  assign add_955085 = sel_955082 + 8'h01;
  assign sel_955086 = array_index_954721 == array_index_949033 ? add_955085 : sel_955082;
  assign add_955089 = sel_955086 + 8'h01;
  assign sel_955090 = array_index_954721 == array_index_949039 ? add_955089 : sel_955086;
  assign add_955093 = sel_955090 + 8'h01;
  assign sel_955094 = array_index_954721 == array_index_949045 ? add_955093 : sel_955090;
  assign add_955097 = sel_955094 + 8'h01;
  assign sel_955098 = array_index_954721 == array_index_949051 ? add_955097 : sel_955094;
  assign add_955101 = sel_955098 + 8'h01;
  assign sel_955102 = array_index_954721 == array_index_949057 ? add_955101 : sel_955098;
  assign add_955105 = sel_955102 + 8'h01;
  assign sel_955106 = array_index_954721 == array_index_949063 ? add_955105 : sel_955102;
  assign add_955109 = sel_955106 + 8'h01;
  assign sel_955110 = array_index_954721 == array_index_949069 ? add_955109 : sel_955106;
  assign add_955113 = sel_955110 + 8'h01;
  assign sel_955114 = array_index_954721 == array_index_949075 ? add_955113 : sel_955110;
  assign add_955117 = sel_955114 + 8'h01;
  assign sel_955118 = array_index_954721 == array_index_949081 ? add_955117 : sel_955114;
  assign add_955122 = sel_955118 + 8'h01;
  assign array_index_955123 = set1_unflattened[7'h10];
  assign sel_955124 = array_index_954721 == array_index_949087 ? add_955122 : sel_955118;
  assign add_955127 = sel_955124 + 8'h01;
  assign sel_955128 = array_index_955123 == array_index_948483 ? add_955127 : sel_955124;
  assign add_955131 = sel_955128 + 8'h01;
  assign sel_955132 = array_index_955123 == array_index_948487 ? add_955131 : sel_955128;
  assign add_955135 = sel_955132 + 8'h01;
  assign sel_955136 = array_index_955123 == array_index_948495 ? add_955135 : sel_955132;
  assign add_955139 = sel_955136 + 8'h01;
  assign sel_955140 = array_index_955123 == array_index_948503 ? add_955139 : sel_955136;
  assign add_955143 = sel_955140 + 8'h01;
  assign sel_955144 = array_index_955123 == array_index_948511 ? add_955143 : sel_955140;
  assign add_955147 = sel_955144 + 8'h01;
  assign sel_955148 = array_index_955123 == array_index_948519 ? add_955147 : sel_955144;
  assign add_955151 = sel_955148 + 8'h01;
  assign sel_955152 = array_index_955123 == array_index_948527 ? add_955151 : sel_955148;
  assign add_955155 = sel_955152 + 8'h01;
  assign sel_955156 = array_index_955123 == array_index_948535 ? add_955155 : sel_955152;
  assign add_955159 = sel_955156 + 8'h01;
  assign sel_955160 = array_index_955123 == array_index_948541 ? add_955159 : sel_955156;
  assign add_955163 = sel_955160 + 8'h01;
  assign sel_955164 = array_index_955123 == array_index_948547 ? add_955163 : sel_955160;
  assign add_955167 = sel_955164 + 8'h01;
  assign sel_955168 = array_index_955123 == array_index_948553 ? add_955167 : sel_955164;
  assign add_955171 = sel_955168 + 8'h01;
  assign sel_955172 = array_index_955123 == array_index_948559 ? add_955171 : sel_955168;
  assign add_955175 = sel_955172 + 8'h01;
  assign sel_955176 = array_index_955123 == array_index_948565 ? add_955175 : sel_955172;
  assign add_955179 = sel_955176 + 8'h01;
  assign sel_955180 = array_index_955123 == array_index_948571 ? add_955179 : sel_955176;
  assign add_955183 = sel_955180 + 8'h01;
  assign sel_955184 = array_index_955123 == array_index_948577 ? add_955183 : sel_955180;
  assign add_955187 = sel_955184 + 8'h01;
  assign sel_955188 = array_index_955123 == array_index_948583 ? add_955187 : sel_955184;
  assign add_955191 = sel_955188 + 8'h01;
  assign sel_955192 = array_index_955123 == array_index_948589 ? add_955191 : sel_955188;
  assign add_955195 = sel_955192 + 8'h01;
  assign sel_955196 = array_index_955123 == array_index_948595 ? add_955195 : sel_955192;
  assign add_955199 = sel_955196 + 8'h01;
  assign sel_955200 = array_index_955123 == array_index_948601 ? add_955199 : sel_955196;
  assign add_955203 = sel_955200 + 8'h01;
  assign sel_955204 = array_index_955123 == array_index_948607 ? add_955203 : sel_955200;
  assign add_955207 = sel_955204 + 8'h01;
  assign sel_955208 = array_index_955123 == array_index_948613 ? add_955207 : sel_955204;
  assign add_955211 = sel_955208 + 8'h01;
  assign sel_955212 = array_index_955123 == array_index_948619 ? add_955211 : sel_955208;
  assign add_955215 = sel_955212 + 8'h01;
  assign sel_955216 = array_index_955123 == array_index_948625 ? add_955215 : sel_955212;
  assign add_955219 = sel_955216 + 8'h01;
  assign sel_955220 = array_index_955123 == array_index_948631 ? add_955219 : sel_955216;
  assign add_955223 = sel_955220 + 8'h01;
  assign sel_955224 = array_index_955123 == array_index_948637 ? add_955223 : sel_955220;
  assign add_955227 = sel_955224 + 8'h01;
  assign sel_955228 = array_index_955123 == array_index_948643 ? add_955227 : sel_955224;
  assign add_955231 = sel_955228 + 8'h01;
  assign sel_955232 = array_index_955123 == array_index_948649 ? add_955231 : sel_955228;
  assign add_955235 = sel_955232 + 8'h01;
  assign sel_955236 = array_index_955123 == array_index_948655 ? add_955235 : sel_955232;
  assign add_955239 = sel_955236 + 8'h01;
  assign sel_955240 = array_index_955123 == array_index_948661 ? add_955239 : sel_955236;
  assign add_955243 = sel_955240 + 8'h01;
  assign sel_955244 = array_index_955123 == array_index_948667 ? add_955243 : sel_955240;
  assign add_955247 = sel_955244 + 8'h01;
  assign sel_955248 = array_index_955123 == array_index_948673 ? add_955247 : sel_955244;
  assign add_955251 = sel_955248 + 8'h01;
  assign sel_955252 = array_index_955123 == array_index_948679 ? add_955251 : sel_955248;
  assign add_955255 = sel_955252 + 8'h01;
  assign sel_955256 = array_index_955123 == array_index_948685 ? add_955255 : sel_955252;
  assign add_955259 = sel_955256 + 8'h01;
  assign sel_955260 = array_index_955123 == array_index_948691 ? add_955259 : sel_955256;
  assign add_955263 = sel_955260 + 8'h01;
  assign sel_955264 = array_index_955123 == array_index_948697 ? add_955263 : sel_955260;
  assign add_955267 = sel_955264 + 8'h01;
  assign sel_955268 = array_index_955123 == array_index_948703 ? add_955267 : sel_955264;
  assign add_955271 = sel_955268 + 8'h01;
  assign sel_955272 = array_index_955123 == array_index_948709 ? add_955271 : sel_955268;
  assign add_955275 = sel_955272 + 8'h01;
  assign sel_955276 = array_index_955123 == array_index_948715 ? add_955275 : sel_955272;
  assign add_955279 = sel_955276 + 8'h01;
  assign sel_955280 = array_index_955123 == array_index_948721 ? add_955279 : sel_955276;
  assign add_955283 = sel_955280 + 8'h01;
  assign sel_955284 = array_index_955123 == array_index_948727 ? add_955283 : sel_955280;
  assign add_955287 = sel_955284 + 8'h01;
  assign sel_955288 = array_index_955123 == array_index_948733 ? add_955287 : sel_955284;
  assign add_955291 = sel_955288 + 8'h01;
  assign sel_955292 = array_index_955123 == array_index_948739 ? add_955291 : sel_955288;
  assign add_955295 = sel_955292 + 8'h01;
  assign sel_955296 = array_index_955123 == array_index_948745 ? add_955295 : sel_955292;
  assign add_955299 = sel_955296 + 8'h01;
  assign sel_955300 = array_index_955123 == array_index_948751 ? add_955299 : sel_955296;
  assign add_955303 = sel_955300 + 8'h01;
  assign sel_955304 = array_index_955123 == array_index_948757 ? add_955303 : sel_955300;
  assign add_955307 = sel_955304 + 8'h01;
  assign sel_955308 = array_index_955123 == array_index_948763 ? add_955307 : sel_955304;
  assign add_955311 = sel_955308 + 8'h01;
  assign sel_955312 = array_index_955123 == array_index_948769 ? add_955311 : sel_955308;
  assign add_955315 = sel_955312 + 8'h01;
  assign sel_955316 = array_index_955123 == array_index_948775 ? add_955315 : sel_955312;
  assign add_955319 = sel_955316 + 8'h01;
  assign sel_955320 = array_index_955123 == array_index_948781 ? add_955319 : sel_955316;
  assign add_955323 = sel_955320 + 8'h01;
  assign sel_955324 = array_index_955123 == array_index_948787 ? add_955323 : sel_955320;
  assign add_955327 = sel_955324 + 8'h01;
  assign sel_955328 = array_index_955123 == array_index_948793 ? add_955327 : sel_955324;
  assign add_955331 = sel_955328 + 8'h01;
  assign sel_955332 = array_index_955123 == array_index_948799 ? add_955331 : sel_955328;
  assign add_955335 = sel_955332 + 8'h01;
  assign sel_955336 = array_index_955123 == array_index_948805 ? add_955335 : sel_955332;
  assign add_955339 = sel_955336 + 8'h01;
  assign sel_955340 = array_index_955123 == array_index_948811 ? add_955339 : sel_955336;
  assign add_955343 = sel_955340 + 8'h01;
  assign sel_955344 = array_index_955123 == array_index_948817 ? add_955343 : sel_955340;
  assign add_955347 = sel_955344 + 8'h01;
  assign sel_955348 = array_index_955123 == array_index_948823 ? add_955347 : sel_955344;
  assign add_955351 = sel_955348 + 8'h01;
  assign sel_955352 = array_index_955123 == array_index_948829 ? add_955351 : sel_955348;
  assign add_955355 = sel_955352 + 8'h01;
  assign sel_955356 = array_index_955123 == array_index_948835 ? add_955355 : sel_955352;
  assign add_955359 = sel_955356 + 8'h01;
  assign sel_955360 = array_index_955123 == array_index_948841 ? add_955359 : sel_955356;
  assign add_955363 = sel_955360 + 8'h01;
  assign sel_955364 = array_index_955123 == array_index_948847 ? add_955363 : sel_955360;
  assign add_955367 = sel_955364 + 8'h01;
  assign sel_955368 = array_index_955123 == array_index_948853 ? add_955367 : sel_955364;
  assign add_955371 = sel_955368 + 8'h01;
  assign sel_955372 = array_index_955123 == array_index_948859 ? add_955371 : sel_955368;
  assign add_955375 = sel_955372 + 8'h01;
  assign sel_955376 = array_index_955123 == array_index_948865 ? add_955375 : sel_955372;
  assign add_955379 = sel_955376 + 8'h01;
  assign sel_955380 = array_index_955123 == array_index_948871 ? add_955379 : sel_955376;
  assign add_955383 = sel_955380 + 8'h01;
  assign sel_955384 = array_index_955123 == array_index_948877 ? add_955383 : sel_955380;
  assign add_955387 = sel_955384 + 8'h01;
  assign sel_955388 = array_index_955123 == array_index_948883 ? add_955387 : sel_955384;
  assign add_955391 = sel_955388 + 8'h01;
  assign sel_955392 = array_index_955123 == array_index_948889 ? add_955391 : sel_955388;
  assign add_955395 = sel_955392 + 8'h01;
  assign sel_955396 = array_index_955123 == array_index_948895 ? add_955395 : sel_955392;
  assign add_955399 = sel_955396 + 8'h01;
  assign sel_955400 = array_index_955123 == array_index_948901 ? add_955399 : sel_955396;
  assign add_955403 = sel_955400 + 8'h01;
  assign sel_955404 = array_index_955123 == array_index_948907 ? add_955403 : sel_955400;
  assign add_955407 = sel_955404 + 8'h01;
  assign sel_955408 = array_index_955123 == array_index_948913 ? add_955407 : sel_955404;
  assign add_955411 = sel_955408 + 8'h01;
  assign sel_955412 = array_index_955123 == array_index_948919 ? add_955411 : sel_955408;
  assign add_955415 = sel_955412 + 8'h01;
  assign sel_955416 = array_index_955123 == array_index_948925 ? add_955415 : sel_955412;
  assign add_955419 = sel_955416 + 8'h01;
  assign sel_955420 = array_index_955123 == array_index_948931 ? add_955419 : sel_955416;
  assign add_955423 = sel_955420 + 8'h01;
  assign sel_955424 = array_index_955123 == array_index_948937 ? add_955423 : sel_955420;
  assign add_955427 = sel_955424 + 8'h01;
  assign sel_955428 = array_index_955123 == array_index_948943 ? add_955427 : sel_955424;
  assign add_955431 = sel_955428 + 8'h01;
  assign sel_955432 = array_index_955123 == array_index_948949 ? add_955431 : sel_955428;
  assign add_955435 = sel_955432 + 8'h01;
  assign sel_955436 = array_index_955123 == array_index_948955 ? add_955435 : sel_955432;
  assign add_955439 = sel_955436 + 8'h01;
  assign sel_955440 = array_index_955123 == array_index_948961 ? add_955439 : sel_955436;
  assign add_955443 = sel_955440 + 8'h01;
  assign sel_955444 = array_index_955123 == array_index_948967 ? add_955443 : sel_955440;
  assign add_955447 = sel_955444 + 8'h01;
  assign sel_955448 = array_index_955123 == array_index_948973 ? add_955447 : sel_955444;
  assign add_955451 = sel_955448 + 8'h01;
  assign sel_955452 = array_index_955123 == array_index_948979 ? add_955451 : sel_955448;
  assign add_955455 = sel_955452 + 8'h01;
  assign sel_955456 = array_index_955123 == array_index_948985 ? add_955455 : sel_955452;
  assign add_955459 = sel_955456 + 8'h01;
  assign sel_955460 = array_index_955123 == array_index_948991 ? add_955459 : sel_955456;
  assign add_955463 = sel_955460 + 8'h01;
  assign sel_955464 = array_index_955123 == array_index_948997 ? add_955463 : sel_955460;
  assign add_955467 = sel_955464 + 8'h01;
  assign sel_955468 = array_index_955123 == array_index_949003 ? add_955467 : sel_955464;
  assign add_955471 = sel_955468 + 8'h01;
  assign sel_955472 = array_index_955123 == array_index_949009 ? add_955471 : sel_955468;
  assign add_955475 = sel_955472 + 8'h01;
  assign sel_955476 = array_index_955123 == array_index_949015 ? add_955475 : sel_955472;
  assign add_955479 = sel_955476 + 8'h01;
  assign sel_955480 = array_index_955123 == array_index_949021 ? add_955479 : sel_955476;
  assign add_955483 = sel_955480 + 8'h01;
  assign sel_955484 = array_index_955123 == array_index_949027 ? add_955483 : sel_955480;
  assign add_955487 = sel_955484 + 8'h01;
  assign sel_955488 = array_index_955123 == array_index_949033 ? add_955487 : sel_955484;
  assign add_955491 = sel_955488 + 8'h01;
  assign sel_955492 = array_index_955123 == array_index_949039 ? add_955491 : sel_955488;
  assign add_955495 = sel_955492 + 8'h01;
  assign sel_955496 = array_index_955123 == array_index_949045 ? add_955495 : sel_955492;
  assign add_955499 = sel_955496 + 8'h01;
  assign sel_955500 = array_index_955123 == array_index_949051 ? add_955499 : sel_955496;
  assign add_955503 = sel_955500 + 8'h01;
  assign sel_955504 = array_index_955123 == array_index_949057 ? add_955503 : sel_955500;
  assign add_955507 = sel_955504 + 8'h01;
  assign sel_955508 = array_index_955123 == array_index_949063 ? add_955507 : sel_955504;
  assign add_955511 = sel_955508 + 8'h01;
  assign sel_955512 = array_index_955123 == array_index_949069 ? add_955511 : sel_955508;
  assign add_955515 = sel_955512 + 8'h01;
  assign sel_955516 = array_index_955123 == array_index_949075 ? add_955515 : sel_955512;
  assign add_955519 = sel_955516 + 8'h01;
  assign sel_955520 = array_index_955123 == array_index_949081 ? add_955519 : sel_955516;
  assign add_955524 = sel_955520 + 8'h01;
  assign array_index_955525 = set1_unflattened[7'h11];
  assign sel_955526 = array_index_955123 == array_index_949087 ? add_955524 : sel_955520;
  assign add_955529 = sel_955526 + 8'h01;
  assign sel_955530 = array_index_955525 == array_index_948483 ? add_955529 : sel_955526;
  assign add_955533 = sel_955530 + 8'h01;
  assign sel_955534 = array_index_955525 == array_index_948487 ? add_955533 : sel_955530;
  assign add_955537 = sel_955534 + 8'h01;
  assign sel_955538 = array_index_955525 == array_index_948495 ? add_955537 : sel_955534;
  assign add_955541 = sel_955538 + 8'h01;
  assign sel_955542 = array_index_955525 == array_index_948503 ? add_955541 : sel_955538;
  assign add_955545 = sel_955542 + 8'h01;
  assign sel_955546 = array_index_955525 == array_index_948511 ? add_955545 : sel_955542;
  assign add_955549 = sel_955546 + 8'h01;
  assign sel_955550 = array_index_955525 == array_index_948519 ? add_955549 : sel_955546;
  assign add_955553 = sel_955550 + 8'h01;
  assign sel_955554 = array_index_955525 == array_index_948527 ? add_955553 : sel_955550;
  assign add_955557 = sel_955554 + 8'h01;
  assign sel_955558 = array_index_955525 == array_index_948535 ? add_955557 : sel_955554;
  assign add_955561 = sel_955558 + 8'h01;
  assign sel_955562 = array_index_955525 == array_index_948541 ? add_955561 : sel_955558;
  assign add_955565 = sel_955562 + 8'h01;
  assign sel_955566 = array_index_955525 == array_index_948547 ? add_955565 : sel_955562;
  assign add_955569 = sel_955566 + 8'h01;
  assign sel_955570 = array_index_955525 == array_index_948553 ? add_955569 : sel_955566;
  assign add_955573 = sel_955570 + 8'h01;
  assign sel_955574 = array_index_955525 == array_index_948559 ? add_955573 : sel_955570;
  assign add_955577 = sel_955574 + 8'h01;
  assign sel_955578 = array_index_955525 == array_index_948565 ? add_955577 : sel_955574;
  assign add_955581 = sel_955578 + 8'h01;
  assign sel_955582 = array_index_955525 == array_index_948571 ? add_955581 : sel_955578;
  assign add_955585 = sel_955582 + 8'h01;
  assign sel_955586 = array_index_955525 == array_index_948577 ? add_955585 : sel_955582;
  assign add_955589 = sel_955586 + 8'h01;
  assign sel_955590 = array_index_955525 == array_index_948583 ? add_955589 : sel_955586;
  assign add_955593 = sel_955590 + 8'h01;
  assign sel_955594 = array_index_955525 == array_index_948589 ? add_955593 : sel_955590;
  assign add_955597 = sel_955594 + 8'h01;
  assign sel_955598 = array_index_955525 == array_index_948595 ? add_955597 : sel_955594;
  assign add_955601 = sel_955598 + 8'h01;
  assign sel_955602 = array_index_955525 == array_index_948601 ? add_955601 : sel_955598;
  assign add_955605 = sel_955602 + 8'h01;
  assign sel_955606 = array_index_955525 == array_index_948607 ? add_955605 : sel_955602;
  assign add_955609 = sel_955606 + 8'h01;
  assign sel_955610 = array_index_955525 == array_index_948613 ? add_955609 : sel_955606;
  assign add_955613 = sel_955610 + 8'h01;
  assign sel_955614 = array_index_955525 == array_index_948619 ? add_955613 : sel_955610;
  assign add_955617 = sel_955614 + 8'h01;
  assign sel_955618 = array_index_955525 == array_index_948625 ? add_955617 : sel_955614;
  assign add_955621 = sel_955618 + 8'h01;
  assign sel_955622 = array_index_955525 == array_index_948631 ? add_955621 : sel_955618;
  assign add_955625 = sel_955622 + 8'h01;
  assign sel_955626 = array_index_955525 == array_index_948637 ? add_955625 : sel_955622;
  assign add_955629 = sel_955626 + 8'h01;
  assign sel_955630 = array_index_955525 == array_index_948643 ? add_955629 : sel_955626;
  assign add_955633 = sel_955630 + 8'h01;
  assign sel_955634 = array_index_955525 == array_index_948649 ? add_955633 : sel_955630;
  assign add_955637 = sel_955634 + 8'h01;
  assign sel_955638 = array_index_955525 == array_index_948655 ? add_955637 : sel_955634;
  assign add_955641 = sel_955638 + 8'h01;
  assign sel_955642 = array_index_955525 == array_index_948661 ? add_955641 : sel_955638;
  assign add_955645 = sel_955642 + 8'h01;
  assign sel_955646 = array_index_955525 == array_index_948667 ? add_955645 : sel_955642;
  assign add_955649 = sel_955646 + 8'h01;
  assign sel_955650 = array_index_955525 == array_index_948673 ? add_955649 : sel_955646;
  assign add_955653 = sel_955650 + 8'h01;
  assign sel_955654 = array_index_955525 == array_index_948679 ? add_955653 : sel_955650;
  assign add_955657 = sel_955654 + 8'h01;
  assign sel_955658 = array_index_955525 == array_index_948685 ? add_955657 : sel_955654;
  assign add_955661 = sel_955658 + 8'h01;
  assign sel_955662 = array_index_955525 == array_index_948691 ? add_955661 : sel_955658;
  assign add_955665 = sel_955662 + 8'h01;
  assign sel_955666 = array_index_955525 == array_index_948697 ? add_955665 : sel_955662;
  assign add_955669 = sel_955666 + 8'h01;
  assign sel_955670 = array_index_955525 == array_index_948703 ? add_955669 : sel_955666;
  assign add_955673 = sel_955670 + 8'h01;
  assign sel_955674 = array_index_955525 == array_index_948709 ? add_955673 : sel_955670;
  assign add_955677 = sel_955674 + 8'h01;
  assign sel_955678 = array_index_955525 == array_index_948715 ? add_955677 : sel_955674;
  assign add_955681 = sel_955678 + 8'h01;
  assign sel_955682 = array_index_955525 == array_index_948721 ? add_955681 : sel_955678;
  assign add_955685 = sel_955682 + 8'h01;
  assign sel_955686 = array_index_955525 == array_index_948727 ? add_955685 : sel_955682;
  assign add_955689 = sel_955686 + 8'h01;
  assign sel_955690 = array_index_955525 == array_index_948733 ? add_955689 : sel_955686;
  assign add_955693 = sel_955690 + 8'h01;
  assign sel_955694 = array_index_955525 == array_index_948739 ? add_955693 : sel_955690;
  assign add_955697 = sel_955694 + 8'h01;
  assign sel_955698 = array_index_955525 == array_index_948745 ? add_955697 : sel_955694;
  assign add_955701 = sel_955698 + 8'h01;
  assign sel_955702 = array_index_955525 == array_index_948751 ? add_955701 : sel_955698;
  assign add_955705 = sel_955702 + 8'h01;
  assign sel_955706 = array_index_955525 == array_index_948757 ? add_955705 : sel_955702;
  assign add_955709 = sel_955706 + 8'h01;
  assign sel_955710 = array_index_955525 == array_index_948763 ? add_955709 : sel_955706;
  assign add_955713 = sel_955710 + 8'h01;
  assign sel_955714 = array_index_955525 == array_index_948769 ? add_955713 : sel_955710;
  assign add_955717 = sel_955714 + 8'h01;
  assign sel_955718 = array_index_955525 == array_index_948775 ? add_955717 : sel_955714;
  assign add_955721 = sel_955718 + 8'h01;
  assign sel_955722 = array_index_955525 == array_index_948781 ? add_955721 : sel_955718;
  assign add_955725 = sel_955722 + 8'h01;
  assign sel_955726 = array_index_955525 == array_index_948787 ? add_955725 : sel_955722;
  assign add_955729 = sel_955726 + 8'h01;
  assign sel_955730 = array_index_955525 == array_index_948793 ? add_955729 : sel_955726;
  assign add_955733 = sel_955730 + 8'h01;
  assign sel_955734 = array_index_955525 == array_index_948799 ? add_955733 : sel_955730;
  assign add_955737 = sel_955734 + 8'h01;
  assign sel_955738 = array_index_955525 == array_index_948805 ? add_955737 : sel_955734;
  assign add_955741 = sel_955738 + 8'h01;
  assign sel_955742 = array_index_955525 == array_index_948811 ? add_955741 : sel_955738;
  assign add_955745 = sel_955742 + 8'h01;
  assign sel_955746 = array_index_955525 == array_index_948817 ? add_955745 : sel_955742;
  assign add_955749 = sel_955746 + 8'h01;
  assign sel_955750 = array_index_955525 == array_index_948823 ? add_955749 : sel_955746;
  assign add_955753 = sel_955750 + 8'h01;
  assign sel_955754 = array_index_955525 == array_index_948829 ? add_955753 : sel_955750;
  assign add_955757 = sel_955754 + 8'h01;
  assign sel_955758 = array_index_955525 == array_index_948835 ? add_955757 : sel_955754;
  assign add_955761 = sel_955758 + 8'h01;
  assign sel_955762 = array_index_955525 == array_index_948841 ? add_955761 : sel_955758;
  assign add_955765 = sel_955762 + 8'h01;
  assign sel_955766 = array_index_955525 == array_index_948847 ? add_955765 : sel_955762;
  assign add_955769 = sel_955766 + 8'h01;
  assign sel_955770 = array_index_955525 == array_index_948853 ? add_955769 : sel_955766;
  assign add_955773 = sel_955770 + 8'h01;
  assign sel_955774 = array_index_955525 == array_index_948859 ? add_955773 : sel_955770;
  assign add_955777 = sel_955774 + 8'h01;
  assign sel_955778 = array_index_955525 == array_index_948865 ? add_955777 : sel_955774;
  assign add_955781 = sel_955778 + 8'h01;
  assign sel_955782 = array_index_955525 == array_index_948871 ? add_955781 : sel_955778;
  assign add_955785 = sel_955782 + 8'h01;
  assign sel_955786 = array_index_955525 == array_index_948877 ? add_955785 : sel_955782;
  assign add_955789 = sel_955786 + 8'h01;
  assign sel_955790 = array_index_955525 == array_index_948883 ? add_955789 : sel_955786;
  assign add_955793 = sel_955790 + 8'h01;
  assign sel_955794 = array_index_955525 == array_index_948889 ? add_955793 : sel_955790;
  assign add_955797 = sel_955794 + 8'h01;
  assign sel_955798 = array_index_955525 == array_index_948895 ? add_955797 : sel_955794;
  assign add_955801 = sel_955798 + 8'h01;
  assign sel_955802 = array_index_955525 == array_index_948901 ? add_955801 : sel_955798;
  assign add_955805 = sel_955802 + 8'h01;
  assign sel_955806 = array_index_955525 == array_index_948907 ? add_955805 : sel_955802;
  assign add_955809 = sel_955806 + 8'h01;
  assign sel_955810 = array_index_955525 == array_index_948913 ? add_955809 : sel_955806;
  assign add_955813 = sel_955810 + 8'h01;
  assign sel_955814 = array_index_955525 == array_index_948919 ? add_955813 : sel_955810;
  assign add_955817 = sel_955814 + 8'h01;
  assign sel_955818 = array_index_955525 == array_index_948925 ? add_955817 : sel_955814;
  assign add_955821 = sel_955818 + 8'h01;
  assign sel_955822 = array_index_955525 == array_index_948931 ? add_955821 : sel_955818;
  assign add_955825 = sel_955822 + 8'h01;
  assign sel_955826 = array_index_955525 == array_index_948937 ? add_955825 : sel_955822;
  assign add_955829 = sel_955826 + 8'h01;
  assign sel_955830 = array_index_955525 == array_index_948943 ? add_955829 : sel_955826;
  assign add_955833 = sel_955830 + 8'h01;
  assign sel_955834 = array_index_955525 == array_index_948949 ? add_955833 : sel_955830;
  assign add_955837 = sel_955834 + 8'h01;
  assign sel_955838 = array_index_955525 == array_index_948955 ? add_955837 : sel_955834;
  assign add_955841 = sel_955838 + 8'h01;
  assign sel_955842 = array_index_955525 == array_index_948961 ? add_955841 : sel_955838;
  assign add_955845 = sel_955842 + 8'h01;
  assign sel_955846 = array_index_955525 == array_index_948967 ? add_955845 : sel_955842;
  assign add_955849 = sel_955846 + 8'h01;
  assign sel_955850 = array_index_955525 == array_index_948973 ? add_955849 : sel_955846;
  assign add_955853 = sel_955850 + 8'h01;
  assign sel_955854 = array_index_955525 == array_index_948979 ? add_955853 : sel_955850;
  assign add_955857 = sel_955854 + 8'h01;
  assign sel_955858 = array_index_955525 == array_index_948985 ? add_955857 : sel_955854;
  assign add_955861 = sel_955858 + 8'h01;
  assign sel_955862 = array_index_955525 == array_index_948991 ? add_955861 : sel_955858;
  assign add_955865 = sel_955862 + 8'h01;
  assign sel_955866 = array_index_955525 == array_index_948997 ? add_955865 : sel_955862;
  assign add_955869 = sel_955866 + 8'h01;
  assign sel_955870 = array_index_955525 == array_index_949003 ? add_955869 : sel_955866;
  assign add_955873 = sel_955870 + 8'h01;
  assign sel_955874 = array_index_955525 == array_index_949009 ? add_955873 : sel_955870;
  assign add_955877 = sel_955874 + 8'h01;
  assign sel_955878 = array_index_955525 == array_index_949015 ? add_955877 : sel_955874;
  assign add_955881 = sel_955878 + 8'h01;
  assign sel_955882 = array_index_955525 == array_index_949021 ? add_955881 : sel_955878;
  assign add_955885 = sel_955882 + 8'h01;
  assign sel_955886 = array_index_955525 == array_index_949027 ? add_955885 : sel_955882;
  assign add_955889 = sel_955886 + 8'h01;
  assign sel_955890 = array_index_955525 == array_index_949033 ? add_955889 : sel_955886;
  assign add_955893 = sel_955890 + 8'h01;
  assign sel_955894 = array_index_955525 == array_index_949039 ? add_955893 : sel_955890;
  assign add_955897 = sel_955894 + 8'h01;
  assign sel_955898 = array_index_955525 == array_index_949045 ? add_955897 : sel_955894;
  assign add_955901 = sel_955898 + 8'h01;
  assign sel_955902 = array_index_955525 == array_index_949051 ? add_955901 : sel_955898;
  assign add_955905 = sel_955902 + 8'h01;
  assign sel_955906 = array_index_955525 == array_index_949057 ? add_955905 : sel_955902;
  assign add_955909 = sel_955906 + 8'h01;
  assign sel_955910 = array_index_955525 == array_index_949063 ? add_955909 : sel_955906;
  assign add_955913 = sel_955910 + 8'h01;
  assign sel_955914 = array_index_955525 == array_index_949069 ? add_955913 : sel_955910;
  assign add_955917 = sel_955914 + 8'h01;
  assign sel_955918 = array_index_955525 == array_index_949075 ? add_955917 : sel_955914;
  assign add_955921 = sel_955918 + 8'h01;
  assign sel_955922 = array_index_955525 == array_index_949081 ? add_955921 : sel_955918;
  assign add_955926 = sel_955922 + 8'h01;
  assign array_index_955927 = set1_unflattened[7'h12];
  assign sel_955928 = array_index_955525 == array_index_949087 ? add_955926 : sel_955922;
  assign add_955931 = sel_955928 + 8'h01;
  assign sel_955932 = array_index_955927 == array_index_948483 ? add_955931 : sel_955928;
  assign add_955935 = sel_955932 + 8'h01;
  assign sel_955936 = array_index_955927 == array_index_948487 ? add_955935 : sel_955932;
  assign add_955939 = sel_955936 + 8'h01;
  assign sel_955940 = array_index_955927 == array_index_948495 ? add_955939 : sel_955936;
  assign add_955943 = sel_955940 + 8'h01;
  assign sel_955944 = array_index_955927 == array_index_948503 ? add_955943 : sel_955940;
  assign add_955947 = sel_955944 + 8'h01;
  assign sel_955948 = array_index_955927 == array_index_948511 ? add_955947 : sel_955944;
  assign add_955951 = sel_955948 + 8'h01;
  assign sel_955952 = array_index_955927 == array_index_948519 ? add_955951 : sel_955948;
  assign add_955955 = sel_955952 + 8'h01;
  assign sel_955956 = array_index_955927 == array_index_948527 ? add_955955 : sel_955952;
  assign add_955959 = sel_955956 + 8'h01;
  assign sel_955960 = array_index_955927 == array_index_948535 ? add_955959 : sel_955956;
  assign add_955963 = sel_955960 + 8'h01;
  assign sel_955964 = array_index_955927 == array_index_948541 ? add_955963 : sel_955960;
  assign add_955967 = sel_955964 + 8'h01;
  assign sel_955968 = array_index_955927 == array_index_948547 ? add_955967 : sel_955964;
  assign add_955971 = sel_955968 + 8'h01;
  assign sel_955972 = array_index_955927 == array_index_948553 ? add_955971 : sel_955968;
  assign add_955975 = sel_955972 + 8'h01;
  assign sel_955976 = array_index_955927 == array_index_948559 ? add_955975 : sel_955972;
  assign add_955979 = sel_955976 + 8'h01;
  assign sel_955980 = array_index_955927 == array_index_948565 ? add_955979 : sel_955976;
  assign add_955983 = sel_955980 + 8'h01;
  assign sel_955984 = array_index_955927 == array_index_948571 ? add_955983 : sel_955980;
  assign add_955987 = sel_955984 + 8'h01;
  assign sel_955988 = array_index_955927 == array_index_948577 ? add_955987 : sel_955984;
  assign add_955991 = sel_955988 + 8'h01;
  assign sel_955992 = array_index_955927 == array_index_948583 ? add_955991 : sel_955988;
  assign add_955995 = sel_955992 + 8'h01;
  assign sel_955996 = array_index_955927 == array_index_948589 ? add_955995 : sel_955992;
  assign add_955999 = sel_955996 + 8'h01;
  assign sel_956000 = array_index_955927 == array_index_948595 ? add_955999 : sel_955996;
  assign add_956003 = sel_956000 + 8'h01;
  assign sel_956004 = array_index_955927 == array_index_948601 ? add_956003 : sel_956000;
  assign add_956007 = sel_956004 + 8'h01;
  assign sel_956008 = array_index_955927 == array_index_948607 ? add_956007 : sel_956004;
  assign add_956011 = sel_956008 + 8'h01;
  assign sel_956012 = array_index_955927 == array_index_948613 ? add_956011 : sel_956008;
  assign add_956015 = sel_956012 + 8'h01;
  assign sel_956016 = array_index_955927 == array_index_948619 ? add_956015 : sel_956012;
  assign add_956019 = sel_956016 + 8'h01;
  assign sel_956020 = array_index_955927 == array_index_948625 ? add_956019 : sel_956016;
  assign add_956023 = sel_956020 + 8'h01;
  assign sel_956024 = array_index_955927 == array_index_948631 ? add_956023 : sel_956020;
  assign add_956027 = sel_956024 + 8'h01;
  assign sel_956028 = array_index_955927 == array_index_948637 ? add_956027 : sel_956024;
  assign add_956031 = sel_956028 + 8'h01;
  assign sel_956032 = array_index_955927 == array_index_948643 ? add_956031 : sel_956028;
  assign add_956035 = sel_956032 + 8'h01;
  assign sel_956036 = array_index_955927 == array_index_948649 ? add_956035 : sel_956032;
  assign add_956039 = sel_956036 + 8'h01;
  assign sel_956040 = array_index_955927 == array_index_948655 ? add_956039 : sel_956036;
  assign add_956043 = sel_956040 + 8'h01;
  assign sel_956044 = array_index_955927 == array_index_948661 ? add_956043 : sel_956040;
  assign add_956047 = sel_956044 + 8'h01;
  assign sel_956048 = array_index_955927 == array_index_948667 ? add_956047 : sel_956044;
  assign add_956051 = sel_956048 + 8'h01;
  assign sel_956052 = array_index_955927 == array_index_948673 ? add_956051 : sel_956048;
  assign add_956055 = sel_956052 + 8'h01;
  assign sel_956056 = array_index_955927 == array_index_948679 ? add_956055 : sel_956052;
  assign add_956059 = sel_956056 + 8'h01;
  assign sel_956060 = array_index_955927 == array_index_948685 ? add_956059 : sel_956056;
  assign add_956063 = sel_956060 + 8'h01;
  assign sel_956064 = array_index_955927 == array_index_948691 ? add_956063 : sel_956060;
  assign add_956067 = sel_956064 + 8'h01;
  assign sel_956068 = array_index_955927 == array_index_948697 ? add_956067 : sel_956064;
  assign add_956071 = sel_956068 + 8'h01;
  assign sel_956072 = array_index_955927 == array_index_948703 ? add_956071 : sel_956068;
  assign add_956075 = sel_956072 + 8'h01;
  assign sel_956076 = array_index_955927 == array_index_948709 ? add_956075 : sel_956072;
  assign add_956079 = sel_956076 + 8'h01;
  assign sel_956080 = array_index_955927 == array_index_948715 ? add_956079 : sel_956076;
  assign add_956083 = sel_956080 + 8'h01;
  assign sel_956084 = array_index_955927 == array_index_948721 ? add_956083 : sel_956080;
  assign add_956087 = sel_956084 + 8'h01;
  assign sel_956088 = array_index_955927 == array_index_948727 ? add_956087 : sel_956084;
  assign add_956091 = sel_956088 + 8'h01;
  assign sel_956092 = array_index_955927 == array_index_948733 ? add_956091 : sel_956088;
  assign add_956095 = sel_956092 + 8'h01;
  assign sel_956096 = array_index_955927 == array_index_948739 ? add_956095 : sel_956092;
  assign add_956099 = sel_956096 + 8'h01;
  assign sel_956100 = array_index_955927 == array_index_948745 ? add_956099 : sel_956096;
  assign add_956103 = sel_956100 + 8'h01;
  assign sel_956104 = array_index_955927 == array_index_948751 ? add_956103 : sel_956100;
  assign add_956107 = sel_956104 + 8'h01;
  assign sel_956108 = array_index_955927 == array_index_948757 ? add_956107 : sel_956104;
  assign add_956111 = sel_956108 + 8'h01;
  assign sel_956112 = array_index_955927 == array_index_948763 ? add_956111 : sel_956108;
  assign add_956115 = sel_956112 + 8'h01;
  assign sel_956116 = array_index_955927 == array_index_948769 ? add_956115 : sel_956112;
  assign add_956119 = sel_956116 + 8'h01;
  assign sel_956120 = array_index_955927 == array_index_948775 ? add_956119 : sel_956116;
  assign add_956123 = sel_956120 + 8'h01;
  assign sel_956124 = array_index_955927 == array_index_948781 ? add_956123 : sel_956120;
  assign add_956127 = sel_956124 + 8'h01;
  assign sel_956128 = array_index_955927 == array_index_948787 ? add_956127 : sel_956124;
  assign add_956131 = sel_956128 + 8'h01;
  assign sel_956132 = array_index_955927 == array_index_948793 ? add_956131 : sel_956128;
  assign add_956135 = sel_956132 + 8'h01;
  assign sel_956136 = array_index_955927 == array_index_948799 ? add_956135 : sel_956132;
  assign add_956139 = sel_956136 + 8'h01;
  assign sel_956140 = array_index_955927 == array_index_948805 ? add_956139 : sel_956136;
  assign add_956143 = sel_956140 + 8'h01;
  assign sel_956144 = array_index_955927 == array_index_948811 ? add_956143 : sel_956140;
  assign add_956147 = sel_956144 + 8'h01;
  assign sel_956148 = array_index_955927 == array_index_948817 ? add_956147 : sel_956144;
  assign add_956151 = sel_956148 + 8'h01;
  assign sel_956152 = array_index_955927 == array_index_948823 ? add_956151 : sel_956148;
  assign add_956155 = sel_956152 + 8'h01;
  assign sel_956156 = array_index_955927 == array_index_948829 ? add_956155 : sel_956152;
  assign add_956159 = sel_956156 + 8'h01;
  assign sel_956160 = array_index_955927 == array_index_948835 ? add_956159 : sel_956156;
  assign add_956163 = sel_956160 + 8'h01;
  assign sel_956164 = array_index_955927 == array_index_948841 ? add_956163 : sel_956160;
  assign add_956167 = sel_956164 + 8'h01;
  assign sel_956168 = array_index_955927 == array_index_948847 ? add_956167 : sel_956164;
  assign add_956171 = sel_956168 + 8'h01;
  assign sel_956172 = array_index_955927 == array_index_948853 ? add_956171 : sel_956168;
  assign add_956175 = sel_956172 + 8'h01;
  assign sel_956176 = array_index_955927 == array_index_948859 ? add_956175 : sel_956172;
  assign add_956179 = sel_956176 + 8'h01;
  assign sel_956180 = array_index_955927 == array_index_948865 ? add_956179 : sel_956176;
  assign add_956183 = sel_956180 + 8'h01;
  assign sel_956184 = array_index_955927 == array_index_948871 ? add_956183 : sel_956180;
  assign add_956187 = sel_956184 + 8'h01;
  assign sel_956188 = array_index_955927 == array_index_948877 ? add_956187 : sel_956184;
  assign add_956191 = sel_956188 + 8'h01;
  assign sel_956192 = array_index_955927 == array_index_948883 ? add_956191 : sel_956188;
  assign add_956195 = sel_956192 + 8'h01;
  assign sel_956196 = array_index_955927 == array_index_948889 ? add_956195 : sel_956192;
  assign add_956199 = sel_956196 + 8'h01;
  assign sel_956200 = array_index_955927 == array_index_948895 ? add_956199 : sel_956196;
  assign add_956203 = sel_956200 + 8'h01;
  assign sel_956204 = array_index_955927 == array_index_948901 ? add_956203 : sel_956200;
  assign add_956207 = sel_956204 + 8'h01;
  assign sel_956208 = array_index_955927 == array_index_948907 ? add_956207 : sel_956204;
  assign add_956211 = sel_956208 + 8'h01;
  assign sel_956212 = array_index_955927 == array_index_948913 ? add_956211 : sel_956208;
  assign add_956215 = sel_956212 + 8'h01;
  assign sel_956216 = array_index_955927 == array_index_948919 ? add_956215 : sel_956212;
  assign add_956219 = sel_956216 + 8'h01;
  assign sel_956220 = array_index_955927 == array_index_948925 ? add_956219 : sel_956216;
  assign add_956223 = sel_956220 + 8'h01;
  assign sel_956224 = array_index_955927 == array_index_948931 ? add_956223 : sel_956220;
  assign add_956227 = sel_956224 + 8'h01;
  assign sel_956228 = array_index_955927 == array_index_948937 ? add_956227 : sel_956224;
  assign add_956231 = sel_956228 + 8'h01;
  assign sel_956232 = array_index_955927 == array_index_948943 ? add_956231 : sel_956228;
  assign add_956235 = sel_956232 + 8'h01;
  assign sel_956236 = array_index_955927 == array_index_948949 ? add_956235 : sel_956232;
  assign add_956239 = sel_956236 + 8'h01;
  assign sel_956240 = array_index_955927 == array_index_948955 ? add_956239 : sel_956236;
  assign add_956243 = sel_956240 + 8'h01;
  assign sel_956244 = array_index_955927 == array_index_948961 ? add_956243 : sel_956240;
  assign add_956247 = sel_956244 + 8'h01;
  assign sel_956248 = array_index_955927 == array_index_948967 ? add_956247 : sel_956244;
  assign add_956251 = sel_956248 + 8'h01;
  assign sel_956252 = array_index_955927 == array_index_948973 ? add_956251 : sel_956248;
  assign add_956255 = sel_956252 + 8'h01;
  assign sel_956256 = array_index_955927 == array_index_948979 ? add_956255 : sel_956252;
  assign add_956259 = sel_956256 + 8'h01;
  assign sel_956260 = array_index_955927 == array_index_948985 ? add_956259 : sel_956256;
  assign add_956263 = sel_956260 + 8'h01;
  assign sel_956264 = array_index_955927 == array_index_948991 ? add_956263 : sel_956260;
  assign add_956267 = sel_956264 + 8'h01;
  assign sel_956268 = array_index_955927 == array_index_948997 ? add_956267 : sel_956264;
  assign add_956271 = sel_956268 + 8'h01;
  assign sel_956272 = array_index_955927 == array_index_949003 ? add_956271 : sel_956268;
  assign add_956275 = sel_956272 + 8'h01;
  assign sel_956276 = array_index_955927 == array_index_949009 ? add_956275 : sel_956272;
  assign add_956279 = sel_956276 + 8'h01;
  assign sel_956280 = array_index_955927 == array_index_949015 ? add_956279 : sel_956276;
  assign add_956283 = sel_956280 + 8'h01;
  assign sel_956284 = array_index_955927 == array_index_949021 ? add_956283 : sel_956280;
  assign add_956287 = sel_956284 + 8'h01;
  assign sel_956288 = array_index_955927 == array_index_949027 ? add_956287 : sel_956284;
  assign add_956291 = sel_956288 + 8'h01;
  assign sel_956292 = array_index_955927 == array_index_949033 ? add_956291 : sel_956288;
  assign add_956295 = sel_956292 + 8'h01;
  assign sel_956296 = array_index_955927 == array_index_949039 ? add_956295 : sel_956292;
  assign add_956299 = sel_956296 + 8'h01;
  assign sel_956300 = array_index_955927 == array_index_949045 ? add_956299 : sel_956296;
  assign add_956303 = sel_956300 + 8'h01;
  assign sel_956304 = array_index_955927 == array_index_949051 ? add_956303 : sel_956300;
  assign add_956307 = sel_956304 + 8'h01;
  assign sel_956308 = array_index_955927 == array_index_949057 ? add_956307 : sel_956304;
  assign add_956311 = sel_956308 + 8'h01;
  assign sel_956312 = array_index_955927 == array_index_949063 ? add_956311 : sel_956308;
  assign add_956315 = sel_956312 + 8'h01;
  assign sel_956316 = array_index_955927 == array_index_949069 ? add_956315 : sel_956312;
  assign add_956319 = sel_956316 + 8'h01;
  assign sel_956320 = array_index_955927 == array_index_949075 ? add_956319 : sel_956316;
  assign add_956323 = sel_956320 + 8'h01;
  assign sel_956324 = array_index_955927 == array_index_949081 ? add_956323 : sel_956320;
  assign add_956328 = sel_956324 + 8'h01;
  assign array_index_956329 = set1_unflattened[7'h13];
  assign sel_956330 = array_index_955927 == array_index_949087 ? add_956328 : sel_956324;
  assign add_956333 = sel_956330 + 8'h01;
  assign sel_956334 = array_index_956329 == array_index_948483 ? add_956333 : sel_956330;
  assign add_956337 = sel_956334 + 8'h01;
  assign sel_956338 = array_index_956329 == array_index_948487 ? add_956337 : sel_956334;
  assign add_956341 = sel_956338 + 8'h01;
  assign sel_956342 = array_index_956329 == array_index_948495 ? add_956341 : sel_956338;
  assign add_956345 = sel_956342 + 8'h01;
  assign sel_956346 = array_index_956329 == array_index_948503 ? add_956345 : sel_956342;
  assign add_956349 = sel_956346 + 8'h01;
  assign sel_956350 = array_index_956329 == array_index_948511 ? add_956349 : sel_956346;
  assign add_956353 = sel_956350 + 8'h01;
  assign sel_956354 = array_index_956329 == array_index_948519 ? add_956353 : sel_956350;
  assign add_956357 = sel_956354 + 8'h01;
  assign sel_956358 = array_index_956329 == array_index_948527 ? add_956357 : sel_956354;
  assign add_956361 = sel_956358 + 8'h01;
  assign sel_956362 = array_index_956329 == array_index_948535 ? add_956361 : sel_956358;
  assign add_956365 = sel_956362 + 8'h01;
  assign sel_956366 = array_index_956329 == array_index_948541 ? add_956365 : sel_956362;
  assign add_956369 = sel_956366 + 8'h01;
  assign sel_956370 = array_index_956329 == array_index_948547 ? add_956369 : sel_956366;
  assign add_956373 = sel_956370 + 8'h01;
  assign sel_956374 = array_index_956329 == array_index_948553 ? add_956373 : sel_956370;
  assign add_956377 = sel_956374 + 8'h01;
  assign sel_956378 = array_index_956329 == array_index_948559 ? add_956377 : sel_956374;
  assign add_956381 = sel_956378 + 8'h01;
  assign sel_956382 = array_index_956329 == array_index_948565 ? add_956381 : sel_956378;
  assign add_956385 = sel_956382 + 8'h01;
  assign sel_956386 = array_index_956329 == array_index_948571 ? add_956385 : sel_956382;
  assign add_956389 = sel_956386 + 8'h01;
  assign sel_956390 = array_index_956329 == array_index_948577 ? add_956389 : sel_956386;
  assign add_956393 = sel_956390 + 8'h01;
  assign sel_956394 = array_index_956329 == array_index_948583 ? add_956393 : sel_956390;
  assign add_956397 = sel_956394 + 8'h01;
  assign sel_956398 = array_index_956329 == array_index_948589 ? add_956397 : sel_956394;
  assign add_956401 = sel_956398 + 8'h01;
  assign sel_956402 = array_index_956329 == array_index_948595 ? add_956401 : sel_956398;
  assign add_956405 = sel_956402 + 8'h01;
  assign sel_956406 = array_index_956329 == array_index_948601 ? add_956405 : sel_956402;
  assign add_956409 = sel_956406 + 8'h01;
  assign sel_956410 = array_index_956329 == array_index_948607 ? add_956409 : sel_956406;
  assign add_956413 = sel_956410 + 8'h01;
  assign sel_956414 = array_index_956329 == array_index_948613 ? add_956413 : sel_956410;
  assign add_956417 = sel_956414 + 8'h01;
  assign sel_956418 = array_index_956329 == array_index_948619 ? add_956417 : sel_956414;
  assign add_956421 = sel_956418 + 8'h01;
  assign sel_956422 = array_index_956329 == array_index_948625 ? add_956421 : sel_956418;
  assign add_956425 = sel_956422 + 8'h01;
  assign sel_956426 = array_index_956329 == array_index_948631 ? add_956425 : sel_956422;
  assign add_956429 = sel_956426 + 8'h01;
  assign sel_956430 = array_index_956329 == array_index_948637 ? add_956429 : sel_956426;
  assign add_956433 = sel_956430 + 8'h01;
  assign sel_956434 = array_index_956329 == array_index_948643 ? add_956433 : sel_956430;
  assign add_956437 = sel_956434 + 8'h01;
  assign sel_956438 = array_index_956329 == array_index_948649 ? add_956437 : sel_956434;
  assign add_956441 = sel_956438 + 8'h01;
  assign sel_956442 = array_index_956329 == array_index_948655 ? add_956441 : sel_956438;
  assign add_956445 = sel_956442 + 8'h01;
  assign sel_956446 = array_index_956329 == array_index_948661 ? add_956445 : sel_956442;
  assign add_956449 = sel_956446 + 8'h01;
  assign sel_956450 = array_index_956329 == array_index_948667 ? add_956449 : sel_956446;
  assign add_956453 = sel_956450 + 8'h01;
  assign sel_956454 = array_index_956329 == array_index_948673 ? add_956453 : sel_956450;
  assign add_956457 = sel_956454 + 8'h01;
  assign sel_956458 = array_index_956329 == array_index_948679 ? add_956457 : sel_956454;
  assign add_956461 = sel_956458 + 8'h01;
  assign sel_956462 = array_index_956329 == array_index_948685 ? add_956461 : sel_956458;
  assign add_956465 = sel_956462 + 8'h01;
  assign sel_956466 = array_index_956329 == array_index_948691 ? add_956465 : sel_956462;
  assign add_956469 = sel_956466 + 8'h01;
  assign sel_956470 = array_index_956329 == array_index_948697 ? add_956469 : sel_956466;
  assign add_956473 = sel_956470 + 8'h01;
  assign sel_956474 = array_index_956329 == array_index_948703 ? add_956473 : sel_956470;
  assign add_956477 = sel_956474 + 8'h01;
  assign sel_956478 = array_index_956329 == array_index_948709 ? add_956477 : sel_956474;
  assign add_956481 = sel_956478 + 8'h01;
  assign sel_956482 = array_index_956329 == array_index_948715 ? add_956481 : sel_956478;
  assign add_956485 = sel_956482 + 8'h01;
  assign sel_956486 = array_index_956329 == array_index_948721 ? add_956485 : sel_956482;
  assign add_956489 = sel_956486 + 8'h01;
  assign sel_956490 = array_index_956329 == array_index_948727 ? add_956489 : sel_956486;
  assign add_956493 = sel_956490 + 8'h01;
  assign sel_956494 = array_index_956329 == array_index_948733 ? add_956493 : sel_956490;
  assign add_956497 = sel_956494 + 8'h01;
  assign sel_956498 = array_index_956329 == array_index_948739 ? add_956497 : sel_956494;
  assign add_956501 = sel_956498 + 8'h01;
  assign sel_956502 = array_index_956329 == array_index_948745 ? add_956501 : sel_956498;
  assign add_956505 = sel_956502 + 8'h01;
  assign sel_956506 = array_index_956329 == array_index_948751 ? add_956505 : sel_956502;
  assign add_956509 = sel_956506 + 8'h01;
  assign sel_956510 = array_index_956329 == array_index_948757 ? add_956509 : sel_956506;
  assign add_956513 = sel_956510 + 8'h01;
  assign sel_956514 = array_index_956329 == array_index_948763 ? add_956513 : sel_956510;
  assign add_956517 = sel_956514 + 8'h01;
  assign sel_956518 = array_index_956329 == array_index_948769 ? add_956517 : sel_956514;
  assign add_956521 = sel_956518 + 8'h01;
  assign sel_956522 = array_index_956329 == array_index_948775 ? add_956521 : sel_956518;
  assign add_956525 = sel_956522 + 8'h01;
  assign sel_956526 = array_index_956329 == array_index_948781 ? add_956525 : sel_956522;
  assign add_956529 = sel_956526 + 8'h01;
  assign sel_956530 = array_index_956329 == array_index_948787 ? add_956529 : sel_956526;
  assign add_956533 = sel_956530 + 8'h01;
  assign sel_956534 = array_index_956329 == array_index_948793 ? add_956533 : sel_956530;
  assign add_956537 = sel_956534 + 8'h01;
  assign sel_956538 = array_index_956329 == array_index_948799 ? add_956537 : sel_956534;
  assign add_956541 = sel_956538 + 8'h01;
  assign sel_956542 = array_index_956329 == array_index_948805 ? add_956541 : sel_956538;
  assign add_956545 = sel_956542 + 8'h01;
  assign sel_956546 = array_index_956329 == array_index_948811 ? add_956545 : sel_956542;
  assign add_956549 = sel_956546 + 8'h01;
  assign sel_956550 = array_index_956329 == array_index_948817 ? add_956549 : sel_956546;
  assign add_956553 = sel_956550 + 8'h01;
  assign sel_956554 = array_index_956329 == array_index_948823 ? add_956553 : sel_956550;
  assign add_956557 = sel_956554 + 8'h01;
  assign sel_956558 = array_index_956329 == array_index_948829 ? add_956557 : sel_956554;
  assign add_956561 = sel_956558 + 8'h01;
  assign sel_956562 = array_index_956329 == array_index_948835 ? add_956561 : sel_956558;
  assign add_956565 = sel_956562 + 8'h01;
  assign sel_956566 = array_index_956329 == array_index_948841 ? add_956565 : sel_956562;
  assign add_956569 = sel_956566 + 8'h01;
  assign sel_956570 = array_index_956329 == array_index_948847 ? add_956569 : sel_956566;
  assign add_956573 = sel_956570 + 8'h01;
  assign sel_956574 = array_index_956329 == array_index_948853 ? add_956573 : sel_956570;
  assign add_956577 = sel_956574 + 8'h01;
  assign sel_956578 = array_index_956329 == array_index_948859 ? add_956577 : sel_956574;
  assign add_956581 = sel_956578 + 8'h01;
  assign sel_956582 = array_index_956329 == array_index_948865 ? add_956581 : sel_956578;
  assign add_956585 = sel_956582 + 8'h01;
  assign sel_956586 = array_index_956329 == array_index_948871 ? add_956585 : sel_956582;
  assign add_956589 = sel_956586 + 8'h01;
  assign sel_956590 = array_index_956329 == array_index_948877 ? add_956589 : sel_956586;
  assign add_956593 = sel_956590 + 8'h01;
  assign sel_956594 = array_index_956329 == array_index_948883 ? add_956593 : sel_956590;
  assign add_956597 = sel_956594 + 8'h01;
  assign sel_956598 = array_index_956329 == array_index_948889 ? add_956597 : sel_956594;
  assign add_956601 = sel_956598 + 8'h01;
  assign sel_956602 = array_index_956329 == array_index_948895 ? add_956601 : sel_956598;
  assign add_956605 = sel_956602 + 8'h01;
  assign sel_956606 = array_index_956329 == array_index_948901 ? add_956605 : sel_956602;
  assign add_956609 = sel_956606 + 8'h01;
  assign sel_956610 = array_index_956329 == array_index_948907 ? add_956609 : sel_956606;
  assign add_956613 = sel_956610 + 8'h01;
  assign sel_956614 = array_index_956329 == array_index_948913 ? add_956613 : sel_956610;
  assign add_956617 = sel_956614 + 8'h01;
  assign sel_956618 = array_index_956329 == array_index_948919 ? add_956617 : sel_956614;
  assign add_956621 = sel_956618 + 8'h01;
  assign sel_956622 = array_index_956329 == array_index_948925 ? add_956621 : sel_956618;
  assign add_956625 = sel_956622 + 8'h01;
  assign sel_956626 = array_index_956329 == array_index_948931 ? add_956625 : sel_956622;
  assign add_956629 = sel_956626 + 8'h01;
  assign sel_956630 = array_index_956329 == array_index_948937 ? add_956629 : sel_956626;
  assign add_956633 = sel_956630 + 8'h01;
  assign sel_956634 = array_index_956329 == array_index_948943 ? add_956633 : sel_956630;
  assign add_956637 = sel_956634 + 8'h01;
  assign sel_956638 = array_index_956329 == array_index_948949 ? add_956637 : sel_956634;
  assign add_956641 = sel_956638 + 8'h01;
  assign sel_956642 = array_index_956329 == array_index_948955 ? add_956641 : sel_956638;
  assign add_956645 = sel_956642 + 8'h01;
  assign sel_956646 = array_index_956329 == array_index_948961 ? add_956645 : sel_956642;
  assign add_956649 = sel_956646 + 8'h01;
  assign sel_956650 = array_index_956329 == array_index_948967 ? add_956649 : sel_956646;
  assign add_956653 = sel_956650 + 8'h01;
  assign sel_956654 = array_index_956329 == array_index_948973 ? add_956653 : sel_956650;
  assign add_956657 = sel_956654 + 8'h01;
  assign sel_956658 = array_index_956329 == array_index_948979 ? add_956657 : sel_956654;
  assign add_956661 = sel_956658 + 8'h01;
  assign sel_956662 = array_index_956329 == array_index_948985 ? add_956661 : sel_956658;
  assign add_956665 = sel_956662 + 8'h01;
  assign sel_956666 = array_index_956329 == array_index_948991 ? add_956665 : sel_956662;
  assign add_956669 = sel_956666 + 8'h01;
  assign sel_956670 = array_index_956329 == array_index_948997 ? add_956669 : sel_956666;
  assign add_956673 = sel_956670 + 8'h01;
  assign sel_956674 = array_index_956329 == array_index_949003 ? add_956673 : sel_956670;
  assign add_956677 = sel_956674 + 8'h01;
  assign sel_956678 = array_index_956329 == array_index_949009 ? add_956677 : sel_956674;
  assign add_956681 = sel_956678 + 8'h01;
  assign sel_956682 = array_index_956329 == array_index_949015 ? add_956681 : sel_956678;
  assign add_956685 = sel_956682 + 8'h01;
  assign sel_956686 = array_index_956329 == array_index_949021 ? add_956685 : sel_956682;
  assign add_956689 = sel_956686 + 8'h01;
  assign sel_956690 = array_index_956329 == array_index_949027 ? add_956689 : sel_956686;
  assign add_956693 = sel_956690 + 8'h01;
  assign sel_956694 = array_index_956329 == array_index_949033 ? add_956693 : sel_956690;
  assign add_956697 = sel_956694 + 8'h01;
  assign sel_956698 = array_index_956329 == array_index_949039 ? add_956697 : sel_956694;
  assign add_956701 = sel_956698 + 8'h01;
  assign sel_956702 = array_index_956329 == array_index_949045 ? add_956701 : sel_956698;
  assign add_956705 = sel_956702 + 8'h01;
  assign sel_956706 = array_index_956329 == array_index_949051 ? add_956705 : sel_956702;
  assign add_956709 = sel_956706 + 8'h01;
  assign sel_956710 = array_index_956329 == array_index_949057 ? add_956709 : sel_956706;
  assign add_956713 = sel_956710 + 8'h01;
  assign sel_956714 = array_index_956329 == array_index_949063 ? add_956713 : sel_956710;
  assign add_956717 = sel_956714 + 8'h01;
  assign sel_956718 = array_index_956329 == array_index_949069 ? add_956717 : sel_956714;
  assign add_956721 = sel_956718 + 8'h01;
  assign sel_956722 = array_index_956329 == array_index_949075 ? add_956721 : sel_956718;
  assign add_956725 = sel_956722 + 8'h01;
  assign sel_956726 = array_index_956329 == array_index_949081 ? add_956725 : sel_956722;
  assign add_956730 = sel_956726 + 8'h01;
  assign array_index_956731 = set1_unflattened[7'h14];
  assign sel_956732 = array_index_956329 == array_index_949087 ? add_956730 : sel_956726;
  assign add_956735 = sel_956732 + 8'h01;
  assign sel_956736 = array_index_956731 == array_index_948483 ? add_956735 : sel_956732;
  assign add_956739 = sel_956736 + 8'h01;
  assign sel_956740 = array_index_956731 == array_index_948487 ? add_956739 : sel_956736;
  assign add_956743 = sel_956740 + 8'h01;
  assign sel_956744 = array_index_956731 == array_index_948495 ? add_956743 : sel_956740;
  assign add_956747 = sel_956744 + 8'h01;
  assign sel_956748 = array_index_956731 == array_index_948503 ? add_956747 : sel_956744;
  assign add_956751 = sel_956748 + 8'h01;
  assign sel_956752 = array_index_956731 == array_index_948511 ? add_956751 : sel_956748;
  assign add_956755 = sel_956752 + 8'h01;
  assign sel_956756 = array_index_956731 == array_index_948519 ? add_956755 : sel_956752;
  assign add_956759 = sel_956756 + 8'h01;
  assign sel_956760 = array_index_956731 == array_index_948527 ? add_956759 : sel_956756;
  assign add_956763 = sel_956760 + 8'h01;
  assign sel_956764 = array_index_956731 == array_index_948535 ? add_956763 : sel_956760;
  assign add_956767 = sel_956764 + 8'h01;
  assign sel_956768 = array_index_956731 == array_index_948541 ? add_956767 : sel_956764;
  assign add_956771 = sel_956768 + 8'h01;
  assign sel_956772 = array_index_956731 == array_index_948547 ? add_956771 : sel_956768;
  assign add_956775 = sel_956772 + 8'h01;
  assign sel_956776 = array_index_956731 == array_index_948553 ? add_956775 : sel_956772;
  assign add_956779 = sel_956776 + 8'h01;
  assign sel_956780 = array_index_956731 == array_index_948559 ? add_956779 : sel_956776;
  assign add_956783 = sel_956780 + 8'h01;
  assign sel_956784 = array_index_956731 == array_index_948565 ? add_956783 : sel_956780;
  assign add_956787 = sel_956784 + 8'h01;
  assign sel_956788 = array_index_956731 == array_index_948571 ? add_956787 : sel_956784;
  assign add_956791 = sel_956788 + 8'h01;
  assign sel_956792 = array_index_956731 == array_index_948577 ? add_956791 : sel_956788;
  assign add_956795 = sel_956792 + 8'h01;
  assign sel_956796 = array_index_956731 == array_index_948583 ? add_956795 : sel_956792;
  assign add_956799 = sel_956796 + 8'h01;
  assign sel_956800 = array_index_956731 == array_index_948589 ? add_956799 : sel_956796;
  assign add_956803 = sel_956800 + 8'h01;
  assign sel_956804 = array_index_956731 == array_index_948595 ? add_956803 : sel_956800;
  assign add_956807 = sel_956804 + 8'h01;
  assign sel_956808 = array_index_956731 == array_index_948601 ? add_956807 : sel_956804;
  assign add_956811 = sel_956808 + 8'h01;
  assign sel_956812 = array_index_956731 == array_index_948607 ? add_956811 : sel_956808;
  assign add_956815 = sel_956812 + 8'h01;
  assign sel_956816 = array_index_956731 == array_index_948613 ? add_956815 : sel_956812;
  assign add_956819 = sel_956816 + 8'h01;
  assign sel_956820 = array_index_956731 == array_index_948619 ? add_956819 : sel_956816;
  assign add_956823 = sel_956820 + 8'h01;
  assign sel_956824 = array_index_956731 == array_index_948625 ? add_956823 : sel_956820;
  assign add_956827 = sel_956824 + 8'h01;
  assign sel_956828 = array_index_956731 == array_index_948631 ? add_956827 : sel_956824;
  assign add_956831 = sel_956828 + 8'h01;
  assign sel_956832 = array_index_956731 == array_index_948637 ? add_956831 : sel_956828;
  assign add_956835 = sel_956832 + 8'h01;
  assign sel_956836 = array_index_956731 == array_index_948643 ? add_956835 : sel_956832;
  assign add_956839 = sel_956836 + 8'h01;
  assign sel_956840 = array_index_956731 == array_index_948649 ? add_956839 : sel_956836;
  assign add_956843 = sel_956840 + 8'h01;
  assign sel_956844 = array_index_956731 == array_index_948655 ? add_956843 : sel_956840;
  assign add_956847 = sel_956844 + 8'h01;
  assign sel_956848 = array_index_956731 == array_index_948661 ? add_956847 : sel_956844;
  assign add_956851 = sel_956848 + 8'h01;
  assign sel_956852 = array_index_956731 == array_index_948667 ? add_956851 : sel_956848;
  assign add_956855 = sel_956852 + 8'h01;
  assign sel_956856 = array_index_956731 == array_index_948673 ? add_956855 : sel_956852;
  assign add_956859 = sel_956856 + 8'h01;
  assign sel_956860 = array_index_956731 == array_index_948679 ? add_956859 : sel_956856;
  assign add_956863 = sel_956860 + 8'h01;
  assign sel_956864 = array_index_956731 == array_index_948685 ? add_956863 : sel_956860;
  assign add_956867 = sel_956864 + 8'h01;
  assign sel_956868 = array_index_956731 == array_index_948691 ? add_956867 : sel_956864;
  assign add_956871 = sel_956868 + 8'h01;
  assign sel_956872 = array_index_956731 == array_index_948697 ? add_956871 : sel_956868;
  assign add_956875 = sel_956872 + 8'h01;
  assign sel_956876 = array_index_956731 == array_index_948703 ? add_956875 : sel_956872;
  assign add_956879 = sel_956876 + 8'h01;
  assign sel_956880 = array_index_956731 == array_index_948709 ? add_956879 : sel_956876;
  assign add_956883 = sel_956880 + 8'h01;
  assign sel_956884 = array_index_956731 == array_index_948715 ? add_956883 : sel_956880;
  assign add_956887 = sel_956884 + 8'h01;
  assign sel_956888 = array_index_956731 == array_index_948721 ? add_956887 : sel_956884;
  assign add_956891 = sel_956888 + 8'h01;
  assign sel_956892 = array_index_956731 == array_index_948727 ? add_956891 : sel_956888;
  assign add_956895 = sel_956892 + 8'h01;
  assign sel_956896 = array_index_956731 == array_index_948733 ? add_956895 : sel_956892;
  assign add_956899 = sel_956896 + 8'h01;
  assign sel_956900 = array_index_956731 == array_index_948739 ? add_956899 : sel_956896;
  assign add_956903 = sel_956900 + 8'h01;
  assign sel_956904 = array_index_956731 == array_index_948745 ? add_956903 : sel_956900;
  assign add_956907 = sel_956904 + 8'h01;
  assign sel_956908 = array_index_956731 == array_index_948751 ? add_956907 : sel_956904;
  assign add_956911 = sel_956908 + 8'h01;
  assign sel_956912 = array_index_956731 == array_index_948757 ? add_956911 : sel_956908;
  assign add_956915 = sel_956912 + 8'h01;
  assign sel_956916 = array_index_956731 == array_index_948763 ? add_956915 : sel_956912;
  assign add_956919 = sel_956916 + 8'h01;
  assign sel_956920 = array_index_956731 == array_index_948769 ? add_956919 : sel_956916;
  assign add_956923 = sel_956920 + 8'h01;
  assign sel_956924 = array_index_956731 == array_index_948775 ? add_956923 : sel_956920;
  assign add_956927 = sel_956924 + 8'h01;
  assign sel_956928 = array_index_956731 == array_index_948781 ? add_956927 : sel_956924;
  assign add_956931 = sel_956928 + 8'h01;
  assign sel_956932 = array_index_956731 == array_index_948787 ? add_956931 : sel_956928;
  assign add_956935 = sel_956932 + 8'h01;
  assign sel_956936 = array_index_956731 == array_index_948793 ? add_956935 : sel_956932;
  assign add_956939 = sel_956936 + 8'h01;
  assign sel_956940 = array_index_956731 == array_index_948799 ? add_956939 : sel_956936;
  assign add_956943 = sel_956940 + 8'h01;
  assign sel_956944 = array_index_956731 == array_index_948805 ? add_956943 : sel_956940;
  assign add_956947 = sel_956944 + 8'h01;
  assign sel_956948 = array_index_956731 == array_index_948811 ? add_956947 : sel_956944;
  assign add_956951 = sel_956948 + 8'h01;
  assign sel_956952 = array_index_956731 == array_index_948817 ? add_956951 : sel_956948;
  assign add_956955 = sel_956952 + 8'h01;
  assign sel_956956 = array_index_956731 == array_index_948823 ? add_956955 : sel_956952;
  assign add_956959 = sel_956956 + 8'h01;
  assign sel_956960 = array_index_956731 == array_index_948829 ? add_956959 : sel_956956;
  assign add_956963 = sel_956960 + 8'h01;
  assign sel_956964 = array_index_956731 == array_index_948835 ? add_956963 : sel_956960;
  assign add_956967 = sel_956964 + 8'h01;
  assign sel_956968 = array_index_956731 == array_index_948841 ? add_956967 : sel_956964;
  assign add_956971 = sel_956968 + 8'h01;
  assign sel_956972 = array_index_956731 == array_index_948847 ? add_956971 : sel_956968;
  assign add_956975 = sel_956972 + 8'h01;
  assign sel_956976 = array_index_956731 == array_index_948853 ? add_956975 : sel_956972;
  assign add_956979 = sel_956976 + 8'h01;
  assign sel_956980 = array_index_956731 == array_index_948859 ? add_956979 : sel_956976;
  assign add_956983 = sel_956980 + 8'h01;
  assign sel_956984 = array_index_956731 == array_index_948865 ? add_956983 : sel_956980;
  assign add_956987 = sel_956984 + 8'h01;
  assign sel_956988 = array_index_956731 == array_index_948871 ? add_956987 : sel_956984;
  assign add_956991 = sel_956988 + 8'h01;
  assign sel_956992 = array_index_956731 == array_index_948877 ? add_956991 : sel_956988;
  assign add_956995 = sel_956992 + 8'h01;
  assign sel_956996 = array_index_956731 == array_index_948883 ? add_956995 : sel_956992;
  assign add_956999 = sel_956996 + 8'h01;
  assign sel_957000 = array_index_956731 == array_index_948889 ? add_956999 : sel_956996;
  assign add_957003 = sel_957000 + 8'h01;
  assign sel_957004 = array_index_956731 == array_index_948895 ? add_957003 : sel_957000;
  assign add_957007 = sel_957004 + 8'h01;
  assign sel_957008 = array_index_956731 == array_index_948901 ? add_957007 : sel_957004;
  assign add_957011 = sel_957008 + 8'h01;
  assign sel_957012 = array_index_956731 == array_index_948907 ? add_957011 : sel_957008;
  assign add_957015 = sel_957012 + 8'h01;
  assign sel_957016 = array_index_956731 == array_index_948913 ? add_957015 : sel_957012;
  assign add_957019 = sel_957016 + 8'h01;
  assign sel_957020 = array_index_956731 == array_index_948919 ? add_957019 : sel_957016;
  assign add_957023 = sel_957020 + 8'h01;
  assign sel_957024 = array_index_956731 == array_index_948925 ? add_957023 : sel_957020;
  assign add_957027 = sel_957024 + 8'h01;
  assign sel_957028 = array_index_956731 == array_index_948931 ? add_957027 : sel_957024;
  assign add_957031 = sel_957028 + 8'h01;
  assign sel_957032 = array_index_956731 == array_index_948937 ? add_957031 : sel_957028;
  assign add_957035 = sel_957032 + 8'h01;
  assign sel_957036 = array_index_956731 == array_index_948943 ? add_957035 : sel_957032;
  assign add_957039 = sel_957036 + 8'h01;
  assign sel_957040 = array_index_956731 == array_index_948949 ? add_957039 : sel_957036;
  assign add_957043 = sel_957040 + 8'h01;
  assign sel_957044 = array_index_956731 == array_index_948955 ? add_957043 : sel_957040;
  assign add_957047 = sel_957044 + 8'h01;
  assign sel_957048 = array_index_956731 == array_index_948961 ? add_957047 : sel_957044;
  assign add_957051 = sel_957048 + 8'h01;
  assign sel_957052 = array_index_956731 == array_index_948967 ? add_957051 : sel_957048;
  assign add_957055 = sel_957052 + 8'h01;
  assign sel_957056 = array_index_956731 == array_index_948973 ? add_957055 : sel_957052;
  assign add_957059 = sel_957056 + 8'h01;
  assign sel_957060 = array_index_956731 == array_index_948979 ? add_957059 : sel_957056;
  assign add_957063 = sel_957060 + 8'h01;
  assign sel_957064 = array_index_956731 == array_index_948985 ? add_957063 : sel_957060;
  assign add_957067 = sel_957064 + 8'h01;
  assign sel_957068 = array_index_956731 == array_index_948991 ? add_957067 : sel_957064;
  assign add_957071 = sel_957068 + 8'h01;
  assign sel_957072 = array_index_956731 == array_index_948997 ? add_957071 : sel_957068;
  assign add_957075 = sel_957072 + 8'h01;
  assign sel_957076 = array_index_956731 == array_index_949003 ? add_957075 : sel_957072;
  assign add_957079 = sel_957076 + 8'h01;
  assign sel_957080 = array_index_956731 == array_index_949009 ? add_957079 : sel_957076;
  assign add_957083 = sel_957080 + 8'h01;
  assign sel_957084 = array_index_956731 == array_index_949015 ? add_957083 : sel_957080;
  assign add_957087 = sel_957084 + 8'h01;
  assign sel_957088 = array_index_956731 == array_index_949021 ? add_957087 : sel_957084;
  assign add_957091 = sel_957088 + 8'h01;
  assign sel_957092 = array_index_956731 == array_index_949027 ? add_957091 : sel_957088;
  assign add_957095 = sel_957092 + 8'h01;
  assign sel_957096 = array_index_956731 == array_index_949033 ? add_957095 : sel_957092;
  assign add_957099 = sel_957096 + 8'h01;
  assign sel_957100 = array_index_956731 == array_index_949039 ? add_957099 : sel_957096;
  assign add_957103 = sel_957100 + 8'h01;
  assign sel_957104 = array_index_956731 == array_index_949045 ? add_957103 : sel_957100;
  assign add_957107 = sel_957104 + 8'h01;
  assign sel_957108 = array_index_956731 == array_index_949051 ? add_957107 : sel_957104;
  assign add_957111 = sel_957108 + 8'h01;
  assign sel_957112 = array_index_956731 == array_index_949057 ? add_957111 : sel_957108;
  assign add_957115 = sel_957112 + 8'h01;
  assign sel_957116 = array_index_956731 == array_index_949063 ? add_957115 : sel_957112;
  assign add_957119 = sel_957116 + 8'h01;
  assign sel_957120 = array_index_956731 == array_index_949069 ? add_957119 : sel_957116;
  assign add_957123 = sel_957120 + 8'h01;
  assign sel_957124 = array_index_956731 == array_index_949075 ? add_957123 : sel_957120;
  assign add_957127 = sel_957124 + 8'h01;
  assign sel_957128 = array_index_956731 == array_index_949081 ? add_957127 : sel_957124;
  assign add_957132 = sel_957128 + 8'h01;
  assign array_index_957133 = set1_unflattened[7'h15];
  assign sel_957134 = array_index_956731 == array_index_949087 ? add_957132 : sel_957128;
  assign add_957137 = sel_957134 + 8'h01;
  assign sel_957138 = array_index_957133 == array_index_948483 ? add_957137 : sel_957134;
  assign add_957141 = sel_957138 + 8'h01;
  assign sel_957142 = array_index_957133 == array_index_948487 ? add_957141 : sel_957138;
  assign add_957145 = sel_957142 + 8'h01;
  assign sel_957146 = array_index_957133 == array_index_948495 ? add_957145 : sel_957142;
  assign add_957149 = sel_957146 + 8'h01;
  assign sel_957150 = array_index_957133 == array_index_948503 ? add_957149 : sel_957146;
  assign add_957153 = sel_957150 + 8'h01;
  assign sel_957154 = array_index_957133 == array_index_948511 ? add_957153 : sel_957150;
  assign add_957157 = sel_957154 + 8'h01;
  assign sel_957158 = array_index_957133 == array_index_948519 ? add_957157 : sel_957154;
  assign add_957161 = sel_957158 + 8'h01;
  assign sel_957162 = array_index_957133 == array_index_948527 ? add_957161 : sel_957158;
  assign add_957165 = sel_957162 + 8'h01;
  assign sel_957166 = array_index_957133 == array_index_948535 ? add_957165 : sel_957162;
  assign add_957169 = sel_957166 + 8'h01;
  assign sel_957170 = array_index_957133 == array_index_948541 ? add_957169 : sel_957166;
  assign add_957173 = sel_957170 + 8'h01;
  assign sel_957174 = array_index_957133 == array_index_948547 ? add_957173 : sel_957170;
  assign add_957177 = sel_957174 + 8'h01;
  assign sel_957178 = array_index_957133 == array_index_948553 ? add_957177 : sel_957174;
  assign add_957181 = sel_957178 + 8'h01;
  assign sel_957182 = array_index_957133 == array_index_948559 ? add_957181 : sel_957178;
  assign add_957185 = sel_957182 + 8'h01;
  assign sel_957186 = array_index_957133 == array_index_948565 ? add_957185 : sel_957182;
  assign add_957189 = sel_957186 + 8'h01;
  assign sel_957190 = array_index_957133 == array_index_948571 ? add_957189 : sel_957186;
  assign add_957193 = sel_957190 + 8'h01;
  assign sel_957194 = array_index_957133 == array_index_948577 ? add_957193 : sel_957190;
  assign add_957197 = sel_957194 + 8'h01;
  assign sel_957198 = array_index_957133 == array_index_948583 ? add_957197 : sel_957194;
  assign add_957201 = sel_957198 + 8'h01;
  assign sel_957202 = array_index_957133 == array_index_948589 ? add_957201 : sel_957198;
  assign add_957205 = sel_957202 + 8'h01;
  assign sel_957206 = array_index_957133 == array_index_948595 ? add_957205 : sel_957202;
  assign add_957209 = sel_957206 + 8'h01;
  assign sel_957210 = array_index_957133 == array_index_948601 ? add_957209 : sel_957206;
  assign add_957213 = sel_957210 + 8'h01;
  assign sel_957214 = array_index_957133 == array_index_948607 ? add_957213 : sel_957210;
  assign add_957217 = sel_957214 + 8'h01;
  assign sel_957218 = array_index_957133 == array_index_948613 ? add_957217 : sel_957214;
  assign add_957221 = sel_957218 + 8'h01;
  assign sel_957222 = array_index_957133 == array_index_948619 ? add_957221 : sel_957218;
  assign add_957225 = sel_957222 + 8'h01;
  assign sel_957226 = array_index_957133 == array_index_948625 ? add_957225 : sel_957222;
  assign add_957229 = sel_957226 + 8'h01;
  assign sel_957230 = array_index_957133 == array_index_948631 ? add_957229 : sel_957226;
  assign add_957233 = sel_957230 + 8'h01;
  assign sel_957234 = array_index_957133 == array_index_948637 ? add_957233 : sel_957230;
  assign add_957237 = sel_957234 + 8'h01;
  assign sel_957238 = array_index_957133 == array_index_948643 ? add_957237 : sel_957234;
  assign add_957241 = sel_957238 + 8'h01;
  assign sel_957242 = array_index_957133 == array_index_948649 ? add_957241 : sel_957238;
  assign add_957245 = sel_957242 + 8'h01;
  assign sel_957246 = array_index_957133 == array_index_948655 ? add_957245 : sel_957242;
  assign add_957249 = sel_957246 + 8'h01;
  assign sel_957250 = array_index_957133 == array_index_948661 ? add_957249 : sel_957246;
  assign add_957253 = sel_957250 + 8'h01;
  assign sel_957254 = array_index_957133 == array_index_948667 ? add_957253 : sel_957250;
  assign add_957257 = sel_957254 + 8'h01;
  assign sel_957258 = array_index_957133 == array_index_948673 ? add_957257 : sel_957254;
  assign add_957261 = sel_957258 + 8'h01;
  assign sel_957262 = array_index_957133 == array_index_948679 ? add_957261 : sel_957258;
  assign add_957265 = sel_957262 + 8'h01;
  assign sel_957266 = array_index_957133 == array_index_948685 ? add_957265 : sel_957262;
  assign add_957269 = sel_957266 + 8'h01;
  assign sel_957270 = array_index_957133 == array_index_948691 ? add_957269 : sel_957266;
  assign add_957273 = sel_957270 + 8'h01;
  assign sel_957274 = array_index_957133 == array_index_948697 ? add_957273 : sel_957270;
  assign add_957277 = sel_957274 + 8'h01;
  assign sel_957278 = array_index_957133 == array_index_948703 ? add_957277 : sel_957274;
  assign add_957281 = sel_957278 + 8'h01;
  assign sel_957282 = array_index_957133 == array_index_948709 ? add_957281 : sel_957278;
  assign add_957285 = sel_957282 + 8'h01;
  assign sel_957286 = array_index_957133 == array_index_948715 ? add_957285 : sel_957282;
  assign add_957289 = sel_957286 + 8'h01;
  assign sel_957290 = array_index_957133 == array_index_948721 ? add_957289 : sel_957286;
  assign add_957293 = sel_957290 + 8'h01;
  assign sel_957294 = array_index_957133 == array_index_948727 ? add_957293 : sel_957290;
  assign add_957297 = sel_957294 + 8'h01;
  assign sel_957298 = array_index_957133 == array_index_948733 ? add_957297 : sel_957294;
  assign add_957301 = sel_957298 + 8'h01;
  assign sel_957302 = array_index_957133 == array_index_948739 ? add_957301 : sel_957298;
  assign add_957305 = sel_957302 + 8'h01;
  assign sel_957306 = array_index_957133 == array_index_948745 ? add_957305 : sel_957302;
  assign add_957309 = sel_957306 + 8'h01;
  assign sel_957310 = array_index_957133 == array_index_948751 ? add_957309 : sel_957306;
  assign add_957313 = sel_957310 + 8'h01;
  assign sel_957314 = array_index_957133 == array_index_948757 ? add_957313 : sel_957310;
  assign add_957317 = sel_957314 + 8'h01;
  assign sel_957318 = array_index_957133 == array_index_948763 ? add_957317 : sel_957314;
  assign add_957321 = sel_957318 + 8'h01;
  assign sel_957322 = array_index_957133 == array_index_948769 ? add_957321 : sel_957318;
  assign add_957325 = sel_957322 + 8'h01;
  assign sel_957326 = array_index_957133 == array_index_948775 ? add_957325 : sel_957322;
  assign add_957329 = sel_957326 + 8'h01;
  assign sel_957330 = array_index_957133 == array_index_948781 ? add_957329 : sel_957326;
  assign add_957333 = sel_957330 + 8'h01;
  assign sel_957334 = array_index_957133 == array_index_948787 ? add_957333 : sel_957330;
  assign add_957337 = sel_957334 + 8'h01;
  assign sel_957338 = array_index_957133 == array_index_948793 ? add_957337 : sel_957334;
  assign add_957341 = sel_957338 + 8'h01;
  assign sel_957342 = array_index_957133 == array_index_948799 ? add_957341 : sel_957338;
  assign add_957345 = sel_957342 + 8'h01;
  assign sel_957346 = array_index_957133 == array_index_948805 ? add_957345 : sel_957342;
  assign add_957349 = sel_957346 + 8'h01;
  assign sel_957350 = array_index_957133 == array_index_948811 ? add_957349 : sel_957346;
  assign add_957353 = sel_957350 + 8'h01;
  assign sel_957354 = array_index_957133 == array_index_948817 ? add_957353 : sel_957350;
  assign add_957357 = sel_957354 + 8'h01;
  assign sel_957358 = array_index_957133 == array_index_948823 ? add_957357 : sel_957354;
  assign add_957361 = sel_957358 + 8'h01;
  assign sel_957362 = array_index_957133 == array_index_948829 ? add_957361 : sel_957358;
  assign add_957365 = sel_957362 + 8'h01;
  assign sel_957366 = array_index_957133 == array_index_948835 ? add_957365 : sel_957362;
  assign add_957369 = sel_957366 + 8'h01;
  assign sel_957370 = array_index_957133 == array_index_948841 ? add_957369 : sel_957366;
  assign add_957373 = sel_957370 + 8'h01;
  assign sel_957374 = array_index_957133 == array_index_948847 ? add_957373 : sel_957370;
  assign add_957377 = sel_957374 + 8'h01;
  assign sel_957378 = array_index_957133 == array_index_948853 ? add_957377 : sel_957374;
  assign add_957381 = sel_957378 + 8'h01;
  assign sel_957382 = array_index_957133 == array_index_948859 ? add_957381 : sel_957378;
  assign add_957385 = sel_957382 + 8'h01;
  assign sel_957386 = array_index_957133 == array_index_948865 ? add_957385 : sel_957382;
  assign add_957389 = sel_957386 + 8'h01;
  assign sel_957390 = array_index_957133 == array_index_948871 ? add_957389 : sel_957386;
  assign add_957393 = sel_957390 + 8'h01;
  assign sel_957394 = array_index_957133 == array_index_948877 ? add_957393 : sel_957390;
  assign add_957397 = sel_957394 + 8'h01;
  assign sel_957398 = array_index_957133 == array_index_948883 ? add_957397 : sel_957394;
  assign add_957401 = sel_957398 + 8'h01;
  assign sel_957402 = array_index_957133 == array_index_948889 ? add_957401 : sel_957398;
  assign add_957405 = sel_957402 + 8'h01;
  assign sel_957406 = array_index_957133 == array_index_948895 ? add_957405 : sel_957402;
  assign add_957409 = sel_957406 + 8'h01;
  assign sel_957410 = array_index_957133 == array_index_948901 ? add_957409 : sel_957406;
  assign add_957413 = sel_957410 + 8'h01;
  assign sel_957414 = array_index_957133 == array_index_948907 ? add_957413 : sel_957410;
  assign add_957417 = sel_957414 + 8'h01;
  assign sel_957418 = array_index_957133 == array_index_948913 ? add_957417 : sel_957414;
  assign add_957421 = sel_957418 + 8'h01;
  assign sel_957422 = array_index_957133 == array_index_948919 ? add_957421 : sel_957418;
  assign add_957425 = sel_957422 + 8'h01;
  assign sel_957426 = array_index_957133 == array_index_948925 ? add_957425 : sel_957422;
  assign add_957429 = sel_957426 + 8'h01;
  assign sel_957430 = array_index_957133 == array_index_948931 ? add_957429 : sel_957426;
  assign add_957433 = sel_957430 + 8'h01;
  assign sel_957434 = array_index_957133 == array_index_948937 ? add_957433 : sel_957430;
  assign add_957437 = sel_957434 + 8'h01;
  assign sel_957438 = array_index_957133 == array_index_948943 ? add_957437 : sel_957434;
  assign add_957441 = sel_957438 + 8'h01;
  assign sel_957442 = array_index_957133 == array_index_948949 ? add_957441 : sel_957438;
  assign add_957445 = sel_957442 + 8'h01;
  assign sel_957446 = array_index_957133 == array_index_948955 ? add_957445 : sel_957442;
  assign add_957449 = sel_957446 + 8'h01;
  assign sel_957450 = array_index_957133 == array_index_948961 ? add_957449 : sel_957446;
  assign add_957453 = sel_957450 + 8'h01;
  assign sel_957454 = array_index_957133 == array_index_948967 ? add_957453 : sel_957450;
  assign add_957457 = sel_957454 + 8'h01;
  assign sel_957458 = array_index_957133 == array_index_948973 ? add_957457 : sel_957454;
  assign add_957461 = sel_957458 + 8'h01;
  assign sel_957462 = array_index_957133 == array_index_948979 ? add_957461 : sel_957458;
  assign add_957465 = sel_957462 + 8'h01;
  assign sel_957466 = array_index_957133 == array_index_948985 ? add_957465 : sel_957462;
  assign add_957469 = sel_957466 + 8'h01;
  assign sel_957470 = array_index_957133 == array_index_948991 ? add_957469 : sel_957466;
  assign add_957473 = sel_957470 + 8'h01;
  assign sel_957474 = array_index_957133 == array_index_948997 ? add_957473 : sel_957470;
  assign add_957477 = sel_957474 + 8'h01;
  assign sel_957478 = array_index_957133 == array_index_949003 ? add_957477 : sel_957474;
  assign add_957481 = sel_957478 + 8'h01;
  assign sel_957482 = array_index_957133 == array_index_949009 ? add_957481 : sel_957478;
  assign add_957485 = sel_957482 + 8'h01;
  assign sel_957486 = array_index_957133 == array_index_949015 ? add_957485 : sel_957482;
  assign add_957489 = sel_957486 + 8'h01;
  assign sel_957490 = array_index_957133 == array_index_949021 ? add_957489 : sel_957486;
  assign add_957493 = sel_957490 + 8'h01;
  assign sel_957494 = array_index_957133 == array_index_949027 ? add_957493 : sel_957490;
  assign add_957497 = sel_957494 + 8'h01;
  assign sel_957498 = array_index_957133 == array_index_949033 ? add_957497 : sel_957494;
  assign add_957501 = sel_957498 + 8'h01;
  assign sel_957502 = array_index_957133 == array_index_949039 ? add_957501 : sel_957498;
  assign add_957505 = sel_957502 + 8'h01;
  assign sel_957506 = array_index_957133 == array_index_949045 ? add_957505 : sel_957502;
  assign add_957509 = sel_957506 + 8'h01;
  assign sel_957510 = array_index_957133 == array_index_949051 ? add_957509 : sel_957506;
  assign add_957513 = sel_957510 + 8'h01;
  assign sel_957514 = array_index_957133 == array_index_949057 ? add_957513 : sel_957510;
  assign add_957517 = sel_957514 + 8'h01;
  assign sel_957518 = array_index_957133 == array_index_949063 ? add_957517 : sel_957514;
  assign add_957521 = sel_957518 + 8'h01;
  assign sel_957522 = array_index_957133 == array_index_949069 ? add_957521 : sel_957518;
  assign add_957525 = sel_957522 + 8'h01;
  assign sel_957526 = array_index_957133 == array_index_949075 ? add_957525 : sel_957522;
  assign add_957529 = sel_957526 + 8'h01;
  assign sel_957530 = array_index_957133 == array_index_949081 ? add_957529 : sel_957526;
  assign add_957534 = sel_957530 + 8'h01;
  assign array_index_957535 = set1_unflattened[7'h16];
  assign sel_957536 = array_index_957133 == array_index_949087 ? add_957534 : sel_957530;
  assign add_957539 = sel_957536 + 8'h01;
  assign sel_957540 = array_index_957535 == array_index_948483 ? add_957539 : sel_957536;
  assign add_957543 = sel_957540 + 8'h01;
  assign sel_957544 = array_index_957535 == array_index_948487 ? add_957543 : sel_957540;
  assign add_957547 = sel_957544 + 8'h01;
  assign sel_957548 = array_index_957535 == array_index_948495 ? add_957547 : sel_957544;
  assign add_957551 = sel_957548 + 8'h01;
  assign sel_957552 = array_index_957535 == array_index_948503 ? add_957551 : sel_957548;
  assign add_957555 = sel_957552 + 8'h01;
  assign sel_957556 = array_index_957535 == array_index_948511 ? add_957555 : sel_957552;
  assign add_957559 = sel_957556 + 8'h01;
  assign sel_957560 = array_index_957535 == array_index_948519 ? add_957559 : sel_957556;
  assign add_957563 = sel_957560 + 8'h01;
  assign sel_957564 = array_index_957535 == array_index_948527 ? add_957563 : sel_957560;
  assign add_957567 = sel_957564 + 8'h01;
  assign sel_957568 = array_index_957535 == array_index_948535 ? add_957567 : sel_957564;
  assign add_957571 = sel_957568 + 8'h01;
  assign sel_957572 = array_index_957535 == array_index_948541 ? add_957571 : sel_957568;
  assign add_957575 = sel_957572 + 8'h01;
  assign sel_957576 = array_index_957535 == array_index_948547 ? add_957575 : sel_957572;
  assign add_957579 = sel_957576 + 8'h01;
  assign sel_957580 = array_index_957535 == array_index_948553 ? add_957579 : sel_957576;
  assign add_957583 = sel_957580 + 8'h01;
  assign sel_957584 = array_index_957535 == array_index_948559 ? add_957583 : sel_957580;
  assign add_957587 = sel_957584 + 8'h01;
  assign sel_957588 = array_index_957535 == array_index_948565 ? add_957587 : sel_957584;
  assign add_957591 = sel_957588 + 8'h01;
  assign sel_957592 = array_index_957535 == array_index_948571 ? add_957591 : sel_957588;
  assign add_957595 = sel_957592 + 8'h01;
  assign sel_957596 = array_index_957535 == array_index_948577 ? add_957595 : sel_957592;
  assign add_957599 = sel_957596 + 8'h01;
  assign sel_957600 = array_index_957535 == array_index_948583 ? add_957599 : sel_957596;
  assign add_957603 = sel_957600 + 8'h01;
  assign sel_957604 = array_index_957535 == array_index_948589 ? add_957603 : sel_957600;
  assign add_957607 = sel_957604 + 8'h01;
  assign sel_957608 = array_index_957535 == array_index_948595 ? add_957607 : sel_957604;
  assign add_957611 = sel_957608 + 8'h01;
  assign sel_957612 = array_index_957535 == array_index_948601 ? add_957611 : sel_957608;
  assign add_957615 = sel_957612 + 8'h01;
  assign sel_957616 = array_index_957535 == array_index_948607 ? add_957615 : sel_957612;
  assign add_957619 = sel_957616 + 8'h01;
  assign sel_957620 = array_index_957535 == array_index_948613 ? add_957619 : sel_957616;
  assign add_957623 = sel_957620 + 8'h01;
  assign sel_957624 = array_index_957535 == array_index_948619 ? add_957623 : sel_957620;
  assign add_957627 = sel_957624 + 8'h01;
  assign sel_957628 = array_index_957535 == array_index_948625 ? add_957627 : sel_957624;
  assign add_957631 = sel_957628 + 8'h01;
  assign sel_957632 = array_index_957535 == array_index_948631 ? add_957631 : sel_957628;
  assign add_957635 = sel_957632 + 8'h01;
  assign sel_957636 = array_index_957535 == array_index_948637 ? add_957635 : sel_957632;
  assign add_957639 = sel_957636 + 8'h01;
  assign sel_957640 = array_index_957535 == array_index_948643 ? add_957639 : sel_957636;
  assign add_957643 = sel_957640 + 8'h01;
  assign sel_957644 = array_index_957535 == array_index_948649 ? add_957643 : sel_957640;
  assign add_957647 = sel_957644 + 8'h01;
  assign sel_957648 = array_index_957535 == array_index_948655 ? add_957647 : sel_957644;
  assign add_957651 = sel_957648 + 8'h01;
  assign sel_957652 = array_index_957535 == array_index_948661 ? add_957651 : sel_957648;
  assign add_957655 = sel_957652 + 8'h01;
  assign sel_957656 = array_index_957535 == array_index_948667 ? add_957655 : sel_957652;
  assign add_957659 = sel_957656 + 8'h01;
  assign sel_957660 = array_index_957535 == array_index_948673 ? add_957659 : sel_957656;
  assign add_957663 = sel_957660 + 8'h01;
  assign sel_957664 = array_index_957535 == array_index_948679 ? add_957663 : sel_957660;
  assign add_957667 = sel_957664 + 8'h01;
  assign sel_957668 = array_index_957535 == array_index_948685 ? add_957667 : sel_957664;
  assign add_957671 = sel_957668 + 8'h01;
  assign sel_957672 = array_index_957535 == array_index_948691 ? add_957671 : sel_957668;
  assign add_957675 = sel_957672 + 8'h01;
  assign sel_957676 = array_index_957535 == array_index_948697 ? add_957675 : sel_957672;
  assign add_957679 = sel_957676 + 8'h01;
  assign sel_957680 = array_index_957535 == array_index_948703 ? add_957679 : sel_957676;
  assign add_957683 = sel_957680 + 8'h01;
  assign sel_957684 = array_index_957535 == array_index_948709 ? add_957683 : sel_957680;
  assign add_957687 = sel_957684 + 8'h01;
  assign sel_957688 = array_index_957535 == array_index_948715 ? add_957687 : sel_957684;
  assign add_957691 = sel_957688 + 8'h01;
  assign sel_957692 = array_index_957535 == array_index_948721 ? add_957691 : sel_957688;
  assign add_957695 = sel_957692 + 8'h01;
  assign sel_957696 = array_index_957535 == array_index_948727 ? add_957695 : sel_957692;
  assign add_957699 = sel_957696 + 8'h01;
  assign sel_957700 = array_index_957535 == array_index_948733 ? add_957699 : sel_957696;
  assign add_957703 = sel_957700 + 8'h01;
  assign sel_957704 = array_index_957535 == array_index_948739 ? add_957703 : sel_957700;
  assign add_957707 = sel_957704 + 8'h01;
  assign sel_957708 = array_index_957535 == array_index_948745 ? add_957707 : sel_957704;
  assign add_957711 = sel_957708 + 8'h01;
  assign sel_957712 = array_index_957535 == array_index_948751 ? add_957711 : sel_957708;
  assign add_957715 = sel_957712 + 8'h01;
  assign sel_957716 = array_index_957535 == array_index_948757 ? add_957715 : sel_957712;
  assign add_957719 = sel_957716 + 8'h01;
  assign sel_957720 = array_index_957535 == array_index_948763 ? add_957719 : sel_957716;
  assign add_957723 = sel_957720 + 8'h01;
  assign sel_957724 = array_index_957535 == array_index_948769 ? add_957723 : sel_957720;
  assign add_957727 = sel_957724 + 8'h01;
  assign sel_957728 = array_index_957535 == array_index_948775 ? add_957727 : sel_957724;
  assign add_957731 = sel_957728 + 8'h01;
  assign sel_957732 = array_index_957535 == array_index_948781 ? add_957731 : sel_957728;
  assign add_957735 = sel_957732 + 8'h01;
  assign sel_957736 = array_index_957535 == array_index_948787 ? add_957735 : sel_957732;
  assign add_957739 = sel_957736 + 8'h01;
  assign sel_957740 = array_index_957535 == array_index_948793 ? add_957739 : sel_957736;
  assign add_957743 = sel_957740 + 8'h01;
  assign sel_957744 = array_index_957535 == array_index_948799 ? add_957743 : sel_957740;
  assign add_957747 = sel_957744 + 8'h01;
  assign sel_957748 = array_index_957535 == array_index_948805 ? add_957747 : sel_957744;
  assign add_957751 = sel_957748 + 8'h01;
  assign sel_957752 = array_index_957535 == array_index_948811 ? add_957751 : sel_957748;
  assign add_957755 = sel_957752 + 8'h01;
  assign sel_957756 = array_index_957535 == array_index_948817 ? add_957755 : sel_957752;
  assign add_957759 = sel_957756 + 8'h01;
  assign sel_957760 = array_index_957535 == array_index_948823 ? add_957759 : sel_957756;
  assign add_957763 = sel_957760 + 8'h01;
  assign sel_957764 = array_index_957535 == array_index_948829 ? add_957763 : sel_957760;
  assign add_957767 = sel_957764 + 8'h01;
  assign sel_957768 = array_index_957535 == array_index_948835 ? add_957767 : sel_957764;
  assign add_957771 = sel_957768 + 8'h01;
  assign sel_957772 = array_index_957535 == array_index_948841 ? add_957771 : sel_957768;
  assign add_957775 = sel_957772 + 8'h01;
  assign sel_957776 = array_index_957535 == array_index_948847 ? add_957775 : sel_957772;
  assign add_957779 = sel_957776 + 8'h01;
  assign sel_957780 = array_index_957535 == array_index_948853 ? add_957779 : sel_957776;
  assign add_957783 = sel_957780 + 8'h01;
  assign sel_957784 = array_index_957535 == array_index_948859 ? add_957783 : sel_957780;
  assign add_957787 = sel_957784 + 8'h01;
  assign sel_957788 = array_index_957535 == array_index_948865 ? add_957787 : sel_957784;
  assign add_957791 = sel_957788 + 8'h01;
  assign sel_957792 = array_index_957535 == array_index_948871 ? add_957791 : sel_957788;
  assign add_957795 = sel_957792 + 8'h01;
  assign sel_957796 = array_index_957535 == array_index_948877 ? add_957795 : sel_957792;
  assign add_957799 = sel_957796 + 8'h01;
  assign sel_957800 = array_index_957535 == array_index_948883 ? add_957799 : sel_957796;
  assign add_957803 = sel_957800 + 8'h01;
  assign sel_957804 = array_index_957535 == array_index_948889 ? add_957803 : sel_957800;
  assign add_957807 = sel_957804 + 8'h01;
  assign sel_957808 = array_index_957535 == array_index_948895 ? add_957807 : sel_957804;
  assign add_957811 = sel_957808 + 8'h01;
  assign sel_957812 = array_index_957535 == array_index_948901 ? add_957811 : sel_957808;
  assign add_957815 = sel_957812 + 8'h01;
  assign sel_957816 = array_index_957535 == array_index_948907 ? add_957815 : sel_957812;
  assign add_957819 = sel_957816 + 8'h01;
  assign sel_957820 = array_index_957535 == array_index_948913 ? add_957819 : sel_957816;
  assign add_957823 = sel_957820 + 8'h01;
  assign sel_957824 = array_index_957535 == array_index_948919 ? add_957823 : sel_957820;
  assign add_957827 = sel_957824 + 8'h01;
  assign sel_957828 = array_index_957535 == array_index_948925 ? add_957827 : sel_957824;
  assign add_957831 = sel_957828 + 8'h01;
  assign sel_957832 = array_index_957535 == array_index_948931 ? add_957831 : sel_957828;
  assign add_957835 = sel_957832 + 8'h01;
  assign sel_957836 = array_index_957535 == array_index_948937 ? add_957835 : sel_957832;
  assign add_957839 = sel_957836 + 8'h01;
  assign sel_957840 = array_index_957535 == array_index_948943 ? add_957839 : sel_957836;
  assign add_957843 = sel_957840 + 8'h01;
  assign sel_957844 = array_index_957535 == array_index_948949 ? add_957843 : sel_957840;
  assign add_957847 = sel_957844 + 8'h01;
  assign sel_957848 = array_index_957535 == array_index_948955 ? add_957847 : sel_957844;
  assign add_957851 = sel_957848 + 8'h01;
  assign sel_957852 = array_index_957535 == array_index_948961 ? add_957851 : sel_957848;
  assign add_957855 = sel_957852 + 8'h01;
  assign sel_957856 = array_index_957535 == array_index_948967 ? add_957855 : sel_957852;
  assign add_957859 = sel_957856 + 8'h01;
  assign sel_957860 = array_index_957535 == array_index_948973 ? add_957859 : sel_957856;
  assign add_957863 = sel_957860 + 8'h01;
  assign sel_957864 = array_index_957535 == array_index_948979 ? add_957863 : sel_957860;
  assign add_957867 = sel_957864 + 8'h01;
  assign sel_957868 = array_index_957535 == array_index_948985 ? add_957867 : sel_957864;
  assign add_957871 = sel_957868 + 8'h01;
  assign sel_957872 = array_index_957535 == array_index_948991 ? add_957871 : sel_957868;
  assign add_957875 = sel_957872 + 8'h01;
  assign sel_957876 = array_index_957535 == array_index_948997 ? add_957875 : sel_957872;
  assign add_957879 = sel_957876 + 8'h01;
  assign sel_957880 = array_index_957535 == array_index_949003 ? add_957879 : sel_957876;
  assign add_957883 = sel_957880 + 8'h01;
  assign sel_957884 = array_index_957535 == array_index_949009 ? add_957883 : sel_957880;
  assign add_957887 = sel_957884 + 8'h01;
  assign sel_957888 = array_index_957535 == array_index_949015 ? add_957887 : sel_957884;
  assign add_957891 = sel_957888 + 8'h01;
  assign sel_957892 = array_index_957535 == array_index_949021 ? add_957891 : sel_957888;
  assign add_957895 = sel_957892 + 8'h01;
  assign sel_957896 = array_index_957535 == array_index_949027 ? add_957895 : sel_957892;
  assign add_957899 = sel_957896 + 8'h01;
  assign sel_957900 = array_index_957535 == array_index_949033 ? add_957899 : sel_957896;
  assign add_957903 = sel_957900 + 8'h01;
  assign sel_957904 = array_index_957535 == array_index_949039 ? add_957903 : sel_957900;
  assign add_957907 = sel_957904 + 8'h01;
  assign sel_957908 = array_index_957535 == array_index_949045 ? add_957907 : sel_957904;
  assign add_957911 = sel_957908 + 8'h01;
  assign sel_957912 = array_index_957535 == array_index_949051 ? add_957911 : sel_957908;
  assign add_957915 = sel_957912 + 8'h01;
  assign sel_957916 = array_index_957535 == array_index_949057 ? add_957915 : sel_957912;
  assign add_957919 = sel_957916 + 8'h01;
  assign sel_957920 = array_index_957535 == array_index_949063 ? add_957919 : sel_957916;
  assign add_957923 = sel_957920 + 8'h01;
  assign sel_957924 = array_index_957535 == array_index_949069 ? add_957923 : sel_957920;
  assign add_957927 = sel_957924 + 8'h01;
  assign sel_957928 = array_index_957535 == array_index_949075 ? add_957927 : sel_957924;
  assign add_957931 = sel_957928 + 8'h01;
  assign sel_957932 = array_index_957535 == array_index_949081 ? add_957931 : sel_957928;
  assign add_957936 = sel_957932 + 8'h01;
  assign array_index_957937 = set1_unflattened[7'h17];
  assign sel_957938 = array_index_957535 == array_index_949087 ? add_957936 : sel_957932;
  assign add_957941 = sel_957938 + 8'h01;
  assign sel_957942 = array_index_957937 == array_index_948483 ? add_957941 : sel_957938;
  assign add_957945 = sel_957942 + 8'h01;
  assign sel_957946 = array_index_957937 == array_index_948487 ? add_957945 : sel_957942;
  assign add_957949 = sel_957946 + 8'h01;
  assign sel_957950 = array_index_957937 == array_index_948495 ? add_957949 : sel_957946;
  assign add_957953 = sel_957950 + 8'h01;
  assign sel_957954 = array_index_957937 == array_index_948503 ? add_957953 : sel_957950;
  assign add_957957 = sel_957954 + 8'h01;
  assign sel_957958 = array_index_957937 == array_index_948511 ? add_957957 : sel_957954;
  assign add_957961 = sel_957958 + 8'h01;
  assign sel_957962 = array_index_957937 == array_index_948519 ? add_957961 : sel_957958;
  assign add_957965 = sel_957962 + 8'h01;
  assign sel_957966 = array_index_957937 == array_index_948527 ? add_957965 : sel_957962;
  assign add_957969 = sel_957966 + 8'h01;
  assign sel_957970 = array_index_957937 == array_index_948535 ? add_957969 : sel_957966;
  assign add_957973 = sel_957970 + 8'h01;
  assign sel_957974 = array_index_957937 == array_index_948541 ? add_957973 : sel_957970;
  assign add_957977 = sel_957974 + 8'h01;
  assign sel_957978 = array_index_957937 == array_index_948547 ? add_957977 : sel_957974;
  assign add_957981 = sel_957978 + 8'h01;
  assign sel_957982 = array_index_957937 == array_index_948553 ? add_957981 : sel_957978;
  assign add_957985 = sel_957982 + 8'h01;
  assign sel_957986 = array_index_957937 == array_index_948559 ? add_957985 : sel_957982;
  assign add_957989 = sel_957986 + 8'h01;
  assign sel_957990 = array_index_957937 == array_index_948565 ? add_957989 : sel_957986;
  assign add_957993 = sel_957990 + 8'h01;
  assign sel_957994 = array_index_957937 == array_index_948571 ? add_957993 : sel_957990;
  assign add_957997 = sel_957994 + 8'h01;
  assign sel_957998 = array_index_957937 == array_index_948577 ? add_957997 : sel_957994;
  assign add_958001 = sel_957998 + 8'h01;
  assign sel_958002 = array_index_957937 == array_index_948583 ? add_958001 : sel_957998;
  assign add_958005 = sel_958002 + 8'h01;
  assign sel_958006 = array_index_957937 == array_index_948589 ? add_958005 : sel_958002;
  assign add_958009 = sel_958006 + 8'h01;
  assign sel_958010 = array_index_957937 == array_index_948595 ? add_958009 : sel_958006;
  assign add_958013 = sel_958010 + 8'h01;
  assign sel_958014 = array_index_957937 == array_index_948601 ? add_958013 : sel_958010;
  assign add_958017 = sel_958014 + 8'h01;
  assign sel_958018 = array_index_957937 == array_index_948607 ? add_958017 : sel_958014;
  assign add_958021 = sel_958018 + 8'h01;
  assign sel_958022 = array_index_957937 == array_index_948613 ? add_958021 : sel_958018;
  assign add_958025 = sel_958022 + 8'h01;
  assign sel_958026 = array_index_957937 == array_index_948619 ? add_958025 : sel_958022;
  assign add_958029 = sel_958026 + 8'h01;
  assign sel_958030 = array_index_957937 == array_index_948625 ? add_958029 : sel_958026;
  assign add_958033 = sel_958030 + 8'h01;
  assign sel_958034 = array_index_957937 == array_index_948631 ? add_958033 : sel_958030;
  assign add_958037 = sel_958034 + 8'h01;
  assign sel_958038 = array_index_957937 == array_index_948637 ? add_958037 : sel_958034;
  assign add_958041 = sel_958038 + 8'h01;
  assign sel_958042 = array_index_957937 == array_index_948643 ? add_958041 : sel_958038;
  assign add_958045 = sel_958042 + 8'h01;
  assign sel_958046 = array_index_957937 == array_index_948649 ? add_958045 : sel_958042;
  assign add_958049 = sel_958046 + 8'h01;
  assign sel_958050 = array_index_957937 == array_index_948655 ? add_958049 : sel_958046;
  assign add_958053 = sel_958050 + 8'h01;
  assign sel_958054 = array_index_957937 == array_index_948661 ? add_958053 : sel_958050;
  assign add_958057 = sel_958054 + 8'h01;
  assign sel_958058 = array_index_957937 == array_index_948667 ? add_958057 : sel_958054;
  assign add_958061 = sel_958058 + 8'h01;
  assign sel_958062 = array_index_957937 == array_index_948673 ? add_958061 : sel_958058;
  assign add_958065 = sel_958062 + 8'h01;
  assign sel_958066 = array_index_957937 == array_index_948679 ? add_958065 : sel_958062;
  assign add_958069 = sel_958066 + 8'h01;
  assign sel_958070 = array_index_957937 == array_index_948685 ? add_958069 : sel_958066;
  assign add_958073 = sel_958070 + 8'h01;
  assign sel_958074 = array_index_957937 == array_index_948691 ? add_958073 : sel_958070;
  assign add_958077 = sel_958074 + 8'h01;
  assign sel_958078 = array_index_957937 == array_index_948697 ? add_958077 : sel_958074;
  assign add_958081 = sel_958078 + 8'h01;
  assign sel_958082 = array_index_957937 == array_index_948703 ? add_958081 : sel_958078;
  assign add_958085 = sel_958082 + 8'h01;
  assign sel_958086 = array_index_957937 == array_index_948709 ? add_958085 : sel_958082;
  assign add_958089 = sel_958086 + 8'h01;
  assign sel_958090 = array_index_957937 == array_index_948715 ? add_958089 : sel_958086;
  assign add_958093 = sel_958090 + 8'h01;
  assign sel_958094 = array_index_957937 == array_index_948721 ? add_958093 : sel_958090;
  assign add_958097 = sel_958094 + 8'h01;
  assign sel_958098 = array_index_957937 == array_index_948727 ? add_958097 : sel_958094;
  assign add_958101 = sel_958098 + 8'h01;
  assign sel_958102 = array_index_957937 == array_index_948733 ? add_958101 : sel_958098;
  assign add_958105 = sel_958102 + 8'h01;
  assign sel_958106 = array_index_957937 == array_index_948739 ? add_958105 : sel_958102;
  assign add_958109 = sel_958106 + 8'h01;
  assign sel_958110 = array_index_957937 == array_index_948745 ? add_958109 : sel_958106;
  assign add_958113 = sel_958110 + 8'h01;
  assign sel_958114 = array_index_957937 == array_index_948751 ? add_958113 : sel_958110;
  assign add_958117 = sel_958114 + 8'h01;
  assign sel_958118 = array_index_957937 == array_index_948757 ? add_958117 : sel_958114;
  assign add_958121 = sel_958118 + 8'h01;
  assign sel_958122 = array_index_957937 == array_index_948763 ? add_958121 : sel_958118;
  assign add_958125 = sel_958122 + 8'h01;
  assign sel_958126 = array_index_957937 == array_index_948769 ? add_958125 : sel_958122;
  assign add_958129 = sel_958126 + 8'h01;
  assign sel_958130 = array_index_957937 == array_index_948775 ? add_958129 : sel_958126;
  assign add_958133 = sel_958130 + 8'h01;
  assign sel_958134 = array_index_957937 == array_index_948781 ? add_958133 : sel_958130;
  assign add_958137 = sel_958134 + 8'h01;
  assign sel_958138 = array_index_957937 == array_index_948787 ? add_958137 : sel_958134;
  assign add_958141 = sel_958138 + 8'h01;
  assign sel_958142 = array_index_957937 == array_index_948793 ? add_958141 : sel_958138;
  assign add_958145 = sel_958142 + 8'h01;
  assign sel_958146 = array_index_957937 == array_index_948799 ? add_958145 : sel_958142;
  assign add_958149 = sel_958146 + 8'h01;
  assign sel_958150 = array_index_957937 == array_index_948805 ? add_958149 : sel_958146;
  assign add_958153 = sel_958150 + 8'h01;
  assign sel_958154 = array_index_957937 == array_index_948811 ? add_958153 : sel_958150;
  assign add_958157 = sel_958154 + 8'h01;
  assign sel_958158 = array_index_957937 == array_index_948817 ? add_958157 : sel_958154;
  assign add_958161 = sel_958158 + 8'h01;
  assign sel_958162 = array_index_957937 == array_index_948823 ? add_958161 : sel_958158;
  assign add_958165 = sel_958162 + 8'h01;
  assign sel_958166 = array_index_957937 == array_index_948829 ? add_958165 : sel_958162;
  assign add_958169 = sel_958166 + 8'h01;
  assign sel_958170 = array_index_957937 == array_index_948835 ? add_958169 : sel_958166;
  assign add_958173 = sel_958170 + 8'h01;
  assign sel_958174 = array_index_957937 == array_index_948841 ? add_958173 : sel_958170;
  assign add_958177 = sel_958174 + 8'h01;
  assign sel_958178 = array_index_957937 == array_index_948847 ? add_958177 : sel_958174;
  assign add_958181 = sel_958178 + 8'h01;
  assign sel_958182 = array_index_957937 == array_index_948853 ? add_958181 : sel_958178;
  assign add_958185 = sel_958182 + 8'h01;
  assign sel_958186 = array_index_957937 == array_index_948859 ? add_958185 : sel_958182;
  assign add_958189 = sel_958186 + 8'h01;
  assign sel_958190 = array_index_957937 == array_index_948865 ? add_958189 : sel_958186;
  assign add_958193 = sel_958190 + 8'h01;
  assign sel_958194 = array_index_957937 == array_index_948871 ? add_958193 : sel_958190;
  assign add_958197 = sel_958194 + 8'h01;
  assign sel_958198 = array_index_957937 == array_index_948877 ? add_958197 : sel_958194;
  assign add_958201 = sel_958198 + 8'h01;
  assign sel_958202 = array_index_957937 == array_index_948883 ? add_958201 : sel_958198;
  assign add_958205 = sel_958202 + 8'h01;
  assign sel_958206 = array_index_957937 == array_index_948889 ? add_958205 : sel_958202;
  assign add_958209 = sel_958206 + 8'h01;
  assign sel_958210 = array_index_957937 == array_index_948895 ? add_958209 : sel_958206;
  assign add_958213 = sel_958210 + 8'h01;
  assign sel_958214 = array_index_957937 == array_index_948901 ? add_958213 : sel_958210;
  assign add_958217 = sel_958214 + 8'h01;
  assign sel_958218 = array_index_957937 == array_index_948907 ? add_958217 : sel_958214;
  assign add_958221 = sel_958218 + 8'h01;
  assign sel_958222 = array_index_957937 == array_index_948913 ? add_958221 : sel_958218;
  assign add_958225 = sel_958222 + 8'h01;
  assign sel_958226 = array_index_957937 == array_index_948919 ? add_958225 : sel_958222;
  assign add_958229 = sel_958226 + 8'h01;
  assign sel_958230 = array_index_957937 == array_index_948925 ? add_958229 : sel_958226;
  assign add_958233 = sel_958230 + 8'h01;
  assign sel_958234 = array_index_957937 == array_index_948931 ? add_958233 : sel_958230;
  assign add_958237 = sel_958234 + 8'h01;
  assign sel_958238 = array_index_957937 == array_index_948937 ? add_958237 : sel_958234;
  assign add_958241 = sel_958238 + 8'h01;
  assign sel_958242 = array_index_957937 == array_index_948943 ? add_958241 : sel_958238;
  assign add_958245 = sel_958242 + 8'h01;
  assign sel_958246 = array_index_957937 == array_index_948949 ? add_958245 : sel_958242;
  assign add_958249 = sel_958246 + 8'h01;
  assign sel_958250 = array_index_957937 == array_index_948955 ? add_958249 : sel_958246;
  assign add_958253 = sel_958250 + 8'h01;
  assign sel_958254 = array_index_957937 == array_index_948961 ? add_958253 : sel_958250;
  assign add_958257 = sel_958254 + 8'h01;
  assign sel_958258 = array_index_957937 == array_index_948967 ? add_958257 : sel_958254;
  assign add_958261 = sel_958258 + 8'h01;
  assign sel_958262 = array_index_957937 == array_index_948973 ? add_958261 : sel_958258;
  assign add_958265 = sel_958262 + 8'h01;
  assign sel_958266 = array_index_957937 == array_index_948979 ? add_958265 : sel_958262;
  assign add_958269 = sel_958266 + 8'h01;
  assign sel_958270 = array_index_957937 == array_index_948985 ? add_958269 : sel_958266;
  assign add_958273 = sel_958270 + 8'h01;
  assign sel_958274 = array_index_957937 == array_index_948991 ? add_958273 : sel_958270;
  assign add_958277 = sel_958274 + 8'h01;
  assign sel_958278 = array_index_957937 == array_index_948997 ? add_958277 : sel_958274;
  assign add_958281 = sel_958278 + 8'h01;
  assign sel_958282 = array_index_957937 == array_index_949003 ? add_958281 : sel_958278;
  assign add_958285 = sel_958282 + 8'h01;
  assign sel_958286 = array_index_957937 == array_index_949009 ? add_958285 : sel_958282;
  assign add_958289 = sel_958286 + 8'h01;
  assign sel_958290 = array_index_957937 == array_index_949015 ? add_958289 : sel_958286;
  assign add_958293 = sel_958290 + 8'h01;
  assign sel_958294 = array_index_957937 == array_index_949021 ? add_958293 : sel_958290;
  assign add_958297 = sel_958294 + 8'h01;
  assign sel_958298 = array_index_957937 == array_index_949027 ? add_958297 : sel_958294;
  assign add_958301 = sel_958298 + 8'h01;
  assign sel_958302 = array_index_957937 == array_index_949033 ? add_958301 : sel_958298;
  assign add_958305 = sel_958302 + 8'h01;
  assign sel_958306 = array_index_957937 == array_index_949039 ? add_958305 : sel_958302;
  assign add_958309 = sel_958306 + 8'h01;
  assign sel_958310 = array_index_957937 == array_index_949045 ? add_958309 : sel_958306;
  assign add_958313 = sel_958310 + 8'h01;
  assign sel_958314 = array_index_957937 == array_index_949051 ? add_958313 : sel_958310;
  assign add_958317 = sel_958314 + 8'h01;
  assign sel_958318 = array_index_957937 == array_index_949057 ? add_958317 : sel_958314;
  assign add_958321 = sel_958318 + 8'h01;
  assign sel_958322 = array_index_957937 == array_index_949063 ? add_958321 : sel_958318;
  assign add_958325 = sel_958322 + 8'h01;
  assign sel_958326 = array_index_957937 == array_index_949069 ? add_958325 : sel_958322;
  assign add_958329 = sel_958326 + 8'h01;
  assign sel_958330 = array_index_957937 == array_index_949075 ? add_958329 : sel_958326;
  assign add_958333 = sel_958330 + 8'h01;
  assign sel_958334 = array_index_957937 == array_index_949081 ? add_958333 : sel_958330;
  assign add_958338 = sel_958334 + 8'h01;
  assign array_index_958339 = set1_unflattened[7'h18];
  assign sel_958340 = array_index_957937 == array_index_949087 ? add_958338 : sel_958334;
  assign add_958343 = sel_958340 + 8'h01;
  assign sel_958344 = array_index_958339 == array_index_948483 ? add_958343 : sel_958340;
  assign add_958347 = sel_958344 + 8'h01;
  assign sel_958348 = array_index_958339 == array_index_948487 ? add_958347 : sel_958344;
  assign add_958351 = sel_958348 + 8'h01;
  assign sel_958352 = array_index_958339 == array_index_948495 ? add_958351 : sel_958348;
  assign add_958355 = sel_958352 + 8'h01;
  assign sel_958356 = array_index_958339 == array_index_948503 ? add_958355 : sel_958352;
  assign add_958359 = sel_958356 + 8'h01;
  assign sel_958360 = array_index_958339 == array_index_948511 ? add_958359 : sel_958356;
  assign add_958363 = sel_958360 + 8'h01;
  assign sel_958364 = array_index_958339 == array_index_948519 ? add_958363 : sel_958360;
  assign add_958367 = sel_958364 + 8'h01;
  assign sel_958368 = array_index_958339 == array_index_948527 ? add_958367 : sel_958364;
  assign add_958371 = sel_958368 + 8'h01;
  assign sel_958372 = array_index_958339 == array_index_948535 ? add_958371 : sel_958368;
  assign add_958375 = sel_958372 + 8'h01;
  assign sel_958376 = array_index_958339 == array_index_948541 ? add_958375 : sel_958372;
  assign add_958379 = sel_958376 + 8'h01;
  assign sel_958380 = array_index_958339 == array_index_948547 ? add_958379 : sel_958376;
  assign add_958383 = sel_958380 + 8'h01;
  assign sel_958384 = array_index_958339 == array_index_948553 ? add_958383 : sel_958380;
  assign add_958387 = sel_958384 + 8'h01;
  assign sel_958388 = array_index_958339 == array_index_948559 ? add_958387 : sel_958384;
  assign add_958391 = sel_958388 + 8'h01;
  assign sel_958392 = array_index_958339 == array_index_948565 ? add_958391 : sel_958388;
  assign add_958395 = sel_958392 + 8'h01;
  assign sel_958396 = array_index_958339 == array_index_948571 ? add_958395 : sel_958392;
  assign add_958399 = sel_958396 + 8'h01;
  assign sel_958400 = array_index_958339 == array_index_948577 ? add_958399 : sel_958396;
  assign add_958403 = sel_958400 + 8'h01;
  assign sel_958404 = array_index_958339 == array_index_948583 ? add_958403 : sel_958400;
  assign add_958407 = sel_958404 + 8'h01;
  assign sel_958408 = array_index_958339 == array_index_948589 ? add_958407 : sel_958404;
  assign add_958411 = sel_958408 + 8'h01;
  assign sel_958412 = array_index_958339 == array_index_948595 ? add_958411 : sel_958408;
  assign add_958415 = sel_958412 + 8'h01;
  assign sel_958416 = array_index_958339 == array_index_948601 ? add_958415 : sel_958412;
  assign add_958419 = sel_958416 + 8'h01;
  assign sel_958420 = array_index_958339 == array_index_948607 ? add_958419 : sel_958416;
  assign add_958423 = sel_958420 + 8'h01;
  assign sel_958424 = array_index_958339 == array_index_948613 ? add_958423 : sel_958420;
  assign add_958427 = sel_958424 + 8'h01;
  assign sel_958428 = array_index_958339 == array_index_948619 ? add_958427 : sel_958424;
  assign add_958431 = sel_958428 + 8'h01;
  assign sel_958432 = array_index_958339 == array_index_948625 ? add_958431 : sel_958428;
  assign add_958435 = sel_958432 + 8'h01;
  assign sel_958436 = array_index_958339 == array_index_948631 ? add_958435 : sel_958432;
  assign add_958439 = sel_958436 + 8'h01;
  assign sel_958440 = array_index_958339 == array_index_948637 ? add_958439 : sel_958436;
  assign add_958443 = sel_958440 + 8'h01;
  assign sel_958444 = array_index_958339 == array_index_948643 ? add_958443 : sel_958440;
  assign add_958447 = sel_958444 + 8'h01;
  assign sel_958448 = array_index_958339 == array_index_948649 ? add_958447 : sel_958444;
  assign add_958451 = sel_958448 + 8'h01;
  assign sel_958452 = array_index_958339 == array_index_948655 ? add_958451 : sel_958448;
  assign add_958455 = sel_958452 + 8'h01;
  assign sel_958456 = array_index_958339 == array_index_948661 ? add_958455 : sel_958452;
  assign add_958459 = sel_958456 + 8'h01;
  assign sel_958460 = array_index_958339 == array_index_948667 ? add_958459 : sel_958456;
  assign add_958463 = sel_958460 + 8'h01;
  assign sel_958464 = array_index_958339 == array_index_948673 ? add_958463 : sel_958460;
  assign add_958467 = sel_958464 + 8'h01;
  assign sel_958468 = array_index_958339 == array_index_948679 ? add_958467 : sel_958464;
  assign add_958471 = sel_958468 + 8'h01;
  assign sel_958472 = array_index_958339 == array_index_948685 ? add_958471 : sel_958468;
  assign add_958475 = sel_958472 + 8'h01;
  assign sel_958476 = array_index_958339 == array_index_948691 ? add_958475 : sel_958472;
  assign add_958479 = sel_958476 + 8'h01;
  assign sel_958480 = array_index_958339 == array_index_948697 ? add_958479 : sel_958476;
  assign add_958483 = sel_958480 + 8'h01;
  assign sel_958484 = array_index_958339 == array_index_948703 ? add_958483 : sel_958480;
  assign add_958487 = sel_958484 + 8'h01;
  assign sel_958488 = array_index_958339 == array_index_948709 ? add_958487 : sel_958484;
  assign add_958491 = sel_958488 + 8'h01;
  assign sel_958492 = array_index_958339 == array_index_948715 ? add_958491 : sel_958488;
  assign add_958495 = sel_958492 + 8'h01;
  assign sel_958496 = array_index_958339 == array_index_948721 ? add_958495 : sel_958492;
  assign add_958499 = sel_958496 + 8'h01;
  assign sel_958500 = array_index_958339 == array_index_948727 ? add_958499 : sel_958496;
  assign add_958503 = sel_958500 + 8'h01;
  assign sel_958504 = array_index_958339 == array_index_948733 ? add_958503 : sel_958500;
  assign add_958507 = sel_958504 + 8'h01;
  assign sel_958508 = array_index_958339 == array_index_948739 ? add_958507 : sel_958504;
  assign add_958511 = sel_958508 + 8'h01;
  assign sel_958512 = array_index_958339 == array_index_948745 ? add_958511 : sel_958508;
  assign add_958515 = sel_958512 + 8'h01;
  assign sel_958516 = array_index_958339 == array_index_948751 ? add_958515 : sel_958512;
  assign add_958519 = sel_958516 + 8'h01;
  assign sel_958520 = array_index_958339 == array_index_948757 ? add_958519 : sel_958516;
  assign add_958523 = sel_958520 + 8'h01;
  assign sel_958524 = array_index_958339 == array_index_948763 ? add_958523 : sel_958520;
  assign add_958527 = sel_958524 + 8'h01;
  assign sel_958528 = array_index_958339 == array_index_948769 ? add_958527 : sel_958524;
  assign add_958531 = sel_958528 + 8'h01;
  assign sel_958532 = array_index_958339 == array_index_948775 ? add_958531 : sel_958528;
  assign add_958535 = sel_958532 + 8'h01;
  assign sel_958536 = array_index_958339 == array_index_948781 ? add_958535 : sel_958532;
  assign add_958539 = sel_958536 + 8'h01;
  assign sel_958540 = array_index_958339 == array_index_948787 ? add_958539 : sel_958536;
  assign add_958543 = sel_958540 + 8'h01;
  assign sel_958544 = array_index_958339 == array_index_948793 ? add_958543 : sel_958540;
  assign add_958547 = sel_958544 + 8'h01;
  assign sel_958548 = array_index_958339 == array_index_948799 ? add_958547 : sel_958544;
  assign add_958551 = sel_958548 + 8'h01;
  assign sel_958552 = array_index_958339 == array_index_948805 ? add_958551 : sel_958548;
  assign add_958555 = sel_958552 + 8'h01;
  assign sel_958556 = array_index_958339 == array_index_948811 ? add_958555 : sel_958552;
  assign add_958559 = sel_958556 + 8'h01;
  assign sel_958560 = array_index_958339 == array_index_948817 ? add_958559 : sel_958556;
  assign add_958563 = sel_958560 + 8'h01;
  assign sel_958564 = array_index_958339 == array_index_948823 ? add_958563 : sel_958560;
  assign add_958567 = sel_958564 + 8'h01;
  assign sel_958568 = array_index_958339 == array_index_948829 ? add_958567 : sel_958564;
  assign add_958571 = sel_958568 + 8'h01;
  assign sel_958572 = array_index_958339 == array_index_948835 ? add_958571 : sel_958568;
  assign add_958575 = sel_958572 + 8'h01;
  assign sel_958576 = array_index_958339 == array_index_948841 ? add_958575 : sel_958572;
  assign add_958579 = sel_958576 + 8'h01;
  assign sel_958580 = array_index_958339 == array_index_948847 ? add_958579 : sel_958576;
  assign add_958583 = sel_958580 + 8'h01;
  assign sel_958584 = array_index_958339 == array_index_948853 ? add_958583 : sel_958580;
  assign add_958587 = sel_958584 + 8'h01;
  assign sel_958588 = array_index_958339 == array_index_948859 ? add_958587 : sel_958584;
  assign add_958591 = sel_958588 + 8'h01;
  assign sel_958592 = array_index_958339 == array_index_948865 ? add_958591 : sel_958588;
  assign add_958595 = sel_958592 + 8'h01;
  assign sel_958596 = array_index_958339 == array_index_948871 ? add_958595 : sel_958592;
  assign add_958599 = sel_958596 + 8'h01;
  assign sel_958600 = array_index_958339 == array_index_948877 ? add_958599 : sel_958596;
  assign add_958603 = sel_958600 + 8'h01;
  assign sel_958604 = array_index_958339 == array_index_948883 ? add_958603 : sel_958600;
  assign add_958607 = sel_958604 + 8'h01;
  assign sel_958608 = array_index_958339 == array_index_948889 ? add_958607 : sel_958604;
  assign add_958611 = sel_958608 + 8'h01;
  assign sel_958612 = array_index_958339 == array_index_948895 ? add_958611 : sel_958608;
  assign add_958615 = sel_958612 + 8'h01;
  assign sel_958616 = array_index_958339 == array_index_948901 ? add_958615 : sel_958612;
  assign add_958619 = sel_958616 + 8'h01;
  assign sel_958620 = array_index_958339 == array_index_948907 ? add_958619 : sel_958616;
  assign add_958623 = sel_958620 + 8'h01;
  assign sel_958624 = array_index_958339 == array_index_948913 ? add_958623 : sel_958620;
  assign add_958627 = sel_958624 + 8'h01;
  assign sel_958628 = array_index_958339 == array_index_948919 ? add_958627 : sel_958624;
  assign add_958631 = sel_958628 + 8'h01;
  assign sel_958632 = array_index_958339 == array_index_948925 ? add_958631 : sel_958628;
  assign add_958635 = sel_958632 + 8'h01;
  assign sel_958636 = array_index_958339 == array_index_948931 ? add_958635 : sel_958632;
  assign add_958639 = sel_958636 + 8'h01;
  assign sel_958640 = array_index_958339 == array_index_948937 ? add_958639 : sel_958636;
  assign add_958643 = sel_958640 + 8'h01;
  assign sel_958644 = array_index_958339 == array_index_948943 ? add_958643 : sel_958640;
  assign add_958647 = sel_958644 + 8'h01;
  assign sel_958648 = array_index_958339 == array_index_948949 ? add_958647 : sel_958644;
  assign add_958651 = sel_958648 + 8'h01;
  assign sel_958652 = array_index_958339 == array_index_948955 ? add_958651 : sel_958648;
  assign add_958655 = sel_958652 + 8'h01;
  assign sel_958656 = array_index_958339 == array_index_948961 ? add_958655 : sel_958652;
  assign add_958659 = sel_958656 + 8'h01;
  assign sel_958660 = array_index_958339 == array_index_948967 ? add_958659 : sel_958656;
  assign add_958663 = sel_958660 + 8'h01;
  assign sel_958664 = array_index_958339 == array_index_948973 ? add_958663 : sel_958660;
  assign add_958667 = sel_958664 + 8'h01;
  assign sel_958668 = array_index_958339 == array_index_948979 ? add_958667 : sel_958664;
  assign add_958671 = sel_958668 + 8'h01;
  assign sel_958672 = array_index_958339 == array_index_948985 ? add_958671 : sel_958668;
  assign add_958675 = sel_958672 + 8'h01;
  assign sel_958676 = array_index_958339 == array_index_948991 ? add_958675 : sel_958672;
  assign add_958679 = sel_958676 + 8'h01;
  assign sel_958680 = array_index_958339 == array_index_948997 ? add_958679 : sel_958676;
  assign add_958683 = sel_958680 + 8'h01;
  assign sel_958684 = array_index_958339 == array_index_949003 ? add_958683 : sel_958680;
  assign add_958687 = sel_958684 + 8'h01;
  assign sel_958688 = array_index_958339 == array_index_949009 ? add_958687 : sel_958684;
  assign add_958691 = sel_958688 + 8'h01;
  assign sel_958692 = array_index_958339 == array_index_949015 ? add_958691 : sel_958688;
  assign add_958695 = sel_958692 + 8'h01;
  assign sel_958696 = array_index_958339 == array_index_949021 ? add_958695 : sel_958692;
  assign add_958699 = sel_958696 + 8'h01;
  assign sel_958700 = array_index_958339 == array_index_949027 ? add_958699 : sel_958696;
  assign add_958703 = sel_958700 + 8'h01;
  assign sel_958704 = array_index_958339 == array_index_949033 ? add_958703 : sel_958700;
  assign add_958707 = sel_958704 + 8'h01;
  assign sel_958708 = array_index_958339 == array_index_949039 ? add_958707 : sel_958704;
  assign add_958711 = sel_958708 + 8'h01;
  assign sel_958712 = array_index_958339 == array_index_949045 ? add_958711 : sel_958708;
  assign add_958715 = sel_958712 + 8'h01;
  assign sel_958716 = array_index_958339 == array_index_949051 ? add_958715 : sel_958712;
  assign add_958719 = sel_958716 + 8'h01;
  assign sel_958720 = array_index_958339 == array_index_949057 ? add_958719 : sel_958716;
  assign add_958723 = sel_958720 + 8'h01;
  assign sel_958724 = array_index_958339 == array_index_949063 ? add_958723 : sel_958720;
  assign add_958727 = sel_958724 + 8'h01;
  assign sel_958728 = array_index_958339 == array_index_949069 ? add_958727 : sel_958724;
  assign add_958731 = sel_958728 + 8'h01;
  assign sel_958732 = array_index_958339 == array_index_949075 ? add_958731 : sel_958728;
  assign add_958735 = sel_958732 + 8'h01;
  assign sel_958736 = array_index_958339 == array_index_949081 ? add_958735 : sel_958732;
  assign add_958740 = sel_958736 + 8'h01;
  assign array_index_958741 = set1_unflattened[7'h19];
  assign sel_958742 = array_index_958339 == array_index_949087 ? add_958740 : sel_958736;
  assign add_958745 = sel_958742 + 8'h01;
  assign sel_958746 = array_index_958741 == array_index_948483 ? add_958745 : sel_958742;
  assign add_958749 = sel_958746 + 8'h01;
  assign sel_958750 = array_index_958741 == array_index_948487 ? add_958749 : sel_958746;
  assign add_958753 = sel_958750 + 8'h01;
  assign sel_958754 = array_index_958741 == array_index_948495 ? add_958753 : sel_958750;
  assign add_958757 = sel_958754 + 8'h01;
  assign sel_958758 = array_index_958741 == array_index_948503 ? add_958757 : sel_958754;
  assign add_958761 = sel_958758 + 8'h01;
  assign sel_958762 = array_index_958741 == array_index_948511 ? add_958761 : sel_958758;
  assign add_958765 = sel_958762 + 8'h01;
  assign sel_958766 = array_index_958741 == array_index_948519 ? add_958765 : sel_958762;
  assign add_958769 = sel_958766 + 8'h01;
  assign sel_958770 = array_index_958741 == array_index_948527 ? add_958769 : sel_958766;
  assign add_958773 = sel_958770 + 8'h01;
  assign sel_958774 = array_index_958741 == array_index_948535 ? add_958773 : sel_958770;
  assign add_958777 = sel_958774 + 8'h01;
  assign sel_958778 = array_index_958741 == array_index_948541 ? add_958777 : sel_958774;
  assign add_958781 = sel_958778 + 8'h01;
  assign sel_958782 = array_index_958741 == array_index_948547 ? add_958781 : sel_958778;
  assign add_958785 = sel_958782 + 8'h01;
  assign sel_958786 = array_index_958741 == array_index_948553 ? add_958785 : sel_958782;
  assign add_958789 = sel_958786 + 8'h01;
  assign sel_958790 = array_index_958741 == array_index_948559 ? add_958789 : sel_958786;
  assign add_958793 = sel_958790 + 8'h01;
  assign sel_958794 = array_index_958741 == array_index_948565 ? add_958793 : sel_958790;
  assign add_958797 = sel_958794 + 8'h01;
  assign sel_958798 = array_index_958741 == array_index_948571 ? add_958797 : sel_958794;
  assign add_958801 = sel_958798 + 8'h01;
  assign sel_958802 = array_index_958741 == array_index_948577 ? add_958801 : sel_958798;
  assign add_958805 = sel_958802 + 8'h01;
  assign sel_958806 = array_index_958741 == array_index_948583 ? add_958805 : sel_958802;
  assign add_958809 = sel_958806 + 8'h01;
  assign sel_958810 = array_index_958741 == array_index_948589 ? add_958809 : sel_958806;
  assign add_958813 = sel_958810 + 8'h01;
  assign sel_958814 = array_index_958741 == array_index_948595 ? add_958813 : sel_958810;
  assign add_958817 = sel_958814 + 8'h01;
  assign sel_958818 = array_index_958741 == array_index_948601 ? add_958817 : sel_958814;
  assign add_958821 = sel_958818 + 8'h01;
  assign sel_958822 = array_index_958741 == array_index_948607 ? add_958821 : sel_958818;
  assign add_958825 = sel_958822 + 8'h01;
  assign sel_958826 = array_index_958741 == array_index_948613 ? add_958825 : sel_958822;
  assign add_958829 = sel_958826 + 8'h01;
  assign sel_958830 = array_index_958741 == array_index_948619 ? add_958829 : sel_958826;
  assign add_958833 = sel_958830 + 8'h01;
  assign sel_958834 = array_index_958741 == array_index_948625 ? add_958833 : sel_958830;
  assign add_958837 = sel_958834 + 8'h01;
  assign sel_958838 = array_index_958741 == array_index_948631 ? add_958837 : sel_958834;
  assign add_958841 = sel_958838 + 8'h01;
  assign sel_958842 = array_index_958741 == array_index_948637 ? add_958841 : sel_958838;
  assign add_958845 = sel_958842 + 8'h01;
  assign sel_958846 = array_index_958741 == array_index_948643 ? add_958845 : sel_958842;
  assign add_958849 = sel_958846 + 8'h01;
  assign sel_958850 = array_index_958741 == array_index_948649 ? add_958849 : sel_958846;
  assign add_958853 = sel_958850 + 8'h01;
  assign sel_958854 = array_index_958741 == array_index_948655 ? add_958853 : sel_958850;
  assign add_958857 = sel_958854 + 8'h01;
  assign sel_958858 = array_index_958741 == array_index_948661 ? add_958857 : sel_958854;
  assign add_958861 = sel_958858 + 8'h01;
  assign sel_958862 = array_index_958741 == array_index_948667 ? add_958861 : sel_958858;
  assign add_958865 = sel_958862 + 8'h01;
  assign sel_958866 = array_index_958741 == array_index_948673 ? add_958865 : sel_958862;
  assign add_958869 = sel_958866 + 8'h01;
  assign sel_958870 = array_index_958741 == array_index_948679 ? add_958869 : sel_958866;
  assign add_958873 = sel_958870 + 8'h01;
  assign sel_958874 = array_index_958741 == array_index_948685 ? add_958873 : sel_958870;
  assign add_958877 = sel_958874 + 8'h01;
  assign sel_958878 = array_index_958741 == array_index_948691 ? add_958877 : sel_958874;
  assign add_958881 = sel_958878 + 8'h01;
  assign sel_958882 = array_index_958741 == array_index_948697 ? add_958881 : sel_958878;
  assign add_958885 = sel_958882 + 8'h01;
  assign sel_958886 = array_index_958741 == array_index_948703 ? add_958885 : sel_958882;
  assign add_958889 = sel_958886 + 8'h01;
  assign sel_958890 = array_index_958741 == array_index_948709 ? add_958889 : sel_958886;
  assign add_958893 = sel_958890 + 8'h01;
  assign sel_958894 = array_index_958741 == array_index_948715 ? add_958893 : sel_958890;
  assign add_958897 = sel_958894 + 8'h01;
  assign sel_958898 = array_index_958741 == array_index_948721 ? add_958897 : sel_958894;
  assign add_958901 = sel_958898 + 8'h01;
  assign sel_958902 = array_index_958741 == array_index_948727 ? add_958901 : sel_958898;
  assign add_958905 = sel_958902 + 8'h01;
  assign sel_958906 = array_index_958741 == array_index_948733 ? add_958905 : sel_958902;
  assign add_958909 = sel_958906 + 8'h01;
  assign sel_958910 = array_index_958741 == array_index_948739 ? add_958909 : sel_958906;
  assign add_958913 = sel_958910 + 8'h01;
  assign sel_958914 = array_index_958741 == array_index_948745 ? add_958913 : sel_958910;
  assign add_958917 = sel_958914 + 8'h01;
  assign sel_958918 = array_index_958741 == array_index_948751 ? add_958917 : sel_958914;
  assign add_958921 = sel_958918 + 8'h01;
  assign sel_958922 = array_index_958741 == array_index_948757 ? add_958921 : sel_958918;
  assign add_958925 = sel_958922 + 8'h01;
  assign sel_958926 = array_index_958741 == array_index_948763 ? add_958925 : sel_958922;
  assign add_958929 = sel_958926 + 8'h01;
  assign sel_958930 = array_index_958741 == array_index_948769 ? add_958929 : sel_958926;
  assign add_958933 = sel_958930 + 8'h01;
  assign sel_958934 = array_index_958741 == array_index_948775 ? add_958933 : sel_958930;
  assign add_958937 = sel_958934 + 8'h01;
  assign sel_958938 = array_index_958741 == array_index_948781 ? add_958937 : sel_958934;
  assign add_958941 = sel_958938 + 8'h01;
  assign sel_958942 = array_index_958741 == array_index_948787 ? add_958941 : sel_958938;
  assign add_958945 = sel_958942 + 8'h01;
  assign sel_958946 = array_index_958741 == array_index_948793 ? add_958945 : sel_958942;
  assign add_958949 = sel_958946 + 8'h01;
  assign sel_958950 = array_index_958741 == array_index_948799 ? add_958949 : sel_958946;
  assign add_958953 = sel_958950 + 8'h01;
  assign sel_958954 = array_index_958741 == array_index_948805 ? add_958953 : sel_958950;
  assign add_958957 = sel_958954 + 8'h01;
  assign sel_958958 = array_index_958741 == array_index_948811 ? add_958957 : sel_958954;
  assign add_958961 = sel_958958 + 8'h01;
  assign sel_958962 = array_index_958741 == array_index_948817 ? add_958961 : sel_958958;
  assign add_958965 = sel_958962 + 8'h01;
  assign sel_958966 = array_index_958741 == array_index_948823 ? add_958965 : sel_958962;
  assign add_958969 = sel_958966 + 8'h01;
  assign sel_958970 = array_index_958741 == array_index_948829 ? add_958969 : sel_958966;
  assign add_958973 = sel_958970 + 8'h01;
  assign sel_958974 = array_index_958741 == array_index_948835 ? add_958973 : sel_958970;
  assign add_958977 = sel_958974 + 8'h01;
  assign sel_958978 = array_index_958741 == array_index_948841 ? add_958977 : sel_958974;
  assign add_958981 = sel_958978 + 8'h01;
  assign sel_958982 = array_index_958741 == array_index_948847 ? add_958981 : sel_958978;
  assign add_958985 = sel_958982 + 8'h01;
  assign sel_958986 = array_index_958741 == array_index_948853 ? add_958985 : sel_958982;
  assign add_958989 = sel_958986 + 8'h01;
  assign sel_958990 = array_index_958741 == array_index_948859 ? add_958989 : sel_958986;
  assign add_958993 = sel_958990 + 8'h01;
  assign sel_958994 = array_index_958741 == array_index_948865 ? add_958993 : sel_958990;
  assign add_958997 = sel_958994 + 8'h01;
  assign sel_958998 = array_index_958741 == array_index_948871 ? add_958997 : sel_958994;
  assign add_959001 = sel_958998 + 8'h01;
  assign sel_959002 = array_index_958741 == array_index_948877 ? add_959001 : sel_958998;
  assign add_959005 = sel_959002 + 8'h01;
  assign sel_959006 = array_index_958741 == array_index_948883 ? add_959005 : sel_959002;
  assign add_959009 = sel_959006 + 8'h01;
  assign sel_959010 = array_index_958741 == array_index_948889 ? add_959009 : sel_959006;
  assign add_959013 = sel_959010 + 8'h01;
  assign sel_959014 = array_index_958741 == array_index_948895 ? add_959013 : sel_959010;
  assign add_959017 = sel_959014 + 8'h01;
  assign sel_959018 = array_index_958741 == array_index_948901 ? add_959017 : sel_959014;
  assign add_959021 = sel_959018 + 8'h01;
  assign sel_959022 = array_index_958741 == array_index_948907 ? add_959021 : sel_959018;
  assign add_959025 = sel_959022 + 8'h01;
  assign sel_959026 = array_index_958741 == array_index_948913 ? add_959025 : sel_959022;
  assign add_959029 = sel_959026 + 8'h01;
  assign sel_959030 = array_index_958741 == array_index_948919 ? add_959029 : sel_959026;
  assign add_959033 = sel_959030 + 8'h01;
  assign sel_959034 = array_index_958741 == array_index_948925 ? add_959033 : sel_959030;
  assign add_959037 = sel_959034 + 8'h01;
  assign sel_959038 = array_index_958741 == array_index_948931 ? add_959037 : sel_959034;
  assign add_959041 = sel_959038 + 8'h01;
  assign sel_959042 = array_index_958741 == array_index_948937 ? add_959041 : sel_959038;
  assign add_959045 = sel_959042 + 8'h01;
  assign sel_959046 = array_index_958741 == array_index_948943 ? add_959045 : sel_959042;
  assign add_959049 = sel_959046 + 8'h01;
  assign sel_959050 = array_index_958741 == array_index_948949 ? add_959049 : sel_959046;
  assign add_959053 = sel_959050 + 8'h01;
  assign sel_959054 = array_index_958741 == array_index_948955 ? add_959053 : sel_959050;
  assign add_959057 = sel_959054 + 8'h01;
  assign sel_959058 = array_index_958741 == array_index_948961 ? add_959057 : sel_959054;
  assign add_959061 = sel_959058 + 8'h01;
  assign sel_959062 = array_index_958741 == array_index_948967 ? add_959061 : sel_959058;
  assign add_959065 = sel_959062 + 8'h01;
  assign sel_959066 = array_index_958741 == array_index_948973 ? add_959065 : sel_959062;
  assign add_959069 = sel_959066 + 8'h01;
  assign sel_959070 = array_index_958741 == array_index_948979 ? add_959069 : sel_959066;
  assign add_959073 = sel_959070 + 8'h01;
  assign sel_959074 = array_index_958741 == array_index_948985 ? add_959073 : sel_959070;
  assign add_959077 = sel_959074 + 8'h01;
  assign sel_959078 = array_index_958741 == array_index_948991 ? add_959077 : sel_959074;
  assign add_959081 = sel_959078 + 8'h01;
  assign sel_959082 = array_index_958741 == array_index_948997 ? add_959081 : sel_959078;
  assign add_959085 = sel_959082 + 8'h01;
  assign sel_959086 = array_index_958741 == array_index_949003 ? add_959085 : sel_959082;
  assign add_959089 = sel_959086 + 8'h01;
  assign sel_959090 = array_index_958741 == array_index_949009 ? add_959089 : sel_959086;
  assign add_959093 = sel_959090 + 8'h01;
  assign sel_959094 = array_index_958741 == array_index_949015 ? add_959093 : sel_959090;
  assign add_959097 = sel_959094 + 8'h01;
  assign sel_959098 = array_index_958741 == array_index_949021 ? add_959097 : sel_959094;
  assign add_959101 = sel_959098 + 8'h01;
  assign sel_959102 = array_index_958741 == array_index_949027 ? add_959101 : sel_959098;
  assign add_959105 = sel_959102 + 8'h01;
  assign sel_959106 = array_index_958741 == array_index_949033 ? add_959105 : sel_959102;
  assign add_959109 = sel_959106 + 8'h01;
  assign sel_959110 = array_index_958741 == array_index_949039 ? add_959109 : sel_959106;
  assign add_959113 = sel_959110 + 8'h01;
  assign sel_959114 = array_index_958741 == array_index_949045 ? add_959113 : sel_959110;
  assign add_959117 = sel_959114 + 8'h01;
  assign sel_959118 = array_index_958741 == array_index_949051 ? add_959117 : sel_959114;
  assign add_959121 = sel_959118 + 8'h01;
  assign sel_959122 = array_index_958741 == array_index_949057 ? add_959121 : sel_959118;
  assign add_959125 = sel_959122 + 8'h01;
  assign sel_959126 = array_index_958741 == array_index_949063 ? add_959125 : sel_959122;
  assign add_959129 = sel_959126 + 8'h01;
  assign sel_959130 = array_index_958741 == array_index_949069 ? add_959129 : sel_959126;
  assign add_959133 = sel_959130 + 8'h01;
  assign sel_959134 = array_index_958741 == array_index_949075 ? add_959133 : sel_959130;
  assign add_959137 = sel_959134 + 8'h01;
  assign sel_959138 = array_index_958741 == array_index_949081 ? add_959137 : sel_959134;
  assign add_959142 = sel_959138 + 8'h01;
  assign array_index_959143 = set1_unflattened[7'h1a];
  assign sel_959144 = array_index_958741 == array_index_949087 ? add_959142 : sel_959138;
  assign add_959147 = sel_959144 + 8'h01;
  assign sel_959148 = array_index_959143 == array_index_948483 ? add_959147 : sel_959144;
  assign add_959151 = sel_959148 + 8'h01;
  assign sel_959152 = array_index_959143 == array_index_948487 ? add_959151 : sel_959148;
  assign add_959155 = sel_959152 + 8'h01;
  assign sel_959156 = array_index_959143 == array_index_948495 ? add_959155 : sel_959152;
  assign add_959159 = sel_959156 + 8'h01;
  assign sel_959160 = array_index_959143 == array_index_948503 ? add_959159 : sel_959156;
  assign add_959163 = sel_959160 + 8'h01;
  assign sel_959164 = array_index_959143 == array_index_948511 ? add_959163 : sel_959160;
  assign add_959167 = sel_959164 + 8'h01;
  assign sel_959168 = array_index_959143 == array_index_948519 ? add_959167 : sel_959164;
  assign add_959171 = sel_959168 + 8'h01;
  assign sel_959172 = array_index_959143 == array_index_948527 ? add_959171 : sel_959168;
  assign add_959175 = sel_959172 + 8'h01;
  assign sel_959176 = array_index_959143 == array_index_948535 ? add_959175 : sel_959172;
  assign add_959179 = sel_959176 + 8'h01;
  assign sel_959180 = array_index_959143 == array_index_948541 ? add_959179 : sel_959176;
  assign add_959183 = sel_959180 + 8'h01;
  assign sel_959184 = array_index_959143 == array_index_948547 ? add_959183 : sel_959180;
  assign add_959187 = sel_959184 + 8'h01;
  assign sel_959188 = array_index_959143 == array_index_948553 ? add_959187 : sel_959184;
  assign add_959191 = sel_959188 + 8'h01;
  assign sel_959192 = array_index_959143 == array_index_948559 ? add_959191 : sel_959188;
  assign add_959195 = sel_959192 + 8'h01;
  assign sel_959196 = array_index_959143 == array_index_948565 ? add_959195 : sel_959192;
  assign add_959199 = sel_959196 + 8'h01;
  assign sel_959200 = array_index_959143 == array_index_948571 ? add_959199 : sel_959196;
  assign add_959203 = sel_959200 + 8'h01;
  assign sel_959204 = array_index_959143 == array_index_948577 ? add_959203 : sel_959200;
  assign add_959207 = sel_959204 + 8'h01;
  assign sel_959208 = array_index_959143 == array_index_948583 ? add_959207 : sel_959204;
  assign add_959211 = sel_959208 + 8'h01;
  assign sel_959212 = array_index_959143 == array_index_948589 ? add_959211 : sel_959208;
  assign add_959215 = sel_959212 + 8'h01;
  assign sel_959216 = array_index_959143 == array_index_948595 ? add_959215 : sel_959212;
  assign add_959219 = sel_959216 + 8'h01;
  assign sel_959220 = array_index_959143 == array_index_948601 ? add_959219 : sel_959216;
  assign add_959223 = sel_959220 + 8'h01;
  assign sel_959224 = array_index_959143 == array_index_948607 ? add_959223 : sel_959220;
  assign add_959227 = sel_959224 + 8'h01;
  assign sel_959228 = array_index_959143 == array_index_948613 ? add_959227 : sel_959224;
  assign add_959231 = sel_959228 + 8'h01;
  assign sel_959232 = array_index_959143 == array_index_948619 ? add_959231 : sel_959228;
  assign add_959235 = sel_959232 + 8'h01;
  assign sel_959236 = array_index_959143 == array_index_948625 ? add_959235 : sel_959232;
  assign add_959239 = sel_959236 + 8'h01;
  assign sel_959240 = array_index_959143 == array_index_948631 ? add_959239 : sel_959236;
  assign add_959243 = sel_959240 + 8'h01;
  assign sel_959244 = array_index_959143 == array_index_948637 ? add_959243 : sel_959240;
  assign add_959247 = sel_959244 + 8'h01;
  assign sel_959248 = array_index_959143 == array_index_948643 ? add_959247 : sel_959244;
  assign add_959251 = sel_959248 + 8'h01;
  assign sel_959252 = array_index_959143 == array_index_948649 ? add_959251 : sel_959248;
  assign add_959255 = sel_959252 + 8'h01;
  assign sel_959256 = array_index_959143 == array_index_948655 ? add_959255 : sel_959252;
  assign add_959259 = sel_959256 + 8'h01;
  assign sel_959260 = array_index_959143 == array_index_948661 ? add_959259 : sel_959256;
  assign add_959263 = sel_959260 + 8'h01;
  assign sel_959264 = array_index_959143 == array_index_948667 ? add_959263 : sel_959260;
  assign add_959267 = sel_959264 + 8'h01;
  assign sel_959268 = array_index_959143 == array_index_948673 ? add_959267 : sel_959264;
  assign add_959271 = sel_959268 + 8'h01;
  assign sel_959272 = array_index_959143 == array_index_948679 ? add_959271 : sel_959268;
  assign add_959275 = sel_959272 + 8'h01;
  assign sel_959276 = array_index_959143 == array_index_948685 ? add_959275 : sel_959272;
  assign add_959279 = sel_959276 + 8'h01;
  assign sel_959280 = array_index_959143 == array_index_948691 ? add_959279 : sel_959276;
  assign add_959283 = sel_959280 + 8'h01;
  assign sel_959284 = array_index_959143 == array_index_948697 ? add_959283 : sel_959280;
  assign add_959287 = sel_959284 + 8'h01;
  assign sel_959288 = array_index_959143 == array_index_948703 ? add_959287 : sel_959284;
  assign add_959291 = sel_959288 + 8'h01;
  assign sel_959292 = array_index_959143 == array_index_948709 ? add_959291 : sel_959288;
  assign add_959295 = sel_959292 + 8'h01;
  assign sel_959296 = array_index_959143 == array_index_948715 ? add_959295 : sel_959292;
  assign add_959299 = sel_959296 + 8'h01;
  assign sel_959300 = array_index_959143 == array_index_948721 ? add_959299 : sel_959296;
  assign add_959303 = sel_959300 + 8'h01;
  assign sel_959304 = array_index_959143 == array_index_948727 ? add_959303 : sel_959300;
  assign add_959307 = sel_959304 + 8'h01;
  assign sel_959308 = array_index_959143 == array_index_948733 ? add_959307 : sel_959304;
  assign add_959311 = sel_959308 + 8'h01;
  assign sel_959312 = array_index_959143 == array_index_948739 ? add_959311 : sel_959308;
  assign add_959315 = sel_959312 + 8'h01;
  assign sel_959316 = array_index_959143 == array_index_948745 ? add_959315 : sel_959312;
  assign add_959319 = sel_959316 + 8'h01;
  assign sel_959320 = array_index_959143 == array_index_948751 ? add_959319 : sel_959316;
  assign add_959323 = sel_959320 + 8'h01;
  assign sel_959324 = array_index_959143 == array_index_948757 ? add_959323 : sel_959320;
  assign add_959327 = sel_959324 + 8'h01;
  assign sel_959328 = array_index_959143 == array_index_948763 ? add_959327 : sel_959324;
  assign add_959331 = sel_959328 + 8'h01;
  assign sel_959332 = array_index_959143 == array_index_948769 ? add_959331 : sel_959328;
  assign add_959335 = sel_959332 + 8'h01;
  assign sel_959336 = array_index_959143 == array_index_948775 ? add_959335 : sel_959332;
  assign add_959339 = sel_959336 + 8'h01;
  assign sel_959340 = array_index_959143 == array_index_948781 ? add_959339 : sel_959336;
  assign add_959343 = sel_959340 + 8'h01;
  assign sel_959344 = array_index_959143 == array_index_948787 ? add_959343 : sel_959340;
  assign add_959347 = sel_959344 + 8'h01;
  assign sel_959348 = array_index_959143 == array_index_948793 ? add_959347 : sel_959344;
  assign add_959351 = sel_959348 + 8'h01;
  assign sel_959352 = array_index_959143 == array_index_948799 ? add_959351 : sel_959348;
  assign add_959355 = sel_959352 + 8'h01;
  assign sel_959356 = array_index_959143 == array_index_948805 ? add_959355 : sel_959352;
  assign add_959359 = sel_959356 + 8'h01;
  assign sel_959360 = array_index_959143 == array_index_948811 ? add_959359 : sel_959356;
  assign add_959363 = sel_959360 + 8'h01;
  assign sel_959364 = array_index_959143 == array_index_948817 ? add_959363 : sel_959360;
  assign add_959367 = sel_959364 + 8'h01;
  assign sel_959368 = array_index_959143 == array_index_948823 ? add_959367 : sel_959364;
  assign add_959371 = sel_959368 + 8'h01;
  assign sel_959372 = array_index_959143 == array_index_948829 ? add_959371 : sel_959368;
  assign add_959375 = sel_959372 + 8'h01;
  assign sel_959376 = array_index_959143 == array_index_948835 ? add_959375 : sel_959372;
  assign add_959379 = sel_959376 + 8'h01;
  assign sel_959380 = array_index_959143 == array_index_948841 ? add_959379 : sel_959376;
  assign add_959383 = sel_959380 + 8'h01;
  assign sel_959384 = array_index_959143 == array_index_948847 ? add_959383 : sel_959380;
  assign add_959387 = sel_959384 + 8'h01;
  assign sel_959388 = array_index_959143 == array_index_948853 ? add_959387 : sel_959384;
  assign add_959391 = sel_959388 + 8'h01;
  assign sel_959392 = array_index_959143 == array_index_948859 ? add_959391 : sel_959388;
  assign add_959395 = sel_959392 + 8'h01;
  assign sel_959396 = array_index_959143 == array_index_948865 ? add_959395 : sel_959392;
  assign add_959399 = sel_959396 + 8'h01;
  assign sel_959400 = array_index_959143 == array_index_948871 ? add_959399 : sel_959396;
  assign add_959403 = sel_959400 + 8'h01;
  assign sel_959404 = array_index_959143 == array_index_948877 ? add_959403 : sel_959400;
  assign add_959407 = sel_959404 + 8'h01;
  assign sel_959408 = array_index_959143 == array_index_948883 ? add_959407 : sel_959404;
  assign add_959411 = sel_959408 + 8'h01;
  assign sel_959412 = array_index_959143 == array_index_948889 ? add_959411 : sel_959408;
  assign add_959415 = sel_959412 + 8'h01;
  assign sel_959416 = array_index_959143 == array_index_948895 ? add_959415 : sel_959412;
  assign add_959419 = sel_959416 + 8'h01;
  assign sel_959420 = array_index_959143 == array_index_948901 ? add_959419 : sel_959416;
  assign add_959423 = sel_959420 + 8'h01;
  assign sel_959424 = array_index_959143 == array_index_948907 ? add_959423 : sel_959420;
  assign add_959427 = sel_959424 + 8'h01;
  assign sel_959428 = array_index_959143 == array_index_948913 ? add_959427 : sel_959424;
  assign add_959431 = sel_959428 + 8'h01;
  assign sel_959432 = array_index_959143 == array_index_948919 ? add_959431 : sel_959428;
  assign add_959435 = sel_959432 + 8'h01;
  assign sel_959436 = array_index_959143 == array_index_948925 ? add_959435 : sel_959432;
  assign add_959439 = sel_959436 + 8'h01;
  assign sel_959440 = array_index_959143 == array_index_948931 ? add_959439 : sel_959436;
  assign add_959443 = sel_959440 + 8'h01;
  assign sel_959444 = array_index_959143 == array_index_948937 ? add_959443 : sel_959440;
  assign add_959447 = sel_959444 + 8'h01;
  assign sel_959448 = array_index_959143 == array_index_948943 ? add_959447 : sel_959444;
  assign add_959451 = sel_959448 + 8'h01;
  assign sel_959452 = array_index_959143 == array_index_948949 ? add_959451 : sel_959448;
  assign add_959455 = sel_959452 + 8'h01;
  assign sel_959456 = array_index_959143 == array_index_948955 ? add_959455 : sel_959452;
  assign add_959459 = sel_959456 + 8'h01;
  assign sel_959460 = array_index_959143 == array_index_948961 ? add_959459 : sel_959456;
  assign add_959463 = sel_959460 + 8'h01;
  assign sel_959464 = array_index_959143 == array_index_948967 ? add_959463 : sel_959460;
  assign add_959467 = sel_959464 + 8'h01;
  assign sel_959468 = array_index_959143 == array_index_948973 ? add_959467 : sel_959464;
  assign add_959471 = sel_959468 + 8'h01;
  assign sel_959472 = array_index_959143 == array_index_948979 ? add_959471 : sel_959468;
  assign add_959475 = sel_959472 + 8'h01;
  assign sel_959476 = array_index_959143 == array_index_948985 ? add_959475 : sel_959472;
  assign add_959479 = sel_959476 + 8'h01;
  assign sel_959480 = array_index_959143 == array_index_948991 ? add_959479 : sel_959476;
  assign add_959483 = sel_959480 + 8'h01;
  assign sel_959484 = array_index_959143 == array_index_948997 ? add_959483 : sel_959480;
  assign add_959487 = sel_959484 + 8'h01;
  assign sel_959488 = array_index_959143 == array_index_949003 ? add_959487 : sel_959484;
  assign add_959491 = sel_959488 + 8'h01;
  assign sel_959492 = array_index_959143 == array_index_949009 ? add_959491 : sel_959488;
  assign add_959495 = sel_959492 + 8'h01;
  assign sel_959496 = array_index_959143 == array_index_949015 ? add_959495 : sel_959492;
  assign add_959499 = sel_959496 + 8'h01;
  assign sel_959500 = array_index_959143 == array_index_949021 ? add_959499 : sel_959496;
  assign add_959503 = sel_959500 + 8'h01;
  assign sel_959504 = array_index_959143 == array_index_949027 ? add_959503 : sel_959500;
  assign add_959507 = sel_959504 + 8'h01;
  assign sel_959508 = array_index_959143 == array_index_949033 ? add_959507 : sel_959504;
  assign add_959511 = sel_959508 + 8'h01;
  assign sel_959512 = array_index_959143 == array_index_949039 ? add_959511 : sel_959508;
  assign add_959515 = sel_959512 + 8'h01;
  assign sel_959516 = array_index_959143 == array_index_949045 ? add_959515 : sel_959512;
  assign add_959519 = sel_959516 + 8'h01;
  assign sel_959520 = array_index_959143 == array_index_949051 ? add_959519 : sel_959516;
  assign add_959523 = sel_959520 + 8'h01;
  assign sel_959524 = array_index_959143 == array_index_949057 ? add_959523 : sel_959520;
  assign add_959527 = sel_959524 + 8'h01;
  assign sel_959528 = array_index_959143 == array_index_949063 ? add_959527 : sel_959524;
  assign add_959531 = sel_959528 + 8'h01;
  assign sel_959532 = array_index_959143 == array_index_949069 ? add_959531 : sel_959528;
  assign add_959535 = sel_959532 + 8'h01;
  assign sel_959536 = array_index_959143 == array_index_949075 ? add_959535 : sel_959532;
  assign add_959539 = sel_959536 + 8'h01;
  assign sel_959540 = array_index_959143 == array_index_949081 ? add_959539 : sel_959536;
  assign add_959544 = sel_959540 + 8'h01;
  assign array_index_959545 = set1_unflattened[7'h1b];
  assign sel_959546 = array_index_959143 == array_index_949087 ? add_959544 : sel_959540;
  assign add_959549 = sel_959546 + 8'h01;
  assign sel_959550 = array_index_959545 == array_index_948483 ? add_959549 : sel_959546;
  assign add_959553 = sel_959550 + 8'h01;
  assign sel_959554 = array_index_959545 == array_index_948487 ? add_959553 : sel_959550;
  assign add_959557 = sel_959554 + 8'h01;
  assign sel_959558 = array_index_959545 == array_index_948495 ? add_959557 : sel_959554;
  assign add_959561 = sel_959558 + 8'h01;
  assign sel_959562 = array_index_959545 == array_index_948503 ? add_959561 : sel_959558;
  assign add_959565 = sel_959562 + 8'h01;
  assign sel_959566 = array_index_959545 == array_index_948511 ? add_959565 : sel_959562;
  assign add_959569 = sel_959566 + 8'h01;
  assign sel_959570 = array_index_959545 == array_index_948519 ? add_959569 : sel_959566;
  assign add_959573 = sel_959570 + 8'h01;
  assign sel_959574 = array_index_959545 == array_index_948527 ? add_959573 : sel_959570;
  assign add_959577 = sel_959574 + 8'h01;
  assign sel_959578 = array_index_959545 == array_index_948535 ? add_959577 : sel_959574;
  assign add_959581 = sel_959578 + 8'h01;
  assign sel_959582 = array_index_959545 == array_index_948541 ? add_959581 : sel_959578;
  assign add_959585 = sel_959582 + 8'h01;
  assign sel_959586 = array_index_959545 == array_index_948547 ? add_959585 : sel_959582;
  assign add_959589 = sel_959586 + 8'h01;
  assign sel_959590 = array_index_959545 == array_index_948553 ? add_959589 : sel_959586;
  assign add_959593 = sel_959590 + 8'h01;
  assign sel_959594 = array_index_959545 == array_index_948559 ? add_959593 : sel_959590;
  assign add_959597 = sel_959594 + 8'h01;
  assign sel_959598 = array_index_959545 == array_index_948565 ? add_959597 : sel_959594;
  assign add_959601 = sel_959598 + 8'h01;
  assign sel_959602 = array_index_959545 == array_index_948571 ? add_959601 : sel_959598;
  assign add_959605 = sel_959602 + 8'h01;
  assign sel_959606 = array_index_959545 == array_index_948577 ? add_959605 : sel_959602;
  assign add_959609 = sel_959606 + 8'h01;
  assign sel_959610 = array_index_959545 == array_index_948583 ? add_959609 : sel_959606;
  assign add_959613 = sel_959610 + 8'h01;
  assign sel_959614 = array_index_959545 == array_index_948589 ? add_959613 : sel_959610;
  assign add_959617 = sel_959614 + 8'h01;
  assign sel_959618 = array_index_959545 == array_index_948595 ? add_959617 : sel_959614;
  assign add_959621 = sel_959618 + 8'h01;
  assign sel_959622 = array_index_959545 == array_index_948601 ? add_959621 : sel_959618;
  assign add_959625 = sel_959622 + 8'h01;
  assign sel_959626 = array_index_959545 == array_index_948607 ? add_959625 : sel_959622;
  assign add_959629 = sel_959626 + 8'h01;
  assign sel_959630 = array_index_959545 == array_index_948613 ? add_959629 : sel_959626;
  assign add_959633 = sel_959630 + 8'h01;
  assign sel_959634 = array_index_959545 == array_index_948619 ? add_959633 : sel_959630;
  assign add_959637 = sel_959634 + 8'h01;
  assign sel_959638 = array_index_959545 == array_index_948625 ? add_959637 : sel_959634;
  assign add_959641 = sel_959638 + 8'h01;
  assign sel_959642 = array_index_959545 == array_index_948631 ? add_959641 : sel_959638;
  assign add_959645 = sel_959642 + 8'h01;
  assign sel_959646 = array_index_959545 == array_index_948637 ? add_959645 : sel_959642;
  assign add_959649 = sel_959646 + 8'h01;
  assign sel_959650 = array_index_959545 == array_index_948643 ? add_959649 : sel_959646;
  assign add_959653 = sel_959650 + 8'h01;
  assign sel_959654 = array_index_959545 == array_index_948649 ? add_959653 : sel_959650;
  assign add_959657 = sel_959654 + 8'h01;
  assign sel_959658 = array_index_959545 == array_index_948655 ? add_959657 : sel_959654;
  assign add_959661 = sel_959658 + 8'h01;
  assign sel_959662 = array_index_959545 == array_index_948661 ? add_959661 : sel_959658;
  assign add_959665 = sel_959662 + 8'h01;
  assign sel_959666 = array_index_959545 == array_index_948667 ? add_959665 : sel_959662;
  assign add_959669 = sel_959666 + 8'h01;
  assign sel_959670 = array_index_959545 == array_index_948673 ? add_959669 : sel_959666;
  assign add_959673 = sel_959670 + 8'h01;
  assign sel_959674 = array_index_959545 == array_index_948679 ? add_959673 : sel_959670;
  assign add_959677 = sel_959674 + 8'h01;
  assign sel_959678 = array_index_959545 == array_index_948685 ? add_959677 : sel_959674;
  assign add_959681 = sel_959678 + 8'h01;
  assign sel_959682 = array_index_959545 == array_index_948691 ? add_959681 : sel_959678;
  assign add_959685 = sel_959682 + 8'h01;
  assign sel_959686 = array_index_959545 == array_index_948697 ? add_959685 : sel_959682;
  assign add_959689 = sel_959686 + 8'h01;
  assign sel_959690 = array_index_959545 == array_index_948703 ? add_959689 : sel_959686;
  assign add_959693 = sel_959690 + 8'h01;
  assign sel_959694 = array_index_959545 == array_index_948709 ? add_959693 : sel_959690;
  assign add_959697 = sel_959694 + 8'h01;
  assign sel_959698 = array_index_959545 == array_index_948715 ? add_959697 : sel_959694;
  assign add_959701 = sel_959698 + 8'h01;
  assign sel_959702 = array_index_959545 == array_index_948721 ? add_959701 : sel_959698;
  assign add_959705 = sel_959702 + 8'h01;
  assign sel_959706 = array_index_959545 == array_index_948727 ? add_959705 : sel_959702;
  assign add_959709 = sel_959706 + 8'h01;
  assign sel_959710 = array_index_959545 == array_index_948733 ? add_959709 : sel_959706;
  assign add_959713 = sel_959710 + 8'h01;
  assign sel_959714 = array_index_959545 == array_index_948739 ? add_959713 : sel_959710;
  assign add_959717 = sel_959714 + 8'h01;
  assign sel_959718 = array_index_959545 == array_index_948745 ? add_959717 : sel_959714;
  assign add_959721 = sel_959718 + 8'h01;
  assign sel_959722 = array_index_959545 == array_index_948751 ? add_959721 : sel_959718;
  assign add_959725 = sel_959722 + 8'h01;
  assign sel_959726 = array_index_959545 == array_index_948757 ? add_959725 : sel_959722;
  assign add_959729 = sel_959726 + 8'h01;
  assign sel_959730 = array_index_959545 == array_index_948763 ? add_959729 : sel_959726;
  assign add_959733 = sel_959730 + 8'h01;
  assign sel_959734 = array_index_959545 == array_index_948769 ? add_959733 : sel_959730;
  assign add_959737 = sel_959734 + 8'h01;
  assign sel_959738 = array_index_959545 == array_index_948775 ? add_959737 : sel_959734;
  assign add_959741 = sel_959738 + 8'h01;
  assign sel_959742 = array_index_959545 == array_index_948781 ? add_959741 : sel_959738;
  assign add_959745 = sel_959742 + 8'h01;
  assign sel_959746 = array_index_959545 == array_index_948787 ? add_959745 : sel_959742;
  assign add_959749 = sel_959746 + 8'h01;
  assign sel_959750 = array_index_959545 == array_index_948793 ? add_959749 : sel_959746;
  assign add_959753 = sel_959750 + 8'h01;
  assign sel_959754 = array_index_959545 == array_index_948799 ? add_959753 : sel_959750;
  assign add_959757 = sel_959754 + 8'h01;
  assign sel_959758 = array_index_959545 == array_index_948805 ? add_959757 : sel_959754;
  assign add_959761 = sel_959758 + 8'h01;
  assign sel_959762 = array_index_959545 == array_index_948811 ? add_959761 : sel_959758;
  assign add_959765 = sel_959762 + 8'h01;
  assign sel_959766 = array_index_959545 == array_index_948817 ? add_959765 : sel_959762;
  assign add_959769 = sel_959766 + 8'h01;
  assign sel_959770 = array_index_959545 == array_index_948823 ? add_959769 : sel_959766;
  assign add_959773 = sel_959770 + 8'h01;
  assign sel_959774 = array_index_959545 == array_index_948829 ? add_959773 : sel_959770;
  assign add_959777 = sel_959774 + 8'h01;
  assign sel_959778 = array_index_959545 == array_index_948835 ? add_959777 : sel_959774;
  assign add_959781 = sel_959778 + 8'h01;
  assign sel_959782 = array_index_959545 == array_index_948841 ? add_959781 : sel_959778;
  assign add_959785 = sel_959782 + 8'h01;
  assign sel_959786 = array_index_959545 == array_index_948847 ? add_959785 : sel_959782;
  assign add_959789 = sel_959786 + 8'h01;
  assign sel_959790 = array_index_959545 == array_index_948853 ? add_959789 : sel_959786;
  assign add_959793 = sel_959790 + 8'h01;
  assign sel_959794 = array_index_959545 == array_index_948859 ? add_959793 : sel_959790;
  assign add_959797 = sel_959794 + 8'h01;
  assign sel_959798 = array_index_959545 == array_index_948865 ? add_959797 : sel_959794;
  assign add_959801 = sel_959798 + 8'h01;
  assign sel_959802 = array_index_959545 == array_index_948871 ? add_959801 : sel_959798;
  assign add_959805 = sel_959802 + 8'h01;
  assign sel_959806 = array_index_959545 == array_index_948877 ? add_959805 : sel_959802;
  assign add_959809 = sel_959806 + 8'h01;
  assign sel_959810 = array_index_959545 == array_index_948883 ? add_959809 : sel_959806;
  assign add_959813 = sel_959810 + 8'h01;
  assign sel_959814 = array_index_959545 == array_index_948889 ? add_959813 : sel_959810;
  assign add_959817 = sel_959814 + 8'h01;
  assign sel_959818 = array_index_959545 == array_index_948895 ? add_959817 : sel_959814;
  assign add_959821 = sel_959818 + 8'h01;
  assign sel_959822 = array_index_959545 == array_index_948901 ? add_959821 : sel_959818;
  assign add_959825 = sel_959822 + 8'h01;
  assign sel_959826 = array_index_959545 == array_index_948907 ? add_959825 : sel_959822;
  assign add_959829 = sel_959826 + 8'h01;
  assign sel_959830 = array_index_959545 == array_index_948913 ? add_959829 : sel_959826;
  assign add_959833 = sel_959830 + 8'h01;
  assign sel_959834 = array_index_959545 == array_index_948919 ? add_959833 : sel_959830;
  assign add_959837 = sel_959834 + 8'h01;
  assign sel_959838 = array_index_959545 == array_index_948925 ? add_959837 : sel_959834;
  assign add_959841 = sel_959838 + 8'h01;
  assign sel_959842 = array_index_959545 == array_index_948931 ? add_959841 : sel_959838;
  assign add_959845 = sel_959842 + 8'h01;
  assign sel_959846 = array_index_959545 == array_index_948937 ? add_959845 : sel_959842;
  assign add_959849 = sel_959846 + 8'h01;
  assign sel_959850 = array_index_959545 == array_index_948943 ? add_959849 : sel_959846;
  assign add_959853 = sel_959850 + 8'h01;
  assign sel_959854 = array_index_959545 == array_index_948949 ? add_959853 : sel_959850;
  assign add_959857 = sel_959854 + 8'h01;
  assign sel_959858 = array_index_959545 == array_index_948955 ? add_959857 : sel_959854;
  assign add_959861 = sel_959858 + 8'h01;
  assign sel_959862 = array_index_959545 == array_index_948961 ? add_959861 : sel_959858;
  assign add_959865 = sel_959862 + 8'h01;
  assign sel_959866 = array_index_959545 == array_index_948967 ? add_959865 : sel_959862;
  assign add_959869 = sel_959866 + 8'h01;
  assign sel_959870 = array_index_959545 == array_index_948973 ? add_959869 : sel_959866;
  assign add_959873 = sel_959870 + 8'h01;
  assign sel_959874 = array_index_959545 == array_index_948979 ? add_959873 : sel_959870;
  assign add_959877 = sel_959874 + 8'h01;
  assign sel_959878 = array_index_959545 == array_index_948985 ? add_959877 : sel_959874;
  assign add_959881 = sel_959878 + 8'h01;
  assign sel_959882 = array_index_959545 == array_index_948991 ? add_959881 : sel_959878;
  assign add_959885 = sel_959882 + 8'h01;
  assign sel_959886 = array_index_959545 == array_index_948997 ? add_959885 : sel_959882;
  assign add_959889 = sel_959886 + 8'h01;
  assign sel_959890 = array_index_959545 == array_index_949003 ? add_959889 : sel_959886;
  assign add_959893 = sel_959890 + 8'h01;
  assign sel_959894 = array_index_959545 == array_index_949009 ? add_959893 : sel_959890;
  assign add_959897 = sel_959894 + 8'h01;
  assign sel_959898 = array_index_959545 == array_index_949015 ? add_959897 : sel_959894;
  assign add_959901 = sel_959898 + 8'h01;
  assign sel_959902 = array_index_959545 == array_index_949021 ? add_959901 : sel_959898;
  assign add_959905 = sel_959902 + 8'h01;
  assign sel_959906 = array_index_959545 == array_index_949027 ? add_959905 : sel_959902;
  assign add_959909 = sel_959906 + 8'h01;
  assign sel_959910 = array_index_959545 == array_index_949033 ? add_959909 : sel_959906;
  assign add_959913 = sel_959910 + 8'h01;
  assign sel_959914 = array_index_959545 == array_index_949039 ? add_959913 : sel_959910;
  assign add_959917 = sel_959914 + 8'h01;
  assign sel_959918 = array_index_959545 == array_index_949045 ? add_959917 : sel_959914;
  assign add_959921 = sel_959918 + 8'h01;
  assign sel_959922 = array_index_959545 == array_index_949051 ? add_959921 : sel_959918;
  assign add_959925 = sel_959922 + 8'h01;
  assign sel_959926 = array_index_959545 == array_index_949057 ? add_959925 : sel_959922;
  assign add_959929 = sel_959926 + 8'h01;
  assign sel_959930 = array_index_959545 == array_index_949063 ? add_959929 : sel_959926;
  assign add_959933 = sel_959930 + 8'h01;
  assign sel_959934 = array_index_959545 == array_index_949069 ? add_959933 : sel_959930;
  assign add_959937 = sel_959934 + 8'h01;
  assign sel_959938 = array_index_959545 == array_index_949075 ? add_959937 : sel_959934;
  assign add_959941 = sel_959938 + 8'h01;
  assign sel_959942 = array_index_959545 == array_index_949081 ? add_959941 : sel_959938;
  assign add_959946 = sel_959942 + 8'h01;
  assign array_index_959947 = set1_unflattened[7'h1c];
  assign sel_959948 = array_index_959545 == array_index_949087 ? add_959946 : sel_959942;
  assign add_959951 = sel_959948 + 8'h01;
  assign sel_959952 = array_index_959947 == array_index_948483 ? add_959951 : sel_959948;
  assign add_959955 = sel_959952 + 8'h01;
  assign sel_959956 = array_index_959947 == array_index_948487 ? add_959955 : sel_959952;
  assign add_959959 = sel_959956 + 8'h01;
  assign sel_959960 = array_index_959947 == array_index_948495 ? add_959959 : sel_959956;
  assign add_959963 = sel_959960 + 8'h01;
  assign sel_959964 = array_index_959947 == array_index_948503 ? add_959963 : sel_959960;
  assign add_959967 = sel_959964 + 8'h01;
  assign sel_959968 = array_index_959947 == array_index_948511 ? add_959967 : sel_959964;
  assign add_959971 = sel_959968 + 8'h01;
  assign sel_959972 = array_index_959947 == array_index_948519 ? add_959971 : sel_959968;
  assign add_959975 = sel_959972 + 8'h01;
  assign sel_959976 = array_index_959947 == array_index_948527 ? add_959975 : sel_959972;
  assign add_959979 = sel_959976 + 8'h01;
  assign sel_959980 = array_index_959947 == array_index_948535 ? add_959979 : sel_959976;
  assign add_959983 = sel_959980 + 8'h01;
  assign sel_959984 = array_index_959947 == array_index_948541 ? add_959983 : sel_959980;
  assign add_959987 = sel_959984 + 8'h01;
  assign sel_959988 = array_index_959947 == array_index_948547 ? add_959987 : sel_959984;
  assign add_959991 = sel_959988 + 8'h01;
  assign sel_959992 = array_index_959947 == array_index_948553 ? add_959991 : sel_959988;
  assign add_959995 = sel_959992 + 8'h01;
  assign sel_959996 = array_index_959947 == array_index_948559 ? add_959995 : sel_959992;
  assign add_959999 = sel_959996 + 8'h01;
  assign sel_960000 = array_index_959947 == array_index_948565 ? add_959999 : sel_959996;
  assign add_960003 = sel_960000 + 8'h01;
  assign sel_960004 = array_index_959947 == array_index_948571 ? add_960003 : sel_960000;
  assign add_960007 = sel_960004 + 8'h01;
  assign sel_960008 = array_index_959947 == array_index_948577 ? add_960007 : sel_960004;
  assign add_960011 = sel_960008 + 8'h01;
  assign sel_960012 = array_index_959947 == array_index_948583 ? add_960011 : sel_960008;
  assign add_960015 = sel_960012 + 8'h01;
  assign sel_960016 = array_index_959947 == array_index_948589 ? add_960015 : sel_960012;
  assign add_960019 = sel_960016 + 8'h01;
  assign sel_960020 = array_index_959947 == array_index_948595 ? add_960019 : sel_960016;
  assign add_960023 = sel_960020 + 8'h01;
  assign sel_960024 = array_index_959947 == array_index_948601 ? add_960023 : sel_960020;
  assign add_960027 = sel_960024 + 8'h01;
  assign sel_960028 = array_index_959947 == array_index_948607 ? add_960027 : sel_960024;
  assign add_960031 = sel_960028 + 8'h01;
  assign sel_960032 = array_index_959947 == array_index_948613 ? add_960031 : sel_960028;
  assign add_960035 = sel_960032 + 8'h01;
  assign sel_960036 = array_index_959947 == array_index_948619 ? add_960035 : sel_960032;
  assign add_960039 = sel_960036 + 8'h01;
  assign sel_960040 = array_index_959947 == array_index_948625 ? add_960039 : sel_960036;
  assign add_960043 = sel_960040 + 8'h01;
  assign sel_960044 = array_index_959947 == array_index_948631 ? add_960043 : sel_960040;
  assign add_960047 = sel_960044 + 8'h01;
  assign sel_960048 = array_index_959947 == array_index_948637 ? add_960047 : sel_960044;
  assign add_960051 = sel_960048 + 8'h01;
  assign sel_960052 = array_index_959947 == array_index_948643 ? add_960051 : sel_960048;
  assign add_960055 = sel_960052 + 8'h01;
  assign sel_960056 = array_index_959947 == array_index_948649 ? add_960055 : sel_960052;
  assign add_960059 = sel_960056 + 8'h01;
  assign sel_960060 = array_index_959947 == array_index_948655 ? add_960059 : sel_960056;
  assign add_960063 = sel_960060 + 8'h01;
  assign sel_960064 = array_index_959947 == array_index_948661 ? add_960063 : sel_960060;
  assign add_960067 = sel_960064 + 8'h01;
  assign sel_960068 = array_index_959947 == array_index_948667 ? add_960067 : sel_960064;
  assign add_960071 = sel_960068 + 8'h01;
  assign sel_960072 = array_index_959947 == array_index_948673 ? add_960071 : sel_960068;
  assign add_960075 = sel_960072 + 8'h01;
  assign sel_960076 = array_index_959947 == array_index_948679 ? add_960075 : sel_960072;
  assign add_960079 = sel_960076 + 8'h01;
  assign sel_960080 = array_index_959947 == array_index_948685 ? add_960079 : sel_960076;
  assign add_960083 = sel_960080 + 8'h01;
  assign sel_960084 = array_index_959947 == array_index_948691 ? add_960083 : sel_960080;
  assign add_960087 = sel_960084 + 8'h01;
  assign sel_960088 = array_index_959947 == array_index_948697 ? add_960087 : sel_960084;
  assign add_960091 = sel_960088 + 8'h01;
  assign sel_960092 = array_index_959947 == array_index_948703 ? add_960091 : sel_960088;
  assign add_960095 = sel_960092 + 8'h01;
  assign sel_960096 = array_index_959947 == array_index_948709 ? add_960095 : sel_960092;
  assign add_960099 = sel_960096 + 8'h01;
  assign sel_960100 = array_index_959947 == array_index_948715 ? add_960099 : sel_960096;
  assign add_960103 = sel_960100 + 8'h01;
  assign sel_960104 = array_index_959947 == array_index_948721 ? add_960103 : sel_960100;
  assign add_960107 = sel_960104 + 8'h01;
  assign sel_960108 = array_index_959947 == array_index_948727 ? add_960107 : sel_960104;
  assign add_960111 = sel_960108 + 8'h01;
  assign sel_960112 = array_index_959947 == array_index_948733 ? add_960111 : sel_960108;
  assign add_960115 = sel_960112 + 8'h01;
  assign sel_960116 = array_index_959947 == array_index_948739 ? add_960115 : sel_960112;
  assign add_960119 = sel_960116 + 8'h01;
  assign sel_960120 = array_index_959947 == array_index_948745 ? add_960119 : sel_960116;
  assign add_960123 = sel_960120 + 8'h01;
  assign sel_960124 = array_index_959947 == array_index_948751 ? add_960123 : sel_960120;
  assign add_960127 = sel_960124 + 8'h01;
  assign sel_960128 = array_index_959947 == array_index_948757 ? add_960127 : sel_960124;
  assign add_960131 = sel_960128 + 8'h01;
  assign sel_960132 = array_index_959947 == array_index_948763 ? add_960131 : sel_960128;
  assign add_960135 = sel_960132 + 8'h01;
  assign sel_960136 = array_index_959947 == array_index_948769 ? add_960135 : sel_960132;
  assign add_960139 = sel_960136 + 8'h01;
  assign sel_960140 = array_index_959947 == array_index_948775 ? add_960139 : sel_960136;
  assign add_960143 = sel_960140 + 8'h01;
  assign sel_960144 = array_index_959947 == array_index_948781 ? add_960143 : sel_960140;
  assign add_960147 = sel_960144 + 8'h01;
  assign sel_960148 = array_index_959947 == array_index_948787 ? add_960147 : sel_960144;
  assign add_960151 = sel_960148 + 8'h01;
  assign sel_960152 = array_index_959947 == array_index_948793 ? add_960151 : sel_960148;
  assign add_960155 = sel_960152 + 8'h01;
  assign sel_960156 = array_index_959947 == array_index_948799 ? add_960155 : sel_960152;
  assign add_960159 = sel_960156 + 8'h01;
  assign sel_960160 = array_index_959947 == array_index_948805 ? add_960159 : sel_960156;
  assign add_960163 = sel_960160 + 8'h01;
  assign sel_960164 = array_index_959947 == array_index_948811 ? add_960163 : sel_960160;
  assign add_960167 = sel_960164 + 8'h01;
  assign sel_960168 = array_index_959947 == array_index_948817 ? add_960167 : sel_960164;
  assign add_960171 = sel_960168 + 8'h01;
  assign sel_960172 = array_index_959947 == array_index_948823 ? add_960171 : sel_960168;
  assign add_960175 = sel_960172 + 8'h01;
  assign sel_960176 = array_index_959947 == array_index_948829 ? add_960175 : sel_960172;
  assign add_960179 = sel_960176 + 8'h01;
  assign sel_960180 = array_index_959947 == array_index_948835 ? add_960179 : sel_960176;
  assign add_960183 = sel_960180 + 8'h01;
  assign sel_960184 = array_index_959947 == array_index_948841 ? add_960183 : sel_960180;
  assign add_960187 = sel_960184 + 8'h01;
  assign sel_960188 = array_index_959947 == array_index_948847 ? add_960187 : sel_960184;
  assign add_960191 = sel_960188 + 8'h01;
  assign sel_960192 = array_index_959947 == array_index_948853 ? add_960191 : sel_960188;
  assign add_960195 = sel_960192 + 8'h01;
  assign sel_960196 = array_index_959947 == array_index_948859 ? add_960195 : sel_960192;
  assign add_960199 = sel_960196 + 8'h01;
  assign sel_960200 = array_index_959947 == array_index_948865 ? add_960199 : sel_960196;
  assign add_960203 = sel_960200 + 8'h01;
  assign sel_960204 = array_index_959947 == array_index_948871 ? add_960203 : sel_960200;
  assign add_960207 = sel_960204 + 8'h01;
  assign sel_960208 = array_index_959947 == array_index_948877 ? add_960207 : sel_960204;
  assign add_960211 = sel_960208 + 8'h01;
  assign sel_960212 = array_index_959947 == array_index_948883 ? add_960211 : sel_960208;
  assign add_960215 = sel_960212 + 8'h01;
  assign sel_960216 = array_index_959947 == array_index_948889 ? add_960215 : sel_960212;
  assign add_960219 = sel_960216 + 8'h01;
  assign sel_960220 = array_index_959947 == array_index_948895 ? add_960219 : sel_960216;
  assign add_960223 = sel_960220 + 8'h01;
  assign sel_960224 = array_index_959947 == array_index_948901 ? add_960223 : sel_960220;
  assign add_960227 = sel_960224 + 8'h01;
  assign sel_960228 = array_index_959947 == array_index_948907 ? add_960227 : sel_960224;
  assign add_960231 = sel_960228 + 8'h01;
  assign sel_960232 = array_index_959947 == array_index_948913 ? add_960231 : sel_960228;
  assign add_960235 = sel_960232 + 8'h01;
  assign sel_960236 = array_index_959947 == array_index_948919 ? add_960235 : sel_960232;
  assign add_960239 = sel_960236 + 8'h01;
  assign sel_960240 = array_index_959947 == array_index_948925 ? add_960239 : sel_960236;
  assign add_960243 = sel_960240 + 8'h01;
  assign sel_960244 = array_index_959947 == array_index_948931 ? add_960243 : sel_960240;
  assign add_960247 = sel_960244 + 8'h01;
  assign sel_960248 = array_index_959947 == array_index_948937 ? add_960247 : sel_960244;
  assign add_960251 = sel_960248 + 8'h01;
  assign sel_960252 = array_index_959947 == array_index_948943 ? add_960251 : sel_960248;
  assign add_960255 = sel_960252 + 8'h01;
  assign sel_960256 = array_index_959947 == array_index_948949 ? add_960255 : sel_960252;
  assign add_960259 = sel_960256 + 8'h01;
  assign sel_960260 = array_index_959947 == array_index_948955 ? add_960259 : sel_960256;
  assign add_960263 = sel_960260 + 8'h01;
  assign sel_960264 = array_index_959947 == array_index_948961 ? add_960263 : sel_960260;
  assign add_960267 = sel_960264 + 8'h01;
  assign sel_960268 = array_index_959947 == array_index_948967 ? add_960267 : sel_960264;
  assign add_960271 = sel_960268 + 8'h01;
  assign sel_960272 = array_index_959947 == array_index_948973 ? add_960271 : sel_960268;
  assign add_960275 = sel_960272 + 8'h01;
  assign sel_960276 = array_index_959947 == array_index_948979 ? add_960275 : sel_960272;
  assign add_960279 = sel_960276 + 8'h01;
  assign sel_960280 = array_index_959947 == array_index_948985 ? add_960279 : sel_960276;
  assign add_960283 = sel_960280 + 8'h01;
  assign sel_960284 = array_index_959947 == array_index_948991 ? add_960283 : sel_960280;
  assign add_960287 = sel_960284 + 8'h01;
  assign sel_960288 = array_index_959947 == array_index_948997 ? add_960287 : sel_960284;
  assign add_960291 = sel_960288 + 8'h01;
  assign sel_960292 = array_index_959947 == array_index_949003 ? add_960291 : sel_960288;
  assign add_960295 = sel_960292 + 8'h01;
  assign sel_960296 = array_index_959947 == array_index_949009 ? add_960295 : sel_960292;
  assign add_960299 = sel_960296 + 8'h01;
  assign sel_960300 = array_index_959947 == array_index_949015 ? add_960299 : sel_960296;
  assign add_960303 = sel_960300 + 8'h01;
  assign sel_960304 = array_index_959947 == array_index_949021 ? add_960303 : sel_960300;
  assign add_960307 = sel_960304 + 8'h01;
  assign sel_960308 = array_index_959947 == array_index_949027 ? add_960307 : sel_960304;
  assign add_960311 = sel_960308 + 8'h01;
  assign sel_960312 = array_index_959947 == array_index_949033 ? add_960311 : sel_960308;
  assign add_960315 = sel_960312 + 8'h01;
  assign sel_960316 = array_index_959947 == array_index_949039 ? add_960315 : sel_960312;
  assign add_960319 = sel_960316 + 8'h01;
  assign sel_960320 = array_index_959947 == array_index_949045 ? add_960319 : sel_960316;
  assign add_960323 = sel_960320 + 8'h01;
  assign sel_960324 = array_index_959947 == array_index_949051 ? add_960323 : sel_960320;
  assign add_960327 = sel_960324 + 8'h01;
  assign sel_960328 = array_index_959947 == array_index_949057 ? add_960327 : sel_960324;
  assign add_960331 = sel_960328 + 8'h01;
  assign sel_960332 = array_index_959947 == array_index_949063 ? add_960331 : sel_960328;
  assign add_960335 = sel_960332 + 8'h01;
  assign sel_960336 = array_index_959947 == array_index_949069 ? add_960335 : sel_960332;
  assign add_960339 = sel_960336 + 8'h01;
  assign sel_960340 = array_index_959947 == array_index_949075 ? add_960339 : sel_960336;
  assign add_960343 = sel_960340 + 8'h01;
  assign sel_960344 = array_index_959947 == array_index_949081 ? add_960343 : sel_960340;
  assign add_960348 = sel_960344 + 8'h01;
  assign array_index_960349 = set1_unflattened[7'h1d];
  assign sel_960350 = array_index_959947 == array_index_949087 ? add_960348 : sel_960344;
  assign add_960353 = sel_960350 + 8'h01;
  assign sel_960354 = array_index_960349 == array_index_948483 ? add_960353 : sel_960350;
  assign add_960357 = sel_960354 + 8'h01;
  assign sel_960358 = array_index_960349 == array_index_948487 ? add_960357 : sel_960354;
  assign add_960361 = sel_960358 + 8'h01;
  assign sel_960362 = array_index_960349 == array_index_948495 ? add_960361 : sel_960358;
  assign add_960365 = sel_960362 + 8'h01;
  assign sel_960366 = array_index_960349 == array_index_948503 ? add_960365 : sel_960362;
  assign add_960369 = sel_960366 + 8'h01;
  assign sel_960370 = array_index_960349 == array_index_948511 ? add_960369 : sel_960366;
  assign add_960373 = sel_960370 + 8'h01;
  assign sel_960374 = array_index_960349 == array_index_948519 ? add_960373 : sel_960370;
  assign add_960377 = sel_960374 + 8'h01;
  assign sel_960378 = array_index_960349 == array_index_948527 ? add_960377 : sel_960374;
  assign add_960381 = sel_960378 + 8'h01;
  assign sel_960382 = array_index_960349 == array_index_948535 ? add_960381 : sel_960378;
  assign add_960385 = sel_960382 + 8'h01;
  assign sel_960386 = array_index_960349 == array_index_948541 ? add_960385 : sel_960382;
  assign add_960389 = sel_960386 + 8'h01;
  assign sel_960390 = array_index_960349 == array_index_948547 ? add_960389 : sel_960386;
  assign add_960393 = sel_960390 + 8'h01;
  assign sel_960394 = array_index_960349 == array_index_948553 ? add_960393 : sel_960390;
  assign add_960397 = sel_960394 + 8'h01;
  assign sel_960398 = array_index_960349 == array_index_948559 ? add_960397 : sel_960394;
  assign add_960401 = sel_960398 + 8'h01;
  assign sel_960402 = array_index_960349 == array_index_948565 ? add_960401 : sel_960398;
  assign add_960405 = sel_960402 + 8'h01;
  assign sel_960406 = array_index_960349 == array_index_948571 ? add_960405 : sel_960402;
  assign add_960409 = sel_960406 + 8'h01;
  assign sel_960410 = array_index_960349 == array_index_948577 ? add_960409 : sel_960406;
  assign add_960413 = sel_960410 + 8'h01;
  assign sel_960414 = array_index_960349 == array_index_948583 ? add_960413 : sel_960410;
  assign add_960417 = sel_960414 + 8'h01;
  assign sel_960418 = array_index_960349 == array_index_948589 ? add_960417 : sel_960414;
  assign add_960421 = sel_960418 + 8'h01;
  assign sel_960422 = array_index_960349 == array_index_948595 ? add_960421 : sel_960418;
  assign add_960425 = sel_960422 + 8'h01;
  assign sel_960426 = array_index_960349 == array_index_948601 ? add_960425 : sel_960422;
  assign add_960429 = sel_960426 + 8'h01;
  assign sel_960430 = array_index_960349 == array_index_948607 ? add_960429 : sel_960426;
  assign add_960433 = sel_960430 + 8'h01;
  assign sel_960434 = array_index_960349 == array_index_948613 ? add_960433 : sel_960430;
  assign add_960437 = sel_960434 + 8'h01;
  assign sel_960438 = array_index_960349 == array_index_948619 ? add_960437 : sel_960434;
  assign add_960441 = sel_960438 + 8'h01;
  assign sel_960442 = array_index_960349 == array_index_948625 ? add_960441 : sel_960438;
  assign add_960445 = sel_960442 + 8'h01;
  assign sel_960446 = array_index_960349 == array_index_948631 ? add_960445 : sel_960442;
  assign add_960449 = sel_960446 + 8'h01;
  assign sel_960450 = array_index_960349 == array_index_948637 ? add_960449 : sel_960446;
  assign add_960453 = sel_960450 + 8'h01;
  assign sel_960454 = array_index_960349 == array_index_948643 ? add_960453 : sel_960450;
  assign add_960457 = sel_960454 + 8'h01;
  assign sel_960458 = array_index_960349 == array_index_948649 ? add_960457 : sel_960454;
  assign add_960461 = sel_960458 + 8'h01;
  assign sel_960462 = array_index_960349 == array_index_948655 ? add_960461 : sel_960458;
  assign add_960465 = sel_960462 + 8'h01;
  assign sel_960466 = array_index_960349 == array_index_948661 ? add_960465 : sel_960462;
  assign add_960469 = sel_960466 + 8'h01;
  assign sel_960470 = array_index_960349 == array_index_948667 ? add_960469 : sel_960466;
  assign add_960473 = sel_960470 + 8'h01;
  assign sel_960474 = array_index_960349 == array_index_948673 ? add_960473 : sel_960470;
  assign add_960477 = sel_960474 + 8'h01;
  assign sel_960478 = array_index_960349 == array_index_948679 ? add_960477 : sel_960474;
  assign add_960481 = sel_960478 + 8'h01;
  assign sel_960482 = array_index_960349 == array_index_948685 ? add_960481 : sel_960478;
  assign add_960485 = sel_960482 + 8'h01;
  assign sel_960486 = array_index_960349 == array_index_948691 ? add_960485 : sel_960482;
  assign add_960489 = sel_960486 + 8'h01;
  assign sel_960490 = array_index_960349 == array_index_948697 ? add_960489 : sel_960486;
  assign add_960493 = sel_960490 + 8'h01;
  assign sel_960494 = array_index_960349 == array_index_948703 ? add_960493 : sel_960490;
  assign add_960497 = sel_960494 + 8'h01;
  assign sel_960498 = array_index_960349 == array_index_948709 ? add_960497 : sel_960494;
  assign add_960501 = sel_960498 + 8'h01;
  assign sel_960502 = array_index_960349 == array_index_948715 ? add_960501 : sel_960498;
  assign add_960505 = sel_960502 + 8'h01;
  assign sel_960506 = array_index_960349 == array_index_948721 ? add_960505 : sel_960502;
  assign add_960509 = sel_960506 + 8'h01;
  assign sel_960510 = array_index_960349 == array_index_948727 ? add_960509 : sel_960506;
  assign add_960513 = sel_960510 + 8'h01;
  assign sel_960514 = array_index_960349 == array_index_948733 ? add_960513 : sel_960510;
  assign add_960517 = sel_960514 + 8'h01;
  assign sel_960518 = array_index_960349 == array_index_948739 ? add_960517 : sel_960514;
  assign add_960521 = sel_960518 + 8'h01;
  assign sel_960522 = array_index_960349 == array_index_948745 ? add_960521 : sel_960518;
  assign add_960525 = sel_960522 + 8'h01;
  assign sel_960526 = array_index_960349 == array_index_948751 ? add_960525 : sel_960522;
  assign add_960529 = sel_960526 + 8'h01;
  assign sel_960530 = array_index_960349 == array_index_948757 ? add_960529 : sel_960526;
  assign add_960533 = sel_960530 + 8'h01;
  assign sel_960534 = array_index_960349 == array_index_948763 ? add_960533 : sel_960530;
  assign add_960537 = sel_960534 + 8'h01;
  assign sel_960538 = array_index_960349 == array_index_948769 ? add_960537 : sel_960534;
  assign add_960541 = sel_960538 + 8'h01;
  assign sel_960542 = array_index_960349 == array_index_948775 ? add_960541 : sel_960538;
  assign add_960545 = sel_960542 + 8'h01;
  assign sel_960546 = array_index_960349 == array_index_948781 ? add_960545 : sel_960542;
  assign add_960549 = sel_960546 + 8'h01;
  assign sel_960550 = array_index_960349 == array_index_948787 ? add_960549 : sel_960546;
  assign add_960553 = sel_960550 + 8'h01;
  assign sel_960554 = array_index_960349 == array_index_948793 ? add_960553 : sel_960550;
  assign add_960557 = sel_960554 + 8'h01;
  assign sel_960558 = array_index_960349 == array_index_948799 ? add_960557 : sel_960554;
  assign add_960561 = sel_960558 + 8'h01;
  assign sel_960562 = array_index_960349 == array_index_948805 ? add_960561 : sel_960558;
  assign add_960565 = sel_960562 + 8'h01;
  assign sel_960566 = array_index_960349 == array_index_948811 ? add_960565 : sel_960562;
  assign add_960569 = sel_960566 + 8'h01;
  assign sel_960570 = array_index_960349 == array_index_948817 ? add_960569 : sel_960566;
  assign add_960573 = sel_960570 + 8'h01;
  assign sel_960574 = array_index_960349 == array_index_948823 ? add_960573 : sel_960570;
  assign add_960577 = sel_960574 + 8'h01;
  assign sel_960578 = array_index_960349 == array_index_948829 ? add_960577 : sel_960574;
  assign add_960581 = sel_960578 + 8'h01;
  assign sel_960582 = array_index_960349 == array_index_948835 ? add_960581 : sel_960578;
  assign add_960585 = sel_960582 + 8'h01;
  assign sel_960586 = array_index_960349 == array_index_948841 ? add_960585 : sel_960582;
  assign add_960589 = sel_960586 + 8'h01;
  assign sel_960590 = array_index_960349 == array_index_948847 ? add_960589 : sel_960586;
  assign add_960593 = sel_960590 + 8'h01;
  assign sel_960594 = array_index_960349 == array_index_948853 ? add_960593 : sel_960590;
  assign add_960597 = sel_960594 + 8'h01;
  assign sel_960598 = array_index_960349 == array_index_948859 ? add_960597 : sel_960594;
  assign add_960601 = sel_960598 + 8'h01;
  assign sel_960602 = array_index_960349 == array_index_948865 ? add_960601 : sel_960598;
  assign add_960605 = sel_960602 + 8'h01;
  assign sel_960606 = array_index_960349 == array_index_948871 ? add_960605 : sel_960602;
  assign add_960609 = sel_960606 + 8'h01;
  assign sel_960610 = array_index_960349 == array_index_948877 ? add_960609 : sel_960606;
  assign add_960613 = sel_960610 + 8'h01;
  assign sel_960614 = array_index_960349 == array_index_948883 ? add_960613 : sel_960610;
  assign add_960617 = sel_960614 + 8'h01;
  assign sel_960618 = array_index_960349 == array_index_948889 ? add_960617 : sel_960614;
  assign add_960621 = sel_960618 + 8'h01;
  assign sel_960622 = array_index_960349 == array_index_948895 ? add_960621 : sel_960618;
  assign add_960625 = sel_960622 + 8'h01;
  assign sel_960626 = array_index_960349 == array_index_948901 ? add_960625 : sel_960622;
  assign add_960629 = sel_960626 + 8'h01;
  assign sel_960630 = array_index_960349 == array_index_948907 ? add_960629 : sel_960626;
  assign add_960633 = sel_960630 + 8'h01;
  assign sel_960634 = array_index_960349 == array_index_948913 ? add_960633 : sel_960630;
  assign add_960637 = sel_960634 + 8'h01;
  assign sel_960638 = array_index_960349 == array_index_948919 ? add_960637 : sel_960634;
  assign add_960641 = sel_960638 + 8'h01;
  assign sel_960642 = array_index_960349 == array_index_948925 ? add_960641 : sel_960638;
  assign add_960645 = sel_960642 + 8'h01;
  assign sel_960646 = array_index_960349 == array_index_948931 ? add_960645 : sel_960642;
  assign add_960649 = sel_960646 + 8'h01;
  assign sel_960650 = array_index_960349 == array_index_948937 ? add_960649 : sel_960646;
  assign add_960653 = sel_960650 + 8'h01;
  assign sel_960654 = array_index_960349 == array_index_948943 ? add_960653 : sel_960650;
  assign add_960657 = sel_960654 + 8'h01;
  assign sel_960658 = array_index_960349 == array_index_948949 ? add_960657 : sel_960654;
  assign add_960661 = sel_960658 + 8'h01;
  assign sel_960662 = array_index_960349 == array_index_948955 ? add_960661 : sel_960658;
  assign add_960665 = sel_960662 + 8'h01;
  assign sel_960666 = array_index_960349 == array_index_948961 ? add_960665 : sel_960662;
  assign add_960669 = sel_960666 + 8'h01;
  assign sel_960670 = array_index_960349 == array_index_948967 ? add_960669 : sel_960666;
  assign add_960673 = sel_960670 + 8'h01;
  assign sel_960674 = array_index_960349 == array_index_948973 ? add_960673 : sel_960670;
  assign add_960677 = sel_960674 + 8'h01;
  assign sel_960678 = array_index_960349 == array_index_948979 ? add_960677 : sel_960674;
  assign add_960681 = sel_960678 + 8'h01;
  assign sel_960682 = array_index_960349 == array_index_948985 ? add_960681 : sel_960678;
  assign add_960685 = sel_960682 + 8'h01;
  assign sel_960686 = array_index_960349 == array_index_948991 ? add_960685 : sel_960682;
  assign add_960689 = sel_960686 + 8'h01;
  assign sel_960690 = array_index_960349 == array_index_948997 ? add_960689 : sel_960686;
  assign add_960693 = sel_960690 + 8'h01;
  assign sel_960694 = array_index_960349 == array_index_949003 ? add_960693 : sel_960690;
  assign add_960697 = sel_960694 + 8'h01;
  assign sel_960698 = array_index_960349 == array_index_949009 ? add_960697 : sel_960694;
  assign add_960701 = sel_960698 + 8'h01;
  assign sel_960702 = array_index_960349 == array_index_949015 ? add_960701 : sel_960698;
  assign add_960705 = sel_960702 + 8'h01;
  assign sel_960706 = array_index_960349 == array_index_949021 ? add_960705 : sel_960702;
  assign add_960709 = sel_960706 + 8'h01;
  assign sel_960710 = array_index_960349 == array_index_949027 ? add_960709 : sel_960706;
  assign add_960713 = sel_960710 + 8'h01;
  assign sel_960714 = array_index_960349 == array_index_949033 ? add_960713 : sel_960710;
  assign add_960717 = sel_960714 + 8'h01;
  assign sel_960718 = array_index_960349 == array_index_949039 ? add_960717 : sel_960714;
  assign add_960721 = sel_960718 + 8'h01;
  assign sel_960722 = array_index_960349 == array_index_949045 ? add_960721 : sel_960718;
  assign add_960725 = sel_960722 + 8'h01;
  assign sel_960726 = array_index_960349 == array_index_949051 ? add_960725 : sel_960722;
  assign add_960729 = sel_960726 + 8'h01;
  assign sel_960730 = array_index_960349 == array_index_949057 ? add_960729 : sel_960726;
  assign add_960733 = sel_960730 + 8'h01;
  assign sel_960734 = array_index_960349 == array_index_949063 ? add_960733 : sel_960730;
  assign add_960737 = sel_960734 + 8'h01;
  assign sel_960738 = array_index_960349 == array_index_949069 ? add_960737 : sel_960734;
  assign add_960741 = sel_960738 + 8'h01;
  assign sel_960742 = array_index_960349 == array_index_949075 ? add_960741 : sel_960738;
  assign add_960745 = sel_960742 + 8'h01;
  assign sel_960746 = array_index_960349 == array_index_949081 ? add_960745 : sel_960742;
  assign add_960750 = sel_960746 + 8'h01;
  assign array_index_960751 = set1_unflattened[7'h1e];
  assign sel_960752 = array_index_960349 == array_index_949087 ? add_960750 : sel_960746;
  assign add_960755 = sel_960752 + 8'h01;
  assign sel_960756 = array_index_960751 == array_index_948483 ? add_960755 : sel_960752;
  assign add_960759 = sel_960756 + 8'h01;
  assign sel_960760 = array_index_960751 == array_index_948487 ? add_960759 : sel_960756;
  assign add_960763 = sel_960760 + 8'h01;
  assign sel_960764 = array_index_960751 == array_index_948495 ? add_960763 : sel_960760;
  assign add_960767 = sel_960764 + 8'h01;
  assign sel_960768 = array_index_960751 == array_index_948503 ? add_960767 : sel_960764;
  assign add_960771 = sel_960768 + 8'h01;
  assign sel_960772 = array_index_960751 == array_index_948511 ? add_960771 : sel_960768;
  assign add_960775 = sel_960772 + 8'h01;
  assign sel_960776 = array_index_960751 == array_index_948519 ? add_960775 : sel_960772;
  assign add_960779 = sel_960776 + 8'h01;
  assign sel_960780 = array_index_960751 == array_index_948527 ? add_960779 : sel_960776;
  assign add_960783 = sel_960780 + 8'h01;
  assign sel_960784 = array_index_960751 == array_index_948535 ? add_960783 : sel_960780;
  assign add_960787 = sel_960784 + 8'h01;
  assign sel_960788 = array_index_960751 == array_index_948541 ? add_960787 : sel_960784;
  assign add_960791 = sel_960788 + 8'h01;
  assign sel_960792 = array_index_960751 == array_index_948547 ? add_960791 : sel_960788;
  assign add_960795 = sel_960792 + 8'h01;
  assign sel_960796 = array_index_960751 == array_index_948553 ? add_960795 : sel_960792;
  assign add_960799 = sel_960796 + 8'h01;
  assign sel_960800 = array_index_960751 == array_index_948559 ? add_960799 : sel_960796;
  assign add_960803 = sel_960800 + 8'h01;
  assign sel_960804 = array_index_960751 == array_index_948565 ? add_960803 : sel_960800;
  assign add_960807 = sel_960804 + 8'h01;
  assign sel_960808 = array_index_960751 == array_index_948571 ? add_960807 : sel_960804;
  assign add_960811 = sel_960808 + 8'h01;
  assign sel_960812 = array_index_960751 == array_index_948577 ? add_960811 : sel_960808;
  assign add_960815 = sel_960812 + 8'h01;
  assign sel_960816 = array_index_960751 == array_index_948583 ? add_960815 : sel_960812;
  assign add_960819 = sel_960816 + 8'h01;
  assign sel_960820 = array_index_960751 == array_index_948589 ? add_960819 : sel_960816;
  assign add_960823 = sel_960820 + 8'h01;
  assign sel_960824 = array_index_960751 == array_index_948595 ? add_960823 : sel_960820;
  assign add_960827 = sel_960824 + 8'h01;
  assign sel_960828 = array_index_960751 == array_index_948601 ? add_960827 : sel_960824;
  assign add_960831 = sel_960828 + 8'h01;
  assign sel_960832 = array_index_960751 == array_index_948607 ? add_960831 : sel_960828;
  assign add_960835 = sel_960832 + 8'h01;
  assign sel_960836 = array_index_960751 == array_index_948613 ? add_960835 : sel_960832;
  assign add_960839 = sel_960836 + 8'h01;
  assign sel_960840 = array_index_960751 == array_index_948619 ? add_960839 : sel_960836;
  assign add_960843 = sel_960840 + 8'h01;
  assign sel_960844 = array_index_960751 == array_index_948625 ? add_960843 : sel_960840;
  assign add_960847 = sel_960844 + 8'h01;
  assign sel_960848 = array_index_960751 == array_index_948631 ? add_960847 : sel_960844;
  assign add_960851 = sel_960848 + 8'h01;
  assign sel_960852 = array_index_960751 == array_index_948637 ? add_960851 : sel_960848;
  assign add_960855 = sel_960852 + 8'h01;
  assign sel_960856 = array_index_960751 == array_index_948643 ? add_960855 : sel_960852;
  assign add_960859 = sel_960856 + 8'h01;
  assign sel_960860 = array_index_960751 == array_index_948649 ? add_960859 : sel_960856;
  assign add_960863 = sel_960860 + 8'h01;
  assign sel_960864 = array_index_960751 == array_index_948655 ? add_960863 : sel_960860;
  assign add_960867 = sel_960864 + 8'h01;
  assign sel_960868 = array_index_960751 == array_index_948661 ? add_960867 : sel_960864;
  assign add_960871 = sel_960868 + 8'h01;
  assign sel_960872 = array_index_960751 == array_index_948667 ? add_960871 : sel_960868;
  assign add_960875 = sel_960872 + 8'h01;
  assign sel_960876 = array_index_960751 == array_index_948673 ? add_960875 : sel_960872;
  assign add_960879 = sel_960876 + 8'h01;
  assign sel_960880 = array_index_960751 == array_index_948679 ? add_960879 : sel_960876;
  assign add_960883 = sel_960880 + 8'h01;
  assign sel_960884 = array_index_960751 == array_index_948685 ? add_960883 : sel_960880;
  assign add_960887 = sel_960884 + 8'h01;
  assign sel_960888 = array_index_960751 == array_index_948691 ? add_960887 : sel_960884;
  assign add_960891 = sel_960888 + 8'h01;
  assign sel_960892 = array_index_960751 == array_index_948697 ? add_960891 : sel_960888;
  assign add_960895 = sel_960892 + 8'h01;
  assign sel_960896 = array_index_960751 == array_index_948703 ? add_960895 : sel_960892;
  assign add_960899 = sel_960896 + 8'h01;
  assign sel_960900 = array_index_960751 == array_index_948709 ? add_960899 : sel_960896;
  assign add_960903 = sel_960900 + 8'h01;
  assign sel_960904 = array_index_960751 == array_index_948715 ? add_960903 : sel_960900;
  assign add_960907 = sel_960904 + 8'h01;
  assign sel_960908 = array_index_960751 == array_index_948721 ? add_960907 : sel_960904;
  assign add_960911 = sel_960908 + 8'h01;
  assign sel_960912 = array_index_960751 == array_index_948727 ? add_960911 : sel_960908;
  assign add_960915 = sel_960912 + 8'h01;
  assign sel_960916 = array_index_960751 == array_index_948733 ? add_960915 : sel_960912;
  assign add_960919 = sel_960916 + 8'h01;
  assign sel_960920 = array_index_960751 == array_index_948739 ? add_960919 : sel_960916;
  assign add_960923 = sel_960920 + 8'h01;
  assign sel_960924 = array_index_960751 == array_index_948745 ? add_960923 : sel_960920;
  assign add_960927 = sel_960924 + 8'h01;
  assign sel_960928 = array_index_960751 == array_index_948751 ? add_960927 : sel_960924;
  assign add_960931 = sel_960928 + 8'h01;
  assign sel_960932 = array_index_960751 == array_index_948757 ? add_960931 : sel_960928;
  assign add_960935 = sel_960932 + 8'h01;
  assign sel_960936 = array_index_960751 == array_index_948763 ? add_960935 : sel_960932;
  assign add_960939 = sel_960936 + 8'h01;
  assign sel_960940 = array_index_960751 == array_index_948769 ? add_960939 : sel_960936;
  assign add_960943 = sel_960940 + 8'h01;
  assign sel_960944 = array_index_960751 == array_index_948775 ? add_960943 : sel_960940;
  assign add_960947 = sel_960944 + 8'h01;
  assign sel_960948 = array_index_960751 == array_index_948781 ? add_960947 : sel_960944;
  assign add_960951 = sel_960948 + 8'h01;
  assign sel_960952 = array_index_960751 == array_index_948787 ? add_960951 : sel_960948;
  assign add_960955 = sel_960952 + 8'h01;
  assign sel_960956 = array_index_960751 == array_index_948793 ? add_960955 : sel_960952;
  assign add_960959 = sel_960956 + 8'h01;
  assign sel_960960 = array_index_960751 == array_index_948799 ? add_960959 : sel_960956;
  assign add_960963 = sel_960960 + 8'h01;
  assign sel_960964 = array_index_960751 == array_index_948805 ? add_960963 : sel_960960;
  assign add_960967 = sel_960964 + 8'h01;
  assign sel_960968 = array_index_960751 == array_index_948811 ? add_960967 : sel_960964;
  assign add_960971 = sel_960968 + 8'h01;
  assign sel_960972 = array_index_960751 == array_index_948817 ? add_960971 : sel_960968;
  assign add_960975 = sel_960972 + 8'h01;
  assign sel_960976 = array_index_960751 == array_index_948823 ? add_960975 : sel_960972;
  assign add_960979 = sel_960976 + 8'h01;
  assign sel_960980 = array_index_960751 == array_index_948829 ? add_960979 : sel_960976;
  assign add_960983 = sel_960980 + 8'h01;
  assign sel_960984 = array_index_960751 == array_index_948835 ? add_960983 : sel_960980;
  assign add_960987 = sel_960984 + 8'h01;
  assign sel_960988 = array_index_960751 == array_index_948841 ? add_960987 : sel_960984;
  assign add_960991 = sel_960988 + 8'h01;
  assign sel_960992 = array_index_960751 == array_index_948847 ? add_960991 : sel_960988;
  assign add_960995 = sel_960992 + 8'h01;
  assign sel_960996 = array_index_960751 == array_index_948853 ? add_960995 : sel_960992;
  assign add_960999 = sel_960996 + 8'h01;
  assign sel_961000 = array_index_960751 == array_index_948859 ? add_960999 : sel_960996;
  assign add_961003 = sel_961000 + 8'h01;
  assign sel_961004 = array_index_960751 == array_index_948865 ? add_961003 : sel_961000;
  assign add_961007 = sel_961004 + 8'h01;
  assign sel_961008 = array_index_960751 == array_index_948871 ? add_961007 : sel_961004;
  assign add_961011 = sel_961008 + 8'h01;
  assign sel_961012 = array_index_960751 == array_index_948877 ? add_961011 : sel_961008;
  assign add_961015 = sel_961012 + 8'h01;
  assign sel_961016 = array_index_960751 == array_index_948883 ? add_961015 : sel_961012;
  assign add_961019 = sel_961016 + 8'h01;
  assign sel_961020 = array_index_960751 == array_index_948889 ? add_961019 : sel_961016;
  assign add_961023 = sel_961020 + 8'h01;
  assign sel_961024 = array_index_960751 == array_index_948895 ? add_961023 : sel_961020;
  assign add_961027 = sel_961024 + 8'h01;
  assign sel_961028 = array_index_960751 == array_index_948901 ? add_961027 : sel_961024;
  assign add_961031 = sel_961028 + 8'h01;
  assign sel_961032 = array_index_960751 == array_index_948907 ? add_961031 : sel_961028;
  assign add_961035 = sel_961032 + 8'h01;
  assign sel_961036 = array_index_960751 == array_index_948913 ? add_961035 : sel_961032;
  assign add_961039 = sel_961036 + 8'h01;
  assign sel_961040 = array_index_960751 == array_index_948919 ? add_961039 : sel_961036;
  assign add_961043 = sel_961040 + 8'h01;
  assign sel_961044 = array_index_960751 == array_index_948925 ? add_961043 : sel_961040;
  assign add_961047 = sel_961044 + 8'h01;
  assign sel_961048 = array_index_960751 == array_index_948931 ? add_961047 : sel_961044;
  assign add_961051 = sel_961048 + 8'h01;
  assign sel_961052 = array_index_960751 == array_index_948937 ? add_961051 : sel_961048;
  assign add_961055 = sel_961052 + 8'h01;
  assign sel_961056 = array_index_960751 == array_index_948943 ? add_961055 : sel_961052;
  assign add_961059 = sel_961056 + 8'h01;
  assign sel_961060 = array_index_960751 == array_index_948949 ? add_961059 : sel_961056;
  assign add_961063 = sel_961060 + 8'h01;
  assign sel_961064 = array_index_960751 == array_index_948955 ? add_961063 : sel_961060;
  assign add_961067 = sel_961064 + 8'h01;
  assign sel_961068 = array_index_960751 == array_index_948961 ? add_961067 : sel_961064;
  assign add_961071 = sel_961068 + 8'h01;
  assign sel_961072 = array_index_960751 == array_index_948967 ? add_961071 : sel_961068;
  assign add_961075 = sel_961072 + 8'h01;
  assign sel_961076 = array_index_960751 == array_index_948973 ? add_961075 : sel_961072;
  assign add_961079 = sel_961076 + 8'h01;
  assign sel_961080 = array_index_960751 == array_index_948979 ? add_961079 : sel_961076;
  assign add_961083 = sel_961080 + 8'h01;
  assign sel_961084 = array_index_960751 == array_index_948985 ? add_961083 : sel_961080;
  assign add_961087 = sel_961084 + 8'h01;
  assign sel_961088 = array_index_960751 == array_index_948991 ? add_961087 : sel_961084;
  assign add_961091 = sel_961088 + 8'h01;
  assign sel_961092 = array_index_960751 == array_index_948997 ? add_961091 : sel_961088;
  assign add_961095 = sel_961092 + 8'h01;
  assign sel_961096 = array_index_960751 == array_index_949003 ? add_961095 : sel_961092;
  assign add_961099 = sel_961096 + 8'h01;
  assign sel_961100 = array_index_960751 == array_index_949009 ? add_961099 : sel_961096;
  assign add_961103 = sel_961100 + 8'h01;
  assign sel_961104 = array_index_960751 == array_index_949015 ? add_961103 : sel_961100;
  assign add_961107 = sel_961104 + 8'h01;
  assign sel_961108 = array_index_960751 == array_index_949021 ? add_961107 : sel_961104;
  assign add_961111 = sel_961108 + 8'h01;
  assign sel_961112 = array_index_960751 == array_index_949027 ? add_961111 : sel_961108;
  assign add_961115 = sel_961112 + 8'h01;
  assign sel_961116 = array_index_960751 == array_index_949033 ? add_961115 : sel_961112;
  assign add_961119 = sel_961116 + 8'h01;
  assign sel_961120 = array_index_960751 == array_index_949039 ? add_961119 : sel_961116;
  assign add_961123 = sel_961120 + 8'h01;
  assign sel_961124 = array_index_960751 == array_index_949045 ? add_961123 : sel_961120;
  assign add_961127 = sel_961124 + 8'h01;
  assign sel_961128 = array_index_960751 == array_index_949051 ? add_961127 : sel_961124;
  assign add_961131 = sel_961128 + 8'h01;
  assign sel_961132 = array_index_960751 == array_index_949057 ? add_961131 : sel_961128;
  assign add_961135 = sel_961132 + 8'h01;
  assign sel_961136 = array_index_960751 == array_index_949063 ? add_961135 : sel_961132;
  assign add_961139 = sel_961136 + 8'h01;
  assign sel_961140 = array_index_960751 == array_index_949069 ? add_961139 : sel_961136;
  assign add_961143 = sel_961140 + 8'h01;
  assign sel_961144 = array_index_960751 == array_index_949075 ? add_961143 : sel_961140;
  assign add_961147 = sel_961144 + 8'h01;
  assign sel_961148 = array_index_960751 == array_index_949081 ? add_961147 : sel_961144;
  assign add_961152 = sel_961148 + 8'h01;
  assign array_index_961153 = set1_unflattened[7'h1f];
  assign sel_961154 = array_index_960751 == array_index_949087 ? add_961152 : sel_961148;
  assign add_961157 = sel_961154 + 8'h01;
  assign sel_961158 = array_index_961153 == array_index_948483 ? add_961157 : sel_961154;
  assign add_961161 = sel_961158 + 8'h01;
  assign sel_961162 = array_index_961153 == array_index_948487 ? add_961161 : sel_961158;
  assign add_961165 = sel_961162 + 8'h01;
  assign sel_961166 = array_index_961153 == array_index_948495 ? add_961165 : sel_961162;
  assign add_961169 = sel_961166 + 8'h01;
  assign sel_961170 = array_index_961153 == array_index_948503 ? add_961169 : sel_961166;
  assign add_961173 = sel_961170 + 8'h01;
  assign sel_961174 = array_index_961153 == array_index_948511 ? add_961173 : sel_961170;
  assign add_961177 = sel_961174 + 8'h01;
  assign sel_961178 = array_index_961153 == array_index_948519 ? add_961177 : sel_961174;
  assign add_961181 = sel_961178 + 8'h01;
  assign sel_961182 = array_index_961153 == array_index_948527 ? add_961181 : sel_961178;
  assign add_961185 = sel_961182 + 8'h01;
  assign sel_961186 = array_index_961153 == array_index_948535 ? add_961185 : sel_961182;
  assign add_961189 = sel_961186 + 8'h01;
  assign sel_961190 = array_index_961153 == array_index_948541 ? add_961189 : sel_961186;
  assign add_961193 = sel_961190 + 8'h01;
  assign sel_961194 = array_index_961153 == array_index_948547 ? add_961193 : sel_961190;
  assign add_961197 = sel_961194 + 8'h01;
  assign sel_961198 = array_index_961153 == array_index_948553 ? add_961197 : sel_961194;
  assign add_961201 = sel_961198 + 8'h01;
  assign sel_961202 = array_index_961153 == array_index_948559 ? add_961201 : sel_961198;
  assign add_961205 = sel_961202 + 8'h01;
  assign sel_961206 = array_index_961153 == array_index_948565 ? add_961205 : sel_961202;
  assign add_961209 = sel_961206 + 8'h01;
  assign sel_961210 = array_index_961153 == array_index_948571 ? add_961209 : sel_961206;
  assign add_961213 = sel_961210 + 8'h01;
  assign sel_961214 = array_index_961153 == array_index_948577 ? add_961213 : sel_961210;
  assign add_961217 = sel_961214 + 8'h01;
  assign sel_961218 = array_index_961153 == array_index_948583 ? add_961217 : sel_961214;
  assign add_961221 = sel_961218 + 8'h01;
  assign sel_961222 = array_index_961153 == array_index_948589 ? add_961221 : sel_961218;
  assign add_961225 = sel_961222 + 8'h01;
  assign sel_961226 = array_index_961153 == array_index_948595 ? add_961225 : sel_961222;
  assign add_961229 = sel_961226 + 8'h01;
  assign sel_961230 = array_index_961153 == array_index_948601 ? add_961229 : sel_961226;
  assign add_961233 = sel_961230 + 8'h01;
  assign sel_961234 = array_index_961153 == array_index_948607 ? add_961233 : sel_961230;
  assign add_961237 = sel_961234 + 8'h01;
  assign sel_961238 = array_index_961153 == array_index_948613 ? add_961237 : sel_961234;
  assign add_961241 = sel_961238 + 8'h01;
  assign sel_961242 = array_index_961153 == array_index_948619 ? add_961241 : sel_961238;
  assign add_961245 = sel_961242 + 8'h01;
  assign sel_961246 = array_index_961153 == array_index_948625 ? add_961245 : sel_961242;
  assign add_961249 = sel_961246 + 8'h01;
  assign sel_961250 = array_index_961153 == array_index_948631 ? add_961249 : sel_961246;
  assign add_961253 = sel_961250 + 8'h01;
  assign sel_961254 = array_index_961153 == array_index_948637 ? add_961253 : sel_961250;
  assign add_961257 = sel_961254 + 8'h01;
  assign sel_961258 = array_index_961153 == array_index_948643 ? add_961257 : sel_961254;
  assign add_961261 = sel_961258 + 8'h01;
  assign sel_961262 = array_index_961153 == array_index_948649 ? add_961261 : sel_961258;
  assign add_961265 = sel_961262 + 8'h01;
  assign sel_961266 = array_index_961153 == array_index_948655 ? add_961265 : sel_961262;
  assign add_961269 = sel_961266 + 8'h01;
  assign sel_961270 = array_index_961153 == array_index_948661 ? add_961269 : sel_961266;
  assign add_961273 = sel_961270 + 8'h01;
  assign sel_961274 = array_index_961153 == array_index_948667 ? add_961273 : sel_961270;
  assign add_961277 = sel_961274 + 8'h01;
  assign sel_961278 = array_index_961153 == array_index_948673 ? add_961277 : sel_961274;
  assign add_961281 = sel_961278 + 8'h01;
  assign sel_961282 = array_index_961153 == array_index_948679 ? add_961281 : sel_961278;
  assign add_961285 = sel_961282 + 8'h01;
  assign sel_961286 = array_index_961153 == array_index_948685 ? add_961285 : sel_961282;
  assign add_961289 = sel_961286 + 8'h01;
  assign sel_961290 = array_index_961153 == array_index_948691 ? add_961289 : sel_961286;
  assign add_961293 = sel_961290 + 8'h01;
  assign sel_961294 = array_index_961153 == array_index_948697 ? add_961293 : sel_961290;
  assign add_961297 = sel_961294 + 8'h01;
  assign sel_961298 = array_index_961153 == array_index_948703 ? add_961297 : sel_961294;
  assign add_961301 = sel_961298 + 8'h01;
  assign sel_961302 = array_index_961153 == array_index_948709 ? add_961301 : sel_961298;
  assign add_961305 = sel_961302 + 8'h01;
  assign sel_961306 = array_index_961153 == array_index_948715 ? add_961305 : sel_961302;
  assign add_961309 = sel_961306 + 8'h01;
  assign sel_961310 = array_index_961153 == array_index_948721 ? add_961309 : sel_961306;
  assign add_961313 = sel_961310 + 8'h01;
  assign sel_961314 = array_index_961153 == array_index_948727 ? add_961313 : sel_961310;
  assign add_961317 = sel_961314 + 8'h01;
  assign sel_961318 = array_index_961153 == array_index_948733 ? add_961317 : sel_961314;
  assign add_961321 = sel_961318 + 8'h01;
  assign sel_961322 = array_index_961153 == array_index_948739 ? add_961321 : sel_961318;
  assign add_961325 = sel_961322 + 8'h01;
  assign sel_961326 = array_index_961153 == array_index_948745 ? add_961325 : sel_961322;
  assign add_961329 = sel_961326 + 8'h01;
  assign sel_961330 = array_index_961153 == array_index_948751 ? add_961329 : sel_961326;
  assign add_961333 = sel_961330 + 8'h01;
  assign sel_961334 = array_index_961153 == array_index_948757 ? add_961333 : sel_961330;
  assign add_961337 = sel_961334 + 8'h01;
  assign sel_961338 = array_index_961153 == array_index_948763 ? add_961337 : sel_961334;
  assign add_961341 = sel_961338 + 8'h01;
  assign sel_961342 = array_index_961153 == array_index_948769 ? add_961341 : sel_961338;
  assign add_961345 = sel_961342 + 8'h01;
  assign sel_961346 = array_index_961153 == array_index_948775 ? add_961345 : sel_961342;
  assign add_961349 = sel_961346 + 8'h01;
  assign sel_961350 = array_index_961153 == array_index_948781 ? add_961349 : sel_961346;
  assign add_961353 = sel_961350 + 8'h01;
  assign sel_961354 = array_index_961153 == array_index_948787 ? add_961353 : sel_961350;
  assign add_961357 = sel_961354 + 8'h01;
  assign sel_961358 = array_index_961153 == array_index_948793 ? add_961357 : sel_961354;
  assign add_961361 = sel_961358 + 8'h01;
  assign sel_961362 = array_index_961153 == array_index_948799 ? add_961361 : sel_961358;
  assign add_961365 = sel_961362 + 8'h01;
  assign sel_961366 = array_index_961153 == array_index_948805 ? add_961365 : sel_961362;
  assign add_961369 = sel_961366 + 8'h01;
  assign sel_961370 = array_index_961153 == array_index_948811 ? add_961369 : sel_961366;
  assign add_961373 = sel_961370 + 8'h01;
  assign sel_961374 = array_index_961153 == array_index_948817 ? add_961373 : sel_961370;
  assign add_961377 = sel_961374 + 8'h01;
  assign sel_961378 = array_index_961153 == array_index_948823 ? add_961377 : sel_961374;
  assign add_961381 = sel_961378 + 8'h01;
  assign sel_961382 = array_index_961153 == array_index_948829 ? add_961381 : sel_961378;
  assign add_961385 = sel_961382 + 8'h01;
  assign sel_961386 = array_index_961153 == array_index_948835 ? add_961385 : sel_961382;
  assign add_961389 = sel_961386 + 8'h01;
  assign sel_961390 = array_index_961153 == array_index_948841 ? add_961389 : sel_961386;
  assign add_961393 = sel_961390 + 8'h01;
  assign sel_961394 = array_index_961153 == array_index_948847 ? add_961393 : sel_961390;
  assign add_961397 = sel_961394 + 8'h01;
  assign sel_961398 = array_index_961153 == array_index_948853 ? add_961397 : sel_961394;
  assign add_961401 = sel_961398 + 8'h01;
  assign sel_961402 = array_index_961153 == array_index_948859 ? add_961401 : sel_961398;
  assign add_961405 = sel_961402 + 8'h01;
  assign sel_961406 = array_index_961153 == array_index_948865 ? add_961405 : sel_961402;
  assign add_961409 = sel_961406 + 8'h01;
  assign sel_961410 = array_index_961153 == array_index_948871 ? add_961409 : sel_961406;
  assign add_961413 = sel_961410 + 8'h01;
  assign sel_961414 = array_index_961153 == array_index_948877 ? add_961413 : sel_961410;
  assign add_961417 = sel_961414 + 8'h01;
  assign sel_961418 = array_index_961153 == array_index_948883 ? add_961417 : sel_961414;
  assign add_961421 = sel_961418 + 8'h01;
  assign sel_961422 = array_index_961153 == array_index_948889 ? add_961421 : sel_961418;
  assign add_961425 = sel_961422 + 8'h01;
  assign sel_961426 = array_index_961153 == array_index_948895 ? add_961425 : sel_961422;
  assign add_961429 = sel_961426 + 8'h01;
  assign sel_961430 = array_index_961153 == array_index_948901 ? add_961429 : sel_961426;
  assign add_961433 = sel_961430 + 8'h01;
  assign sel_961434 = array_index_961153 == array_index_948907 ? add_961433 : sel_961430;
  assign add_961437 = sel_961434 + 8'h01;
  assign sel_961438 = array_index_961153 == array_index_948913 ? add_961437 : sel_961434;
  assign add_961441 = sel_961438 + 8'h01;
  assign sel_961442 = array_index_961153 == array_index_948919 ? add_961441 : sel_961438;
  assign add_961445 = sel_961442 + 8'h01;
  assign sel_961446 = array_index_961153 == array_index_948925 ? add_961445 : sel_961442;
  assign add_961449 = sel_961446 + 8'h01;
  assign sel_961450 = array_index_961153 == array_index_948931 ? add_961449 : sel_961446;
  assign add_961453 = sel_961450 + 8'h01;
  assign sel_961454 = array_index_961153 == array_index_948937 ? add_961453 : sel_961450;
  assign add_961457 = sel_961454 + 8'h01;
  assign sel_961458 = array_index_961153 == array_index_948943 ? add_961457 : sel_961454;
  assign add_961461 = sel_961458 + 8'h01;
  assign sel_961462 = array_index_961153 == array_index_948949 ? add_961461 : sel_961458;
  assign add_961465 = sel_961462 + 8'h01;
  assign sel_961466 = array_index_961153 == array_index_948955 ? add_961465 : sel_961462;
  assign add_961469 = sel_961466 + 8'h01;
  assign sel_961470 = array_index_961153 == array_index_948961 ? add_961469 : sel_961466;
  assign add_961473 = sel_961470 + 8'h01;
  assign sel_961474 = array_index_961153 == array_index_948967 ? add_961473 : sel_961470;
  assign add_961477 = sel_961474 + 8'h01;
  assign sel_961478 = array_index_961153 == array_index_948973 ? add_961477 : sel_961474;
  assign add_961481 = sel_961478 + 8'h01;
  assign sel_961482 = array_index_961153 == array_index_948979 ? add_961481 : sel_961478;
  assign add_961485 = sel_961482 + 8'h01;
  assign sel_961486 = array_index_961153 == array_index_948985 ? add_961485 : sel_961482;
  assign add_961489 = sel_961486 + 8'h01;
  assign sel_961490 = array_index_961153 == array_index_948991 ? add_961489 : sel_961486;
  assign add_961493 = sel_961490 + 8'h01;
  assign sel_961494 = array_index_961153 == array_index_948997 ? add_961493 : sel_961490;
  assign add_961497 = sel_961494 + 8'h01;
  assign sel_961498 = array_index_961153 == array_index_949003 ? add_961497 : sel_961494;
  assign add_961501 = sel_961498 + 8'h01;
  assign sel_961502 = array_index_961153 == array_index_949009 ? add_961501 : sel_961498;
  assign add_961505 = sel_961502 + 8'h01;
  assign sel_961506 = array_index_961153 == array_index_949015 ? add_961505 : sel_961502;
  assign add_961509 = sel_961506 + 8'h01;
  assign sel_961510 = array_index_961153 == array_index_949021 ? add_961509 : sel_961506;
  assign add_961513 = sel_961510 + 8'h01;
  assign sel_961514 = array_index_961153 == array_index_949027 ? add_961513 : sel_961510;
  assign add_961517 = sel_961514 + 8'h01;
  assign sel_961518 = array_index_961153 == array_index_949033 ? add_961517 : sel_961514;
  assign add_961521 = sel_961518 + 8'h01;
  assign sel_961522 = array_index_961153 == array_index_949039 ? add_961521 : sel_961518;
  assign add_961525 = sel_961522 + 8'h01;
  assign sel_961526 = array_index_961153 == array_index_949045 ? add_961525 : sel_961522;
  assign add_961529 = sel_961526 + 8'h01;
  assign sel_961530 = array_index_961153 == array_index_949051 ? add_961529 : sel_961526;
  assign add_961533 = sel_961530 + 8'h01;
  assign sel_961534 = array_index_961153 == array_index_949057 ? add_961533 : sel_961530;
  assign add_961537 = sel_961534 + 8'h01;
  assign sel_961538 = array_index_961153 == array_index_949063 ? add_961537 : sel_961534;
  assign add_961541 = sel_961538 + 8'h01;
  assign sel_961542 = array_index_961153 == array_index_949069 ? add_961541 : sel_961538;
  assign add_961545 = sel_961542 + 8'h01;
  assign sel_961546 = array_index_961153 == array_index_949075 ? add_961545 : sel_961542;
  assign add_961549 = sel_961546 + 8'h01;
  assign sel_961550 = array_index_961153 == array_index_949081 ? add_961549 : sel_961546;
  assign add_961554 = sel_961550 + 8'h01;
  assign array_index_961555 = set1_unflattened[7'h20];
  assign sel_961556 = array_index_961153 == array_index_949087 ? add_961554 : sel_961550;
  assign add_961559 = sel_961556 + 8'h01;
  assign sel_961560 = array_index_961555 == array_index_948483 ? add_961559 : sel_961556;
  assign add_961563 = sel_961560 + 8'h01;
  assign sel_961564 = array_index_961555 == array_index_948487 ? add_961563 : sel_961560;
  assign add_961567 = sel_961564 + 8'h01;
  assign sel_961568 = array_index_961555 == array_index_948495 ? add_961567 : sel_961564;
  assign add_961571 = sel_961568 + 8'h01;
  assign sel_961572 = array_index_961555 == array_index_948503 ? add_961571 : sel_961568;
  assign add_961575 = sel_961572 + 8'h01;
  assign sel_961576 = array_index_961555 == array_index_948511 ? add_961575 : sel_961572;
  assign add_961579 = sel_961576 + 8'h01;
  assign sel_961580 = array_index_961555 == array_index_948519 ? add_961579 : sel_961576;
  assign add_961583 = sel_961580 + 8'h01;
  assign sel_961584 = array_index_961555 == array_index_948527 ? add_961583 : sel_961580;
  assign add_961587 = sel_961584 + 8'h01;
  assign sel_961588 = array_index_961555 == array_index_948535 ? add_961587 : sel_961584;
  assign add_961591 = sel_961588 + 8'h01;
  assign sel_961592 = array_index_961555 == array_index_948541 ? add_961591 : sel_961588;
  assign add_961595 = sel_961592 + 8'h01;
  assign sel_961596 = array_index_961555 == array_index_948547 ? add_961595 : sel_961592;
  assign add_961599 = sel_961596 + 8'h01;
  assign sel_961600 = array_index_961555 == array_index_948553 ? add_961599 : sel_961596;
  assign add_961603 = sel_961600 + 8'h01;
  assign sel_961604 = array_index_961555 == array_index_948559 ? add_961603 : sel_961600;
  assign add_961607 = sel_961604 + 8'h01;
  assign sel_961608 = array_index_961555 == array_index_948565 ? add_961607 : sel_961604;
  assign add_961611 = sel_961608 + 8'h01;
  assign sel_961612 = array_index_961555 == array_index_948571 ? add_961611 : sel_961608;
  assign add_961615 = sel_961612 + 8'h01;
  assign sel_961616 = array_index_961555 == array_index_948577 ? add_961615 : sel_961612;
  assign add_961619 = sel_961616 + 8'h01;
  assign sel_961620 = array_index_961555 == array_index_948583 ? add_961619 : sel_961616;
  assign add_961623 = sel_961620 + 8'h01;
  assign sel_961624 = array_index_961555 == array_index_948589 ? add_961623 : sel_961620;
  assign add_961627 = sel_961624 + 8'h01;
  assign sel_961628 = array_index_961555 == array_index_948595 ? add_961627 : sel_961624;
  assign add_961631 = sel_961628 + 8'h01;
  assign sel_961632 = array_index_961555 == array_index_948601 ? add_961631 : sel_961628;
  assign add_961635 = sel_961632 + 8'h01;
  assign sel_961636 = array_index_961555 == array_index_948607 ? add_961635 : sel_961632;
  assign add_961639 = sel_961636 + 8'h01;
  assign sel_961640 = array_index_961555 == array_index_948613 ? add_961639 : sel_961636;
  assign add_961643 = sel_961640 + 8'h01;
  assign sel_961644 = array_index_961555 == array_index_948619 ? add_961643 : sel_961640;
  assign add_961647 = sel_961644 + 8'h01;
  assign sel_961648 = array_index_961555 == array_index_948625 ? add_961647 : sel_961644;
  assign add_961651 = sel_961648 + 8'h01;
  assign sel_961652 = array_index_961555 == array_index_948631 ? add_961651 : sel_961648;
  assign add_961655 = sel_961652 + 8'h01;
  assign sel_961656 = array_index_961555 == array_index_948637 ? add_961655 : sel_961652;
  assign add_961659 = sel_961656 + 8'h01;
  assign sel_961660 = array_index_961555 == array_index_948643 ? add_961659 : sel_961656;
  assign add_961663 = sel_961660 + 8'h01;
  assign sel_961664 = array_index_961555 == array_index_948649 ? add_961663 : sel_961660;
  assign add_961667 = sel_961664 + 8'h01;
  assign sel_961668 = array_index_961555 == array_index_948655 ? add_961667 : sel_961664;
  assign add_961671 = sel_961668 + 8'h01;
  assign sel_961672 = array_index_961555 == array_index_948661 ? add_961671 : sel_961668;
  assign add_961675 = sel_961672 + 8'h01;
  assign sel_961676 = array_index_961555 == array_index_948667 ? add_961675 : sel_961672;
  assign add_961679 = sel_961676 + 8'h01;
  assign sel_961680 = array_index_961555 == array_index_948673 ? add_961679 : sel_961676;
  assign add_961683 = sel_961680 + 8'h01;
  assign sel_961684 = array_index_961555 == array_index_948679 ? add_961683 : sel_961680;
  assign add_961687 = sel_961684 + 8'h01;
  assign sel_961688 = array_index_961555 == array_index_948685 ? add_961687 : sel_961684;
  assign add_961691 = sel_961688 + 8'h01;
  assign sel_961692 = array_index_961555 == array_index_948691 ? add_961691 : sel_961688;
  assign add_961695 = sel_961692 + 8'h01;
  assign sel_961696 = array_index_961555 == array_index_948697 ? add_961695 : sel_961692;
  assign add_961699 = sel_961696 + 8'h01;
  assign sel_961700 = array_index_961555 == array_index_948703 ? add_961699 : sel_961696;
  assign add_961703 = sel_961700 + 8'h01;
  assign sel_961704 = array_index_961555 == array_index_948709 ? add_961703 : sel_961700;
  assign add_961707 = sel_961704 + 8'h01;
  assign sel_961708 = array_index_961555 == array_index_948715 ? add_961707 : sel_961704;
  assign add_961711 = sel_961708 + 8'h01;
  assign sel_961712 = array_index_961555 == array_index_948721 ? add_961711 : sel_961708;
  assign add_961715 = sel_961712 + 8'h01;
  assign sel_961716 = array_index_961555 == array_index_948727 ? add_961715 : sel_961712;
  assign add_961719 = sel_961716 + 8'h01;
  assign sel_961720 = array_index_961555 == array_index_948733 ? add_961719 : sel_961716;
  assign add_961723 = sel_961720 + 8'h01;
  assign sel_961724 = array_index_961555 == array_index_948739 ? add_961723 : sel_961720;
  assign add_961727 = sel_961724 + 8'h01;
  assign sel_961728 = array_index_961555 == array_index_948745 ? add_961727 : sel_961724;
  assign add_961731 = sel_961728 + 8'h01;
  assign sel_961732 = array_index_961555 == array_index_948751 ? add_961731 : sel_961728;
  assign add_961735 = sel_961732 + 8'h01;
  assign sel_961736 = array_index_961555 == array_index_948757 ? add_961735 : sel_961732;
  assign add_961739 = sel_961736 + 8'h01;
  assign sel_961740 = array_index_961555 == array_index_948763 ? add_961739 : sel_961736;
  assign add_961743 = sel_961740 + 8'h01;
  assign sel_961744 = array_index_961555 == array_index_948769 ? add_961743 : sel_961740;
  assign add_961747 = sel_961744 + 8'h01;
  assign sel_961748 = array_index_961555 == array_index_948775 ? add_961747 : sel_961744;
  assign add_961751 = sel_961748 + 8'h01;
  assign sel_961752 = array_index_961555 == array_index_948781 ? add_961751 : sel_961748;
  assign add_961755 = sel_961752 + 8'h01;
  assign sel_961756 = array_index_961555 == array_index_948787 ? add_961755 : sel_961752;
  assign add_961759 = sel_961756 + 8'h01;
  assign sel_961760 = array_index_961555 == array_index_948793 ? add_961759 : sel_961756;
  assign add_961763 = sel_961760 + 8'h01;
  assign sel_961764 = array_index_961555 == array_index_948799 ? add_961763 : sel_961760;
  assign add_961767 = sel_961764 + 8'h01;
  assign sel_961768 = array_index_961555 == array_index_948805 ? add_961767 : sel_961764;
  assign add_961771 = sel_961768 + 8'h01;
  assign sel_961772 = array_index_961555 == array_index_948811 ? add_961771 : sel_961768;
  assign add_961775 = sel_961772 + 8'h01;
  assign sel_961776 = array_index_961555 == array_index_948817 ? add_961775 : sel_961772;
  assign add_961779 = sel_961776 + 8'h01;
  assign sel_961780 = array_index_961555 == array_index_948823 ? add_961779 : sel_961776;
  assign add_961783 = sel_961780 + 8'h01;
  assign sel_961784 = array_index_961555 == array_index_948829 ? add_961783 : sel_961780;
  assign add_961787 = sel_961784 + 8'h01;
  assign sel_961788 = array_index_961555 == array_index_948835 ? add_961787 : sel_961784;
  assign add_961791 = sel_961788 + 8'h01;
  assign sel_961792 = array_index_961555 == array_index_948841 ? add_961791 : sel_961788;
  assign add_961795 = sel_961792 + 8'h01;
  assign sel_961796 = array_index_961555 == array_index_948847 ? add_961795 : sel_961792;
  assign add_961799 = sel_961796 + 8'h01;
  assign sel_961800 = array_index_961555 == array_index_948853 ? add_961799 : sel_961796;
  assign add_961803 = sel_961800 + 8'h01;
  assign sel_961804 = array_index_961555 == array_index_948859 ? add_961803 : sel_961800;
  assign add_961807 = sel_961804 + 8'h01;
  assign sel_961808 = array_index_961555 == array_index_948865 ? add_961807 : sel_961804;
  assign add_961811 = sel_961808 + 8'h01;
  assign sel_961812 = array_index_961555 == array_index_948871 ? add_961811 : sel_961808;
  assign add_961815 = sel_961812 + 8'h01;
  assign sel_961816 = array_index_961555 == array_index_948877 ? add_961815 : sel_961812;
  assign add_961819 = sel_961816 + 8'h01;
  assign sel_961820 = array_index_961555 == array_index_948883 ? add_961819 : sel_961816;
  assign add_961823 = sel_961820 + 8'h01;
  assign sel_961824 = array_index_961555 == array_index_948889 ? add_961823 : sel_961820;
  assign add_961827 = sel_961824 + 8'h01;
  assign sel_961828 = array_index_961555 == array_index_948895 ? add_961827 : sel_961824;
  assign add_961831 = sel_961828 + 8'h01;
  assign sel_961832 = array_index_961555 == array_index_948901 ? add_961831 : sel_961828;
  assign add_961835 = sel_961832 + 8'h01;
  assign sel_961836 = array_index_961555 == array_index_948907 ? add_961835 : sel_961832;
  assign add_961839 = sel_961836 + 8'h01;
  assign sel_961840 = array_index_961555 == array_index_948913 ? add_961839 : sel_961836;
  assign add_961843 = sel_961840 + 8'h01;
  assign sel_961844 = array_index_961555 == array_index_948919 ? add_961843 : sel_961840;
  assign add_961847 = sel_961844 + 8'h01;
  assign sel_961848 = array_index_961555 == array_index_948925 ? add_961847 : sel_961844;
  assign add_961851 = sel_961848 + 8'h01;
  assign sel_961852 = array_index_961555 == array_index_948931 ? add_961851 : sel_961848;
  assign add_961855 = sel_961852 + 8'h01;
  assign sel_961856 = array_index_961555 == array_index_948937 ? add_961855 : sel_961852;
  assign add_961859 = sel_961856 + 8'h01;
  assign sel_961860 = array_index_961555 == array_index_948943 ? add_961859 : sel_961856;
  assign add_961863 = sel_961860 + 8'h01;
  assign sel_961864 = array_index_961555 == array_index_948949 ? add_961863 : sel_961860;
  assign add_961867 = sel_961864 + 8'h01;
  assign sel_961868 = array_index_961555 == array_index_948955 ? add_961867 : sel_961864;
  assign add_961871 = sel_961868 + 8'h01;
  assign sel_961872 = array_index_961555 == array_index_948961 ? add_961871 : sel_961868;
  assign add_961875 = sel_961872 + 8'h01;
  assign sel_961876 = array_index_961555 == array_index_948967 ? add_961875 : sel_961872;
  assign add_961879 = sel_961876 + 8'h01;
  assign sel_961880 = array_index_961555 == array_index_948973 ? add_961879 : sel_961876;
  assign add_961883 = sel_961880 + 8'h01;
  assign sel_961884 = array_index_961555 == array_index_948979 ? add_961883 : sel_961880;
  assign add_961887 = sel_961884 + 8'h01;
  assign sel_961888 = array_index_961555 == array_index_948985 ? add_961887 : sel_961884;
  assign add_961891 = sel_961888 + 8'h01;
  assign sel_961892 = array_index_961555 == array_index_948991 ? add_961891 : sel_961888;
  assign add_961895 = sel_961892 + 8'h01;
  assign sel_961896 = array_index_961555 == array_index_948997 ? add_961895 : sel_961892;
  assign add_961899 = sel_961896 + 8'h01;
  assign sel_961900 = array_index_961555 == array_index_949003 ? add_961899 : sel_961896;
  assign add_961903 = sel_961900 + 8'h01;
  assign sel_961904 = array_index_961555 == array_index_949009 ? add_961903 : sel_961900;
  assign add_961907 = sel_961904 + 8'h01;
  assign sel_961908 = array_index_961555 == array_index_949015 ? add_961907 : sel_961904;
  assign add_961911 = sel_961908 + 8'h01;
  assign sel_961912 = array_index_961555 == array_index_949021 ? add_961911 : sel_961908;
  assign add_961915 = sel_961912 + 8'h01;
  assign sel_961916 = array_index_961555 == array_index_949027 ? add_961915 : sel_961912;
  assign add_961919 = sel_961916 + 8'h01;
  assign sel_961920 = array_index_961555 == array_index_949033 ? add_961919 : sel_961916;
  assign add_961923 = sel_961920 + 8'h01;
  assign sel_961924 = array_index_961555 == array_index_949039 ? add_961923 : sel_961920;
  assign add_961927 = sel_961924 + 8'h01;
  assign sel_961928 = array_index_961555 == array_index_949045 ? add_961927 : sel_961924;
  assign add_961931 = sel_961928 + 8'h01;
  assign sel_961932 = array_index_961555 == array_index_949051 ? add_961931 : sel_961928;
  assign add_961935 = sel_961932 + 8'h01;
  assign sel_961936 = array_index_961555 == array_index_949057 ? add_961935 : sel_961932;
  assign add_961939 = sel_961936 + 8'h01;
  assign sel_961940 = array_index_961555 == array_index_949063 ? add_961939 : sel_961936;
  assign add_961943 = sel_961940 + 8'h01;
  assign sel_961944 = array_index_961555 == array_index_949069 ? add_961943 : sel_961940;
  assign add_961947 = sel_961944 + 8'h01;
  assign sel_961948 = array_index_961555 == array_index_949075 ? add_961947 : sel_961944;
  assign add_961951 = sel_961948 + 8'h01;
  assign sel_961952 = array_index_961555 == array_index_949081 ? add_961951 : sel_961948;
  assign add_961956 = sel_961952 + 8'h01;
  assign array_index_961957 = set1_unflattened[7'h21];
  assign sel_961958 = array_index_961555 == array_index_949087 ? add_961956 : sel_961952;
  assign add_961961 = sel_961958 + 8'h01;
  assign sel_961962 = array_index_961957 == array_index_948483 ? add_961961 : sel_961958;
  assign add_961965 = sel_961962 + 8'h01;
  assign sel_961966 = array_index_961957 == array_index_948487 ? add_961965 : sel_961962;
  assign add_961969 = sel_961966 + 8'h01;
  assign sel_961970 = array_index_961957 == array_index_948495 ? add_961969 : sel_961966;
  assign add_961973 = sel_961970 + 8'h01;
  assign sel_961974 = array_index_961957 == array_index_948503 ? add_961973 : sel_961970;
  assign add_961977 = sel_961974 + 8'h01;
  assign sel_961978 = array_index_961957 == array_index_948511 ? add_961977 : sel_961974;
  assign add_961981 = sel_961978 + 8'h01;
  assign sel_961982 = array_index_961957 == array_index_948519 ? add_961981 : sel_961978;
  assign add_961985 = sel_961982 + 8'h01;
  assign sel_961986 = array_index_961957 == array_index_948527 ? add_961985 : sel_961982;
  assign add_961989 = sel_961986 + 8'h01;
  assign sel_961990 = array_index_961957 == array_index_948535 ? add_961989 : sel_961986;
  assign add_961993 = sel_961990 + 8'h01;
  assign sel_961994 = array_index_961957 == array_index_948541 ? add_961993 : sel_961990;
  assign add_961997 = sel_961994 + 8'h01;
  assign sel_961998 = array_index_961957 == array_index_948547 ? add_961997 : sel_961994;
  assign add_962001 = sel_961998 + 8'h01;
  assign sel_962002 = array_index_961957 == array_index_948553 ? add_962001 : sel_961998;
  assign add_962005 = sel_962002 + 8'h01;
  assign sel_962006 = array_index_961957 == array_index_948559 ? add_962005 : sel_962002;
  assign add_962009 = sel_962006 + 8'h01;
  assign sel_962010 = array_index_961957 == array_index_948565 ? add_962009 : sel_962006;
  assign add_962013 = sel_962010 + 8'h01;
  assign sel_962014 = array_index_961957 == array_index_948571 ? add_962013 : sel_962010;
  assign add_962017 = sel_962014 + 8'h01;
  assign sel_962018 = array_index_961957 == array_index_948577 ? add_962017 : sel_962014;
  assign add_962021 = sel_962018 + 8'h01;
  assign sel_962022 = array_index_961957 == array_index_948583 ? add_962021 : sel_962018;
  assign add_962025 = sel_962022 + 8'h01;
  assign sel_962026 = array_index_961957 == array_index_948589 ? add_962025 : sel_962022;
  assign add_962029 = sel_962026 + 8'h01;
  assign sel_962030 = array_index_961957 == array_index_948595 ? add_962029 : sel_962026;
  assign add_962033 = sel_962030 + 8'h01;
  assign sel_962034 = array_index_961957 == array_index_948601 ? add_962033 : sel_962030;
  assign add_962037 = sel_962034 + 8'h01;
  assign sel_962038 = array_index_961957 == array_index_948607 ? add_962037 : sel_962034;
  assign add_962041 = sel_962038 + 8'h01;
  assign sel_962042 = array_index_961957 == array_index_948613 ? add_962041 : sel_962038;
  assign add_962045 = sel_962042 + 8'h01;
  assign sel_962046 = array_index_961957 == array_index_948619 ? add_962045 : sel_962042;
  assign add_962049 = sel_962046 + 8'h01;
  assign sel_962050 = array_index_961957 == array_index_948625 ? add_962049 : sel_962046;
  assign add_962053 = sel_962050 + 8'h01;
  assign sel_962054 = array_index_961957 == array_index_948631 ? add_962053 : sel_962050;
  assign add_962057 = sel_962054 + 8'h01;
  assign sel_962058 = array_index_961957 == array_index_948637 ? add_962057 : sel_962054;
  assign add_962061 = sel_962058 + 8'h01;
  assign sel_962062 = array_index_961957 == array_index_948643 ? add_962061 : sel_962058;
  assign add_962065 = sel_962062 + 8'h01;
  assign sel_962066 = array_index_961957 == array_index_948649 ? add_962065 : sel_962062;
  assign add_962069 = sel_962066 + 8'h01;
  assign sel_962070 = array_index_961957 == array_index_948655 ? add_962069 : sel_962066;
  assign add_962073 = sel_962070 + 8'h01;
  assign sel_962074 = array_index_961957 == array_index_948661 ? add_962073 : sel_962070;
  assign add_962077 = sel_962074 + 8'h01;
  assign sel_962078 = array_index_961957 == array_index_948667 ? add_962077 : sel_962074;
  assign add_962081 = sel_962078 + 8'h01;
  assign sel_962082 = array_index_961957 == array_index_948673 ? add_962081 : sel_962078;
  assign add_962085 = sel_962082 + 8'h01;
  assign sel_962086 = array_index_961957 == array_index_948679 ? add_962085 : sel_962082;
  assign add_962089 = sel_962086 + 8'h01;
  assign sel_962090 = array_index_961957 == array_index_948685 ? add_962089 : sel_962086;
  assign add_962093 = sel_962090 + 8'h01;
  assign sel_962094 = array_index_961957 == array_index_948691 ? add_962093 : sel_962090;
  assign add_962097 = sel_962094 + 8'h01;
  assign sel_962098 = array_index_961957 == array_index_948697 ? add_962097 : sel_962094;
  assign add_962101 = sel_962098 + 8'h01;
  assign sel_962102 = array_index_961957 == array_index_948703 ? add_962101 : sel_962098;
  assign add_962105 = sel_962102 + 8'h01;
  assign sel_962106 = array_index_961957 == array_index_948709 ? add_962105 : sel_962102;
  assign add_962109 = sel_962106 + 8'h01;
  assign sel_962110 = array_index_961957 == array_index_948715 ? add_962109 : sel_962106;
  assign add_962113 = sel_962110 + 8'h01;
  assign sel_962114 = array_index_961957 == array_index_948721 ? add_962113 : sel_962110;
  assign add_962117 = sel_962114 + 8'h01;
  assign sel_962118 = array_index_961957 == array_index_948727 ? add_962117 : sel_962114;
  assign add_962121 = sel_962118 + 8'h01;
  assign sel_962122 = array_index_961957 == array_index_948733 ? add_962121 : sel_962118;
  assign add_962125 = sel_962122 + 8'h01;
  assign sel_962126 = array_index_961957 == array_index_948739 ? add_962125 : sel_962122;
  assign add_962129 = sel_962126 + 8'h01;
  assign sel_962130 = array_index_961957 == array_index_948745 ? add_962129 : sel_962126;
  assign add_962133 = sel_962130 + 8'h01;
  assign sel_962134 = array_index_961957 == array_index_948751 ? add_962133 : sel_962130;
  assign add_962137 = sel_962134 + 8'h01;
  assign sel_962138 = array_index_961957 == array_index_948757 ? add_962137 : sel_962134;
  assign add_962141 = sel_962138 + 8'h01;
  assign sel_962142 = array_index_961957 == array_index_948763 ? add_962141 : sel_962138;
  assign add_962145 = sel_962142 + 8'h01;
  assign sel_962146 = array_index_961957 == array_index_948769 ? add_962145 : sel_962142;
  assign add_962149 = sel_962146 + 8'h01;
  assign sel_962150 = array_index_961957 == array_index_948775 ? add_962149 : sel_962146;
  assign add_962153 = sel_962150 + 8'h01;
  assign sel_962154 = array_index_961957 == array_index_948781 ? add_962153 : sel_962150;
  assign add_962157 = sel_962154 + 8'h01;
  assign sel_962158 = array_index_961957 == array_index_948787 ? add_962157 : sel_962154;
  assign add_962161 = sel_962158 + 8'h01;
  assign sel_962162 = array_index_961957 == array_index_948793 ? add_962161 : sel_962158;
  assign add_962165 = sel_962162 + 8'h01;
  assign sel_962166 = array_index_961957 == array_index_948799 ? add_962165 : sel_962162;
  assign add_962169 = sel_962166 + 8'h01;
  assign sel_962170 = array_index_961957 == array_index_948805 ? add_962169 : sel_962166;
  assign add_962173 = sel_962170 + 8'h01;
  assign sel_962174 = array_index_961957 == array_index_948811 ? add_962173 : sel_962170;
  assign add_962177 = sel_962174 + 8'h01;
  assign sel_962178 = array_index_961957 == array_index_948817 ? add_962177 : sel_962174;
  assign add_962181 = sel_962178 + 8'h01;
  assign sel_962182 = array_index_961957 == array_index_948823 ? add_962181 : sel_962178;
  assign add_962185 = sel_962182 + 8'h01;
  assign sel_962186 = array_index_961957 == array_index_948829 ? add_962185 : sel_962182;
  assign add_962189 = sel_962186 + 8'h01;
  assign sel_962190 = array_index_961957 == array_index_948835 ? add_962189 : sel_962186;
  assign add_962193 = sel_962190 + 8'h01;
  assign sel_962194 = array_index_961957 == array_index_948841 ? add_962193 : sel_962190;
  assign add_962197 = sel_962194 + 8'h01;
  assign sel_962198 = array_index_961957 == array_index_948847 ? add_962197 : sel_962194;
  assign add_962201 = sel_962198 + 8'h01;
  assign sel_962202 = array_index_961957 == array_index_948853 ? add_962201 : sel_962198;
  assign add_962205 = sel_962202 + 8'h01;
  assign sel_962206 = array_index_961957 == array_index_948859 ? add_962205 : sel_962202;
  assign add_962209 = sel_962206 + 8'h01;
  assign sel_962210 = array_index_961957 == array_index_948865 ? add_962209 : sel_962206;
  assign add_962213 = sel_962210 + 8'h01;
  assign sel_962214 = array_index_961957 == array_index_948871 ? add_962213 : sel_962210;
  assign add_962217 = sel_962214 + 8'h01;
  assign sel_962218 = array_index_961957 == array_index_948877 ? add_962217 : sel_962214;
  assign add_962221 = sel_962218 + 8'h01;
  assign sel_962222 = array_index_961957 == array_index_948883 ? add_962221 : sel_962218;
  assign add_962225 = sel_962222 + 8'h01;
  assign sel_962226 = array_index_961957 == array_index_948889 ? add_962225 : sel_962222;
  assign add_962229 = sel_962226 + 8'h01;
  assign sel_962230 = array_index_961957 == array_index_948895 ? add_962229 : sel_962226;
  assign add_962233 = sel_962230 + 8'h01;
  assign sel_962234 = array_index_961957 == array_index_948901 ? add_962233 : sel_962230;
  assign add_962237 = sel_962234 + 8'h01;
  assign sel_962238 = array_index_961957 == array_index_948907 ? add_962237 : sel_962234;
  assign add_962241 = sel_962238 + 8'h01;
  assign sel_962242 = array_index_961957 == array_index_948913 ? add_962241 : sel_962238;
  assign add_962245 = sel_962242 + 8'h01;
  assign sel_962246 = array_index_961957 == array_index_948919 ? add_962245 : sel_962242;
  assign add_962249 = sel_962246 + 8'h01;
  assign sel_962250 = array_index_961957 == array_index_948925 ? add_962249 : sel_962246;
  assign add_962253 = sel_962250 + 8'h01;
  assign sel_962254 = array_index_961957 == array_index_948931 ? add_962253 : sel_962250;
  assign add_962257 = sel_962254 + 8'h01;
  assign sel_962258 = array_index_961957 == array_index_948937 ? add_962257 : sel_962254;
  assign add_962261 = sel_962258 + 8'h01;
  assign sel_962262 = array_index_961957 == array_index_948943 ? add_962261 : sel_962258;
  assign add_962265 = sel_962262 + 8'h01;
  assign sel_962266 = array_index_961957 == array_index_948949 ? add_962265 : sel_962262;
  assign add_962269 = sel_962266 + 8'h01;
  assign sel_962270 = array_index_961957 == array_index_948955 ? add_962269 : sel_962266;
  assign add_962273 = sel_962270 + 8'h01;
  assign sel_962274 = array_index_961957 == array_index_948961 ? add_962273 : sel_962270;
  assign add_962277 = sel_962274 + 8'h01;
  assign sel_962278 = array_index_961957 == array_index_948967 ? add_962277 : sel_962274;
  assign add_962281 = sel_962278 + 8'h01;
  assign sel_962282 = array_index_961957 == array_index_948973 ? add_962281 : sel_962278;
  assign add_962285 = sel_962282 + 8'h01;
  assign sel_962286 = array_index_961957 == array_index_948979 ? add_962285 : sel_962282;
  assign add_962289 = sel_962286 + 8'h01;
  assign sel_962290 = array_index_961957 == array_index_948985 ? add_962289 : sel_962286;
  assign add_962293 = sel_962290 + 8'h01;
  assign sel_962294 = array_index_961957 == array_index_948991 ? add_962293 : sel_962290;
  assign add_962297 = sel_962294 + 8'h01;
  assign sel_962298 = array_index_961957 == array_index_948997 ? add_962297 : sel_962294;
  assign add_962301 = sel_962298 + 8'h01;
  assign sel_962302 = array_index_961957 == array_index_949003 ? add_962301 : sel_962298;
  assign add_962305 = sel_962302 + 8'h01;
  assign sel_962306 = array_index_961957 == array_index_949009 ? add_962305 : sel_962302;
  assign add_962309 = sel_962306 + 8'h01;
  assign sel_962310 = array_index_961957 == array_index_949015 ? add_962309 : sel_962306;
  assign add_962313 = sel_962310 + 8'h01;
  assign sel_962314 = array_index_961957 == array_index_949021 ? add_962313 : sel_962310;
  assign add_962317 = sel_962314 + 8'h01;
  assign sel_962318 = array_index_961957 == array_index_949027 ? add_962317 : sel_962314;
  assign add_962321 = sel_962318 + 8'h01;
  assign sel_962322 = array_index_961957 == array_index_949033 ? add_962321 : sel_962318;
  assign add_962325 = sel_962322 + 8'h01;
  assign sel_962326 = array_index_961957 == array_index_949039 ? add_962325 : sel_962322;
  assign add_962329 = sel_962326 + 8'h01;
  assign sel_962330 = array_index_961957 == array_index_949045 ? add_962329 : sel_962326;
  assign add_962333 = sel_962330 + 8'h01;
  assign sel_962334 = array_index_961957 == array_index_949051 ? add_962333 : sel_962330;
  assign add_962337 = sel_962334 + 8'h01;
  assign sel_962338 = array_index_961957 == array_index_949057 ? add_962337 : sel_962334;
  assign add_962341 = sel_962338 + 8'h01;
  assign sel_962342 = array_index_961957 == array_index_949063 ? add_962341 : sel_962338;
  assign add_962345 = sel_962342 + 8'h01;
  assign sel_962346 = array_index_961957 == array_index_949069 ? add_962345 : sel_962342;
  assign add_962349 = sel_962346 + 8'h01;
  assign sel_962350 = array_index_961957 == array_index_949075 ? add_962349 : sel_962346;
  assign add_962353 = sel_962350 + 8'h01;
  assign sel_962354 = array_index_961957 == array_index_949081 ? add_962353 : sel_962350;
  assign add_962358 = sel_962354 + 8'h01;
  assign array_index_962359 = set1_unflattened[7'h22];
  assign sel_962360 = array_index_961957 == array_index_949087 ? add_962358 : sel_962354;
  assign add_962363 = sel_962360 + 8'h01;
  assign sel_962364 = array_index_962359 == array_index_948483 ? add_962363 : sel_962360;
  assign add_962367 = sel_962364 + 8'h01;
  assign sel_962368 = array_index_962359 == array_index_948487 ? add_962367 : sel_962364;
  assign add_962371 = sel_962368 + 8'h01;
  assign sel_962372 = array_index_962359 == array_index_948495 ? add_962371 : sel_962368;
  assign add_962375 = sel_962372 + 8'h01;
  assign sel_962376 = array_index_962359 == array_index_948503 ? add_962375 : sel_962372;
  assign add_962379 = sel_962376 + 8'h01;
  assign sel_962380 = array_index_962359 == array_index_948511 ? add_962379 : sel_962376;
  assign add_962383 = sel_962380 + 8'h01;
  assign sel_962384 = array_index_962359 == array_index_948519 ? add_962383 : sel_962380;
  assign add_962387 = sel_962384 + 8'h01;
  assign sel_962388 = array_index_962359 == array_index_948527 ? add_962387 : sel_962384;
  assign add_962391 = sel_962388 + 8'h01;
  assign sel_962392 = array_index_962359 == array_index_948535 ? add_962391 : sel_962388;
  assign add_962395 = sel_962392 + 8'h01;
  assign sel_962396 = array_index_962359 == array_index_948541 ? add_962395 : sel_962392;
  assign add_962399 = sel_962396 + 8'h01;
  assign sel_962400 = array_index_962359 == array_index_948547 ? add_962399 : sel_962396;
  assign add_962403 = sel_962400 + 8'h01;
  assign sel_962404 = array_index_962359 == array_index_948553 ? add_962403 : sel_962400;
  assign add_962407 = sel_962404 + 8'h01;
  assign sel_962408 = array_index_962359 == array_index_948559 ? add_962407 : sel_962404;
  assign add_962411 = sel_962408 + 8'h01;
  assign sel_962412 = array_index_962359 == array_index_948565 ? add_962411 : sel_962408;
  assign add_962415 = sel_962412 + 8'h01;
  assign sel_962416 = array_index_962359 == array_index_948571 ? add_962415 : sel_962412;
  assign add_962419 = sel_962416 + 8'h01;
  assign sel_962420 = array_index_962359 == array_index_948577 ? add_962419 : sel_962416;
  assign add_962423 = sel_962420 + 8'h01;
  assign sel_962424 = array_index_962359 == array_index_948583 ? add_962423 : sel_962420;
  assign add_962427 = sel_962424 + 8'h01;
  assign sel_962428 = array_index_962359 == array_index_948589 ? add_962427 : sel_962424;
  assign add_962431 = sel_962428 + 8'h01;
  assign sel_962432 = array_index_962359 == array_index_948595 ? add_962431 : sel_962428;
  assign add_962435 = sel_962432 + 8'h01;
  assign sel_962436 = array_index_962359 == array_index_948601 ? add_962435 : sel_962432;
  assign add_962439 = sel_962436 + 8'h01;
  assign sel_962440 = array_index_962359 == array_index_948607 ? add_962439 : sel_962436;
  assign add_962443 = sel_962440 + 8'h01;
  assign sel_962444 = array_index_962359 == array_index_948613 ? add_962443 : sel_962440;
  assign add_962447 = sel_962444 + 8'h01;
  assign sel_962448 = array_index_962359 == array_index_948619 ? add_962447 : sel_962444;
  assign add_962451 = sel_962448 + 8'h01;
  assign sel_962452 = array_index_962359 == array_index_948625 ? add_962451 : sel_962448;
  assign add_962455 = sel_962452 + 8'h01;
  assign sel_962456 = array_index_962359 == array_index_948631 ? add_962455 : sel_962452;
  assign add_962459 = sel_962456 + 8'h01;
  assign sel_962460 = array_index_962359 == array_index_948637 ? add_962459 : sel_962456;
  assign add_962463 = sel_962460 + 8'h01;
  assign sel_962464 = array_index_962359 == array_index_948643 ? add_962463 : sel_962460;
  assign add_962467 = sel_962464 + 8'h01;
  assign sel_962468 = array_index_962359 == array_index_948649 ? add_962467 : sel_962464;
  assign add_962471 = sel_962468 + 8'h01;
  assign sel_962472 = array_index_962359 == array_index_948655 ? add_962471 : sel_962468;
  assign add_962475 = sel_962472 + 8'h01;
  assign sel_962476 = array_index_962359 == array_index_948661 ? add_962475 : sel_962472;
  assign add_962479 = sel_962476 + 8'h01;
  assign sel_962480 = array_index_962359 == array_index_948667 ? add_962479 : sel_962476;
  assign add_962483 = sel_962480 + 8'h01;
  assign sel_962484 = array_index_962359 == array_index_948673 ? add_962483 : sel_962480;
  assign add_962487 = sel_962484 + 8'h01;
  assign sel_962488 = array_index_962359 == array_index_948679 ? add_962487 : sel_962484;
  assign add_962491 = sel_962488 + 8'h01;
  assign sel_962492 = array_index_962359 == array_index_948685 ? add_962491 : sel_962488;
  assign add_962495 = sel_962492 + 8'h01;
  assign sel_962496 = array_index_962359 == array_index_948691 ? add_962495 : sel_962492;
  assign add_962499 = sel_962496 + 8'h01;
  assign sel_962500 = array_index_962359 == array_index_948697 ? add_962499 : sel_962496;
  assign add_962503 = sel_962500 + 8'h01;
  assign sel_962504 = array_index_962359 == array_index_948703 ? add_962503 : sel_962500;
  assign add_962507 = sel_962504 + 8'h01;
  assign sel_962508 = array_index_962359 == array_index_948709 ? add_962507 : sel_962504;
  assign add_962511 = sel_962508 + 8'h01;
  assign sel_962512 = array_index_962359 == array_index_948715 ? add_962511 : sel_962508;
  assign add_962515 = sel_962512 + 8'h01;
  assign sel_962516 = array_index_962359 == array_index_948721 ? add_962515 : sel_962512;
  assign add_962519 = sel_962516 + 8'h01;
  assign sel_962520 = array_index_962359 == array_index_948727 ? add_962519 : sel_962516;
  assign add_962523 = sel_962520 + 8'h01;
  assign sel_962524 = array_index_962359 == array_index_948733 ? add_962523 : sel_962520;
  assign add_962527 = sel_962524 + 8'h01;
  assign sel_962528 = array_index_962359 == array_index_948739 ? add_962527 : sel_962524;
  assign add_962531 = sel_962528 + 8'h01;
  assign sel_962532 = array_index_962359 == array_index_948745 ? add_962531 : sel_962528;
  assign add_962535 = sel_962532 + 8'h01;
  assign sel_962536 = array_index_962359 == array_index_948751 ? add_962535 : sel_962532;
  assign add_962539 = sel_962536 + 8'h01;
  assign sel_962540 = array_index_962359 == array_index_948757 ? add_962539 : sel_962536;
  assign add_962543 = sel_962540 + 8'h01;
  assign sel_962544 = array_index_962359 == array_index_948763 ? add_962543 : sel_962540;
  assign add_962547 = sel_962544 + 8'h01;
  assign sel_962548 = array_index_962359 == array_index_948769 ? add_962547 : sel_962544;
  assign add_962551 = sel_962548 + 8'h01;
  assign sel_962552 = array_index_962359 == array_index_948775 ? add_962551 : sel_962548;
  assign add_962555 = sel_962552 + 8'h01;
  assign sel_962556 = array_index_962359 == array_index_948781 ? add_962555 : sel_962552;
  assign add_962559 = sel_962556 + 8'h01;
  assign sel_962560 = array_index_962359 == array_index_948787 ? add_962559 : sel_962556;
  assign add_962563 = sel_962560 + 8'h01;
  assign sel_962564 = array_index_962359 == array_index_948793 ? add_962563 : sel_962560;
  assign add_962567 = sel_962564 + 8'h01;
  assign sel_962568 = array_index_962359 == array_index_948799 ? add_962567 : sel_962564;
  assign add_962571 = sel_962568 + 8'h01;
  assign sel_962572 = array_index_962359 == array_index_948805 ? add_962571 : sel_962568;
  assign add_962575 = sel_962572 + 8'h01;
  assign sel_962576 = array_index_962359 == array_index_948811 ? add_962575 : sel_962572;
  assign add_962579 = sel_962576 + 8'h01;
  assign sel_962580 = array_index_962359 == array_index_948817 ? add_962579 : sel_962576;
  assign add_962583 = sel_962580 + 8'h01;
  assign sel_962584 = array_index_962359 == array_index_948823 ? add_962583 : sel_962580;
  assign add_962587 = sel_962584 + 8'h01;
  assign sel_962588 = array_index_962359 == array_index_948829 ? add_962587 : sel_962584;
  assign add_962591 = sel_962588 + 8'h01;
  assign sel_962592 = array_index_962359 == array_index_948835 ? add_962591 : sel_962588;
  assign add_962595 = sel_962592 + 8'h01;
  assign sel_962596 = array_index_962359 == array_index_948841 ? add_962595 : sel_962592;
  assign add_962599 = sel_962596 + 8'h01;
  assign sel_962600 = array_index_962359 == array_index_948847 ? add_962599 : sel_962596;
  assign add_962603 = sel_962600 + 8'h01;
  assign sel_962604 = array_index_962359 == array_index_948853 ? add_962603 : sel_962600;
  assign add_962607 = sel_962604 + 8'h01;
  assign sel_962608 = array_index_962359 == array_index_948859 ? add_962607 : sel_962604;
  assign add_962611 = sel_962608 + 8'h01;
  assign sel_962612 = array_index_962359 == array_index_948865 ? add_962611 : sel_962608;
  assign add_962615 = sel_962612 + 8'h01;
  assign sel_962616 = array_index_962359 == array_index_948871 ? add_962615 : sel_962612;
  assign add_962619 = sel_962616 + 8'h01;
  assign sel_962620 = array_index_962359 == array_index_948877 ? add_962619 : sel_962616;
  assign add_962623 = sel_962620 + 8'h01;
  assign sel_962624 = array_index_962359 == array_index_948883 ? add_962623 : sel_962620;
  assign add_962627 = sel_962624 + 8'h01;
  assign sel_962628 = array_index_962359 == array_index_948889 ? add_962627 : sel_962624;
  assign add_962631 = sel_962628 + 8'h01;
  assign sel_962632 = array_index_962359 == array_index_948895 ? add_962631 : sel_962628;
  assign add_962635 = sel_962632 + 8'h01;
  assign sel_962636 = array_index_962359 == array_index_948901 ? add_962635 : sel_962632;
  assign add_962639 = sel_962636 + 8'h01;
  assign sel_962640 = array_index_962359 == array_index_948907 ? add_962639 : sel_962636;
  assign add_962643 = sel_962640 + 8'h01;
  assign sel_962644 = array_index_962359 == array_index_948913 ? add_962643 : sel_962640;
  assign add_962647 = sel_962644 + 8'h01;
  assign sel_962648 = array_index_962359 == array_index_948919 ? add_962647 : sel_962644;
  assign add_962651 = sel_962648 + 8'h01;
  assign sel_962652 = array_index_962359 == array_index_948925 ? add_962651 : sel_962648;
  assign add_962655 = sel_962652 + 8'h01;
  assign sel_962656 = array_index_962359 == array_index_948931 ? add_962655 : sel_962652;
  assign add_962659 = sel_962656 + 8'h01;
  assign sel_962660 = array_index_962359 == array_index_948937 ? add_962659 : sel_962656;
  assign add_962663 = sel_962660 + 8'h01;
  assign sel_962664 = array_index_962359 == array_index_948943 ? add_962663 : sel_962660;
  assign add_962667 = sel_962664 + 8'h01;
  assign sel_962668 = array_index_962359 == array_index_948949 ? add_962667 : sel_962664;
  assign add_962671 = sel_962668 + 8'h01;
  assign sel_962672 = array_index_962359 == array_index_948955 ? add_962671 : sel_962668;
  assign add_962675 = sel_962672 + 8'h01;
  assign sel_962676 = array_index_962359 == array_index_948961 ? add_962675 : sel_962672;
  assign add_962679 = sel_962676 + 8'h01;
  assign sel_962680 = array_index_962359 == array_index_948967 ? add_962679 : sel_962676;
  assign add_962683 = sel_962680 + 8'h01;
  assign sel_962684 = array_index_962359 == array_index_948973 ? add_962683 : sel_962680;
  assign add_962687 = sel_962684 + 8'h01;
  assign sel_962688 = array_index_962359 == array_index_948979 ? add_962687 : sel_962684;
  assign add_962691 = sel_962688 + 8'h01;
  assign sel_962692 = array_index_962359 == array_index_948985 ? add_962691 : sel_962688;
  assign add_962695 = sel_962692 + 8'h01;
  assign sel_962696 = array_index_962359 == array_index_948991 ? add_962695 : sel_962692;
  assign add_962699 = sel_962696 + 8'h01;
  assign sel_962700 = array_index_962359 == array_index_948997 ? add_962699 : sel_962696;
  assign add_962703 = sel_962700 + 8'h01;
  assign sel_962704 = array_index_962359 == array_index_949003 ? add_962703 : sel_962700;
  assign add_962707 = sel_962704 + 8'h01;
  assign sel_962708 = array_index_962359 == array_index_949009 ? add_962707 : sel_962704;
  assign add_962711 = sel_962708 + 8'h01;
  assign sel_962712 = array_index_962359 == array_index_949015 ? add_962711 : sel_962708;
  assign add_962715 = sel_962712 + 8'h01;
  assign sel_962716 = array_index_962359 == array_index_949021 ? add_962715 : sel_962712;
  assign add_962719 = sel_962716 + 8'h01;
  assign sel_962720 = array_index_962359 == array_index_949027 ? add_962719 : sel_962716;
  assign add_962723 = sel_962720 + 8'h01;
  assign sel_962724 = array_index_962359 == array_index_949033 ? add_962723 : sel_962720;
  assign add_962727 = sel_962724 + 8'h01;
  assign sel_962728 = array_index_962359 == array_index_949039 ? add_962727 : sel_962724;
  assign add_962731 = sel_962728 + 8'h01;
  assign sel_962732 = array_index_962359 == array_index_949045 ? add_962731 : sel_962728;
  assign add_962735 = sel_962732 + 8'h01;
  assign sel_962736 = array_index_962359 == array_index_949051 ? add_962735 : sel_962732;
  assign add_962739 = sel_962736 + 8'h01;
  assign sel_962740 = array_index_962359 == array_index_949057 ? add_962739 : sel_962736;
  assign add_962743 = sel_962740 + 8'h01;
  assign sel_962744 = array_index_962359 == array_index_949063 ? add_962743 : sel_962740;
  assign add_962747 = sel_962744 + 8'h01;
  assign sel_962748 = array_index_962359 == array_index_949069 ? add_962747 : sel_962744;
  assign add_962751 = sel_962748 + 8'h01;
  assign sel_962752 = array_index_962359 == array_index_949075 ? add_962751 : sel_962748;
  assign add_962755 = sel_962752 + 8'h01;
  assign sel_962756 = array_index_962359 == array_index_949081 ? add_962755 : sel_962752;
  assign add_962760 = sel_962756 + 8'h01;
  assign array_index_962761 = set1_unflattened[7'h23];
  assign sel_962762 = array_index_962359 == array_index_949087 ? add_962760 : sel_962756;
  assign add_962765 = sel_962762 + 8'h01;
  assign sel_962766 = array_index_962761 == array_index_948483 ? add_962765 : sel_962762;
  assign add_962769 = sel_962766 + 8'h01;
  assign sel_962770 = array_index_962761 == array_index_948487 ? add_962769 : sel_962766;
  assign add_962773 = sel_962770 + 8'h01;
  assign sel_962774 = array_index_962761 == array_index_948495 ? add_962773 : sel_962770;
  assign add_962777 = sel_962774 + 8'h01;
  assign sel_962778 = array_index_962761 == array_index_948503 ? add_962777 : sel_962774;
  assign add_962781 = sel_962778 + 8'h01;
  assign sel_962782 = array_index_962761 == array_index_948511 ? add_962781 : sel_962778;
  assign add_962785 = sel_962782 + 8'h01;
  assign sel_962786 = array_index_962761 == array_index_948519 ? add_962785 : sel_962782;
  assign add_962789 = sel_962786 + 8'h01;
  assign sel_962790 = array_index_962761 == array_index_948527 ? add_962789 : sel_962786;
  assign add_962793 = sel_962790 + 8'h01;
  assign sel_962794 = array_index_962761 == array_index_948535 ? add_962793 : sel_962790;
  assign add_962797 = sel_962794 + 8'h01;
  assign sel_962798 = array_index_962761 == array_index_948541 ? add_962797 : sel_962794;
  assign add_962801 = sel_962798 + 8'h01;
  assign sel_962802 = array_index_962761 == array_index_948547 ? add_962801 : sel_962798;
  assign add_962805 = sel_962802 + 8'h01;
  assign sel_962806 = array_index_962761 == array_index_948553 ? add_962805 : sel_962802;
  assign add_962809 = sel_962806 + 8'h01;
  assign sel_962810 = array_index_962761 == array_index_948559 ? add_962809 : sel_962806;
  assign add_962813 = sel_962810 + 8'h01;
  assign sel_962814 = array_index_962761 == array_index_948565 ? add_962813 : sel_962810;
  assign add_962817 = sel_962814 + 8'h01;
  assign sel_962818 = array_index_962761 == array_index_948571 ? add_962817 : sel_962814;
  assign add_962821 = sel_962818 + 8'h01;
  assign sel_962822 = array_index_962761 == array_index_948577 ? add_962821 : sel_962818;
  assign add_962825 = sel_962822 + 8'h01;
  assign sel_962826 = array_index_962761 == array_index_948583 ? add_962825 : sel_962822;
  assign add_962829 = sel_962826 + 8'h01;
  assign sel_962830 = array_index_962761 == array_index_948589 ? add_962829 : sel_962826;
  assign add_962833 = sel_962830 + 8'h01;
  assign sel_962834 = array_index_962761 == array_index_948595 ? add_962833 : sel_962830;
  assign add_962837 = sel_962834 + 8'h01;
  assign sel_962838 = array_index_962761 == array_index_948601 ? add_962837 : sel_962834;
  assign add_962841 = sel_962838 + 8'h01;
  assign sel_962842 = array_index_962761 == array_index_948607 ? add_962841 : sel_962838;
  assign add_962845 = sel_962842 + 8'h01;
  assign sel_962846 = array_index_962761 == array_index_948613 ? add_962845 : sel_962842;
  assign add_962849 = sel_962846 + 8'h01;
  assign sel_962850 = array_index_962761 == array_index_948619 ? add_962849 : sel_962846;
  assign add_962853 = sel_962850 + 8'h01;
  assign sel_962854 = array_index_962761 == array_index_948625 ? add_962853 : sel_962850;
  assign add_962857 = sel_962854 + 8'h01;
  assign sel_962858 = array_index_962761 == array_index_948631 ? add_962857 : sel_962854;
  assign add_962861 = sel_962858 + 8'h01;
  assign sel_962862 = array_index_962761 == array_index_948637 ? add_962861 : sel_962858;
  assign add_962865 = sel_962862 + 8'h01;
  assign sel_962866 = array_index_962761 == array_index_948643 ? add_962865 : sel_962862;
  assign add_962869 = sel_962866 + 8'h01;
  assign sel_962870 = array_index_962761 == array_index_948649 ? add_962869 : sel_962866;
  assign add_962873 = sel_962870 + 8'h01;
  assign sel_962874 = array_index_962761 == array_index_948655 ? add_962873 : sel_962870;
  assign add_962877 = sel_962874 + 8'h01;
  assign sel_962878 = array_index_962761 == array_index_948661 ? add_962877 : sel_962874;
  assign add_962881 = sel_962878 + 8'h01;
  assign sel_962882 = array_index_962761 == array_index_948667 ? add_962881 : sel_962878;
  assign add_962885 = sel_962882 + 8'h01;
  assign sel_962886 = array_index_962761 == array_index_948673 ? add_962885 : sel_962882;
  assign add_962889 = sel_962886 + 8'h01;
  assign sel_962890 = array_index_962761 == array_index_948679 ? add_962889 : sel_962886;
  assign add_962893 = sel_962890 + 8'h01;
  assign sel_962894 = array_index_962761 == array_index_948685 ? add_962893 : sel_962890;
  assign add_962897 = sel_962894 + 8'h01;
  assign sel_962898 = array_index_962761 == array_index_948691 ? add_962897 : sel_962894;
  assign add_962901 = sel_962898 + 8'h01;
  assign sel_962902 = array_index_962761 == array_index_948697 ? add_962901 : sel_962898;
  assign add_962905 = sel_962902 + 8'h01;
  assign sel_962906 = array_index_962761 == array_index_948703 ? add_962905 : sel_962902;
  assign add_962909 = sel_962906 + 8'h01;
  assign sel_962910 = array_index_962761 == array_index_948709 ? add_962909 : sel_962906;
  assign add_962913 = sel_962910 + 8'h01;
  assign sel_962914 = array_index_962761 == array_index_948715 ? add_962913 : sel_962910;
  assign add_962917 = sel_962914 + 8'h01;
  assign sel_962918 = array_index_962761 == array_index_948721 ? add_962917 : sel_962914;
  assign add_962921 = sel_962918 + 8'h01;
  assign sel_962922 = array_index_962761 == array_index_948727 ? add_962921 : sel_962918;
  assign add_962925 = sel_962922 + 8'h01;
  assign sel_962926 = array_index_962761 == array_index_948733 ? add_962925 : sel_962922;
  assign add_962929 = sel_962926 + 8'h01;
  assign sel_962930 = array_index_962761 == array_index_948739 ? add_962929 : sel_962926;
  assign add_962933 = sel_962930 + 8'h01;
  assign sel_962934 = array_index_962761 == array_index_948745 ? add_962933 : sel_962930;
  assign add_962937 = sel_962934 + 8'h01;
  assign sel_962938 = array_index_962761 == array_index_948751 ? add_962937 : sel_962934;
  assign add_962941 = sel_962938 + 8'h01;
  assign sel_962942 = array_index_962761 == array_index_948757 ? add_962941 : sel_962938;
  assign add_962945 = sel_962942 + 8'h01;
  assign sel_962946 = array_index_962761 == array_index_948763 ? add_962945 : sel_962942;
  assign add_962949 = sel_962946 + 8'h01;
  assign sel_962950 = array_index_962761 == array_index_948769 ? add_962949 : sel_962946;
  assign add_962953 = sel_962950 + 8'h01;
  assign sel_962954 = array_index_962761 == array_index_948775 ? add_962953 : sel_962950;
  assign add_962957 = sel_962954 + 8'h01;
  assign sel_962958 = array_index_962761 == array_index_948781 ? add_962957 : sel_962954;
  assign add_962961 = sel_962958 + 8'h01;
  assign sel_962962 = array_index_962761 == array_index_948787 ? add_962961 : sel_962958;
  assign add_962965 = sel_962962 + 8'h01;
  assign sel_962966 = array_index_962761 == array_index_948793 ? add_962965 : sel_962962;
  assign add_962969 = sel_962966 + 8'h01;
  assign sel_962970 = array_index_962761 == array_index_948799 ? add_962969 : sel_962966;
  assign add_962973 = sel_962970 + 8'h01;
  assign sel_962974 = array_index_962761 == array_index_948805 ? add_962973 : sel_962970;
  assign add_962977 = sel_962974 + 8'h01;
  assign sel_962978 = array_index_962761 == array_index_948811 ? add_962977 : sel_962974;
  assign add_962981 = sel_962978 + 8'h01;
  assign sel_962982 = array_index_962761 == array_index_948817 ? add_962981 : sel_962978;
  assign add_962985 = sel_962982 + 8'h01;
  assign sel_962986 = array_index_962761 == array_index_948823 ? add_962985 : sel_962982;
  assign add_962989 = sel_962986 + 8'h01;
  assign sel_962990 = array_index_962761 == array_index_948829 ? add_962989 : sel_962986;
  assign add_962993 = sel_962990 + 8'h01;
  assign sel_962994 = array_index_962761 == array_index_948835 ? add_962993 : sel_962990;
  assign add_962997 = sel_962994 + 8'h01;
  assign sel_962998 = array_index_962761 == array_index_948841 ? add_962997 : sel_962994;
  assign add_963001 = sel_962998 + 8'h01;
  assign sel_963002 = array_index_962761 == array_index_948847 ? add_963001 : sel_962998;
  assign add_963005 = sel_963002 + 8'h01;
  assign sel_963006 = array_index_962761 == array_index_948853 ? add_963005 : sel_963002;
  assign add_963009 = sel_963006 + 8'h01;
  assign sel_963010 = array_index_962761 == array_index_948859 ? add_963009 : sel_963006;
  assign add_963013 = sel_963010 + 8'h01;
  assign sel_963014 = array_index_962761 == array_index_948865 ? add_963013 : sel_963010;
  assign add_963017 = sel_963014 + 8'h01;
  assign sel_963018 = array_index_962761 == array_index_948871 ? add_963017 : sel_963014;
  assign add_963021 = sel_963018 + 8'h01;
  assign sel_963022 = array_index_962761 == array_index_948877 ? add_963021 : sel_963018;
  assign add_963025 = sel_963022 + 8'h01;
  assign sel_963026 = array_index_962761 == array_index_948883 ? add_963025 : sel_963022;
  assign add_963029 = sel_963026 + 8'h01;
  assign sel_963030 = array_index_962761 == array_index_948889 ? add_963029 : sel_963026;
  assign add_963033 = sel_963030 + 8'h01;
  assign sel_963034 = array_index_962761 == array_index_948895 ? add_963033 : sel_963030;
  assign add_963037 = sel_963034 + 8'h01;
  assign sel_963038 = array_index_962761 == array_index_948901 ? add_963037 : sel_963034;
  assign add_963041 = sel_963038 + 8'h01;
  assign sel_963042 = array_index_962761 == array_index_948907 ? add_963041 : sel_963038;
  assign add_963045 = sel_963042 + 8'h01;
  assign sel_963046 = array_index_962761 == array_index_948913 ? add_963045 : sel_963042;
  assign add_963049 = sel_963046 + 8'h01;
  assign sel_963050 = array_index_962761 == array_index_948919 ? add_963049 : sel_963046;
  assign add_963053 = sel_963050 + 8'h01;
  assign sel_963054 = array_index_962761 == array_index_948925 ? add_963053 : sel_963050;
  assign add_963057 = sel_963054 + 8'h01;
  assign sel_963058 = array_index_962761 == array_index_948931 ? add_963057 : sel_963054;
  assign add_963061 = sel_963058 + 8'h01;
  assign sel_963062 = array_index_962761 == array_index_948937 ? add_963061 : sel_963058;
  assign add_963065 = sel_963062 + 8'h01;
  assign sel_963066 = array_index_962761 == array_index_948943 ? add_963065 : sel_963062;
  assign add_963069 = sel_963066 + 8'h01;
  assign sel_963070 = array_index_962761 == array_index_948949 ? add_963069 : sel_963066;
  assign add_963073 = sel_963070 + 8'h01;
  assign sel_963074 = array_index_962761 == array_index_948955 ? add_963073 : sel_963070;
  assign add_963077 = sel_963074 + 8'h01;
  assign sel_963078 = array_index_962761 == array_index_948961 ? add_963077 : sel_963074;
  assign add_963081 = sel_963078 + 8'h01;
  assign sel_963082 = array_index_962761 == array_index_948967 ? add_963081 : sel_963078;
  assign add_963085 = sel_963082 + 8'h01;
  assign sel_963086 = array_index_962761 == array_index_948973 ? add_963085 : sel_963082;
  assign add_963089 = sel_963086 + 8'h01;
  assign sel_963090 = array_index_962761 == array_index_948979 ? add_963089 : sel_963086;
  assign add_963093 = sel_963090 + 8'h01;
  assign sel_963094 = array_index_962761 == array_index_948985 ? add_963093 : sel_963090;
  assign add_963097 = sel_963094 + 8'h01;
  assign sel_963098 = array_index_962761 == array_index_948991 ? add_963097 : sel_963094;
  assign add_963101 = sel_963098 + 8'h01;
  assign sel_963102 = array_index_962761 == array_index_948997 ? add_963101 : sel_963098;
  assign add_963105 = sel_963102 + 8'h01;
  assign sel_963106 = array_index_962761 == array_index_949003 ? add_963105 : sel_963102;
  assign add_963109 = sel_963106 + 8'h01;
  assign sel_963110 = array_index_962761 == array_index_949009 ? add_963109 : sel_963106;
  assign add_963113 = sel_963110 + 8'h01;
  assign sel_963114 = array_index_962761 == array_index_949015 ? add_963113 : sel_963110;
  assign add_963117 = sel_963114 + 8'h01;
  assign sel_963118 = array_index_962761 == array_index_949021 ? add_963117 : sel_963114;
  assign add_963121 = sel_963118 + 8'h01;
  assign sel_963122 = array_index_962761 == array_index_949027 ? add_963121 : sel_963118;
  assign add_963125 = sel_963122 + 8'h01;
  assign sel_963126 = array_index_962761 == array_index_949033 ? add_963125 : sel_963122;
  assign add_963129 = sel_963126 + 8'h01;
  assign sel_963130 = array_index_962761 == array_index_949039 ? add_963129 : sel_963126;
  assign add_963133 = sel_963130 + 8'h01;
  assign sel_963134 = array_index_962761 == array_index_949045 ? add_963133 : sel_963130;
  assign add_963137 = sel_963134 + 8'h01;
  assign sel_963138 = array_index_962761 == array_index_949051 ? add_963137 : sel_963134;
  assign add_963141 = sel_963138 + 8'h01;
  assign sel_963142 = array_index_962761 == array_index_949057 ? add_963141 : sel_963138;
  assign add_963145 = sel_963142 + 8'h01;
  assign sel_963146 = array_index_962761 == array_index_949063 ? add_963145 : sel_963142;
  assign add_963149 = sel_963146 + 8'h01;
  assign sel_963150 = array_index_962761 == array_index_949069 ? add_963149 : sel_963146;
  assign add_963153 = sel_963150 + 8'h01;
  assign sel_963154 = array_index_962761 == array_index_949075 ? add_963153 : sel_963150;
  assign add_963157 = sel_963154 + 8'h01;
  assign sel_963158 = array_index_962761 == array_index_949081 ? add_963157 : sel_963154;
  assign add_963162 = sel_963158 + 8'h01;
  assign array_index_963163 = set1_unflattened[7'h24];
  assign sel_963164 = array_index_962761 == array_index_949087 ? add_963162 : sel_963158;
  assign add_963167 = sel_963164 + 8'h01;
  assign sel_963168 = array_index_963163 == array_index_948483 ? add_963167 : sel_963164;
  assign add_963171 = sel_963168 + 8'h01;
  assign sel_963172 = array_index_963163 == array_index_948487 ? add_963171 : sel_963168;
  assign add_963175 = sel_963172 + 8'h01;
  assign sel_963176 = array_index_963163 == array_index_948495 ? add_963175 : sel_963172;
  assign add_963179 = sel_963176 + 8'h01;
  assign sel_963180 = array_index_963163 == array_index_948503 ? add_963179 : sel_963176;
  assign add_963183 = sel_963180 + 8'h01;
  assign sel_963184 = array_index_963163 == array_index_948511 ? add_963183 : sel_963180;
  assign add_963187 = sel_963184 + 8'h01;
  assign sel_963188 = array_index_963163 == array_index_948519 ? add_963187 : sel_963184;
  assign add_963191 = sel_963188 + 8'h01;
  assign sel_963192 = array_index_963163 == array_index_948527 ? add_963191 : sel_963188;
  assign add_963195 = sel_963192 + 8'h01;
  assign sel_963196 = array_index_963163 == array_index_948535 ? add_963195 : sel_963192;
  assign add_963199 = sel_963196 + 8'h01;
  assign sel_963200 = array_index_963163 == array_index_948541 ? add_963199 : sel_963196;
  assign add_963203 = sel_963200 + 8'h01;
  assign sel_963204 = array_index_963163 == array_index_948547 ? add_963203 : sel_963200;
  assign add_963207 = sel_963204 + 8'h01;
  assign sel_963208 = array_index_963163 == array_index_948553 ? add_963207 : sel_963204;
  assign add_963211 = sel_963208 + 8'h01;
  assign sel_963212 = array_index_963163 == array_index_948559 ? add_963211 : sel_963208;
  assign add_963215 = sel_963212 + 8'h01;
  assign sel_963216 = array_index_963163 == array_index_948565 ? add_963215 : sel_963212;
  assign add_963219 = sel_963216 + 8'h01;
  assign sel_963220 = array_index_963163 == array_index_948571 ? add_963219 : sel_963216;
  assign add_963223 = sel_963220 + 8'h01;
  assign sel_963224 = array_index_963163 == array_index_948577 ? add_963223 : sel_963220;
  assign add_963227 = sel_963224 + 8'h01;
  assign sel_963228 = array_index_963163 == array_index_948583 ? add_963227 : sel_963224;
  assign add_963231 = sel_963228 + 8'h01;
  assign sel_963232 = array_index_963163 == array_index_948589 ? add_963231 : sel_963228;
  assign add_963235 = sel_963232 + 8'h01;
  assign sel_963236 = array_index_963163 == array_index_948595 ? add_963235 : sel_963232;
  assign add_963239 = sel_963236 + 8'h01;
  assign sel_963240 = array_index_963163 == array_index_948601 ? add_963239 : sel_963236;
  assign add_963243 = sel_963240 + 8'h01;
  assign sel_963244 = array_index_963163 == array_index_948607 ? add_963243 : sel_963240;
  assign add_963247 = sel_963244 + 8'h01;
  assign sel_963248 = array_index_963163 == array_index_948613 ? add_963247 : sel_963244;
  assign add_963251 = sel_963248 + 8'h01;
  assign sel_963252 = array_index_963163 == array_index_948619 ? add_963251 : sel_963248;
  assign add_963255 = sel_963252 + 8'h01;
  assign sel_963256 = array_index_963163 == array_index_948625 ? add_963255 : sel_963252;
  assign add_963259 = sel_963256 + 8'h01;
  assign sel_963260 = array_index_963163 == array_index_948631 ? add_963259 : sel_963256;
  assign add_963263 = sel_963260 + 8'h01;
  assign sel_963264 = array_index_963163 == array_index_948637 ? add_963263 : sel_963260;
  assign add_963267 = sel_963264 + 8'h01;
  assign sel_963268 = array_index_963163 == array_index_948643 ? add_963267 : sel_963264;
  assign add_963271 = sel_963268 + 8'h01;
  assign sel_963272 = array_index_963163 == array_index_948649 ? add_963271 : sel_963268;
  assign add_963275 = sel_963272 + 8'h01;
  assign sel_963276 = array_index_963163 == array_index_948655 ? add_963275 : sel_963272;
  assign add_963279 = sel_963276 + 8'h01;
  assign sel_963280 = array_index_963163 == array_index_948661 ? add_963279 : sel_963276;
  assign add_963283 = sel_963280 + 8'h01;
  assign sel_963284 = array_index_963163 == array_index_948667 ? add_963283 : sel_963280;
  assign add_963287 = sel_963284 + 8'h01;
  assign sel_963288 = array_index_963163 == array_index_948673 ? add_963287 : sel_963284;
  assign add_963291 = sel_963288 + 8'h01;
  assign sel_963292 = array_index_963163 == array_index_948679 ? add_963291 : sel_963288;
  assign add_963295 = sel_963292 + 8'h01;
  assign sel_963296 = array_index_963163 == array_index_948685 ? add_963295 : sel_963292;
  assign add_963299 = sel_963296 + 8'h01;
  assign sel_963300 = array_index_963163 == array_index_948691 ? add_963299 : sel_963296;
  assign add_963303 = sel_963300 + 8'h01;
  assign sel_963304 = array_index_963163 == array_index_948697 ? add_963303 : sel_963300;
  assign add_963307 = sel_963304 + 8'h01;
  assign sel_963308 = array_index_963163 == array_index_948703 ? add_963307 : sel_963304;
  assign add_963311 = sel_963308 + 8'h01;
  assign sel_963312 = array_index_963163 == array_index_948709 ? add_963311 : sel_963308;
  assign add_963315 = sel_963312 + 8'h01;
  assign sel_963316 = array_index_963163 == array_index_948715 ? add_963315 : sel_963312;
  assign add_963319 = sel_963316 + 8'h01;
  assign sel_963320 = array_index_963163 == array_index_948721 ? add_963319 : sel_963316;
  assign add_963323 = sel_963320 + 8'h01;
  assign sel_963324 = array_index_963163 == array_index_948727 ? add_963323 : sel_963320;
  assign add_963327 = sel_963324 + 8'h01;
  assign sel_963328 = array_index_963163 == array_index_948733 ? add_963327 : sel_963324;
  assign add_963331 = sel_963328 + 8'h01;
  assign sel_963332 = array_index_963163 == array_index_948739 ? add_963331 : sel_963328;
  assign add_963335 = sel_963332 + 8'h01;
  assign sel_963336 = array_index_963163 == array_index_948745 ? add_963335 : sel_963332;
  assign add_963339 = sel_963336 + 8'h01;
  assign sel_963340 = array_index_963163 == array_index_948751 ? add_963339 : sel_963336;
  assign add_963343 = sel_963340 + 8'h01;
  assign sel_963344 = array_index_963163 == array_index_948757 ? add_963343 : sel_963340;
  assign add_963347 = sel_963344 + 8'h01;
  assign sel_963348 = array_index_963163 == array_index_948763 ? add_963347 : sel_963344;
  assign add_963351 = sel_963348 + 8'h01;
  assign sel_963352 = array_index_963163 == array_index_948769 ? add_963351 : sel_963348;
  assign add_963355 = sel_963352 + 8'h01;
  assign sel_963356 = array_index_963163 == array_index_948775 ? add_963355 : sel_963352;
  assign add_963359 = sel_963356 + 8'h01;
  assign sel_963360 = array_index_963163 == array_index_948781 ? add_963359 : sel_963356;
  assign add_963363 = sel_963360 + 8'h01;
  assign sel_963364 = array_index_963163 == array_index_948787 ? add_963363 : sel_963360;
  assign add_963367 = sel_963364 + 8'h01;
  assign sel_963368 = array_index_963163 == array_index_948793 ? add_963367 : sel_963364;
  assign add_963371 = sel_963368 + 8'h01;
  assign sel_963372 = array_index_963163 == array_index_948799 ? add_963371 : sel_963368;
  assign add_963375 = sel_963372 + 8'h01;
  assign sel_963376 = array_index_963163 == array_index_948805 ? add_963375 : sel_963372;
  assign add_963379 = sel_963376 + 8'h01;
  assign sel_963380 = array_index_963163 == array_index_948811 ? add_963379 : sel_963376;
  assign add_963383 = sel_963380 + 8'h01;
  assign sel_963384 = array_index_963163 == array_index_948817 ? add_963383 : sel_963380;
  assign add_963387 = sel_963384 + 8'h01;
  assign sel_963388 = array_index_963163 == array_index_948823 ? add_963387 : sel_963384;
  assign add_963391 = sel_963388 + 8'h01;
  assign sel_963392 = array_index_963163 == array_index_948829 ? add_963391 : sel_963388;
  assign add_963395 = sel_963392 + 8'h01;
  assign sel_963396 = array_index_963163 == array_index_948835 ? add_963395 : sel_963392;
  assign add_963399 = sel_963396 + 8'h01;
  assign sel_963400 = array_index_963163 == array_index_948841 ? add_963399 : sel_963396;
  assign add_963403 = sel_963400 + 8'h01;
  assign sel_963404 = array_index_963163 == array_index_948847 ? add_963403 : sel_963400;
  assign add_963407 = sel_963404 + 8'h01;
  assign sel_963408 = array_index_963163 == array_index_948853 ? add_963407 : sel_963404;
  assign add_963411 = sel_963408 + 8'h01;
  assign sel_963412 = array_index_963163 == array_index_948859 ? add_963411 : sel_963408;
  assign add_963415 = sel_963412 + 8'h01;
  assign sel_963416 = array_index_963163 == array_index_948865 ? add_963415 : sel_963412;
  assign add_963419 = sel_963416 + 8'h01;
  assign sel_963420 = array_index_963163 == array_index_948871 ? add_963419 : sel_963416;
  assign add_963423 = sel_963420 + 8'h01;
  assign sel_963424 = array_index_963163 == array_index_948877 ? add_963423 : sel_963420;
  assign add_963427 = sel_963424 + 8'h01;
  assign sel_963428 = array_index_963163 == array_index_948883 ? add_963427 : sel_963424;
  assign add_963431 = sel_963428 + 8'h01;
  assign sel_963432 = array_index_963163 == array_index_948889 ? add_963431 : sel_963428;
  assign add_963435 = sel_963432 + 8'h01;
  assign sel_963436 = array_index_963163 == array_index_948895 ? add_963435 : sel_963432;
  assign add_963439 = sel_963436 + 8'h01;
  assign sel_963440 = array_index_963163 == array_index_948901 ? add_963439 : sel_963436;
  assign add_963443 = sel_963440 + 8'h01;
  assign sel_963444 = array_index_963163 == array_index_948907 ? add_963443 : sel_963440;
  assign add_963447 = sel_963444 + 8'h01;
  assign sel_963448 = array_index_963163 == array_index_948913 ? add_963447 : sel_963444;
  assign add_963451 = sel_963448 + 8'h01;
  assign sel_963452 = array_index_963163 == array_index_948919 ? add_963451 : sel_963448;
  assign add_963455 = sel_963452 + 8'h01;
  assign sel_963456 = array_index_963163 == array_index_948925 ? add_963455 : sel_963452;
  assign add_963459 = sel_963456 + 8'h01;
  assign sel_963460 = array_index_963163 == array_index_948931 ? add_963459 : sel_963456;
  assign add_963463 = sel_963460 + 8'h01;
  assign sel_963464 = array_index_963163 == array_index_948937 ? add_963463 : sel_963460;
  assign add_963467 = sel_963464 + 8'h01;
  assign sel_963468 = array_index_963163 == array_index_948943 ? add_963467 : sel_963464;
  assign add_963471 = sel_963468 + 8'h01;
  assign sel_963472 = array_index_963163 == array_index_948949 ? add_963471 : sel_963468;
  assign add_963475 = sel_963472 + 8'h01;
  assign sel_963476 = array_index_963163 == array_index_948955 ? add_963475 : sel_963472;
  assign add_963479 = sel_963476 + 8'h01;
  assign sel_963480 = array_index_963163 == array_index_948961 ? add_963479 : sel_963476;
  assign add_963483 = sel_963480 + 8'h01;
  assign sel_963484 = array_index_963163 == array_index_948967 ? add_963483 : sel_963480;
  assign add_963487 = sel_963484 + 8'h01;
  assign sel_963488 = array_index_963163 == array_index_948973 ? add_963487 : sel_963484;
  assign add_963491 = sel_963488 + 8'h01;
  assign sel_963492 = array_index_963163 == array_index_948979 ? add_963491 : sel_963488;
  assign add_963495 = sel_963492 + 8'h01;
  assign sel_963496 = array_index_963163 == array_index_948985 ? add_963495 : sel_963492;
  assign add_963499 = sel_963496 + 8'h01;
  assign sel_963500 = array_index_963163 == array_index_948991 ? add_963499 : sel_963496;
  assign add_963503 = sel_963500 + 8'h01;
  assign sel_963504 = array_index_963163 == array_index_948997 ? add_963503 : sel_963500;
  assign add_963507 = sel_963504 + 8'h01;
  assign sel_963508 = array_index_963163 == array_index_949003 ? add_963507 : sel_963504;
  assign add_963511 = sel_963508 + 8'h01;
  assign sel_963512 = array_index_963163 == array_index_949009 ? add_963511 : sel_963508;
  assign add_963515 = sel_963512 + 8'h01;
  assign sel_963516 = array_index_963163 == array_index_949015 ? add_963515 : sel_963512;
  assign add_963519 = sel_963516 + 8'h01;
  assign sel_963520 = array_index_963163 == array_index_949021 ? add_963519 : sel_963516;
  assign add_963523 = sel_963520 + 8'h01;
  assign sel_963524 = array_index_963163 == array_index_949027 ? add_963523 : sel_963520;
  assign add_963527 = sel_963524 + 8'h01;
  assign sel_963528 = array_index_963163 == array_index_949033 ? add_963527 : sel_963524;
  assign add_963531 = sel_963528 + 8'h01;
  assign sel_963532 = array_index_963163 == array_index_949039 ? add_963531 : sel_963528;
  assign add_963535 = sel_963532 + 8'h01;
  assign sel_963536 = array_index_963163 == array_index_949045 ? add_963535 : sel_963532;
  assign add_963539 = sel_963536 + 8'h01;
  assign sel_963540 = array_index_963163 == array_index_949051 ? add_963539 : sel_963536;
  assign add_963543 = sel_963540 + 8'h01;
  assign sel_963544 = array_index_963163 == array_index_949057 ? add_963543 : sel_963540;
  assign add_963547 = sel_963544 + 8'h01;
  assign sel_963548 = array_index_963163 == array_index_949063 ? add_963547 : sel_963544;
  assign add_963551 = sel_963548 + 8'h01;
  assign sel_963552 = array_index_963163 == array_index_949069 ? add_963551 : sel_963548;
  assign add_963555 = sel_963552 + 8'h01;
  assign sel_963556 = array_index_963163 == array_index_949075 ? add_963555 : sel_963552;
  assign add_963559 = sel_963556 + 8'h01;
  assign sel_963560 = array_index_963163 == array_index_949081 ? add_963559 : sel_963556;
  assign add_963564 = sel_963560 + 8'h01;
  assign array_index_963565 = set1_unflattened[7'h25];
  assign sel_963566 = array_index_963163 == array_index_949087 ? add_963564 : sel_963560;
  assign add_963569 = sel_963566 + 8'h01;
  assign sel_963570 = array_index_963565 == array_index_948483 ? add_963569 : sel_963566;
  assign add_963573 = sel_963570 + 8'h01;
  assign sel_963574 = array_index_963565 == array_index_948487 ? add_963573 : sel_963570;
  assign add_963577 = sel_963574 + 8'h01;
  assign sel_963578 = array_index_963565 == array_index_948495 ? add_963577 : sel_963574;
  assign add_963581 = sel_963578 + 8'h01;
  assign sel_963582 = array_index_963565 == array_index_948503 ? add_963581 : sel_963578;
  assign add_963585 = sel_963582 + 8'h01;
  assign sel_963586 = array_index_963565 == array_index_948511 ? add_963585 : sel_963582;
  assign add_963589 = sel_963586 + 8'h01;
  assign sel_963590 = array_index_963565 == array_index_948519 ? add_963589 : sel_963586;
  assign add_963593 = sel_963590 + 8'h01;
  assign sel_963594 = array_index_963565 == array_index_948527 ? add_963593 : sel_963590;
  assign add_963597 = sel_963594 + 8'h01;
  assign sel_963598 = array_index_963565 == array_index_948535 ? add_963597 : sel_963594;
  assign add_963601 = sel_963598 + 8'h01;
  assign sel_963602 = array_index_963565 == array_index_948541 ? add_963601 : sel_963598;
  assign add_963605 = sel_963602 + 8'h01;
  assign sel_963606 = array_index_963565 == array_index_948547 ? add_963605 : sel_963602;
  assign add_963609 = sel_963606 + 8'h01;
  assign sel_963610 = array_index_963565 == array_index_948553 ? add_963609 : sel_963606;
  assign add_963613 = sel_963610 + 8'h01;
  assign sel_963614 = array_index_963565 == array_index_948559 ? add_963613 : sel_963610;
  assign add_963617 = sel_963614 + 8'h01;
  assign sel_963618 = array_index_963565 == array_index_948565 ? add_963617 : sel_963614;
  assign add_963621 = sel_963618 + 8'h01;
  assign sel_963622 = array_index_963565 == array_index_948571 ? add_963621 : sel_963618;
  assign add_963625 = sel_963622 + 8'h01;
  assign sel_963626 = array_index_963565 == array_index_948577 ? add_963625 : sel_963622;
  assign add_963629 = sel_963626 + 8'h01;
  assign sel_963630 = array_index_963565 == array_index_948583 ? add_963629 : sel_963626;
  assign add_963633 = sel_963630 + 8'h01;
  assign sel_963634 = array_index_963565 == array_index_948589 ? add_963633 : sel_963630;
  assign add_963637 = sel_963634 + 8'h01;
  assign sel_963638 = array_index_963565 == array_index_948595 ? add_963637 : sel_963634;
  assign add_963641 = sel_963638 + 8'h01;
  assign sel_963642 = array_index_963565 == array_index_948601 ? add_963641 : sel_963638;
  assign add_963645 = sel_963642 + 8'h01;
  assign sel_963646 = array_index_963565 == array_index_948607 ? add_963645 : sel_963642;
  assign add_963649 = sel_963646 + 8'h01;
  assign sel_963650 = array_index_963565 == array_index_948613 ? add_963649 : sel_963646;
  assign add_963653 = sel_963650 + 8'h01;
  assign sel_963654 = array_index_963565 == array_index_948619 ? add_963653 : sel_963650;
  assign add_963657 = sel_963654 + 8'h01;
  assign sel_963658 = array_index_963565 == array_index_948625 ? add_963657 : sel_963654;
  assign add_963661 = sel_963658 + 8'h01;
  assign sel_963662 = array_index_963565 == array_index_948631 ? add_963661 : sel_963658;
  assign add_963665 = sel_963662 + 8'h01;
  assign sel_963666 = array_index_963565 == array_index_948637 ? add_963665 : sel_963662;
  assign add_963669 = sel_963666 + 8'h01;
  assign sel_963670 = array_index_963565 == array_index_948643 ? add_963669 : sel_963666;
  assign add_963673 = sel_963670 + 8'h01;
  assign sel_963674 = array_index_963565 == array_index_948649 ? add_963673 : sel_963670;
  assign add_963677 = sel_963674 + 8'h01;
  assign sel_963678 = array_index_963565 == array_index_948655 ? add_963677 : sel_963674;
  assign add_963681 = sel_963678 + 8'h01;
  assign sel_963682 = array_index_963565 == array_index_948661 ? add_963681 : sel_963678;
  assign add_963685 = sel_963682 + 8'h01;
  assign sel_963686 = array_index_963565 == array_index_948667 ? add_963685 : sel_963682;
  assign add_963689 = sel_963686 + 8'h01;
  assign sel_963690 = array_index_963565 == array_index_948673 ? add_963689 : sel_963686;
  assign add_963693 = sel_963690 + 8'h01;
  assign sel_963694 = array_index_963565 == array_index_948679 ? add_963693 : sel_963690;
  assign add_963697 = sel_963694 + 8'h01;
  assign sel_963698 = array_index_963565 == array_index_948685 ? add_963697 : sel_963694;
  assign add_963701 = sel_963698 + 8'h01;
  assign sel_963702 = array_index_963565 == array_index_948691 ? add_963701 : sel_963698;
  assign add_963705 = sel_963702 + 8'h01;
  assign sel_963706 = array_index_963565 == array_index_948697 ? add_963705 : sel_963702;
  assign add_963709 = sel_963706 + 8'h01;
  assign sel_963710 = array_index_963565 == array_index_948703 ? add_963709 : sel_963706;
  assign add_963713 = sel_963710 + 8'h01;
  assign sel_963714 = array_index_963565 == array_index_948709 ? add_963713 : sel_963710;
  assign add_963717 = sel_963714 + 8'h01;
  assign sel_963718 = array_index_963565 == array_index_948715 ? add_963717 : sel_963714;
  assign add_963721 = sel_963718 + 8'h01;
  assign sel_963722 = array_index_963565 == array_index_948721 ? add_963721 : sel_963718;
  assign add_963725 = sel_963722 + 8'h01;
  assign sel_963726 = array_index_963565 == array_index_948727 ? add_963725 : sel_963722;
  assign add_963729 = sel_963726 + 8'h01;
  assign sel_963730 = array_index_963565 == array_index_948733 ? add_963729 : sel_963726;
  assign add_963733 = sel_963730 + 8'h01;
  assign sel_963734 = array_index_963565 == array_index_948739 ? add_963733 : sel_963730;
  assign add_963737 = sel_963734 + 8'h01;
  assign sel_963738 = array_index_963565 == array_index_948745 ? add_963737 : sel_963734;
  assign add_963741 = sel_963738 + 8'h01;
  assign sel_963742 = array_index_963565 == array_index_948751 ? add_963741 : sel_963738;
  assign add_963745 = sel_963742 + 8'h01;
  assign sel_963746 = array_index_963565 == array_index_948757 ? add_963745 : sel_963742;
  assign add_963749 = sel_963746 + 8'h01;
  assign sel_963750 = array_index_963565 == array_index_948763 ? add_963749 : sel_963746;
  assign add_963753 = sel_963750 + 8'h01;
  assign sel_963754 = array_index_963565 == array_index_948769 ? add_963753 : sel_963750;
  assign add_963757 = sel_963754 + 8'h01;
  assign sel_963758 = array_index_963565 == array_index_948775 ? add_963757 : sel_963754;
  assign add_963761 = sel_963758 + 8'h01;
  assign sel_963762 = array_index_963565 == array_index_948781 ? add_963761 : sel_963758;
  assign add_963765 = sel_963762 + 8'h01;
  assign sel_963766 = array_index_963565 == array_index_948787 ? add_963765 : sel_963762;
  assign add_963769 = sel_963766 + 8'h01;
  assign sel_963770 = array_index_963565 == array_index_948793 ? add_963769 : sel_963766;
  assign add_963773 = sel_963770 + 8'h01;
  assign sel_963774 = array_index_963565 == array_index_948799 ? add_963773 : sel_963770;
  assign add_963777 = sel_963774 + 8'h01;
  assign sel_963778 = array_index_963565 == array_index_948805 ? add_963777 : sel_963774;
  assign add_963781 = sel_963778 + 8'h01;
  assign sel_963782 = array_index_963565 == array_index_948811 ? add_963781 : sel_963778;
  assign add_963785 = sel_963782 + 8'h01;
  assign sel_963786 = array_index_963565 == array_index_948817 ? add_963785 : sel_963782;
  assign add_963789 = sel_963786 + 8'h01;
  assign sel_963790 = array_index_963565 == array_index_948823 ? add_963789 : sel_963786;
  assign add_963793 = sel_963790 + 8'h01;
  assign sel_963794 = array_index_963565 == array_index_948829 ? add_963793 : sel_963790;
  assign add_963797 = sel_963794 + 8'h01;
  assign sel_963798 = array_index_963565 == array_index_948835 ? add_963797 : sel_963794;
  assign add_963801 = sel_963798 + 8'h01;
  assign sel_963802 = array_index_963565 == array_index_948841 ? add_963801 : sel_963798;
  assign add_963805 = sel_963802 + 8'h01;
  assign sel_963806 = array_index_963565 == array_index_948847 ? add_963805 : sel_963802;
  assign add_963809 = sel_963806 + 8'h01;
  assign sel_963810 = array_index_963565 == array_index_948853 ? add_963809 : sel_963806;
  assign add_963813 = sel_963810 + 8'h01;
  assign sel_963814 = array_index_963565 == array_index_948859 ? add_963813 : sel_963810;
  assign add_963817 = sel_963814 + 8'h01;
  assign sel_963818 = array_index_963565 == array_index_948865 ? add_963817 : sel_963814;
  assign add_963821 = sel_963818 + 8'h01;
  assign sel_963822 = array_index_963565 == array_index_948871 ? add_963821 : sel_963818;
  assign add_963825 = sel_963822 + 8'h01;
  assign sel_963826 = array_index_963565 == array_index_948877 ? add_963825 : sel_963822;
  assign add_963829 = sel_963826 + 8'h01;
  assign sel_963830 = array_index_963565 == array_index_948883 ? add_963829 : sel_963826;
  assign add_963833 = sel_963830 + 8'h01;
  assign sel_963834 = array_index_963565 == array_index_948889 ? add_963833 : sel_963830;
  assign add_963837 = sel_963834 + 8'h01;
  assign sel_963838 = array_index_963565 == array_index_948895 ? add_963837 : sel_963834;
  assign add_963841 = sel_963838 + 8'h01;
  assign sel_963842 = array_index_963565 == array_index_948901 ? add_963841 : sel_963838;
  assign add_963845 = sel_963842 + 8'h01;
  assign sel_963846 = array_index_963565 == array_index_948907 ? add_963845 : sel_963842;
  assign add_963849 = sel_963846 + 8'h01;
  assign sel_963850 = array_index_963565 == array_index_948913 ? add_963849 : sel_963846;
  assign add_963853 = sel_963850 + 8'h01;
  assign sel_963854 = array_index_963565 == array_index_948919 ? add_963853 : sel_963850;
  assign add_963857 = sel_963854 + 8'h01;
  assign sel_963858 = array_index_963565 == array_index_948925 ? add_963857 : sel_963854;
  assign add_963861 = sel_963858 + 8'h01;
  assign sel_963862 = array_index_963565 == array_index_948931 ? add_963861 : sel_963858;
  assign add_963865 = sel_963862 + 8'h01;
  assign sel_963866 = array_index_963565 == array_index_948937 ? add_963865 : sel_963862;
  assign add_963869 = sel_963866 + 8'h01;
  assign sel_963870 = array_index_963565 == array_index_948943 ? add_963869 : sel_963866;
  assign add_963873 = sel_963870 + 8'h01;
  assign sel_963874 = array_index_963565 == array_index_948949 ? add_963873 : sel_963870;
  assign add_963877 = sel_963874 + 8'h01;
  assign sel_963878 = array_index_963565 == array_index_948955 ? add_963877 : sel_963874;
  assign add_963881 = sel_963878 + 8'h01;
  assign sel_963882 = array_index_963565 == array_index_948961 ? add_963881 : sel_963878;
  assign add_963885 = sel_963882 + 8'h01;
  assign sel_963886 = array_index_963565 == array_index_948967 ? add_963885 : sel_963882;
  assign add_963889 = sel_963886 + 8'h01;
  assign sel_963890 = array_index_963565 == array_index_948973 ? add_963889 : sel_963886;
  assign add_963893 = sel_963890 + 8'h01;
  assign sel_963894 = array_index_963565 == array_index_948979 ? add_963893 : sel_963890;
  assign add_963897 = sel_963894 + 8'h01;
  assign sel_963898 = array_index_963565 == array_index_948985 ? add_963897 : sel_963894;
  assign add_963901 = sel_963898 + 8'h01;
  assign sel_963902 = array_index_963565 == array_index_948991 ? add_963901 : sel_963898;
  assign add_963905 = sel_963902 + 8'h01;
  assign sel_963906 = array_index_963565 == array_index_948997 ? add_963905 : sel_963902;
  assign add_963909 = sel_963906 + 8'h01;
  assign sel_963910 = array_index_963565 == array_index_949003 ? add_963909 : sel_963906;
  assign add_963913 = sel_963910 + 8'h01;
  assign sel_963914 = array_index_963565 == array_index_949009 ? add_963913 : sel_963910;
  assign add_963917 = sel_963914 + 8'h01;
  assign sel_963918 = array_index_963565 == array_index_949015 ? add_963917 : sel_963914;
  assign add_963921 = sel_963918 + 8'h01;
  assign sel_963922 = array_index_963565 == array_index_949021 ? add_963921 : sel_963918;
  assign add_963925 = sel_963922 + 8'h01;
  assign sel_963926 = array_index_963565 == array_index_949027 ? add_963925 : sel_963922;
  assign add_963929 = sel_963926 + 8'h01;
  assign sel_963930 = array_index_963565 == array_index_949033 ? add_963929 : sel_963926;
  assign add_963933 = sel_963930 + 8'h01;
  assign sel_963934 = array_index_963565 == array_index_949039 ? add_963933 : sel_963930;
  assign add_963937 = sel_963934 + 8'h01;
  assign sel_963938 = array_index_963565 == array_index_949045 ? add_963937 : sel_963934;
  assign add_963941 = sel_963938 + 8'h01;
  assign sel_963942 = array_index_963565 == array_index_949051 ? add_963941 : sel_963938;
  assign add_963945 = sel_963942 + 8'h01;
  assign sel_963946 = array_index_963565 == array_index_949057 ? add_963945 : sel_963942;
  assign add_963949 = sel_963946 + 8'h01;
  assign sel_963950 = array_index_963565 == array_index_949063 ? add_963949 : sel_963946;
  assign add_963953 = sel_963950 + 8'h01;
  assign sel_963954 = array_index_963565 == array_index_949069 ? add_963953 : sel_963950;
  assign add_963957 = sel_963954 + 8'h01;
  assign sel_963958 = array_index_963565 == array_index_949075 ? add_963957 : sel_963954;
  assign add_963961 = sel_963958 + 8'h01;
  assign sel_963962 = array_index_963565 == array_index_949081 ? add_963961 : sel_963958;
  assign add_963966 = sel_963962 + 8'h01;
  assign array_index_963967 = set1_unflattened[7'h26];
  assign sel_963968 = array_index_963565 == array_index_949087 ? add_963966 : sel_963962;
  assign add_963971 = sel_963968 + 8'h01;
  assign sel_963972 = array_index_963967 == array_index_948483 ? add_963971 : sel_963968;
  assign add_963975 = sel_963972 + 8'h01;
  assign sel_963976 = array_index_963967 == array_index_948487 ? add_963975 : sel_963972;
  assign add_963979 = sel_963976 + 8'h01;
  assign sel_963980 = array_index_963967 == array_index_948495 ? add_963979 : sel_963976;
  assign add_963983 = sel_963980 + 8'h01;
  assign sel_963984 = array_index_963967 == array_index_948503 ? add_963983 : sel_963980;
  assign add_963987 = sel_963984 + 8'h01;
  assign sel_963988 = array_index_963967 == array_index_948511 ? add_963987 : sel_963984;
  assign add_963991 = sel_963988 + 8'h01;
  assign sel_963992 = array_index_963967 == array_index_948519 ? add_963991 : sel_963988;
  assign add_963995 = sel_963992 + 8'h01;
  assign sel_963996 = array_index_963967 == array_index_948527 ? add_963995 : sel_963992;
  assign add_963999 = sel_963996 + 8'h01;
  assign sel_964000 = array_index_963967 == array_index_948535 ? add_963999 : sel_963996;
  assign add_964003 = sel_964000 + 8'h01;
  assign sel_964004 = array_index_963967 == array_index_948541 ? add_964003 : sel_964000;
  assign add_964007 = sel_964004 + 8'h01;
  assign sel_964008 = array_index_963967 == array_index_948547 ? add_964007 : sel_964004;
  assign add_964011 = sel_964008 + 8'h01;
  assign sel_964012 = array_index_963967 == array_index_948553 ? add_964011 : sel_964008;
  assign add_964015 = sel_964012 + 8'h01;
  assign sel_964016 = array_index_963967 == array_index_948559 ? add_964015 : sel_964012;
  assign add_964019 = sel_964016 + 8'h01;
  assign sel_964020 = array_index_963967 == array_index_948565 ? add_964019 : sel_964016;
  assign add_964023 = sel_964020 + 8'h01;
  assign sel_964024 = array_index_963967 == array_index_948571 ? add_964023 : sel_964020;
  assign add_964027 = sel_964024 + 8'h01;
  assign sel_964028 = array_index_963967 == array_index_948577 ? add_964027 : sel_964024;
  assign add_964031 = sel_964028 + 8'h01;
  assign sel_964032 = array_index_963967 == array_index_948583 ? add_964031 : sel_964028;
  assign add_964035 = sel_964032 + 8'h01;
  assign sel_964036 = array_index_963967 == array_index_948589 ? add_964035 : sel_964032;
  assign add_964039 = sel_964036 + 8'h01;
  assign sel_964040 = array_index_963967 == array_index_948595 ? add_964039 : sel_964036;
  assign add_964043 = sel_964040 + 8'h01;
  assign sel_964044 = array_index_963967 == array_index_948601 ? add_964043 : sel_964040;
  assign add_964047 = sel_964044 + 8'h01;
  assign sel_964048 = array_index_963967 == array_index_948607 ? add_964047 : sel_964044;
  assign add_964051 = sel_964048 + 8'h01;
  assign sel_964052 = array_index_963967 == array_index_948613 ? add_964051 : sel_964048;
  assign add_964055 = sel_964052 + 8'h01;
  assign sel_964056 = array_index_963967 == array_index_948619 ? add_964055 : sel_964052;
  assign add_964059 = sel_964056 + 8'h01;
  assign sel_964060 = array_index_963967 == array_index_948625 ? add_964059 : sel_964056;
  assign add_964063 = sel_964060 + 8'h01;
  assign sel_964064 = array_index_963967 == array_index_948631 ? add_964063 : sel_964060;
  assign add_964067 = sel_964064 + 8'h01;
  assign sel_964068 = array_index_963967 == array_index_948637 ? add_964067 : sel_964064;
  assign add_964071 = sel_964068 + 8'h01;
  assign sel_964072 = array_index_963967 == array_index_948643 ? add_964071 : sel_964068;
  assign add_964075 = sel_964072 + 8'h01;
  assign sel_964076 = array_index_963967 == array_index_948649 ? add_964075 : sel_964072;
  assign add_964079 = sel_964076 + 8'h01;
  assign sel_964080 = array_index_963967 == array_index_948655 ? add_964079 : sel_964076;
  assign add_964083 = sel_964080 + 8'h01;
  assign sel_964084 = array_index_963967 == array_index_948661 ? add_964083 : sel_964080;
  assign add_964087 = sel_964084 + 8'h01;
  assign sel_964088 = array_index_963967 == array_index_948667 ? add_964087 : sel_964084;
  assign add_964091 = sel_964088 + 8'h01;
  assign sel_964092 = array_index_963967 == array_index_948673 ? add_964091 : sel_964088;
  assign add_964095 = sel_964092 + 8'h01;
  assign sel_964096 = array_index_963967 == array_index_948679 ? add_964095 : sel_964092;
  assign add_964099 = sel_964096 + 8'h01;
  assign sel_964100 = array_index_963967 == array_index_948685 ? add_964099 : sel_964096;
  assign add_964103 = sel_964100 + 8'h01;
  assign sel_964104 = array_index_963967 == array_index_948691 ? add_964103 : sel_964100;
  assign add_964107 = sel_964104 + 8'h01;
  assign sel_964108 = array_index_963967 == array_index_948697 ? add_964107 : sel_964104;
  assign add_964111 = sel_964108 + 8'h01;
  assign sel_964112 = array_index_963967 == array_index_948703 ? add_964111 : sel_964108;
  assign add_964115 = sel_964112 + 8'h01;
  assign sel_964116 = array_index_963967 == array_index_948709 ? add_964115 : sel_964112;
  assign add_964119 = sel_964116 + 8'h01;
  assign sel_964120 = array_index_963967 == array_index_948715 ? add_964119 : sel_964116;
  assign add_964123 = sel_964120 + 8'h01;
  assign sel_964124 = array_index_963967 == array_index_948721 ? add_964123 : sel_964120;
  assign add_964127 = sel_964124 + 8'h01;
  assign sel_964128 = array_index_963967 == array_index_948727 ? add_964127 : sel_964124;
  assign add_964131 = sel_964128 + 8'h01;
  assign sel_964132 = array_index_963967 == array_index_948733 ? add_964131 : sel_964128;
  assign add_964135 = sel_964132 + 8'h01;
  assign sel_964136 = array_index_963967 == array_index_948739 ? add_964135 : sel_964132;
  assign add_964139 = sel_964136 + 8'h01;
  assign sel_964140 = array_index_963967 == array_index_948745 ? add_964139 : sel_964136;
  assign add_964143 = sel_964140 + 8'h01;
  assign sel_964144 = array_index_963967 == array_index_948751 ? add_964143 : sel_964140;
  assign add_964147 = sel_964144 + 8'h01;
  assign sel_964148 = array_index_963967 == array_index_948757 ? add_964147 : sel_964144;
  assign add_964151 = sel_964148 + 8'h01;
  assign sel_964152 = array_index_963967 == array_index_948763 ? add_964151 : sel_964148;
  assign add_964155 = sel_964152 + 8'h01;
  assign sel_964156 = array_index_963967 == array_index_948769 ? add_964155 : sel_964152;
  assign add_964159 = sel_964156 + 8'h01;
  assign sel_964160 = array_index_963967 == array_index_948775 ? add_964159 : sel_964156;
  assign add_964163 = sel_964160 + 8'h01;
  assign sel_964164 = array_index_963967 == array_index_948781 ? add_964163 : sel_964160;
  assign add_964167 = sel_964164 + 8'h01;
  assign sel_964168 = array_index_963967 == array_index_948787 ? add_964167 : sel_964164;
  assign add_964171 = sel_964168 + 8'h01;
  assign sel_964172 = array_index_963967 == array_index_948793 ? add_964171 : sel_964168;
  assign add_964175 = sel_964172 + 8'h01;
  assign sel_964176 = array_index_963967 == array_index_948799 ? add_964175 : sel_964172;
  assign add_964179 = sel_964176 + 8'h01;
  assign sel_964180 = array_index_963967 == array_index_948805 ? add_964179 : sel_964176;
  assign add_964183 = sel_964180 + 8'h01;
  assign sel_964184 = array_index_963967 == array_index_948811 ? add_964183 : sel_964180;
  assign add_964187 = sel_964184 + 8'h01;
  assign sel_964188 = array_index_963967 == array_index_948817 ? add_964187 : sel_964184;
  assign add_964191 = sel_964188 + 8'h01;
  assign sel_964192 = array_index_963967 == array_index_948823 ? add_964191 : sel_964188;
  assign add_964195 = sel_964192 + 8'h01;
  assign sel_964196 = array_index_963967 == array_index_948829 ? add_964195 : sel_964192;
  assign add_964199 = sel_964196 + 8'h01;
  assign sel_964200 = array_index_963967 == array_index_948835 ? add_964199 : sel_964196;
  assign add_964203 = sel_964200 + 8'h01;
  assign sel_964204 = array_index_963967 == array_index_948841 ? add_964203 : sel_964200;
  assign add_964207 = sel_964204 + 8'h01;
  assign sel_964208 = array_index_963967 == array_index_948847 ? add_964207 : sel_964204;
  assign add_964211 = sel_964208 + 8'h01;
  assign sel_964212 = array_index_963967 == array_index_948853 ? add_964211 : sel_964208;
  assign add_964215 = sel_964212 + 8'h01;
  assign sel_964216 = array_index_963967 == array_index_948859 ? add_964215 : sel_964212;
  assign add_964219 = sel_964216 + 8'h01;
  assign sel_964220 = array_index_963967 == array_index_948865 ? add_964219 : sel_964216;
  assign add_964223 = sel_964220 + 8'h01;
  assign sel_964224 = array_index_963967 == array_index_948871 ? add_964223 : sel_964220;
  assign add_964227 = sel_964224 + 8'h01;
  assign sel_964228 = array_index_963967 == array_index_948877 ? add_964227 : sel_964224;
  assign add_964231 = sel_964228 + 8'h01;
  assign sel_964232 = array_index_963967 == array_index_948883 ? add_964231 : sel_964228;
  assign add_964235 = sel_964232 + 8'h01;
  assign sel_964236 = array_index_963967 == array_index_948889 ? add_964235 : sel_964232;
  assign add_964239 = sel_964236 + 8'h01;
  assign sel_964240 = array_index_963967 == array_index_948895 ? add_964239 : sel_964236;
  assign add_964243 = sel_964240 + 8'h01;
  assign sel_964244 = array_index_963967 == array_index_948901 ? add_964243 : sel_964240;
  assign add_964247 = sel_964244 + 8'h01;
  assign sel_964248 = array_index_963967 == array_index_948907 ? add_964247 : sel_964244;
  assign add_964251 = sel_964248 + 8'h01;
  assign sel_964252 = array_index_963967 == array_index_948913 ? add_964251 : sel_964248;
  assign add_964255 = sel_964252 + 8'h01;
  assign sel_964256 = array_index_963967 == array_index_948919 ? add_964255 : sel_964252;
  assign add_964259 = sel_964256 + 8'h01;
  assign sel_964260 = array_index_963967 == array_index_948925 ? add_964259 : sel_964256;
  assign add_964263 = sel_964260 + 8'h01;
  assign sel_964264 = array_index_963967 == array_index_948931 ? add_964263 : sel_964260;
  assign add_964267 = sel_964264 + 8'h01;
  assign sel_964268 = array_index_963967 == array_index_948937 ? add_964267 : sel_964264;
  assign add_964271 = sel_964268 + 8'h01;
  assign sel_964272 = array_index_963967 == array_index_948943 ? add_964271 : sel_964268;
  assign add_964275 = sel_964272 + 8'h01;
  assign sel_964276 = array_index_963967 == array_index_948949 ? add_964275 : sel_964272;
  assign add_964279 = sel_964276 + 8'h01;
  assign sel_964280 = array_index_963967 == array_index_948955 ? add_964279 : sel_964276;
  assign add_964283 = sel_964280 + 8'h01;
  assign sel_964284 = array_index_963967 == array_index_948961 ? add_964283 : sel_964280;
  assign add_964287 = sel_964284 + 8'h01;
  assign sel_964288 = array_index_963967 == array_index_948967 ? add_964287 : sel_964284;
  assign add_964291 = sel_964288 + 8'h01;
  assign sel_964292 = array_index_963967 == array_index_948973 ? add_964291 : sel_964288;
  assign add_964295 = sel_964292 + 8'h01;
  assign sel_964296 = array_index_963967 == array_index_948979 ? add_964295 : sel_964292;
  assign add_964299 = sel_964296 + 8'h01;
  assign sel_964300 = array_index_963967 == array_index_948985 ? add_964299 : sel_964296;
  assign add_964303 = sel_964300 + 8'h01;
  assign sel_964304 = array_index_963967 == array_index_948991 ? add_964303 : sel_964300;
  assign add_964307 = sel_964304 + 8'h01;
  assign sel_964308 = array_index_963967 == array_index_948997 ? add_964307 : sel_964304;
  assign add_964311 = sel_964308 + 8'h01;
  assign sel_964312 = array_index_963967 == array_index_949003 ? add_964311 : sel_964308;
  assign add_964315 = sel_964312 + 8'h01;
  assign sel_964316 = array_index_963967 == array_index_949009 ? add_964315 : sel_964312;
  assign add_964319 = sel_964316 + 8'h01;
  assign sel_964320 = array_index_963967 == array_index_949015 ? add_964319 : sel_964316;
  assign add_964323 = sel_964320 + 8'h01;
  assign sel_964324 = array_index_963967 == array_index_949021 ? add_964323 : sel_964320;
  assign add_964327 = sel_964324 + 8'h01;
  assign sel_964328 = array_index_963967 == array_index_949027 ? add_964327 : sel_964324;
  assign add_964331 = sel_964328 + 8'h01;
  assign sel_964332 = array_index_963967 == array_index_949033 ? add_964331 : sel_964328;
  assign add_964335 = sel_964332 + 8'h01;
  assign sel_964336 = array_index_963967 == array_index_949039 ? add_964335 : sel_964332;
  assign add_964339 = sel_964336 + 8'h01;
  assign sel_964340 = array_index_963967 == array_index_949045 ? add_964339 : sel_964336;
  assign add_964343 = sel_964340 + 8'h01;
  assign sel_964344 = array_index_963967 == array_index_949051 ? add_964343 : sel_964340;
  assign add_964347 = sel_964344 + 8'h01;
  assign sel_964348 = array_index_963967 == array_index_949057 ? add_964347 : sel_964344;
  assign add_964351 = sel_964348 + 8'h01;
  assign sel_964352 = array_index_963967 == array_index_949063 ? add_964351 : sel_964348;
  assign add_964355 = sel_964352 + 8'h01;
  assign sel_964356 = array_index_963967 == array_index_949069 ? add_964355 : sel_964352;
  assign add_964359 = sel_964356 + 8'h01;
  assign sel_964360 = array_index_963967 == array_index_949075 ? add_964359 : sel_964356;
  assign add_964363 = sel_964360 + 8'h01;
  assign sel_964364 = array_index_963967 == array_index_949081 ? add_964363 : sel_964360;
  assign add_964368 = sel_964364 + 8'h01;
  assign array_index_964369 = set1_unflattened[7'h27];
  assign sel_964370 = array_index_963967 == array_index_949087 ? add_964368 : sel_964364;
  assign add_964373 = sel_964370 + 8'h01;
  assign sel_964374 = array_index_964369 == array_index_948483 ? add_964373 : sel_964370;
  assign add_964377 = sel_964374 + 8'h01;
  assign sel_964378 = array_index_964369 == array_index_948487 ? add_964377 : sel_964374;
  assign add_964381 = sel_964378 + 8'h01;
  assign sel_964382 = array_index_964369 == array_index_948495 ? add_964381 : sel_964378;
  assign add_964385 = sel_964382 + 8'h01;
  assign sel_964386 = array_index_964369 == array_index_948503 ? add_964385 : sel_964382;
  assign add_964389 = sel_964386 + 8'h01;
  assign sel_964390 = array_index_964369 == array_index_948511 ? add_964389 : sel_964386;
  assign add_964393 = sel_964390 + 8'h01;
  assign sel_964394 = array_index_964369 == array_index_948519 ? add_964393 : sel_964390;
  assign add_964397 = sel_964394 + 8'h01;
  assign sel_964398 = array_index_964369 == array_index_948527 ? add_964397 : sel_964394;
  assign add_964401 = sel_964398 + 8'h01;
  assign sel_964402 = array_index_964369 == array_index_948535 ? add_964401 : sel_964398;
  assign add_964405 = sel_964402 + 8'h01;
  assign sel_964406 = array_index_964369 == array_index_948541 ? add_964405 : sel_964402;
  assign add_964409 = sel_964406 + 8'h01;
  assign sel_964410 = array_index_964369 == array_index_948547 ? add_964409 : sel_964406;
  assign add_964413 = sel_964410 + 8'h01;
  assign sel_964414 = array_index_964369 == array_index_948553 ? add_964413 : sel_964410;
  assign add_964417 = sel_964414 + 8'h01;
  assign sel_964418 = array_index_964369 == array_index_948559 ? add_964417 : sel_964414;
  assign add_964421 = sel_964418 + 8'h01;
  assign sel_964422 = array_index_964369 == array_index_948565 ? add_964421 : sel_964418;
  assign add_964425 = sel_964422 + 8'h01;
  assign sel_964426 = array_index_964369 == array_index_948571 ? add_964425 : sel_964422;
  assign add_964429 = sel_964426 + 8'h01;
  assign sel_964430 = array_index_964369 == array_index_948577 ? add_964429 : sel_964426;
  assign add_964433 = sel_964430 + 8'h01;
  assign sel_964434 = array_index_964369 == array_index_948583 ? add_964433 : sel_964430;
  assign add_964437 = sel_964434 + 8'h01;
  assign sel_964438 = array_index_964369 == array_index_948589 ? add_964437 : sel_964434;
  assign add_964441 = sel_964438 + 8'h01;
  assign sel_964442 = array_index_964369 == array_index_948595 ? add_964441 : sel_964438;
  assign add_964445 = sel_964442 + 8'h01;
  assign sel_964446 = array_index_964369 == array_index_948601 ? add_964445 : sel_964442;
  assign add_964449 = sel_964446 + 8'h01;
  assign sel_964450 = array_index_964369 == array_index_948607 ? add_964449 : sel_964446;
  assign add_964453 = sel_964450 + 8'h01;
  assign sel_964454 = array_index_964369 == array_index_948613 ? add_964453 : sel_964450;
  assign add_964457 = sel_964454 + 8'h01;
  assign sel_964458 = array_index_964369 == array_index_948619 ? add_964457 : sel_964454;
  assign add_964461 = sel_964458 + 8'h01;
  assign sel_964462 = array_index_964369 == array_index_948625 ? add_964461 : sel_964458;
  assign add_964465 = sel_964462 + 8'h01;
  assign sel_964466 = array_index_964369 == array_index_948631 ? add_964465 : sel_964462;
  assign add_964469 = sel_964466 + 8'h01;
  assign sel_964470 = array_index_964369 == array_index_948637 ? add_964469 : sel_964466;
  assign add_964473 = sel_964470 + 8'h01;
  assign sel_964474 = array_index_964369 == array_index_948643 ? add_964473 : sel_964470;
  assign add_964477 = sel_964474 + 8'h01;
  assign sel_964478 = array_index_964369 == array_index_948649 ? add_964477 : sel_964474;
  assign add_964481 = sel_964478 + 8'h01;
  assign sel_964482 = array_index_964369 == array_index_948655 ? add_964481 : sel_964478;
  assign add_964485 = sel_964482 + 8'h01;
  assign sel_964486 = array_index_964369 == array_index_948661 ? add_964485 : sel_964482;
  assign add_964489 = sel_964486 + 8'h01;
  assign sel_964490 = array_index_964369 == array_index_948667 ? add_964489 : sel_964486;
  assign add_964493 = sel_964490 + 8'h01;
  assign sel_964494 = array_index_964369 == array_index_948673 ? add_964493 : sel_964490;
  assign add_964497 = sel_964494 + 8'h01;
  assign sel_964498 = array_index_964369 == array_index_948679 ? add_964497 : sel_964494;
  assign add_964501 = sel_964498 + 8'h01;
  assign sel_964502 = array_index_964369 == array_index_948685 ? add_964501 : sel_964498;
  assign add_964505 = sel_964502 + 8'h01;
  assign sel_964506 = array_index_964369 == array_index_948691 ? add_964505 : sel_964502;
  assign add_964509 = sel_964506 + 8'h01;
  assign sel_964510 = array_index_964369 == array_index_948697 ? add_964509 : sel_964506;
  assign add_964513 = sel_964510 + 8'h01;
  assign sel_964514 = array_index_964369 == array_index_948703 ? add_964513 : sel_964510;
  assign add_964517 = sel_964514 + 8'h01;
  assign sel_964518 = array_index_964369 == array_index_948709 ? add_964517 : sel_964514;
  assign add_964521 = sel_964518 + 8'h01;
  assign sel_964522 = array_index_964369 == array_index_948715 ? add_964521 : sel_964518;
  assign add_964525 = sel_964522 + 8'h01;
  assign sel_964526 = array_index_964369 == array_index_948721 ? add_964525 : sel_964522;
  assign add_964529 = sel_964526 + 8'h01;
  assign sel_964530 = array_index_964369 == array_index_948727 ? add_964529 : sel_964526;
  assign add_964533 = sel_964530 + 8'h01;
  assign sel_964534 = array_index_964369 == array_index_948733 ? add_964533 : sel_964530;
  assign add_964537 = sel_964534 + 8'h01;
  assign sel_964538 = array_index_964369 == array_index_948739 ? add_964537 : sel_964534;
  assign add_964541 = sel_964538 + 8'h01;
  assign sel_964542 = array_index_964369 == array_index_948745 ? add_964541 : sel_964538;
  assign add_964545 = sel_964542 + 8'h01;
  assign sel_964546 = array_index_964369 == array_index_948751 ? add_964545 : sel_964542;
  assign add_964549 = sel_964546 + 8'h01;
  assign sel_964550 = array_index_964369 == array_index_948757 ? add_964549 : sel_964546;
  assign add_964553 = sel_964550 + 8'h01;
  assign sel_964554 = array_index_964369 == array_index_948763 ? add_964553 : sel_964550;
  assign add_964557 = sel_964554 + 8'h01;
  assign sel_964558 = array_index_964369 == array_index_948769 ? add_964557 : sel_964554;
  assign add_964561 = sel_964558 + 8'h01;
  assign sel_964562 = array_index_964369 == array_index_948775 ? add_964561 : sel_964558;
  assign add_964565 = sel_964562 + 8'h01;
  assign sel_964566 = array_index_964369 == array_index_948781 ? add_964565 : sel_964562;
  assign add_964569 = sel_964566 + 8'h01;
  assign sel_964570 = array_index_964369 == array_index_948787 ? add_964569 : sel_964566;
  assign add_964573 = sel_964570 + 8'h01;
  assign sel_964574 = array_index_964369 == array_index_948793 ? add_964573 : sel_964570;
  assign add_964577 = sel_964574 + 8'h01;
  assign sel_964578 = array_index_964369 == array_index_948799 ? add_964577 : sel_964574;
  assign add_964581 = sel_964578 + 8'h01;
  assign sel_964582 = array_index_964369 == array_index_948805 ? add_964581 : sel_964578;
  assign add_964585 = sel_964582 + 8'h01;
  assign sel_964586 = array_index_964369 == array_index_948811 ? add_964585 : sel_964582;
  assign add_964589 = sel_964586 + 8'h01;
  assign sel_964590 = array_index_964369 == array_index_948817 ? add_964589 : sel_964586;
  assign add_964593 = sel_964590 + 8'h01;
  assign sel_964594 = array_index_964369 == array_index_948823 ? add_964593 : sel_964590;
  assign add_964597 = sel_964594 + 8'h01;
  assign sel_964598 = array_index_964369 == array_index_948829 ? add_964597 : sel_964594;
  assign add_964601 = sel_964598 + 8'h01;
  assign sel_964602 = array_index_964369 == array_index_948835 ? add_964601 : sel_964598;
  assign add_964605 = sel_964602 + 8'h01;
  assign sel_964606 = array_index_964369 == array_index_948841 ? add_964605 : sel_964602;
  assign add_964609 = sel_964606 + 8'h01;
  assign sel_964610 = array_index_964369 == array_index_948847 ? add_964609 : sel_964606;
  assign add_964613 = sel_964610 + 8'h01;
  assign sel_964614 = array_index_964369 == array_index_948853 ? add_964613 : sel_964610;
  assign add_964617 = sel_964614 + 8'h01;
  assign sel_964618 = array_index_964369 == array_index_948859 ? add_964617 : sel_964614;
  assign add_964621 = sel_964618 + 8'h01;
  assign sel_964622 = array_index_964369 == array_index_948865 ? add_964621 : sel_964618;
  assign add_964625 = sel_964622 + 8'h01;
  assign sel_964626 = array_index_964369 == array_index_948871 ? add_964625 : sel_964622;
  assign add_964629 = sel_964626 + 8'h01;
  assign sel_964630 = array_index_964369 == array_index_948877 ? add_964629 : sel_964626;
  assign add_964633 = sel_964630 + 8'h01;
  assign sel_964634 = array_index_964369 == array_index_948883 ? add_964633 : sel_964630;
  assign add_964637 = sel_964634 + 8'h01;
  assign sel_964638 = array_index_964369 == array_index_948889 ? add_964637 : sel_964634;
  assign add_964641 = sel_964638 + 8'h01;
  assign sel_964642 = array_index_964369 == array_index_948895 ? add_964641 : sel_964638;
  assign add_964645 = sel_964642 + 8'h01;
  assign sel_964646 = array_index_964369 == array_index_948901 ? add_964645 : sel_964642;
  assign add_964649 = sel_964646 + 8'h01;
  assign sel_964650 = array_index_964369 == array_index_948907 ? add_964649 : sel_964646;
  assign add_964653 = sel_964650 + 8'h01;
  assign sel_964654 = array_index_964369 == array_index_948913 ? add_964653 : sel_964650;
  assign add_964657 = sel_964654 + 8'h01;
  assign sel_964658 = array_index_964369 == array_index_948919 ? add_964657 : sel_964654;
  assign add_964661 = sel_964658 + 8'h01;
  assign sel_964662 = array_index_964369 == array_index_948925 ? add_964661 : sel_964658;
  assign add_964665 = sel_964662 + 8'h01;
  assign sel_964666 = array_index_964369 == array_index_948931 ? add_964665 : sel_964662;
  assign add_964669 = sel_964666 + 8'h01;
  assign sel_964670 = array_index_964369 == array_index_948937 ? add_964669 : sel_964666;
  assign add_964673 = sel_964670 + 8'h01;
  assign sel_964674 = array_index_964369 == array_index_948943 ? add_964673 : sel_964670;
  assign add_964677 = sel_964674 + 8'h01;
  assign sel_964678 = array_index_964369 == array_index_948949 ? add_964677 : sel_964674;
  assign add_964681 = sel_964678 + 8'h01;
  assign sel_964682 = array_index_964369 == array_index_948955 ? add_964681 : sel_964678;
  assign add_964685 = sel_964682 + 8'h01;
  assign sel_964686 = array_index_964369 == array_index_948961 ? add_964685 : sel_964682;
  assign add_964689 = sel_964686 + 8'h01;
  assign sel_964690 = array_index_964369 == array_index_948967 ? add_964689 : sel_964686;
  assign add_964693 = sel_964690 + 8'h01;
  assign sel_964694 = array_index_964369 == array_index_948973 ? add_964693 : sel_964690;
  assign add_964697 = sel_964694 + 8'h01;
  assign sel_964698 = array_index_964369 == array_index_948979 ? add_964697 : sel_964694;
  assign add_964701 = sel_964698 + 8'h01;
  assign sel_964702 = array_index_964369 == array_index_948985 ? add_964701 : sel_964698;
  assign add_964705 = sel_964702 + 8'h01;
  assign sel_964706 = array_index_964369 == array_index_948991 ? add_964705 : sel_964702;
  assign add_964709 = sel_964706 + 8'h01;
  assign sel_964710 = array_index_964369 == array_index_948997 ? add_964709 : sel_964706;
  assign add_964713 = sel_964710 + 8'h01;
  assign sel_964714 = array_index_964369 == array_index_949003 ? add_964713 : sel_964710;
  assign add_964717 = sel_964714 + 8'h01;
  assign sel_964718 = array_index_964369 == array_index_949009 ? add_964717 : sel_964714;
  assign add_964721 = sel_964718 + 8'h01;
  assign sel_964722 = array_index_964369 == array_index_949015 ? add_964721 : sel_964718;
  assign add_964725 = sel_964722 + 8'h01;
  assign sel_964726 = array_index_964369 == array_index_949021 ? add_964725 : sel_964722;
  assign add_964729 = sel_964726 + 8'h01;
  assign sel_964730 = array_index_964369 == array_index_949027 ? add_964729 : sel_964726;
  assign add_964733 = sel_964730 + 8'h01;
  assign sel_964734 = array_index_964369 == array_index_949033 ? add_964733 : sel_964730;
  assign add_964737 = sel_964734 + 8'h01;
  assign sel_964738 = array_index_964369 == array_index_949039 ? add_964737 : sel_964734;
  assign add_964741 = sel_964738 + 8'h01;
  assign sel_964742 = array_index_964369 == array_index_949045 ? add_964741 : sel_964738;
  assign add_964745 = sel_964742 + 8'h01;
  assign sel_964746 = array_index_964369 == array_index_949051 ? add_964745 : sel_964742;
  assign add_964749 = sel_964746 + 8'h01;
  assign sel_964750 = array_index_964369 == array_index_949057 ? add_964749 : sel_964746;
  assign add_964753 = sel_964750 + 8'h01;
  assign sel_964754 = array_index_964369 == array_index_949063 ? add_964753 : sel_964750;
  assign add_964757 = sel_964754 + 8'h01;
  assign sel_964758 = array_index_964369 == array_index_949069 ? add_964757 : sel_964754;
  assign add_964761 = sel_964758 + 8'h01;
  assign sel_964762 = array_index_964369 == array_index_949075 ? add_964761 : sel_964758;
  assign add_964765 = sel_964762 + 8'h01;
  assign sel_964766 = array_index_964369 == array_index_949081 ? add_964765 : sel_964762;
  assign add_964770 = sel_964766 + 8'h01;
  assign array_index_964771 = set1_unflattened[7'h28];
  assign sel_964772 = array_index_964369 == array_index_949087 ? add_964770 : sel_964766;
  assign add_964775 = sel_964772 + 8'h01;
  assign sel_964776 = array_index_964771 == array_index_948483 ? add_964775 : sel_964772;
  assign add_964779 = sel_964776 + 8'h01;
  assign sel_964780 = array_index_964771 == array_index_948487 ? add_964779 : sel_964776;
  assign add_964783 = sel_964780 + 8'h01;
  assign sel_964784 = array_index_964771 == array_index_948495 ? add_964783 : sel_964780;
  assign add_964787 = sel_964784 + 8'h01;
  assign sel_964788 = array_index_964771 == array_index_948503 ? add_964787 : sel_964784;
  assign add_964791 = sel_964788 + 8'h01;
  assign sel_964792 = array_index_964771 == array_index_948511 ? add_964791 : sel_964788;
  assign add_964795 = sel_964792 + 8'h01;
  assign sel_964796 = array_index_964771 == array_index_948519 ? add_964795 : sel_964792;
  assign add_964799 = sel_964796 + 8'h01;
  assign sel_964800 = array_index_964771 == array_index_948527 ? add_964799 : sel_964796;
  assign add_964803 = sel_964800 + 8'h01;
  assign sel_964804 = array_index_964771 == array_index_948535 ? add_964803 : sel_964800;
  assign add_964807 = sel_964804 + 8'h01;
  assign sel_964808 = array_index_964771 == array_index_948541 ? add_964807 : sel_964804;
  assign add_964811 = sel_964808 + 8'h01;
  assign sel_964812 = array_index_964771 == array_index_948547 ? add_964811 : sel_964808;
  assign add_964815 = sel_964812 + 8'h01;
  assign sel_964816 = array_index_964771 == array_index_948553 ? add_964815 : sel_964812;
  assign add_964819 = sel_964816 + 8'h01;
  assign sel_964820 = array_index_964771 == array_index_948559 ? add_964819 : sel_964816;
  assign add_964823 = sel_964820 + 8'h01;
  assign sel_964824 = array_index_964771 == array_index_948565 ? add_964823 : sel_964820;
  assign add_964827 = sel_964824 + 8'h01;
  assign sel_964828 = array_index_964771 == array_index_948571 ? add_964827 : sel_964824;
  assign add_964831 = sel_964828 + 8'h01;
  assign sel_964832 = array_index_964771 == array_index_948577 ? add_964831 : sel_964828;
  assign add_964835 = sel_964832 + 8'h01;
  assign sel_964836 = array_index_964771 == array_index_948583 ? add_964835 : sel_964832;
  assign add_964839 = sel_964836 + 8'h01;
  assign sel_964840 = array_index_964771 == array_index_948589 ? add_964839 : sel_964836;
  assign add_964843 = sel_964840 + 8'h01;
  assign sel_964844 = array_index_964771 == array_index_948595 ? add_964843 : sel_964840;
  assign add_964847 = sel_964844 + 8'h01;
  assign sel_964848 = array_index_964771 == array_index_948601 ? add_964847 : sel_964844;
  assign add_964851 = sel_964848 + 8'h01;
  assign sel_964852 = array_index_964771 == array_index_948607 ? add_964851 : sel_964848;
  assign add_964855 = sel_964852 + 8'h01;
  assign sel_964856 = array_index_964771 == array_index_948613 ? add_964855 : sel_964852;
  assign add_964859 = sel_964856 + 8'h01;
  assign sel_964860 = array_index_964771 == array_index_948619 ? add_964859 : sel_964856;
  assign add_964863 = sel_964860 + 8'h01;
  assign sel_964864 = array_index_964771 == array_index_948625 ? add_964863 : sel_964860;
  assign add_964867 = sel_964864 + 8'h01;
  assign sel_964868 = array_index_964771 == array_index_948631 ? add_964867 : sel_964864;
  assign add_964871 = sel_964868 + 8'h01;
  assign sel_964872 = array_index_964771 == array_index_948637 ? add_964871 : sel_964868;
  assign add_964875 = sel_964872 + 8'h01;
  assign sel_964876 = array_index_964771 == array_index_948643 ? add_964875 : sel_964872;
  assign add_964879 = sel_964876 + 8'h01;
  assign sel_964880 = array_index_964771 == array_index_948649 ? add_964879 : sel_964876;
  assign add_964883 = sel_964880 + 8'h01;
  assign sel_964884 = array_index_964771 == array_index_948655 ? add_964883 : sel_964880;
  assign add_964887 = sel_964884 + 8'h01;
  assign sel_964888 = array_index_964771 == array_index_948661 ? add_964887 : sel_964884;
  assign add_964891 = sel_964888 + 8'h01;
  assign sel_964892 = array_index_964771 == array_index_948667 ? add_964891 : sel_964888;
  assign add_964895 = sel_964892 + 8'h01;
  assign sel_964896 = array_index_964771 == array_index_948673 ? add_964895 : sel_964892;
  assign add_964899 = sel_964896 + 8'h01;
  assign sel_964900 = array_index_964771 == array_index_948679 ? add_964899 : sel_964896;
  assign add_964903 = sel_964900 + 8'h01;
  assign sel_964904 = array_index_964771 == array_index_948685 ? add_964903 : sel_964900;
  assign add_964907 = sel_964904 + 8'h01;
  assign sel_964908 = array_index_964771 == array_index_948691 ? add_964907 : sel_964904;
  assign add_964911 = sel_964908 + 8'h01;
  assign sel_964912 = array_index_964771 == array_index_948697 ? add_964911 : sel_964908;
  assign add_964915 = sel_964912 + 8'h01;
  assign sel_964916 = array_index_964771 == array_index_948703 ? add_964915 : sel_964912;
  assign add_964919 = sel_964916 + 8'h01;
  assign sel_964920 = array_index_964771 == array_index_948709 ? add_964919 : sel_964916;
  assign add_964923 = sel_964920 + 8'h01;
  assign sel_964924 = array_index_964771 == array_index_948715 ? add_964923 : sel_964920;
  assign add_964927 = sel_964924 + 8'h01;
  assign sel_964928 = array_index_964771 == array_index_948721 ? add_964927 : sel_964924;
  assign add_964931 = sel_964928 + 8'h01;
  assign sel_964932 = array_index_964771 == array_index_948727 ? add_964931 : sel_964928;
  assign add_964935 = sel_964932 + 8'h01;
  assign sel_964936 = array_index_964771 == array_index_948733 ? add_964935 : sel_964932;
  assign add_964939 = sel_964936 + 8'h01;
  assign sel_964940 = array_index_964771 == array_index_948739 ? add_964939 : sel_964936;
  assign add_964943 = sel_964940 + 8'h01;
  assign sel_964944 = array_index_964771 == array_index_948745 ? add_964943 : sel_964940;
  assign add_964947 = sel_964944 + 8'h01;
  assign sel_964948 = array_index_964771 == array_index_948751 ? add_964947 : sel_964944;
  assign add_964951 = sel_964948 + 8'h01;
  assign sel_964952 = array_index_964771 == array_index_948757 ? add_964951 : sel_964948;
  assign add_964955 = sel_964952 + 8'h01;
  assign sel_964956 = array_index_964771 == array_index_948763 ? add_964955 : sel_964952;
  assign add_964959 = sel_964956 + 8'h01;
  assign sel_964960 = array_index_964771 == array_index_948769 ? add_964959 : sel_964956;
  assign add_964963 = sel_964960 + 8'h01;
  assign sel_964964 = array_index_964771 == array_index_948775 ? add_964963 : sel_964960;
  assign add_964967 = sel_964964 + 8'h01;
  assign sel_964968 = array_index_964771 == array_index_948781 ? add_964967 : sel_964964;
  assign add_964971 = sel_964968 + 8'h01;
  assign sel_964972 = array_index_964771 == array_index_948787 ? add_964971 : sel_964968;
  assign add_964975 = sel_964972 + 8'h01;
  assign sel_964976 = array_index_964771 == array_index_948793 ? add_964975 : sel_964972;
  assign add_964979 = sel_964976 + 8'h01;
  assign sel_964980 = array_index_964771 == array_index_948799 ? add_964979 : sel_964976;
  assign add_964983 = sel_964980 + 8'h01;
  assign sel_964984 = array_index_964771 == array_index_948805 ? add_964983 : sel_964980;
  assign add_964987 = sel_964984 + 8'h01;
  assign sel_964988 = array_index_964771 == array_index_948811 ? add_964987 : sel_964984;
  assign add_964991 = sel_964988 + 8'h01;
  assign sel_964992 = array_index_964771 == array_index_948817 ? add_964991 : sel_964988;
  assign add_964995 = sel_964992 + 8'h01;
  assign sel_964996 = array_index_964771 == array_index_948823 ? add_964995 : sel_964992;
  assign add_964999 = sel_964996 + 8'h01;
  assign sel_965000 = array_index_964771 == array_index_948829 ? add_964999 : sel_964996;
  assign add_965003 = sel_965000 + 8'h01;
  assign sel_965004 = array_index_964771 == array_index_948835 ? add_965003 : sel_965000;
  assign add_965007 = sel_965004 + 8'h01;
  assign sel_965008 = array_index_964771 == array_index_948841 ? add_965007 : sel_965004;
  assign add_965011 = sel_965008 + 8'h01;
  assign sel_965012 = array_index_964771 == array_index_948847 ? add_965011 : sel_965008;
  assign add_965015 = sel_965012 + 8'h01;
  assign sel_965016 = array_index_964771 == array_index_948853 ? add_965015 : sel_965012;
  assign add_965019 = sel_965016 + 8'h01;
  assign sel_965020 = array_index_964771 == array_index_948859 ? add_965019 : sel_965016;
  assign add_965023 = sel_965020 + 8'h01;
  assign sel_965024 = array_index_964771 == array_index_948865 ? add_965023 : sel_965020;
  assign add_965027 = sel_965024 + 8'h01;
  assign sel_965028 = array_index_964771 == array_index_948871 ? add_965027 : sel_965024;
  assign add_965031 = sel_965028 + 8'h01;
  assign sel_965032 = array_index_964771 == array_index_948877 ? add_965031 : sel_965028;
  assign add_965035 = sel_965032 + 8'h01;
  assign sel_965036 = array_index_964771 == array_index_948883 ? add_965035 : sel_965032;
  assign add_965039 = sel_965036 + 8'h01;
  assign sel_965040 = array_index_964771 == array_index_948889 ? add_965039 : sel_965036;
  assign add_965043 = sel_965040 + 8'h01;
  assign sel_965044 = array_index_964771 == array_index_948895 ? add_965043 : sel_965040;
  assign add_965047 = sel_965044 + 8'h01;
  assign sel_965048 = array_index_964771 == array_index_948901 ? add_965047 : sel_965044;
  assign add_965051 = sel_965048 + 8'h01;
  assign sel_965052 = array_index_964771 == array_index_948907 ? add_965051 : sel_965048;
  assign add_965055 = sel_965052 + 8'h01;
  assign sel_965056 = array_index_964771 == array_index_948913 ? add_965055 : sel_965052;
  assign add_965059 = sel_965056 + 8'h01;
  assign sel_965060 = array_index_964771 == array_index_948919 ? add_965059 : sel_965056;
  assign add_965063 = sel_965060 + 8'h01;
  assign sel_965064 = array_index_964771 == array_index_948925 ? add_965063 : sel_965060;
  assign add_965067 = sel_965064 + 8'h01;
  assign sel_965068 = array_index_964771 == array_index_948931 ? add_965067 : sel_965064;
  assign add_965071 = sel_965068 + 8'h01;
  assign sel_965072 = array_index_964771 == array_index_948937 ? add_965071 : sel_965068;
  assign add_965075 = sel_965072 + 8'h01;
  assign sel_965076 = array_index_964771 == array_index_948943 ? add_965075 : sel_965072;
  assign add_965079 = sel_965076 + 8'h01;
  assign sel_965080 = array_index_964771 == array_index_948949 ? add_965079 : sel_965076;
  assign add_965083 = sel_965080 + 8'h01;
  assign sel_965084 = array_index_964771 == array_index_948955 ? add_965083 : sel_965080;
  assign add_965087 = sel_965084 + 8'h01;
  assign sel_965088 = array_index_964771 == array_index_948961 ? add_965087 : sel_965084;
  assign add_965091 = sel_965088 + 8'h01;
  assign sel_965092 = array_index_964771 == array_index_948967 ? add_965091 : sel_965088;
  assign add_965095 = sel_965092 + 8'h01;
  assign sel_965096 = array_index_964771 == array_index_948973 ? add_965095 : sel_965092;
  assign add_965099 = sel_965096 + 8'h01;
  assign sel_965100 = array_index_964771 == array_index_948979 ? add_965099 : sel_965096;
  assign add_965103 = sel_965100 + 8'h01;
  assign sel_965104 = array_index_964771 == array_index_948985 ? add_965103 : sel_965100;
  assign add_965107 = sel_965104 + 8'h01;
  assign sel_965108 = array_index_964771 == array_index_948991 ? add_965107 : sel_965104;
  assign add_965111 = sel_965108 + 8'h01;
  assign sel_965112 = array_index_964771 == array_index_948997 ? add_965111 : sel_965108;
  assign add_965115 = sel_965112 + 8'h01;
  assign sel_965116 = array_index_964771 == array_index_949003 ? add_965115 : sel_965112;
  assign add_965119 = sel_965116 + 8'h01;
  assign sel_965120 = array_index_964771 == array_index_949009 ? add_965119 : sel_965116;
  assign add_965123 = sel_965120 + 8'h01;
  assign sel_965124 = array_index_964771 == array_index_949015 ? add_965123 : sel_965120;
  assign add_965127 = sel_965124 + 8'h01;
  assign sel_965128 = array_index_964771 == array_index_949021 ? add_965127 : sel_965124;
  assign add_965131 = sel_965128 + 8'h01;
  assign sel_965132 = array_index_964771 == array_index_949027 ? add_965131 : sel_965128;
  assign add_965135 = sel_965132 + 8'h01;
  assign sel_965136 = array_index_964771 == array_index_949033 ? add_965135 : sel_965132;
  assign add_965139 = sel_965136 + 8'h01;
  assign sel_965140 = array_index_964771 == array_index_949039 ? add_965139 : sel_965136;
  assign add_965143 = sel_965140 + 8'h01;
  assign sel_965144 = array_index_964771 == array_index_949045 ? add_965143 : sel_965140;
  assign add_965147 = sel_965144 + 8'h01;
  assign sel_965148 = array_index_964771 == array_index_949051 ? add_965147 : sel_965144;
  assign add_965151 = sel_965148 + 8'h01;
  assign sel_965152 = array_index_964771 == array_index_949057 ? add_965151 : sel_965148;
  assign add_965155 = sel_965152 + 8'h01;
  assign sel_965156 = array_index_964771 == array_index_949063 ? add_965155 : sel_965152;
  assign add_965159 = sel_965156 + 8'h01;
  assign sel_965160 = array_index_964771 == array_index_949069 ? add_965159 : sel_965156;
  assign add_965163 = sel_965160 + 8'h01;
  assign sel_965164 = array_index_964771 == array_index_949075 ? add_965163 : sel_965160;
  assign add_965167 = sel_965164 + 8'h01;
  assign sel_965168 = array_index_964771 == array_index_949081 ? add_965167 : sel_965164;
  assign add_965172 = sel_965168 + 8'h01;
  assign array_index_965173 = set1_unflattened[7'h29];
  assign sel_965174 = array_index_964771 == array_index_949087 ? add_965172 : sel_965168;
  assign add_965177 = sel_965174 + 8'h01;
  assign sel_965178 = array_index_965173 == array_index_948483 ? add_965177 : sel_965174;
  assign add_965181 = sel_965178 + 8'h01;
  assign sel_965182 = array_index_965173 == array_index_948487 ? add_965181 : sel_965178;
  assign add_965185 = sel_965182 + 8'h01;
  assign sel_965186 = array_index_965173 == array_index_948495 ? add_965185 : sel_965182;
  assign add_965189 = sel_965186 + 8'h01;
  assign sel_965190 = array_index_965173 == array_index_948503 ? add_965189 : sel_965186;
  assign add_965193 = sel_965190 + 8'h01;
  assign sel_965194 = array_index_965173 == array_index_948511 ? add_965193 : sel_965190;
  assign add_965197 = sel_965194 + 8'h01;
  assign sel_965198 = array_index_965173 == array_index_948519 ? add_965197 : sel_965194;
  assign add_965201 = sel_965198 + 8'h01;
  assign sel_965202 = array_index_965173 == array_index_948527 ? add_965201 : sel_965198;
  assign add_965205 = sel_965202 + 8'h01;
  assign sel_965206 = array_index_965173 == array_index_948535 ? add_965205 : sel_965202;
  assign add_965209 = sel_965206 + 8'h01;
  assign sel_965210 = array_index_965173 == array_index_948541 ? add_965209 : sel_965206;
  assign add_965213 = sel_965210 + 8'h01;
  assign sel_965214 = array_index_965173 == array_index_948547 ? add_965213 : sel_965210;
  assign add_965217 = sel_965214 + 8'h01;
  assign sel_965218 = array_index_965173 == array_index_948553 ? add_965217 : sel_965214;
  assign add_965221 = sel_965218 + 8'h01;
  assign sel_965222 = array_index_965173 == array_index_948559 ? add_965221 : sel_965218;
  assign add_965225 = sel_965222 + 8'h01;
  assign sel_965226 = array_index_965173 == array_index_948565 ? add_965225 : sel_965222;
  assign add_965229 = sel_965226 + 8'h01;
  assign sel_965230 = array_index_965173 == array_index_948571 ? add_965229 : sel_965226;
  assign add_965233 = sel_965230 + 8'h01;
  assign sel_965234 = array_index_965173 == array_index_948577 ? add_965233 : sel_965230;
  assign add_965237 = sel_965234 + 8'h01;
  assign sel_965238 = array_index_965173 == array_index_948583 ? add_965237 : sel_965234;
  assign add_965241 = sel_965238 + 8'h01;
  assign sel_965242 = array_index_965173 == array_index_948589 ? add_965241 : sel_965238;
  assign add_965245 = sel_965242 + 8'h01;
  assign sel_965246 = array_index_965173 == array_index_948595 ? add_965245 : sel_965242;
  assign add_965249 = sel_965246 + 8'h01;
  assign sel_965250 = array_index_965173 == array_index_948601 ? add_965249 : sel_965246;
  assign add_965253 = sel_965250 + 8'h01;
  assign sel_965254 = array_index_965173 == array_index_948607 ? add_965253 : sel_965250;
  assign add_965257 = sel_965254 + 8'h01;
  assign sel_965258 = array_index_965173 == array_index_948613 ? add_965257 : sel_965254;
  assign add_965261 = sel_965258 + 8'h01;
  assign sel_965262 = array_index_965173 == array_index_948619 ? add_965261 : sel_965258;
  assign add_965265 = sel_965262 + 8'h01;
  assign sel_965266 = array_index_965173 == array_index_948625 ? add_965265 : sel_965262;
  assign add_965269 = sel_965266 + 8'h01;
  assign sel_965270 = array_index_965173 == array_index_948631 ? add_965269 : sel_965266;
  assign add_965273 = sel_965270 + 8'h01;
  assign sel_965274 = array_index_965173 == array_index_948637 ? add_965273 : sel_965270;
  assign add_965277 = sel_965274 + 8'h01;
  assign sel_965278 = array_index_965173 == array_index_948643 ? add_965277 : sel_965274;
  assign add_965281 = sel_965278 + 8'h01;
  assign sel_965282 = array_index_965173 == array_index_948649 ? add_965281 : sel_965278;
  assign add_965285 = sel_965282 + 8'h01;
  assign sel_965286 = array_index_965173 == array_index_948655 ? add_965285 : sel_965282;
  assign add_965289 = sel_965286 + 8'h01;
  assign sel_965290 = array_index_965173 == array_index_948661 ? add_965289 : sel_965286;
  assign add_965293 = sel_965290 + 8'h01;
  assign sel_965294 = array_index_965173 == array_index_948667 ? add_965293 : sel_965290;
  assign add_965297 = sel_965294 + 8'h01;
  assign sel_965298 = array_index_965173 == array_index_948673 ? add_965297 : sel_965294;
  assign add_965301 = sel_965298 + 8'h01;
  assign sel_965302 = array_index_965173 == array_index_948679 ? add_965301 : sel_965298;
  assign add_965305 = sel_965302 + 8'h01;
  assign sel_965306 = array_index_965173 == array_index_948685 ? add_965305 : sel_965302;
  assign add_965309 = sel_965306 + 8'h01;
  assign sel_965310 = array_index_965173 == array_index_948691 ? add_965309 : sel_965306;
  assign add_965313 = sel_965310 + 8'h01;
  assign sel_965314 = array_index_965173 == array_index_948697 ? add_965313 : sel_965310;
  assign add_965317 = sel_965314 + 8'h01;
  assign sel_965318 = array_index_965173 == array_index_948703 ? add_965317 : sel_965314;
  assign add_965321 = sel_965318 + 8'h01;
  assign sel_965322 = array_index_965173 == array_index_948709 ? add_965321 : sel_965318;
  assign add_965325 = sel_965322 + 8'h01;
  assign sel_965326 = array_index_965173 == array_index_948715 ? add_965325 : sel_965322;
  assign add_965329 = sel_965326 + 8'h01;
  assign sel_965330 = array_index_965173 == array_index_948721 ? add_965329 : sel_965326;
  assign add_965333 = sel_965330 + 8'h01;
  assign sel_965334 = array_index_965173 == array_index_948727 ? add_965333 : sel_965330;
  assign add_965337 = sel_965334 + 8'h01;
  assign sel_965338 = array_index_965173 == array_index_948733 ? add_965337 : sel_965334;
  assign add_965341 = sel_965338 + 8'h01;
  assign sel_965342 = array_index_965173 == array_index_948739 ? add_965341 : sel_965338;
  assign add_965345 = sel_965342 + 8'h01;
  assign sel_965346 = array_index_965173 == array_index_948745 ? add_965345 : sel_965342;
  assign add_965349 = sel_965346 + 8'h01;
  assign sel_965350 = array_index_965173 == array_index_948751 ? add_965349 : sel_965346;
  assign add_965353 = sel_965350 + 8'h01;
  assign sel_965354 = array_index_965173 == array_index_948757 ? add_965353 : sel_965350;
  assign add_965357 = sel_965354 + 8'h01;
  assign sel_965358 = array_index_965173 == array_index_948763 ? add_965357 : sel_965354;
  assign add_965361 = sel_965358 + 8'h01;
  assign sel_965362 = array_index_965173 == array_index_948769 ? add_965361 : sel_965358;
  assign add_965365 = sel_965362 + 8'h01;
  assign sel_965366 = array_index_965173 == array_index_948775 ? add_965365 : sel_965362;
  assign add_965369 = sel_965366 + 8'h01;
  assign sel_965370 = array_index_965173 == array_index_948781 ? add_965369 : sel_965366;
  assign add_965373 = sel_965370 + 8'h01;
  assign sel_965374 = array_index_965173 == array_index_948787 ? add_965373 : sel_965370;
  assign add_965377 = sel_965374 + 8'h01;
  assign sel_965378 = array_index_965173 == array_index_948793 ? add_965377 : sel_965374;
  assign add_965381 = sel_965378 + 8'h01;
  assign sel_965382 = array_index_965173 == array_index_948799 ? add_965381 : sel_965378;
  assign add_965385 = sel_965382 + 8'h01;
  assign sel_965386 = array_index_965173 == array_index_948805 ? add_965385 : sel_965382;
  assign add_965389 = sel_965386 + 8'h01;
  assign sel_965390 = array_index_965173 == array_index_948811 ? add_965389 : sel_965386;
  assign add_965393 = sel_965390 + 8'h01;
  assign sel_965394 = array_index_965173 == array_index_948817 ? add_965393 : sel_965390;
  assign add_965397 = sel_965394 + 8'h01;
  assign sel_965398 = array_index_965173 == array_index_948823 ? add_965397 : sel_965394;
  assign add_965401 = sel_965398 + 8'h01;
  assign sel_965402 = array_index_965173 == array_index_948829 ? add_965401 : sel_965398;
  assign add_965405 = sel_965402 + 8'h01;
  assign sel_965406 = array_index_965173 == array_index_948835 ? add_965405 : sel_965402;
  assign add_965409 = sel_965406 + 8'h01;
  assign sel_965410 = array_index_965173 == array_index_948841 ? add_965409 : sel_965406;
  assign add_965413 = sel_965410 + 8'h01;
  assign sel_965414 = array_index_965173 == array_index_948847 ? add_965413 : sel_965410;
  assign add_965417 = sel_965414 + 8'h01;
  assign sel_965418 = array_index_965173 == array_index_948853 ? add_965417 : sel_965414;
  assign add_965421 = sel_965418 + 8'h01;
  assign sel_965422 = array_index_965173 == array_index_948859 ? add_965421 : sel_965418;
  assign add_965425 = sel_965422 + 8'h01;
  assign sel_965426 = array_index_965173 == array_index_948865 ? add_965425 : sel_965422;
  assign add_965429 = sel_965426 + 8'h01;
  assign sel_965430 = array_index_965173 == array_index_948871 ? add_965429 : sel_965426;
  assign add_965433 = sel_965430 + 8'h01;
  assign sel_965434 = array_index_965173 == array_index_948877 ? add_965433 : sel_965430;
  assign add_965437 = sel_965434 + 8'h01;
  assign sel_965438 = array_index_965173 == array_index_948883 ? add_965437 : sel_965434;
  assign add_965441 = sel_965438 + 8'h01;
  assign sel_965442 = array_index_965173 == array_index_948889 ? add_965441 : sel_965438;
  assign add_965445 = sel_965442 + 8'h01;
  assign sel_965446 = array_index_965173 == array_index_948895 ? add_965445 : sel_965442;
  assign add_965449 = sel_965446 + 8'h01;
  assign sel_965450 = array_index_965173 == array_index_948901 ? add_965449 : sel_965446;
  assign add_965453 = sel_965450 + 8'h01;
  assign sel_965454 = array_index_965173 == array_index_948907 ? add_965453 : sel_965450;
  assign add_965457 = sel_965454 + 8'h01;
  assign sel_965458 = array_index_965173 == array_index_948913 ? add_965457 : sel_965454;
  assign add_965461 = sel_965458 + 8'h01;
  assign sel_965462 = array_index_965173 == array_index_948919 ? add_965461 : sel_965458;
  assign add_965465 = sel_965462 + 8'h01;
  assign sel_965466 = array_index_965173 == array_index_948925 ? add_965465 : sel_965462;
  assign add_965469 = sel_965466 + 8'h01;
  assign sel_965470 = array_index_965173 == array_index_948931 ? add_965469 : sel_965466;
  assign add_965473 = sel_965470 + 8'h01;
  assign sel_965474 = array_index_965173 == array_index_948937 ? add_965473 : sel_965470;
  assign add_965477 = sel_965474 + 8'h01;
  assign sel_965478 = array_index_965173 == array_index_948943 ? add_965477 : sel_965474;
  assign add_965481 = sel_965478 + 8'h01;
  assign sel_965482 = array_index_965173 == array_index_948949 ? add_965481 : sel_965478;
  assign add_965485 = sel_965482 + 8'h01;
  assign sel_965486 = array_index_965173 == array_index_948955 ? add_965485 : sel_965482;
  assign add_965489 = sel_965486 + 8'h01;
  assign sel_965490 = array_index_965173 == array_index_948961 ? add_965489 : sel_965486;
  assign add_965493 = sel_965490 + 8'h01;
  assign sel_965494 = array_index_965173 == array_index_948967 ? add_965493 : sel_965490;
  assign add_965497 = sel_965494 + 8'h01;
  assign sel_965498 = array_index_965173 == array_index_948973 ? add_965497 : sel_965494;
  assign add_965501 = sel_965498 + 8'h01;
  assign sel_965502 = array_index_965173 == array_index_948979 ? add_965501 : sel_965498;
  assign add_965505 = sel_965502 + 8'h01;
  assign sel_965506 = array_index_965173 == array_index_948985 ? add_965505 : sel_965502;
  assign add_965509 = sel_965506 + 8'h01;
  assign sel_965510 = array_index_965173 == array_index_948991 ? add_965509 : sel_965506;
  assign add_965513 = sel_965510 + 8'h01;
  assign sel_965514 = array_index_965173 == array_index_948997 ? add_965513 : sel_965510;
  assign add_965517 = sel_965514 + 8'h01;
  assign sel_965518 = array_index_965173 == array_index_949003 ? add_965517 : sel_965514;
  assign add_965521 = sel_965518 + 8'h01;
  assign sel_965522 = array_index_965173 == array_index_949009 ? add_965521 : sel_965518;
  assign add_965525 = sel_965522 + 8'h01;
  assign sel_965526 = array_index_965173 == array_index_949015 ? add_965525 : sel_965522;
  assign add_965529 = sel_965526 + 8'h01;
  assign sel_965530 = array_index_965173 == array_index_949021 ? add_965529 : sel_965526;
  assign add_965533 = sel_965530 + 8'h01;
  assign sel_965534 = array_index_965173 == array_index_949027 ? add_965533 : sel_965530;
  assign add_965537 = sel_965534 + 8'h01;
  assign sel_965538 = array_index_965173 == array_index_949033 ? add_965537 : sel_965534;
  assign add_965541 = sel_965538 + 8'h01;
  assign sel_965542 = array_index_965173 == array_index_949039 ? add_965541 : sel_965538;
  assign add_965545 = sel_965542 + 8'h01;
  assign sel_965546 = array_index_965173 == array_index_949045 ? add_965545 : sel_965542;
  assign add_965549 = sel_965546 + 8'h01;
  assign sel_965550 = array_index_965173 == array_index_949051 ? add_965549 : sel_965546;
  assign add_965553 = sel_965550 + 8'h01;
  assign sel_965554 = array_index_965173 == array_index_949057 ? add_965553 : sel_965550;
  assign add_965557 = sel_965554 + 8'h01;
  assign sel_965558 = array_index_965173 == array_index_949063 ? add_965557 : sel_965554;
  assign add_965561 = sel_965558 + 8'h01;
  assign sel_965562 = array_index_965173 == array_index_949069 ? add_965561 : sel_965558;
  assign add_965565 = sel_965562 + 8'h01;
  assign sel_965566 = array_index_965173 == array_index_949075 ? add_965565 : sel_965562;
  assign add_965569 = sel_965566 + 8'h01;
  assign sel_965570 = array_index_965173 == array_index_949081 ? add_965569 : sel_965566;
  assign add_965574 = sel_965570 + 8'h01;
  assign array_index_965575 = set1_unflattened[7'h2a];
  assign sel_965576 = array_index_965173 == array_index_949087 ? add_965574 : sel_965570;
  assign add_965579 = sel_965576 + 8'h01;
  assign sel_965580 = array_index_965575 == array_index_948483 ? add_965579 : sel_965576;
  assign add_965583 = sel_965580 + 8'h01;
  assign sel_965584 = array_index_965575 == array_index_948487 ? add_965583 : sel_965580;
  assign add_965587 = sel_965584 + 8'h01;
  assign sel_965588 = array_index_965575 == array_index_948495 ? add_965587 : sel_965584;
  assign add_965591 = sel_965588 + 8'h01;
  assign sel_965592 = array_index_965575 == array_index_948503 ? add_965591 : sel_965588;
  assign add_965595 = sel_965592 + 8'h01;
  assign sel_965596 = array_index_965575 == array_index_948511 ? add_965595 : sel_965592;
  assign add_965599 = sel_965596 + 8'h01;
  assign sel_965600 = array_index_965575 == array_index_948519 ? add_965599 : sel_965596;
  assign add_965603 = sel_965600 + 8'h01;
  assign sel_965604 = array_index_965575 == array_index_948527 ? add_965603 : sel_965600;
  assign add_965607 = sel_965604 + 8'h01;
  assign sel_965608 = array_index_965575 == array_index_948535 ? add_965607 : sel_965604;
  assign add_965611 = sel_965608 + 8'h01;
  assign sel_965612 = array_index_965575 == array_index_948541 ? add_965611 : sel_965608;
  assign add_965615 = sel_965612 + 8'h01;
  assign sel_965616 = array_index_965575 == array_index_948547 ? add_965615 : sel_965612;
  assign add_965619 = sel_965616 + 8'h01;
  assign sel_965620 = array_index_965575 == array_index_948553 ? add_965619 : sel_965616;
  assign add_965623 = sel_965620 + 8'h01;
  assign sel_965624 = array_index_965575 == array_index_948559 ? add_965623 : sel_965620;
  assign add_965627 = sel_965624 + 8'h01;
  assign sel_965628 = array_index_965575 == array_index_948565 ? add_965627 : sel_965624;
  assign add_965631 = sel_965628 + 8'h01;
  assign sel_965632 = array_index_965575 == array_index_948571 ? add_965631 : sel_965628;
  assign add_965635 = sel_965632 + 8'h01;
  assign sel_965636 = array_index_965575 == array_index_948577 ? add_965635 : sel_965632;
  assign add_965639 = sel_965636 + 8'h01;
  assign sel_965640 = array_index_965575 == array_index_948583 ? add_965639 : sel_965636;
  assign add_965643 = sel_965640 + 8'h01;
  assign sel_965644 = array_index_965575 == array_index_948589 ? add_965643 : sel_965640;
  assign add_965647 = sel_965644 + 8'h01;
  assign sel_965648 = array_index_965575 == array_index_948595 ? add_965647 : sel_965644;
  assign add_965651 = sel_965648 + 8'h01;
  assign sel_965652 = array_index_965575 == array_index_948601 ? add_965651 : sel_965648;
  assign add_965655 = sel_965652 + 8'h01;
  assign sel_965656 = array_index_965575 == array_index_948607 ? add_965655 : sel_965652;
  assign add_965659 = sel_965656 + 8'h01;
  assign sel_965660 = array_index_965575 == array_index_948613 ? add_965659 : sel_965656;
  assign add_965663 = sel_965660 + 8'h01;
  assign sel_965664 = array_index_965575 == array_index_948619 ? add_965663 : sel_965660;
  assign add_965667 = sel_965664 + 8'h01;
  assign sel_965668 = array_index_965575 == array_index_948625 ? add_965667 : sel_965664;
  assign add_965671 = sel_965668 + 8'h01;
  assign sel_965672 = array_index_965575 == array_index_948631 ? add_965671 : sel_965668;
  assign add_965675 = sel_965672 + 8'h01;
  assign sel_965676 = array_index_965575 == array_index_948637 ? add_965675 : sel_965672;
  assign add_965679 = sel_965676 + 8'h01;
  assign sel_965680 = array_index_965575 == array_index_948643 ? add_965679 : sel_965676;
  assign add_965683 = sel_965680 + 8'h01;
  assign sel_965684 = array_index_965575 == array_index_948649 ? add_965683 : sel_965680;
  assign add_965687 = sel_965684 + 8'h01;
  assign sel_965688 = array_index_965575 == array_index_948655 ? add_965687 : sel_965684;
  assign add_965691 = sel_965688 + 8'h01;
  assign sel_965692 = array_index_965575 == array_index_948661 ? add_965691 : sel_965688;
  assign add_965695 = sel_965692 + 8'h01;
  assign sel_965696 = array_index_965575 == array_index_948667 ? add_965695 : sel_965692;
  assign add_965699 = sel_965696 + 8'h01;
  assign sel_965700 = array_index_965575 == array_index_948673 ? add_965699 : sel_965696;
  assign add_965703 = sel_965700 + 8'h01;
  assign sel_965704 = array_index_965575 == array_index_948679 ? add_965703 : sel_965700;
  assign add_965707 = sel_965704 + 8'h01;
  assign sel_965708 = array_index_965575 == array_index_948685 ? add_965707 : sel_965704;
  assign add_965711 = sel_965708 + 8'h01;
  assign sel_965712 = array_index_965575 == array_index_948691 ? add_965711 : sel_965708;
  assign add_965715 = sel_965712 + 8'h01;
  assign sel_965716 = array_index_965575 == array_index_948697 ? add_965715 : sel_965712;
  assign add_965719 = sel_965716 + 8'h01;
  assign sel_965720 = array_index_965575 == array_index_948703 ? add_965719 : sel_965716;
  assign add_965723 = sel_965720 + 8'h01;
  assign sel_965724 = array_index_965575 == array_index_948709 ? add_965723 : sel_965720;
  assign add_965727 = sel_965724 + 8'h01;
  assign sel_965728 = array_index_965575 == array_index_948715 ? add_965727 : sel_965724;
  assign add_965731 = sel_965728 + 8'h01;
  assign sel_965732 = array_index_965575 == array_index_948721 ? add_965731 : sel_965728;
  assign add_965735 = sel_965732 + 8'h01;
  assign sel_965736 = array_index_965575 == array_index_948727 ? add_965735 : sel_965732;
  assign add_965739 = sel_965736 + 8'h01;
  assign sel_965740 = array_index_965575 == array_index_948733 ? add_965739 : sel_965736;
  assign add_965743 = sel_965740 + 8'h01;
  assign sel_965744 = array_index_965575 == array_index_948739 ? add_965743 : sel_965740;
  assign add_965747 = sel_965744 + 8'h01;
  assign sel_965748 = array_index_965575 == array_index_948745 ? add_965747 : sel_965744;
  assign add_965751 = sel_965748 + 8'h01;
  assign sel_965752 = array_index_965575 == array_index_948751 ? add_965751 : sel_965748;
  assign add_965755 = sel_965752 + 8'h01;
  assign sel_965756 = array_index_965575 == array_index_948757 ? add_965755 : sel_965752;
  assign add_965759 = sel_965756 + 8'h01;
  assign sel_965760 = array_index_965575 == array_index_948763 ? add_965759 : sel_965756;
  assign add_965763 = sel_965760 + 8'h01;
  assign sel_965764 = array_index_965575 == array_index_948769 ? add_965763 : sel_965760;
  assign add_965767 = sel_965764 + 8'h01;
  assign sel_965768 = array_index_965575 == array_index_948775 ? add_965767 : sel_965764;
  assign add_965771 = sel_965768 + 8'h01;
  assign sel_965772 = array_index_965575 == array_index_948781 ? add_965771 : sel_965768;
  assign add_965775 = sel_965772 + 8'h01;
  assign sel_965776 = array_index_965575 == array_index_948787 ? add_965775 : sel_965772;
  assign add_965779 = sel_965776 + 8'h01;
  assign sel_965780 = array_index_965575 == array_index_948793 ? add_965779 : sel_965776;
  assign add_965783 = sel_965780 + 8'h01;
  assign sel_965784 = array_index_965575 == array_index_948799 ? add_965783 : sel_965780;
  assign add_965787 = sel_965784 + 8'h01;
  assign sel_965788 = array_index_965575 == array_index_948805 ? add_965787 : sel_965784;
  assign add_965791 = sel_965788 + 8'h01;
  assign sel_965792 = array_index_965575 == array_index_948811 ? add_965791 : sel_965788;
  assign add_965795 = sel_965792 + 8'h01;
  assign sel_965796 = array_index_965575 == array_index_948817 ? add_965795 : sel_965792;
  assign add_965799 = sel_965796 + 8'h01;
  assign sel_965800 = array_index_965575 == array_index_948823 ? add_965799 : sel_965796;
  assign add_965803 = sel_965800 + 8'h01;
  assign sel_965804 = array_index_965575 == array_index_948829 ? add_965803 : sel_965800;
  assign add_965807 = sel_965804 + 8'h01;
  assign sel_965808 = array_index_965575 == array_index_948835 ? add_965807 : sel_965804;
  assign add_965811 = sel_965808 + 8'h01;
  assign sel_965812 = array_index_965575 == array_index_948841 ? add_965811 : sel_965808;
  assign add_965815 = sel_965812 + 8'h01;
  assign sel_965816 = array_index_965575 == array_index_948847 ? add_965815 : sel_965812;
  assign add_965819 = sel_965816 + 8'h01;
  assign sel_965820 = array_index_965575 == array_index_948853 ? add_965819 : sel_965816;
  assign add_965823 = sel_965820 + 8'h01;
  assign sel_965824 = array_index_965575 == array_index_948859 ? add_965823 : sel_965820;
  assign add_965827 = sel_965824 + 8'h01;
  assign sel_965828 = array_index_965575 == array_index_948865 ? add_965827 : sel_965824;
  assign add_965831 = sel_965828 + 8'h01;
  assign sel_965832 = array_index_965575 == array_index_948871 ? add_965831 : sel_965828;
  assign add_965835 = sel_965832 + 8'h01;
  assign sel_965836 = array_index_965575 == array_index_948877 ? add_965835 : sel_965832;
  assign add_965839 = sel_965836 + 8'h01;
  assign sel_965840 = array_index_965575 == array_index_948883 ? add_965839 : sel_965836;
  assign add_965843 = sel_965840 + 8'h01;
  assign sel_965844 = array_index_965575 == array_index_948889 ? add_965843 : sel_965840;
  assign add_965847 = sel_965844 + 8'h01;
  assign sel_965848 = array_index_965575 == array_index_948895 ? add_965847 : sel_965844;
  assign add_965851 = sel_965848 + 8'h01;
  assign sel_965852 = array_index_965575 == array_index_948901 ? add_965851 : sel_965848;
  assign add_965855 = sel_965852 + 8'h01;
  assign sel_965856 = array_index_965575 == array_index_948907 ? add_965855 : sel_965852;
  assign add_965859 = sel_965856 + 8'h01;
  assign sel_965860 = array_index_965575 == array_index_948913 ? add_965859 : sel_965856;
  assign add_965863 = sel_965860 + 8'h01;
  assign sel_965864 = array_index_965575 == array_index_948919 ? add_965863 : sel_965860;
  assign add_965867 = sel_965864 + 8'h01;
  assign sel_965868 = array_index_965575 == array_index_948925 ? add_965867 : sel_965864;
  assign add_965871 = sel_965868 + 8'h01;
  assign sel_965872 = array_index_965575 == array_index_948931 ? add_965871 : sel_965868;
  assign add_965875 = sel_965872 + 8'h01;
  assign sel_965876 = array_index_965575 == array_index_948937 ? add_965875 : sel_965872;
  assign add_965879 = sel_965876 + 8'h01;
  assign sel_965880 = array_index_965575 == array_index_948943 ? add_965879 : sel_965876;
  assign add_965883 = sel_965880 + 8'h01;
  assign sel_965884 = array_index_965575 == array_index_948949 ? add_965883 : sel_965880;
  assign add_965887 = sel_965884 + 8'h01;
  assign sel_965888 = array_index_965575 == array_index_948955 ? add_965887 : sel_965884;
  assign add_965891 = sel_965888 + 8'h01;
  assign sel_965892 = array_index_965575 == array_index_948961 ? add_965891 : sel_965888;
  assign add_965895 = sel_965892 + 8'h01;
  assign sel_965896 = array_index_965575 == array_index_948967 ? add_965895 : sel_965892;
  assign add_965899 = sel_965896 + 8'h01;
  assign sel_965900 = array_index_965575 == array_index_948973 ? add_965899 : sel_965896;
  assign add_965903 = sel_965900 + 8'h01;
  assign sel_965904 = array_index_965575 == array_index_948979 ? add_965903 : sel_965900;
  assign add_965907 = sel_965904 + 8'h01;
  assign sel_965908 = array_index_965575 == array_index_948985 ? add_965907 : sel_965904;
  assign add_965911 = sel_965908 + 8'h01;
  assign sel_965912 = array_index_965575 == array_index_948991 ? add_965911 : sel_965908;
  assign add_965915 = sel_965912 + 8'h01;
  assign sel_965916 = array_index_965575 == array_index_948997 ? add_965915 : sel_965912;
  assign add_965919 = sel_965916 + 8'h01;
  assign sel_965920 = array_index_965575 == array_index_949003 ? add_965919 : sel_965916;
  assign add_965923 = sel_965920 + 8'h01;
  assign sel_965924 = array_index_965575 == array_index_949009 ? add_965923 : sel_965920;
  assign add_965927 = sel_965924 + 8'h01;
  assign sel_965928 = array_index_965575 == array_index_949015 ? add_965927 : sel_965924;
  assign add_965931 = sel_965928 + 8'h01;
  assign sel_965932 = array_index_965575 == array_index_949021 ? add_965931 : sel_965928;
  assign add_965935 = sel_965932 + 8'h01;
  assign sel_965936 = array_index_965575 == array_index_949027 ? add_965935 : sel_965932;
  assign add_965939 = sel_965936 + 8'h01;
  assign sel_965940 = array_index_965575 == array_index_949033 ? add_965939 : sel_965936;
  assign add_965943 = sel_965940 + 8'h01;
  assign sel_965944 = array_index_965575 == array_index_949039 ? add_965943 : sel_965940;
  assign add_965947 = sel_965944 + 8'h01;
  assign sel_965948 = array_index_965575 == array_index_949045 ? add_965947 : sel_965944;
  assign add_965951 = sel_965948 + 8'h01;
  assign sel_965952 = array_index_965575 == array_index_949051 ? add_965951 : sel_965948;
  assign add_965955 = sel_965952 + 8'h01;
  assign sel_965956 = array_index_965575 == array_index_949057 ? add_965955 : sel_965952;
  assign add_965959 = sel_965956 + 8'h01;
  assign sel_965960 = array_index_965575 == array_index_949063 ? add_965959 : sel_965956;
  assign add_965963 = sel_965960 + 8'h01;
  assign sel_965964 = array_index_965575 == array_index_949069 ? add_965963 : sel_965960;
  assign add_965967 = sel_965964 + 8'h01;
  assign sel_965968 = array_index_965575 == array_index_949075 ? add_965967 : sel_965964;
  assign add_965971 = sel_965968 + 8'h01;
  assign sel_965972 = array_index_965575 == array_index_949081 ? add_965971 : sel_965968;
  assign add_965976 = sel_965972 + 8'h01;
  assign array_index_965977 = set1_unflattened[7'h2b];
  assign sel_965978 = array_index_965575 == array_index_949087 ? add_965976 : sel_965972;
  assign add_965981 = sel_965978 + 8'h01;
  assign sel_965982 = array_index_965977 == array_index_948483 ? add_965981 : sel_965978;
  assign add_965985 = sel_965982 + 8'h01;
  assign sel_965986 = array_index_965977 == array_index_948487 ? add_965985 : sel_965982;
  assign add_965989 = sel_965986 + 8'h01;
  assign sel_965990 = array_index_965977 == array_index_948495 ? add_965989 : sel_965986;
  assign add_965993 = sel_965990 + 8'h01;
  assign sel_965994 = array_index_965977 == array_index_948503 ? add_965993 : sel_965990;
  assign add_965997 = sel_965994 + 8'h01;
  assign sel_965998 = array_index_965977 == array_index_948511 ? add_965997 : sel_965994;
  assign add_966001 = sel_965998 + 8'h01;
  assign sel_966002 = array_index_965977 == array_index_948519 ? add_966001 : sel_965998;
  assign add_966005 = sel_966002 + 8'h01;
  assign sel_966006 = array_index_965977 == array_index_948527 ? add_966005 : sel_966002;
  assign add_966009 = sel_966006 + 8'h01;
  assign sel_966010 = array_index_965977 == array_index_948535 ? add_966009 : sel_966006;
  assign add_966013 = sel_966010 + 8'h01;
  assign sel_966014 = array_index_965977 == array_index_948541 ? add_966013 : sel_966010;
  assign add_966017 = sel_966014 + 8'h01;
  assign sel_966018 = array_index_965977 == array_index_948547 ? add_966017 : sel_966014;
  assign add_966021 = sel_966018 + 8'h01;
  assign sel_966022 = array_index_965977 == array_index_948553 ? add_966021 : sel_966018;
  assign add_966025 = sel_966022 + 8'h01;
  assign sel_966026 = array_index_965977 == array_index_948559 ? add_966025 : sel_966022;
  assign add_966029 = sel_966026 + 8'h01;
  assign sel_966030 = array_index_965977 == array_index_948565 ? add_966029 : sel_966026;
  assign add_966033 = sel_966030 + 8'h01;
  assign sel_966034 = array_index_965977 == array_index_948571 ? add_966033 : sel_966030;
  assign add_966037 = sel_966034 + 8'h01;
  assign sel_966038 = array_index_965977 == array_index_948577 ? add_966037 : sel_966034;
  assign add_966041 = sel_966038 + 8'h01;
  assign sel_966042 = array_index_965977 == array_index_948583 ? add_966041 : sel_966038;
  assign add_966045 = sel_966042 + 8'h01;
  assign sel_966046 = array_index_965977 == array_index_948589 ? add_966045 : sel_966042;
  assign add_966049 = sel_966046 + 8'h01;
  assign sel_966050 = array_index_965977 == array_index_948595 ? add_966049 : sel_966046;
  assign add_966053 = sel_966050 + 8'h01;
  assign sel_966054 = array_index_965977 == array_index_948601 ? add_966053 : sel_966050;
  assign add_966057 = sel_966054 + 8'h01;
  assign sel_966058 = array_index_965977 == array_index_948607 ? add_966057 : sel_966054;
  assign add_966061 = sel_966058 + 8'h01;
  assign sel_966062 = array_index_965977 == array_index_948613 ? add_966061 : sel_966058;
  assign add_966065 = sel_966062 + 8'h01;
  assign sel_966066 = array_index_965977 == array_index_948619 ? add_966065 : sel_966062;
  assign add_966069 = sel_966066 + 8'h01;
  assign sel_966070 = array_index_965977 == array_index_948625 ? add_966069 : sel_966066;
  assign add_966073 = sel_966070 + 8'h01;
  assign sel_966074 = array_index_965977 == array_index_948631 ? add_966073 : sel_966070;
  assign add_966077 = sel_966074 + 8'h01;
  assign sel_966078 = array_index_965977 == array_index_948637 ? add_966077 : sel_966074;
  assign add_966081 = sel_966078 + 8'h01;
  assign sel_966082 = array_index_965977 == array_index_948643 ? add_966081 : sel_966078;
  assign add_966085 = sel_966082 + 8'h01;
  assign sel_966086 = array_index_965977 == array_index_948649 ? add_966085 : sel_966082;
  assign add_966089 = sel_966086 + 8'h01;
  assign sel_966090 = array_index_965977 == array_index_948655 ? add_966089 : sel_966086;
  assign add_966093 = sel_966090 + 8'h01;
  assign sel_966094 = array_index_965977 == array_index_948661 ? add_966093 : sel_966090;
  assign add_966097 = sel_966094 + 8'h01;
  assign sel_966098 = array_index_965977 == array_index_948667 ? add_966097 : sel_966094;
  assign add_966101 = sel_966098 + 8'h01;
  assign sel_966102 = array_index_965977 == array_index_948673 ? add_966101 : sel_966098;
  assign add_966105 = sel_966102 + 8'h01;
  assign sel_966106 = array_index_965977 == array_index_948679 ? add_966105 : sel_966102;
  assign add_966109 = sel_966106 + 8'h01;
  assign sel_966110 = array_index_965977 == array_index_948685 ? add_966109 : sel_966106;
  assign add_966113 = sel_966110 + 8'h01;
  assign sel_966114 = array_index_965977 == array_index_948691 ? add_966113 : sel_966110;
  assign add_966117 = sel_966114 + 8'h01;
  assign sel_966118 = array_index_965977 == array_index_948697 ? add_966117 : sel_966114;
  assign add_966121 = sel_966118 + 8'h01;
  assign sel_966122 = array_index_965977 == array_index_948703 ? add_966121 : sel_966118;
  assign add_966125 = sel_966122 + 8'h01;
  assign sel_966126 = array_index_965977 == array_index_948709 ? add_966125 : sel_966122;
  assign add_966129 = sel_966126 + 8'h01;
  assign sel_966130 = array_index_965977 == array_index_948715 ? add_966129 : sel_966126;
  assign add_966133 = sel_966130 + 8'h01;
  assign sel_966134 = array_index_965977 == array_index_948721 ? add_966133 : sel_966130;
  assign add_966137 = sel_966134 + 8'h01;
  assign sel_966138 = array_index_965977 == array_index_948727 ? add_966137 : sel_966134;
  assign add_966141 = sel_966138 + 8'h01;
  assign sel_966142 = array_index_965977 == array_index_948733 ? add_966141 : sel_966138;
  assign add_966145 = sel_966142 + 8'h01;
  assign sel_966146 = array_index_965977 == array_index_948739 ? add_966145 : sel_966142;
  assign add_966149 = sel_966146 + 8'h01;
  assign sel_966150 = array_index_965977 == array_index_948745 ? add_966149 : sel_966146;
  assign add_966153 = sel_966150 + 8'h01;
  assign sel_966154 = array_index_965977 == array_index_948751 ? add_966153 : sel_966150;
  assign add_966157 = sel_966154 + 8'h01;
  assign sel_966158 = array_index_965977 == array_index_948757 ? add_966157 : sel_966154;
  assign add_966161 = sel_966158 + 8'h01;
  assign sel_966162 = array_index_965977 == array_index_948763 ? add_966161 : sel_966158;
  assign add_966165 = sel_966162 + 8'h01;
  assign sel_966166 = array_index_965977 == array_index_948769 ? add_966165 : sel_966162;
  assign add_966169 = sel_966166 + 8'h01;
  assign sel_966170 = array_index_965977 == array_index_948775 ? add_966169 : sel_966166;
  assign add_966173 = sel_966170 + 8'h01;
  assign sel_966174 = array_index_965977 == array_index_948781 ? add_966173 : sel_966170;
  assign add_966177 = sel_966174 + 8'h01;
  assign sel_966178 = array_index_965977 == array_index_948787 ? add_966177 : sel_966174;
  assign add_966181 = sel_966178 + 8'h01;
  assign sel_966182 = array_index_965977 == array_index_948793 ? add_966181 : sel_966178;
  assign add_966185 = sel_966182 + 8'h01;
  assign sel_966186 = array_index_965977 == array_index_948799 ? add_966185 : sel_966182;
  assign add_966189 = sel_966186 + 8'h01;
  assign sel_966190 = array_index_965977 == array_index_948805 ? add_966189 : sel_966186;
  assign add_966193 = sel_966190 + 8'h01;
  assign sel_966194 = array_index_965977 == array_index_948811 ? add_966193 : sel_966190;
  assign add_966197 = sel_966194 + 8'h01;
  assign sel_966198 = array_index_965977 == array_index_948817 ? add_966197 : sel_966194;
  assign add_966201 = sel_966198 + 8'h01;
  assign sel_966202 = array_index_965977 == array_index_948823 ? add_966201 : sel_966198;
  assign add_966205 = sel_966202 + 8'h01;
  assign sel_966206 = array_index_965977 == array_index_948829 ? add_966205 : sel_966202;
  assign add_966209 = sel_966206 + 8'h01;
  assign sel_966210 = array_index_965977 == array_index_948835 ? add_966209 : sel_966206;
  assign add_966213 = sel_966210 + 8'h01;
  assign sel_966214 = array_index_965977 == array_index_948841 ? add_966213 : sel_966210;
  assign add_966217 = sel_966214 + 8'h01;
  assign sel_966218 = array_index_965977 == array_index_948847 ? add_966217 : sel_966214;
  assign add_966221 = sel_966218 + 8'h01;
  assign sel_966222 = array_index_965977 == array_index_948853 ? add_966221 : sel_966218;
  assign add_966225 = sel_966222 + 8'h01;
  assign sel_966226 = array_index_965977 == array_index_948859 ? add_966225 : sel_966222;
  assign add_966229 = sel_966226 + 8'h01;
  assign sel_966230 = array_index_965977 == array_index_948865 ? add_966229 : sel_966226;
  assign add_966233 = sel_966230 + 8'h01;
  assign sel_966234 = array_index_965977 == array_index_948871 ? add_966233 : sel_966230;
  assign add_966237 = sel_966234 + 8'h01;
  assign sel_966238 = array_index_965977 == array_index_948877 ? add_966237 : sel_966234;
  assign add_966241 = sel_966238 + 8'h01;
  assign sel_966242 = array_index_965977 == array_index_948883 ? add_966241 : sel_966238;
  assign add_966245 = sel_966242 + 8'h01;
  assign sel_966246 = array_index_965977 == array_index_948889 ? add_966245 : sel_966242;
  assign add_966249 = sel_966246 + 8'h01;
  assign sel_966250 = array_index_965977 == array_index_948895 ? add_966249 : sel_966246;
  assign add_966253 = sel_966250 + 8'h01;
  assign sel_966254 = array_index_965977 == array_index_948901 ? add_966253 : sel_966250;
  assign add_966257 = sel_966254 + 8'h01;
  assign sel_966258 = array_index_965977 == array_index_948907 ? add_966257 : sel_966254;
  assign add_966261 = sel_966258 + 8'h01;
  assign sel_966262 = array_index_965977 == array_index_948913 ? add_966261 : sel_966258;
  assign add_966265 = sel_966262 + 8'h01;
  assign sel_966266 = array_index_965977 == array_index_948919 ? add_966265 : sel_966262;
  assign add_966269 = sel_966266 + 8'h01;
  assign sel_966270 = array_index_965977 == array_index_948925 ? add_966269 : sel_966266;
  assign add_966273 = sel_966270 + 8'h01;
  assign sel_966274 = array_index_965977 == array_index_948931 ? add_966273 : sel_966270;
  assign add_966277 = sel_966274 + 8'h01;
  assign sel_966278 = array_index_965977 == array_index_948937 ? add_966277 : sel_966274;
  assign add_966281 = sel_966278 + 8'h01;
  assign sel_966282 = array_index_965977 == array_index_948943 ? add_966281 : sel_966278;
  assign add_966285 = sel_966282 + 8'h01;
  assign sel_966286 = array_index_965977 == array_index_948949 ? add_966285 : sel_966282;
  assign add_966289 = sel_966286 + 8'h01;
  assign sel_966290 = array_index_965977 == array_index_948955 ? add_966289 : sel_966286;
  assign add_966293 = sel_966290 + 8'h01;
  assign sel_966294 = array_index_965977 == array_index_948961 ? add_966293 : sel_966290;
  assign add_966297 = sel_966294 + 8'h01;
  assign sel_966298 = array_index_965977 == array_index_948967 ? add_966297 : sel_966294;
  assign add_966301 = sel_966298 + 8'h01;
  assign sel_966302 = array_index_965977 == array_index_948973 ? add_966301 : sel_966298;
  assign add_966305 = sel_966302 + 8'h01;
  assign sel_966306 = array_index_965977 == array_index_948979 ? add_966305 : sel_966302;
  assign add_966309 = sel_966306 + 8'h01;
  assign sel_966310 = array_index_965977 == array_index_948985 ? add_966309 : sel_966306;
  assign add_966313 = sel_966310 + 8'h01;
  assign sel_966314 = array_index_965977 == array_index_948991 ? add_966313 : sel_966310;
  assign add_966317 = sel_966314 + 8'h01;
  assign sel_966318 = array_index_965977 == array_index_948997 ? add_966317 : sel_966314;
  assign add_966321 = sel_966318 + 8'h01;
  assign sel_966322 = array_index_965977 == array_index_949003 ? add_966321 : sel_966318;
  assign add_966325 = sel_966322 + 8'h01;
  assign sel_966326 = array_index_965977 == array_index_949009 ? add_966325 : sel_966322;
  assign add_966329 = sel_966326 + 8'h01;
  assign sel_966330 = array_index_965977 == array_index_949015 ? add_966329 : sel_966326;
  assign add_966333 = sel_966330 + 8'h01;
  assign sel_966334 = array_index_965977 == array_index_949021 ? add_966333 : sel_966330;
  assign add_966337 = sel_966334 + 8'h01;
  assign sel_966338 = array_index_965977 == array_index_949027 ? add_966337 : sel_966334;
  assign add_966341 = sel_966338 + 8'h01;
  assign sel_966342 = array_index_965977 == array_index_949033 ? add_966341 : sel_966338;
  assign add_966345 = sel_966342 + 8'h01;
  assign sel_966346 = array_index_965977 == array_index_949039 ? add_966345 : sel_966342;
  assign add_966349 = sel_966346 + 8'h01;
  assign sel_966350 = array_index_965977 == array_index_949045 ? add_966349 : sel_966346;
  assign add_966353 = sel_966350 + 8'h01;
  assign sel_966354 = array_index_965977 == array_index_949051 ? add_966353 : sel_966350;
  assign add_966357 = sel_966354 + 8'h01;
  assign sel_966358 = array_index_965977 == array_index_949057 ? add_966357 : sel_966354;
  assign add_966361 = sel_966358 + 8'h01;
  assign sel_966362 = array_index_965977 == array_index_949063 ? add_966361 : sel_966358;
  assign add_966365 = sel_966362 + 8'h01;
  assign sel_966366 = array_index_965977 == array_index_949069 ? add_966365 : sel_966362;
  assign add_966369 = sel_966366 + 8'h01;
  assign sel_966370 = array_index_965977 == array_index_949075 ? add_966369 : sel_966366;
  assign add_966373 = sel_966370 + 8'h01;
  assign sel_966374 = array_index_965977 == array_index_949081 ? add_966373 : sel_966370;
  assign add_966378 = sel_966374 + 8'h01;
  assign array_index_966379 = set1_unflattened[7'h2c];
  assign sel_966380 = array_index_965977 == array_index_949087 ? add_966378 : sel_966374;
  assign add_966383 = sel_966380 + 8'h01;
  assign sel_966384 = array_index_966379 == array_index_948483 ? add_966383 : sel_966380;
  assign add_966387 = sel_966384 + 8'h01;
  assign sel_966388 = array_index_966379 == array_index_948487 ? add_966387 : sel_966384;
  assign add_966391 = sel_966388 + 8'h01;
  assign sel_966392 = array_index_966379 == array_index_948495 ? add_966391 : sel_966388;
  assign add_966395 = sel_966392 + 8'h01;
  assign sel_966396 = array_index_966379 == array_index_948503 ? add_966395 : sel_966392;
  assign add_966399 = sel_966396 + 8'h01;
  assign sel_966400 = array_index_966379 == array_index_948511 ? add_966399 : sel_966396;
  assign add_966403 = sel_966400 + 8'h01;
  assign sel_966404 = array_index_966379 == array_index_948519 ? add_966403 : sel_966400;
  assign add_966407 = sel_966404 + 8'h01;
  assign sel_966408 = array_index_966379 == array_index_948527 ? add_966407 : sel_966404;
  assign add_966411 = sel_966408 + 8'h01;
  assign sel_966412 = array_index_966379 == array_index_948535 ? add_966411 : sel_966408;
  assign add_966415 = sel_966412 + 8'h01;
  assign sel_966416 = array_index_966379 == array_index_948541 ? add_966415 : sel_966412;
  assign add_966419 = sel_966416 + 8'h01;
  assign sel_966420 = array_index_966379 == array_index_948547 ? add_966419 : sel_966416;
  assign add_966423 = sel_966420 + 8'h01;
  assign sel_966424 = array_index_966379 == array_index_948553 ? add_966423 : sel_966420;
  assign add_966427 = sel_966424 + 8'h01;
  assign sel_966428 = array_index_966379 == array_index_948559 ? add_966427 : sel_966424;
  assign add_966431 = sel_966428 + 8'h01;
  assign sel_966432 = array_index_966379 == array_index_948565 ? add_966431 : sel_966428;
  assign add_966435 = sel_966432 + 8'h01;
  assign sel_966436 = array_index_966379 == array_index_948571 ? add_966435 : sel_966432;
  assign add_966439 = sel_966436 + 8'h01;
  assign sel_966440 = array_index_966379 == array_index_948577 ? add_966439 : sel_966436;
  assign add_966443 = sel_966440 + 8'h01;
  assign sel_966444 = array_index_966379 == array_index_948583 ? add_966443 : sel_966440;
  assign add_966447 = sel_966444 + 8'h01;
  assign sel_966448 = array_index_966379 == array_index_948589 ? add_966447 : sel_966444;
  assign add_966451 = sel_966448 + 8'h01;
  assign sel_966452 = array_index_966379 == array_index_948595 ? add_966451 : sel_966448;
  assign add_966455 = sel_966452 + 8'h01;
  assign sel_966456 = array_index_966379 == array_index_948601 ? add_966455 : sel_966452;
  assign add_966459 = sel_966456 + 8'h01;
  assign sel_966460 = array_index_966379 == array_index_948607 ? add_966459 : sel_966456;
  assign add_966463 = sel_966460 + 8'h01;
  assign sel_966464 = array_index_966379 == array_index_948613 ? add_966463 : sel_966460;
  assign add_966467 = sel_966464 + 8'h01;
  assign sel_966468 = array_index_966379 == array_index_948619 ? add_966467 : sel_966464;
  assign add_966471 = sel_966468 + 8'h01;
  assign sel_966472 = array_index_966379 == array_index_948625 ? add_966471 : sel_966468;
  assign add_966475 = sel_966472 + 8'h01;
  assign sel_966476 = array_index_966379 == array_index_948631 ? add_966475 : sel_966472;
  assign add_966479 = sel_966476 + 8'h01;
  assign sel_966480 = array_index_966379 == array_index_948637 ? add_966479 : sel_966476;
  assign add_966483 = sel_966480 + 8'h01;
  assign sel_966484 = array_index_966379 == array_index_948643 ? add_966483 : sel_966480;
  assign add_966487 = sel_966484 + 8'h01;
  assign sel_966488 = array_index_966379 == array_index_948649 ? add_966487 : sel_966484;
  assign add_966491 = sel_966488 + 8'h01;
  assign sel_966492 = array_index_966379 == array_index_948655 ? add_966491 : sel_966488;
  assign add_966495 = sel_966492 + 8'h01;
  assign sel_966496 = array_index_966379 == array_index_948661 ? add_966495 : sel_966492;
  assign add_966499 = sel_966496 + 8'h01;
  assign sel_966500 = array_index_966379 == array_index_948667 ? add_966499 : sel_966496;
  assign add_966503 = sel_966500 + 8'h01;
  assign sel_966504 = array_index_966379 == array_index_948673 ? add_966503 : sel_966500;
  assign add_966507 = sel_966504 + 8'h01;
  assign sel_966508 = array_index_966379 == array_index_948679 ? add_966507 : sel_966504;
  assign add_966511 = sel_966508 + 8'h01;
  assign sel_966512 = array_index_966379 == array_index_948685 ? add_966511 : sel_966508;
  assign add_966515 = sel_966512 + 8'h01;
  assign sel_966516 = array_index_966379 == array_index_948691 ? add_966515 : sel_966512;
  assign add_966519 = sel_966516 + 8'h01;
  assign sel_966520 = array_index_966379 == array_index_948697 ? add_966519 : sel_966516;
  assign add_966523 = sel_966520 + 8'h01;
  assign sel_966524 = array_index_966379 == array_index_948703 ? add_966523 : sel_966520;
  assign add_966527 = sel_966524 + 8'h01;
  assign sel_966528 = array_index_966379 == array_index_948709 ? add_966527 : sel_966524;
  assign add_966531 = sel_966528 + 8'h01;
  assign sel_966532 = array_index_966379 == array_index_948715 ? add_966531 : sel_966528;
  assign add_966535 = sel_966532 + 8'h01;
  assign sel_966536 = array_index_966379 == array_index_948721 ? add_966535 : sel_966532;
  assign add_966539 = sel_966536 + 8'h01;
  assign sel_966540 = array_index_966379 == array_index_948727 ? add_966539 : sel_966536;
  assign add_966543 = sel_966540 + 8'h01;
  assign sel_966544 = array_index_966379 == array_index_948733 ? add_966543 : sel_966540;
  assign add_966547 = sel_966544 + 8'h01;
  assign sel_966548 = array_index_966379 == array_index_948739 ? add_966547 : sel_966544;
  assign add_966551 = sel_966548 + 8'h01;
  assign sel_966552 = array_index_966379 == array_index_948745 ? add_966551 : sel_966548;
  assign add_966555 = sel_966552 + 8'h01;
  assign sel_966556 = array_index_966379 == array_index_948751 ? add_966555 : sel_966552;
  assign add_966559 = sel_966556 + 8'h01;
  assign sel_966560 = array_index_966379 == array_index_948757 ? add_966559 : sel_966556;
  assign add_966563 = sel_966560 + 8'h01;
  assign sel_966564 = array_index_966379 == array_index_948763 ? add_966563 : sel_966560;
  assign add_966567 = sel_966564 + 8'h01;
  assign sel_966568 = array_index_966379 == array_index_948769 ? add_966567 : sel_966564;
  assign add_966571 = sel_966568 + 8'h01;
  assign sel_966572 = array_index_966379 == array_index_948775 ? add_966571 : sel_966568;
  assign add_966575 = sel_966572 + 8'h01;
  assign sel_966576 = array_index_966379 == array_index_948781 ? add_966575 : sel_966572;
  assign add_966579 = sel_966576 + 8'h01;
  assign sel_966580 = array_index_966379 == array_index_948787 ? add_966579 : sel_966576;
  assign add_966583 = sel_966580 + 8'h01;
  assign sel_966584 = array_index_966379 == array_index_948793 ? add_966583 : sel_966580;
  assign add_966587 = sel_966584 + 8'h01;
  assign sel_966588 = array_index_966379 == array_index_948799 ? add_966587 : sel_966584;
  assign add_966591 = sel_966588 + 8'h01;
  assign sel_966592 = array_index_966379 == array_index_948805 ? add_966591 : sel_966588;
  assign add_966595 = sel_966592 + 8'h01;
  assign sel_966596 = array_index_966379 == array_index_948811 ? add_966595 : sel_966592;
  assign add_966599 = sel_966596 + 8'h01;
  assign sel_966600 = array_index_966379 == array_index_948817 ? add_966599 : sel_966596;
  assign add_966603 = sel_966600 + 8'h01;
  assign sel_966604 = array_index_966379 == array_index_948823 ? add_966603 : sel_966600;
  assign add_966607 = sel_966604 + 8'h01;
  assign sel_966608 = array_index_966379 == array_index_948829 ? add_966607 : sel_966604;
  assign add_966611 = sel_966608 + 8'h01;
  assign sel_966612 = array_index_966379 == array_index_948835 ? add_966611 : sel_966608;
  assign add_966615 = sel_966612 + 8'h01;
  assign sel_966616 = array_index_966379 == array_index_948841 ? add_966615 : sel_966612;
  assign add_966619 = sel_966616 + 8'h01;
  assign sel_966620 = array_index_966379 == array_index_948847 ? add_966619 : sel_966616;
  assign add_966623 = sel_966620 + 8'h01;
  assign sel_966624 = array_index_966379 == array_index_948853 ? add_966623 : sel_966620;
  assign add_966627 = sel_966624 + 8'h01;
  assign sel_966628 = array_index_966379 == array_index_948859 ? add_966627 : sel_966624;
  assign add_966631 = sel_966628 + 8'h01;
  assign sel_966632 = array_index_966379 == array_index_948865 ? add_966631 : sel_966628;
  assign add_966635 = sel_966632 + 8'h01;
  assign sel_966636 = array_index_966379 == array_index_948871 ? add_966635 : sel_966632;
  assign add_966639 = sel_966636 + 8'h01;
  assign sel_966640 = array_index_966379 == array_index_948877 ? add_966639 : sel_966636;
  assign add_966643 = sel_966640 + 8'h01;
  assign sel_966644 = array_index_966379 == array_index_948883 ? add_966643 : sel_966640;
  assign add_966647 = sel_966644 + 8'h01;
  assign sel_966648 = array_index_966379 == array_index_948889 ? add_966647 : sel_966644;
  assign add_966651 = sel_966648 + 8'h01;
  assign sel_966652 = array_index_966379 == array_index_948895 ? add_966651 : sel_966648;
  assign add_966655 = sel_966652 + 8'h01;
  assign sel_966656 = array_index_966379 == array_index_948901 ? add_966655 : sel_966652;
  assign add_966659 = sel_966656 + 8'h01;
  assign sel_966660 = array_index_966379 == array_index_948907 ? add_966659 : sel_966656;
  assign add_966663 = sel_966660 + 8'h01;
  assign sel_966664 = array_index_966379 == array_index_948913 ? add_966663 : sel_966660;
  assign add_966667 = sel_966664 + 8'h01;
  assign sel_966668 = array_index_966379 == array_index_948919 ? add_966667 : sel_966664;
  assign add_966671 = sel_966668 + 8'h01;
  assign sel_966672 = array_index_966379 == array_index_948925 ? add_966671 : sel_966668;
  assign add_966675 = sel_966672 + 8'h01;
  assign sel_966676 = array_index_966379 == array_index_948931 ? add_966675 : sel_966672;
  assign add_966679 = sel_966676 + 8'h01;
  assign sel_966680 = array_index_966379 == array_index_948937 ? add_966679 : sel_966676;
  assign add_966683 = sel_966680 + 8'h01;
  assign sel_966684 = array_index_966379 == array_index_948943 ? add_966683 : sel_966680;
  assign add_966687 = sel_966684 + 8'h01;
  assign sel_966688 = array_index_966379 == array_index_948949 ? add_966687 : sel_966684;
  assign add_966691 = sel_966688 + 8'h01;
  assign sel_966692 = array_index_966379 == array_index_948955 ? add_966691 : sel_966688;
  assign add_966695 = sel_966692 + 8'h01;
  assign sel_966696 = array_index_966379 == array_index_948961 ? add_966695 : sel_966692;
  assign add_966699 = sel_966696 + 8'h01;
  assign sel_966700 = array_index_966379 == array_index_948967 ? add_966699 : sel_966696;
  assign add_966703 = sel_966700 + 8'h01;
  assign sel_966704 = array_index_966379 == array_index_948973 ? add_966703 : sel_966700;
  assign add_966707 = sel_966704 + 8'h01;
  assign sel_966708 = array_index_966379 == array_index_948979 ? add_966707 : sel_966704;
  assign add_966711 = sel_966708 + 8'h01;
  assign sel_966712 = array_index_966379 == array_index_948985 ? add_966711 : sel_966708;
  assign add_966715 = sel_966712 + 8'h01;
  assign sel_966716 = array_index_966379 == array_index_948991 ? add_966715 : sel_966712;
  assign add_966719 = sel_966716 + 8'h01;
  assign sel_966720 = array_index_966379 == array_index_948997 ? add_966719 : sel_966716;
  assign add_966723 = sel_966720 + 8'h01;
  assign sel_966724 = array_index_966379 == array_index_949003 ? add_966723 : sel_966720;
  assign add_966727 = sel_966724 + 8'h01;
  assign sel_966728 = array_index_966379 == array_index_949009 ? add_966727 : sel_966724;
  assign add_966731 = sel_966728 + 8'h01;
  assign sel_966732 = array_index_966379 == array_index_949015 ? add_966731 : sel_966728;
  assign add_966735 = sel_966732 + 8'h01;
  assign sel_966736 = array_index_966379 == array_index_949021 ? add_966735 : sel_966732;
  assign add_966739 = sel_966736 + 8'h01;
  assign sel_966740 = array_index_966379 == array_index_949027 ? add_966739 : sel_966736;
  assign add_966743 = sel_966740 + 8'h01;
  assign sel_966744 = array_index_966379 == array_index_949033 ? add_966743 : sel_966740;
  assign add_966747 = sel_966744 + 8'h01;
  assign sel_966748 = array_index_966379 == array_index_949039 ? add_966747 : sel_966744;
  assign add_966751 = sel_966748 + 8'h01;
  assign sel_966752 = array_index_966379 == array_index_949045 ? add_966751 : sel_966748;
  assign add_966755 = sel_966752 + 8'h01;
  assign sel_966756 = array_index_966379 == array_index_949051 ? add_966755 : sel_966752;
  assign add_966759 = sel_966756 + 8'h01;
  assign sel_966760 = array_index_966379 == array_index_949057 ? add_966759 : sel_966756;
  assign add_966763 = sel_966760 + 8'h01;
  assign sel_966764 = array_index_966379 == array_index_949063 ? add_966763 : sel_966760;
  assign add_966767 = sel_966764 + 8'h01;
  assign sel_966768 = array_index_966379 == array_index_949069 ? add_966767 : sel_966764;
  assign add_966771 = sel_966768 + 8'h01;
  assign sel_966772 = array_index_966379 == array_index_949075 ? add_966771 : sel_966768;
  assign add_966775 = sel_966772 + 8'h01;
  assign sel_966776 = array_index_966379 == array_index_949081 ? add_966775 : sel_966772;
  assign add_966780 = sel_966776 + 8'h01;
  assign array_index_966781 = set1_unflattened[7'h2d];
  assign sel_966782 = array_index_966379 == array_index_949087 ? add_966780 : sel_966776;
  assign add_966785 = sel_966782 + 8'h01;
  assign sel_966786 = array_index_966781 == array_index_948483 ? add_966785 : sel_966782;
  assign add_966789 = sel_966786 + 8'h01;
  assign sel_966790 = array_index_966781 == array_index_948487 ? add_966789 : sel_966786;
  assign add_966793 = sel_966790 + 8'h01;
  assign sel_966794 = array_index_966781 == array_index_948495 ? add_966793 : sel_966790;
  assign add_966797 = sel_966794 + 8'h01;
  assign sel_966798 = array_index_966781 == array_index_948503 ? add_966797 : sel_966794;
  assign add_966801 = sel_966798 + 8'h01;
  assign sel_966802 = array_index_966781 == array_index_948511 ? add_966801 : sel_966798;
  assign add_966805 = sel_966802 + 8'h01;
  assign sel_966806 = array_index_966781 == array_index_948519 ? add_966805 : sel_966802;
  assign add_966809 = sel_966806 + 8'h01;
  assign sel_966810 = array_index_966781 == array_index_948527 ? add_966809 : sel_966806;
  assign add_966813 = sel_966810 + 8'h01;
  assign sel_966814 = array_index_966781 == array_index_948535 ? add_966813 : sel_966810;
  assign add_966817 = sel_966814 + 8'h01;
  assign sel_966818 = array_index_966781 == array_index_948541 ? add_966817 : sel_966814;
  assign add_966821 = sel_966818 + 8'h01;
  assign sel_966822 = array_index_966781 == array_index_948547 ? add_966821 : sel_966818;
  assign add_966825 = sel_966822 + 8'h01;
  assign sel_966826 = array_index_966781 == array_index_948553 ? add_966825 : sel_966822;
  assign add_966829 = sel_966826 + 8'h01;
  assign sel_966830 = array_index_966781 == array_index_948559 ? add_966829 : sel_966826;
  assign add_966833 = sel_966830 + 8'h01;
  assign sel_966834 = array_index_966781 == array_index_948565 ? add_966833 : sel_966830;
  assign add_966837 = sel_966834 + 8'h01;
  assign sel_966838 = array_index_966781 == array_index_948571 ? add_966837 : sel_966834;
  assign add_966841 = sel_966838 + 8'h01;
  assign sel_966842 = array_index_966781 == array_index_948577 ? add_966841 : sel_966838;
  assign add_966845 = sel_966842 + 8'h01;
  assign sel_966846 = array_index_966781 == array_index_948583 ? add_966845 : sel_966842;
  assign add_966849 = sel_966846 + 8'h01;
  assign sel_966850 = array_index_966781 == array_index_948589 ? add_966849 : sel_966846;
  assign add_966853 = sel_966850 + 8'h01;
  assign sel_966854 = array_index_966781 == array_index_948595 ? add_966853 : sel_966850;
  assign add_966857 = sel_966854 + 8'h01;
  assign sel_966858 = array_index_966781 == array_index_948601 ? add_966857 : sel_966854;
  assign add_966861 = sel_966858 + 8'h01;
  assign sel_966862 = array_index_966781 == array_index_948607 ? add_966861 : sel_966858;
  assign add_966865 = sel_966862 + 8'h01;
  assign sel_966866 = array_index_966781 == array_index_948613 ? add_966865 : sel_966862;
  assign add_966869 = sel_966866 + 8'h01;
  assign sel_966870 = array_index_966781 == array_index_948619 ? add_966869 : sel_966866;
  assign add_966873 = sel_966870 + 8'h01;
  assign sel_966874 = array_index_966781 == array_index_948625 ? add_966873 : sel_966870;
  assign add_966877 = sel_966874 + 8'h01;
  assign sel_966878 = array_index_966781 == array_index_948631 ? add_966877 : sel_966874;
  assign add_966881 = sel_966878 + 8'h01;
  assign sel_966882 = array_index_966781 == array_index_948637 ? add_966881 : sel_966878;
  assign add_966885 = sel_966882 + 8'h01;
  assign sel_966886 = array_index_966781 == array_index_948643 ? add_966885 : sel_966882;
  assign add_966889 = sel_966886 + 8'h01;
  assign sel_966890 = array_index_966781 == array_index_948649 ? add_966889 : sel_966886;
  assign add_966893 = sel_966890 + 8'h01;
  assign sel_966894 = array_index_966781 == array_index_948655 ? add_966893 : sel_966890;
  assign add_966897 = sel_966894 + 8'h01;
  assign sel_966898 = array_index_966781 == array_index_948661 ? add_966897 : sel_966894;
  assign add_966901 = sel_966898 + 8'h01;
  assign sel_966902 = array_index_966781 == array_index_948667 ? add_966901 : sel_966898;
  assign add_966905 = sel_966902 + 8'h01;
  assign sel_966906 = array_index_966781 == array_index_948673 ? add_966905 : sel_966902;
  assign add_966909 = sel_966906 + 8'h01;
  assign sel_966910 = array_index_966781 == array_index_948679 ? add_966909 : sel_966906;
  assign add_966913 = sel_966910 + 8'h01;
  assign sel_966914 = array_index_966781 == array_index_948685 ? add_966913 : sel_966910;
  assign add_966917 = sel_966914 + 8'h01;
  assign sel_966918 = array_index_966781 == array_index_948691 ? add_966917 : sel_966914;
  assign add_966921 = sel_966918 + 8'h01;
  assign sel_966922 = array_index_966781 == array_index_948697 ? add_966921 : sel_966918;
  assign add_966925 = sel_966922 + 8'h01;
  assign sel_966926 = array_index_966781 == array_index_948703 ? add_966925 : sel_966922;
  assign add_966929 = sel_966926 + 8'h01;
  assign sel_966930 = array_index_966781 == array_index_948709 ? add_966929 : sel_966926;
  assign add_966933 = sel_966930 + 8'h01;
  assign sel_966934 = array_index_966781 == array_index_948715 ? add_966933 : sel_966930;
  assign add_966937 = sel_966934 + 8'h01;
  assign sel_966938 = array_index_966781 == array_index_948721 ? add_966937 : sel_966934;
  assign add_966941 = sel_966938 + 8'h01;
  assign sel_966942 = array_index_966781 == array_index_948727 ? add_966941 : sel_966938;
  assign add_966945 = sel_966942 + 8'h01;
  assign sel_966946 = array_index_966781 == array_index_948733 ? add_966945 : sel_966942;
  assign add_966949 = sel_966946 + 8'h01;
  assign sel_966950 = array_index_966781 == array_index_948739 ? add_966949 : sel_966946;
  assign add_966953 = sel_966950 + 8'h01;
  assign sel_966954 = array_index_966781 == array_index_948745 ? add_966953 : sel_966950;
  assign add_966957 = sel_966954 + 8'h01;
  assign sel_966958 = array_index_966781 == array_index_948751 ? add_966957 : sel_966954;
  assign add_966961 = sel_966958 + 8'h01;
  assign sel_966962 = array_index_966781 == array_index_948757 ? add_966961 : sel_966958;
  assign add_966965 = sel_966962 + 8'h01;
  assign sel_966966 = array_index_966781 == array_index_948763 ? add_966965 : sel_966962;
  assign add_966969 = sel_966966 + 8'h01;
  assign sel_966970 = array_index_966781 == array_index_948769 ? add_966969 : sel_966966;
  assign add_966973 = sel_966970 + 8'h01;
  assign sel_966974 = array_index_966781 == array_index_948775 ? add_966973 : sel_966970;
  assign add_966977 = sel_966974 + 8'h01;
  assign sel_966978 = array_index_966781 == array_index_948781 ? add_966977 : sel_966974;
  assign add_966981 = sel_966978 + 8'h01;
  assign sel_966982 = array_index_966781 == array_index_948787 ? add_966981 : sel_966978;
  assign add_966985 = sel_966982 + 8'h01;
  assign sel_966986 = array_index_966781 == array_index_948793 ? add_966985 : sel_966982;
  assign add_966989 = sel_966986 + 8'h01;
  assign sel_966990 = array_index_966781 == array_index_948799 ? add_966989 : sel_966986;
  assign add_966993 = sel_966990 + 8'h01;
  assign sel_966994 = array_index_966781 == array_index_948805 ? add_966993 : sel_966990;
  assign add_966997 = sel_966994 + 8'h01;
  assign sel_966998 = array_index_966781 == array_index_948811 ? add_966997 : sel_966994;
  assign add_967001 = sel_966998 + 8'h01;
  assign sel_967002 = array_index_966781 == array_index_948817 ? add_967001 : sel_966998;
  assign add_967005 = sel_967002 + 8'h01;
  assign sel_967006 = array_index_966781 == array_index_948823 ? add_967005 : sel_967002;
  assign add_967009 = sel_967006 + 8'h01;
  assign sel_967010 = array_index_966781 == array_index_948829 ? add_967009 : sel_967006;
  assign add_967013 = sel_967010 + 8'h01;
  assign sel_967014 = array_index_966781 == array_index_948835 ? add_967013 : sel_967010;
  assign add_967017 = sel_967014 + 8'h01;
  assign sel_967018 = array_index_966781 == array_index_948841 ? add_967017 : sel_967014;
  assign add_967021 = sel_967018 + 8'h01;
  assign sel_967022 = array_index_966781 == array_index_948847 ? add_967021 : sel_967018;
  assign add_967025 = sel_967022 + 8'h01;
  assign sel_967026 = array_index_966781 == array_index_948853 ? add_967025 : sel_967022;
  assign add_967029 = sel_967026 + 8'h01;
  assign sel_967030 = array_index_966781 == array_index_948859 ? add_967029 : sel_967026;
  assign add_967033 = sel_967030 + 8'h01;
  assign sel_967034 = array_index_966781 == array_index_948865 ? add_967033 : sel_967030;
  assign add_967037 = sel_967034 + 8'h01;
  assign sel_967038 = array_index_966781 == array_index_948871 ? add_967037 : sel_967034;
  assign add_967041 = sel_967038 + 8'h01;
  assign sel_967042 = array_index_966781 == array_index_948877 ? add_967041 : sel_967038;
  assign add_967045 = sel_967042 + 8'h01;
  assign sel_967046 = array_index_966781 == array_index_948883 ? add_967045 : sel_967042;
  assign add_967049 = sel_967046 + 8'h01;
  assign sel_967050 = array_index_966781 == array_index_948889 ? add_967049 : sel_967046;
  assign add_967053 = sel_967050 + 8'h01;
  assign sel_967054 = array_index_966781 == array_index_948895 ? add_967053 : sel_967050;
  assign add_967057 = sel_967054 + 8'h01;
  assign sel_967058 = array_index_966781 == array_index_948901 ? add_967057 : sel_967054;
  assign add_967061 = sel_967058 + 8'h01;
  assign sel_967062 = array_index_966781 == array_index_948907 ? add_967061 : sel_967058;
  assign add_967065 = sel_967062 + 8'h01;
  assign sel_967066 = array_index_966781 == array_index_948913 ? add_967065 : sel_967062;
  assign add_967069 = sel_967066 + 8'h01;
  assign sel_967070 = array_index_966781 == array_index_948919 ? add_967069 : sel_967066;
  assign add_967073 = sel_967070 + 8'h01;
  assign sel_967074 = array_index_966781 == array_index_948925 ? add_967073 : sel_967070;
  assign add_967077 = sel_967074 + 8'h01;
  assign sel_967078 = array_index_966781 == array_index_948931 ? add_967077 : sel_967074;
  assign add_967081 = sel_967078 + 8'h01;
  assign sel_967082 = array_index_966781 == array_index_948937 ? add_967081 : sel_967078;
  assign add_967085 = sel_967082 + 8'h01;
  assign sel_967086 = array_index_966781 == array_index_948943 ? add_967085 : sel_967082;
  assign add_967089 = sel_967086 + 8'h01;
  assign sel_967090 = array_index_966781 == array_index_948949 ? add_967089 : sel_967086;
  assign add_967093 = sel_967090 + 8'h01;
  assign sel_967094 = array_index_966781 == array_index_948955 ? add_967093 : sel_967090;
  assign add_967097 = sel_967094 + 8'h01;
  assign sel_967098 = array_index_966781 == array_index_948961 ? add_967097 : sel_967094;
  assign add_967101 = sel_967098 + 8'h01;
  assign sel_967102 = array_index_966781 == array_index_948967 ? add_967101 : sel_967098;
  assign add_967105 = sel_967102 + 8'h01;
  assign sel_967106 = array_index_966781 == array_index_948973 ? add_967105 : sel_967102;
  assign add_967109 = sel_967106 + 8'h01;
  assign sel_967110 = array_index_966781 == array_index_948979 ? add_967109 : sel_967106;
  assign add_967113 = sel_967110 + 8'h01;
  assign sel_967114 = array_index_966781 == array_index_948985 ? add_967113 : sel_967110;
  assign add_967117 = sel_967114 + 8'h01;
  assign sel_967118 = array_index_966781 == array_index_948991 ? add_967117 : sel_967114;
  assign add_967121 = sel_967118 + 8'h01;
  assign sel_967122 = array_index_966781 == array_index_948997 ? add_967121 : sel_967118;
  assign add_967125 = sel_967122 + 8'h01;
  assign sel_967126 = array_index_966781 == array_index_949003 ? add_967125 : sel_967122;
  assign add_967129 = sel_967126 + 8'h01;
  assign sel_967130 = array_index_966781 == array_index_949009 ? add_967129 : sel_967126;
  assign add_967133 = sel_967130 + 8'h01;
  assign sel_967134 = array_index_966781 == array_index_949015 ? add_967133 : sel_967130;
  assign add_967137 = sel_967134 + 8'h01;
  assign sel_967138 = array_index_966781 == array_index_949021 ? add_967137 : sel_967134;
  assign add_967141 = sel_967138 + 8'h01;
  assign sel_967142 = array_index_966781 == array_index_949027 ? add_967141 : sel_967138;
  assign add_967145 = sel_967142 + 8'h01;
  assign sel_967146 = array_index_966781 == array_index_949033 ? add_967145 : sel_967142;
  assign add_967149 = sel_967146 + 8'h01;
  assign sel_967150 = array_index_966781 == array_index_949039 ? add_967149 : sel_967146;
  assign add_967153 = sel_967150 + 8'h01;
  assign sel_967154 = array_index_966781 == array_index_949045 ? add_967153 : sel_967150;
  assign add_967157 = sel_967154 + 8'h01;
  assign sel_967158 = array_index_966781 == array_index_949051 ? add_967157 : sel_967154;
  assign add_967161 = sel_967158 + 8'h01;
  assign sel_967162 = array_index_966781 == array_index_949057 ? add_967161 : sel_967158;
  assign add_967165 = sel_967162 + 8'h01;
  assign sel_967166 = array_index_966781 == array_index_949063 ? add_967165 : sel_967162;
  assign add_967169 = sel_967166 + 8'h01;
  assign sel_967170 = array_index_966781 == array_index_949069 ? add_967169 : sel_967166;
  assign add_967173 = sel_967170 + 8'h01;
  assign sel_967174 = array_index_966781 == array_index_949075 ? add_967173 : sel_967170;
  assign add_967177 = sel_967174 + 8'h01;
  assign sel_967178 = array_index_966781 == array_index_949081 ? add_967177 : sel_967174;
  assign add_967182 = sel_967178 + 8'h01;
  assign array_index_967183 = set1_unflattened[7'h2e];
  assign sel_967184 = array_index_966781 == array_index_949087 ? add_967182 : sel_967178;
  assign add_967187 = sel_967184 + 8'h01;
  assign sel_967188 = array_index_967183 == array_index_948483 ? add_967187 : sel_967184;
  assign add_967191 = sel_967188 + 8'h01;
  assign sel_967192 = array_index_967183 == array_index_948487 ? add_967191 : sel_967188;
  assign add_967195 = sel_967192 + 8'h01;
  assign sel_967196 = array_index_967183 == array_index_948495 ? add_967195 : sel_967192;
  assign add_967199 = sel_967196 + 8'h01;
  assign sel_967200 = array_index_967183 == array_index_948503 ? add_967199 : sel_967196;
  assign add_967203 = sel_967200 + 8'h01;
  assign sel_967204 = array_index_967183 == array_index_948511 ? add_967203 : sel_967200;
  assign add_967207 = sel_967204 + 8'h01;
  assign sel_967208 = array_index_967183 == array_index_948519 ? add_967207 : sel_967204;
  assign add_967211 = sel_967208 + 8'h01;
  assign sel_967212 = array_index_967183 == array_index_948527 ? add_967211 : sel_967208;
  assign add_967215 = sel_967212 + 8'h01;
  assign sel_967216 = array_index_967183 == array_index_948535 ? add_967215 : sel_967212;
  assign add_967219 = sel_967216 + 8'h01;
  assign sel_967220 = array_index_967183 == array_index_948541 ? add_967219 : sel_967216;
  assign add_967223 = sel_967220 + 8'h01;
  assign sel_967224 = array_index_967183 == array_index_948547 ? add_967223 : sel_967220;
  assign add_967227 = sel_967224 + 8'h01;
  assign sel_967228 = array_index_967183 == array_index_948553 ? add_967227 : sel_967224;
  assign add_967231 = sel_967228 + 8'h01;
  assign sel_967232 = array_index_967183 == array_index_948559 ? add_967231 : sel_967228;
  assign add_967235 = sel_967232 + 8'h01;
  assign sel_967236 = array_index_967183 == array_index_948565 ? add_967235 : sel_967232;
  assign add_967239 = sel_967236 + 8'h01;
  assign sel_967240 = array_index_967183 == array_index_948571 ? add_967239 : sel_967236;
  assign add_967243 = sel_967240 + 8'h01;
  assign sel_967244 = array_index_967183 == array_index_948577 ? add_967243 : sel_967240;
  assign add_967247 = sel_967244 + 8'h01;
  assign sel_967248 = array_index_967183 == array_index_948583 ? add_967247 : sel_967244;
  assign add_967251 = sel_967248 + 8'h01;
  assign sel_967252 = array_index_967183 == array_index_948589 ? add_967251 : sel_967248;
  assign add_967255 = sel_967252 + 8'h01;
  assign sel_967256 = array_index_967183 == array_index_948595 ? add_967255 : sel_967252;
  assign add_967259 = sel_967256 + 8'h01;
  assign sel_967260 = array_index_967183 == array_index_948601 ? add_967259 : sel_967256;
  assign add_967263 = sel_967260 + 8'h01;
  assign sel_967264 = array_index_967183 == array_index_948607 ? add_967263 : sel_967260;
  assign add_967267 = sel_967264 + 8'h01;
  assign sel_967268 = array_index_967183 == array_index_948613 ? add_967267 : sel_967264;
  assign add_967271 = sel_967268 + 8'h01;
  assign sel_967272 = array_index_967183 == array_index_948619 ? add_967271 : sel_967268;
  assign add_967275 = sel_967272 + 8'h01;
  assign sel_967276 = array_index_967183 == array_index_948625 ? add_967275 : sel_967272;
  assign add_967279 = sel_967276 + 8'h01;
  assign sel_967280 = array_index_967183 == array_index_948631 ? add_967279 : sel_967276;
  assign add_967283 = sel_967280 + 8'h01;
  assign sel_967284 = array_index_967183 == array_index_948637 ? add_967283 : sel_967280;
  assign add_967287 = sel_967284 + 8'h01;
  assign sel_967288 = array_index_967183 == array_index_948643 ? add_967287 : sel_967284;
  assign add_967291 = sel_967288 + 8'h01;
  assign sel_967292 = array_index_967183 == array_index_948649 ? add_967291 : sel_967288;
  assign add_967295 = sel_967292 + 8'h01;
  assign sel_967296 = array_index_967183 == array_index_948655 ? add_967295 : sel_967292;
  assign add_967299 = sel_967296 + 8'h01;
  assign sel_967300 = array_index_967183 == array_index_948661 ? add_967299 : sel_967296;
  assign add_967303 = sel_967300 + 8'h01;
  assign sel_967304 = array_index_967183 == array_index_948667 ? add_967303 : sel_967300;
  assign add_967307 = sel_967304 + 8'h01;
  assign sel_967308 = array_index_967183 == array_index_948673 ? add_967307 : sel_967304;
  assign add_967311 = sel_967308 + 8'h01;
  assign sel_967312 = array_index_967183 == array_index_948679 ? add_967311 : sel_967308;
  assign add_967315 = sel_967312 + 8'h01;
  assign sel_967316 = array_index_967183 == array_index_948685 ? add_967315 : sel_967312;
  assign add_967319 = sel_967316 + 8'h01;
  assign sel_967320 = array_index_967183 == array_index_948691 ? add_967319 : sel_967316;
  assign add_967323 = sel_967320 + 8'h01;
  assign sel_967324 = array_index_967183 == array_index_948697 ? add_967323 : sel_967320;
  assign add_967327 = sel_967324 + 8'h01;
  assign sel_967328 = array_index_967183 == array_index_948703 ? add_967327 : sel_967324;
  assign add_967331 = sel_967328 + 8'h01;
  assign sel_967332 = array_index_967183 == array_index_948709 ? add_967331 : sel_967328;
  assign add_967335 = sel_967332 + 8'h01;
  assign sel_967336 = array_index_967183 == array_index_948715 ? add_967335 : sel_967332;
  assign add_967339 = sel_967336 + 8'h01;
  assign sel_967340 = array_index_967183 == array_index_948721 ? add_967339 : sel_967336;
  assign add_967343 = sel_967340 + 8'h01;
  assign sel_967344 = array_index_967183 == array_index_948727 ? add_967343 : sel_967340;
  assign add_967347 = sel_967344 + 8'h01;
  assign sel_967348 = array_index_967183 == array_index_948733 ? add_967347 : sel_967344;
  assign add_967351 = sel_967348 + 8'h01;
  assign sel_967352 = array_index_967183 == array_index_948739 ? add_967351 : sel_967348;
  assign add_967355 = sel_967352 + 8'h01;
  assign sel_967356 = array_index_967183 == array_index_948745 ? add_967355 : sel_967352;
  assign add_967359 = sel_967356 + 8'h01;
  assign sel_967360 = array_index_967183 == array_index_948751 ? add_967359 : sel_967356;
  assign add_967363 = sel_967360 + 8'h01;
  assign sel_967364 = array_index_967183 == array_index_948757 ? add_967363 : sel_967360;
  assign add_967367 = sel_967364 + 8'h01;
  assign sel_967368 = array_index_967183 == array_index_948763 ? add_967367 : sel_967364;
  assign add_967371 = sel_967368 + 8'h01;
  assign sel_967372 = array_index_967183 == array_index_948769 ? add_967371 : sel_967368;
  assign add_967375 = sel_967372 + 8'h01;
  assign sel_967376 = array_index_967183 == array_index_948775 ? add_967375 : sel_967372;
  assign add_967379 = sel_967376 + 8'h01;
  assign sel_967380 = array_index_967183 == array_index_948781 ? add_967379 : sel_967376;
  assign add_967383 = sel_967380 + 8'h01;
  assign sel_967384 = array_index_967183 == array_index_948787 ? add_967383 : sel_967380;
  assign add_967387 = sel_967384 + 8'h01;
  assign sel_967388 = array_index_967183 == array_index_948793 ? add_967387 : sel_967384;
  assign add_967391 = sel_967388 + 8'h01;
  assign sel_967392 = array_index_967183 == array_index_948799 ? add_967391 : sel_967388;
  assign add_967395 = sel_967392 + 8'h01;
  assign sel_967396 = array_index_967183 == array_index_948805 ? add_967395 : sel_967392;
  assign add_967399 = sel_967396 + 8'h01;
  assign sel_967400 = array_index_967183 == array_index_948811 ? add_967399 : sel_967396;
  assign add_967403 = sel_967400 + 8'h01;
  assign sel_967404 = array_index_967183 == array_index_948817 ? add_967403 : sel_967400;
  assign add_967407 = sel_967404 + 8'h01;
  assign sel_967408 = array_index_967183 == array_index_948823 ? add_967407 : sel_967404;
  assign add_967411 = sel_967408 + 8'h01;
  assign sel_967412 = array_index_967183 == array_index_948829 ? add_967411 : sel_967408;
  assign add_967415 = sel_967412 + 8'h01;
  assign sel_967416 = array_index_967183 == array_index_948835 ? add_967415 : sel_967412;
  assign add_967419 = sel_967416 + 8'h01;
  assign sel_967420 = array_index_967183 == array_index_948841 ? add_967419 : sel_967416;
  assign add_967423 = sel_967420 + 8'h01;
  assign sel_967424 = array_index_967183 == array_index_948847 ? add_967423 : sel_967420;
  assign add_967427 = sel_967424 + 8'h01;
  assign sel_967428 = array_index_967183 == array_index_948853 ? add_967427 : sel_967424;
  assign add_967431 = sel_967428 + 8'h01;
  assign sel_967432 = array_index_967183 == array_index_948859 ? add_967431 : sel_967428;
  assign add_967435 = sel_967432 + 8'h01;
  assign sel_967436 = array_index_967183 == array_index_948865 ? add_967435 : sel_967432;
  assign add_967439 = sel_967436 + 8'h01;
  assign sel_967440 = array_index_967183 == array_index_948871 ? add_967439 : sel_967436;
  assign add_967443 = sel_967440 + 8'h01;
  assign sel_967444 = array_index_967183 == array_index_948877 ? add_967443 : sel_967440;
  assign add_967447 = sel_967444 + 8'h01;
  assign sel_967448 = array_index_967183 == array_index_948883 ? add_967447 : sel_967444;
  assign add_967451 = sel_967448 + 8'h01;
  assign sel_967452 = array_index_967183 == array_index_948889 ? add_967451 : sel_967448;
  assign add_967455 = sel_967452 + 8'h01;
  assign sel_967456 = array_index_967183 == array_index_948895 ? add_967455 : sel_967452;
  assign add_967459 = sel_967456 + 8'h01;
  assign sel_967460 = array_index_967183 == array_index_948901 ? add_967459 : sel_967456;
  assign add_967463 = sel_967460 + 8'h01;
  assign sel_967464 = array_index_967183 == array_index_948907 ? add_967463 : sel_967460;
  assign add_967467 = sel_967464 + 8'h01;
  assign sel_967468 = array_index_967183 == array_index_948913 ? add_967467 : sel_967464;
  assign add_967471 = sel_967468 + 8'h01;
  assign sel_967472 = array_index_967183 == array_index_948919 ? add_967471 : sel_967468;
  assign add_967475 = sel_967472 + 8'h01;
  assign sel_967476 = array_index_967183 == array_index_948925 ? add_967475 : sel_967472;
  assign add_967479 = sel_967476 + 8'h01;
  assign sel_967480 = array_index_967183 == array_index_948931 ? add_967479 : sel_967476;
  assign add_967483 = sel_967480 + 8'h01;
  assign sel_967484 = array_index_967183 == array_index_948937 ? add_967483 : sel_967480;
  assign add_967487 = sel_967484 + 8'h01;
  assign sel_967488 = array_index_967183 == array_index_948943 ? add_967487 : sel_967484;
  assign add_967491 = sel_967488 + 8'h01;
  assign sel_967492 = array_index_967183 == array_index_948949 ? add_967491 : sel_967488;
  assign add_967495 = sel_967492 + 8'h01;
  assign sel_967496 = array_index_967183 == array_index_948955 ? add_967495 : sel_967492;
  assign add_967499 = sel_967496 + 8'h01;
  assign sel_967500 = array_index_967183 == array_index_948961 ? add_967499 : sel_967496;
  assign add_967503 = sel_967500 + 8'h01;
  assign sel_967504 = array_index_967183 == array_index_948967 ? add_967503 : sel_967500;
  assign add_967507 = sel_967504 + 8'h01;
  assign sel_967508 = array_index_967183 == array_index_948973 ? add_967507 : sel_967504;
  assign add_967511 = sel_967508 + 8'h01;
  assign sel_967512 = array_index_967183 == array_index_948979 ? add_967511 : sel_967508;
  assign add_967515 = sel_967512 + 8'h01;
  assign sel_967516 = array_index_967183 == array_index_948985 ? add_967515 : sel_967512;
  assign add_967519 = sel_967516 + 8'h01;
  assign sel_967520 = array_index_967183 == array_index_948991 ? add_967519 : sel_967516;
  assign add_967523 = sel_967520 + 8'h01;
  assign sel_967524 = array_index_967183 == array_index_948997 ? add_967523 : sel_967520;
  assign add_967527 = sel_967524 + 8'h01;
  assign sel_967528 = array_index_967183 == array_index_949003 ? add_967527 : sel_967524;
  assign add_967531 = sel_967528 + 8'h01;
  assign sel_967532 = array_index_967183 == array_index_949009 ? add_967531 : sel_967528;
  assign add_967535 = sel_967532 + 8'h01;
  assign sel_967536 = array_index_967183 == array_index_949015 ? add_967535 : sel_967532;
  assign add_967539 = sel_967536 + 8'h01;
  assign sel_967540 = array_index_967183 == array_index_949021 ? add_967539 : sel_967536;
  assign add_967543 = sel_967540 + 8'h01;
  assign sel_967544 = array_index_967183 == array_index_949027 ? add_967543 : sel_967540;
  assign add_967547 = sel_967544 + 8'h01;
  assign sel_967548 = array_index_967183 == array_index_949033 ? add_967547 : sel_967544;
  assign add_967551 = sel_967548 + 8'h01;
  assign sel_967552 = array_index_967183 == array_index_949039 ? add_967551 : sel_967548;
  assign add_967555 = sel_967552 + 8'h01;
  assign sel_967556 = array_index_967183 == array_index_949045 ? add_967555 : sel_967552;
  assign add_967559 = sel_967556 + 8'h01;
  assign sel_967560 = array_index_967183 == array_index_949051 ? add_967559 : sel_967556;
  assign add_967563 = sel_967560 + 8'h01;
  assign sel_967564 = array_index_967183 == array_index_949057 ? add_967563 : sel_967560;
  assign add_967567 = sel_967564 + 8'h01;
  assign sel_967568 = array_index_967183 == array_index_949063 ? add_967567 : sel_967564;
  assign add_967571 = sel_967568 + 8'h01;
  assign sel_967572 = array_index_967183 == array_index_949069 ? add_967571 : sel_967568;
  assign add_967575 = sel_967572 + 8'h01;
  assign sel_967576 = array_index_967183 == array_index_949075 ? add_967575 : sel_967572;
  assign add_967579 = sel_967576 + 8'h01;
  assign sel_967580 = array_index_967183 == array_index_949081 ? add_967579 : sel_967576;
  assign add_967584 = sel_967580 + 8'h01;
  assign array_index_967585 = set1_unflattened[7'h2f];
  assign sel_967586 = array_index_967183 == array_index_949087 ? add_967584 : sel_967580;
  assign add_967589 = sel_967586 + 8'h01;
  assign sel_967590 = array_index_967585 == array_index_948483 ? add_967589 : sel_967586;
  assign add_967593 = sel_967590 + 8'h01;
  assign sel_967594 = array_index_967585 == array_index_948487 ? add_967593 : sel_967590;
  assign add_967597 = sel_967594 + 8'h01;
  assign sel_967598 = array_index_967585 == array_index_948495 ? add_967597 : sel_967594;
  assign add_967601 = sel_967598 + 8'h01;
  assign sel_967602 = array_index_967585 == array_index_948503 ? add_967601 : sel_967598;
  assign add_967605 = sel_967602 + 8'h01;
  assign sel_967606 = array_index_967585 == array_index_948511 ? add_967605 : sel_967602;
  assign add_967609 = sel_967606 + 8'h01;
  assign sel_967610 = array_index_967585 == array_index_948519 ? add_967609 : sel_967606;
  assign add_967613 = sel_967610 + 8'h01;
  assign sel_967614 = array_index_967585 == array_index_948527 ? add_967613 : sel_967610;
  assign add_967617 = sel_967614 + 8'h01;
  assign sel_967618 = array_index_967585 == array_index_948535 ? add_967617 : sel_967614;
  assign add_967621 = sel_967618 + 8'h01;
  assign sel_967622 = array_index_967585 == array_index_948541 ? add_967621 : sel_967618;
  assign add_967625 = sel_967622 + 8'h01;
  assign sel_967626 = array_index_967585 == array_index_948547 ? add_967625 : sel_967622;
  assign add_967629 = sel_967626 + 8'h01;
  assign sel_967630 = array_index_967585 == array_index_948553 ? add_967629 : sel_967626;
  assign add_967633 = sel_967630 + 8'h01;
  assign sel_967634 = array_index_967585 == array_index_948559 ? add_967633 : sel_967630;
  assign add_967637 = sel_967634 + 8'h01;
  assign sel_967638 = array_index_967585 == array_index_948565 ? add_967637 : sel_967634;
  assign add_967641 = sel_967638 + 8'h01;
  assign sel_967642 = array_index_967585 == array_index_948571 ? add_967641 : sel_967638;
  assign add_967645 = sel_967642 + 8'h01;
  assign sel_967646 = array_index_967585 == array_index_948577 ? add_967645 : sel_967642;
  assign add_967649 = sel_967646 + 8'h01;
  assign sel_967650 = array_index_967585 == array_index_948583 ? add_967649 : sel_967646;
  assign add_967653 = sel_967650 + 8'h01;
  assign sel_967654 = array_index_967585 == array_index_948589 ? add_967653 : sel_967650;
  assign add_967657 = sel_967654 + 8'h01;
  assign sel_967658 = array_index_967585 == array_index_948595 ? add_967657 : sel_967654;
  assign add_967661 = sel_967658 + 8'h01;
  assign sel_967662 = array_index_967585 == array_index_948601 ? add_967661 : sel_967658;
  assign add_967665 = sel_967662 + 8'h01;
  assign sel_967666 = array_index_967585 == array_index_948607 ? add_967665 : sel_967662;
  assign add_967669 = sel_967666 + 8'h01;
  assign sel_967670 = array_index_967585 == array_index_948613 ? add_967669 : sel_967666;
  assign add_967673 = sel_967670 + 8'h01;
  assign sel_967674 = array_index_967585 == array_index_948619 ? add_967673 : sel_967670;
  assign add_967677 = sel_967674 + 8'h01;
  assign sel_967678 = array_index_967585 == array_index_948625 ? add_967677 : sel_967674;
  assign add_967681 = sel_967678 + 8'h01;
  assign sel_967682 = array_index_967585 == array_index_948631 ? add_967681 : sel_967678;
  assign add_967685 = sel_967682 + 8'h01;
  assign sel_967686 = array_index_967585 == array_index_948637 ? add_967685 : sel_967682;
  assign add_967689 = sel_967686 + 8'h01;
  assign sel_967690 = array_index_967585 == array_index_948643 ? add_967689 : sel_967686;
  assign add_967693 = sel_967690 + 8'h01;
  assign sel_967694 = array_index_967585 == array_index_948649 ? add_967693 : sel_967690;
  assign add_967697 = sel_967694 + 8'h01;
  assign sel_967698 = array_index_967585 == array_index_948655 ? add_967697 : sel_967694;
  assign add_967701 = sel_967698 + 8'h01;
  assign sel_967702 = array_index_967585 == array_index_948661 ? add_967701 : sel_967698;
  assign add_967705 = sel_967702 + 8'h01;
  assign sel_967706 = array_index_967585 == array_index_948667 ? add_967705 : sel_967702;
  assign add_967709 = sel_967706 + 8'h01;
  assign sel_967710 = array_index_967585 == array_index_948673 ? add_967709 : sel_967706;
  assign add_967713 = sel_967710 + 8'h01;
  assign sel_967714 = array_index_967585 == array_index_948679 ? add_967713 : sel_967710;
  assign add_967717 = sel_967714 + 8'h01;
  assign sel_967718 = array_index_967585 == array_index_948685 ? add_967717 : sel_967714;
  assign add_967721 = sel_967718 + 8'h01;
  assign sel_967722 = array_index_967585 == array_index_948691 ? add_967721 : sel_967718;
  assign add_967725 = sel_967722 + 8'h01;
  assign sel_967726 = array_index_967585 == array_index_948697 ? add_967725 : sel_967722;
  assign add_967729 = sel_967726 + 8'h01;
  assign sel_967730 = array_index_967585 == array_index_948703 ? add_967729 : sel_967726;
  assign add_967733 = sel_967730 + 8'h01;
  assign sel_967734 = array_index_967585 == array_index_948709 ? add_967733 : sel_967730;
  assign add_967737 = sel_967734 + 8'h01;
  assign sel_967738 = array_index_967585 == array_index_948715 ? add_967737 : sel_967734;
  assign add_967741 = sel_967738 + 8'h01;
  assign sel_967742 = array_index_967585 == array_index_948721 ? add_967741 : sel_967738;
  assign add_967745 = sel_967742 + 8'h01;
  assign sel_967746 = array_index_967585 == array_index_948727 ? add_967745 : sel_967742;
  assign add_967749 = sel_967746 + 8'h01;
  assign sel_967750 = array_index_967585 == array_index_948733 ? add_967749 : sel_967746;
  assign add_967753 = sel_967750 + 8'h01;
  assign sel_967754 = array_index_967585 == array_index_948739 ? add_967753 : sel_967750;
  assign add_967757 = sel_967754 + 8'h01;
  assign sel_967758 = array_index_967585 == array_index_948745 ? add_967757 : sel_967754;
  assign add_967761 = sel_967758 + 8'h01;
  assign sel_967762 = array_index_967585 == array_index_948751 ? add_967761 : sel_967758;
  assign add_967765 = sel_967762 + 8'h01;
  assign sel_967766 = array_index_967585 == array_index_948757 ? add_967765 : sel_967762;
  assign add_967769 = sel_967766 + 8'h01;
  assign sel_967770 = array_index_967585 == array_index_948763 ? add_967769 : sel_967766;
  assign add_967773 = sel_967770 + 8'h01;
  assign sel_967774 = array_index_967585 == array_index_948769 ? add_967773 : sel_967770;
  assign add_967777 = sel_967774 + 8'h01;
  assign sel_967778 = array_index_967585 == array_index_948775 ? add_967777 : sel_967774;
  assign add_967781 = sel_967778 + 8'h01;
  assign sel_967782 = array_index_967585 == array_index_948781 ? add_967781 : sel_967778;
  assign add_967785 = sel_967782 + 8'h01;
  assign sel_967786 = array_index_967585 == array_index_948787 ? add_967785 : sel_967782;
  assign add_967789 = sel_967786 + 8'h01;
  assign sel_967790 = array_index_967585 == array_index_948793 ? add_967789 : sel_967786;
  assign add_967793 = sel_967790 + 8'h01;
  assign sel_967794 = array_index_967585 == array_index_948799 ? add_967793 : sel_967790;
  assign add_967797 = sel_967794 + 8'h01;
  assign sel_967798 = array_index_967585 == array_index_948805 ? add_967797 : sel_967794;
  assign add_967801 = sel_967798 + 8'h01;
  assign sel_967802 = array_index_967585 == array_index_948811 ? add_967801 : sel_967798;
  assign add_967805 = sel_967802 + 8'h01;
  assign sel_967806 = array_index_967585 == array_index_948817 ? add_967805 : sel_967802;
  assign add_967809 = sel_967806 + 8'h01;
  assign sel_967810 = array_index_967585 == array_index_948823 ? add_967809 : sel_967806;
  assign add_967813 = sel_967810 + 8'h01;
  assign sel_967814 = array_index_967585 == array_index_948829 ? add_967813 : sel_967810;
  assign add_967817 = sel_967814 + 8'h01;
  assign sel_967818 = array_index_967585 == array_index_948835 ? add_967817 : sel_967814;
  assign add_967821 = sel_967818 + 8'h01;
  assign sel_967822 = array_index_967585 == array_index_948841 ? add_967821 : sel_967818;
  assign add_967825 = sel_967822 + 8'h01;
  assign sel_967826 = array_index_967585 == array_index_948847 ? add_967825 : sel_967822;
  assign add_967829 = sel_967826 + 8'h01;
  assign sel_967830 = array_index_967585 == array_index_948853 ? add_967829 : sel_967826;
  assign add_967833 = sel_967830 + 8'h01;
  assign sel_967834 = array_index_967585 == array_index_948859 ? add_967833 : sel_967830;
  assign add_967837 = sel_967834 + 8'h01;
  assign sel_967838 = array_index_967585 == array_index_948865 ? add_967837 : sel_967834;
  assign add_967841 = sel_967838 + 8'h01;
  assign sel_967842 = array_index_967585 == array_index_948871 ? add_967841 : sel_967838;
  assign add_967845 = sel_967842 + 8'h01;
  assign sel_967846 = array_index_967585 == array_index_948877 ? add_967845 : sel_967842;
  assign add_967849 = sel_967846 + 8'h01;
  assign sel_967850 = array_index_967585 == array_index_948883 ? add_967849 : sel_967846;
  assign add_967853 = sel_967850 + 8'h01;
  assign sel_967854 = array_index_967585 == array_index_948889 ? add_967853 : sel_967850;
  assign add_967857 = sel_967854 + 8'h01;
  assign sel_967858 = array_index_967585 == array_index_948895 ? add_967857 : sel_967854;
  assign add_967861 = sel_967858 + 8'h01;
  assign sel_967862 = array_index_967585 == array_index_948901 ? add_967861 : sel_967858;
  assign add_967865 = sel_967862 + 8'h01;
  assign sel_967866 = array_index_967585 == array_index_948907 ? add_967865 : sel_967862;
  assign add_967869 = sel_967866 + 8'h01;
  assign sel_967870 = array_index_967585 == array_index_948913 ? add_967869 : sel_967866;
  assign add_967873 = sel_967870 + 8'h01;
  assign sel_967874 = array_index_967585 == array_index_948919 ? add_967873 : sel_967870;
  assign add_967877 = sel_967874 + 8'h01;
  assign sel_967878 = array_index_967585 == array_index_948925 ? add_967877 : sel_967874;
  assign add_967881 = sel_967878 + 8'h01;
  assign sel_967882 = array_index_967585 == array_index_948931 ? add_967881 : sel_967878;
  assign add_967885 = sel_967882 + 8'h01;
  assign sel_967886 = array_index_967585 == array_index_948937 ? add_967885 : sel_967882;
  assign add_967889 = sel_967886 + 8'h01;
  assign sel_967890 = array_index_967585 == array_index_948943 ? add_967889 : sel_967886;
  assign add_967893 = sel_967890 + 8'h01;
  assign sel_967894 = array_index_967585 == array_index_948949 ? add_967893 : sel_967890;
  assign add_967897 = sel_967894 + 8'h01;
  assign sel_967898 = array_index_967585 == array_index_948955 ? add_967897 : sel_967894;
  assign add_967901 = sel_967898 + 8'h01;
  assign sel_967902 = array_index_967585 == array_index_948961 ? add_967901 : sel_967898;
  assign add_967905 = sel_967902 + 8'h01;
  assign sel_967906 = array_index_967585 == array_index_948967 ? add_967905 : sel_967902;
  assign add_967909 = sel_967906 + 8'h01;
  assign sel_967910 = array_index_967585 == array_index_948973 ? add_967909 : sel_967906;
  assign add_967913 = sel_967910 + 8'h01;
  assign sel_967914 = array_index_967585 == array_index_948979 ? add_967913 : sel_967910;
  assign add_967917 = sel_967914 + 8'h01;
  assign sel_967918 = array_index_967585 == array_index_948985 ? add_967917 : sel_967914;
  assign add_967921 = sel_967918 + 8'h01;
  assign sel_967922 = array_index_967585 == array_index_948991 ? add_967921 : sel_967918;
  assign add_967925 = sel_967922 + 8'h01;
  assign sel_967926 = array_index_967585 == array_index_948997 ? add_967925 : sel_967922;
  assign add_967929 = sel_967926 + 8'h01;
  assign sel_967930 = array_index_967585 == array_index_949003 ? add_967929 : sel_967926;
  assign add_967933 = sel_967930 + 8'h01;
  assign sel_967934 = array_index_967585 == array_index_949009 ? add_967933 : sel_967930;
  assign add_967937 = sel_967934 + 8'h01;
  assign sel_967938 = array_index_967585 == array_index_949015 ? add_967937 : sel_967934;
  assign add_967941 = sel_967938 + 8'h01;
  assign sel_967942 = array_index_967585 == array_index_949021 ? add_967941 : sel_967938;
  assign add_967945 = sel_967942 + 8'h01;
  assign sel_967946 = array_index_967585 == array_index_949027 ? add_967945 : sel_967942;
  assign add_967949 = sel_967946 + 8'h01;
  assign sel_967950 = array_index_967585 == array_index_949033 ? add_967949 : sel_967946;
  assign add_967953 = sel_967950 + 8'h01;
  assign sel_967954 = array_index_967585 == array_index_949039 ? add_967953 : sel_967950;
  assign add_967957 = sel_967954 + 8'h01;
  assign sel_967958 = array_index_967585 == array_index_949045 ? add_967957 : sel_967954;
  assign add_967961 = sel_967958 + 8'h01;
  assign sel_967962 = array_index_967585 == array_index_949051 ? add_967961 : sel_967958;
  assign add_967965 = sel_967962 + 8'h01;
  assign sel_967966 = array_index_967585 == array_index_949057 ? add_967965 : sel_967962;
  assign add_967969 = sel_967966 + 8'h01;
  assign sel_967970 = array_index_967585 == array_index_949063 ? add_967969 : sel_967966;
  assign add_967973 = sel_967970 + 8'h01;
  assign sel_967974 = array_index_967585 == array_index_949069 ? add_967973 : sel_967970;
  assign add_967977 = sel_967974 + 8'h01;
  assign sel_967978 = array_index_967585 == array_index_949075 ? add_967977 : sel_967974;
  assign add_967981 = sel_967978 + 8'h01;
  assign sel_967982 = array_index_967585 == array_index_949081 ? add_967981 : sel_967978;
  assign add_967986 = sel_967982 + 8'h01;
  assign array_index_967987 = set1_unflattened[7'h30];
  assign sel_967988 = array_index_967585 == array_index_949087 ? add_967986 : sel_967982;
  assign add_967991 = sel_967988 + 8'h01;
  assign sel_967992 = array_index_967987 == array_index_948483 ? add_967991 : sel_967988;
  assign add_967995 = sel_967992 + 8'h01;
  assign sel_967996 = array_index_967987 == array_index_948487 ? add_967995 : sel_967992;
  assign add_967999 = sel_967996 + 8'h01;
  assign sel_968000 = array_index_967987 == array_index_948495 ? add_967999 : sel_967996;
  assign add_968003 = sel_968000 + 8'h01;
  assign sel_968004 = array_index_967987 == array_index_948503 ? add_968003 : sel_968000;
  assign add_968007 = sel_968004 + 8'h01;
  assign sel_968008 = array_index_967987 == array_index_948511 ? add_968007 : sel_968004;
  assign add_968011 = sel_968008 + 8'h01;
  assign sel_968012 = array_index_967987 == array_index_948519 ? add_968011 : sel_968008;
  assign add_968015 = sel_968012 + 8'h01;
  assign sel_968016 = array_index_967987 == array_index_948527 ? add_968015 : sel_968012;
  assign add_968019 = sel_968016 + 8'h01;
  assign sel_968020 = array_index_967987 == array_index_948535 ? add_968019 : sel_968016;
  assign add_968023 = sel_968020 + 8'h01;
  assign sel_968024 = array_index_967987 == array_index_948541 ? add_968023 : sel_968020;
  assign add_968027 = sel_968024 + 8'h01;
  assign sel_968028 = array_index_967987 == array_index_948547 ? add_968027 : sel_968024;
  assign add_968031 = sel_968028 + 8'h01;
  assign sel_968032 = array_index_967987 == array_index_948553 ? add_968031 : sel_968028;
  assign add_968035 = sel_968032 + 8'h01;
  assign sel_968036 = array_index_967987 == array_index_948559 ? add_968035 : sel_968032;
  assign add_968039 = sel_968036 + 8'h01;
  assign sel_968040 = array_index_967987 == array_index_948565 ? add_968039 : sel_968036;
  assign add_968043 = sel_968040 + 8'h01;
  assign sel_968044 = array_index_967987 == array_index_948571 ? add_968043 : sel_968040;
  assign add_968047 = sel_968044 + 8'h01;
  assign sel_968048 = array_index_967987 == array_index_948577 ? add_968047 : sel_968044;
  assign add_968051 = sel_968048 + 8'h01;
  assign sel_968052 = array_index_967987 == array_index_948583 ? add_968051 : sel_968048;
  assign add_968055 = sel_968052 + 8'h01;
  assign sel_968056 = array_index_967987 == array_index_948589 ? add_968055 : sel_968052;
  assign add_968059 = sel_968056 + 8'h01;
  assign sel_968060 = array_index_967987 == array_index_948595 ? add_968059 : sel_968056;
  assign add_968063 = sel_968060 + 8'h01;
  assign sel_968064 = array_index_967987 == array_index_948601 ? add_968063 : sel_968060;
  assign add_968067 = sel_968064 + 8'h01;
  assign sel_968068 = array_index_967987 == array_index_948607 ? add_968067 : sel_968064;
  assign add_968071 = sel_968068 + 8'h01;
  assign sel_968072 = array_index_967987 == array_index_948613 ? add_968071 : sel_968068;
  assign add_968075 = sel_968072 + 8'h01;
  assign sel_968076 = array_index_967987 == array_index_948619 ? add_968075 : sel_968072;
  assign add_968079 = sel_968076 + 8'h01;
  assign sel_968080 = array_index_967987 == array_index_948625 ? add_968079 : sel_968076;
  assign add_968083 = sel_968080 + 8'h01;
  assign sel_968084 = array_index_967987 == array_index_948631 ? add_968083 : sel_968080;
  assign add_968087 = sel_968084 + 8'h01;
  assign sel_968088 = array_index_967987 == array_index_948637 ? add_968087 : sel_968084;
  assign add_968091 = sel_968088 + 8'h01;
  assign sel_968092 = array_index_967987 == array_index_948643 ? add_968091 : sel_968088;
  assign add_968095 = sel_968092 + 8'h01;
  assign sel_968096 = array_index_967987 == array_index_948649 ? add_968095 : sel_968092;
  assign add_968099 = sel_968096 + 8'h01;
  assign sel_968100 = array_index_967987 == array_index_948655 ? add_968099 : sel_968096;
  assign add_968103 = sel_968100 + 8'h01;
  assign sel_968104 = array_index_967987 == array_index_948661 ? add_968103 : sel_968100;
  assign add_968107 = sel_968104 + 8'h01;
  assign sel_968108 = array_index_967987 == array_index_948667 ? add_968107 : sel_968104;
  assign add_968111 = sel_968108 + 8'h01;
  assign sel_968112 = array_index_967987 == array_index_948673 ? add_968111 : sel_968108;
  assign add_968115 = sel_968112 + 8'h01;
  assign sel_968116 = array_index_967987 == array_index_948679 ? add_968115 : sel_968112;
  assign add_968119 = sel_968116 + 8'h01;
  assign sel_968120 = array_index_967987 == array_index_948685 ? add_968119 : sel_968116;
  assign add_968123 = sel_968120 + 8'h01;
  assign sel_968124 = array_index_967987 == array_index_948691 ? add_968123 : sel_968120;
  assign add_968127 = sel_968124 + 8'h01;
  assign sel_968128 = array_index_967987 == array_index_948697 ? add_968127 : sel_968124;
  assign add_968131 = sel_968128 + 8'h01;
  assign sel_968132 = array_index_967987 == array_index_948703 ? add_968131 : sel_968128;
  assign add_968135 = sel_968132 + 8'h01;
  assign sel_968136 = array_index_967987 == array_index_948709 ? add_968135 : sel_968132;
  assign add_968139 = sel_968136 + 8'h01;
  assign sel_968140 = array_index_967987 == array_index_948715 ? add_968139 : sel_968136;
  assign add_968143 = sel_968140 + 8'h01;
  assign sel_968144 = array_index_967987 == array_index_948721 ? add_968143 : sel_968140;
  assign add_968147 = sel_968144 + 8'h01;
  assign sel_968148 = array_index_967987 == array_index_948727 ? add_968147 : sel_968144;
  assign add_968151 = sel_968148 + 8'h01;
  assign sel_968152 = array_index_967987 == array_index_948733 ? add_968151 : sel_968148;
  assign add_968155 = sel_968152 + 8'h01;
  assign sel_968156 = array_index_967987 == array_index_948739 ? add_968155 : sel_968152;
  assign add_968159 = sel_968156 + 8'h01;
  assign sel_968160 = array_index_967987 == array_index_948745 ? add_968159 : sel_968156;
  assign add_968163 = sel_968160 + 8'h01;
  assign sel_968164 = array_index_967987 == array_index_948751 ? add_968163 : sel_968160;
  assign add_968167 = sel_968164 + 8'h01;
  assign sel_968168 = array_index_967987 == array_index_948757 ? add_968167 : sel_968164;
  assign add_968171 = sel_968168 + 8'h01;
  assign sel_968172 = array_index_967987 == array_index_948763 ? add_968171 : sel_968168;
  assign add_968175 = sel_968172 + 8'h01;
  assign sel_968176 = array_index_967987 == array_index_948769 ? add_968175 : sel_968172;
  assign add_968179 = sel_968176 + 8'h01;
  assign sel_968180 = array_index_967987 == array_index_948775 ? add_968179 : sel_968176;
  assign add_968183 = sel_968180 + 8'h01;
  assign sel_968184 = array_index_967987 == array_index_948781 ? add_968183 : sel_968180;
  assign add_968187 = sel_968184 + 8'h01;
  assign sel_968188 = array_index_967987 == array_index_948787 ? add_968187 : sel_968184;
  assign add_968191 = sel_968188 + 8'h01;
  assign sel_968192 = array_index_967987 == array_index_948793 ? add_968191 : sel_968188;
  assign add_968195 = sel_968192 + 8'h01;
  assign sel_968196 = array_index_967987 == array_index_948799 ? add_968195 : sel_968192;
  assign add_968199 = sel_968196 + 8'h01;
  assign sel_968200 = array_index_967987 == array_index_948805 ? add_968199 : sel_968196;
  assign add_968203 = sel_968200 + 8'h01;
  assign sel_968204 = array_index_967987 == array_index_948811 ? add_968203 : sel_968200;
  assign add_968207 = sel_968204 + 8'h01;
  assign sel_968208 = array_index_967987 == array_index_948817 ? add_968207 : sel_968204;
  assign add_968211 = sel_968208 + 8'h01;
  assign sel_968212 = array_index_967987 == array_index_948823 ? add_968211 : sel_968208;
  assign add_968215 = sel_968212 + 8'h01;
  assign sel_968216 = array_index_967987 == array_index_948829 ? add_968215 : sel_968212;
  assign add_968219 = sel_968216 + 8'h01;
  assign sel_968220 = array_index_967987 == array_index_948835 ? add_968219 : sel_968216;
  assign add_968223 = sel_968220 + 8'h01;
  assign sel_968224 = array_index_967987 == array_index_948841 ? add_968223 : sel_968220;
  assign add_968227 = sel_968224 + 8'h01;
  assign sel_968228 = array_index_967987 == array_index_948847 ? add_968227 : sel_968224;
  assign add_968231 = sel_968228 + 8'h01;
  assign sel_968232 = array_index_967987 == array_index_948853 ? add_968231 : sel_968228;
  assign add_968235 = sel_968232 + 8'h01;
  assign sel_968236 = array_index_967987 == array_index_948859 ? add_968235 : sel_968232;
  assign add_968239 = sel_968236 + 8'h01;
  assign sel_968240 = array_index_967987 == array_index_948865 ? add_968239 : sel_968236;
  assign add_968243 = sel_968240 + 8'h01;
  assign sel_968244 = array_index_967987 == array_index_948871 ? add_968243 : sel_968240;
  assign add_968247 = sel_968244 + 8'h01;
  assign sel_968248 = array_index_967987 == array_index_948877 ? add_968247 : sel_968244;
  assign add_968251 = sel_968248 + 8'h01;
  assign sel_968252 = array_index_967987 == array_index_948883 ? add_968251 : sel_968248;
  assign add_968255 = sel_968252 + 8'h01;
  assign sel_968256 = array_index_967987 == array_index_948889 ? add_968255 : sel_968252;
  assign add_968259 = sel_968256 + 8'h01;
  assign sel_968260 = array_index_967987 == array_index_948895 ? add_968259 : sel_968256;
  assign add_968263 = sel_968260 + 8'h01;
  assign sel_968264 = array_index_967987 == array_index_948901 ? add_968263 : sel_968260;
  assign add_968267 = sel_968264 + 8'h01;
  assign sel_968268 = array_index_967987 == array_index_948907 ? add_968267 : sel_968264;
  assign add_968271 = sel_968268 + 8'h01;
  assign sel_968272 = array_index_967987 == array_index_948913 ? add_968271 : sel_968268;
  assign add_968275 = sel_968272 + 8'h01;
  assign sel_968276 = array_index_967987 == array_index_948919 ? add_968275 : sel_968272;
  assign add_968279 = sel_968276 + 8'h01;
  assign sel_968280 = array_index_967987 == array_index_948925 ? add_968279 : sel_968276;
  assign add_968283 = sel_968280 + 8'h01;
  assign sel_968284 = array_index_967987 == array_index_948931 ? add_968283 : sel_968280;
  assign add_968287 = sel_968284 + 8'h01;
  assign sel_968288 = array_index_967987 == array_index_948937 ? add_968287 : sel_968284;
  assign add_968291 = sel_968288 + 8'h01;
  assign sel_968292 = array_index_967987 == array_index_948943 ? add_968291 : sel_968288;
  assign add_968295 = sel_968292 + 8'h01;
  assign sel_968296 = array_index_967987 == array_index_948949 ? add_968295 : sel_968292;
  assign add_968299 = sel_968296 + 8'h01;
  assign sel_968300 = array_index_967987 == array_index_948955 ? add_968299 : sel_968296;
  assign add_968303 = sel_968300 + 8'h01;
  assign sel_968304 = array_index_967987 == array_index_948961 ? add_968303 : sel_968300;
  assign add_968307 = sel_968304 + 8'h01;
  assign sel_968308 = array_index_967987 == array_index_948967 ? add_968307 : sel_968304;
  assign add_968311 = sel_968308 + 8'h01;
  assign sel_968312 = array_index_967987 == array_index_948973 ? add_968311 : sel_968308;
  assign add_968315 = sel_968312 + 8'h01;
  assign sel_968316 = array_index_967987 == array_index_948979 ? add_968315 : sel_968312;
  assign add_968319 = sel_968316 + 8'h01;
  assign sel_968320 = array_index_967987 == array_index_948985 ? add_968319 : sel_968316;
  assign add_968323 = sel_968320 + 8'h01;
  assign sel_968324 = array_index_967987 == array_index_948991 ? add_968323 : sel_968320;
  assign add_968327 = sel_968324 + 8'h01;
  assign sel_968328 = array_index_967987 == array_index_948997 ? add_968327 : sel_968324;
  assign add_968331 = sel_968328 + 8'h01;
  assign sel_968332 = array_index_967987 == array_index_949003 ? add_968331 : sel_968328;
  assign add_968335 = sel_968332 + 8'h01;
  assign sel_968336 = array_index_967987 == array_index_949009 ? add_968335 : sel_968332;
  assign add_968339 = sel_968336 + 8'h01;
  assign sel_968340 = array_index_967987 == array_index_949015 ? add_968339 : sel_968336;
  assign add_968343 = sel_968340 + 8'h01;
  assign sel_968344 = array_index_967987 == array_index_949021 ? add_968343 : sel_968340;
  assign add_968347 = sel_968344 + 8'h01;
  assign sel_968348 = array_index_967987 == array_index_949027 ? add_968347 : sel_968344;
  assign add_968351 = sel_968348 + 8'h01;
  assign sel_968352 = array_index_967987 == array_index_949033 ? add_968351 : sel_968348;
  assign add_968355 = sel_968352 + 8'h01;
  assign sel_968356 = array_index_967987 == array_index_949039 ? add_968355 : sel_968352;
  assign add_968359 = sel_968356 + 8'h01;
  assign sel_968360 = array_index_967987 == array_index_949045 ? add_968359 : sel_968356;
  assign add_968363 = sel_968360 + 8'h01;
  assign sel_968364 = array_index_967987 == array_index_949051 ? add_968363 : sel_968360;
  assign add_968367 = sel_968364 + 8'h01;
  assign sel_968368 = array_index_967987 == array_index_949057 ? add_968367 : sel_968364;
  assign add_968371 = sel_968368 + 8'h01;
  assign sel_968372 = array_index_967987 == array_index_949063 ? add_968371 : sel_968368;
  assign add_968375 = sel_968372 + 8'h01;
  assign sel_968376 = array_index_967987 == array_index_949069 ? add_968375 : sel_968372;
  assign add_968379 = sel_968376 + 8'h01;
  assign sel_968380 = array_index_967987 == array_index_949075 ? add_968379 : sel_968376;
  assign add_968383 = sel_968380 + 8'h01;
  assign sel_968384 = array_index_967987 == array_index_949081 ? add_968383 : sel_968380;
  assign add_968388 = sel_968384 + 8'h01;
  assign array_index_968389 = set1_unflattened[7'h31];
  assign sel_968390 = array_index_967987 == array_index_949087 ? add_968388 : sel_968384;
  assign add_968393 = sel_968390 + 8'h01;
  assign sel_968394 = array_index_968389 == array_index_948483 ? add_968393 : sel_968390;
  assign add_968397 = sel_968394 + 8'h01;
  assign sel_968398 = array_index_968389 == array_index_948487 ? add_968397 : sel_968394;
  assign add_968401 = sel_968398 + 8'h01;
  assign sel_968402 = array_index_968389 == array_index_948495 ? add_968401 : sel_968398;
  assign add_968405 = sel_968402 + 8'h01;
  assign sel_968406 = array_index_968389 == array_index_948503 ? add_968405 : sel_968402;
  assign add_968409 = sel_968406 + 8'h01;
  assign sel_968410 = array_index_968389 == array_index_948511 ? add_968409 : sel_968406;
  assign add_968413 = sel_968410 + 8'h01;
  assign sel_968414 = array_index_968389 == array_index_948519 ? add_968413 : sel_968410;
  assign add_968417 = sel_968414 + 8'h01;
  assign sel_968418 = array_index_968389 == array_index_948527 ? add_968417 : sel_968414;
  assign add_968421 = sel_968418 + 8'h01;
  assign sel_968422 = array_index_968389 == array_index_948535 ? add_968421 : sel_968418;
  assign add_968425 = sel_968422 + 8'h01;
  assign sel_968426 = array_index_968389 == array_index_948541 ? add_968425 : sel_968422;
  assign add_968429 = sel_968426 + 8'h01;
  assign sel_968430 = array_index_968389 == array_index_948547 ? add_968429 : sel_968426;
  assign add_968433 = sel_968430 + 8'h01;
  assign sel_968434 = array_index_968389 == array_index_948553 ? add_968433 : sel_968430;
  assign add_968437 = sel_968434 + 8'h01;
  assign sel_968438 = array_index_968389 == array_index_948559 ? add_968437 : sel_968434;
  assign add_968441 = sel_968438 + 8'h01;
  assign sel_968442 = array_index_968389 == array_index_948565 ? add_968441 : sel_968438;
  assign add_968445 = sel_968442 + 8'h01;
  assign sel_968446 = array_index_968389 == array_index_948571 ? add_968445 : sel_968442;
  assign add_968449 = sel_968446 + 8'h01;
  assign sel_968450 = array_index_968389 == array_index_948577 ? add_968449 : sel_968446;
  assign add_968453 = sel_968450 + 8'h01;
  assign sel_968454 = array_index_968389 == array_index_948583 ? add_968453 : sel_968450;
  assign add_968457 = sel_968454 + 8'h01;
  assign sel_968458 = array_index_968389 == array_index_948589 ? add_968457 : sel_968454;
  assign add_968461 = sel_968458 + 8'h01;
  assign sel_968462 = array_index_968389 == array_index_948595 ? add_968461 : sel_968458;
  assign add_968465 = sel_968462 + 8'h01;
  assign sel_968466 = array_index_968389 == array_index_948601 ? add_968465 : sel_968462;
  assign add_968469 = sel_968466 + 8'h01;
  assign sel_968470 = array_index_968389 == array_index_948607 ? add_968469 : sel_968466;
  assign add_968473 = sel_968470 + 8'h01;
  assign sel_968474 = array_index_968389 == array_index_948613 ? add_968473 : sel_968470;
  assign add_968477 = sel_968474 + 8'h01;
  assign sel_968478 = array_index_968389 == array_index_948619 ? add_968477 : sel_968474;
  assign add_968481 = sel_968478 + 8'h01;
  assign sel_968482 = array_index_968389 == array_index_948625 ? add_968481 : sel_968478;
  assign add_968485 = sel_968482 + 8'h01;
  assign sel_968486 = array_index_968389 == array_index_948631 ? add_968485 : sel_968482;
  assign add_968489 = sel_968486 + 8'h01;
  assign sel_968490 = array_index_968389 == array_index_948637 ? add_968489 : sel_968486;
  assign add_968493 = sel_968490 + 8'h01;
  assign sel_968494 = array_index_968389 == array_index_948643 ? add_968493 : sel_968490;
  assign add_968497 = sel_968494 + 8'h01;
  assign sel_968498 = array_index_968389 == array_index_948649 ? add_968497 : sel_968494;
  assign add_968501 = sel_968498 + 8'h01;
  assign sel_968502 = array_index_968389 == array_index_948655 ? add_968501 : sel_968498;
  assign add_968505 = sel_968502 + 8'h01;
  assign sel_968506 = array_index_968389 == array_index_948661 ? add_968505 : sel_968502;
  assign add_968509 = sel_968506 + 8'h01;
  assign sel_968510 = array_index_968389 == array_index_948667 ? add_968509 : sel_968506;
  assign add_968513 = sel_968510 + 8'h01;
  assign sel_968514 = array_index_968389 == array_index_948673 ? add_968513 : sel_968510;
  assign add_968517 = sel_968514 + 8'h01;
  assign sel_968518 = array_index_968389 == array_index_948679 ? add_968517 : sel_968514;
  assign add_968521 = sel_968518 + 8'h01;
  assign sel_968522 = array_index_968389 == array_index_948685 ? add_968521 : sel_968518;
  assign add_968525 = sel_968522 + 8'h01;
  assign sel_968526 = array_index_968389 == array_index_948691 ? add_968525 : sel_968522;
  assign add_968529 = sel_968526 + 8'h01;
  assign sel_968530 = array_index_968389 == array_index_948697 ? add_968529 : sel_968526;
  assign add_968533 = sel_968530 + 8'h01;
  assign sel_968534 = array_index_968389 == array_index_948703 ? add_968533 : sel_968530;
  assign add_968537 = sel_968534 + 8'h01;
  assign sel_968538 = array_index_968389 == array_index_948709 ? add_968537 : sel_968534;
  assign add_968541 = sel_968538 + 8'h01;
  assign sel_968542 = array_index_968389 == array_index_948715 ? add_968541 : sel_968538;
  assign add_968545 = sel_968542 + 8'h01;
  assign sel_968546 = array_index_968389 == array_index_948721 ? add_968545 : sel_968542;
  assign add_968549 = sel_968546 + 8'h01;
  assign sel_968550 = array_index_968389 == array_index_948727 ? add_968549 : sel_968546;
  assign add_968553 = sel_968550 + 8'h01;
  assign sel_968554 = array_index_968389 == array_index_948733 ? add_968553 : sel_968550;
  assign add_968557 = sel_968554 + 8'h01;
  assign sel_968558 = array_index_968389 == array_index_948739 ? add_968557 : sel_968554;
  assign add_968561 = sel_968558 + 8'h01;
  assign sel_968562 = array_index_968389 == array_index_948745 ? add_968561 : sel_968558;
  assign add_968565 = sel_968562 + 8'h01;
  assign sel_968566 = array_index_968389 == array_index_948751 ? add_968565 : sel_968562;
  assign add_968569 = sel_968566 + 8'h01;
  assign sel_968570 = array_index_968389 == array_index_948757 ? add_968569 : sel_968566;
  assign add_968573 = sel_968570 + 8'h01;
  assign sel_968574 = array_index_968389 == array_index_948763 ? add_968573 : sel_968570;
  assign add_968577 = sel_968574 + 8'h01;
  assign sel_968578 = array_index_968389 == array_index_948769 ? add_968577 : sel_968574;
  assign add_968581 = sel_968578 + 8'h01;
  assign sel_968582 = array_index_968389 == array_index_948775 ? add_968581 : sel_968578;
  assign add_968585 = sel_968582 + 8'h01;
  assign sel_968586 = array_index_968389 == array_index_948781 ? add_968585 : sel_968582;
  assign add_968589 = sel_968586 + 8'h01;
  assign sel_968590 = array_index_968389 == array_index_948787 ? add_968589 : sel_968586;
  assign add_968593 = sel_968590 + 8'h01;
  assign sel_968594 = array_index_968389 == array_index_948793 ? add_968593 : sel_968590;
  assign add_968597 = sel_968594 + 8'h01;
  assign sel_968598 = array_index_968389 == array_index_948799 ? add_968597 : sel_968594;
  assign add_968601 = sel_968598 + 8'h01;
  assign sel_968602 = array_index_968389 == array_index_948805 ? add_968601 : sel_968598;
  assign add_968605 = sel_968602 + 8'h01;
  assign sel_968606 = array_index_968389 == array_index_948811 ? add_968605 : sel_968602;
  assign add_968609 = sel_968606 + 8'h01;
  assign sel_968610 = array_index_968389 == array_index_948817 ? add_968609 : sel_968606;
  assign add_968613 = sel_968610 + 8'h01;
  assign sel_968614 = array_index_968389 == array_index_948823 ? add_968613 : sel_968610;
  assign add_968617 = sel_968614 + 8'h01;
  assign sel_968618 = array_index_968389 == array_index_948829 ? add_968617 : sel_968614;
  assign add_968621 = sel_968618 + 8'h01;
  assign sel_968622 = array_index_968389 == array_index_948835 ? add_968621 : sel_968618;
  assign add_968625 = sel_968622 + 8'h01;
  assign sel_968626 = array_index_968389 == array_index_948841 ? add_968625 : sel_968622;
  assign add_968629 = sel_968626 + 8'h01;
  assign sel_968630 = array_index_968389 == array_index_948847 ? add_968629 : sel_968626;
  assign add_968633 = sel_968630 + 8'h01;
  assign sel_968634 = array_index_968389 == array_index_948853 ? add_968633 : sel_968630;
  assign add_968637 = sel_968634 + 8'h01;
  assign sel_968638 = array_index_968389 == array_index_948859 ? add_968637 : sel_968634;
  assign add_968641 = sel_968638 + 8'h01;
  assign sel_968642 = array_index_968389 == array_index_948865 ? add_968641 : sel_968638;
  assign add_968645 = sel_968642 + 8'h01;
  assign sel_968646 = array_index_968389 == array_index_948871 ? add_968645 : sel_968642;
  assign add_968649 = sel_968646 + 8'h01;
  assign sel_968650 = array_index_968389 == array_index_948877 ? add_968649 : sel_968646;
  assign add_968653 = sel_968650 + 8'h01;
  assign sel_968654 = array_index_968389 == array_index_948883 ? add_968653 : sel_968650;
  assign add_968657 = sel_968654 + 8'h01;
  assign sel_968658 = array_index_968389 == array_index_948889 ? add_968657 : sel_968654;
  assign add_968661 = sel_968658 + 8'h01;
  assign sel_968662 = array_index_968389 == array_index_948895 ? add_968661 : sel_968658;
  assign add_968665 = sel_968662 + 8'h01;
  assign sel_968666 = array_index_968389 == array_index_948901 ? add_968665 : sel_968662;
  assign add_968669 = sel_968666 + 8'h01;
  assign sel_968670 = array_index_968389 == array_index_948907 ? add_968669 : sel_968666;
  assign add_968673 = sel_968670 + 8'h01;
  assign sel_968674 = array_index_968389 == array_index_948913 ? add_968673 : sel_968670;
  assign add_968677 = sel_968674 + 8'h01;
  assign sel_968678 = array_index_968389 == array_index_948919 ? add_968677 : sel_968674;
  assign add_968681 = sel_968678 + 8'h01;
  assign sel_968682 = array_index_968389 == array_index_948925 ? add_968681 : sel_968678;
  assign add_968685 = sel_968682 + 8'h01;
  assign sel_968686 = array_index_968389 == array_index_948931 ? add_968685 : sel_968682;
  assign add_968689 = sel_968686 + 8'h01;
  assign sel_968690 = array_index_968389 == array_index_948937 ? add_968689 : sel_968686;
  assign add_968693 = sel_968690 + 8'h01;
  assign sel_968694 = array_index_968389 == array_index_948943 ? add_968693 : sel_968690;
  assign add_968697 = sel_968694 + 8'h01;
  assign sel_968698 = array_index_968389 == array_index_948949 ? add_968697 : sel_968694;
  assign add_968701 = sel_968698 + 8'h01;
  assign sel_968702 = array_index_968389 == array_index_948955 ? add_968701 : sel_968698;
  assign add_968705 = sel_968702 + 8'h01;
  assign sel_968706 = array_index_968389 == array_index_948961 ? add_968705 : sel_968702;
  assign add_968709 = sel_968706 + 8'h01;
  assign sel_968710 = array_index_968389 == array_index_948967 ? add_968709 : sel_968706;
  assign add_968713 = sel_968710 + 8'h01;
  assign sel_968714 = array_index_968389 == array_index_948973 ? add_968713 : sel_968710;
  assign add_968717 = sel_968714 + 8'h01;
  assign sel_968718 = array_index_968389 == array_index_948979 ? add_968717 : sel_968714;
  assign add_968721 = sel_968718 + 8'h01;
  assign sel_968722 = array_index_968389 == array_index_948985 ? add_968721 : sel_968718;
  assign add_968725 = sel_968722 + 8'h01;
  assign sel_968726 = array_index_968389 == array_index_948991 ? add_968725 : sel_968722;
  assign add_968729 = sel_968726 + 8'h01;
  assign sel_968730 = array_index_968389 == array_index_948997 ? add_968729 : sel_968726;
  assign add_968733 = sel_968730 + 8'h01;
  assign sel_968734 = array_index_968389 == array_index_949003 ? add_968733 : sel_968730;
  assign add_968737 = sel_968734 + 8'h01;
  assign sel_968738 = array_index_968389 == array_index_949009 ? add_968737 : sel_968734;
  assign add_968741 = sel_968738 + 8'h01;
  assign sel_968742 = array_index_968389 == array_index_949015 ? add_968741 : sel_968738;
  assign add_968745 = sel_968742 + 8'h01;
  assign sel_968746 = array_index_968389 == array_index_949021 ? add_968745 : sel_968742;
  assign add_968749 = sel_968746 + 8'h01;
  assign sel_968750 = array_index_968389 == array_index_949027 ? add_968749 : sel_968746;
  assign add_968753 = sel_968750 + 8'h01;
  assign sel_968754 = array_index_968389 == array_index_949033 ? add_968753 : sel_968750;
  assign add_968757 = sel_968754 + 8'h01;
  assign sel_968758 = array_index_968389 == array_index_949039 ? add_968757 : sel_968754;
  assign add_968761 = sel_968758 + 8'h01;
  assign sel_968762 = array_index_968389 == array_index_949045 ? add_968761 : sel_968758;
  assign add_968765 = sel_968762 + 8'h01;
  assign sel_968766 = array_index_968389 == array_index_949051 ? add_968765 : sel_968762;
  assign add_968769 = sel_968766 + 8'h01;
  assign sel_968770 = array_index_968389 == array_index_949057 ? add_968769 : sel_968766;
  assign add_968773 = sel_968770 + 8'h01;
  assign sel_968774 = array_index_968389 == array_index_949063 ? add_968773 : sel_968770;
  assign add_968777 = sel_968774 + 8'h01;
  assign sel_968778 = array_index_968389 == array_index_949069 ? add_968777 : sel_968774;
  assign add_968781 = sel_968778 + 8'h01;
  assign sel_968782 = array_index_968389 == array_index_949075 ? add_968781 : sel_968778;
  assign add_968785 = sel_968782 + 8'h01;
  assign sel_968786 = array_index_968389 == array_index_949081 ? add_968785 : sel_968782;
  assign add_968790 = sel_968786 + 8'h01;
  assign array_index_968791 = set1_unflattened[7'h32];
  assign sel_968792 = array_index_968389 == array_index_949087 ? add_968790 : sel_968786;
  assign add_968795 = sel_968792 + 8'h01;
  assign sel_968796 = array_index_968791 == array_index_948483 ? add_968795 : sel_968792;
  assign add_968799 = sel_968796 + 8'h01;
  assign sel_968800 = array_index_968791 == array_index_948487 ? add_968799 : sel_968796;
  assign add_968803 = sel_968800 + 8'h01;
  assign sel_968804 = array_index_968791 == array_index_948495 ? add_968803 : sel_968800;
  assign add_968807 = sel_968804 + 8'h01;
  assign sel_968808 = array_index_968791 == array_index_948503 ? add_968807 : sel_968804;
  assign add_968811 = sel_968808 + 8'h01;
  assign sel_968812 = array_index_968791 == array_index_948511 ? add_968811 : sel_968808;
  assign add_968815 = sel_968812 + 8'h01;
  assign sel_968816 = array_index_968791 == array_index_948519 ? add_968815 : sel_968812;
  assign add_968819 = sel_968816 + 8'h01;
  assign sel_968820 = array_index_968791 == array_index_948527 ? add_968819 : sel_968816;
  assign add_968823 = sel_968820 + 8'h01;
  assign sel_968824 = array_index_968791 == array_index_948535 ? add_968823 : sel_968820;
  assign add_968827 = sel_968824 + 8'h01;
  assign sel_968828 = array_index_968791 == array_index_948541 ? add_968827 : sel_968824;
  assign add_968831 = sel_968828 + 8'h01;
  assign sel_968832 = array_index_968791 == array_index_948547 ? add_968831 : sel_968828;
  assign add_968835 = sel_968832 + 8'h01;
  assign sel_968836 = array_index_968791 == array_index_948553 ? add_968835 : sel_968832;
  assign add_968839 = sel_968836 + 8'h01;
  assign sel_968840 = array_index_968791 == array_index_948559 ? add_968839 : sel_968836;
  assign add_968843 = sel_968840 + 8'h01;
  assign sel_968844 = array_index_968791 == array_index_948565 ? add_968843 : sel_968840;
  assign add_968847 = sel_968844 + 8'h01;
  assign sel_968848 = array_index_968791 == array_index_948571 ? add_968847 : sel_968844;
  assign add_968851 = sel_968848 + 8'h01;
  assign sel_968852 = array_index_968791 == array_index_948577 ? add_968851 : sel_968848;
  assign add_968855 = sel_968852 + 8'h01;
  assign sel_968856 = array_index_968791 == array_index_948583 ? add_968855 : sel_968852;
  assign add_968859 = sel_968856 + 8'h01;
  assign sel_968860 = array_index_968791 == array_index_948589 ? add_968859 : sel_968856;
  assign add_968863 = sel_968860 + 8'h01;
  assign sel_968864 = array_index_968791 == array_index_948595 ? add_968863 : sel_968860;
  assign add_968867 = sel_968864 + 8'h01;
  assign sel_968868 = array_index_968791 == array_index_948601 ? add_968867 : sel_968864;
  assign add_968871 = sel_968868 + 8'h01;
  assign sel_968872 = array_index_968791 == array_index_948607 ? add_968871 : sel_968868;
  assign add_968875 = sel_968872 + 8'h01;
  assign sel_968876 = array_index_968791 == array_index_948613 ? add_968875 : sel_968872;
  assign add_968879 = sel_968876 + 8'h01;
  assign sel_968880 = array_index_968791 == array_index_948619 ? add_968879 : sel_968876;
  assign add_968883 = sel_968880 + 8'h01;
  assign sel_968884 = array_index_968791 == array_index_948625 ? add_968883 : sel_968880;
  assign add_968887 = sel_968884 + 8'h01;
  assign sel_968888 = array_index_968791 == array_index_948631 ? add_968887 : sel_968884;
  assign add_968891 = sel_968888 + 8'h01;
  assign sel_968892 = array_index_968791 == array_index_948637 ? add_968891 : sel_968888;
  assign add_968895 = sel_968892 + 8'h01;
  assign sel_968896 = array_index_968791 == array_index_948643 ? add_968895 : sel_968892;
  assign add_968899 = sel_968896 + 8'h01;
  assign sel_968900 = array_index_968791 == array_index_948649 ? add_968899 : sel_968896;
  assign add_968903 = sel_968900 + 8'h01;
  assign sel_968904 = array_index_968791 == array_index_948655 ? add_968903 : sel_968900;
  assign add_968907 = sel_968904 + 8'h01;
  assign sel_968908 = array_index_968791 == array_index_948661 ? add_968907 : sel_968904;
  assign add_968911 = sel_968908 + 8'h01;
  assign sel_968912 = array_index_968791 == array_index_948667 ? add_968911 : sel_968908;
  assign add_968915 = sel_968912 + 8'h01;
  assign sel_968916 = array_index_968791 == array_index_948673 ? add_968915 : sel_968912;
  assign add_968919 = sel_968916 + 8'h01;
  assign sel_968920 = array_index_968791 == array_index_948679 ? add_968919 : sel_968916;
  assign add_968923 = sel_968920 + 8'h01;
  assign sel_968924 = array_index_968791 == array_index_948685 ? add_968923 : sel_968920;
  assign add_968927 = sel_968924 + 8'h01;
  assign sel_968928 = array_index_968791 == array_index_948691 ? add_968927 : sel_968924;
  assign add_968931 = sel_968928 + 8'h01;
  assign sel_968932 = array_index_968791 == array_index_948697 ? add_968931 : sel_968928;
  assign add_968935 = sel_968932 + 8'h01;
  assign sel_968936 = array_index_968791 == array_index_948703 ? add_968935 : sel_968932;
  assign add_968939 = sel_968936 + 8'h01;
  assign sel_968940 = array_index_968791 == array_index_948709 ? add_968939 : sel_968936;
  assign add_968943 = sel_968940 + 8'h01;
  assign sel_968944 = array_index_968791 == array_index_948715 ? add_968943 : sel_968940;
  assign add_968947 = sel_968944 + 8'h01;
  assign sel_968948 = array_index_968791 == array_index_948721 ? add_968947 : sel_968944;
  assign add_968951 = sel_968948 + 8'h01;
  assign sel_968952 = array_index_968791 == array_index_948727 ? add_968951 : sel_968948;
  assign add_968955 = sel_968952 + 8'h01;
  assign sel_968956 = array_index_968791 == array_index_948733 ? add_968955 : sel_968952;
  assign add_968959 = sel_968956 + 8'h01;
  assign sel_968960 = array_index_968791 == array_index_948739 ? add_968959 : sel_968956;
  assign add_968963 = sel_968960 + 8'h01;
  assign sel_968964 = array_index_968791 == array_index_948745 ? add_968963 : sel_968960;
  assign add_968967 = sel_968964 + 8'h01;
  assign sel_968968 = array_index_968791 == array_index_948751 ? add_968967 : sel_968964;
  assign add_968971 = sel_968968 + 8'h01;
  assign sel_968972 = array_index_968791 == array_index_948757 ? add_968971 : sel_968968;
  assign add_968975 = sel_968972 + 8'h01;
  assign sel_968976 = array_index_968791 == array_index_948763 ? add_968975 : sel_968972;
  assign add_968979 = sel_968976 + 8'h01;
  assign sel_968980 = array_index_968791 == array_index_948769 ? add_968979 : sel_968976;
  assign add_968983 = sel_968980 + 8'h01;
  assign sel_968984 = array_index_968791 == array_index_948775 ? add_968983 : sel_968980;
  assign add_968987 = sel_968984 + 8'h01;
  assign sel_968988 = array_index_968791 == array_index_948781 ? add_968987 : sel_968984;
  assign add_968991 = sel_968988 + 8'h01;
  assign sel_968992 = array_index_968791 == array_index_948787 ? add_968991 : sel_968988;
  assign add_968995 = sel_968992 + 8'h01;
  assign sel_968996 = array_index_968791 == array_index_948793 ? add_968995 : sel_968992;
  assign add_968999 = sel_968996 + 8'h01;
  assign sel_969000 = array_index_968791 == array_index_948799 ? add_968999 : sel_968996;
  assign add_969003 = sel_969000 + 8'h01;
  assign sel_969004 = array_index_968791 == array_index_948805 ? add_969003 : sel_969000;
  assign add_969007 = sel_969004 + 8'h01;
  assign sel_969008 = array_index_968791 == array_index_948811 ? add_969007 : sel_969004;
  assign add_969011 = sel_969008 + 8'h01;
  assign sel_969012 = array_index_968791 == array_index_948817 ? add_969011 : sel_969008;
  assign add_969015 = sel_969012 + 8'h01;
  assign sel_969016 = array_index_968791 == array_index_948823 ? add_969015 : sel_969012;
  assign add_969019 = sel_969016 + 8'h01;
  assign sel_969020 = array_index_968791 == array_index_948829 ? add_969019 : sel_969016;
  assign add_969023 = sel_969020 + 8'h01;
  assign sel_969024 = array_index_968791 == array_index_948835 ? add_969023 : sel_969020;
  assign add_969027 = sel_969024 + 8'h01;
  assign sel_969028 = array_index_968791 == array_index_948841 ? add_969027 : sel_969024;
  assign add_969031 = sel_969028 + 8'h01;
  assign sel_969032 = array_index_968791 == array_index_948847 ? add_969031 : sel_969028;
  assign add_969035 = sel_969032 + 8'h01;
  assign sel_969036 = array_index_968791 == array_index_948853 ? add_969035 : sel_969032;
  assign add_969039 = sel_969036 + 8'h01;
  assign sel_969040 = array_index_968791 == array_index_948859 ? add_969039 : sel_969036;
  assign add_969043 = sel_969040 + 8'h01;
  assign sel_969044 = array_index_968791 == array_index_948865 ? add_969043 : sel_969040;
  assign add_969047 = sel_969044 + 8'h01;
  assign sel_969048 = array_index_968791 == array_index_948871 ? add_969047 : sel_969044;
  assign add_969051 = sel_969048 + 8'h01;
  assign sel_969052 = array_index_968791 == array_index_948877 ? add_969051 : sel_969048;
  assign add_969055 = sel_969052 + 8'h01;
  assign sel_969056 = array_index_968791 == array_index_948883 ? add_969055 : sel_969052;
  assign add_969059 = sel_969056 + 8'h01;
  assign sel_969060 = array_index_968791 == array_index_948889 ? add_969059 : sel_969056;
  assign add_969063 = sel_969060 + 8'h01;
  assign sel_969064 = array_index_968791 == array_index_948895 ? add_969063 : sel_969060;
  assign add_969067 = sel_969064 + 8'h01;
  assign sel_969068 = array_index_968791 == array_index_948901 ? add_969067 : sel_969064;
  assign add_969071 = sel_969068 + 8'h01;
  assign sel_969072 = array_index_968791 == array_index_948907 ? add_969071 : sel_969068;
  assign add_969075 = sel_969072 + 8'h01;
  assign sel_969076 = array_index_968791 == array_index_948913 ? add_969075 : sel_969072;
  assign add_969079 = sel_969076 + 8'h01;
  assign sel_969080 = array_index_968791 == array_index_948919 ? add_969079 : sel_969076;
  assign add_969083 = sel_969080 + 8'h01;
  assign sel_969084 = array_index_968791 == array_index_948925 ? add_969083 : sel_969080;
  assign add_969087 = sel_969084 + 8'h01;
  assign sel_969088 = array_index_968791 == array_index_948931 ? add_969087 : sel_969084;
  assign add_969091 = sel_969088 + 8'h01;
  assign sel_969092 = array_index_968791 == array_index_948937 ? add_969091 : sel_969088;
  assign add_969095 = sel_969092 + 8'h01;
  assign sel_969096 = array_index_968791 == array_index_948943 ? add_969095 : sel_969092;
  assign add_969099 = sel_969096 + 8'h01;
  assign sel_969100 = array_index_968791 == array_index_948949 ? add_969099 : sel_969096;
  assign add_969103 = sel_969100 + 8'h01;
  assign sel_969104 = array_index_968791 == array_index_948955 ? add_969103 : sel_969100;
  assign add_969107 = sel_969104 + 8'h01;
  assign sel_969108 = array_index_968791 == array_index_948961 ? add_969107 : sel_969104;
  assign add_969111 = sel_969108 + 8'h01;
  assign sel_969112 = array_index_968791 == array_index_948967 ? add_969111 : sel_969108;
  assign add_969115 = sel_969112 + 8'h01;
  assign sel_969116 = array_index_968791 == array_index_948973 ? add_969115 : sel_969112;
  assign add_969119 = sel_969116 + 8'h01;
  assign sel_969120 = array_index_968791 == array_index_948979 ? add_969119 : sel_969116;
  assign add_969123 = sel_969120 + 8'h01;
  assign sel_969124 = array_index_968791 == array_index_948985 ? add_969123 : sel_969120;
  assign add_969127 = sel_969124 + 8'h01;
  assign sel_969128 = array_index_968791 == array_index_948991 ? add_969127 : sel_969124;
  assign add_969131 = sel_969128 + 8'h01;
  assign sel_969132 = array_index_968791 == array_index_948997 ? add_969131 : sel_969128;
  assign add_969135 = sel_969132 + 8'h01;
  assign sel_969136 = array_index_968791 == array_index_949003 ? add_969135 : sel_969132;
  assign add_969139 = sel_969136 + 8'h01;
  assign sel_969140 = array_index_968791 == array_index_949009 ? add_969139 : sel_969136;
  assign add_969143 = sel_969140 + 8'h01;
  assign sel_969144 = array_index_968791 == array_index_949015 ? add_969143 : sel_969140;
  assign add_969147 = sel_969144 + 8'h01;
  assign sel_969148 = array_index_968791 == array_index_949021 ? add_969147 : sel_969144;
  assign add_969151 = sel_969148 + 8'h01;
  assign sel_969152 = array_index_968791 == array_index_949027 ? add_969151 : sel_969148;
  assign add_969155 = sel_969152 + 8'h01;
  assign sel_969156 = array_index_968791 == array_index_949033 ? add_969155 : sel_969152;
  assign add_969159 = sel_969156 + 8'h01;
  assign sel_969160 = array_index_968791 == array_index_949039 ? add_969159 : sel_969156;
  assign add_969163 = sel_969160 + 8'h01;
  assign sel_969164 = array_index_968791 == array_index_949045 ? add_969163 : sel_969160;
  assign add_969167 = sel_969164 + 8'h01;
  assign sel_969168 = array_index_968791 == array_index_949051 ? add_969167 : sel_969164;
  assign add_969171 = sel_969168 + 8'h01;
  assign sel_969172 = array_index_968791 == array_index_949057 ? add_969171 : sel_969168;
  assign add_969175 = sel_969172 + 8'h01;
  assign sel_969176 = array_index_968791 == array_index_949063 ? add_969175 : sel_969172;
  assign add_969179 = sel_969176 + 8'h01;
  assign sel_969180 = array_index_968791 == array_index_949069 ? add_969179 : sel_969176;
  assign add_969183 = sel_969180 + 8'h01;
  assign sel_969184 = array_index_968791 == array_index_949075 ? add_969183 : sel_969180;
  assign add_969187 = sel_969184 + 8'h01;
  assign sel_969188 = array_index_968791 == array_index_949081 ? add_969187 : sel_969184;
  assign add_969192 = sel_969188 + 8'h01;
  assign array_index_969193 = set1_unflattened[7'h33];
  assign sel_969194 = array_index_968791 == array_index_949087 ? add_969192 : sel_969188;
  assign add_969197 = sel_969194 + 8'h01;
  assign sel_969198 = array_index_969193 == array_index_948483 ? add_969197 : sel_969194;
  assign add_969201 = sel_969198 + 8'h01;
  assign sel_969202 = array_index_969193 == array_index_948487 ? add_969201 : sel_969198;
  assign add_969205 = sel_969202 + 8'h01;
  assign sel_969206 = array_index_969193 == array_index_948495 ? add_969205 : sel_969202;
  assign add_969209 = sel_969206 + 8'h01;
  assign sel_969210 = array_index_969193 == array_index_948503 ? add_969209 : sel_969206;
  assign add_969213 = sel_969210 + 8'h01;
  assign sel_969214 = array_index_969193 == array_index_948511 ? add_969213 : sel_969210;
  assign add_969217 = sel_969214 + 8'h01;
  assign sel_969218 = array_index_969193 == array_index_948519 ? add_969217 : sel_969214;
  assign add_969221 = sel_969218 + 8'h01;
  assign sel_969222 = array_index_969193 == array_index_948527 ? add_969221 : sel_969218;
  assign add_969225 = sel_969222 + 8'h01;
  assign sel_969226 = array_index_969193 == array_index_948535 ? add_969225 : sel_969222;
  assign add_969229 = sel_969226 + 8'h01;
  assign sel_969230 = array_index_969193 == array_index_948541 ? add_969229 : sel_969226;
  assign add_969233 = sel_969230 + 8'h01;
  assign sel_969234 = array_index_969193 == array_index_948547 ? add_969233 : sel_969230;
  assign add_969237 = sel_969234 + 8'h01;
  assign sel_969238 = array_index_969193 == array_index_948553 ? add_969237 : sel_969234;
  assign add_969241 = sel_969238 + 8'h01;
  assign sel_969242 = array_index_969193 == array_index_948559 ? add_969241 : sel_969238;
  assign add_969245 = sel_969242 + 8'h01;
  assign sel_969246 = array_index_969193 == array_index_948565 ? add_969245 : sel_969242;
  assign add_969249 = sel_969246 + 8'h01;
  assign sel_969250 = array_index_969193 == array_index_948571 ? add_969249 : sel_969246;
  assign add_969253 = sel_969250 + 8'h01;
  assign sel_969254 = array_index_969193 == array_index_948577 ? add_969253 : sel_969250;
  assign add_969257 = sel_969254 + 8'h01;
  assign sel_969258 = array_index_969193 == array_index_948583 ? add_969257 : sel_969254;
  assign add_969261 = sel_969258 + 8'h01;
  assign sel_969262 = array_index_969193 == array_index_948589 ? add_969261 : sel_969258;
  assign add_969265 = sel_969262 + 8'h01;
  assign sel_969266 = array_index_969193 == array_index_948595 ? add_969265 : sel_969262;
  assign add_969269 = sel_969266 + 8'h01;
  assign sel_969270 = array_index_969193 == array_index_948601 ? add_969269 : sel_969266;
  assign add_969273 = sel_969270 + 8'h01;
  assign sel_969274 = array_index_969193 == array_index_948607 ? add_969273 : sel_969270;
  assign add_969277 = sel_969274 + 8'h01;
  assign sel_969278 = array_index_969193 == array_index_948613 ? add_969277 : sel_969274;
  assign add_969281 = sel_969278 + 8'h01;
  assign sel_969282 = array_index_969193 == array_index_948619 ? add_969281 : sel_969278;
  assign add_969285 = sel_969282 + 8'h01;
  assign sel_969286 = array_index_969193 == array_index_948625 ? add_969285 : sel_969282;
  assign add_969289 = sel_969286 + 8'h01;
  assign sel_969290 = array_index_969193 == array_index_948631 ? add_969289 : sel_969286;
  assign add_969293 = sel_969290 + 8'h01;
  assign sel_969294 = array_index_969193 == array_index_948637 ? add_969293 : sel_969290;
  assign add_969297 = sel_969294 + 8'h01;
  assign sel_969298 = array_index_969193 == array_index_948643 ? add_969297 : sel_969294;
  assign add_969301 = sel_969298 + 8'h01;
  assign sel_969302 = array_index_969193 == array_index_948649 ? add_969301 : sel_969298;
  assign add_969305 = sel_969302 + 8'h01;
  assign sel_969306 = array_index_969193 == array_index_948655 ? add_969305 : sel_969302;
  assign add_969309 = sel_969306 + 8'h01;
  assign sel_969310 = array_index_969193 == array_index_948661 ? add_969309 : sel_969306;
  assign add_969313 = sel_969310 + 8'h01;
  assign sel_969314 = array_index_969193 == array_index_948667 ? add_969313 : sel_969310;
  assign add_969317 = sel_969314 + 8'h01;
  assign sel_969318 = array_index_969193 == array_index_948673 ? add_969317 : sel_969314;
  assign add_969321 = sel_969318 + 8'h01;
  assign sel_969322 = array_index_969193 == array_index_948679 ? add_969321 : sel_969318;
  assign add_969325 = sel_969322 + 8'h01;
  assign sel_969326 = array_index_969193 == array_index_948685 ? add_969325 : sel_969322;
  assign add_969329 = sel_969326 + 8'h01;
  assign sel_969330 = array_index_969193 == array_index_948691 ? add_969329 : sel_969326;
  assign add_969333 = sel_969330 + 8'h01;
  assign sel_969334 = array_index_969193 == array_index_948697 ? add_969333 : sel_969330;
  assign add_969337 = sel_969334 + 8'h01;
  assign sel_969338 = array_index_969193 == array_index_948703 ? add_969337 : sel_969334;
  assign add_969341 = sel_969338 + 8'h01;
  assign sel_969342 = array_index_969193 == array_index_948709 ? add_969341 : sel_969338;
  assign add_969345 = sel_969342 + 8'h01;
  assign sel_969346 = array_index_969193 == array_index_948715 ? add_969345 : sel_969342;
  assign add_969349 = sel_969346 + 8'h01;
  assign sel_969350 = array_index_969193 == array_index_948721 ? add_969349 : sel_969346;
  assign add_969353 = sel_969350 + 8'h01;
  assign sel_969354 = array_index_969193 == array_index_948727 ? add_969353 : sel_969350;
  assign add_969357 = sel_969354 + 8'h01;
  assign sel_969358 = array_index_969193 == array_index_948733 ? add_969357 : sel_969354;
  assign add_969361 = sel_969358 + 8'h01;
  assign sel_969362 = array_index_969193 == array_index_948739 ? add_969361 : sel_969358;
  assign add_969365 = sel_969362 + 8'h01;
  assign sel_969366 = array_index_969193 == array_index_948745 ? add_969365 : sel_969362;
  assign add_969369 = sel_969366 + 8'h01;
  assign sel_969370 = array_index_969193 == array_index_948751 ? add_969369 : sel_969366;
  assign add_969373 = sel_969370 + 8'h01;
  assign sel_969374 = array_index_969193 == array_index_948757 ? add_969373 : sel_969370;
  assign add_969377 = sel_969374 + 8'h01;
  assign sel_969378 = array_index_969193 == array_index_948763 ? add_969377 : sel_969374;
  assign add_969381 = sel_969378 + 8'h01;
  assign sel_969382 = array_index_969193 == array_index_948769 ? add_969381 : sel_969378;
  assign add_969385 = sel_969382 + 8'h01;
  assign sel_969386 = array_index_969193 == array_index_948775 ? add_969385 : sel_969382;
  assign add_969389 = sel_969386 + 8'h01;
  assign sel_969390 = array_index_969193 == array_index_948781 ? add_969389 : sel_969386;
  assign add_969393 = sel_969390 + 8'h01;
  assign sel_969394 = array_index_969193 == array_index_948787 ? add_969393 : sel_969390;
  assign add_969397 = sel_969394 + 8'h01;
  assign sel_969398 = array_index_969193 == array_index_948793 ? add_969397 : sel_969394;
  assign add_969401 = sel_969398 + 8'h01;
  assign sel_969402 = array_index_969193 == array_index_948799 ? add_969401 : sel_969398;
  assign add_969405 = sel_969402 + 8'h01;
  assign sel_969406 = array_index_969193 == array_index_948805 ? add_969405 : sel_969402;
  assign add_969409 = sel_969406 + 8'h01;
  assign sel_969410 = array_index_969193 == array_index_948811 ? add_969409 : sel_969406;
  assign add_969413 = sel_969410 + 8'h01;
  assign sel_969414 = array_index_969193 == array_index_948817 ? add_969413 : sel_969410;
  assign add_969417 = sel_969414 + 8'h01;
  assign sel_969418 = array_index_969193 == array_index_948823 ? add_969417 : sel_969414;
  assign add_969421 = sel_969418 + 8'h01;
  assign sel_969422 = array_index_969193 == array_index_948829 ? add_969421 : sel_969418;
  assign add_969425 = sel_969422 + 8'h01;
  assign sel_969426 = array_index_969193 == array_index_948835 ? add_969425 : sel_969422;
  assign add_969429 = sel_969426 + 8'h01;
  assign sel_969430 = array_index_969193 == array_index_948841 ? add_969429 : sel_969426;
  assign add_969433 = sel_969430 + 8'h01;
  assign sel_969434 = array_index_969193 == array_index_948847 ? add_969433 : sel_969430;
  assign add_969437 = sel_969434 + 8'h01;
  assign sel_969438 = array_index_969193 == array_index_948853 ? add_969437 : sel_969434;
  assign add_969441 = sel_969438 + 8'h01;
  assign sel_969442 = array_index_969193 == array_index_948859 ? add_969441 : sel_969438;
  assign add_969445 = sel_969442 + 8'h01;
  assign sel_969446 = array_index_969193 == array_index_948865 ? add_969445 : sel_969442;
  assign add_969449 = sel_969446 + 8'h01;
  assign sel_969450 = array_index_969193 == array_index_948871 ? add_969449 : sel_969446;
  assign add_969453 = sel_969450 + 8'h01;
  assign sel_969454 = array_index_969193 == array_index_948877 ? add_969453 : sel_969450;
  assign add_969457 = sel_969454 + 8'h01;
  assign sel_969458 = array_index_969193 == array_index_948883 ? add_969457 : sel_969454;
  assign add_969461 = sel_969458 + 8'h01;
  assign sel_969462 = array_index_969193 == array_index_948889 ? add_969461 : sel_969458;
  assign add_969465 = sel_969462 + 8'h01;
  assign sel_969466 = array_index_969193 == array_index_948895 ? add_969465 : sel_969462;
  assign add_969469 = sel_969466 + 8'h01;
  assign sel_969470 = array_index_969193 == array_index_948901 ? add_969469 : sel_969466;
  assign add_969473 = sel_969470 + 8'h01;
  assign sel_969474 = array_index_969193 == array_index_948907 ? add_969473 : sel_969470;
  assign add_969477 = sel_969474 + 8'h01;
  assign sel_969478 = array_index_969193 == array_index_948913 ? add_969477 : sel_969474;
  assign add_969481 = sel_969478 + 8'h01;
  assign sel_969482 = array_index_969193 == array_index_948919 ? add_969481 : sel_969478;
  assign add_969485 = sel_969482 + 8'h01;
  assign sel_969486 = array_index_969193 == array_index_948925 ? add_969485 : sel_969482;
  assign add_969489 = sel_969486 + 8'h01;
  assign sel_969490 = array_index_969193 == array_index_948931 ? add_969489 : sel_969486;
  assign add_969493 = sel_969490 + 8'h01;
  assign sel_969494 = array_index_969193 == array_index_948937 ? add_969493 : sel_969490;
  assign add_969497 = sel_969494 + 8'h01;
  assign sel_969498 = array_index_969193 == array_index_948943 ? add_969497 : sel_969494;
  assign add_969501 = sel_969498 + 8'h01;
  assign sel_969502 = array_index_969193 == array_index_948949 ? add_969501 : sel_969498;
  assign add_969505 = sel_969502 + 8'h01;
  assign sel_969506 = array_index_969193 == array_index_948955 ? add_969505 : sel_969502;
  assign add_969509 = sel_969506 + 8'h01;
  assign sel_969510 = array_index_969193 == array_index_948961 ? add_969509 : sel_969506;
  assign add_969513 = sel_969510 + 8'h01;
  assign sel_969514 = array_index_969193 == array_index_948967 ? add_969513 : sel_969510;
  assign add_969517 = sel_969514 + 8'h01;
  assign sel_969518 = array_index_969193 == array_index_948973 ? add_969517 : sel_969514;
  assign add_969521 = sel_969518 + 8'h01;
  assign sel_969522 = array_index_969193 == array_index_948979 ? add_969521 : sel_969518;
  assign add_969525 = sel_969522 + 8'h01;
  assign sel_969526 = array_index_969193 == array_index_948985 ? add_969525 : sel_969522;
  assign add_969529 = sel_969526 + 8'h01;
  assign sel_969530 = array_index_969193 == array_index_948991 ? add_969529 : sel_969526;
  assign add_969533 = sel_969530 + 8'h01;
  assign sel_969534 = array_index_969193 == array_index_948997 ? add_969533 : sel_969530;
  assign add_969537 = sel_969534 + 8'h01;
  assign sel_969538 = array_index_969193 == array_index_949003 ? add_969537 : sel_969534;
  assign add_969541 = sel_969538 + 8'h01;
  assign sel_969542 = array_index_969193 == array_index_949009 ? add_969541 : sel_969538;
  assign add_969545 = sel_969542 + 8'h01;
  assign sel_969546 = array_index_969193 == array_index_949015 ? add_969545 : sel_969542;
  assign add_969549 = sel_969546 + 8'h01;
  assign sel_969550 = array_index_969193 == array_index_949021 ? add_969549 : sel_969546;
  assign add_969553 = sel_969550 + 8'h01;
  assign sel_969554 = array_index_969193 == array_index_949027 ? add_969553 : sel_969550;
  assign add_969557 = sel_969554 + 8'h01;
  assign sel_969558 = array_index_969193 == array_index_949033 ? add_969557 : sel_969554;
  assign add_969561 = sel_969558 + 8'h01;
  assign sel_969562 = array_index_969193 == array_index_949039 ? add_969561 : sel_969558;
  assign add_969565 = sel_969562 + 8'h01;
  assign sel_969566 = array_index_969193 == array_index_949045 ? add_969565 : sel_969562;
  assign add_969569 = sel_969566 + 8'h01;
  assign sel_969570 = array_index_969193 == array_index_949051 ? add_969569 : sel_969566;
  assign add_969573 = sel_969570 + 8'h01;
  assign sel_969574 = array_index_969193 == array_index_949057 ? add_969573 : sel_969570;
  assign add_969577 = sel_969574 + 8'h01;
  assign sel_969578 = array_index_969193 == array_index_949063 ? add_969577 : sel_969574;
  assign add_969581 = sel_969578 + 8'h01;
  assign sel_969582 = array_index_969193 == array_index_949069 ? add_969581 : sel_969578;
  assign add_969585 = sel_969582 + 8'h01;
  assign sel_969586 = array_index_969193 == array_index_949075 ? add_969585 : sel_969582;
  assign add_969589 = sel_969586 + 8'h01;
  assign sel_969590 = array_index_969193 == array_index_949081 ? add_969589 : sel_969586;
  assign add_969594 = sel_969590 + 8'h01;
  assign array_index_969595 = set1_unflattened[7'h34];
  assign sel_969596 = array_index_969193 == array_index_949087 ? add_969594 : sel_969590;
  assign add_969599 = sel_969596 + 8'h01;
  assign sel_969600 = array_index_969595 == array_index_948483 ? add_969599 : sel_969596;
  assign add_969603 = sel_969600 + 8'h01;
  assign sel_969604 = array_index_969595 == array_index_948487 ? add_969603 : sel_969600;
  assign add_969607 = sel_969604 + 8'h01;
  assign sel_969608 = array_index_969595 == array_index_948495 ? add_969607 : sel_969604;
  assign add_969611 = sel_969608 + 8'h01;
  assign sel_969612 = array_index_969595 == array_index_948503 ? add_969611 : sel_969608;
  assign add_969615 = sel_969612 + 8'h01;
  assign sel_969616 = array_index_969595 == array_index_948511 ? add_969615 : sel_969612;
  assign add_969619 = sel_969616 + 8'h01;
  assign sel_969620 = array_index_969595 == array_index_948519 ? add_969619 : sel_969616;
  assign add_969623 = sel_969620 + 8'h01;
  assign sel_969624 = array_index_969595 == array_index_948527 ? add_969623 : sel_969620;
  assign add_969627 = sel_969624 + 8'h01;
  assign sel_969628 = array_index_969595 == array_index_948535 ? add_969627 : sel_969624;
  assign add_969631 = sel_969628 + 8'h01;
  assign sel_969632 = array_index_969595 == array_index_948541 ? add_969631 : sel_969628;
  assign add_969635 = sel_969632 + 8'h01;
  assign sel_969636 = array_index_969595 == array_index_948547 ? add_969635 : sel_969632;
  assign add_969639 = sel_969636 + 8'h01;
  assign sel_969640 = array_index_969595 == array_index_948553 ? add_969639 : sel_969636;
  assign add_969643 = sel_969640 + 8'h01;
  assign sel_969644 = array_index_969595 == array_index_948559 ? add_969643 : sel_969640;
  assign add_969647 = sel_969644 + 8'h01;
  assign sel_969648 = array_index_969595 == array_index_948565 ? add_969647 : sel_969644;
  assign add_969651 = sel_969648 + 8'h01;
  assign sel_969652 = array_index_969595 == array_index_948571 ? add_969651 : sel_969648;
  assign add_969655 = sel_969652 + 8'h01;
  assign sel_969656 = array_index_969595 == array_index_948577 ? add_969655 : sel_969652;
  assign add_969659 = sel_969656 + 8'h01;
  assign sel_969660 = array_index_969595 == array_index_948583 ? add_969659 : sel_969656;
  assign add_969663 = sel_969660 + 8'h01;
  assign sel_969664 = array_index_969595 == array_index_948589 ? add_969663 : sel_969660;
  assign add_969667 = sel_969664 + 8'h01;
  assign sel_969668 = array_index_969595 == array_index_948595 ? add_969667 : sel_969664;
  assign add_969671 = sel_969668 + 8'h01;
  assign sel_969672 = array_index_969595 == array_index_948601 ? add_969671 : sel_969668;
  assign add_969675 = sel_969672 + 8'h01;
  assign sel_969676 = array_index_969595 == array_index_948607 ? add_969675 : sel_969672;
  assign add_969679 = sel_969676 + 8'h01;
  assign sel_969680 = array_index_969595 == array_index_948613 ? add_969679 : sel_969676;
  assign add_969683 = sel_969680 + 8'h01;
  assign sel_969684 = array_index_969595 == array_index_948619 ? add_969683 : sel_969680;
  assign add_969687 = sel_969684 + 8'h01;
  assign sel_969688 = array_index_969595 == array_index_948625 ? add_969687 : sel_969684;
  assign add_969691 = sel_969688 + 8'h01;
  assign sel_969692 = array_index_969595 == array_index_948631 ? add_969691 : sel_969688;
  assign add_969695 = sel_969692 + 8'h01;
  assign sel_969696 = array_index_969595 == array_index_948637 ? add_969695 : sel_969692;
  assign add_969699 = sel_969696 + 8'h01;
  assign sel_969700 = array_index_969595 == array_index_948643 ? add_969699 : sel_969696;
  assign add_969703 = sel_969700 + 8'h01;
  assign sel_969704 = array_index_969595 == array_index_948649 ? add_969703 : sel_969700;
  assign add_969707 = sel_969704 + 8'h01;
  assign sel_969708 = array_index_969595 == array_index_948655 ? add_969707 : sel_969704;
  assign add_969711 = sel_969708 + 8'h01;
  assign sel_969712 = array_index_969595 == array_index_948661 ? add_969711 : sel_969708;
  assign add_969715 = sel_969712 + 8'h01;
  assign sel_969716 = array_index_969595 == array_index_948667 ? add_969715 : sel_969712;
  assign add_969719 = sel_969716 + 8'h01;
  assign sel_969720 = array_index_969595 == array_index_948673 ? add_969719 : sel_969716;
  assign add_969723 = sel_969720 + 8'h01;
  assign sel_969724 = array_index_969595 == array_index_948679 ? add_969723 : sel_969720;
  assign add_969727 = sel_969724 + 8'h01;
  assign sel_969728 = array_index_969595 == array_index_948685 ? add_969727 : sel_969724;
  assign add_969731 = sel_969728 + 8'h01;
  assign sel_969732 = array_index_969595 == array_index_948691 ? add_969731 : sel_969728;
  assign add_969735 = sel_969732 + 8'h01;
  assign sel_969736 = array_index_969595 == array_index_948697 ? add_969735 : sel_969732;
  assign add_969739 = sel_969736 + 8'h01;
  assign sel_969740 = array_index_969595 == array_index_948703 ? add_969739 : sel_969736;
  assign add_969743 = sel_969740 + 8'h01;
  assign sel_969744 = array_index_969595 == array_index_948709 ? add_969743 : sel_969740;
  assign add_969747 = sel_969744 + 8'h01;
  assign sel_969748 = array_index_969595 == array_index_948715 ? add_969747 : sel_969744;
  assign add_969751 = sel_969748 + 8'h01;
  assign sel_969752 = array_index_969595 == array_index_948721 ? add_969751 : sel_969748;
  assign add_969755 = sel_969752 + 8'h01;
  assign sel_969756 = array_index_969595 == array_index_948727 ? add_969755 : sel_969752;
  assign add_969759 = sel_969756 + 8'h01;
  assign sel_969760 = array_index_969595 == array_index_948733 ? add_969759 : sel_969756;
  assign add_969763 = sel_969760 + 8'h01;
  assign sel_969764 = array_index_969595 == array_index_948739 ? add_969763 : sel_969760;
  assign add_969767 = sel_969764 + 8'h01;
  assign sel_969768 = array_index_969595 == array_index_948745 ? add_969767 : sel_969764;
  assign add_969771 = sel_969768 + 8'h01;
  assign sel_969772 = array_index_969595 == array_index_948751 ? add_969771 : sel_969768;
  assign add_969775 = sel_969772 + 8'h01;
  assign sel_969776 = array_index_969595 == array_index_948757 ? add_969775 : sel_969772;
  assign add_969779 = sel_969776 + 8'h01;
  assign sel_969780 = array_index_969595 == array_index_948763 ? add_969779 : sel_969776;
  assign add_969783 = sel_969780 + 8'h01;
  assign sel_969784 = array_index_969595 == array_index_948769 ? add_969783 : sel_969780;
  assign add_969787 = sel_969784 + 8'h01;
  assign sel_969788 = array_index_969595 == array_index_948775 ? add_969787 : sel_969784;
  assign add_969791 = sel_969788 + 8'h01;
  assign sel_969792 = array_index_969595 == array_index_948781 ? add_969791 : sel_969788;
  assign add_969795 = sel_969792 + 8'h01;
  assign sel_969796 = array_index_969595 == array_index_948787 ? add_969795 : sel_969792;
  assign add_969799 = sel_969796 + 8'h01;
  assign sel_969800 = array_index_969595 == array_index_948793 ? add_969799 : sel_969796;
  assign add_969803 = sel_969800 + 8'h01;
  assign sel_969804 = array_index_969595 == array_index_948799 ? add_969803 : sel_969800;
  assign add_969807 = sel_969804 + 8'h01;
  assign sel_969808 = array_index_969595 == array_index_948805 ? add_969807 : sel_969804;
  assign add_969811 = sel_969808 + 8'h01;
  assign sel_969812 = array_index_969595 == array_index_948811 ? add_969811 : sel_969808;
  assign add_969815 = sel_969812 + 8'h01;
  assign sel_969816 = array_index_969595 == array_index_948817 ? add_969815 : sel_969812;
  assign add_969819 = sel_969816 + 8'h01;
  assign sel_969820 = array_index_969595 == array_index_948823 ? add_969819 : sel_969816;
  assign add_969823 = sel_969820 + 8'h01;
  assign sel_969824 = array_index_969595 == array_index_948829 ? add_969823 : sel_969820;
  assign add_969827 = sel_969824 + 8'h01;
  assign sel_969828 = array_index_969595 == array_index_948835 ? add_969827 : sel_969824;
  assign add_969831 = sel_969828 + 8'h01;
  assign sel_969832 = array_index_969595 == array_index_948841 ? add_969831 : sel_969828;
  assign add_969835 = sel_969832 + 8'h01;
  assign sel_969836 = array_index_969595 == array_index_948847 ? add_969835 : sel_969832;
  assign add_969839 = sel_969836 + 8'h01;
  assign sel_969840 = array_index_969595 == array_index_948853 ? add_969839 : sel_969836;
  assign add_969843 = sel_969840 + 8'h01;
  assign sel_969844 = array_index_969595 == array_index_948859 ? add_969843 : sel_969840;
  assign add_969847 = sel_969844 + 8'h01;
  assign sel_969848 = array_index_969595 == array_index_948865 ? add_969847 : sel_969844;
  assign add_969851 = sel_969848 + 8'h01;
  assign sel_969852 = array_index_969595 == array_index_948871 ? add_969851 : sel_969848;
  assign add_969855 = sel_969852 + 8'h01;
  assign sel_969856 = array_index_969595 == array_index_948877 ? add_969855 : sel_969852;
  assign add_969859 = sel_969856 + 8'h01;
  assign sel_969860 = array_index_969595 == array_index_948883 ? add_969859 : sel_969856;
  assign add_969863 = sel_969860 + 8'h01;
  assign sel_969864 = array_index_969595 == array_index_948889 ? add_969863 : sel_969860;
  assign add_969867 = sel_969864 + 8'h01;
  assign sel_969868 = array_index_969595 == array_index_948895 ? add_969867 : sel_969864;
  assign add_969871 = sel_969868 + 8'h01;
  assign sel_969872 = array_index_969595 == array_index_948901 ? add_969871 : sel_969868;
  assign add_969875 = sel_969872 + 8'h01;
  assign sel_969876 = array_index_969595 == array_index_948907 ? add_969875 : sel_969872;
  assign add_969879 = sel_969876 + 8'h01;
  assign sel_969880 = array_index_969595 == array_index_948913 ? add_969879 : sel_969876;
  assign add_969883 = sel_969880 + 8'h01;
  assign sel_969884 = array_index_969595 == array_index_948919 ? add_969883 : sel_969880;
  assign add_969887 = sel_969884 + 8'h01;
  assign sel_969888 = array_index_969595 == array_index_948925 ? add_969887 : sel_969884;
  assign add_969891 = sel_969888 + 8'h01;
  assign sel_969892 = array_index_969595 == array_index_948931 ? add_969891 : sel_969888;
  assign add_969895 = sel_969892 + 8'h01;
  assign sel_969896 = array_index_969595 == array_index_948937 ? add_969895 : sel_969892;
  assign add_969899 = sel_969896 + 8'h01;
  assign sel_969900 = array_index_969595 == array_index_948943 ? add_969899 : sel_969896;
  assign add_969903 = sel_969900 + 8'h01;
  assign sel_969904 = array_index_969595 == array_index_948949 ? add_969903 : sel_969900;
  assign add_969907 = sel_969904 + 8'h01;
  assign sel_969908 = array_index_969595 == array_index_948955 ? add_969907 : sel_969904;
  assign add_969911 = sel_969908 + 8'h01;
  assign sel_969912 = array_index_969595 == array_index_948961 ? add_969911 : sel_969908;
  assign add_969915 = sel_969912 + 8'h01;
  assign sel_969916 = array_index_969595 == array_index_948967 ? add_969915 : sel_969912;
  assign add_969919 = sel_969916 + 8'h01;
  assign sel_969920 = array_index_969595 == array_index_948973 ? add_969919 : sel_969916;
  assign add_969923 = sel_969920 + 8'h01;
  assign sel_969924 = array_index_969595 == array_index_948979 ? add_969923 : sel_969920;
  assign add_969927 = sel_969924 + 8'h01;
  assign sel_969928 = array_index_969595 == array_index_948985 ? add_969927 : sel_969924;
  assign add_969931 = sel_969928 + 8'h01;
  assign sel_969932 = array_index_969595 == array_index_948991 ? add_969931 : sel_969928;
  assign add_969935 = sel_969932 + 8'h01;
  assign sel_969936 = array_index_969595 == array_index_948997 ? add_969935 : sel_969932;
  assign add_969939 = sel_969936 + 8'h01;
  assign sel_969940 = array_index_969595 == array_index_949003 ? add_969939 : sel_969936;
  assign add_969943 = sel_969940 + 8'h01;
  assign sel_969944 = array_index_969595 == array_index_949009 ? add_969943 : sel_969940;
  assign add_969947 = sel_969944 + 8'h01;
  assign sel_969948 = array_index_969595 == array_index_949015 ? add_969947 : sel_969944;
  assign add_969951 = sel_969948 + 8'h01;
  assign sel_969952 = array_index_969595 == array_index_949021 ? add_969951 : sel_969948;
  assign add_969955 = sel_969952 + 8'h01;
  assign sel_969956 = array_index_969595 == array_index_949027 ? add_969955 : sel_969952;
  assign add_969959 = sel_969956 + 8'h01;
  assign sel_969960 = array_index_969595 == array_index_949033 ? add_969959 : sel_969956;
  assign add_969963 = sel_969960 + 8'h01;
  assign sel_969964 = array_index_969595 == array_index_949039 ? add_969963 : sel_969960;
  assign add_969967 = sel_969964 + 8'h01;
  assign sel_969968 = array_index_969595 == array_index_949045 ? add_969967 : sel_969964;
  assign add_969971 = sel_969968 + 8'h01;
  assign sel_969972 = array_index_969595 == array_index_949051 ? add_969971 : sel_969968;
  assign add_969975 = sel_969972 + 8'h01;
  assign sel_969976 = array_index_969595 == array_index_949057 ? add_969975 : sel_969972;
  assign add_969979 = sel_969976 + 8'h01;
  assign sel_969980 = array_index_969595 == array_index_949063 ? add_969979 : sel_969976;
  assign add_969983 = sel_969980 + 8'h01;
  assign sel_969984 = array_index_969595 == array_index_949069 ? add_969983 : sel_969980;
  assign add_969987 = sel_969984 + 8'h01;
  assign sel_969988 = array_index_969595 == array_index_949075 ? add_969987 : sel_969984;
  assign add_969991 = sel_969988 + 8'h01;
  assign sel_969992 = array_index_969595 == array_index_949081 ? add_969991 : sel_969988;
  assign add_969996 = sel_969992 + 8'h01;
  assign array_index_969997 = set1_unflattened[7'h35];
  assign sel_969998 = array_index_969595 == array_index_949087 ? add_969996 : sel_969992;
  assign add_970001 = sel_969998 + 8'h01;
  assign sel_970002 = array_index_969997 == array_index_948483 ? add_970001 : sel_969998;
  assign add_970005 = sel_970002 + 8'h01;
  assign sel_970006 = array_index_969997 == array_index_948487 ? add_970005 : sel_970002;
  assign add_970009 = sel_970006 + 8'h01;
  assign sel_970010 = array_index_969997 == array_index_948495 ? add_970009 : sel_970006;
  assign add_970013 = sel_970010 + 8'h01;
  assign sel_970014 = array_index_969997 == array_index_948503 ? add_970013 : sel_970010;
  assign add_970017 = sel_970014 + 8'h01;
  assign sel_970018 = array_index_969997 == array_index_948511 ? add_970017 : sel_970014;
  assign add_970021 = sel_970018 + 8'h01;
  assign sel_970022 = array_index_969997 == array_index_948519 ? add_970021 : sel_970018;
  assign add_970025 = sel_970022 + 8'h01;
  assign sel_970026 = array_index_969997 == array_index_948527 ? add_970025 : sel_970022;
  assign add_970029 = sel_970026 + 8'h01;
  assign sel_970030 = array_index_969997 == array_index_948535 ? add_970029 : sel_970026;
  assign add_970033 = sel_970030 + 8'h01;
  assign sel_970034 = array_index_969997 == array_index_948541 ? add_970033 : sel_970030;
  assign add_970037 = sel_970034 + 8'h01;
  assign sel_970038 = array_index_969997 == array_index_948547 ? add_970037 : sel_970034;
  assign add_970041 = sel_970038 + 8'h01;
  assign sel_970042 = array_index_969997 == array_index_948553 ? add_970041 : sel_970038;
  assign add_970045 = sel_970042 + 8'h01;
  assign sel_970046 = array_index_969997 == array_index_948559 ? add_970045 : sel_970042;
  assign add_970049 = sel_970046 + 8'h01;
  assign sel_970050 = array_index_969997 == array_index_948565 ? add_970049 : sel_970046;
  assign add_970053 = sel_970050 + 8'h01;
  assign sel_970054 = array_index_969997 == array_index_948571 ? add_970053 : sel_970050;
  assign add_970057 = sel_970054 + 8'h01;
  assign sel_970058 = array_index_969997 == array_index_948577 ? add_970057 : sel_970054;
  assign add_970061 = sel_970058 + 8'h01;
  assign sel_970062 = array_index_969997 == array_index_948583 ? add_970061 : sel_970058;
  assign add_970065 = sel_970062 + 8'h01;
  assign sel_970066 = array_index_969997 == array_index_948589 ? add_970065 : sel_970062;
  assign add_970069 = sel_970066 + 8'h01;
  assign sel_970070 = array_index_969997 == array_index_948595 ? add_970069 : sel_970066;
  assign add_970073 = sel_970070 + 8'h01;
  assign sel_970074 = array_index_969997 == array_index_948601 ? add_970073 : sel_970070;
  assign add_970077 = sel_970074 + 8'h01;
  assign sel_970078 = array_index_969997 == array_index_948607 ? add_970077 : sel_970074;
  assign add_970081 = sel_970078 + 8'h01;
  assign sel_970082 = array_index_969997 == array_index_948613 ? add_970081 : sel_970078;
  assign add_970085 = sel_970082 + 8'h01;
  assign sel_970086 = array_index_969997 == array_index_948619 ? add_970085 : sel_970082;
  assign add_970089 = sel_970086 + 8'h01;
  assign sel_970090 = array_index_969997 == array_index_948625 ? add_970089 : sel_970086;
  assign add_970093 = sel_970090 + 8'h01;
  assign sel_970094 = array_index_969997 == array_index_948631 ? add_970093 : sel_970090;
  assign add_970097 = sel_970094 + 8'h01;
  assign sel_970098 = array_index_969997 == array_index_948637 ? add_970097 : sel_970094;
  assign add_970101 = sel_970098 + 8'h01;
  assign sel_970102 = array_index_969997 == array_index_948643 ? add_970101 : sel_970098;
  assign add_970105 = sel_970102 + 8'h01;
  assign sel_970106 = array_index_969997 == array_index_948649 ? add_970105 : sel_970102;
  assign add_970109 = sel_970106 + 8'h01;
  assign sel_970110 = array_index_969997 == array_index_948655 ? add_970109 : sel_970106;
  assign add_970113 = sel_970110 + 8'h01;
  assign sel_970114 = array_index_969997 == array_index_948661 ? add_970113 : sel_970110;
  assign add_970117 = sel_970114 + 8'h01;
  assign sel_970118 = array_index_969997 == array_index_948667 ? add_970117 : sel_970114;
  assign add_970121 = sel_970118 + 8'h01;
  assign sel_970122 = array_index_969997 == array_index_948673 ? add_970121 : sel_970118;
  assign add_970125 = sel_970122 + 8'h01;
  assign sel_970126 = array_index_969997 == array_index_948679 ? add_970125 : sel_970122;
  assign add_970129 = sel_970126 + 8'h01;
  assign sel_970130 = array_index_969997 == array_index_948685 ? add_970129 : sel_970126;
  assign add_970133 = sel_970130 + 8'h01;
  assign sel_970134 = array_index_969997 == array_index_948691 ? add_970133 : sel_970130;
  assign add_970137 = sel_970134 + 8'h01;
  assign sel_970138 = array_index_969997 == array_index_948697 ? add_970137 : sel_970134;
  assign add_970141 = sel_970138 + 8'h01;
  assign sel_970142 = array_index_969997 == array_index_948703 ? add_970141 : sel_970138;
  assign add_970145 = sel_970142 + 8'h01;
  assign sel_970146 = array_index_969997 == array_index_948709 ? add_970145 : sel_970142;
  assign add_970149 = sel_970146 + 8'h01;
  assign sel_970150 = array_index_969997 == array_index_948715 ? add_970149 : sel_970146;
  assign add_970153 = sel_970150 + 8'h01;
  assign sel_970154 = array_index_969997 == array_index_948721 ? add_970153 : sel_970150;
  assign add_970157 = sel_970154 + 8'h01;
  assign sel_970158 = array_index_969997 == array_index_948727 ? add_970157 : sel_970154;
  assign add_970161 = sel_970158 + 8'h01;
  assign sel_970162 = array_index_969997 == array_index_948733 ? add_970161 : sel_970158;
  assign add_970165 = sel_970162 + 8'h01;
  assign sel_970166 = array_index_969997 == array_index_948739 ? add_970165 : sel_970162;
  assign add_970169 = sel_970166 + 8'h01;
  assign sel_970170 = array_index_969997 == array_index_948745 ? add_970169 : sel_970166;
  assign add_970173 = sel_970170 + 8'h01;
  assign sel_970174 = array_index_969997 == array_index_948751 ? add_970173 : sel_970170;
  assign add_970177 = sel_970174 + 8'h01;
  assign sel_970178 = array_index_969997 == array_index_948757 ? add_970177 : sel_970174;
  assign add_970181 = sel_970178 + 8'h01;
  assign sel_970182 = array_index_969997 == array_index_948763 ? add_970181 : sel_970178;
  assign add_970185 = sel_970182 + 8'h01;
  assign sel_970186 = array_index_969997 == array_index_948769 ? add_970185 : sel_970182;
  assign add_970189 = sel_970186 + 8'h01;
  assign sel_970190 = array_index_969997 == array_index_948775 ? add_970189 : sel_970186;
  assign add_970193 = sel_970190 + 8'h01;
  assign sel_970194 = array_index_969997 == array_index_948781 ? add_970193 : sel_970190;
  assign add_970197 = sel_970194 + 8'h01;
  assign sel_970198 = array_index_969997 == array_index_948787 ? add_970197 : sel_970194;
  assign add_970201 = sel_970198 + 8'h01;
  assign sel_970202 = array_index_969997 == array_index_948793 ? add_970201 : sel_970198;
  assign add_970205 = sel_970202 + 8'h01;
  assign sel_970206 = array_index_969997 == array_index_948799 ? add_970205 : sel_970202;
  assign add_970209 = sel_970206 + 8'h01;
  assign sel_970210 = array_index_969997 == array_index_948805 ? add_970209 : sel_970206;
  assign add_970213 = sel_970210 + 8'h01;
  assign sel_970214 = array_index_969997 == array_index_948811 ? add_970213 : sel_970210;
  assign add_970217 = sel_970214 + 8'h01;
  assign sel_970218 = array_index_969997 == array_index_948817 ? add_970217 : sel_970214;
  assign add_970221 = sel_970218 + 8'h01;
  assign sel_970222 = array_index_969997 == array_index_948823 ? add_970221 : sel_970218;
  assign add_970225 = sel_970222 + 8'h01;
  assign sel_970226 = array_index_969997 == array_index_948829 ? add_970225 : sel_970222;
  assign add_970229 = sel_970226 + 8'h01;
  assign sel_970230 = array_index_969997 == array_index_948835 ? add_970229 : sel_970226;
  assign add_970233 = sel_970230 + 8'h01;
  assign sel_970234 = array_index_969997 == array_index_948841 ? add_970233 : sel_970230;
  assign add_970237 = sel_970234 + 8'h01;
  assign sel_970238 = array_index_969997 == array_index_948847 ? add_970237 : sel_970234;
  assign add_970241 = sel_970238 + 8'h01;
  assign sel_970242 = array_index_969997 == array_index_948853 ? add_970241 : sel_970238;
  assign add_970245 = sel_970242 + 8'h01;
  assign sel_970246 = array_index_969997 == array_index_948859 ? add_970245 : sel_970242;
  assign add_970249 = sel_970246 + 8'h01;
  assign sel_970250 = array_index_969997 == array_index_948865 ? add_970249 : sel_970246;
  assign add_970253 = sel_970250 + 8'h01;
  assign sel_970254 = array_index_969997 == array_index_948871 ? add_970253 : sel_970250;
  assign add_970257 = sel_970254 + 8'h01;
  assign sel_970258 = array_index_969997 == array_index_948877 ? add_970257 : sel_970254;
  assign add_970261 = sel_970258 + 8'h01;
  assign sel_970262 = array_index_969997 == array_index_948883 ? add_970261 : sel_970258;
  assign add_970265 = sel_970262 + 8'h01;
  assign sel_970266 = array_index_969997 == array_index_948889 ? add_970265 : sel_970262;
  assign add_970269 = sel_970266 + 8'h01;
  assign sel_970270 = array_index_969997 == array_index_948895 ? add_970269 : sel_970266;
  assign add_970273 = sel_970270 + 8'h01;
  assign sel_970274 = array_index_969997 == array_index_948901 ? add_970273 : sel_970270;
  assign add_970277 = sel_970274 + 8'h01;
  assign sel_970278 = array_index_969997 == array_index_948907 ? add_970277 : sel_970274;
  assign add_970281 = sel_970278 + 8'h01;
  assign sel_970282 = array_index_969997 == array_index_948913 ? add_970281 : sel_970278;
  assign add_970285 = sel_970282 + 8'h01;
  assign sel_970286 = array_index_969997 == array_index_948919 ? add_970285 : sel_970282;
  assign add_970289 = sel_970286 + 8'h01;
  assign sel_970290 = array_index_969997 == array_index_948925 ? add_970289 : sel_970286;
  assign add_970293 = sel_970290 + 8'h01;
  assign sel_970294 = array_index_969997 == array_index_948931 ? add_970293 : sel_970290;
  assign add_970297 = sel_970294 + 8'h01;
  assign sel_970298 = array_index_969997 == array_index_948937 ? add_970297 : sel_970294;
  assign add_970301 = sel_970298 + 8'h01;
  assign sel_970302 = array_index_969997 == array_index_948943 ? add_970301 : sel_970298;
  assign add_970305 = sel_970302 + 8'h01;
  assign sel_970306 = array_index_969997 == array_index_948949 ? add_970305 : sel_970302;
  assign add_970309 = sel_970306 + 8'h01;
  assign sel_970310 = array_index_969997 == array_index_948955 ? add_970309 : sel_970306;
  assign add_970313 = sel_970310 + 8'h01;
  assign sel_970314 = array_index_969997 == array_index_948961 ? add_970313 : sel_970310;
  assign add_970317 = sel_970314 + 8'h01;
  assign sel_970318 = array_index_969997 == array_index_948967 ? add_970317 : sel_970314;
  assign add_970321 = sel_970318 + 8'h01;
  assign sel_970322 = array_index_969997 == array_index_948973 ? add_970321 : sel_970318;
  assign add_970325 = sel_970322 + 8'h01;
  assign sel_970326 = array_index_969997 == array_index_948979 ? add_970325 : sel_970322;
  assign add_970329 = sel_970326 + 8'h01;
  assign sel_970330 = array_index_969997 == array_index_948985 ? add_970329 : sel_970326;
  assign add_970333 = sel_970330 + 8'h01;
  assign sel_970334 = array_index_969997 == array_index_948991 ? add_970333 : sel_970330;
  assign add_970337 = sel_970334 + 8'h01;
  assign sel_970338 = array_index_969997 == array_index_948997 ? add_970337 : sel_970334;
  assign add_970341 = sel_970338 + 8'h01;
  assign sel_970342 = array_index_969997 == array_index_949003 ? add_970341 : sel_970338;
  assign add_970345 = sel_970342 + 8'h01;
  assign sel_970346 = array_index_969997 == array_index_949009 ? add_970345 : sel_970342;
  assign add_970349 = sel_970346 + 8'h01;
  assign sel_970350 = array_index_969997 == array_index_949015 ? add_970349 : sel_970346;
  assign add_970353 = sel_970350 + 8'h01;
  assign sel_970354 = array_index_969997 == array_index_949021 ? add_970353 : sel_970350;
  assign add_970357 = sel_970354 + 8'h01;
  assign sel_970358 = array_index_969997 == array_index_949027 ? add_970357 : sel_970354;
  assign add_970361 = sel_970358 + 8'h01;
  assign sel_970362 = array_index_969997 == array_index_949033 ? add_970361 : sel_970358;
  assign add_970365 = sel_970362 + 8'h01;
  assign sel_970366 = array_index_969997 == array_index_949039 ? add_970365 : sel_970362;
  assign add_970369 = sel_970366 + 8'h01;
  assign sel_970370 = array_index_969997 == array_index_949045 ? add_970369 : sel_970366;
  assign add_970373 = sel_970370 + 8'h01;
  assign sel_970374 = array_index_969997 == array_index_949051 ? add_970373 : sel_970370;
  assign add_970377 = sel_970374 + 8'h01;
  assign sel_970378 = array_index_969997 == array_index_949057 ? add_970377 : sel_970374;
  assign add_970381 = sel_970378 + 8'h01;
  assign sel_970382 = array_index_969997 == array_index_949063 ? add_970381 : sel_970378;
  assign add_970385 = sel_970382 + 8'h01;
  assign sel_970386 = array_index_969997 == array_index_949069 ? add_970385 : sel_970382;
  assign add_970389 = sel_970386 + 8'h01;
  assign sel_970390 = array_index_969997 == array_index_949075 ? add_970389 : sel_970386;
  assign add_970393 = sel_970390 + 8'h01;
  assign sel_970394 = array_index_969997 == array_index_949081 ? add_970393 : sel_970390;
  assign add_970398 = sel_970394 + 8'h01;
  assign array_index_970399 = set1_unflattened[7'h36];
  assign sel_970400 = array_index_969997 == array_index_949087 ? add_970398 : sel_970394;
  assign add_970403 = sel_970400 + 8'h01;
  assign sel_970404 = array_index_970399 == array_index_948483 ? add_970403 : sel_970400;
  assign add_970407 = sel_970404 + 8'h01;
  assign sel_970408 = array_index_970399 == array_index_948487 ? add_970407 : sel_970404;
  assign add_970411 = sel_970408 + 8'h01;
  assign sel_970412 = array_index_970399 == array_index_948495 ? add_970411 : sel_970408;
  assign add_970415 = sel_970412 + 8'h01;
  assign sel_970416 = array_index_970399 == array_index_948503 ? add_970415 : sel_970412;
  assign add_970419 = sel_970416 + 8'h01;
  assign sel_970420 = array_index_970399 == array_index_948511 ? add_970419 : sel_970416;
  assign add_970423 = sel_970420 + 8'h01;
  assign sel_970424 = array_index_970399 == array_index_948519 ? add_970423 : sel_970420;
  assign add_970427 = sel_970424 + 8'h01;
  assign sel_970428 = array_index_970399 == array_index_948527 ? add_970427 : sel_970424;
  assign add_970431 = sel_970428 + 8'h01;
  assign sel_970432 = array_index_970399 == array_index_948535 ? add_970431 : sel_970428;
  assign add_970435 = sel_970432 + 8'h01;
  assign sel_970436 = array_index_970399 == array_index_948541 ? add_970435 : sel_970432;
  assign add_970439 = sel_970436 + 8'h01;
  assign sel_970440 = array_index_970399 == array_index_948547 ? add_970439 : sel_970436;
  assign add_970443 = sel_970440 + 8'h01;
  assign sel_970444 = array_index_970399 == array_index_948553 ? add_970443 : sel_970440;
  assign add_970447 = sel_970444 + 8'h01;
  assign sel_970448 = array_index_970399 == array_index_948559 ? add_970447 : sel_970444;
  assign add_970451 = sel_970448 + 8'h01;
  assign sel_970452 = array_index_970399 == array_index_948565 ? add_970451 : sel_970448;
  assign add_970455 = sel_970452 + 8'h01;
  assign sel_970456 = array_index_970399 == array_index_948571 ? add_970455 : sel_970452;
  assign add_970459 = sel_970456 + 8'h01;
  assign sel_970460 = array_index_970399 == array_index_948577 ? add_970459 : sel_970456;
  assign add_970463 = sel_970460 + 8'h01;
  assign sel_970464 = array_index_970399 == array_index_948583 ? add_970463 : sel_970460;
  assign add_970467 = sel_970464 + 8'h01;
  assign sel_970468 = array_index_970399 == array_index_948589 ? add_970467 : sel_970464;
  assign add_970471 = sel_970468 + 8'h01;
  assign sel_970472 = array_index_970399 == array_index_948595 ? add_970471 : sel_970468;
  assign add_970475 = sel_970472 + 8'h01;
  assign sel_970476 = array_index_970399 == array_index_948601 ? add_970475 : sel_970472;
  assign add_970479 = sel_970476 + 8'h01;
  assign sel_970480 = array_index_970399 == array_index_948607 ? add_970479 : sel_970476;
  assign add_970483 = sel_970480 + 8'h01;
  assign sel_970484 = array_index_970399 == array_index_948613 ? add_970483 : sel_970480;
  assign add_970487 = sel_970484 + 8'h01;
  assign sel_970488 = array_index_970399 == array_index_948619 ? add_970487 : sel_970484;
  assign add_970491 = sel_970488 + 8'h01;
  assign sel_970492 = array_index_970399 == array_index_948625 ? add_970491 : sel_970488;
  assign add_970495 = sel_970492 + 8'h01;
  assign sel_970496 = array_index_970399 == array_index_948631 ? add_970495 : sel_970492;
  assign add_970499 = sel_970496 + 8'h01;
  assign sel_970500 = array_index_970399 == array_index_948637 ? add_970499 : sel_970496;
  assign add_970503 = sel_970500 + 8'h01;
  assign sel_970504 = array_index_970399 == array_index_948643 ? add_970503 : sel_970500;
  assign add_970507 = sel_970504 + 8'h01;
  assign sel_970508 = array_index_970399 == array_index_948649 ? add_970507 : sel_970504;
  assign add_970511 = sel_970508 + 8'h01;
  assign sel_970512 = array_index_970399 == array_index_948655 ? add_970511 : sel_970508;
  assign add_970515 = sel_970512 + 8'h01;
  assign sel_970516 = array_index_970399 == array_index_948661 ? add_970515 : sel_970512;
  assign add_970519 = sel_970516 + 8'h01;
  assign sel_970520 = array_index_970399 == array_index_948667 ? add_970519 : sel_970516;
  assign add_970523 = sel_970520 + 8'h01;
  assign sel_970524 = array_index_970399 == array_index_948673 ? add_970523 : sel_970520;
  assign add_970527 = sel_970524 + 8'h01;
  assign sel_970528 = array_index_970399 == array_index_948679 ? add_970527 : sel_970524;
  assign add_970531 = sel_970528 + 8'h01;
  assign sel_970532 = array_index_970399 == array_index_948685 ? add_970531 : sel_970528;
  assign add_970535 = sel_970532 + 8'h01;
  assign sel_970536 = array_index_970399 == array_index_948691 ? add_970535 : sel_970532;
  assign add_970539 = sel_970536 + 8'h01;
  assign sel_970540 = array_index_970399 == array_index_948697 ? add_970539 : sel_970536;
  assign add_970543 = sel_970540 + 8'h01;
  assign sel_970544 = array_index_970399 == array_index_948703 ? add_970543 : sel_970540;
  assign add_970547 = sel_970544 + 8'h01;
  assign sel_970548 = array_index_970399 == array_index_948709 ? add_970547 : sel_970544;
  assign add_970551 = sel_970548 + 8'h01;
  assign sel_970552 = array_index_970399 == array_index_948715 ? add_970551 : sel_970548;
  assign add_970555 = sel_970552 + 8'h01;
  assign sel_970556 = array_index_970399 == array_index_948721 ? add_970555 : sel_970552;
  assign add_970559 = sel_970556 + 8'h01;
  assign sel_970560 = array_index_970399 == array_index_948727 ? add_970559 : sel_970556;
  assign add_970563 = sel_970560 + 8'h01;
  assign sel_970564 = array_index_970399 == array_index_948733 ? add_970563 : sel_970560;
  assign add_970567 = sel_970564 + 8'h01;
  assign sel_970568 = array_index_970399 == array_index_948739 ? add_970567 : sel_970564;
  assign add_970571 = sel_970568 + 8'h01;
  assign sel_970572 = array_index_970399 == array_index_948745 ? add_970571 : sel_970568;
  assign add_970575 = sel_970572 + 8'h01;
  assign sel_970576 = array_index_970399 == array_index_948751 ? add_970575 : sel_970572;
  assign add_970579 = sel_970576 + 8'h01;
  assign sel_970580 = array_index_970399 == array_index_948757 ? add_970579 : sel_970576;
  assign add_970583 = sel_970580 + 8'h01;
  assign sel_970584 = array_index_970399 == array_index_948763 ? add_970583 : sel_970580;
  assign add_970587 = sel_970584 + 8'h01;
  assign sel_970588 = array_index_970399 == array_index_948769 ? add_970587 : sel_970584;
  assign add_970591 = sel_970588 + 8'h01;
  assign sel_970592 = array_index_970399 == array_index_948775 ? add_970591 : sel_970588;
  assign add_970595 = sel_970592 + 8'h01;
  assign sel_970596 = array_index_970399 == array_index_948781 ? add_970595 : sel_970592;
  assign add_970599 = sel_970596 + 8'h01;
  assign sel_970600 = array_index_970399 == array_index_948787 ? add_970599 : sel_970596;
  assign add_970603 = sel_970600 + 8'h01;
  assign sel_970604 = array_index_970399 == array_index_948793 ? add_970603 : sel_970600;
  assign add_970607 = sel_970604 + 8'h01;
  assign sel_970608 = array_index_970399 == array_index_948799 ? add_970607 : sel_970604;
  assign add_970611 = sel_970608 + 8'h01;
  assign sel_970612 = array_index_970399 == array_index_948805 ? add_970611 : sel_970608;
  assign add_970615 = sel_970612 + 8'h01;
  assign sel_970616 = array_index_970399 == array_index_948811 ? add_970615 : sel_970612;
  assign add_970619 = sel_970616 + 8'h01;
  assign sel_970620 = array_index_970399 == array_index_948817 ? add_970619 : sel_970616;
  assign add_970623 = sel_970620 + 8'h01;
  assign sel_970624 = array_index_970399 == array_index_948823 ? add_970623 : sel_970620;
  assign add_970627 = sel_970624 + 8'h01;
  assign sel_970628 = array_index_970399 == array_index_948829 ? add_970627 : sel_970624;
  assign add_970631 = sel_970628 + 8'h01;
  assign sel_970632 = array_index_970399 == array_index_948835 ? add_970631 : sel_970628;
  assign add_970635 = sel_970632 + 8'h01;
  assign sel_970636 = array_index_970399 == array_index_948841 ? add_970635 : sel_970632;
  assign add_970639 = sel_970636 + 8'h01;
  assign sel_970640 = array_index_970399 == array_index_948847 ? add_970639 : sel_970636;
  assign add_970643 = sel_970640 + 8'h01;
  assign sel_970644 = array_index_970399 == array_index_948853 ? add_970643 : sel_970640;
  assign add_970647 = sel_970644 + 8'h01;
  assign sel_970648 = array_index_970399 == array_index_948859 ? add_970647 : sel_970644;
  assign add_970651 = sel_970648 + 8'h01;
  assign sel_970652 = array_index_970399 == array_index_948865 ? add_970651 : sel_970648;
  assign add_970655 = sel_970652 + 8'h01;
  assign sel_970656 = array_index_970399 == array_index_948871 ? add_970655 : sel_970652;
  assign add_970659 = sel_970656 + 8'h01;
  assign sel_970660 = array_index_970399 == array_index_948877 ? add_970659 : sel_970656;
  assign add_970663 = sel_970660 + 8'h01;
  assign sel_970664 = array_index_970399 == array_index_948883 ? add_970663 : sel_970660;
  assign add_970667 = sel_970664 + 8'h01;
  assign sel_970668 = array_index_970399 == array_index_948889 ? add_970667 : sel_970664;
  assign add_970671 = sel_970668 + 8'h01;
  assign sel_970672 = array_index_970399 == array_index_948895 ? add_970671 : sel_970668;
  assign add_970675 = sel_970672 + 8'h01;
  assign sel_970676 = array_index_970399 == array_index_948901 ? add_970675 : sel_970672;
  assign add_970679 = sel_970676 + 8'h01;
  assign sel_970680 = array_index_970399 == array_index_948907 ? add_970679 : sel_970676;
  assign add_970683 = sel_970680 + 8'h01;
  assign sel_970684 = array_index_970399 == array_index_948913 ? add_970683 : sel_970680;
  assign add_970687 = sel_970684 + 8'h01;
  assign sel_970688 = array_index_970399 == array_index_948919 ? add_970687 : sel_970684;
  assign add_970691 = sel_970688 + 8'h01;
  assign sel_970692 = array_index_970399 == array_index_948925 ? add_970691 : sel_970688;
  assign add_970695 = sel_970692 + 8'h01;
  assign sel_970696 = array_index_970399 == array_index_948931 ? add_970695 : sel_970692;
  assign add_970699 = sel_970696 + 8'h01;
  assign sel_970700 = array_index_970399 == array_index_948937 ? add_970699 : sel_970696;
  assign add_970703 = sel_970700 + 8'h01;
  assign sel_970704 = array_index_970399 == array_index_948943 ? add_970703 : sel_970700;
  assign add_970707 = sel_970704 + 8'h01;
  assign sel_970708 = array_index_970399 == array_index_948949 ? add_970707 : sel_970704;
  assign add_970711 = sel_970708 + 8'h01;
  assign sel_970712 = array_index_970399 == array_index_948955 ? add_970711 : sel_970708;
  assign add_970715 = sel_970712 + 8'h01;
  assign sel_970716 = array_index_970399 == array_index_948961 ? add_970715 : sel_970712;
  assign add_970719 = sel_970716 + 8'h01;
  assign sel_970720 = array_index_970399 == array_index_948967 ? add_970719 : sel_970716;
  assign add_970723 = sel_970720 + 8'h01;
  assign sel_970724 = array_index_970399 == array_index_948973 ? add_970723 : sel_970720;
  assign add_970727 = sel_970724 + 8'h01;
  assign sel_970728 = array_index_970399 == array_index_948979 ? add_970727 : sel_970724;
  assign add_970731 = sel_970728 + 8'h01;
  assign sel_970732 = array_index_970399 == array_index_948985 ? add_970731 : sel_970728;
  assign add_970735 = sel_970732 + 8'h01;
  assign sel_970736 = array_index_970399 == array_index_948991 ? add_970735 : sel_970732;
  assign add_970739 = sel_970736 + 8'h01;
  assign sel_970740 = array_index_970399 == array_index_948997 ? add_970739 : sel_970736;
  assign add_970743 = sel_970740 + 8'h01;
  assign sel_970744 = array_index_970399 == array_index_949003 ? add_970743 : sel_970740;
  assign add_970747 = sel_970744 + 8'h01;
  assign sel_970748 = array_index_970399 == array_index_949009 ? add_970747 : sel_970744;
  assign add_970751 = sel_970748 + 8'h01;
  assign sel_970752 = array_index_970399 == array_index_949015 ? add_970751 : sel_970748;
  assign add_970755 = sel_970752 + 8'h01;
  assign sel_970756 = array_index_970399 == array_index_949021 ? add_970755 : sel_970752;
  assign add_970759 = sel_970756 + 8'h01;
  assign sel_970760 = array_index_970399 == array_index_949027 ? add_970759 : sel_970756;
  assign add_970763 = sel_970760 + 8'h01;
  assign sel_970764 = array_index_970399 == array_index_949033 ? add_970763 : sel_970760;
  assign add_970767 = sel_970764 + 8'h01;
  assign sel_970768 = array_index_970399 == array_index_949039 ? add_970767 : sel_970764;
  assign add_970771 = sel_970768 + 8'h01;
  assign sel_970772 = array_index_970399 == array_index_949045 ? add_970771 : sel_970768;
  assign add_970775 = sel_970772 + 8'h01;
  assign sel_970776 = array_index_970399 == array_index_949051 ? add_970775 : sel_970772;
  assign add_970779 = sel_970776 + 8'h01;
  assign sel_970780 = array_index_970399 == array_index_949057 ? add_970779 : sel_970776;
  assign add_970783 = sel_970780 + 8'h01;
  assign sel_970784 = array_index_970399 == array_index_949063 ? add_970783 : sel_970780;
  assign add_970787 = sel_970784 + 8'h01;
  assign sel_970788 = array_index_970399 == array_index_949069 ? add_970787 : sel_970784;
  assign add_970791 = sel_970788 + 8'h01;
  assign sel_970792 = array_index_970399 == array_index_949075 ? add_970791 : sel_970788;
  assign add_970795 = sel_970792 + 8'h01;
  assign sel_970796 = array_index_970399 == array_index_949081 ? add_970795 : sel_970792;
  assign add_970800 = sel_970796 + 8'h01;
  assign array_index_970801 = set1_unflattened[7'h37];
  assign sel_970802 = array_index_970399 == array_index_949087 ? add_970800 : sel_970796;
  assign add_970805 = sel_970802 + 8'h01;
  assign sel_970806 = array_index_970801 == array_index_948483 ? add_970805 : sel_970802;
  assign add_970809 = sel_970806 + 8'h01;
  assign sel_970810 = array_index_970801 == array_index_948487 ? add_970809 : sel_970806;
  assign add_970813 = sel_970810 + 8'h01;
  assign sel_970814 = array_index_970801 == array_index_948495 ? add_970813 : sel_970810;
  assign add_970817 = sel_970814 + 8'h01;
  assign sel_970818 = array_index_970801 == array_index_948503 ? add_970817 : sel_970814;
  assign add_970821 = sel_970818 + 8'h01;
  assign sel_970822 = array_index_970801 == array_index_948511 ? add_970821 : sel_970818;
  assign add_970825 = sel_970822 + 8'h01;
  assign sel_970826 = array_index_970801 == array_index_948519 ? add_970825 : sel_970822;
  assign add_970829 = sel_970826 + 8'h01;
  assign sel_970830 = array_index_970801 == array_index_948527 ? add_970829 : sel_970826;
  assign add_970833 = sel_970830 + 8'h01;
  assign sel_970834 = array_index_970801 == array_index_948535 ? add_970833 : sel_970830;
  assign add_970837 = sel_970834 + 8'h01;
  assign sel_970838 = array_index_970801 == array_index_948541 ? add_970837 : sel_970834;
  assign add_970841 = sel_970838 + 8'h01;
  assign sel_970842 = array_index_970801 == array_index_948547 ? add_970841 : sel_970838;
  assign add_970845 = sel_970842 + 8'h01;
  assign sel_970846 = array_index_970801 == array_index_948553 ? add_970845 : sel_970842;
  assign add_970849 = sel_970846 + 8'h01;
  assign sel_970850 = array_index_970801 == array_index_948559 ? add_970849 : sel_970846;
  assign add_970853 = sel_970850 + 8'h01;
  assign sel_970854 = array_index_970801 == array_index_948565 ? add_970853 : sel_970850;
  assign add_970857 = sel_970854 + 8'h01;
  assign sel_970858 = array_index_970801 == array_index_948571 ? add_970857 : sel_970854;
  assign add_970861 = sel_970858 + 8'h01;
  assign sel_970862 = array_index_970801 == array_index_948577 ? add_970861 : sel_970858;
  assign add_970865 = sel_970862 + 8'h01;
  assign sel_970866 = array_index_970801 == array_index_948583 ? add_970865 : sel_970862;
  assign add_970869 = sel_970866 + 8'h01;
  assign sel_970870 = array_index_970801 == array_index_948589 ? add_970869 : sel_970866;
  assign add_970873 = sel_970870 + 8'h01;
  assign sel_970874 = array_index_970801 == array_index_948595 ? add_970873 : sel_970870;
  assign add_970877 = sel_970874 + 8'h01;
  assign sel_970878 = array_index_970801 == array_index_948601 ? add_970877 : sel_970874;
  assign add_970881 = sel_970878 + 8'h01;
  assign sel_970882 = array_index_970801 == array_index_948607 ? add_970881 : sel_970878;
  assign add_970885 = sel_970882 + 8'h01;
  assign sel_970886 = array_index_970801 == array_index_948613 ? add_970885 : sel_970882;
  assign add_970889 = sel_970886 + 8'h01;
  assign sel_970890 = array_index_970801 == array_index_948619 ? add_970889 : sel_970886;
  assign add_970893 = sel_970890 + 8'h01;
  assign sel_970894 = array_index_970801 == array_index_948625 ? add_970893 : sel_970890;
  assign add_970897 = sel_970894 + 8'h01;
  assign sel_970898 = array_index_970801 == array_index_948631 ? add_970897 : sel_970894;
  assign add_970901 = sel_970898 + 8'h01;
  assign sel_970902 = array_index_970801 == array_index_948637 ? add_970901 : sel_970898;
  assign add_970905 = sel_970902 + 8'h01;
  assign sel_970906 = array_index_970801 == array_index_948643 ? add_970905 : sel_970902;
  assign add_970909 = sel_970906 + 8'h01;
  assign sel_970910 = array_index_970801 == array_index_948649 ? add_970909 : sel_970906;
  assign add_970913 = sel_970910 + 8'h01;
  assign sel_970914 = array_index_970801 == array_index_948655 ? add_970913 : sel_970910;
  assign add_970917 = sel_970914 + 8'h01;
  assign sel_970918 = array_index_970801 == array_index_948661 ? add_970917 : sel_970914;
  assign add_970921 = sel_970918 + 8'h01;
  assign sel_970922 = array_index_970801 == array_index_948667 ? add_970921 : sel_970918;
  assign add_970925 = sel_970922 + 8'h01;
  assign sel_970926 = array_index_970801 == array_index_948673 ? add_970925 : sel_970922;
  assign add_970929 = sel_970926 + 8'h01;
  assign sel_970930 = array_index_970801 == array_index_948679 ? add_970929 : sel_970926;
  assign add_970933 = sel_970930 + 8'h01;
  assign sel_970934 = array_index_970801 == array_index_948685 ? add_970933 : sel_970930;
  assign add_970937 = sel_970934 + 8'h01;
  assign sel_970938 = array_index_970801 == array_index_948691 ? add_970937 : sel_970934;
  assign add_970941 = sel_970938 + 8'h01;
  assign sel_970942 = array_index_970801 == array_index_948697 ? add_970941 : sel_970938;
  assign add_970945 = sel_970942 + 8'h01;
  assign sel_970946 = array_index_970801 == array_index_948703 ? add_970945 : sel_970942;
  assign add_970949 = sel_970946 + 8'h01;
  assign sel_970950 = array_index_970801 == array_index_948709 ? add_970949 : sel_970946;
  assign add_970953 = sel_970950 + 8'h01;
  assign sel_970954 = array_index_970801 == array_index_948715 ? add_970953 : sel_970950;
  assign add_970957 = sel_970954 + 8'h01;
  assign sel_970958 = array_index_970801 == array_index_948721 ? add_970957 : sel_970954;
  assign add_970961 = sel_970958 + 8'h01;
  assign sel_970962 = array_index_970801 == array_index_948727 ? add_970961 : sel_970958;
  assign add_970965 = sel_970962 + 8'h01;
  assign sel_970966 = array_index_970801 == array_index_948733 ? add_970965 : sel_970962;
  assign add_970969 = sel_970966 + 8'h01;
  assign sel_970970 = array_index_970801 == array_index_948739 ? add_970969 : sel_970966;
  assign add_970973 = sel_970970 + 8'h01;
  assign sel_970974 = array_index_970801 == array_index_948745 ? add_970973 : sel_970970;
  assign add_970977 = sel_970974 + 8'h01;
  assign sel_970978 = array_index_970801 == array_index_948751 ? add_970977 : sel_970974;
  assign add_970981 = sel_970978 + 8'h01;
  assign sel_970982 = array_index_970801 == array_index_948757 ? add_970981 : sel_970978;
  assign add_970985 = sel_970982 + 8'h01;
  assign sel_970986 = array_index_970801 == array_index_948763 ? add_970985 : sel_970982;
  assign add_970989 = sel_970986 + 8'h01;
  assign sel_970990 = array_index_970801 == array_index_948769 ? add_970989 : sel_970986;
  assign add_970993 = sel_970990 + 8'h01;
  assign sel_970994 = array_index_970801 == array_index_948775 ? add_970993 : sel_970990;
  assign add_970997 = sel_970994 + 8'h01;
  assign sel_970998 = array_index_970801 == array_index_948781 ? add_970997 : sel_970994;
  assign add_971001 = sel_970998 + 8'h01;
  assign sel_971002 = array_index_970801 == array_index_948787 ? add_971001 : sel_970998;
  assign add_971005 = sel_971002 + 8'h01;
  assign sel_971006 = array_index_970801 == array_index_948793 ? add_971005 : sel_971002;
  assign add_971009 = sel_971006 + 8'h01;
  assign sel_971010 = array_index_970801 == array_index_948799 ? add_971009 : sel_971006;
  assign add_971013 = sel_971010 + 8'h01;
  assign sel_971014 = array_index_970801 == array_index_948805 ? add_971013 : sel_971010;
  assign add_971017 = sel_971014 + 8'h01;
  assign sel_971018 = array_index_970801 == array_index_948811 ? add_971017 : sel_971014;
  assign add_971021 = sel_971018 + 8'h01;
  assign sel_971022 = array_index_970801 == array_index_948817 ? add_971021 : sel_971018;
  assign add_971025 = sel_971022 + 8'h01;
  assign sel_971026 = array_index_970801 == array_index_948823 ? add_971025 : sel_971022;
  assign add_971029 = sel_971026 + 8'h01;
  assign sel_971030 = array_index_970801 == array_index_948829 ? add_971029 : sel_971026;
  assign add_971033 = sel_971030 + 8'h01;
  assign sel_971034 = array_index_970801 == array_index_948835 ? add_971033 : sel_971030;
  assign add_971037 = sel_971034 + 8'h01;
  assign sel_971038 = array_index_970801 == array_index_948841 ? add_971037 : sel_971034;
  assign add_971041 = sel_971038 + 8'h01;
  assign sel_971042 = array_index_970801 == array_index_948847 ? add_971041 : sel_971038;
  assign add_971045 = sel_971042 + 8'h01;
  assign sel_971046 = array_index_970801 == array_index_948853 ? add_971045 : sel_971042;
  assign add_971049 = sel_971046 + 8'h01;
  assign sel_971050 = array_index_970801 == array_index_948859 ? add_971049 : sel_971046;
  assign add_971053 = sel_971050 + 8'h01;
  assign sel_971054 = array_index_970801 == array_index_948865 ? add_971053 : sel_971050;
  assign add_971057 = sel_971054 + 8'h01;
  assign sel_971058 = array_index_970801 == array_index_948871 ? add_971057 : sel_971054;
  assign add_971061 = sel_971058 + 8'h01;
  assign sel_971062 = array_index_970801 == array_index_948877 ? add_971061 : sel_971058;
  assign add_971065 = sel_971062 + 8'h01;
  assign sel_971066 = array_index_970801 == array_index_948883 ? add_971065 : sel_971062;
  assign add_971069 = sel_971066 + 8'h01;
  assign sel_971070 = array_index_970801 == array_index_948889 ? add_971069 : sel_971066;
  assign add_971073 = sel_971070 + 8'h01;
  assign sel_971074 = array_index_970801 == array_index_948895 ? add_971073 : sel_971070;
  assign add_971077 = sel_971074 + 8'h01;
  assign sel_971078 = array_index_970801 == array_index_948901 ? add_971077 : sel_971074;
  assign add_971081 = sel_971078 + 8'h01;
  assign sel_971082 = array_index_970801 == array_index_948907 ? add_971081 : sel_971078;
  assign add_971085 = sel_971082 + 8'h01;
  assign sel_971086 = array_index_970801 == array_index_948913 ? add_971085 : sel_971082;
  assign add_971089 = sel_971086 + 8'h01;
  assign sel_971090 = array_index_970801 == array_index_948919 ? add_971089 : sel_971086;
  assign add_971093 = sel_971090 + 8'h01;
  assign sel_971094 = array_index_970801 == array_index_948925 ? add_971093 : sel_971090;
  assign add_971097 = sel_971094 + 8'h01;
  assign sel_971098 = array_index_970801 == array_index_948931 ? add_971097 : sel_971094;
  assign add_971101 = sel_971098 + 8'h01;
  assign sel_971102 = array_index_970801 == array_index_948937 ? add_971101 : sel_971098;
  assign add_971105 = sel_971102 + 8'h01;
  assign sel_971106 = array_index_970801 == array_index_948943 ? add_971105 : sel_971102;
  assign add_971109 = sel_971106 + 8'h01;
  assign sel_971110 = array_index_970801 == array_index_948949 ? add_971109 : sel_971106;
  assign add_971113 = sel_971110 + 8'h01;
  assign sel_971114 = array_index_970801 == array_index_948955 ? add_971113 : sel_971110;
  assign add_971117 = sel_971114 + 8'h01;
  assign sel_971118 = array_index_970801 == array_index_948961 ? add_971117 : sel_971114;
  assign add_971121 = sel_971118 + 8'h01;
  assign sel_971122 = array_index_970801 == array_index_948967 ? add_971121 : sel_971118;
  assign add_971125 = sel_971122 + 8'h01;
  assign sel_971126 = array_index_970801 == array_index_948973 ? add_971125 : sel_971122;
  assign add_971129 = sel_971126 + 8'h01;
  assign sel_971130 = array_index_970801 == array_index_948979 ? add_971129 : sel_971126;
  assign add_971133 = sel_971130 + 8'h01;
  assign sel_971134 = array_index_970801 == array_index_948985 ? add_971133 : sel_971130;
  assign add_971137 = sel_971134 + 8'h01;
  assign sel_971138 = array_index_970801 == array_index_948991 ? add_971137 : sel_971134;
  assign add_971141 = sel_971138 + 8'h01;
  assign sel_971142 = array_index_970801 == array_index_948997 ? add_971141 : sel_971138;
  assign add_971145 = sel_971142 + 8'h01;
  assign sel_971146 = array_index_970801 == array_index_949003 ? add_971145 : sel_971142;
  assign add_971149 = sel_971146 + 8'h01;
  assign sel_971150 = array_index_970801 == array_index_949009 ? add_971149 : sel_971146;
  assign add_971153 = sel_971150 + 8'h01;
  assign sel_971154 = array_index_970801 == array_index_949015 ? add_971153 : sel_971150;
  assign add_971157 = sel_971154 + 8'h01;
  assign sel_971158 = array_index_970801 == array_index_949021 ? add_971157 : sel_971154;
  assign add_971161 = sel_971158 + 8'h01;
  assign sel_971162 = array_index_970801 == array_index_949027 ? add_971161 : sel_971158;
  assign add_971165 = sel_971162 + 8'h01;
  assign sel_971166 = array_index_970801 == array_index_949033 ? add_971165 : sel_971162;
  assign add_971169 = sel_971166 + 8'h01;
  assign sel_971170 = array_index_970801 == array_index_949039 ? add_971169 : sel_971166;
  assign add_971173 = sel_971170 + 8'h01;
  assign sel_971174 = array_index_970801 == array_index_949045 ? add_971173 : sel_971170;
  assign add_971177 = sel_971174 + 8'h01;
  assign sel_971178 = array_index_970801 == array_index_949051 ? add_971177 : sel_971174;
  assign add_971181 = sel_971178 + 8'h01;
  assign sel_971182 = array_index_970801 == array_index_949057 ? add_971181 : sel_971178;
  assign add_971185 = sel_971182 + 8'h01;
  assign sel_971186 = array_index_970801 == array_index_949063 ? add_971185 : sel_971182;
  assign add_971189 = sel_971186 + 8'h01;
  assign sel_971190 = array_index_970801 == array_index_949069 ? add_971189 : sel_971186;
  assign add_971193 = sel_971190 + 8'h01;
  assign sel_971194 = array_index_970801 == array_index_949075 ? add_971193 : sel_971190;
  assign add_971197 = sel_971194 + 8'h01;
  assign sel_971198 = array_index_970801 == array_index_949081 ? add_971197 : sel_971194;
  assign add_971202 = sel_971198 + 8'h01;
  assign array_index_971203 = set1_unflattened[7'h38];
  assign sel_971204 = array_index_970801 == array_index_949087 ? add_971202 : sel_971198;
  assign add_971207 = sel_971204 + 8'h01;
  assign sel_971208 = array_index_971203 == array_index_948483 ? add_971207 : sel_971204;
  assign add_971211 = sel_971208 + 8'h01;
  assign sel_971212 = array_index_971203 == array_index_948487 ? add_971211 : sel_971208;
  assign add_971215 = sel_971212 + 8'h01;
  assign sel_971216 = array_index_971203 == array_index_948495 ? add_971215 : sel_971212;
  assign add_971219 = sel_971216 + 8'h01;
  assign sel_971220 = array_index_971203 == array_index_948503 ? add_971219 : sel_971216;
  assign add_971223 = sel_971220 + 8'h01;
  assign sel_971224 = array_index_971203 == array_index_948511 ? add_971223 : sel_971220;
  assign add_971227 = sel_971224 + 8'h01;
  assign sel_971228 = array_index_971203 == array_index_948519 ? add_971227 : sel_971224;
  assign add_971231 = sel_971228 + 8'h01;
  assign sel_971232 = array_index_971203 == array_index_948527 ? add_971231 : sel_971228;
  assign add_971235 = sel_971232 + 8'h01;
  assign sel_971236 = array_index_971203 == array_index_948535 ? add_971235 : sel_971232;
  assign add_971239 = sel_971236 + 8'h01;
  assign sel_971240 = array_index_971203 == array_index_948541 ? add_971239 : sel_971236;
  assign add_971243 = sel_971240 + 8'h01;
  assign sel_971244 = array_index_971203 == array_index_948547 ? add_971243 : sel_971240;
  assign add_971247 = sel_971244 + 8'h01;
  assign sel_971248 = array_index_971203 == array_index_948553 ? add_971247 : sel_971244;
  assign add_971251 = sel_971248 + 8'h01;
  assign sel_971252 = array_index_971203 == array_index_948559 ? add_971251 : sel_971248;
  assign add_971255 = sel_971252 + 8'h01;
  assign sel_971256 = array_index_971203 == array_index_948565 ? add_971255 : sel_971252;
  assign add_971259 = sel_971256 + 8'h01;
  assign sel_971260 = array_index_971203 == array_index_948571 ? add_971259 : sel_971256;
  assign add_971263 = sel_971260 + 8'h01;
  assign sel_971264 = array_index_971203 == array_index_948577 ? add_971263 : sel_971260;
  assign add_971267 = sel_971264 + 8'h01;
  assign sel_971268 = array_index_971203 == array_index_948583 ? add_971267 : sel_971264;
  assign add_971271 = sel_971268 + 8'h01;
  assign sel_971272 = array_index_971203 == array_index_948589 ? add_971271 : sel_971268;
  assign add_971275 = sel_971272 + 8'h01;
  assign sel_971276 = array_index_971203 == array_index_948595 ? add_971275 : sel_971272;
  assign add_971279 = sel_971276 + 8'h01;
  assign sel_971280 = array_index_971203 == array_index_948601 ? add_971279 : sel_971276;
  assign add_971283 = sel_971280 + 8'h01;
  assign sel_971284 = array_index_971203 == array_index_948607 ? add_971283 : sel_971280;
  assign add_971287 = sel_971284 + 8'h01;
  assign sel_971288 = array_index_971203 == array_index_948613 ? add_971287 : sel_971284;
  assign add_971291 = sel_971288 + 8'h01;
  assign sel_971292 = array_index_971203 == array_index_948619 ? add_971291 : sel_971288;
  assign add_971295 = sel_971292 + 8'h01;
  assign sel_971296 = array_index_971203 == array_index_948625 ? add_971295 : sel_971292;
  assign add_971299 = sel_971296 + 8'h01;
  assign sel_971300 = array_index_971203 == array_index_948631 ? add_971299 : sel_971296;
  assign add_971303 = sel_971300 + 8'h01;
  assign sel_971304 = array_index_971203 == array_index_948637 ? add_971303 : sel_971300;
  assign add_971307 = sel_971304 + 8'h01;
  assign sel_971308 = array_index_971203 == array_index_948643 ? add_971307 : sel_971304;
  assign add_971311 = sel_971308 + 8'h01;
  assign sel_971312 = array_index_971203 == array_index_948649 ? add_971311 : sel_971308;
  assign add_971315 = sel_971312 + 8'h01;
  assign sel_971316 = array_index_971203 == array_index_948655 ? add_971315 : sel_971312;
  assign add_971319 = sel_971316 + 8'h01;
  assign sel_971320 = array_index_971203 == array_index_948661 ? add_971319 : sel_971316;
  assign add_971323 = sel_971320 + 8'h01;
  assign sel_971324 = array_index_971203 == array_index_948667 ? add_971323 : sel_971320;
  assign add_971327 = sel_971324 + 8'h01;
  assign sel_971328 = array_index_971203 == array_index_948673 ? add_971327 : sel_971324;
  assign add_971331 = sel_971328 + 8'h01;
  assign sel_971332 = array_index_971203 == array_index_948679 ? add_971331 : sel_971328;
  assign add_971335 = sel_971332 + 8'h01;
  assign sel_971336 = array_index_971203 == array_index_948685 ? add_971335 : sel_971332;
  assign add_971339 = sel_971336 + 8'h01;
  assign sel_971340 = array_index_971203 == array_index_948691 ? add_971339 : sel_971336;
  assign add_971343 = sel_971340 + 8'h01;
  assign sel_971344 = array_index_971203 == array_index_948697 ? add_971343 : sel_971340;
  assign add_971347 = sel_971344 + 8'h01;
  assign sel_971348 = array_index_971203 == array_index_948703 ? add_971347 : sel_971344;
  assign add_971351 = sel_971348 + 8'h01;
  assign sel_971352 = array_index_971203 == array_index_948709 ? add_971351 : sel_971348;
  assign add_971355 = sel_971352 + 8'h01;
  assign sel_971356 = array_index_971203 == array_index_948715 ? add_971355 : sel_971352;
  assign add_971359 = sel_971356 + 8'h01;
  assign sel_971360 = array_index_971203 == array_index_948721 ? add_971359 : sel_971356;
  assign add_971363 = sel_971360 + 8'h01;
  assign sel_971364 = array_index_971203 == array_index_948727 ? add_971363 : sel_971360;
  assign add_971367 = sel_971364 + 8'h01;
  assign sel_971368 = array_index_971203 == array_index_948733 ? add_971367 : sel_971364;
  assign add_971371 = sel_971368 + 8'h01;
  assign sel_971372 = array_index_971203 == array_index_948739 ? add_971371 : sel_971368;
  assign add_971375 = sel_971372 + 8'h01;
  assign sel_971376 = array_index_971203 == array_index_948745 ? add_971375 : sel_971372;
  assign add_971379 = sel_971376 + 8'h01;
  assign sel_971380 = array_index_971203 == array_index_948751 ? add_971379 : sel_971376;
  assign add_971383 = sel_971380 + 8'h01;
  assign sel_971384 = array_index_971203 == array_index_948757 ? add_971383 : sel_971380;
  assign add_971387 = sel_971384 + 8'h01;
  assign sel_971388 = array_index_971203 == array_index_948763 ? add_971387 : sel_971384;
  assign add_971391 = sel_971388 + 8'h01;
  assign sel_971392 = array_index_971203 == array_index_948769 ? add_971391 : sel_971388;
  assign add_971395 = sel_971392 + 8'h01;
  assign sel_971396 = array_index_971203 == array_index_948775 ? add_971395 : sel_971392;
  assign add_971399 = sel_971396 + 8'h01;
  assign sel_971400 = array_index_971203 == array_index_948781 ? add_971399 : sel_971396;
  assign add_971403 = sel_971400 + 8'h01;
  assign sel_971404 = array_index_971203 == array_index_948787 ? add_971403 : sel_971400;
  assign add_971407 = sel_971404 + 8'h01;
  assign sel_971408 = array_index_971203 == array_index_948793 ? add_971407 : sel_971404;
  assign add_971411 = sel_971408 + 8'h01;
  assign sel_971412 = array_index_971203 == array_index_948799 ? add_971411 : sel_971408;
  assign add_971415 = sel_971412 + 8'h01;
  assign sel_971416 = array_index_971203 == array_index_948805 ? add_971415 : sel_971412;
  assign add_971419 = sel_971416 + 8'h01;
  assign sel_971420 = array_index_971203 == array_index_948811 ? add_971419 : sel_971416;
  assign add_971423 = sel_971420 + 8'h01;
  assign sel_971424 = array_index_971203 == array_index_948817 ? add_971423 : sel_971420;
  assign add_971427 = sel_971424 + 8'h01;
  assign sel_971428 = array_index_971203 == array_index_948823 ? add_971427 : sel_971424;
  assign add_971431 = sel_971428 + 8'h01;
  assign sel_971432 = array_index_971203 == array_index_948829 ? add_971431 : sel_971428;
  assign add_971435 = sel_971432 + 8'h01;
  assign sel_971436 = array_index_971203 == array_index_948835 ? add_971435 : sel_971432;
  assign add_971439 = sel_971436 + 8'h01;
  assign sel_971440 = array_index_971203 == array_index_948841 ? add_971439 : sel_971436;
  assign add_971443 = sel_971440 + 8'h01;
  assign sel_971444 = array_index_971203 == array_index_948847 ? add_971443 : sel_971440;
  assign add_971447 = sel_971444 + 8'h01;
  assign sel_971448 = array_index_971203 == array_index_948853 ? add_971447 : sel_971444;
  assign add_971451 = sel_971448 + 8'h01;
  assign sel_971452 = array_index_971203 == array_index_948859 ? add_971451 : sel_971448;
  assign add_971455 = sel_971452 + 8'h01;
  assign sel_971456 = array_index_971203 == array_index_948865 ? add_971455 : sel_971452;
  assign add_971459 = sel_971456 + 8'h01;
  assign sel_971460 = array_index_971203 == array_index_948871 ? add_971459 : sel_971456;
  assign add_971463 = sel_971460 + 8'h01;
  assign sel_971464 = array_index_971203 == array_index_948877 ? add_971463 : sel_971460;
  assign add_971467 = sel_971464 + 8'h01;
  assign sel_971468 = array_index_971203 == array_index_948883 ? add_971467 : sel_971464;
  assign add_971471 = sel_971468 + 8'h01;
  assign sel_971472 = array_index_971203 == array_index_948889 ? add_971471 : sel_971468;
  assign add_971475 = sel_971472 + 8'h01;
  assign sel_971476 = array_index_971203 == array_index_948895 ? add_971475 : sel_971472;
  assign add_971479 = sel_971476 + 8'h01;
  assign sel_971480 = array_index_971203 == array_index_948901 ? add_971479 : sel_971476;
  assign add_971483 = sel_971480 + 8'h01;
  assign sel_971484 = array_index_971203 == array_index_948907 ? add_971483 : sel_971480;
  assign add_971487 = sel_971484 + 8'h01;
  assign sel_971488 = array_index_971203 == array_index_948913 ? add_971487 : sel_971484;
  assign add_971491 = sel_971488 + 8'h01;
  assign sel_971492 = array_index_971203 == array_index_948919 ? add_971491 : sel_971488;
  assign add_971495 = sel_971492 + 8'h01;
  assign sel_971496 = array_index_971203 == array_index_948925 ? add_971495 : sel_971492;
  assign add_971499 = sel_971496 + 8'h01;
  assign sel_971500 = array_index_971203 == array_index_948931 ? add_971499 : sel_971496;
  assign add_971503 = sel_971500 + 8'h01;
  assign sel_971504 = array_index_971203 == array_index_948937 ? add_971503 : sel_971500;
  assign add_971507 = sel_971504 + 8'h01;
  assign sel_971508 = array_index_971203 == array_index_948943 ? add_971507 : sel_971504;
  assign add_971511 = sel_971508 + 8'h01;
  assign sel_971512 = array_index_971203 == array_index_948949 ? add_971511 : sel_971508;
  assign add_971515 = sel_971512 + 8'h01;
  assign sel_971516 = array_index_971203 == array_index_948955 ? add_971515 : sel_971512;
  assign add_971519 = sel_971516 + 8'h01;
  assign sel_971520 = array_index_971203 == array_index_948961 ? add_971519 : sel_971516;
  assign add_971523 = sel_971520 + 8'h01;
  assign sel_971524 = array_index_971203 == array_index_948967 ? add_971523 : sel_971520;
  assign add_971527 = sel_971524 + 8'h01;
  assign sel_971528 = array_index_971203 == array_index_948973 ? add_971527 : sel_971524;
  assign add_971531 = sel_971528 + 8'h01;
  assign sel_971532 = array_index_971203 == array_index_948979 ? add_971531 : sel_971528;
  assign add_971535 = sel_971532 + 8'h01;
  assign sel_971536 = array_index_971203 == array_index_948985 ? add_971535 : sel_971532;
  assign add_971539 = sel_971536 + 8'h01;
  assign sel_971540 = array_index_971203 == array_index_948991 ? add_971539 : sel_971536;
  assign add_971543 = sel_971540 + 8'h01;
  assign sel_971544 = array_index_971203 == array_index_948997 ? add_971543 : sel_971540;
  assign add_971547 = sel_971544 + 8'h01;
  assign sel_971548 = array_index_971203 == array_index_949003 ? add_971547 : sel_971544;
  assign add_971551 = sel_971548 + 8'h01;
  assign sel_971552 = array_index_971203 == array_index_949009 ? add_971551 : sel_971548;
  assign add_971555 = sel_971552 + 8'h01;
  assign sel_971556 = array_index_971203 == array_index_949015 ? add_971555 : sel_971552;
  assign add_971559 = sel_971556 + 8'h01;
  assign sel_971560 = array_index_971203 == array_index_949021 ? add_971559 : sel_971556;
  assign add_971563 = sel_971560 + 8'h01;
  assign sel_971564 = array_index_971203 == array_index_949027 ? add_971563 : sel_971560;
  assign add_971567 = sel_971564 + 8'h01;
  assign sel_971568 = array_index_971203 == array_index_949033 ? add_971567 : sel_971564;
  assign add_971571 = sel_971568 + 8'h01;
  assign sel_971572 = array_index_971203 == array_index_949039 ? add_971571 : sel_971568;
  assign add_971575 = sel_971572 + 8'h01;
  assign sel_971576 = array_index_971203 == array_index_949045 ? add_971575 : sel_971572;
  assign add_971579 = sel_971576 + 8'h01;
  assign sel_971580 = array_index_971203 == array_index_949051 ? add_971579 : sel_971576;
  assign add_971583 = sel_971580 + 8'h01;
  assign sel_971584 = array_index_971203 == array_index_949057 ? add_971583 : sel_971580;
  assign add_971587 = sel_971584 + 8'h01;
  assign sel_971588 = array_index_971203 == array_index_949063 ? add_971587 : sel_971584;
  assign add_971591 = sel_971588 + 8'h01;
  assign sel_971592 = array_index_971203 == array_index_949069 ? add_971591 : sel_971588;
  assign add_971595 = sel_971592 + 8'h01;
  assign sel_971596 = array_index_971203 == array_index_949075 ? add_971595 : sel_971592;
  assign add_971599 = sel_971596 + 8'h01;
  assign sel_971600 = array_index_971203 == array_index_949081 ? add_971599 : sel_971596;
  assign add_971604 = sel_971600 + 8'h01;
  assign array_index_971605 = set1_unflattened[7'h39];
  assign sel_971606 = array_index_971203 == array_index_949087 ? add_971604 : sel_971600;
  assign add_971609 = sel_971606 + 8'h01;
  assign sel_971610 = array_index_971605 == array_index_948483 ? add_971609 : sel_971606;
  assign add_971613 = sel_971610 + 8'h01;
  assign sel_971614 = array_index_971605 == array_index_948487 ? add_971613 : sel_971610;
  assign add_971617 = sel_971614 + 8'h01;
  assign sel_971618 = array_index_971605 == array_index_948495 ? add_971617 : sel_971614;
  assign add_971621 = sel_971618 + 8'h01;
  assign sel_971622 = array_index_971605 == array_index_948503 ? add_971621 : sel_971618;
  assign add_971625 = sel_971622 + 8'h01;
  assign sel_971626 = array_index_971605 == array_index_948511 ? add_971625 : sel_971622;
  assign add_971629 = sel_971626 + 8'h01;
  assign sel_971630 = array_index_971605 == array_index_948519 ? add_971629 : sel_971626;
  assign add_971633 = sel_971630 + 8'h01;
  assign sel_971634 = array_index_971605 == array_index_948527 ? add_971633 : sel_971630;
  assign add_971637 = sel_971634 + 8'h01;
  assign sel_971638 = array_index_971605 == array_index_948535 ? add_971637 : sel_971634;
  assign add_971641 = sel_971638 + 8'h01;
  assign sel_971642 = array_index_971605 == array_index_948541 ? add_971641 : sel_971638;
  assign add_971645 = sel_971642 + 8'h01;
  assign sel_971646 = array_index_971605 == array_index_948547 ? add_971645 : sel_971642;
  assign add_971649 = sel_971646 + 8'h01;
  assign sel_971650 = array_index_971605 == array_index_948553 ? add_971649 : sel_971646;
  assign add_971653 = sel_971650 + 8'h01;
  assign sel_971654 = array_index_971605 == array_index_948559 ? add_971653 : sel_971650;
  assign add_971657 = sel_971654 + 8'h01;
  assign sel_971658 = array_index_971605 == array_index_948565 ? add_971657 : sel_971654;
  assign add_971661 = sel_971658 + 8'h01;
  assign sel_971662 = array_index_971605 == array_index_948571 ? add_971661 : sel_971658;
  assign add_971665 = sel_971662 + 8'h01;
  assign sel_971666 = array_index_971605 == array_index_948577 ? add_971665 : sel_971662;
  assign add_971669 = sel_971666 + 8'h01;
  assign sel_971670 = array_index_971605 == array_index_948583 ? add_971669 : sel_971666;
  assign add_971673 = sel_971670 + 8'h01;
  assign sel_971674 = array_index_971605 == array_index_948589 ? add_971673 : sel_971670;
  assign add_971677 = sel_971674 + 8'h01;
  assign sel_971678 = array_index_971605 == array_index_948595 ? add_971677 : sel_971674;
  assign add_971681 = sel_971678 + 8'h01;
  assign sel_971682 = array_index_971605 == array_index_948601 ? add_971681 : sel_971678;
  assign add_971685 = sel_971682 + 8'h01;
  assign sel_971686 = array_index_971605 == array_index_948607 ? add_971685 : sel_971682;
  assign add_971689 = sel_971686 + 8'h01;
  assign sel_971690 = array_index_971605 == array_index_948613 ? add_971689 : sel_971686;
  assign add_971693 = sel_971690 + 8'h01;
  assign sel_971694 = array_index_971605 == array_index_948619 ? add_971693 : sel_971690;
  assign add_971697 = sel_971694 + 8'h01;
  assign sel_971698 = array_index_971605 == array_index_948625 ? add_971697 : sel_971694;
  assign add_971701 = sel_971698 + 8'h01;
  assign sel_971702 = array_index_971605 == array_index_948631 ? add_971701 : sel_971698;
  assign add_971705 = sel_971702 + 8'h01;
  assign sel_971706 = array_index_971605 == array_index_948637 ? add_971705 : sel_971702;
  assign add_971709 = sel_971706 + 8'h01;
  assign sel_971710 = array_index_971605 == array_index_948643 ? add_971709 : sel_971706;
  assign add_971713 = sel_971710 + 8'h01;
  assign sel_971714 = array_index_971605 == array_index_948649 ? add_971713 : sel_971710;
  assign add_971717 = sel_971714 + 8'h01;
  assign sel_971718 = array_index_971605 == array_index_948655 ? add_971717 : sel_971714;
  assign add_971721 = sel_971718 + 8'h01;
  assign sel_971722 = array_index_971605 == array_index_948661 ? add_971721 : sel_971718;
  assign add_971725 = sel_971722 + 8'h01;
  assign sel_971726 = array_index_971605 == array_index_948667 ? add_971725 : sel_971722;
  assign add_971729 = sel_971726 + 8'h01;
  assign sel_971730 = array_index_971605 == array_index_948673 ? add_971729 : sel_971726;
  assign add_971733 = sel_971730 + 8'h01;
  assign sel_971734 = array_index_971605 == array_index_948679 ? add_971733 : sel_971730;
  assign add_971737 = sel_971734 + 8'h01;
  assign sel_971738 = array_index_971605 == array_index_948685 ? add_971737 : sel_971734;
  assign add_971741 = sel_971738 + 8'h01;
  assign sel_971742 = array_index_971605 == array_index_948691 ? add_971741 : sel_971738;
  assign add_971745 = sel_971742 + 8'h01;
  assign sel_971746 = array_index_971605 == array_index_948697 ? add_971745 : sel_971742;
  assign add_971749 = sel_971746 + 8'h01;
  assign sel_971750 = array_index_971605 == array_index_948703 ? add_971749 : sel_971746;
  assign add_971753 = sel_971750 + 8'h01;
  assign sel_971754 = array_index_971605 == array_index_948709 ? add_971753 : sel_971750;
  assign add_971757 = sel_971754 + 8'h01;
  assign sel_971758 = array_index_971605 == array_index_948715 ? add_971757 : sel_971754;
  assign add_971761 = sel_971758 + 8'h01;
  assign sel_971762 = array_index_971605 == array_index_948721 ? add_971761 : sel_971758;
  assign add_971765 = sel_971762 + 8'h01;
  assign sel_971766 = array_index_971605 == array_index_948727 ? add_971765 : sel_971762;
  assign add_971769 = sel_971766 + 8'h01;
  assign sel_971770 = array_index_971605 == array_index_948733 ? add_971769 : sel_971766;
  assign add_971773 = sel_971770 + 8'h01;
  assign sel_971774 = array_index_971605 == array_index_948739 ? add_971773 : sel_971770;
  assign add_971777 = sel_971774 + 8'h01;
  assign sel_971778 = array_index_971605 == array_index_948745 ? add_971777 : sel_971774;
  assign add_971781 = sel_971778 + 8'h01;
  assign sel_971782 = array_index_971605 == array_index_948751 ? add_971781 : sel_971778;
  assign add_971785 = sel_971782 + 8'h01;
  assign sel_971786 = array_index_971605 == array_index_948757 ? add_971785 : sel_971782;
  assign add_971789 = sel_971786 + 8'h01;
  assign sel_971790 = array_index_971605 == array_index_948763 ? add_971789 : sel_971786;
  assign add_971793 = sel_971790 + 8'h01;
  assign sel_971794 = array_index_971605 == array_index_948769 ? add_971793 : sel_971790;
  assign add_971797 = sel_971794 + 8'h01;
  assign sel_971798 = array_index_971605 == array_index_948775 ? add_971797 : sel_971794;
  assign add_971801 = sel_971798 + 8'h01;
  assign sel_971802 = array_index_971605 == array_index_948781 ? add_971801 : sel_971798;
  assign add_971805 = sel_971802 + 8'h01;
  assign sel_971806 = array_index_971605 == array_index_948787 ? add_971805 : sel_971802;
  assign add_971809 = sel_971806 + 8'h01;
  assign sel_971810 = array_index_971605 == array_index_948793 ? add_971809 : sel_971806;
  assign add_971813 = sel_971810 + 8'h01;
  assign sel_971814 = array_index_971605 == array_index_948799 ? add_971813 : sel_971810;
  assign add_971817 = sel_971814 + 8'h01;
  assign sel_971818 = array_index_971605 == array_index_948805 ? add_971817 : sel_971814;
  assign add_971821 = sel_971818 + 8'h01;
  assign sel_971822 = array_index_971605 == array_index_948811 ? add_971821 : sel_971818;
  assign add_971825 = sel_971822 + 8'h01;
  assign sel_971826 = array_index_971605 == array_index_948817 ? add_971825 : sel_971822;
  assign add_971829 = sel_971826 + 8'h01;
  assign sel_971830 = array_index_971605 == array_index_948823 ? add_971829 : sel_971826;
  assign add_971833 = sel_971830 + 8'h01;
  assign sel_971834 = array_index_971605 == array_index_948829 ? add_971833 : sel_971830;
  assign add_971837 = sel_971834 + 8'h01;
  assign sel_971838 = array_index_971605 == array_index_948835 ? add_971837 : sel_971834;
  assign add_971841 = sel_971838 + 8'h01;
  assign sel_971842 = array_index_971605 == array_index_948841 ? add_971841 : sel_971838;
  assign add_971845 = sel_971842 + 8'h01;
  assign sel_971846 = array_index_971605 == array_index_948847 ? add_971845 : sel_971842;
  assign add_971849 = sel_971846 + 8'h01;
  assign sel_971850 = array_index_971605 == array_index_948853 ? add_971849 : sel_971846;
  assign add_971853 = sel_971850 + 8'h01;
  assign sel_971854 = array_index_971605 == array_index_948859 ? add_971853 : sel_971850;
  assign add_971857 = sel_971854 + 8'h01;
  assign sel_971858 = array_index_971605 == array_index_948865 ? add_971857 : sel_971854;
  assign add_971861 = sel_971858 + 8'h01;
  assign sel_971862 = array_index_971605 == array_index_948871 ? add_971861 : sel_971858;
  assign add_971865 = sel_971862 + 8'h01;
  assign sel_971866 = array_index_971605 == array_index_948877 ? add_971865 : sel_971862;
  assign add_971869 = sel_971866 + 8'h01;
  assign sel_971870 = array_index_971605 == array_index_948883 ? add_971869 : sel_971866;
  assign add_971873 = sel_971870 + 8'h01;
  assign sel_971874 = array_index_971605 == array_index_948889 ? add_971873 : sel_971870;
  assign add_971877 = sel_971874 + 8'h01;
  assign sel_971878 = array_index_971605 == array_index_948895 ? add_971877 : sel_971874;
  assign add_971881 = sel_971878 + 8'h01;
  assign sel_971882 = array_index_971605 == array_index_948901 ? add_971881 : sel_971878;
  assign add_971885 = sel_971882 + 8'h01;
  assign sel_971886 = array_index_971605 == array_index_948907 ? add_971885 : sel_971882;
  assign add_971889 = sel_971886 + 8'h01;
  assign sel_971890 = array_index_971605 == array_index_948913 ? add_971889 : sel_971886;
  assign add_971893 = sel_971890 + 8'h01;
  assign sel_971894 = array_index_971605 == array_index_948919 ? add_971893 : sel_971890;
  assign add_971897 = sel_971894 + 8'h01;
  assign sel_971898 = array_index_971605 == array_index_948925 ? add_971897 : sel_971894;
  assign add_971901 = sel_971898 + 8'h01;
  assign sel_971902 = array_index_971605 == array_index_948931 ? add_971901 : sel_971898;
  assign add_971905 = sel_971902 + 8'h01;
  assign sel_971906 = array_index_971605 == array_index_948937 ? add_971905 : sel_971902;
  assign add_971909 = sel_971906 + 8'h01;
  assign sel_971910 = array_index_971605 == array_index_948943 ? add_971909 : sel_971906;
  assign add_971913 = sel_971910 + 8'h01;
  assign sel_971914 = array_index_971605 == array_index_948949 ? add_971913 : sel_971910;
  assign add_971917 = sel_971914 + 8'h01;
  assign sel_971918 = array_index_971605 == array_index_948955 ? add_971917 : sel_971914;
  assign add_971921 = sel_971918 + 8'h01;
  assign sel_971922 = array_index_971605 == array_index_948961 ? add_971921 : sel_971918;
  assign add_971925 = sel_971922 + 8'h01;
  assign sel_971926 = array_index_971605 == array_index_948967 ? add_971925 : sel_971922;
  assign add_971929 = sel_971926 + 8'h01;
  assign sel_971930 = array_index_971605 == array_index_948973 ? add_971929 : sel_971926;
  assign add_971933 = sel_971930 + 8'h01;
  assign sel_971934 = array_index_971605 == array_index_948979 ? add_971933 : sel_971930;
  assign add_971937 = sel_971934 + 8'h01;
  assign sel_971938 = array_index_971605 == array_index_948985 ? add_971937 : sel_971934;
  assign add_971941 = sel_971938 + 8'h01;
  assign sel_971942 = array_index_971605 == array_index_948991 ? add_971941 : sel_971938;
  assign add_971945 = sel_971942 + 8'h01;
  assign sel_971946 = array_index_971605 == array_index_948997 ? add_971945 : sel_971942;
  assign add_971949 = sel_971946 + 8'h01;
  assign sel_971950 = array_index_971605 == array_index_949003 ? add_971949 : sel_971946;
  assign add_971953 = sel_971950 + 8'h01;
  assign sel_971954 = array_index_971605 == array_index_949009 ? add_971953 : sel_971950;
  assign add_971957 = sel_971954 + 8'h01;
  assign sel_971958 = array_index_971605 == array_index_949015 ? add_971957 : sel_971954;
  assign add_971961 = sel_971958 + 8'h01;
  assign sel_971962 = array_index_971605 == array_index_949021 ? add_971961 : sel_971958;
  assign add_971965 = sel_971962 + 8'h01;
  assign sel_971966 = array_index_971605 == array_index_949027 ? add_971965 : sel_971962;
  assign add_971969 = sel_971966 + 8'h01;
  assign sel_971970 = array_index_971605 == array_index_949033 ? add_971969 : sel_971966;
  assign add_971973 = sel_971970 + 8'h01;
  assign sel_971974 = array_index_971605 == array_index_949039 ? add_971973 : sel_971970;
  assign add_971977 = sel_971974 + 8'h01;
  assign sel_971978 = array_index_971605 == array_index_949045 ? add_971977 : sel_971974;
  assign add_971981 = sel_971978 + 8'h01;
  assign sel_971982 = array_index_971605 == array_index_949051 ? add_971981 : sel_971978;
  assign add_971985 = sel_971982 + 8'h01;
  assign sel_971986 = array_index_971605 == array_index_949057 ? add_971985 : sel_971982;
  assign add_971989 = sel_971986 + 8'h01;
  assign sel_971990 = array_index_971605 == array_index_949063 ? add_971989 : sel_971986;
  assign add_971993 = sel_971990 + 8'h01;
  assign sel_971994 = array_index_971605 == array_index_949069 ? add_971993 : sel_971990;
  assign add_971997 = sel_971994 + 8'h01;
  assign sel_971998 = array_index_971605 == array_index_949075 ? add_971997 : sel_971994;
  assign add_972001 = sel_971998 + 8'h01;
  assign sel_972002 = array_index_971605 == array_index_949081 ? add_972001 : sel_971998;
  assign add_972006 = sel_972002 + 8'h01;
  assign array_index_972007 = set1_unflattened[7'h3a];
  assign sel_972008 = array_index_971605 == array_index_949087 ? add_972006 : sel_972002;
  assign add_972011 = sel_972008 + 8'h01;
  assign sel_972012 = array_index_972007 == array_index_948483 ? add_972011 : sel_972008;
  assign add_972015 = sel_972012 + 8'h01;
  assign sel_972016 = array_index_972007 == array_index_948487 ? add_972015 : sel_972012;
  assign add_972019 = sel_972016 + 8'h01;
  assign sel_972020 = array_index_972007 == array_index_948495 ? add_972019 : sel_972016;
  assign add_972023 = sel_972020 + 8'h01;
  assign sel_972024 = array_index_972007 == array_index_948503 ? add_972023 : sel_972020;
  assign add_972027 = sel_972024 + 8'h01;
  assign sel_972028 = array_index_972007 == array_index_948511 ? add_972027 : sel_972024;
  assign add_972031 = sel_972028 + 8'h01;
  assign sel_972032 = array_index_972007 == array_index_948519 ? add_972031 : sel_972028;
  assign add_972035 = sel_972032 + 8'h01;
  assign sel_972036 = array_index_972007 == array_index_948527 ? add_972035 : sel_972032;
  assign add_972039 = sel_972036 + 8'h01;
  assign sel_972040 = array_index_972007 == array_index_948535 ? add_972039 : sel_972036;
  assign add_972043 = sel_972040 + 8'h01;
  assign sel_972044 = array_index_972007 == array_index_948541 ? add_972043 : sel_972040;
  assign add_972047 = sel_972044 + 8'h01;
  assign sel_972048 = array_index_972007 == array_index_948547 ? add_972047 : sel_972044;
  assign add_972051 = sel_972048 + 8'h01;
  assign sel_972052 = array_index_972007 == array_index_948553 ? add_972051 : sel_972048;
  assign add_972055 = sel_972052 + 8'h01;
  assign sel_972056 = array_index_972007 == array_index_948559 ? add_972055 : sel_972052;
  assign add_972059 = sel_972056 + 8'h01;
  assign sel_972060 = array_index_972007 == array_index_948565 ? add_972059 : sel_972056;
  assign add_972063 = sel_972060 + 8'h01;
  assign sel_972064 = array_index_972007 == array_index_948571 ? add_972063 : sel_972060;
  assign add_972067 = sel_972064 + 8'h01;
  assign sel_972068 = array_index_972007 == array_index_948577 ? add_972067 : sel_972064;
  assign add_972071 = sel_972068 + 8'h01;
  assign sel_972072 = array_index_972007 == array_index_948583 ? add_972071 : sel_972068;
  assign add_972075 = sel_972072 + 8'h01;
  assign sel_972076 = array_index_972007 == array_index_948589 ? add_972075 : sel_972072;
  assign add_972079 = sel_972076 + 8'h01;
  assign sel_972080 = array_index_972007 == array_index_948595 ? add_972079 : sel_972076;
  assign add_972083 = sel_972080 + 8'h01;
  assign sel_972084 = array_index_972007 == array_index_948601 ? add_972083 : sel_972080;
  assign add_972087 = sel_972084 + 8'h01;
  assign sel_972088 = array_index_972007 == array_index_948607 ? add_972087 : sel_972084;
  assign add_972091 = sel_972088 + 8'h01;
  assign sel_972092 = array_index_972007 == array_index_948613 ? add_972091 : sel_972088;
  assign add_972095 = sel_972092 + 8'h01;
  assign sel_972096 = array_index_972007 == array_index_948619 ? add_972095 : sel_972092;
  assign add_972099 = sel_972096 + 8'h01;
  assign sel_972100 = array_index_972007 == array_index_948625 ? add_972099 : sel_972096;
  assign add_972103 = sel_972100 + 8'h01;
  assign sel_972104 = array_index_972007 == array_index_948631 ? add_972103 : sel_972100;
  assign add_972107 = sel_972104 + 8'h01;
  assign sel_972108 = array_index_972007 == array_index_948637 ? add_972107 : sel_972104;
  assign add_972111 = sel_972108 + 8'h01;
  assign sel_972112 = array_index_972007 == array_index_948643 ? add_972111 : sel_972108;
  assign add_972115 = sel_972112 + 8'h01;
  assign sel_972116 = array_index_972007 == array_index_948649 ? add_972115 : sel_972112;
  assign add_972119 = sel_972116 + 8'h01;
  assign sel_972120 = array_index_972007 == array_index_948655 ? add_972119 : sel_972116;
  assign add_972123 = sel_972120 + 8'h01;
  assign sel_972124 = array_index_972007 == array_index_948661 ? add_972123 : sel_972120;
  assign add_972127 = sel_972124 + 8'h01;
  assign sel_972128 = array_index_972007 == array_index_948667 ? add_972127 : sel_972124;
  assign add_972131 = sel_972128 + 8'h01;
  assign sel_972132 = array_index_972007 == array_index_948673 ? add_972131 : sel_972128;
  assign add_972135 = sel_972132 + 8'h01;
  assign sel_972136 = array_index_972007 == array_index_948679 ? add_972135 : sel_972132;
  assign add_972139 = sel_972136 + 8'h01;
  assign sel_972140 = array_index_972007 == array_index_948685 ? add_972139 : sel_972136;
  assign add_972143 = sel_972140 + 8'h01;
  assign sel_972144 = array_index_972007 == array_index_948691 ? add_972143 : sel_972140;
  assign add_972147 = sel_972144 + 8'h01;
  assign sel_972148 = array_index_972007 == array_index_948697 ? add_972147 : sel_972144;
  assign add_972151 = sel_972148 + 8'h01;
  assign sel_972152 = array_index_972007 == array_index_948703 ? add_972151 : sel_972148;
  assign add_972155 = sel_972152 + 8'h01;
  assign sel_972156 = array_index_972007 == array_index_948709 ? add_972155 : sel_972152;
  assign add_972159 = sel_972156 + 8'h01;
  assign sel_972160 = array_index_972007 == array_index_948715 ? add_972159 : sel_972156;
  assign add_972163 = sel_972160 + 8'h01;
  assign sel_972164 = array_index_972007 == array_index_948721 ? add_972163 : sel_972160;
  assign add_972167 = sel_972164 + 8'h01;
  assign sel_972168 = array_index_972007 == array_index_948727 ? add_972167 : sel_972164;
  assign add_972171 = sel_972168 + 8'h01;
  assign sel_972172 = array_index_972007 == array_index_948733 ? add_972171 : sel_972168;
  assign add_972175 = sel_972172 + 8'h01;
  assign sel_972176 = array_index_972007 == array_index_948739 ? add_972175 : sel_972172;
  assign add_972179 = sel_972176 + 8'h01;
  assign sel_972180 = array_index_972007 == array_index_948745 ? add_972179 : sel_972176;
  assign add_972183 = sel_972180 + 8'h01;
  assign sel_972184 = array_index_972007 == array_index_948751 ? add_972183 : sel_972180;
  assign add_972187 = sel_972184 + 8'h01;
  assign sel_972188 = array_index_972007 == array_index_948757 ? add_972187 : sel_972184;
  assign add_972191 = sel_972188 + 8'h01;
  assign sel_972192 = array_index_972007 == array_index_948763 ? add_972191 : sel_972188;
  assign add_972195 = sel_972192 + 8'h01;
  assign sel_972196 = array_index_972007 == array_index_948769 ? add_972195 : sel_972192;
  assign add_972199 = sel_972196 + 8'h01;
  assign sel_972200 = array_index_972007 == array_index_948775 ? add_972199 : sel_972196;
  assign add_972203 = sel_972200 + 8'h01;
  assign sel_972204 = array_index_972007 == array_index_948781 ? add_972203 : sel_972200;
  assign add_972207 = sel_972204 + 8'h01;
  assign sel_972208 = array_index_972007 == array_index_948787 ? add_972207 : sel_972204;
  assign add_972211 = sel_972208 + 8'h01;
  assign sel_972212 = array_index_972007 == array_index_948793 ? add_972211 : sel_972208;
  assign add_972215 = sel_972212 + 8'h01;
  assign sel_972216 = array_index_972007 == array_index_948799 ? add_972215 : sel_972212;
  assign add_972219 = sel_972216 + 8'h01;
  assign sel_972220 = array_index_972007 == array_index_948805 ? add_972219 : sel_972216;
  assign add_972223 = sel_972220 + 8'h01;
  assign sel_972224 = array_index_972007 == array_index_948811 ? add_972223 : sel_972220;
  assign add_972227 = sel_972224 + 8'h01;
  assign sel_972228 = array_index_972007 == array_index_948817 ? add_972227 : sel_972224;
  assign add_972231 = sel_972228 + 8'h01;
  assign sel_972232 = array_index_972007 == array_index_948823 ? add_972231 : sel_972228;
  assign add_972235 = sel_972232 + 8'h01;
  assign sel_972236 = array_index_972007 == array_index_948829 ? add_972235 : sel_972232;
  assign add_972239 = sel_972236 + 8'h01;
  assign sel_972240 = array_index_972007 == array_index_948835 ? add_972239 : sel_972236;
  assign add_972243 = sel_972240 + 8'h01;
  assign sel_972244 = array_index_972007 == array_index_948841 ? add_972243 : sel_972240;
  assign add_972247 = sel_972244 + 8'h01;
  assign sel_972248 = array_index_972007 == array_index_948847 ? add_972247 : sel_972244;
  assign add_972251 = sel_972248 + 8'h01;
  assign sel_972252 = array_index_972007 == array_index_948853 ? add_972251 : sel_972248;
  assign add_972255 = sel_972252 + 8'h01;
  assign sel_972256 = array_index_972007 == array_index_948859 ? add_972255 : sel_972252;
  assign add_972259 = sel_972256 + 8'h01;
  assign sel_972260 = array_index_972007 == array_index_948865 ? add_972259 : sel_972256;
  assign add_972263 = sel_972260 + 8'h01;
  assign sel_972264 = array_index_972007 == array_index_948871 ? add_972263 : sel_972260;
  assign add_972267 = sel_972264 + 8'h01;
  assign sel_972268 = array_index_972007 == array_index_948877 ? add_972267 : sel_972264;
  assign add_972271 = sel_972268 + 8'h01;
  assign sel_972272 = array_index_972007 == array_index_948883 ? add_972271 : sel_972268;
  assign add_972275 = sel_972272 + 8'h01;
  assign sel_972276 = array_index_972007 == array_index_948889 ? add_972275 : sel_972272;
  assign add_972279 = sel_972276 + 8'h01;
  assign sel_972280 = array_index_972007 == array_index_948895 ? add_972279 : sel_972276;
  assign add_972283 = sel_972280 + 8'h01;
  assign sel_972284 = array_index_972007 == array_index_948901 ? add_972283 : sel_972280;
  assign add_972287 = sel_972284 + 8'h01;
  assign sel_972288 = array_index_972007 == array_index_948907 ? add_972287 : sel_972284;
  assign add_972291 = sel_972288 + 8'h01;
  assign sel_972292 = array_index_972007 == array_index_948913 ? add_972291 : sel_972288;
  assign add_972295 = sel_972292 + 8'h01;
  assign sel_972296 = array_index_972007 == array_index_948919 ? add_972295 : sel_972292;
  assign add_972299 = sel_972296 + 8'h01;
  assign sel_972300 = array_index_972007 == array_index_948925 ? add_972299 : sel_972296;
  assign add_972303 = sel_972300 + 8'h01;
  assign sel_972304 = array_index_972007 == array_index_948931 ? add_972303 : sel_972300;
  assign add_972307 = sel_972304 + 8'h01;
  assign sel_972308 = array_index_972007 == array_index_948937 ? add_972307 : sel_972304;
  assign add_972311 = sel_972308 + 8'h01;
  assign sel_972312 = array_index_972007 == array_index_948943 ? add_972311 : sel_972308;
  assign add_972315 = sel_972312 + 8'h01;
  assign sel_972316 = array_index_972007 == array_index_948949 ? add_972315 : sel_972312;
  assign add_972319 = sel_972316 + 8'h01;
  assign sel_972320 = array_index_972007 == array_index_948955 ? add_972319 : sel_972316;
  assign add_972323 = sel_972320 + 8'h01;
  assign sel_972324 = array_index_972007 == array_index_948961 ? add_972323 : sel_972320;
  assign add_972327 = sel_972324 + 8'h01;
  assign sel_972328 = array_index_972007 == array_index_948967 ? add_972327 : sel_972324;
  assign add_972331 = sel_972328 + 8'h01;
  assign sel_972332 = array_index_972007 == array_index_948973 ? add_972331 : sel_972328;
  assign add_972335 = sel_972332 + 8'h01;
  assign sel_972336 = array_index_972007 == array_index_948979 ? add_972335 : sel_972332;
  assign add_972339 = sel_972336 + 8'h01;
  assign sel_972340 = array_index_972007 == array_index_948985 ? add_972339 : sel_972336;
  assign add_972343 = sel_972340 + 8'h01;
  assign sel_972344 = array_index_972007 == array_index_948991 ? add_972343 : sel_972340;
  assign add_972347 = sel_972344 + 8'h01;
  assign sel_972348 = array_index_972007 == array_index_948997 ? add_972347 : sel_972344;
  assign add_972351 = sel_972348 + 8'h01;
  assign sel_972352 = array_index_972007 == array_index_949003 ? add_972351 : sel_972348;
  assign add_972355 = sel_972352 + 8'h01;
  assign sel_972356 = array_index_972007 == array_index_949009 ? add_972355 : sel_972352;
  assign add_972359 = sel_972356 + 8'h01;
  assign sel_972360 = array_index_972007 == array_index_949015 ? add_972359 : sel_972356;
  assign add_972363 = sel_972360 + 8'h01;
  assign sel_972364 = array_index_972007 == array_index_949021 ? add_972363 : sel_972360;
  assign add_972367 = sel_972364 + 8'h01;
  assign sel_972368 = array_index_972007 == array_index_949027 ? add_972367 : sel_972364;
  assign add_972371 = sel_972368 + 8'h01;
  assign sel_972372 = array_index_972007 == array_index_949033 ? add_972371 : sel_972368;
  assign add_972375 = sel_972372 + 8'h01;
  assign sel_972376 = array_index_972007 == array_index_949039 ? add_972375 : sel_972372;
  assign add_972379 = sel_972376 + 8'h01;
  assign sel_972380 = array_index_972007 == array_index_949045 ? add_972379 : sel_972376;
  assign add_972383 = sel_972380 + 8'h01;
  assign sel_972384 = array_index_972007 == array_index_949051 ? add_972383 : sel_972380;
  assign add_972387 = sel_972384 + 8'h01;
  assign sel_972388 = array_index_972007 == array_index_949057 ? add_972387 : sel_972384;
  assign add_972391 = sel_972388 + 8'h01;
  assign sel_972392 = array_index_972007 == array_index_949063 ? add_972391 : sel_972388;
  assign add_972395 = sel_972392 + 8'h01;
  assign sel_972396 = array_index_972007 == array_index_949069 ? add_972395 : sel_972392;
  assign add_972399 = sel_972396 + 8'h01;
  assign sel_972400 = array_index_972007 == array_index_949075 ? add_972399 : sel_972396;
  assign add_972403 = sel_972400 + 8'h01;
  assign sel_972404 = array_index_972007 == array_index_949081 ? add_972403 : sel_972400;
  assign add_972408 = sel_972404 + 8'h01;
  assign array_index_972409 = set1_unflattened[7'h3b];
  assign sel_972410 = array_index_972007 == array_index_949087 ? add_972408 : sel_972404;
  assign add_972413 = sel_972410 + 8'h01;
  assign sel_972414 = array_index_972409 == array_index_948483 ? add_972413 : sel_972410;
  assign add_972417 = sel_972414 + 8'h01;
  assign sel_972418 = array_index_972409 == array_index_948487 ? add_972417 : sel_972414;
  assign add_972421 = sel_972418 + 8'h01;
  assign sel_972422 = array_index_972409 == array_index_948495 ? add_972421 : sel_972418;
  assign add_972425 = sel_972422 + 8'h01;
  assign sel_972426 = array_index_972409 == array_index_948503 ? add_972425 : sel_972422;
  assign add_972429 = sel_972426 + 8'h01;
  assign sel_972430 = array_index_972409 == array_index_948511 ? add_972429 : sel_972426;
  assign add_972433 = sel_972430 + 8'h01;
  assign sel_972434 = array_index_972409 == array_index_948519 ? add_972433 : sel_972430;
  assign add_972437 = sel_972434 + 8'h01;
  assign sel_972438 = array_index_972409 == array_index_948527 ? add_972437 : sel_972434;
  assign add_972441 = sel_972438 + 8'h01;
  assign sel_972442 = array_index_972409 == array_index_948535 ? add_972441 : sel_972438;
  assign add_972445 = sel_972442 + 8'h01;
  assign sel_972446 = array_index_972409 == array_index_948541 ? add_972445 : sel_972442;
  assign add_972449 = sel_972446 + 8'h01;
  assign sel_972450 = array_index_972409 == array_index_948547 ? add_972449 : sel_972446;
  assign add_972453 = sel_972450 + 8'h01;
  assign sel_972454 = array_index_972409 == array_index_948553 ? add_972453 : sel_972450;
  assign add_972457 = sel_972454 + 8'h01;
  assign sel_972458 = array_index_972409 == array_index_948559 ? add_972457 : sel_972454;
  assign add_972461 = sel_972458 + 8'h01;
  assign sel_972462 = array_index_972409 == array_index_948565 ? add_972461 : sel_972458;
  assign add_972465 = sel_972462 + 8'h01;
  assign sel_972466 = array_index_972409 == array_index_948571 ? add_972465 : sel_972462;
  assign add_972469 = sel_972466 + 8'h01;
  assign sel_972470 = array_index_972409 == array_index_948577 ? add_972469 : sel_972466;
  assign add_972473 = sel_972470 + 8'h01;
  assign sel_972474 = array_index_972409 == array_index_948583 ? add_972473 : sel_972470;
  assign add_972477 = sel_972474 + 8'h01;
  assign sel_972478 = array_index_972409 == array_index_948589 ? add_972477 : sel_972474;
  assign add_972481 = sel_972478 + 8'h01;
  assign sel_972482 = array_index_972409 == array_index_948595 ? add_972481 : sel_972478;
  assign add_972485 = sel_972482 + 8'h01;
  assign sel_972486 = array_index_972409 == array_index_948601 ? add_972485 : sel_972482;
  assign add_972489 = sel_972486 + 8'h01;
  assign sel_972490 = array_index_972409 == array_index_948607 ? add_972489 : sel_972486;
  assign add_972493 = sel_972490 + 8'h01;
  assign sel_972494 = array_index_972409 == array_index_948613 ? add_972493 : sel_972490;
  assign add_972497 = sel_972494 + 8'h01;
  assign sel_972498 = array_index_972409 == array_index_948619 ? add_972497 : sel_972494;
  assign add_972501 = sel_972498 + 8'h01;
  assign sel_972502 = array_index_972409 == array_index_948625 ? add_972501 : sel_972498;
  assign add_972505 = sel_972502 + 8'h01;
  assign sel_972506 = array_index_972409 == array_index_948631 ? add_972505 : sel_972502;
  assign add_972509 = sel_972506 + 8'h01;
  assign sel_972510 = array_index_972409 == array_index_948637 ? add_972509 : sel_972506;
  assign add_972513 = sel_972510 + 8'h01;
  assign sel_972514 = array_index_972409 == array_index_948643 ? add_972513 : sel_972510;
  assign add_972517 = sel_972514 + 8'h01;
  assign sel_972518 = array_index_972409 == array_index_948649 ? add_972517 : sel_972514;
  assign add_972521 = sel_972518 + 8'h01;
  assign sel_972522 = array_index_972409 == array_index_948655 ? add_972521 : sel_972518;
  assign add_972525 = sel_972522 + 8'h01;
  assign sel_972526 = array_index_972409 == array_index_948661 ? add_972525 : sel_972522;
  assign add_972529 = sel_972526 + 8'h01;
  assign sel_972530 = array_index_972409 == array_index_948667 ? add_972529 : sel_972526;
  assign add_972533 = sel_972530 + 8'h01;
  assign sel_972534 = array_index_972409 == array_index_948673 ? add_972533 : sel_972530;
  assign add_972537 = sel_972534 + 8'h01;
  assign sel_972538 = array_index_972409 == array_index_948679 ? add_972537 : sel_972534;
  assign add_972541 = sel_972538 + 8'h01;
  assign sel_972542 = array_index_972409 == array_index_948685 ? add_972541 : sel_972538;
  assign add_972545 = sel_972542 + 8'h01;
  assign sel_972546 = array_index_972409 == array_index_948691 ? add_972545 : sel_972542;
  assign add_972549 = sel_972546 + 8'h01;
  assign sel_972550 = array_index_972409 == array_index_948697 ? add_972549 : sel_972546;
  assign add_972553 = sel_972550 + 8'h01;
  assign sel_972554 = array_index_972409 == array_index_948703 ? add_972553 : sel_972550;
  assign add_972557 = sel_972554 + 8'h01;
  assign sel_972558 = array_index_972409 == array_index_948709 ? add_972557 : sel_972554;
  assign add_972561 = sel_972558 + 8'h01;
  assign sel_972562 = array_index_972409 == array_index_948715 ? add_972561 : sel_972558;
  assign add_972565 = sel_972562 + 8'h01;
  assign sel_972566 = array_index_972409 == array_index_948721 ? add_972565 : sel_972562;
  assign add_972569 = sel_972566 + 8'h01;
  assign sel_972570 = array_index_972409 == array_index_948727 ? add_972569 : sel_972566;
  assign add_972573 = sel_972570 + 8'h01;
  assign sel_972574 = array_index_972409 == array_index_948733 ? add_972573 : sel_972570;
  assign add_972577 = sel_972574 + 8'h01;
  assign sel_972578 = array_index_972409 == array_index_948739 ? add_972577 : sel_972574;
  assign add_972581 = sel_972578 + 8'h01;
  assign sel_972582 = array_index_972409 == array_index_948745 ? add_972581 : sel_972578;
  assign add_972585 = sel_972582 + 8'h01;
  assign sel_972586 = array_index_972409 == array_index_948751 ? add_972585 : sel_972582;
  assign add_972589 = sel_972586 + 8'h01;
  assign sel_972590 = array_index_972409 == array_index_948757 ? add_972589 : sel_972586;
  assign add_972593 = sel_972590 + 8'h01;
  assign sel_972594 = array_index_972409 == array_index_948763 ? add_972593 : sel_972590;
  assign add_972597 = sel_972594 + 8'h01;
  assign sel_972598 = array_index_972409 == array_index_948769 ? add_972597 : sel_972594;
  assign add_972601 = sel_972598 + 8'h01;
  assign sel_972602 = array_index_972409 == array_index_948775 ? add_972601 : sel_972598;
  assign add_972605 = sel_972602 + 8'h01;
  assign sel_972606 = array_index_972409 == array_index_948781 ? add_972605 : sel_972602;
  assign add_972609 = sel_972606 + 8'h01;
  assign sel_972610 = array_index_972409 == array_index_948787 ? add_972609 : sel_972606;
  assign add_972613 = sel_972610 + 8'h01;
  assign sel_972614 = array_index_972409 == array_index_948793 ? add_972613 : sel_972610;
  assign add_972617 = sel_972614 + 8'h01;
  assign sel_972618 = array_index_972409 == array_index_948799 ? add_972617 : sel_972614;
  assign add_972621 = sel_972618 + 8'h01;
  assign sel_972622 = array_index_972409 == array_index_948805 ? add_972621 : sel_972618;
  assign add_972625 = sel_972622 + 8'h01;
  assign sel_972626 = array_index_972409 == array_index_948811 ? add_972625 : sel_972622;
  assign add_972629 = sel_972626 + 8'h01;
  assign sel_972630 = array_index_972409 == array_index_948817 ? add_972629 : sel_972626;
  assign add_972633 = sel_972630 + 8'h01;
  assign sel_972634 = array_index_972409 == array_index_948823 ? add_972633 : sel_972630;
  assign add_972637 = sel_972634 + 8'h01;
  assign sel_972638 = array_index_972409 == array_index_948829 ? add_972637 : sel_972634;
  assign add_972641 = sel_972638 + 8'h01;
  assign sel_972642 = array_index_972409 == array_index_948835 ? add_972641 : sel_972638;
  assign add_972645 = sel_972642 + 8'h01;
  assign sel_972646 = array_index_972409 == array_index_948841 ? add_972645 : sel_972642;
  assign add_972649 = sel_972646 + 8'h01;
  assign sel_972650 = array_index_972409 == array_index_948847 ? add_972649 : sel_972646;
  assign add_972653 = sel_972650 + 8'h01;
  assign sel_972654 = array_index_972409 == array_index_948853 ? add_972653 : sel_972650;
  assign add_972657 = sel_972654 + 8'h01;
  assign sel_972658 = array_index_972409 == array_index_948859 ? add_972657 : sel_972654;
  assign add_972661 = sel_972658 + 8'h01;
  assign sel_972662 = array_index_972409 == array_index_948865 ? add_972661 : sel_972658;
  assign add_972665 = sel_972662 + 8'h01;
  assign sel_972666 = array_index_972409 == array_index_948871 ? add_972665 : sel_972662;
  assign add_972669 = sel_972666 + 8'h01;
  assign sel_972670 = array_index_972409 == array_index_948877 ? add_972669 : sel_972666;
  assign add_972673 = sel_972670 + 8'h01;
  assign sel_972674 = array_index_972409 == array_index_948883 ? add_972673 : sel_972670;
  assign add_972677 = sel_972674 + 8'h01;
  assign sel_972678 = array_index_972409 == array_index_948889 ? add_972677 : sel_972674;
  assign add_972681 = sel_972678 + 8'h01;
  assign sel_972682 = array_index_972409 == array_index_948895 ? add_972681 : sel_972678;
  assign add_972685 = sel_972682 + 8'h01;
  assign sel_972686 = array_index_972409 == array_index_948901 ? add_972685 : sel_972682;
  assign add_972689 = sel_972686 + 8'h01;
  assign sel_972690 = array_index_972409 == array_index_948907 ? add_972689 : sel_972686;
  assign add_972693 = sel_972690 + 8'h01;
  assign sel_972694 = array_index_972409 == array_index_948913 ? add_972693 : sel_972690;
  assign add_972697 = sel_972694 + 8'h01;
  assign sel_972698 = array_index_972409 == array_index_948919 ? add_972697 : sel_972694;
  assign add_972701 = sel_972698 + 8'h01;
  assign sel_972702 = array_index_972409 == array_index_948925 ? add_972701 : sel_972698;
  assign add_972705 = sel_972702 + 8'h01;
  assign sel_972706 = array_index_972409 == array_index_948931 ? add_972705 : sel_972702;
  assign add_972709 = sel_972706 + 8'h01;
  assign sel_972710 = array_index_972409 == array_index_948937 ? add_972709 : sel_972706;
  assign add_972713 = sel_972710 + 8'h01;
  assign sel_972714 = array_index_972409 == array_index_948943 ? add_972713 : sel_972710;
  assign add_972717 = sel_972714 + 8'h01;
  assign sel_972718 = array_index_972409 == array_index_948949 ? add_972717 : sel_972714;
  assign add_972721 = sel_972718 + 8'h01;
  assign sel_972722 = array_index_972409 == array_index_948955 ? add_972721 : sel_972718;
  assign add_972725 = sel_972722 + 8'h01;
  assign sel_972726 = array_index_972409 == array_index_948961 ? add_972725 : sel_972722;
  assign add_972729 = sel_972726 + 8'h01;
  assign sel_972730 = array_index_972409 == array_index_948967 ? add_972729 : sel_972726;
  assign add_972733 = sel_972730 + 8'h01;
  assign sel_972734 = array_index_972409 == array_index_948973 ? add_972733 : sel_972730;
  assign add_972737 = sel_972734 + 8'h01;
  assign sel_972738 = array_index_972409 == array_index_948979 ? add_972737 : sel_972734;
  assign add_972741 = sel_972738 + 8'h01;
  assign sel_972742 = array_index_972409 == array_index_948985 ? add_972741 : sel_972738;
  assign add_972745 = sel_972742 + 8'h01;
  assign sel_972746 = array_index_972409 == array_index_948991 ? add_972745 : sel_972742;
  assign add_972749 = sel_972746 + 8'h01;
  assign sel_972750 = array_index_972409 == array_index_948997 ? add_972749 : sel_972746;
  assign add_972753 = sel_972750 + 8'h01;
  assign sel_972754 = array_index_972409 == array_index_949003 ? add_972753 : sel_972750;
  assign add_972757 = sel_972754 + 8'h01;
  assign sel_972758 = array_index_972409 == array_index_949009 ? add_972757 : sel_972754;
  assign add_972761 = sel_972758 + 8'h01;
  assign sel_972762 = array_index_972409 == array_index_949015 ? add_972761 : sel_972758;
  assign add_972765 = sel_972762 + 8'h01;
  assign sel_972766 = array_index_972409 == array_index_949021 ? add_972765 : sel_972762;
  assign add_972769 = sel_972766 + 8'h01;
  assign sel_972770 = array_index_972409 == array_index_949027 ? add_972769 : sel_972766;
  assign add_972773 = sel_972770 + 8'h01;
  assign sel_972774 = array_index_972409 == array_index_949033 ? add_972773 : sel_972770;
  assign add_972777 = sel_972774 + 8'h01;
  assign sel_972778 = array_index_972409 == array_index_949039 ? add_972777 : sel_972774;
  assign add_972781 = sel_972778 + 8'h01;
  assign sel_972782 = array_index_972409 == array_index_949045 ? add_972781 : sel_972778;
  assign add_972785 = sel_972782 + 8'h01;
  assign sel_972786 = array_index_972409 == array_index_949051 ? add_972785 : sel_972782;
  assign add_972789 = sel_972786 + 8'h01;
  assign sel_972790 = array_index_972409 == array_index_949057 ? add_972789 : sel_972786;
  assign add_972793 = sel_972790 + 8'h01;
  assign sel_972794 = array_index_972409 == array_index_949063 ? add_972793 : sel_972790;
  assign add_972797 = sel_972794 + 8'h01;
  assign sel_972798 = array_index_972409 == array_index_949069 ? add_972797 : sel_972794;
  assign add_972801 = sel_972798 + 8'h01;
  assign sel_972802 = array_index_972409 == array_index_949075 ? add_972801 : sel_972798;
  assign add_972805 = sel_972802 + 8'h01;
  assign sel_972806 = array_index_972409 == array_index_949081 ? add_972805 : sel_972802;
  assign add_972810 = sel_972806 + 8'h01;
  assign array_index_972811 = set1_unflattened[7'h3c];
  assign sel_972812 = array_index_972409 == array_index_949087 ? add_972810 : sel_972806;
  assign add_972815 = sel_972812 + 8'h01;
  assign sel_972816 = array_index_972811 == array_index_948483 ? add_972815 : sel_972812;
  assign add_972819 = sel_972816 + 8'h01;
  assign sel_972820 = array_index_972811 == array_index_948487 ? add_972819 : sel_972816;
  assign add_972823 = sel_972820 + 8'h01;
  assign sel_972824 = array_index_972811 == array_index_948495 ? add_972823 : sel_972820;
  assign add_972827 = sel_972824 + 8'h01;
  assign sel_972828 = array_index_972811 == array_index_948503 ? add_972827 : sel_972824;
  assign add_972831 = sel_972828 + 8'h01;
  assign sel_972832 = array_index_972811 == array_index_948511 ? add_972831 : sel_972828;
  assign add_972835 = sel_972832 + 8'h01;
  assign sel_972836 = array_index_972811 == array_index_948519 ? add_972835 : sel_972832;
  assign add_972839 = sel_972836 + 8'h01;
  assign sel_972840 = array_index_972811 == array_index_948527 ? add_972839 : sel_972836;
  assign add_972843 = sel_972840 + 8'h01;
  assign sel_972844 = array_index_972811 == array_index_948535 ? add_972843 : sel_972840;
  assign add_972847 = sel_972844 + 8'h01;
  assign sel_972848 = array_index_972811 == array_index_948541 ? add_972847 : sel_972844;
  assign add_972851 = sel_972848 + 8'h01;
  assign sel_972852 = array_index_972811 == array_index_948547 ? add_972851 : sel_972848;
  assign add_972855 = sel_972852 + 8'h01;
  assign sel_972856 = array_index_972811 == array_index_948553 ? add_972855 : sel_972852;
  assign add_972859 = sel_972856 + 8'h01;
  assign sel_972860 = array_index_972811 == array_index_948559 ? add_972859 : sel_972856;
  assign add_972863 = sel_972860 + 8'h01;
  assign sel_972864 = array_index_972811 == array_index_948565 ? add_972863 : sel_972860;
  assign add_972867 = sel_972864 + 8'h01;
  assign sel_972868 = array_index_972811 == array_index_948571 ? add_972867 : sel_972864;
  assign add_972871 = sel_972868 + 8'h01;
  assign sel_972872 = array_index_972811 == array_index_948577 ? add_972871 : sel_972868;
  assign add_972875 = sel_972872 + 8'h01;
  assign sel_972876 = array_index_972811 == array_index_948583 ? add_972875 : sel_972872;
  assign add_972879 = sel_972876 + 8'h01;
  assign sel_972880 = array_index_972811 == array_index_948589 ? add_972879 : sel_972876;
  assign add_972883 = sel_972880 + 8'h01;
  assign sel_972884 = array_index_972811 == array_index_948595 ? add_972883 : sel_972880;
  assign add_972887 = sel_972884 + 8'h01;
  assign sel_972888 = array_index_972811 == array_index_948601 ? add_972887 : sel_972884;
  assign add_972891 = sel_972888 + 8'h01;
  assign sel_972892 = array_index_972811 == array_index_948607 ? add_972891 : sel_972888;
  assign add_972895 = sel_972892 + 8'h01;
  assign sel_972896 = array_index_972811 == array_index_948613 ? add_972895 : sel_972892;
  assign add_972899 = sel_972896 + 8'h01;
  assign sel_972900 = array_index_972811 == array_index_948619 ? add_972899 : sel_972896;
  assign add_972903 = sel_972900 + 8'h01;
  assign sel_972904 = array_index_972811 == array_index_948625 ? add_972903 : sel_972900;
  assign add_972907 = sel_972904 + 8'h01;
  assign sel_972908 = array_index_972811 == array_index_948631 ? add_972907 : sel_972904;
  assign add_972911 = sel_972908 + 8'h01;
  assign sel_972912 = array_index_972811 == array_index_948637 ? add_972911 : sel_972908;
  assign add_972915 = sel_972912 + 8'h01;
  assign sel_972916 = array_index_972811 == array_index_948643 ? add_972915 : sel_972912;
  assign add_972919 = sel_972916 + 8'h01;
  assign sel_972920 = array_index_972811 == array_index_948649 ? add_972919 : sel_972916;
  assign add_972923 = sel_972920 + 8'h01;
  assign sel_972924 = array_index_972811 == array_index_948655 ? add_972923 : sel_972920;
  assign add_972927 = sel_972924 + 8'h01;
  assign sel_972928 = array_index_972811 == array_index_948661 ? add_972927 : sel_972924;
  assign add_972931 = sel_972928 + 8'h01;
  assign sel_972932 = array_index_972811 == array_index_948667 ? add_972931 : sel_972928;
  assign add_972935 = sel_972932 + 8'h01;
  assign sel_972936 = array_index_972811 == array_index_948673 ? add_972935 : sel_972932;
  assign add_972939 = sel_972936 + 8'h01;
  assign sel_972940 = array_index_972811 == array_index_948679 ? add_972939 : sel_972936;
  assign add_972943 = sel_972940 + 8'h01;
  assign sel_972944 = array_index_972811 == array_index_948685 ? add_972943 : sel_972940;
  assign add_972947 = sel_972944 + 8'h01;
  assign sel_972948 = array_index_972811 == array_index_948691 ? add_972947 : sel_972944;
  assign add_972951 = sel_972948 + 8'h01;
  assign sel_972952 = array_index_972811 == array_index_948697 ? add_972951 : sel_972948;
  assign add_972955 = sel_972952 + 8'h01;
  assign sel_972956 = array_index_972811 == array_index_948703 ? add_972955 : sel_972952;
  assign add_972959 = sel_972956 + 8'h01;
  assign sel_972960 = array_index_972811 == array_index_948709 ? add_972959 : sel_972956;
  assign add_972963 = sel_972960 + 8'h01;
  assign sel_972964 = array_index_972811 == array_index_948715 ? add_972963 : sel_972960;
  assign add_972967 = sel_972964 + 8'h01;
  assign sel_972968 = array_index_972811 == array_index_948721 ? add_972967 : sel_972964;
  assign add_972971 = sel_972968 + 8'h01;
  assign sel_972972 = array_index_972811 == array_index_948727 ? add_972971 : sel_972968;
  assign add_972975 = sel_972972 + 8'h01;
  assign sel_972976 = array_index_972811 == array_index_948733 ? add_972975 : sel_972972;
  assign add_972979 = sel_972976 + 8'h01;
  assign sel_972980 = array_index_972811 == array_index_948739 ? add_972979 : sel_972976;
  assign add_972983 = sel_972980 + 8'h01;
  assign sel_972984 = array_index_972811 == array_index_948745 ? add_972983 : sel_972980;
  assign add_972987 = sel_972984 + 8'h01;
  assign sel_972988 = array_index_972811 == array_index_948751 ? add_972987 : sel_972984;
  assign add_972991 = sel_972988 + 8'h01;
  assign sel_972992 = array_index_972811 == array_index_948757 ? add_972991 : sel_972988;
  assign add_972995 = sel_972992 + 8'h01;
  assign sel_972996 = array_index_972811 == array_index_948763 ? add_972995 : sel_972992;
  assign add_972999 = sel_972996 + 8'h01;
  assign sel_973000 = array_index_972811 == array_index_948769 ? add_972999 : sel_972996;
  assign add_973003 = sel_973000 + 8'h01;
  assign sel_973004 = array_index_972811 == array_index_948775 ? add_973003 : sel_973000;
  assign add_973007 = sel_973004 + 8'h01;
  assign sel_973008 = array_index_972811 == array_index_948781 ? add_973007 : sel_973004;
  assign add_973011 = sel_973008 + 8'h01;
  assign sel_973012 = array_index_972811 == array_index_948787 ? add_973011 : sel_973008;
  assign add_973015 = sel_973012 + 8'h01;
  assign sel_973016 = array_index_972811 == array_index_948793 ? add_973015 : sel_973012;
  assign add_973019 = sel_973016 + 8'h01;
  assign sel_973020 = array_index_972811 == array_index_948799 ? add_973019 : sel_973016;
  assign add_973023 = sel_973020 + 8'h01;
  assign sel_973024 = array_index_972811 == array_index_948805 ? add_973023 : sel_973020;
  assign add_973027 = sel_973024 + 8'h01;
  assign sel_973028 = array_index_972811 == array_index_948811 ? add_973027 : sel_973024;
  assign add_973031 = sel_973028 + 8'h01;
  assign sel_973032 = array_index_972811 == array_index_948817 ? add_973031 : sel_973028;
  assign add_973035 = sel_973032 + 8'h01;
  assign sel_973036 = array_index_972811 == array_index_948823 ? add_973035 : sel_973032;
  assign add_973039 = sel_973036 + 8'h01;
  assign sel_973040 = array_index_972811 == array_index_948829 ? add_973039 : sel_973036;
  assign add_973043 = sel_973040 + 8'h01;
  assign sel_973044 = array_index_972811 == array_index_948835 ? add_973043 : sel_973040;
  assign add_973047 = sel_973044 + 8'h01;
  assign sel_973048 = array_index_972811 == array_index_948841 ? add_973047 : sel_973044;
  assign add_973051 = sel_973048 + 8'h01;
  assign sel_973052 = array_index_972811 == array_index_948847 ? add_973051 : sel_973048;
  assign add_973055 = sel_973052 + 8'h01;
  assign sel_973056 = array_index_972811 == array_index_948853 ? add_973055 : sel_973052;
  assign add_973059 = sel_973056 + 8'h01;
  assign sel_973060 = array_index_972811 == array_index_948859 ? add_973059 : sel_973056;
  assign add_973063 = sel_973060 + 8'h01;
  assign sel_973064 = array_index_972811 == array_index_948865 ? add_973063 : sel_973060;
  assign add_973067 = sel_973064 + 8'h01;
  assign sel_973068 = array_index_972811 == array_index_948871 ? add_973067 : sel_973064;
  assign add_973071 = sel_973068 + 8'h01;
  assign sel_973072 = array_index_972811 == array_index_948877 ? add_973071 : sel_973068;
  assign add_973075 = sel_973072 + 8'h01;
  assign sel_973076 = array_index_972811 == array_index_948883 ? add_973075 : sel_973072;
  assign add_973079 = sel_973076 + 8'h01;
  assign sel_973080 = array_index_972811 == array_index_948889 ? add_973079 : sel_973076;
  assign add_973083 = sel_973080 + 8'h01;
  assign sel_973084 = array_index_972811 == array_index_948895 ? add_973083 : sel_973080;
  assign add_973087 = sel_973084 + 8'h01;
  assign sel_973088 = array_index_972811 == array_index_948901 ? add_973087 : sel_973084;
  assign add_973091 = sel_973088 + 8'h01;
  assign sel_973092 = array_index_972811 == array_index_948907 ? add_973091 : sel_973088;
  assign add_973095 = sel_973092 + 8'h01;
  assign sel_973096 = array_index_972811 == array_index_948913 ? add_973095 : sel_973092;
  assign add_973099 = sel_973096 + 8'h01;
  assign sel_973100 = array_index_972811 == array_index_948919 ? add_973099 : sel_973096;
  assign add_973103 = sel_973100 + 8'h01;
  assign sel_973104 = array_index_972811 == array_index_948925 ? add_973103 : sel_973100;
  assign add_973107 = sel_973104 + 8'h01;
  assign sel_973108 = array_index_972811 == array_index_948931 ? add_973107 : sel_973104;
  assign add_973111 = sel_973108 + 8'h01;
  assign sel_973112 = array_index_972811 == array_index_948937 ? add_973111 : sel_973108;
  assign add_973115 = sel_973112 + 8'h01;
  assign sel_973116 = array_index_972811 == array_index_948943 ? add_973115 : sel_973112;
  assign add_973119 = sel_973116 + 8'h01;
  assign sel_973120 = array_index_972811 == array_index_948949 ? add_973119 : sel_973116;
  assign add_973123 = sel_973120 + 8'h01;
  assign sel_973124 = array_index_972811 == array_index_948955 ? add_973123 : sel_973120;
  assign add_973127 = sel_973124 + 8'h01;
  assign sel_973128 = array_index_972811 == array_index_948961 ? add_973127 : sel_973124;
  assign add_973131 = sel_973128 + 8'h01;
  assign sel_973132 = array_index_972811 == array_index_948967 ? add_973131 : sel_973128;
  assign add_973135 = sel_973132 + 8'h01;
  assign sel_973136 = array_index_972811 == array_index_948973 ? add_973135 : sel_973132;
  assign add_973139 = sel_973136 + 8'h01;
  assign sel_973140 = array_index_972811 == array_index_948979 ? add_973139 : sel_973136;
  assign add_973143 = sel_973140 + 8'h01;
  assign sel_973144 = array_index_972811 == array_index_948985 ? add_973143 : sel_973140;
  assign add_973147 = sel_973144 + 8'h01;
  assign sel_973148 = array_index_972811 == array_index_948991 ? add_973147 : sel_973144;
  assign add_973151 = sel_973148 + 8'h01;
  assign sel_973152 = array_index_972811 == array_index_948997 ? add_973151 : sel_973148;
  assign add_973155 = sel_973152 + 8'h01;
  assign sel_973156 = array_index_972811 == array_index_949003 ? add_973155 : sel_973152;
  assign add_973159 = sel_973156 + 8'h01;
  assign sel_973160 = array_index_972811 == array_index_949009 ? add_973159 : sel_973156;
  assign add_973163 = sel_973160 + 8'h01;
  assign sel_973164 = array_index_972811 == array_index_949015 ? add_973163 : sel_973160;
  assign add_973167 = sel_973164 + 8'h01;
  assign sel_973168 = array_index_972811 == array_index_949021 ? add_973167 : sel_973164;
  assign add_973171 = sel_973168 + 8'h01;
  assign sel_973172 = array_index_972811 == array_index_949027 ? add_973171 : sel_973168;
  assign add_973175 = sel_973172 + 8'h01;
  assign sel_973176 = array_index_972811 == array_index_949033 ? add_973175 : sel_973172;
  assign add_973179 = sel_973176 + 8'h01;
  assign sel_973180 = array_index_972811 == array_index_949039 ? add_973179 : sel_973176;
  assign add_973183 = sel_973180 + 8'h01;
  assign sel_973184 = array_index_972811 == array_index_949045 ? add_973183 : sel_973180;
  assign add_973187 = sel_973184 + 8'h01;
  assign sel_973188 = array_index_972811 == array_index_949051 ? add_973187 : sel_973184;
  assign add_973191 = sel_973188 + 8'h01;
  assign sel_973192 = array_index_972811 == array_index_949057 ? add_973191 : sel_973188;
  assign add_973195 = sel_973192 + 8'h01;
  assign sel_973196 = array_index_972811 == array_index_949063 ? add_973195 : sel_973192;
  assign add_973199 = sel_973196 + 8'h01;
  assign sel_973200 = array_index_972811 == array_index_949069 ? add_973199 : sel_973196;
  assign add_973203 = sel_973200 + 8'h01;
  assign sel_973204 = array_index_972811 == array_index_949075 ? add_973203 : sel_973200;
  assign add_973207 = sel_973204 + 8'h01;
  assign sel_973208 = array_index_972811 == array_index_949081 ? add_973207 : sel_973204;
  assign add_973212 = sel_973208 + 8'h01;
  assign array_index_973213 = set1_unflattened[7'h3d];
  assign sel_973214 = array_index_972811 == array_index_949087 ? add_973212 : sel_973208;
  assign add_973217 = sel_973214 + 8'h01;
  assign sel_973218 = array_index_973213 == array_index_948483 ? add_973217 : sel_973214;
  assign add_973221 = sel_973218 + 8'h01;
  assign sel_973222 = array_index_973213 == array_index_948487 ? add_973221 : sel_973218;
  assign add_973225 = sel_973222 + 8'h01;
  assign sel_973226 = array_index_973213 == array_index_948495 ? add_973225 : sel_973222;
  assign add_973229 = sel_973226 + 8'h01;
  assign sel_973230 = array_index_973213 == array_index_948503 ? add_973229 : sel_973226;
  assign add_973233 = sel_973230 + 8'h01;
  assign sel_973234 = array_index_973213 == array_index_948511 ? add_973233 : sel_973230;
  assign add_973237 = sel_973234 + 8'h01;
  assign sel_973238 = array_index_973213 == array_index_948519 ? add_973237 : sel_973234;
  assign add_973241 = sel_973238 + 8'h01;
  assign sel_973242 = array_index_973213 == array_index_948527 ? add_973241 : sel_973238;
  assign add_973245 = sel_973242 + 8'h01;
  assign sel_973246 = array_index_973213 == array_index_948535 ? add_973245 : sel_973242;
  assign add_973249 = sel_973246 + 8'h01;
  assign sel_973250 = array_index_973213 == array_index_948541 ? add_973249 : sel_973246;
  assign add_973253 = sel_973250 + 8'h01;
  assign sel_973254 = array_index_973213 == array_index_948547 ? add_973253 : sel_973250;
  assign add_973257 = sel_973254 + 8'h01;
  assign sel_973258 = array_index_973213 == array_index_948553 ? add_973257 : sel_973254;
  assign add_973261 = sel_973258 + 8'h01;
  assign sel_973262 = array_index_973213 == array_index_948559 ? add_973261 : sel_973258;
  assign add_973265 = sel_973262 + 8'h01;
  assign sel_973266 = array_index_973213 == array_index_948565 ? add_973265 : sel_973262;
  assign add_973269 = sel_973266 + 8'h01;
  assign sel_973270 = array_index_973213 == array_index_948571 ? add_973269 : sel_973266;
  assign add_973273 = sel_973270 + 8'h01;
  assign sel_973274 = array_index_973213 == array_index_948577 ? add_973273 : sel_973270;
  assign add_973277 = sel_973274 + 8'h01;
  assign sel_973278 = array_index_973213 == array_index_948583 ? add_973277 : sel_973274;
  assign add_973281 = sel_973278 + 8'h01;
  assign sel_973282 = array_index_973213 == array_index_948589 ? add_973281 : sel_973278;
  assign add_973285 = sel_973282 + 8'h01;
  assign sel_973286 = array_index_973213 == array_index_948595 ? add_973285 : sel_973282;
  assign add_973289 = sel_973286 + 8'h01;
  assign sel_973290 = array_index_973213 == array_index_948601 ? add_973289 : sel_973286;
  assign add_973293 = sel_973290 + 8'h01;
  assign sel_973294 = array_index_973213 == array_index_948607 ? add_973293 : sel_973290;
  assign add_973297 = sel_973294 + 8'h01;
  assign sel_973298 = array_index_973213 == array_index_948613 ? add_973297 : sel_973294;
  assign add_973301 = sel_973298 + 8'h01;
  assign sel_973302 = array_index_973213 == array_index_948619 ? add_973301 : sel_973298;
  assign add_973305 = sel_973302 + 8'h01;
  assign sel_973306 = array_index_973213 == array_index_948625 ? add_973305 : sel_973302;
  assign add_973309 = sel_973306 + 8'h01;
  assign sel_973310 = array_index_973213 == array_index_948631 ? add_973309 : sel_973306;
  assign add_973313 = sel_973310 + 8'h01;
  assign sel_973314 = array_index_973213 == array_index_948637 ? add_973313 : sel_973310;
  assign add_973317 = sel_973314 + 8'h01;
  assign sel_973318 = array_index_973213 == array_index_948643 ? add_973317 : sel_973314;
  assign add_973321 = sel_973318 + 8'h01;
  assign sel_973322 = array_index_973213 == array_index_948649 ? add_973321 : sel_973318;
  assign add_973325 = sel_973322 + 8'h01;
  assign sel_973326 = array_index_973213 == array_index_948655 ? add_973325 : sel_973322;
  assign add_973329 = sel_973326 + 8'h01;
  assign sel_973330 = array_index_973213 == array_index_948661 ? add_973329 : sel_973326;
  assign add_973333 = sel_973330 + 8'h01;
  assign sel_973334 = array_index_973213 == array_index_948667 ? add_973333 : sel_973330;
  assign add_973337 = sel_973334 + 8'h01;
  assign sel_973338 = array_index_973213 == array_index_948673 ? add_973337 : sel_973334;
  assign add_973341 = sel_973338 + 8'h01;
  assign sel_973342 = array_index_973213 == array_index_948679 ? add_973341 : sel_973338;
  assign add_973345 = sel_973342 + 8'h01;
  assign sel_973346 = array_index_973213 == array_index_948685 ? add_973345 : sel_973342;
  assign add_973349 = sel_973346 + 8'h01;
  assign sel_973350 = array_index_973213 == array_index_948691 ? add_973349 : sel_973346;
  assign add_973353 = sel_973350 + 8'h01;
  assign sel_973354 = array_index_973213 == array_index_948697 ? add_973353 : sel_973350;
  assign add_973357 = sel_973354 + 8'h01;
  assign sel_973358 = array_index_973213 == array_index_948703 ? add_973357 : sel_973354;
  assign add_973361 = sel_973358 + 8'h01;
  assign sel_973362 = array_index_973213 == array_index_948709 ? add_973361 : sel_973358;
  assign add_973365 = sel_973362 + 8'h01;
  assign sel_973366 = array_index_973213 == array_index_948715 ? add_973365 : sel_973362;
  assign add_973369 = sel_973366 + 8'h01;
  assign sel_973370 = array_index_973213 == array_index_948721 ? add_973369 : sel_973366;
  assign add_973373 = sel_973370 + 8'h01;
  assign sel_973374 = array_index_973213 == array_index_948727 ? add_973373 : sel_973370;
  assign add_973377 = sel_973374 + 8'h01;
  assign sel_973378 = array_index_973213 == array_index_948733 ? add_973377 : sel_973374;
  assign add_973381 = sel_973378 + 8'h01;
  assign sel_973382 = array_index_973213 == array_index_948739 ? add_973381 : sel_973378;
  assign add_973385 = sel_973382 + 8'h01;
  assign sel_973386 = array_index_973213 == array_index_948745 ? add_973385 : sel_973382;
  assign add_973389 = sel_973386 + 8'h01;
  assign sel_973390 = array_index_973213 == array_index_948751 ? add_973389 : sel_973386;
  assign add_973393 = sel_973390 + 8'h01;
  assign sel_973394 = array_index_973213 == array_index_948757 ? add_973393 : sel_973390;
  assign add_973397 = sel_973394 + 8'h01;
  assign sel_973398 = array_index_973213 == array_index_948763 ? add_973397 : sel_973394;
  assign add_973401 = sel_973398 + 8'h01;
  assign sel_973402 = array_index_973213 == array_index_948769 ? add_973401 : sel_973398;
  assign add_973405 = sel_973402 + 8'h01;
  assign sel_973406 = array_index_973213 == array_index_948775 ? add_973405 : sel_973402;
  assign add_973409 = sel_973406 + 8'h01;
  assign sel_973410 = array_index_973213 == array_index_948781 ? add_973409 : sel_973406;
  assign add_973413 = sel_973410 + 8'h01;
  assign sel_973414 = array_index_973213 == array_index_948787 ? add_973413 : sel_973410;
  assign add_973417 = sel_973414 + 8'h01;
  assign sel_973418 = array_index_973213 == array_index_948793 ? add_973417 : sel_973414;
  assign add_973421 = sel_973418 + 8'h01;
  assign sel_973422 = array_index_973213 == array_index_948799 ? add_973421 : sel_973418;
  assign add_973425 = sel_973422 + 8'h01;
  assign sel_973426 = array_index_973213 == array_index_948805 ? add_973425 : sel_973422;
  assign add_973429 = sel_973426 + 8'h01;
  assign sel_973430 = array_index_973213 == array_index_948811 ? add_973429 : sel_973426;
  assign add_973433 = sel_973430 + 8'h01;
  assign sel_973434 = array_index_973213 == array_index_948817 ? add_973433 : sel_973430;
  assign add_973437 = sel_973434 + 8'h01;
  assign sel_973438 = array_index_973213 == array_index_948823 ? add_973437 : sel_973434;
  assign add_973441 = sel_973438 + 8'h01;
  assign sel_973442 = array_index_973213 == array_index_948829 ? add_973441 : sel_973438;
  assign add_973445 = sel_973442 + 8'h01;
  assign sel_973446 = array_index_973213 == array_index_948835 ? add_973445 : sel_973442;
  assign add_973449 = sel_973446 + 8'h01;
  assign sel_973450 = array_index_973213 == array_index_948841 ? add_973449 : sel_973446;
  assign add_973453 = sel_973450 + 8'h01;
  assign sel_973454 = array_index_973213 == array_index_948847 ? add_973453 : sel_973450;
  assign add_973457 = sel_973454 + 8'h01;
  assign sel_973458 = array_index_973213 == array_index_948853 ? add_973457 : sel_973454;
  assign add_973461 = sel_973458 + 8'h01;
  assign sel_973462 = array_index_973213 == array_index_948859 ? add_973461 : sel_973458;
  assign add_973465 = sel_973462 + 8'h01;
  assign sel_973466 = array_index_973213 == array_index_948865 ? add_973465 : sel_973462;
  assign add_973469 = sel_973466 + 8'h01;
  assign sel_973470 = array_index_973213 == array_index_948871 ? add_973469 : sel_973466;
  assign add_973473 = sel_973470 + 8'h01;
  assign sel_973474 = array_index_973213 == array_index_948877 ? add_973473 : sel_973470;
  assign add_973477 = sel_973474 + 8'h01;
  assign sel_973478 = array_index_973213 == array_index_948883 ? add_973477 : sel_973474;
  assign add_973481 = sel_973478 + 8'h01;
  assign sel_973482 = array_index_973213 == array_index_948889 ? add_973481 : sel_973478;
  assign add_973485 = sel_973482 + 8'h01;
  assign sel_973486 = array_index_973213 == array_index_948895 ? add_973485 : sel_973482;
  assign add_973489 = sel_973486 + 8'h01;
  assign sel_973490 = array_index_973213 == array_index_948901 ? add_973489 : sel_973486;
  assign add_973493 = sel_973490 + 8'h01;
  assign sel_973494 = array_index_973213 == array_index_948907 ? add_973493 : sel_973490;
  assign add_973497 = sel_973494 + 8'h01;
  assign sel_973498 = array_index_973213 == array_index_948913 ? add_973497 : sel_973494;
  assign add_973501 = sel_973498 + 8'h01;
  assign sel_973502 = array_index_973213 == array_index_948919 ? add_973501 : sel_973498;
  assign add_973505 = sel_973502 + 8'h01;
  assign sel_973506 = array_index_973213 == array_index_948925 ? add_973505 : sel_973502;
  assign add_973509 = sel_973506 + 8'h01;
  assign sel_973510 = array_index_973213 == array_index_948931 ? add_973509 : sel_973506;
  assign add_973513 = sel_973510 + 8'h01;
  assign sel_973514 = array_index_973213 == array_index_948937 ? add_973513 : sel_973510;
  assign add_973517 = sel_973514 + 8'h01;
  assign sel_973518 = array_index_973213 == array_index_948943 ? add_973517 : sel_973514;
  assign add_973521 = sel_973518 + 8'h01;
  assign sel_973522 = array_index_973213 == array_index_948949 ? add_973521 : sel_973518;
  assign add_973525 = sel_973522 + 8'h01;
  assign sel_973526 = array_index_973213 == array_index_948955 ? add_973525 : sel_973522;
  assign add_973529 = sel_973526 + 8'h01;
  assign sel_973530 = array_index_973213 == array_index_948961 ? add_973529 : sel_973526;
  assign add_973533 = sel_973530 + 8'h01;
  assign sel_973534 = array_index_973213 == array_index_948967 ? add_973533 : sel_973530;
  assign add_973537 = sel_973534 + 8'h01;
  assign sel_973538 = array_index_973213 == array_index_948973 ? add_973537 : sel_973534;
  assign add_973541 = sel_973538 + 8'h01;
  assign sel_973542 = array_index_973213 == array_index_948979 ? add_973541 : sel_973538;
  assign add_973545 = sel_973542 + 8'h01;
  assign sel_973546 = array_index_973213 == array_index_948985 ? add_973545 : sel_973542;
  assign add_973549 = sel_973546 + 8'h01;
  assign sel_973550 = array_index_973213 == array_index_948991 ? add_973549 : sel_973546;
  assign add_973553 = sel_973550 + 8'h01;
  assign sel_973554 = array_index_973213 == array_index_948997 ? add_973553 : sel_973550;
  assign add_973557 = sel_973554 + 8'h01;
  assign sel_973558 = array_index_973213 == array_index_949003 ? add_973557 : sel_973554;
  assign add_973561 = sel_973558 + 8'h01;
  assign sel_973562 = array_index_973213 == array_index_949009 ? add_973561 : sel_973558;
  assign add_973565 = sel_973562 + 8'h01;
  assign sel_973566 = array_index_973213 == array_index_949015 ? add_973565 : sel_973562;
  assign add_973569 = sel_973566 + 8'h01;
  assign sel_973570 = array_index_973213 == array_index_949021 ? add_973569 : sel_973566;
  assign add_973573 = sel_973570 + 8'h01;
  assign sel_973574 = array_index_973213 == array_index_949027 ? add_973573 : sel_973570;
  assign add_973577 = sel_973574 + 8'h01;
  assign sel_973578 = array_index_973213 == array_index_949033 ? add_973577 : sel_973574;
  assign add_973581 = sel_973578 + 8'h01;
  assign sel_973582 = array_index_973213 == array_index_949039 ? add_973581 : sel_973578;
  assign add_973585 = sel_973582 + 8'h01;
  assign sel_973586 = array_index_973213 == array_index_949045 ? add_973585 : sel_973582;
  assign add_973589 = sel_973586 + 8'h01;
  assign sel_973590 = array_index_973213 == array_index_949051 ? add_973589 : sel_973586;
  assign add_973593 = sel_973590 + 8'h01;
  assign sel_973594 = array_index_973213 == array_index_949057 ? add_973593 : sel_973590;
  assign add_973597 = sel_973594 + 8'h01;
  assign sel_973598 = array_index_973213 == array_index_949063 ? add_973597 : sel_973594;
  assign add_973601 = sel_973598 + 8'h01;
  assign sel_973602 = array_index_973213 == array_index_949069 ? add_973601 : sel_973598;
  assign add_973605 = sel_973602 + 8'h01;
  assign sel_973606 = array_index_973213 == array_index_949075 ? add_973605 : sel_973602;
  assign add_973609 = sel_973606 + 8'h01;
  assign sel_973610 = array_index_973213 == array_index_949081 ? add_973609 : sel_973606;
  assign add_973614 = sel_973610 + 8'h01;
  assign array_index_973615 = set1_unflattened[7'h3e];
  assign sel_973616 = array_index_973213 == array_index_949087 ? add_973614 : sel_973610;
  assign add_973619 = sel_973616 + 8'h01;
  assign sel_973620 = array_index_973615 == array_index_948483 ? add_973619 : sel_973616;
  assign add_973623 = sel_973620 + 8'h01;
  assign sel_973624 = array_index_973615 == array_index_948487 ? add_973623 : sel_973620;
  assign add_973627 = sel_973624 + 8'h01;
  assign sel_973628 = array_index_973615 == array_index_948495 ? add_973627 : sel_973624;
  assign add_973631 = sel_973628 + 8'h01;
  assign sel_973632 = array_index_973615 == array_index_948503 ? add_973631 : sel_973628;
  assign add_973635 = sel_973632 + 8'h01;
  assign sel_973636 = array_index_973615 == array_index_948511 ? add_973635 : sel_973632;
  assign add_973639 = sel_973636 + 8'h01;
  assign sel_973640 = array_index_973615 == array_index_948519 ? add_973639 : sel_973636;
  assign add_973643 = sel_973640 + 8'h01;
  assign sel_973644 = array_index_973615 == array_index_948527 ? add_973643 : sel_973640;
  assign add_973647 = sel_973644 + 8'h01;
  assign sel_973648 = array_index_973615 == array_index_948535 ? add_973647 : sel_973644;
  assign add_973651 = sel_973648 + 8'h01;
  assign sel_973652 = array_index_973615 == array_index_948541 ? add_973651 : sel_973648;
  assign add_973655 = sel_973652 + 8'h01;
  assign sel_973656 = array_index_973615 == array_index_948547 ? add_973655 : sel_973652;
  assign add_973659 = sel_973656 + 8'h01;
  assign sel_973660 = array_index_973615 == array_index_948553 ? add_973659 : sel_973656;
  assign add_973663 = sel_973660 + 8'h01;
  assign sel_973664 = array_index_973615 == array_index_948559 ? add_973663 : sel_973660;
  assign add_973667 = sel_973664 + 8'h01;
  assign sel_973668 = array_index_973615 == array_index_948565 ? add_973667 : sel_973664;
  assign add_973671 = sel_973668 + 8'h01;
  assign sel_973672 = array_index_973615 == array_index_948571 ? add_973671 : sel_973668;
  assign add_973675 = sel_973672 + 8'h01;
  assign sel_973676 = array_index_973615 == array_index_948577 ? add_973675 : sel_973672;
  assign add_973679 = sel_973676 + 8'h01;
  assign sel_973680 = array_index_973615 == array_index_948583 ? add_973679 : sel_973676;
  assign add_973683 = sel_973680 + 8'h01;
  assign sel_973684 = array_index_973615 == array_index_948589 ? add_973683 : sel_973680;
  assign add_973687 = sel_973684 + 8'h01;
  assign sel_973688 = array_index_973615 == array_index_948595 ? add_973687 : sel_973684;
  assign add_973691 = sel_973688 + 8'h01;
  assign sel_973692 = array_index_973615 == array_index_948601 ? add_973691 : sel_973688;
  assign add_973695 = sel_973692 + 8'h01;
  assign sel_973696 = array_index_973615 == array_index_948607 ? add_973695 : sel_973692;
  assign add_973699 = sel_973696 + 8'h01;
  assign sel_973700 = array_index_973615 == array_index_948613 ? add_973699 : sel_973696;
  assign add_973703 = sel_973700 + 8'h01;
  assign sel_973704 = array_index_973615 == array_index_948619 ? add_973703 : sel_973700;
  assign add_973707 = sel_973704 + 8'h01;
  assign sel_973708 = array_index_973615 == array_index_948625 ? add_973707 : sel_973704;
  assign add_973711 = sel_973708 + 8'h01;
  assign sel_973712 = array_index_973615 == array_index_948631 ? add_973711 : sel_973708;
  assign add_973715 = sel_973712 + 8'h01;
  assign sel_973716 = array_index_973615 == array_index_948637 ? add_973715 : sel_973712;
  assign add_973719 = sel_973716 + 8'h01;
  assign sel_973720 = array_index_973615 == array_index_948643 ? add_973719 : sel_973716;
  assign add_973723 = sel_973720 + 8'h01;
  assign sel_973724 = array_index_973615 == array_index_948649 ? add_973723 : sel_973720;
  assign add_973727 = sel_973724 + 8'h01;
  assign sel_973728 = array_index_973615 == array_index_948655 ? add_973727 : sel_973724;
  assign add_973731 = sel_973728 + 8'h01;
  assign sel_973732 = array_index_973615 == array_index_948661 ? add_973731 : sel_973728;
  assign add_973735 = sel_973732 + 8'h01;
  assign sel_973736 = array_index_973615 == array_index_948667 ? add_973735 : sel_973732;
  assign add_973739 = sel_973736 + 8'h01;
  assign sel_973740 = array_index_973615 == array_index_948673 ? add_973739 : sel_973736;
  assign add_973743 = sel_973740 + 8'h01;
  assign sel_973744 = array_index_973615 == array_index_948679 ? add_973743 : sel_973740;
  assign add_973747 = sel_973744 + 8'h01;
  assign sel_973748 = array_index_973615 == array_index_948685 ? add_973747 : sel_973744;
  assign add_973751 = sel_973748 + 8'h01;
  assign sel_973752 = array_index_973615 == array_index_948691 ? add_973751 : sel_973748;
  assign add_973755 = sel_973752 + 8'h01;
  assign sel_973756 = array_index_973615 == array_index_948697 ? add_973755 : sel_973752;
  assign add_973759 = sel_973756 + 8'h01;
  assign sel_973760 = array_index_973615 == array_index_948703 ? add_973759 : sel_973756;
  assign add_973763 = sel_973760 + 8'h01;
  assign sel_973764 = array_index_973615 == array_index_948709 ? add_973763 : sel_973760;
  assign add_973767 = sel_973764 + 8'h01;
  assign sel_973768 = array_index_973615 == array_index_948715 ? add_973767 : sel_973764;
  assign add_973771 = sel_973768 + 8'h01;
  assign sel_973772 = array_index_973615 == array_index_948721 ? add_973771 : sel_973768;
  assign add_973775 = sel_973772 + 8'h01;
  assign sel_973776 = array_index_973615 == array_index_948727 ? add_973775 : sel_973772;
  assign add_973779 = sel_973776 + 8'h01;
  assign sel_973780 = array_index_973615 == array_index_948733 ? add_973779 : sel_973776;
  assign add_973783 = sel_973780 + 8'h01;
  assign sel_973784 = array_index_973615 == array_index_948739 ? add_973783 : sel_973780;
  assign add_973787 = sel_973784 + 8'h01;
  assign sel_973788 = array_index_973615 == array_index_948745 ? add_973787 : sel_973784;
  assign add_973791 = sel_973788 + 8'h01;
  assign sel_973792 = array_index_973615 == array_index_948751 ? add_973791 : sel_973788;
  assign add_973795 = sel_973792 + 8'h01;
  assign sel_973796 = array_index_973615 == array_index_948757 ? add_973795 : sel_973792;
  assign add_973799 = sel_973796 + 8'h01;
  assign sel_973800 = array_index_973615 == array_index_948763 ? add_973799 : sel_973796;
  assign add_973803 = sel_973800 + 8'h01;
  assign sel_973804 = array_index_973615 == array_index_948769 ? add_973803 : sel_973800;
  assign add_973807 = sel_973804 + 8'h01;
  assign sel_973808 = array_index_973615 == array_index_948775 ? add_973807 : sel_973804;
  assign add_973811 = sel_973808 + 8'h01;
  assign sel_973812 = array_index_973615 == array_index_948781 ? add_973811 : sel_973808;
  assign add_973815 = sel_973812 + 8'h01;
  assign sel_973816 = array_index_973615 == array_index_948787 ? add_973815 : sel_973812;
  assign add_973819 = sel_973816 + 8'h01;
  assign sel_973820 = array_index_973615 == array_index_948793 ? add_973819 : sel_973816;
  assign add_973823 = sel_973820 + 8'h01;
  assign sel_973824 = array_index_973615 == array_index_948799 ? add_973823 : sel_973820;
  assign add_973827 = sel_973824 + 8'h01;
  assign sel_973828 = array_index_973615 == array_index_948805 ? add_973827 : sel_973824;
  assign add_973831 = sel_973828 + 8'h01;
  assign sel_973832 = array_index_973615 == array_index_948811 ? add_973831 : sel_973828;
  assign add_973835 = sel_973832 + 8'h01;
  assign sel_973836 = array_index_973615 == array_index_948817 ? add_973835 : sel_973832;
  assign add_973839 = sel_973836 + 8'h01;
  assign sel_973840 = array_index_973615 == array_index_948823 ? add_973839 : sel_973836;
  assign add_973843 = sel_973840 + 8'h01;
  assign sel_973844 = array_index_973615 == array_index_948829 ? add_973843 : sel_973840;
  assign add_973847 = sel_973844 + 8'h01;
  assign sel_973848 = array_index_973615 == array_index_948835 ? add_973847 : sel_973844;
  assign add_973851 = sel_973848 + 8'h01;
  assign sel_973852 = array_index_973615 == array_index_948841 ? add_973851 : sel_973848;
  assign add_973855 = sel_973852 + 8'h01;
  assign sel_973856 = array_index_973615 == array_index_948847 ? add_973855 : sel_973852;
  assign add_973859 = sel_973856 + 8'h01;
  assign sel_973860 = array_index_973615 == array_index_948853 ? add_973859 : sel_973856;
  assign add_973863 = sel_973860 + 8'h01;
  assign sel_973864 = array_index_973615 == array_index_948859 ? add_973863 : sel_973860;
  assign add_973867 = sel_973864 + 8'h01;
  assign sel_973868 = array_index_973615 == array_index_948865 ? add_973867 : sel_973864;
  assign add_973871 = sel_973868 + 8'h01;
  assign sel_973872 = array_index_973615 == array_index_948871 ? add_973871 : sel_973868;
  assign add_973875 = sel_973872 + 8'h01;
  assign sel_973876 = array_index_973615 == array_index_948877 ? add_973875 : sel_973872;
  assign add_973879 = sel_973876 + 8'h01;
  assign sel_973880 = array_index_973615 == array_index_948883 ? add_973879 : sel_973876;
  assign add_973883 = sel_973880 + 8'h01;
  assign sel_973884 = array_index_973615 == array_index_948889 ? add_973883 : sel_973880;
  assign add_973887 = sel_973884 + 8'h01;
  assign sel_973888 = array_index_973615 == array_index_948895 ? add_973887 : sel_973884;
  assign add_973891 = sel_973888 + 8'h01;
  assign sel_973892 = array_index_973615 == array_index_948901 ? add_973891 : sel_973888;
  assign add_973895 = sel_973892 + 8'h01;
  assign sel_973896 = array_index_973615 == array_index_948907 ? add_973895 : sel_973892;
  assign add_973899 = sel_973896 + 8'h01;
  assign sel_973900 = array_index_973615 == array_index_948913 ? add_973899 : sel_973896;
  assign add_973903 = sel_973900 + 8'h01;
  assign sel_973904 = array_index_973615 == array_index_948919 ? add_973903 : sel_973900;
  assign add_973907 = sel_973904 + 8'h01;
  assign sel_973908 = array_index_973615 == array_index_948925 ? add_973907 : sel_973904;
  assign add_973911 = sel_973908 + 8'h01;
  assign sel_973912 = array_index_973615 == array_index_948931 ? add_973911 : sel_973908;
  assign add_973915 = sel_973912 + 8'h01;
  assign sel_973916 = array_index_973615 == array_index_948937 ? add_973915 : sel_973912;
  assign add_973919 = sel_973916 + 8'h01;
  assign sel_973920 = array_index_973615 == array_index_948943 ? add_973919 : sel_973916;
  assign add_973923 = sel_973920 + 8'h01;
  assign sel_973924 = array_index_973615 == array_index_948949 ? add_973923 : sel_973920;
  assign add_973927 = sel_973924 + 8'h01;
  assign sel_973928 = array_index_973615 == array_index_948955 ? add_973927 : sel_973924;
  assign add_973931 = sel_973928 + 8'h01;
  assign sel_973932 = array_index_973615 == array_index_948961 ? add_973931 : sel_973928;
  assign add_973935 = sel_973932 + 8'h01;
  assign sel_973936 = array_index_973615 == array_index_948967 ? add_973935 : sel_973932;
  assign add_973939 = sel_973936 + 8'h01;
  assign sel_973940 = array_index_973615 == array_index_948973 ? add_973939 : sel_973936;
  assign add_973943 = sel_973940 + 8'h01;
  assign sel_973944 = array_index_973615 == array_index_948979 ? add_973943 : sel_973940;
  assign add_973947 = sel_973944 + 8'h01;
  assign sel_973948 = array_index_973615 == array_index_948985 ? add_973947 : sel_973944;
  assign add_973951 = sel_973948 + 8'h01;
  assign sel_973952 = array_index_973615 == array_index_948991 ? add_973951 : sel_973948;
  assign add_973955 = sel_973952 + 8'h01;
  assign sel_973956 = array_index_973615 == array_index_948997 ? add_973955 : sel_973952;
  assign add_973959 = sel_973956 + 8'h01;
  assign sel_973960 = array_index_973615 == array_index_949003 ? add_973959 : sel_973956;
  assign add_973963 = sel_973960 + 8'h01;
  assign sel_973964 = array_index_973615 == array_index_949009 ? add_973963 : sel_973960;
  assign add_973967 = sel_973964 + 8'h01;
  assign sel_973968 = array_index_973615 == array_index_949015 ? add_973967 : sel_973964;
  assign add_973971 = sel_973968 + 8'h01;
  assign sel_973972 = array_index_973615 == array_index_949021 ? add_973971 : sel_973968;
  assign add_973975 = sel_973972 + 8'h01;
  assign sel_973976 = array_index_973615 == array_index_949027 ? add_973975 : sel_973972;
  assign add_973979 = sel_973976 + 8'h01;
  assign sel_973980 = array_index_973615 == array_index_949033 ? add_973979 : sel_973976;
  assign add_973983 = sel_973980 + 8'h01;
  assign sel_973984 = array_index_973615 == array_index_949039 ? add_973983 : sel_973980;
  assign add_973987 = sel_973984 + 8'h01;
  assign sel_973988 = array_index_973615 == array_index_949045 ? add_973987 : sel_973984;
  assign add_973991 = sel_973988 + 8'h01;
  assign sel_973992 = array_index_973615 == array_index_949051 ? add_973991 : sel_973988;
  assign add_973995 = sel_973992 + 8'h01;
  assign sel_973996 = array_index_973615 == array_index_949057 ? add_973995 : sel_973992;
  assign add_973999 = sel_973996 + 8'h01;
  assign sel_974000 = array_index_973615 == array_index_949063 ? add_973999 : sel_973996;
  assign add_974003 = sel_974000 + 8'h01;
  assign sel_974004 = array_index_973615 == array_index_949069 ? add_974003 : sel_974000;
  assign add_974007 = sel_974004 + 8'h01;
  assign sel_974008 = array_index_973615 == array_index_949075 ? add_974007 : sel_974004;
  assign add_974011 = sel_974008 + 8'h01;
  assign sel_974012 = array_index_973615 == array_index_949081 ? add_974011 : sel_974008;
  assign add_974016 = sel_974012 + 8'h01;
  assign array_index_974017 = set1_unflattened[7'h3f];
  assign sel_974018 = array_index_973615 == array_index_949087 ? add_974016 : sel_974012;
  assign add_974021 = sel_974018 + 8'h01;
  assign sel_974022 = array_index_974017 == array_index_948483 ? add_974021 : sel_974018;
  assign add_974025 = sel_974022 + 8'h01;
  assign sel_974026 = array_index_974017 == array_index_948487 ? add_974025 : sel_974022;
  assign add_974029 = sel_974026 + 8'h01;
  assign sel_974030 = array_index_974017 == array_index_948495 ? add_974029 : sel_974026;
  assign add_974033 = sel_974030 + 8'h01;
  assign sel_974034 = array_index_974017 == array_index_948503 ? add_974033 : sel_974030;
  assign add_974037 = sel_974034 + 8'h01;
  assign sel_974038 = array_index_974017 == array_index_948511 ? add_974037 : sel_974034;
  assign add_974041 = sel_974038 + 8'h01;
  assign sel_974042 = array_index_974017 == array_index_948519 ? add_974041 : sel_974038;
  assign add_974045 = sel_974042 + 8'h01;
  assign sel_974046 = array_index_974017 == array_index_948527 ? add_974045 : sel_974042;
  assign add_974049 = sel_974046 + 8'h01;
  assign sel_974050 = array_index_974017 == array_index_948535 ? add_974049 : sel_974046;
  assign add_974053 = sel_974050 + 8'h01;
  assign sel_974054 = array_index_974017 == array_index_948541 ? add_974053 : sel_974050;
  assign add_974057 = sel_974054 + 8'h01;
  assign sel_974058 = array_index_974017 == array_index_948547 ? add_974057 : sel_974054;
  assign add_974061 = sel_974058 + 8'h01;
  assign sel_974062 = array_index_974017 == array_index_948553 ? add_974061 : sel_974058;
  assign add_974065 = sel_974062 + 8'h01;
  assign sel_974066 = array_index_974017 == array_index_948559 ? add_974065 : sel_974062;
  assign add_974069 = sel_974066 + 8'h01;
  assign sel_974070 = array_index_974017 == array_index_948565 ? add_974069 : sel_974066;
  assign add_974073 = sel_974070 + 8'h01;
  assign sel_974074 = array_index_974017 == array_index_948571 ? add_974073 : sel_974070;
  assign add_974077 = sel_974074 + 8'h01;
  assign sel_974078 = array_index_974017 == array_index_948577 ? add_974077 : sel_974074;
  assign add_974081 = sel_974078 + 8'h01;
  assign sel_974082 = array_index_974017 == array_index_948583 ? add_974081 : sel_974078;
  assign add_974085 = sel_974082 + 8'h01;
  assign sel_974086 = array_index_974017 == array_index_948589 ? add_974085 : sel_974082;
  assign add_974089 = sel_974086 + 8'h01;
  assign sel_974090 = array_index_974017 == array_index_948595 ? add_974089 : sel_974086;
  assign add_974093 = sel_974090 + 8'h01;
  assign sel_974094 = array_index_974017 == array_index_948601 ? add_974093 : sel_974090;
  assign add_974097 = sel_974094 + 8'h01;
  assign sel_974098 = array_index_974017 == array_index_948607 ? add_974097 : sel_974094;
  assign add_974101 = sel_974098 + 8'h01;
  assign sel_974102 = array_index_974017 == array_index_948613 ? add_974101 : sel_974098;
  assign add_974105 = sel_974102 + 8'h01;
  assign sel_974106 = array_index_974017 == array_index_948619 ? add_974105 : sel_974102;
  assign add_974109 = sel_974106 + 8'h01;
  assign sel_974110 = array_index_974017 == array_index_948625 ? add_974109 : sel_974106;
  assign add_974113 = sel_974110 + 8'h01;
  assign sel_974114 = array_index_974017 == array_index_948631 ? add_974113 : sel_974110;
  assign add_974117 = sel_974114 + 8'h01;
  assign sel_974118 = array_index_974017 == array_index_948637 ? add_974117 : sel_974114;
  assign add_974121 = sel_974118 + 8'h01;
  assign sel_974122 = array_index_974017 == array_index_948643 ? add_974121 : sel_974118;
  assign add_974125 = sel_974122 + 8'h01;
  assign sel_974126 = array_index_974017 == array_index_948649 ? add_974125 : sel_974122;
  assign add_974129 = sel_974126 + 8'h01;
  assign sel_974130 = array_index_974017 == array_index_948655 ? add_974129 : sel_974126;
  assign add_974133 = sel_974130 + 8'h01;
  assign sel_974134 = array_index_974017 == array_index_948661 ? add_974133 : sel_974130;
  assign add_974137 = sel_974134 + 8'h01;
  assign sel_974138 = array_index_974017 == array_index_948667 ? add_974137 : sel_974134;
  assign add_974141 = sel_974138 + 8'h01;
  assign sel_974142 = array_index_974017 == array_index_948673 ? add_974141 : sel_974138;
  assign add_974145 = sel_974142 + 8'h01;
  assign sel_974146 = array_index_974017 == array_index_948679 ? add_974145 : sel_974142;
  assign add_974149 = sel_974146 + 8'h01;
  assign sel_974150 = array_index_974017 == array_index_948685 ? add_974149 : sel_974146;
  assign add_974153 = sel_974150 + 8'h01;
  assign sel_974154 = array_index_974017 == array_index_948691 ? add_974153 : sel_974150;
  assign add_974157 = sel_974154 + 8'h01;
  assign sel_974158 = array_index_974017 == array_index_948697 ? add_974157 : sel_974154;
  assign add_974161 = sel_974158 + 8'h01;
  assign sel_974162 = array_index_974017 == array_index_948703 ? add_974161 : sel_974158;
  assign add_974165 = sel_974162 + 8'h01;
  assign sel_974166 = array_index_974017 == array_index_948709 ? add_974165 : sel_974162;
  assign add_974169 = sel_974166 + 8'h01;
  assign sel_974170 = array_index_974017 == array_index_948715 ? add_974169 : sel_974166;
  assign add_974173 = sel_974170 + 8'h01;
  assign sel_974174 = array_index_974017 == array_index_948721 ? add_974173 : sel_974170;
  assign add_974177 = sel_974174 + 8'h01;
  assign sel_974178 = array_index_974017 == array_index_948727 ? add_974177 : sel_974174;
  assign add_974181 = sel_974178 + 8'h01;
  assign sel_974182 = array_index_974017 == array_index_948733 ? add_974181 : sel_974178;
  assign add_974185 = sel_974182 + 8'h01;
  assign sel_974186 = array_index_974017 == array_index_948739 ? add_974185 : sel_974182;
  assign add_974189 = sel_974186 + 8'h01;
  assign sel_974190 = array_index_974017 == array_index_948745 ? add_974189 : sel_974186;
  assign add_974193 = sel_974190 + 8'h01;
  assign sel_974194 = array_index_974017 == array_index_948751 ? add_974193 : sel_974190;
  assign add_974197 = sel_974194 + 8'h01;
  assign sel_974198 = array_index_974017 == array_index_948757 ? add_974197 : sel_974194;
  assign add_974201 = sel_974198 + 8'h01;
  assign sel_974202 = array_index_974017 == array_index_948763 ? add_974201 : sel_974198;
  assign add_974205 = sel_974202 + 8'h01;
  assign sel_974206 = array_index_974017 == array_index_948769 ? add_974205 : sel_974202;
  assign add_974209 = sel_974206 + 8'h01;
  assign sel_974210 = array_index_974017 == array_index_948775 ? add_974209 : sel_974206;
  assign add_974213 = sel_974210 + 8'h01;
  assign sel_974214 = array_index_974017 == array_index_948781 ? add_974213 : sel_974210;
  assign add_974217 = sel_974214 + 8'h01;
  assign sel_974218 = array_index_974017 == array_index_948787 ? add_974217 : sel_974214;
  assign add_974221 = sel_974218 + 8'h01;
  assign sel_974222 = array_index_974017 == array_index_948793 ? add_974221 : sel_974218;
  assign add_974225 = sel_974222 + 8'h01;
  assign sel_974226 = array_index_974017 == array_index_948799 ? add_974225 : sel_974222;
  assign add_974229 = sel_974226 + 8'h01;
  assign sel_974230 = array_index_974017 == array_index_948805 ? add_974229 : sel_974226;
  assign add_974233 = sel_974230 + 8'h01;
  assign sel_974234 = array_index_974017 == array_index_948811 ? add_974233 : sel_974230;
  assign add_974237 = sel_974234 + 8'h01;
  assign sel_974238 = array_index_974017 == array_index_948817 ? add_974237 : sel_974234;
  assign add_974241 = sel_974238 + 8'h01;
  assign sel_974242 = array_index_974017 == array_index_948823 ? add_974241 : sel_974238;
  assign add_974245 = sel_974242 + 8'h01;
  assign sel_974246 = array_index_974017 == array_index_948829 ? add_974245 : sel_974242;
  assign add_974249 = sel_974246 + 8'h01;
  assign sel_974250 = array_index_974017 == array_index_948835 ? add_974249 : sel_974246;
  assign add_974253 = sel_974250 + 8'h01;
  assign sel_974254 = array_index_974017 == array_index_948841 ? add_974253 : sel_974250;
  assign add_974257 = sel_974254 + 8'h01;
  assign sel_974258 = array_index_974017 == array_index_948847 ? add_974257 : sel_974254;
  assign add_974261 = sel_974258 + 8'h01;
  assign sel_974262 = array_index_974017 == array_index_948853 ? add_974261 : sel_974258;
  assign add_974265 = sel_974262 + 8'h01;
  assign sel_974266 = array_index_974017 == array_index_948859 ? add_974265 : sel_974262;
  assign add_974269 = sel_974266 + 8'h01;
  assign sel_974270 = array_index_974017 == array_index_948865 ? add_974269 : sel_974266;
  assign add_974273 = sel_974270 + 8'h01;
  assign sel_974274 = array_index_974017 == array_index_948871 ? add_974273 : sel_974270;
  assign add_974277 = sel_974274 + 8'h01;
  assign sel_974278 = array_index_974017 == array_index_948877 ? add_974277 : sel_974274;
  assign add_974281 = sel_974278 + 8'h01;
  assign sel_974282 = array_index_974017 == array_index_948883 ? add_974281 : sel_974278;
  assign add_974285 = sel_974282 + 8'h01;
  assign sel_974286 = array_index_974017 == array_index_948889 ? add_974285 : sel_974282;
  assign add_974289 = sel_974286 + 8'h01;
  assign sel_974290 = array_index_974017 == array_index_948895 ? add_974289 : sel_974286;
  assign add_974293 = sel_974290 + 8'h01;
  assign sel_974294 = array_index_974017 == array_index_948901 ? add_974293 : sel_974290;
  assign add_974297 = sel_974294 + 8'h01;
  assign sel_974298 = array_index_974017 == array_index_948907 ? add_974297 : sel_974294;
  assign add_974301 = sel_974298 + 8'h01;
  assign sel_974302 = array_index_974017 == array_index_948913 ? add_974301 : sel_974298;
  assign add_974305 = sel_974302 + 8'h01;
  assign sel_974306 = array_index_974017 == array_index_948919 ? add_974305 : sel_974302;
  assign add_974309 = sel_974306 + 8'h01;
  assign sel_974310 = array_index_974017 == array_index_948925 ? add_974309 : sel_974306;
  assign add_974313 = sel_974310 + 8'h01;
  assign sel_974314 = array_index_974017 == array_index_948931 ? add_974313 : sel_974310;
  assign add_974317 = sel_974314 + 8'h01;
  assign sel_974318 = array_index_974017 == array_index_948937 ? add_974317 : sel_974314;
  assign add_974321 = sel_974318 + 8'h01;
  assign sel_974322 = array_index_974017 == array_index_948943 ? add_974321 : sel_974318;
  assign add_974325 = sel_974322 + 8'h01;
  assign sel_974326 = array_index_974017 == array_index_948949 ? add_974325 : sel_974322;
  assign add_974329 = sel_974326 + 8'h01;
  assign sel_974330 = array_index_974017 == array_index_948955 ? add_974329 : sel_974326;
  assign add_974333 = sel_974330 + 8'h01;
  assign sel_974334 = array_index_974017 == array_index_948961 ? add_974333 : sel_974330;
  assign add_974337 = sel_974334 + 8'h01;
  assign sel_974338 = array_index_974017 == array_index_948967 ? add_974337 : sel_974334;
  assign add_974341 = sel_974338 + 8'h01;
  assign sel_974342 = array_index_974017 == array_index_948973 ? add_974341 : sel_974338;
  assign add_974345 = sel_974342 + 8'h01;
  assign sel_974346 = array_index_974017 == array_index_948979 ? add_974345 : sel_974342;
  assign add_974349 = sel_974346 + 8'h01;
  assign sel_974350 = array_index_974017 == array_index_948985 ? add_974349 : sel_974346;
  assign add_974353 = sel_974350 + 8'h01;
  assign sel_974354 = array_index_974017 == array_index_948991 ? add_974353 : sel_974350;
  assign add_974357 = sel_974354 + 8'h01;
  assign sel_974358 = array_index_974017 == array_index_948997 ? add_974357 : sel_974354;
  assign add_974361 = sel_974358 + 8'h01;
  assign sel_974362 = array_index_974017 == array_index_949003 ? add_974361 : sel_974358;
  assign add_974365 = sel_974362 + 8'h01;
  assign sel_974366 = array_index_974017 == array_index_949009 ? add_974365 : sel_974362;
  assign add_974369 = sel_974366 + 8'h01;
  assign sel_974370 = array_index_974017 == array_index_949015 ? add_974369 : sel_974366;
  assign add_974373 = sel_974370 + 8'h01;
  assign sel_974374 = array_index_974017 == array_index_949021 ? add_974373 : sel_974370;
  assign add_974377 = sel_974374 + 8'h01;
  assign sel_974378 = array_index_974017 == array_index_949027 ? add_974377 : sel_974374;
  assign add_974381 = sel_974378 + 8'h01;
  assign sel_974382 = array_index_974017 == array_index_949033 ? add_974381 : sel_974378;
  assign add_974385 = sel_974382 + 8'h01;
  assign sel_974386 = array_index_974017 == array_index_949039 ? add_974385 : sel_974382;
  assign add_974389 = sel_974386 + 8'h01;
  assign sel_974390 = array_index_974017 == array_index_949045 ? add_974389 : sel_974386;
  assign add_974393 = sel_974390 + 8'h01;
  assign sel_974394 = array_index_974017 == array_index_949051 ? add_974393 : sel_974390;
  assign add_974397 = sel_974394 + 8'h01;
  assign sel_974398 = array_index_974017 == array_index_949057 ? add_974397 : sel_974394;
  assign add_974401 = sel_974398 + 8'h01;
  assign sel_974402 = array_index_974017 == array_index_949063 ? add_974401 : sel_974398;
  assign add_974405 = sel_974402 + 8'h01;
  assign sel_974406 = array_index_974017 == array_index_949069 ? add_974405 : sel_974402;
  assign add_974409 = sel_974406 + 8'h01;
  assign sel_974410 = array_index_974017 == array_index_949075 ? add_974409 : sel_974406;
  assign add_974413 = sel_974410 + 8'h01;
  assign sel_974414 = array_index_974017 == array_index_949081 ? add_974413 : sel_974410;
  assign add_974418 = sel_974414 + 8'h01;
  assign array_index_974419 = set1_unflattened[7'h40];
  assign sel_974420 = array_index_974017 == array_index_949087 ? add_974418 : sel_974414;
  assign add_974423 = sel_974420 + 8'h01;
  assign sel_974424 = array_index_974419 == array_index_948483 ? add_974423 : sel_974420;
  assign add_974427 = sel_974424 + 8'h01;
  assign sel_974428 = array_index_974419 == array_index_948487 ? add_974427 : sel_974424;
  assign add_974431 = sel_974428 + 8'h01;
  assign sel_974432 = array_index_974419 == array_index_948495 ? add_974431 : sel_974428;
  assign add_974435 = sel_974432 + 8'h01;
  assign sel_974436 = array_index_974419 == array_index_948503 ? add_974435 : sel_974432;
  assign add_974439 = sel_974436 + 8'h01;
  assign sel_974440 = array_index_974419 == array_index_948511 ? add_974439 : sel_974436;
  assign add_974443 = sel_974440 + 8'h01;
  assign sel_974444 = array_index_974419 == array_index_948519 ? add_974443 : sel_974440;
  assign add_974447 = sel_974444 + 8'h01;
  assign sel_974448 = array_index_974419 == array_index_948527 ? add_974447 : sel_974444;
  assign add_974451 = sel_974448 + 8'h01;
  assign sel_974452 = array_index_974419 == array_index_948535 ? add_974451 : sel_974448;
  assign add_974455 = sel_974452 + 8'h01;
  assign sel_974456 = array_index_974419 == array_index_948541 ? add_974455 : sel_974452;
  assign add_974459 = sel_974456 + 8'h01;
  assign sel_974460 = array_index_974419 == array_index_948547 ? add_974459 : sel_974456;
  assign add_974463 = sel_974460 + 8'h01;
  assign sel_974464 = array_index_974419 == array_index_948553 ? add_974463 : sel_974460;
  assign add_974467 = sel_974464 + 8'h01;
  assign sel_974468 = array_index_974419 == array_index_948559 ? add_974467 : sel_974464;
  assign add_974471 = sel_974468 + 8'h01;
  assign sel_974472 = array_index_974419 == array_index_948565 ? add_974471 : sel_974468;
  assign add_974475 = sel_974472 + 8'h01;
  assign sel_974476 = array_index_974419 == array_index_948571 ? add_974475 : sel_974472;
  assign add_974479 = sel_974476 + 8'h01;
  assign sel_974480 = array_index_974419 == array_index_948577 ? add_974479 : sel_974476;
  assign add_974483 = sel_974480 + 8'h01;
  assign sel_974484 = array_index_974419 == array_index_948583 ? add_974483 : sel_974480;
  assign add_974487 = sel_974484 + 8'h01;
  assign sel_974488 = array_index_974419 == array_index_948589 ? add_974487 : sel_974484;
  assign add_974491 = sel_974488 + 8'h01;
  assign sel_974492 = array_index_974419 == array_index_948595 ? add_974491 : sel_974488;
  assign add_974495 = sel_974492 + 8'h01;
  assign sel_974496 = array_index_974419 == array_index_948601 ? add_974495 : sel_974492;
  assign add_974499 = sel_974496 + 8'h01;
  assign sel_974500 = array_index_974419 == array_index_948607 ? add_974499 : sel_974496;
  assign add_974503 = sel_974500 + 8'h01;
  assign sel_974504 = array_index_974419 == array_index_948613 ? add_974503 : sel_974500;
  assign add_974507 = sel_974504 + 8'h01;
  assign sel_974508 = array_index_974419 == array_index_948619 ? add_974507 : sel_974504;
  assign add_974511 = sel_974508 + 8'h01;
  assign sel_974512 = array_index_974419 == array_index_948625 ? add_974511 : sel_974508;
  assign add_974515 = sel_974512 + 8'h01;
  assign sel_974516 = array_index_974419 == array_index_948631 ? add_974515 : sel_974512;
  assign add_974519 = sel_974516 + 8'h01;
  assign sel_974520 = array_index_974419 == array_index_948637 ? add_974519 : sel_974516;
  assign add_974523 = sel_974520 + 8'h01;
  assign sel_974524 = array_index_974419 == array_index_948643 ? add_974523 : sel_974520;
  assign add_974527 = sel_974524 + 8'h01;
  assign sel_974528 = array_index_974419 == array_index_948649 ? add_974527 : sel_974524;
  assign add_974531 = sel_974528 + 8'h01;
  assign sel_974532 = array_index_974419 == array_index_948655 ? add_974531 : sel_974528;
  assign add_974535 = sel_974532 + 8'h01;
  assign sel_974536 = array_index_974419 == array_index_948661 ? add_974535 : sel_974532;
  assign add_974539 = sel_974536 + 8'h01;
  assign sel_974540 = array_index_974419 == array_index_948667 ? add_974539 : sel_974536;
  assign add_974543 = sel_974540 + 8'h01;
  assign sel_974544 = array_index_974419 == array_index_948673 ? add_974543 : sel_974540;
  assign add_974547 = sel_974544 + 8'h01;
  assign sel_974548 = array_index_974419 == array_index_948679 ? add_974547 : sel_974544;
  assign add_974551 = sel_974548 + 8'h01;
  assign sel_974552 = array_index_974419 == array_index_948685 ? add_974551 : sel_974548;
  assign add_974555 = sel_974552 + 8'h01;
  assign sel_974556 = array_index_974419 == array_index_948691 ? add_974555 : sel_974552;
  assign add_974559 = sel_974556 + 8'h01;
  assign sel_974560 = array_index_974419 == array_index_948697 ? add_974559 : sel_974556;
  assign add_974563 = sel_974560 + 8'h01;
  assign sel_974564 = array_index_974419 == array_index_948703 ? add_974563 : sel_974560;
  assign add_974567 = sel_974564 + 8'h01;
  assign sel_974568 = array_index_974419 == array_index_948709 ? add_974567 : sel_974564;
  assign add_974571 = sel_974568 + 8'h01;
  assign sel_974572 = array_index_974419 == array_index_948715 ? add_974571 : sel_974568;
  assign add_974575 = sel_974572 + 8'h01;
  assign sel_974576 = array_index_974419 == array_index_948721 ? add_974575 : sel_974572;
  assign add_974579 = sel_974576 + 8'h01;
  assign sel_974580 = array_index_974419 == array_index_948727 ? add_974579 : sel_974576;
  assign add_974583 = sel_974580 + 8'h01;
  assign sel_974584 = array_index_974419 == array_index_948733 ? add_974583 : sel_974580;
  assign add_974587 = sel_974584 + 8'h01;
  assign sel_974588 = array_index_974419 == array_index_948739 ? add_974587 : sel_974584;
  assign add_974591 = sel_974588 + 8'h01;
  assign sel_974592 = array_index_974419 == array_index_948745 ? add_974591 : sel_974588;
  assign add_974595 = sel_974592 + 8'h01;
  assign sel_974596 = array_index_974419 == array_index_948751 ? add_974595 : sel_974592;
  assign add_974599 = sel_974596 + 8'h01;
  assign sel_974600 = array_index_974419 == array_index_948757 ? add_974599 : sel_974596;
  assign add_974603 = sel_974600 + 8'h01;
  assign sel_974604 = array_index_974419 == array_index_948763 ? add_974603 : sel_974600;
  assign add_974607 = sel_974604 + 8'h01;
  assign sel_974608 = array_index_974419 == array_index_948769 ? add_974607 : sel_974604;
  assign add_974611 = sel_974608 + 8'h01;
  assign sel_974612 = array_index_974419 == array_index_948775 ? add_974611 : sel_974608;
  assign add_974615 = sel_974612 + 8'h01;
  assign sel_974616 = array_index_974419 == array_index_948781 ? add_974615 : sel_974612;
  assign add_974619 = sel_974616 + 8'h01;
  assign sel_974620 = array_index_974419 == array_index_948787 ? add_974619 : sel_974616;
  assign add_974623 = sel_974620 + 8'h01;
  assign sel_974624 = array_index_974419 == array_index_948793 ? add_974623 : sel_974620;
  assign add_974627 = sel_974624 + 8'h01;
  assign sel_974628 = array_index_974419 == array_index_948799 ? add_974627 : sel_974624;
  assign add_974631 = sel_974628 + 8'h01;
  assign sel_974632 = array_index_974419 == array_index_948805 ? add_974631 : sel_974628;
  assign add_974635 = sel_974632 + 8'h01;
  assign sel_974636 = array_index_974419 == array_index_948811 ? add_974635 : sel_974632;
  assign add_974639 = sel_974636 + 8'h01;
  assign sel_974640 = array_index_974419 == array_index_948817 ? add_974639 : sel_974636;
  assign add_974643 = sel_974640 + 8'h01;
  assign sel_974644 = array_index_974419 == array_index_948823 ? add_974643 : sel_974640;
  assign add_974647 = sel_974644 + 8'h01;
  assign sel_974648 = array_index_974419 == array_index_948829 ? add_974647 : sel_974644;
  assign add_974651 = sel_974648 + 8'h01;
  assign sel_974652 = array_index_974419 == array_index_948835 ? add_974651 : sel_974648;
  assign add_974655 = sel_974652 + 8'h01;
  assign sel_974656 = array_index_974419 == array_index_948841 ? add_974655 : sel_974652;
  assign add_974659 = sel_974656 + 8'h01;
  assign sel_974660 = array_index_974419 == array_index_948847 ? add_974659 : sel_974656;
  assign add_974663 = sel_974660 + 8'h01;
  assign sel_974664 = array_index_974419 == array_index_948853 ? add_974663 : sel_974660;
  assign add_974667 = sel_974664 + 8'h01;
  assign sel_974668 = array_index_974419 == array_index_948859 ? add_974667 : sel_974664;
  assign add_974671 = sel_974668 + 8'h01;
  assign sel_974672 = array_index_974419 == array_index_948865 ? add_974671 : sel_974668;
  assign add_974675 = sel_974672 + 8'h01;
  assign sel_974676 = array_index_974419 == array_index_948871 ? add_974675 : sel_974672;
  assign add_974679 = sel_974676 + 8'h01;
  assign sel_974680 = array_index_974419 == array_index_948877 ? add_974679 : sel_974676;
  assign add_974683 = sel_974680 + 8'h01;
  assign sel_974684 = array_index_974419 == array_index_948883 ? add_974683 : sel_974680;
  assign add_974687 = sel_974684 + 8'h01;
  assign sel_974688 = array_index_974419 == array_index_948889 ? add_974687 : sel_974684;
  assign add_974691 = sel_974688 + 8'h01;
  assign sel_974692 = array_index_974419 == array_index_948895 ? add_974691 : sel_974688;
  assign add_974695 = sel_974692 + 8'h01;
  assign sel_974696 = array_index_974419 == array_index_948901 ? add_974695 : sel_974692;
  assign add_974699 = sel_974696 + 8'h01;
  assign sel_974700 = array_index_974419 == array_index_948907 ? add_974699 : sel_974696;
  assign add_974703 = sel_974700 + 8'h01;
  assign sel_974704 = array_index_974419 == array_index_948913 ? add_974703 : sel_974700;
  assign add_974707 = sel_974704 + 8'h01;
  assign sel_974708 = array_index_974419 == array_index_948919 ? add_974707 : sel_974704;
  assign add_974711 = sel_974708 + 8'h01;
  assign sel_974712 = array_index_974419 == array_index_948925 ? add_974711 : sel_974708;
  assign add_974715 = sel_974712 + 8'h01;
  assign sel_974716 = array_index_974419 == array_index_948931 ? add_974715 : sel_974712;
  assign add_974719 = sel_974716 + 8'h01;
  assign sel_974720 = array_index_974419 == array_index_948937 ? add_974719 : sel_974716;
  assign add_974723 = sel_974720 + 8'h01;
  assign sel_974724 = array_index_974419 == array_index_948943 ? add_974723 : sel_974720;
  assign add_974727 = sel_974724 + 8'h01;
  assign sel_974728 = array_index_974419 == array_index_948949 ? add_974727 : sel_974724;
  assign add_974731 = sel_974728 + 8'h01;
  assign sel_974732 = array_index_974419 == array_index_948955 ? add_974731 : sel_974728;
  assign add_974735 = sel_974732 + 8'h01;
  assign sel_974736 = array_index_974419 == array_index_948961 ? add_974735 : sel_974732;
  assign add_974739 = sel_974736 + 8'h01;
  assign sel_974740 = array_index_974419 == array_index_948967 ? add_974739 : sel_974736;
  assign add_974743 = sel_974740 + 8'h01;
  assign sel_974744 = array_index_974419 == array_index_948973 ? add_974743 : sel_974740;
  assign add_974747 = sel_974744 + 8'h01;
  assign sel_974748 = array_index_974419 == array_index_948979 ? add_974747 : sel_974744;
  assign add_974751 = sel_974748 + 8'h01;
  assign sel_974752 = array_index_974419 == array_index_948985 ? add_974751 : sel_974748;
  assign add_974755 = sel_974752 + 8'h01;
  assign sel_974756 = array_index_974419 == array_index_948991 ? add_974755 : sel_974752;
  assign add_974759 = sel_974756 + 8'h01;
  assign sel_974760 = array_index_974419 == array_index_948997 ? add_974759 : sel_974756;
  assign add_974763 = sel_974760 + 8'h01;
  assign sel_974764 = array_index_974419 == array_index_949003 ? add_974763 : sel_974760;
  assign add_974767 = sel_974764 + 8'h01;
  assign sel_974768 = array_index_974419 == array_index_949009 ? add_974767 : sel_974764;
  assign add_974771 = sel_974768 + 8'h01;
  assign sel_974772 = array_index_974419 == array_index_949015 ? add_974771 : sel_974768;
  assign add_974775 = sel_974772 + 8'h01;
  assign sel_974776 = array_index_974419 == array_index_949021 ? add_974775 : sel_974772;
  assign add_974779 = sel_974776 + 8'h01;
  assign sel_974780 = array_index_974419 == array_index_949027 ? add_974779 : sel_974776;
  assign add_974783 = sel_974780 + 8'h01;
  assign sel_974784 = array_index_974419 == array_index_949033 ? add_974783 : sel_974780;
  assign add_974787 = sel_974784 + 8'h01;
  assign sel_974788 = array_index_974419 == array_index_949039 ? add_974787 : sel_974784;
  assign add_974791 = sel_974788 + 8'h01;
  assign sel_974792 = array_index_974419 == array_index_949045 ? add_974791 : sel_974788;
  assign add_974795 = sel_974792 + 8'h01;
  assign sel_974796 = array_index_974419 == array_index_949051 ? add_974795 : sel_974792;
  assign add_974799 = sel_974796 + 8'h01;
  assign sel_974800 = array_index_974419 == array_index_949057 ? add_974799 : sel_974796;
  assign add_974803 = sel_974800 + 8'h01;
  assign sel_974804 = array_index_974419 == array_index_949063 ? add_974803 : sel_974800;
  assign add_974807 = sel_974804 + 8'h01;
  assign sel_974808 = array_index_974419 == array_index_949069 ? add_974807 : sel_974804;
  assign add_974811 = sel_974808 + 8'h01;
  assign sel_974812 = array_index_974419 == array_index_949075 ? add_974811 : sel_974808;
  assign add_974815 = sel_974812 + 8'h01;
  assign sel_974816 = array_index_974419 == array_index_949081 ? add_974815 : sel_974812;
  assign add_974820 = sel_974816 + 8'h01;
  assign array_index_974821 = set1_unflattened[7'h41];
  assign sel_974822 = array_index_974419 == array_index_949087 ? add_974820 : sel_974816;
  assign add_974825 = sel_974822 + 8'h01;
  assign sel_974826 = array_index_974821 == array_index_948483 ? add_974825 : sel_974822;
  assign add_974829 = sel_974826 + 8'h01;
  assign sel_974830 = array_index_974821 == array_index_948487 ? add_974829 : sel_974826;
  assign add_974833 = sel_974830 + 8'h01;
  assign sel_974834 = array_index_974821 == array_index_948495 ? add_974833 : sel_974830;
  assign add_974837 = sel_974834 + 8'h01;
  assign sel_974838 = array_index_974821 == array_index_948503 ? add_974837 : sel_974834;
  assign add_974841 = sel_974838 + 8'h01;
  assign sel_974842 = array_index_974821 == array_index_948511 ? add_974841 : sel_974838;
  assign add_974845 = sel_974842 + 8'h01;
  assign sel_974846 = array_index_974821 == array_index_948519 ? add_974845 : sel_974842;
  assign add_974849 = sel_974846 + 8'h01;
  assign sel_974850 = array_index_974821 == array_index_948527 ? add_974849 : sel_974846;
  assign add_974853 = sel_974850 + 8'h01;
  assign sel_974854 = array_index_974821 == array_index_948535 ? add_974853 : sel_974850;
  assign add_974857 = sel_974854 + 8'h01;
  assign sel_974858 = array_index_974821 == array_index_948541 ? add_974857 : sel_974854;
  assign add_974861 = sel_974858 + 8'h01;
  assign sel_974862 = array_index_974821 == array_index_948547 ? add_974861 : sel_974858;
  assign add_974865 = sel_974862 + 8'h01;
  assign sel_974866 = array_index_974821 == array_index_948553 ? add_974865 : sel_974862;
  assign add_974869 = sel_974866 + 8'h01;
  assign sel_974870 = array_index_974821 == array_index_948559 ? add_974869 : sel_974866;
  assign add_974873 = sel_974870 + 8'h01;
  assign sel_974874 = array_index_974821 == array_index_948565 ? add_974873 : sel_974870;
  assign add_974877 = sel_974874 + 8'h01;
  assign sel_974878 = array_index_974821 == array_index_948571 ? add_974877 : sel_974874;
  assign add_974881 = sel_974878 + 8'h01;
  assign sel_974882 = array_index_974821 == array_index_948577 ? add_974881 : sel_974878;
  assign add_974885 = sel_974882 + 8'h01;
  assign sel_974886 = array_index_974821 == array_index_948583 ? add_974885 : sel_974882;
  assign add_974889 = sel_974886 + 8'h01;
  assign sel_974890 = array_index_974821 == array_index_948589 ? add_974889 : sel_974886;
  assign add_974893 = sel_974890 + 8'h01;
  assign sel_974894 = array_index_974821 == array_index_948595 ? add_974893 : sel_974890;
  assign add_974897 = sel_974894 + 8'h01;
  assign sel_974898 = array_index_974821 == array_index_948601 ? add_974897 : sel_974894;
  assign add_974901 = sel_974898 + 8'h01;
  assign sel_974902 = array_index_974821 == array_index_948607 ? add_974901 : sel_974898;
  assign add_974905 = sel_974902 + 8'h01;
  assign sel_974906 = array_index_974821 == array_index_948613 ? add_974905 : sel_974902;
  assign add_974909 = sel_974906 + 8'h01;
  assign sel_974910 = array_index_974821 == array_index_948619 ? add_974909 : sel_974906;
  assign add_974913 = sel_974910 + 8'h01;
  assign sel_974914 = array_index_974821 == array_index_948625 ? add_974913 : sel_974910;
  assign add_974917 = sel_974914 + 8'h01;
  assign sel_974918 = array_index_974821 == array_index_948631 ? add_974917 : sel_974914;
  assign add_974921 = sel_974918 + 8'h01;
  assign sel_974922 = array_index_974821 == array_index_948637 ? add_974921 : sel_974918;
  assign add_974925 = sel_974922 + 8'h01;
  assign sel_974926 = array_index_974821 == array_index_948643 ? add_974925 : sel_974922;
  assign add_974929 = sel_974926 + 8'h01;
  assign sel_974930 = array_index_974821 == array_index_948649 ? add_974929 : sel_974926;
  assign add_974933 = sel_974930 + 8'h01;
  assign sel_974934 = array_index_974821 == array_index_948655 ? add_974933 : sel_974930;
  assign add_974937 = sel_974934 + 8'h01;
  assign sel_974938 = array_index_974821 == array_index_948661 ? add_974937 : sel_974934;
  assign add_974941 = sel_974938 + 8'h01;
  assign sel_974942 = array_index_974821 == array_index_948667 ? add_974941 : sel_974938;
  assign add_974945 = sel_974942 + 8'h01;
  assign sel_974946 = array_index_974821 == array_index_948673 ? add_974945 : sel_974942;
  assign add_974949 = sel_974946 + 8'h01;
  assign sel_974950 = array_index_974821 == array_index_948679 ? add_974949 : sel_974946;
  assign add_974953 = sel_974950 + 8'h01;
  assign sel_974954 = array_index_974821 == array_index_948685 ? add_974953 : sel_974950;
  assign add_974957 = sel_974954 + 8'h01;
  assign sel_974958 = array_index_974821 == array_index_948691 ? add_974957 : sel_974954;
  assign add_974961 = sel_974958 + 8'h01;
  assign sel_974962 = array_index_974821 == array_index_948697 ? add_974961 : sel_974958;
  assign add_974965 = sel_974962 + 8'h01;
  assign sel_974966 = array_index_974821 == array_index_948703 ? add_974965 : sel_974962;
  assign add_974969 = sel_974966 + 8'h01;
  assign sel_974970 = array_index_974821 == array_index_948709 ? add_974969 : sel_974966;
  assign add_974973 = sel_974970 + 8'h01;
  assign sel_974974 = array_index_974821 == array_index_948715 ? add_974973 : sel_974970;
  assign add_974977 = sel_974974 + 8'h01;
  assign sel_974978 = array_index_974821 == array_index_948721 ? add_974977 : sel_974974;
  assign add_974981 = sel_974978 + 8'h01;
  assign sel_974982 = array_index_974821 == array_index_948727 ? add_974981 : sel_974978;
  assign add_974985 = sel_974982 + 8'h01;
  assign sel_974986 = array_index_974821 == array_index_948733 ? add_974985 : sel_974982;
  assign add_974989 = sel_974986 + 8'h01;
  assign sel_974990 = array_index_974821 == array_index_948739 ? add_974989 : sel_974986;
  assign add_974993 = sel_974990 + 8'h01;
  assign sel_974994 = array_index_974821 == array_index_948745 ? add_974993 : sel_974990;
  assign add_974997 = sel_974994 + 8'h01;
  assign sel_974998 = array_index_974821 == array_index_948751 ? add_974997 : sel_974994;
  assign add_975001 = sel_974998 + 8'h01;
  assign sel_975002 = array_index_974821 == array_index_948757 ? add_975001 : sel_974998;
  assign add_975005 = sel_975002 + 8'h01;
  assign sel_975006 = array_index_974821 == array_index_948763 ? add_975005 : sel_975002;
  assign add_975009 = sel_975006 + 8'h01;
  assign sel_975010 = array_index_974821 == array_index_948769 ? add_975009 : sel_975006;
  assign add_975013 = sel_975010 + 8'h01;
  assign sel_975014 = array_index_974821 == array_index_948775 ? add_975013 : sel_975010;
  assign add_975017 = sel_975014 + 8'h01;
  assign sel_975018 = array_index_974821 == array_index_948781 ? add_975017 : sel_975014;
  assign add_975021 = sel_975018 + 8'h01;
  assign sel_975022 = array_index_974821 == array_index_948787 ? add_975021 : sel_975018;
  assign add_975025 = sel_975022 + 8'h01;
  assign sel_975026 = array_index_974821 == array_index_948793 ? add_975025 : sel_975022;
  assign add_975029 = sel_975026 + 8'h01;
  assign sel_975030 = array_index_974821 == array_index_948799 ? add_975029 : sel_975026;
  assign add_975033 = sel_975030 + 8'h01;
  assign sel_975034 = array_index_974821 == array_index_948805 ? add_975033 : sel_975030;
  assign add_975037 = sel_975034 + 8'h01;
  assign sel_975038 = array_index_974821 == array_index_948811 ? add_975037 : sel_975034;
  assign add_975041 = sel_975038 + 8'h01;
  assign sel_975042 = array_index_974821 == array_index_948817 ? add_975041 : sel_975038;
  assign add_975045 = sel_975042 + 8'h01;
  assign sel_975046 = array_index_974821 == array_index_948823 ? add_975045 : sel_975042;
  assign add_975049 = sel_975046 + 8'h01;
  assign sel_975050 = array_index_974821 == array_index_948829 ? add_975049 : sel_975046;
  assign add_975053 = sel_975050 + 8'h01;
  assign sel_975054 = array_index_974821 == array_index_948835 ? add_975053 : sel_975050;
  assign add_975057 = sel_975054 + 8'h01;
  assign sel_975058 = array_index_974821 == array_index_948841 ? add_975057 : sel_975054;
  assign add_975061 = sel_975058 + 8'h01;
  assign sel_975062 = array_index_974821 == array_index_948847 ? add_975061 : sel_975058;
  assign add_975065 = sel_975062 + 8'h01;
  assign sel_975066 = array_index_974821 == array_index_948853 ? add_975065 : sel_975062;
  assign add_975069 = sel_975066 + 8'h01;
  assign sel_975070 = array_index_974821 == array_index_948859 ? add_975069 : sel_975066;
  assign add_975073 = sel_975070 + 8'h01;
  assign sel_975074 = array_index_974821 == array_index_948865 ? add_975073 : sel_975070;
  assign add_975077 = sel_975074 + 8'h01;
  assign sel_975078 = array_index_974821 == array_index_948871 ? add_975077 : sel_975074;
  assign add_975081 = sel_975078 + 8'h01;
  assign sel_975082 = array_index_974821 == array_index_948877 ? add_975081 : sel_975078;
  assign add_975085 = sel_975082 + 8'h01;
  assign sel_975086 = array_index_974821 == array_index_948883 ? add_975085 : sel_975082;
  assign add_975089 = sel_975086 + 8'h01;
  assign sel_975090 = array_index_974821 == array_index_948889 ? add_975089 : sel_975086;
  assign add_975093 = sel_975090 + 8'h01;
  assign sel_975094 = array_index_974821 == array_index_948895 ? add_975093 : sel_975090;
  assign add_975097 = sel_975094 + 8'h01;
  assign sel_975098 = array_index_974821 == array_index_948901 ? add_975097 : sel_975094;
  assign add_975101 = sel_975098 + 8'h01;
  assign sel_975102 = array_index_974821 == array_index_948907 ? add_975101 : sel_975098;
  assign add_975105 = sel_975102 + 8'h01;
  assign sel_975106 = array_index_974821 == array_index_948913 ? add_975105 : sel_975102;
  assign add_975109 = sel_975106 + 8'h01;
  assign sel_975110 = array_index_974821 == array_index_948919 ? add_975109 : sel_975106;
  assign add_975113 = sel_975110 + 8'h01;
  assign sel_975114 = array_index_974821 == array_index_948925 ? add_975113 : sel_975110;
  assign add_975117 = sel_975114 + 8'h01;
  assign sel_975118 = array_index_974821 == array_index_948931 ? add_975117 : sel_975114;
  assign add_975121 = sel_975118 + 8'h01;
  assign sel_975122 = array_index_974821 == array_index_948937 ? add_975121 : sel_975118;
  assign add_975125 = sel_975122 + 8'h01;
  assign sel_975126 = array_index_974821 == array_index_948943 ? add_975125 : sel_975122;
  assign add_975129 = sel_975126 + 8'h01;
  assign sel_975130 = array_index_974821 == array_index_948949 ? add_975129 : sel_975126;
  assign add_975133 = sel_975130 + 8'h01;
  assign sel_975134 = array_index_974821 == array_index_948955 ? add_975133 : sel_975130;
  assign add_975137 = sel_975134 + 8'h01;
  assign sel_975138 = array_index_974821 == array_index_948961 ? add_975137 : sel_975134;
  assign add_975141 = sel_975138 + 8'h01;
  assign sel_975142 = array_index_974821 == array_index_948967 ? add_975141 : sel_975138;
  assign add_975145 = sel_975142 + 8'h01;
  assign sel_975146 = array_index_974821 == array_index_948973 ? add_975145 : sel_975142;
  assign add_975149 = sel_975146 + 8'h01;
  assign sel_975150 = array_index_974821 == array_index_948979 ? add_975149 : sel_975146;
  assign add_975153 = sel_975150 + 8'h01;
  assign sel_975154 = array_index_974821 == array_index_948985 ? add_975153 : sel_975150;
  assign add_975157 = sel_975154 + 8'h01;
  assign sel_975158 = array_index_974821 == array_index_948991 ? add_975157 : sel_975154;
  assign add_975161 = sel_975158 + 8'h01;
  assign sel_975162 = array_index_974821 == array_index_948997 ? add_975161 : sel_975158;
  assign add_975165 = sel_975162 + 8'h01;
  assign sel_975166 = array_index_974821 == array_index_949003 ? add_975165 : sel_975162;
  assign add_975169 = sel_975166 + 8'h01;
  assign sel_975170 = array_index_974821 == array_index_949009 ? add_975169 : sel_975166;
  assign add_975173 = sel_975170 + 8'h01;
  assign sel_975174 = array_index_974821 == array_index_949015 ? add_975173 : sel_975170;
  assign add_975177 = sel_975174 + 8'h01;
  assign sel_975178 = array_index_974821 == array_index_949021 ? add_975177 : sel_975174;
  assign add_975181 = sel_975178 + 8'h01;
  assign sel_975182 = array_index_974821 == array_index_949027 ? add_975181 : sel_975178;
  assign add_975185 = sel_975182 + 8'h01;
  assign sel_975186 = array_index_974821 == array_index_949033 ? add_975185 : sel_975182;
  assign add_975189 = sel_975186 + 8'h01;
  assign sel_975190 = array_index_974821 == array_index_949039 ? add_975189 : sel_975186;
  assign add_975193 = sel_975190 + 8'h01;
  assign sel_975194 = array_index_974821 == array_index_949045 ? add_975193 : sel_975190;
  assign add_975197 = sel_975194 + 8'h01;
  assign sel_975198 = array_index_974821 == array_index_949051 ? add_975197 : sel_975194;
  assign add_975201 = sel_975198 + 8'h01;
  assign sel_975202 = array_index_974821 == array_index_949057 ? add_975201 : sel_975198;
  assign add_975205 = sel_975202 + 8'h01;
  assign sel_975206 = array_index_974821 == array_index_949063 ? add_975205 : sel_975202;
  assign add_975209 = sel_975206 + 8'h01;
  assign sel_975210 = array_index_974821 == array_index_949069 ? add_975209 : sel_975206;
  assign add_975213 = sel_975210 + 8'h01;
  assign sel_975214 = array_index_974821 == array_index_949075 ? add_975213 : sel_975210;
  assign add_975217 = sel_975214 + 8'h01;
  assign sel_975218 = array_index_974821 == array_index_949081 ? add_975217 : sel_975214;
  assign add_975222 = sel_975218 + 8'h01;
  assign array_index_975223 = set1_unflattened[7'h42];
  assign sel_975224 = array_index_974821 == array_index_949087 ? add_975222 : sel_975218;
  assign add_975227 = sel_975224 + 8'h01;
  assign sel_975228 = array_index_975223 == array_index_948483 ? add_975227 : sel_975224;
  assign add_975231 = sel_975228 + 8'h01;
  assign sel_975232 = array_index_975223 == array_index_948487 ? add_975231 : sel_975228;
  assign add_975235 = sel_975232 + 8'h01;
  assign sel_975236 = array_index_975223 == array_index_948495 ? add_975235 : sel_975232;
  assign add_975239 = sel_975236 + 8'h01;
  assign sel_975240 = array_index_975223 == array_index_948503 ? add_975239 : sel_975236;
  assign add_975243 = sel_975240 + 8'h01;
  assign sel_975244 = array_index_975223 == array_index_948511 ? add_975243 : sel_975240;
  assign add_975247 = sel_975244 + 8'h01;
  assign sel_975248 = array_index_975223 == array_index_948519 ? add_975247 : sel_975244;
  assign add_975251 = sel_975248 + 8'h01;
  assign sel_975252 = array_index_975223 == array_index_948527 ? add_975251 : sel_975248;
  assign add_975255 = sel_975252 + 8'h01;
  assign sel_975256 = array_index_975223 == array_index_948535 ? add_975255 : sel_975252;
  assign add_975259 = sel_975256 + 8'h01;
  assign sel_975260 = array_index_975223 == array_index_948541 ? add_975259 : sel_975256;
  assign add_975263 = sel_975260 + 8'h01;
  assign sel_975264 = array_index_975223 == array_index_948547 ? add_975263 : sel_975260;
  assign add_975267 = sel_975264 + 8'h01;
  assign sel_975268 = array_index_975223 == array_index_948553 ? add_975267 : sel_975264;
  assign add_975271 = sel_975268 + 8'h01;
  assign sel_975272 = array_index_975223 == array_index_948559 ? add_975271 : sel_975268;
  assign add_975275 = sel_975272 + 8'h01;
  assign sel_975276 = array_index_975223 == array_index_948565 ? add_975275 : sel_975272;
  assign add_975279 = sel_975276 + 8'h01;
  assign sel_975280 = array_index_975223 == array_index_948571 ? add_975279 : sel_975276;
  assign add_975283 = sel_975280 + 8'h01;
  assign sel_975284 = array_index_975223 == array_index_948577 ? add_975283 : sel_975280;
  assign add_975287 = sel_975284 + 8'h01;
  assign sel_975288 = array_index_975223 == array_index_948583 ? add_975287 : sel_975284;
  assign add_975291 = sel_975288 + 8'h01;
  assign sel_975292 = array_index_975223 == array_index_948589 ? add_975291 : sel_975288;
  assign add_975295 = sel_975292 + 8'h01;
  assign sel_975296 = array_index_975223 == array_index_948595 ? add_975295 : sel_975292;
  assign add_975299 = sel_975296 + 8'h01;
  assign sel_975300 = array_index_975223 == array_index_948601 ? add_975299 : sel_975296;
  assign add_975303 = sel_975300 + 8'h01;
  assign sel_975304 = array_index_975223 == array_index_948607 ? add_975303 : sel_975300;
  assign add_975307 = sel_975304 + 8'h01;
  assign sel_975308 = array_index_975223 == array_index_948613 ? add_975307 : sel_975304;
  assign add_975311 = sel_975308 + 8'h01;
  assign sel_975312 = array_index_975223 == array_index_948619 ? add_975311 : sel_975308;
  assign add_975315 = sel_975312 + 8'h01;
  assign sel_975316 = array_index_975223 == array_index_948625 ? add_975315 : sel_975312;
  assign add_975319 = sel_975316 + 8'h01;
  assign sel_975320 = array_index_975223 == array_index_948631 ? add_975319 : sel_975316;
  assign add_975323 = sel_975320 + 8'h01;
  assign sel_975324 = array_index_975223 == array_index_948637 ? add_975323 : sel_975320;
  assign add_975327 = sel_975324 + 8'h01;
  assign sel_975328 = array_index_975223 == array_index_948643 ? add_975327 : sel_975324;
  assign add_975331 = sel_975328 + 8'h01;
  assign sel_975332 = array_index_975223 == array_index_948649 ? add_975331 : sel_975328;
  assign add_975335 = sel_975332 + 8'h01;
  assign sel_975336 = array_index_975223 == array_index_948655 ? add_975335 : sel_975332;
  assign add_975339 = sel_975336 + 8'h01;
  assign sel_975340 = array_index_975223 == array_index_948661 ? add_975339 : sel_975336;
  assign add_975343 = sel_975340 + 8'h01;
  assign sel_975344 = array_index_975223 == array_index_948667 ? add_975343 : sel_975340;
  assign add_975347 = sel_975344 + 8'h01;
  assign sel_975348 = array_index_975223 == array_index_948673 ? add_975347 : sel_975344;
  assign add_975351 = sel_975348 + 8'h01;
  assign sel_975352 = array_index_975223 == array_index_948679 ? add_975351 : sel_975348;
  assign add_975355 = sel_975352 + 8'h01;
  assign sel_975356 = array_index_975223 == array_index_948685 ? add_975355 : sel_975352;
  assign add_975359 = sel_975356 + 8'h01;
  assign sel_975360 = array_index_975223 == array_index_948691 ? add_975359 : sel_975356;
  assign add_975363 = sel_975360 + 8'h01;
  assign sel_975364 = array_index_975223 == array_index_948697 ? add_975363 : sel_975360;
  assign add_975367 = sel_975364 + 8'h01;
  assign sel_975368 = array_index_975223 == array_index_948703 ? add_975367 : sel_975364;
  assign add_975371 = sel_975368 + 8'h01;
  assign sel_975372 = array_index_975223 == array_index_948709 ? add_975371 : sel_975368;
  assign add_975375 = sel_975372 + 8'h01;
  assign sel_975376 = array_index_975223 == array_index_948715 ? add_975375 : sel_975372;
  assign add_975379 = sel_975376 + 8'h01;
  assign sel_975380 = array_index_975223 == array_index_948721 ? add_975379 : sel_975376;
  assign add_975383 = sel_975380 + 8'h01;
  assign sel_975384 = array_index_975223 == array_index_948727 ? add_975383 : sel_975380;
  assign add_975387 = sel_975384 + 8'h01;
  assign sel_975388 = array_index_975223 == array_index_948733 ? add_975387 : sel_975384;
  assign add_975391 = sel_975388 + 8'h01;
  assign sel_975392 = array_index_975223 == array_index_948739 ? add_975391 : sel_975388;
  assign add_975395 = sel_975392 + 8'h01;
  assign sel_975396 = array_index_975223 == array_index_948745 ? add_975395 : sel_975392;
  assign add_975399 = sel_975396 + 8'h01;
  assign sel_975400 = array_index_975223 == array_index_948751 ? add_975399 : sel_975396;
  assign add_975403 = sel_975400 + 8'h01;
  assign sel_975404 = array_index_975223 == array_index_948757 ? add_975403 : sel_975400;
  assign add_975407 = sel_975404 + 8'h01;
  assign sel_975408 = array_index_975223 == array_index_948763 ? add_975407 : sel_975404;
  assign add_975411 = sel_975408 + 8'h01;
  assign sel_975412 = array_index_975223 == array_index_948769 ? add_975411 : sel_975408;
  assign add_975415 = sel_975412 + 8'h01;
  assign sel_975416 = array_index_975223 == array_index_948775 ? add_975415 : sel_975412;
  assign add_975419 = sel_975416 + 8'h01;
  assign sel_975420 = array_index_975223 == array_index_948781 ? add_975419 : sel_975416;
  assign add_975423 = sel_975420 + 8'h01;
  assign sel_975424 = array_index_975223 == array_index_948787 ? add_975423 : sel_975420;
  assign add_975427 = sel_975424 + 8'h01;
  assign sel_975428 = array_index_975223 == array_index_948793 ? add_975427 : sel_975424;
  assign add_975431 = sel_975428 + 8'h01;
  assign sel_975432 = array_index_975223 == array_index_948799 ? add_975431 : sel_975428;
  assign add_975435 = sel_975432 + 8'h01;
  assign sel_975436 = array_index_975223 == array_index_948805 ? add_975435 : sel_975432;
  assign add_975439 = sel_975436 + 8'h01;
  assign sel_975440 = array_index_975223 == array_index_948811 ? add_975439 : sel_975436;
  assign add_975443 = sel_975440 + 8'h01;
  assign sel_975444 = array_index_975223 == array_index_948817 ? add_975443 : sel_975440;
  assign add_975447 = sel_975444 + 8'h01;
  assign sel_975448 = array_index_975223 == array_index_948823 ? add_975447 : sel_975444;
  assign add_975451 = sel_975448 + 8'h01;
  assign sel_975452 = array_index_975223 == array_index_948829 ? add_975451 : sel_975448;
  assign add_975455 = sel_975452 + 8'h01;
  assign sel_975456 = array_index_975223 == array_index_948835 ? add_975455 : sel_975452;
  assign add_975459 = sel_975456 + 8'h01;
  assign sel_975460 = array_index_975223 == array_index_948841 ? add_975459 : sel_975456;
  assign add_975463 = sel_975460 + 8'h01;
  assign sel_975464 = array_index_975223 == array_index_948847 ? add_975463 : sel_975460;
  assign add_975467 = sel_975464 + 8'h01;
  assign sel_975468 = array_index_975223 == array_index_948853 ? add_975467 : sel_975464;
  assign add_975471 = sel_975468 + 8'h01;
  assign sel_975472 = array_index_975223 == array_index_948859 ? add_975471 : sel_975468;
  assign add_975475 = sel_975472 + 8'h01;
  assign sel_975476 = array_index_975223 == array_index_948865 ? add_975475 : sel_975472;
  assign add_975479 = sel_975476 + 8'h01;
  assign sel_975480 = array_index_975223 == array_index_948871 ? add_975479 : sel_975476;
  assign add_975483 = sel_975480 + 8'h01;
  assign sel_975484 = array_index_975223 == array_index_948877 ? add_975483 : sel_975480;
  assign add_975487 = sel_975484 + 8'h01;
  assign sel_975488 = array_index_975223 == array_index_948883 ? add_975487 : sel_975484;
  assign add_975491 = sel_975488 + 8'h01;
  assign sel_975492 = array_index_975223 == array_index_948889 ? add_975491 : sel_975488;
  assign add_975495 = sel_975492 + 8'h01;
  assign sel_975496 = array_index_975223 == array_index_948895 ? add_975495 : sel_975492;
  assign add_975499 = sel_975496 + 8'h01;
  assign sel_975500 = array_index_975223 == array_index_948901 ? add_975499 : sel_975496;
  assign add_975503 = sel_975500 + 8'h01;
  assign sel_975504 = array_index_975223 == array_index_948907 ? add_975503 : sel_975500;
  assign add_975507 = sel_975504 + 8'h01;
  assign sel_975508 = array_index_975223 == array_index_948913 ? add_975507 : sel_975504;
  assign add_975511 = sel_975508 + 8'h01;
  assign sel_975512 = array_index_975223 == array_index_948919 ? add_975511 : sel_975508;
  assign add_975515 = sel_975512 + 8'h01;
  assign sel_975516 = array_index_975223 == array_index_948925 ? add_975515 : sel_975512;
  assign add_975519 = sel_975516 + 8'h01;
  assign sel_975520 = array_index_975223 == array_index_948931 ? add_975519 : sel_975516;
  assign add_975523 = sel_975520 + 8'h01;
  assign sel_975524 = array_index_975223 == array_index_948937 ? add_975523 : sel_975520;
  assign add_975527 = sel_975524 + 8'h01;
  assign sel_975528 = array_index_975223 == array_index_948943 ? add_975527 : sel_975524;
  assign add_975531 = sel_975528 + 8'h01;
  assign sel_975532 = array_index_975223 == array_index_948949 ? add_975531 : sel_975528;
  assign add_975535 = sel_975532 + 8'h01;
  assign sel_975536 = array_index_975223 == array_index_948955 ? add_975535 : sel_975532;
  assign add_975539 = sel_975536 + 8'h01;
  assign sel_975540 = array_index_975223 == array_index_948961 ? add_975539 : sel_975536;
  assign add_975543 = sel_975540 + 8'h01;
  assign sel_975544 = array_index_975223 == array_index_948967 ? add_975543 : sel_975540;
  assign add_975547 = sel_975544 + 8'h01;
  assign sel_975548 = array_index_975223 == array_index_948973 ? add_975547 : sel_975544;
  assign add_975551 = sel_975548 + 8'h01;
  assign sel_975552 = array_index_975223 == array_index_948979 ? add_975551 : sel_975548;
  assign add_975555 = sel_975552 + 8'h01;
  assign sel_975556 = array_index_975223 == array_index_948985 ? add_975555 : sel_975552;
  assign add_975559 = sel_975556 + 8'h01;
  assign sel_975560 = array_index_975223 == array_index_948991 ? add_975559 : sel_975556;
  assign add_975563 = sel_975560 + 8'h01;
  assign sel_975564 = array_index_975223 == array_index_948997 ? add_975563 : sel_975560;
  assign add_975567 = sel_975564 + 8'h01;
  assign sel_975568 = array_index_975223 == array_index_949003 ? add_975567 : sel_975564;
  assign add_975571 = sel_975568 + 8'h01;
  assign sel_975572 = array_index_975223 == array_index_949009 ? add_975571 : sel_975568;
  assign add_975575 = sel_975572 + 8'h01;
  assign sel_975576 = array_index_975223 == array_index_949015 ? add_975575 : sel_975572;
  assign add_975579 = sel_975576 + 8'h01;
  assign sel_975580 = array_index_975223 == array_index_949021 ? add_975579 : sel_975576;
  assign add_975583 = sel_975580 + 8'h01;
  assign sel_975584 = array_index_975223 == array_index_949027 ? add_975583 : sel_975580;
  assign add_975587 = sel_975584 + 8'h01;
  assign sel_975588 = array_index_975223 == array_index_949033 ? add_975587 : sel_975584;
  assign add_975591 = sel_975588 + 8'h01;
  assign sel_975592 = array_index_975223 == array_index_949039 ? add_975591 : sel_975588;
  assign add_975595 = sel_975592 + 8'h01;
  assign sel_975596 = array_index_975223 == array_index_949045 ? add_975595 : sel_975592;
  assign add_975599 = sel_975596 + 8'h01;
  assign sel_975600 = array_index_975223 == array_index_949051 ? add_975599 : sel_975596;
  assign add_975603 = sel_975600 + 8'h01;
  assign sel_975604 = array_index_975223 == array_index_949057 ? add_975603 : sel_975600;
  assign add_975607 = sel_975604 + 8'h01;
  assign sel_975608 = array_index_975223 == array_index_949063 ? add_975607 : sel_975604;
  assign add_975611 = sel_975608 + 8'h01;
  assign sel_975612 = array_index_975223 == array_index_949069 ? add_975611 : sel_975608;
  assign add_975615 = sel_975612 + 8'h01;
  assign sel_975616 = array_index_975223 == array_index_949075 ? add_975615 : sel_975612;
  assign add_975619 = sel_975616 + 8'h01;
  assign sel_975620 = array_index_975223 == array_index_949081 ? add_975619 : sel_975616;
  assign add_975624 = sel_975620 + 8'h01;
  assign array_index_975625 = set1_unflattened[7'h43];
  assign sel_975626 = array_index_975223 == array_index_949087 ? add_975624 : sel_975620;
  assign add_975629 = sel_975626 + 8'h01;
  assign sel_975630 = array_index_975625 == array_index_948483 ? add_975629 : sel_975626;
  assign add_975633 = sel_975630 + 8'h01;
  assign sel_975634 = array_index_975625 == array_index_948487 ? add_975633 : sel_975630;
  assign add_975637 = sel_975634 + 8'h01;
  assign sel_975638 = array_index_975625 == array_index_948495 ? add_975637 : sel_975634;
  assign add_975641 = sel_975638 + 8'h01;
  assign sel_975642 = array_index_975625 == array_index_948503 ? add_975641 : sel_975638;
  assign add_975645 = sel_975642 + 8'h01;
  assign sel_975646 = array_index_975625 == array_index_948511 ? add_975645 : sel_975642;
  assign add_975649 = sel_975646 + 8'h01;
  assign sel_975650 = array_index_975625 == array_index_948519 ? add_975649 : sel_975646;
  assign add_975653 = sel_975650 + 8'h01;
  assign sel_975654 = array_index_975625 == array_index_948527 ? add_975653 : sel_975650;
  assign add_975657 = sel_975654 + 8'h01;
  assign sel_975658 = array_index_975625 == array_index_948535 ? add_975657 : sel_975654;
  assign add_975661 = sel_975658 + 8'h01;
  assign sel_975662 = array_index_975625 == array_index_948541 ? add_975661 : sel_975658;
  assign add_975665 = sel_975662 + 8'h01;
  assign sel_975666 = array_index_975625 == array_index_948547 ? add_975665 : sel_975662;
  assign add_975669 = sel_975666 + 8'h01;
  assign sel_975670 = array_index_975625 == array_index_948553 ? add_975669 : sel_975666;
  assign add_975673 = sel_975670 + 8'h01;
  assign sel_975674 = array_index_975625 == array_index_948559 ? add_975673 : sel_975670;
  assign add_975677 = sel_975674 + 8'h01;
  assign sel_975678 = array_index_975625 == array_index_948565 ? add_975677 : sel_975674;
  assign add_975681 = sel_975678 + 8'h01;
  assign sel_975682 = array_index_975625 == array_index_948571 ? add_975681 : sel_975678;
  assign add_975685 = sel_975682 + 8'h01;
  assign sel_975686 = array_index_975625 == array_index_948577 ? add_975685 : sel_975682;
  assign add_975689 = sel_975686 + 8'h01;
  assign sel_975690 = array_index_975625 == array_index_948583 ? add_975689 : sel_975686;
  assign add_975693 = sel_975690 + 8'h01;
  assign sel_975694 = array_index_975625 == array_index_948589 ? add_975693 : sel_975690;
  assign add_975697 = sel_975694 + 8'h01;
  assign sel_975698 = array_index_975625 == array_index_948595 ? add_975697 : sel_975694;
  assign add_975701 = sel_975698 + 8'h01;
  assign sel_975702 = array_index_975625 == array_index_948601 ? add_975701 : sel_975698;
  assign add_975705 = sel_975702 + 8'h01;
  assign sel_975706 = array_index_975625 == array_index_948607 ? add_975705 : sel_975702;
  assign add_975709 = sel_975706 + 8'h01;
  assign sel_975710 = array_index_975625 == array_index_948613 ? add_975709 : sel_975706;
  assign add_975713 = sel_975710 + 8'h01;
  assign sel_975714 = array_index_975625 == array_index_948619 ? add_975713 : sel_975710;
  assign add_975717 = sel_975714 + 8'h01;
  assign sel_975718 = array_index_975625 == array_index_948625 ? add_975717 : sel_975714;
  assign add_975721 = sel_975718 + 8'h01;
  assign sel_975722 = array_index_975625 == array_index_948631 ? add_975721 : sel_975718;
  assign add_975725 = sel_975722 + 8'h01;
  assign sel_975726 = array_index_975625 == array_index_948637 ? add_975725 : sel_975722;
  assign add_975729 = sel_975726 + 8'h01;
  assign sel_975730 = array_index_975625 == array_index_948643 ? add_975729 : sel_975726;
  assign add_975733 = sel_975730 + 8'h01;
  assign sel_975734 = array_index_975625 == array_index_948649 ? add_975733 : sel_975730;
  assign add_975737 = sel_975734 + 8'h01;
  assign sel_975738 = array_index_975625 == array_index_948655 ? add_975737 : sel_975734;
  assign add_975741 = sel_975738 + 8'h01;
  assign sel_975742 = array_index_975625 == array_index_948661 ? add_975741 : sel_975738;
  assign add_975745 = sel_975742 + 8'h01;
  assign sel_975746 = array_index_975625 == array_index_948667 ? add_975745 : sel_975742;
  assign add_975749 = sel_975746 + 8'h01;
  assign sel_975750 = array_index_975625 == array_index_948673 ? add_975749 : sel_975746;
  assign add_975753 = sel_975750 + 8'h01;
  assign sel_975754 = array_index_975625 == array_index_948679 ? add_975753 : sel_975750;
  assign add_975757 = sel_975754 + 8'h01;
  assign sel_975758 = array_index_975625 == array_index_948685 ? add_975757 : sel_975754;
  assign add_975761 = sel_975758 + 8'h01;
  assign sel_975762 = array_index_975625 == array_index_948691 ? add_975761 : sel_975758;
  assign add_975765 = sel_975762 + 8'h01;
  assign sel_975766 = array_index_975625 == array_index_948697 ? add_975765 : sel_975762;
  assign add_975769 = sel_975766 + 8'h01;
  assign sel_975770 = array_index_975625 == array_index_948703 ? add_975769 : sel_975766;
  assign add_975773 = sel_975770 + 8'h01;
  assign sel_975774 = array_index_975625 == array_index_948709 ? add_975773 : sel_975770;
  assign add_975777 = sel_975774 + 8'h01;
  assign sel_975778 = array_index_975625 == array_index_948715 ? add_975777 : sel_975774;
  assign add_975781 = sel_975778 + 8'h01;
  assign sel_975782 = array_index_975625 == array_index_948721 ? add_975781 : sel_975778;
  assign add_975785 = sel_975782 + 8'h01;
  assign sel_975786 = array_index_975625 == array_index_948727 ? add_975785 : sel_975782;
  assign add_975789 = sel_975786 + 8'h01;
  assign sel_975790 = array_index_975625 == array_index_948733 ? add_975789 : sel_975786;
  assign add_975793 = sel_975790 + 8'h01;
  assign sel_975794 = array_index_975625 == array_index_948739 ? add_975793 : sel_975790;
  assign add_975797 = sel_975794 + 8'h01;
  assign sel_975798 = array_index_975625 == array_index_948745 ? add_975797 : sel_975794;
  assign add_975801 = sel_975798 + 8'h01;
  assign sel_975802 = array_index_975625 == array_index_948751 ? add_975801 : sel_975798;
  assign add_975805 = sel_975802 + 8'h01;
  assign sel_975806 = array_index_975625 == array_index_948757 ? add_975805 : sel_975802;
  assign add_975809 = sel_975806 + 8'h01;
  assign sel_975810 = array_index_975625 == array_index_948763 ? add_975809 : sel_975806;
  assign add_975813 = sel_975810 + 8'h01;
  assign sel_975814 = array_index_975625 == array_index_948769 ? add_975813 : sel_975810;
  assign add_975817 = sel_975814 + 8'h01;
  assign sel_975818 = array_index_975625 == array_index_948775 ? add_975817 : sel_975814;
  assign add_975821 = sel_975818 + 8'h01;
  assign sel_975822 = array_index_975625 == array_index_948781 ? add_975821 : sel_975818;
  assign add_975825 = sel_975822 + 8'h01;
  assign sel_975826 = array_index_975625 == array_index_948787 ? add_975825 : sel_975822;
  assign add_975829 = sel_975826 + 8'h01;
  assign sel_975830 = array_index_975625 == array_index_948793 ? add_975829 : sel_975826;
  assign add_975833 = sel_975830 + 8'h01;
  assign sel_975834 = array_index_975625 == array_index_948799 ? add_975833 : sel_975830;
  assign add_975837 = sel_975834 + 8'h01;
  assign sel_975838 = array_index_975625 == array_index_948805 ? add_975837 : sel_975834;
  assign add_975841 = sel_975838 + 8'h01;
  assign sel_975842 = array_index_975625 == array_index_948811 ? add_975841 : sel_975838;
  assign add_975845 = sel_975842 + 8'h01;
  assign sel_975846 = array_index_975625 == array_index_948817 ? add_975845 : sel_975842;
  assign add_975849 = sel_975846 + 8'h01;
  assign sel_975850 = array_index_975625 == array_index_948823 ? add_975849 : sel_975846;
  assign add_975853 = sel_975850 + 8'h01;
  assign sel_975854 = array_index_975625 == array_index_948829 ? add_975853 : sel_975850;
  assign add_975857 = sel_975854 + 8'h01;
  assign sel_975858 = array_index_975625 == array_index_948835 ? add_975857 : sel_975854;
  assign add_975861 = sel_975858 + 8'h01;
  assign sel_975862 = array_index_975625 == array_index_948841 ? add_975861 : sel_975858;
  assign add_975865 = sel_975862 + 8'h01;
  assign sel_975866 = array_index_975625 == array_index_948847 ? add_975865 : sel_975862;
  assign add_975869 = sel_975866 + 8'h01;
  assign sel_975870 = array_index_975625 == array_index_948853 ? add_975869 : sel_975866;
  assign add_975873 = sel_975870 + 8'h01;
  assign sel_975874 = array_index_975625 == array_index_948859 ? add_975873 : sel_975870;
  assign add_975877 = sel_975874 + 8'h01;
  assign sel_975878 = array_index_975625 == array_index_948865 ? add_975877 : sel_975874;
  assign add_975881 = sel_975878 + 8'h01;
  assign sel_975882 = array_index_975625 == array_index_948871 ? add_975881 : sel_975878;
  assign add_975885 = sel_975882 + 8'h01;
  assign sel_975886 = array_index_975625 == array_index_948877 ? add_975885 : sel_975882;
  assign add_975889 = sel_975886 + 8'h01;
  assign sel_975890 = array_index_975625 == array_index_948883 ? add_975889 : sel_975886;
  assign add_975893 = sel_975890 + 8'h01;
  assign sel_975894 = array_index_975625 == array_index_948889 ? add_975893 : sel_975890;
  assign add_975897 = sel_975894 + 8'h01;
  assign sel_975898 = array_index_975625 == array_index_948895 ? add_975897 : sel_975894;
  assign add_975901 = sel_975898 + 8'h01;
  assign sel_975902 = array_index_975625 == array_index_948901 ? add_975901 : sel_975898;
  assign add_975905 = sel_975902 + 8'h01;
  assign sel_975906 = array_index_975625 == array_index_948907 ? add_975905 : sel_975902;
  assign add_975909 = sel_975906 + 8'h01;
  assign sel_975910 = array_index_975625 == array_index_948913 ? add_975909 : sel_975906;
  assign add_975913 = sel_975910 + 8'h01;
  assign sel_975914 = array_index_975625 == array_index_948919 ? add_975913 : sel_975910;
  assign add_975917 = sel_975914 + 8'h01;
  assign sel_975918 = array_index_975625 == array_index_948925 ? add_975917 : sel_975914;
  assign add_975921 = sel_975918 + 8'h01;
  assign sel_975922 = array_index_975625 == array_index_948931 ? add_975921 : sel_975918;
  assign add_975925 = sel_975922 + 8'h01;
  assign sel_975926 = array_index_975625 == array_index_948937 ? add_975925 : sel_975922;
  assign add_975929 = sel_975926 + 8'h01;
  assign sel_975930 = array_index_975625 == array_index_948943 ? add_975929 : sel_975926;
  assign add_975933 = sel_975930 + 8'h01;
  assign sel_975934 = array_index_975625 == array_index_948949 ? add_975933 : sel_975930;
  assign add_975937 = sel_975934 + 8'h01;
  assign sel_975938 = array_index_975625 == array_index_948955 ? add_975937 : sel_975934;
  assign add_975941 = sel_975938 + 8'h01;
  assign sel_975942 = array_index_975625 == array_index_948961 ? add_975941 : sel_975938;
  assign add_975945 = sel_975942 + 8'h01;
  assign sel_975946 = array_index_975625 == array_index_948967 ? add_975945 : sel_975942;
  assign add_975949 = sel_975946 + 8'h01;
  assign sel_975950 = array_index_975625 == array_index_948973 ? add_975949 : sel_975946;
  assign add_975953 = sel_975950 + 8'h01;
  assign sel_975954 = array_index_975625 == array_index_948979 ? add_975953 : sel_975950;
  assign add_975957 = sel_975954 + 8'h01;
  assign sel_975958 = array_index_975625 == array_index_948985 ? add_975957 : sel_975954;
  assign add_975961 = sel_975958 + 8'h01;
  assign sel_975962 = array_index_975625 == array_index_948991 ? add_975961 : sel_975958;
  assign add_975965 = sel_975962 + 8'h01;
  assign sel_975966 = array_index_975625 == array_index_948997 ? add_975965 : sel_975962;
  assign add_975969 = sel_975966 + 8'h01;
  assign sel_975970 = array_index_975625 == array_index_949003 ? add_975969 : sel_975966;
  assign add_975973 = sel_975970 + 8'h01;
  assign sel_975974 = array_index_975625 == array_index_949009 ? add_975973 : sel_975970;
  assign add_975977 = sel_975974 + 8'h01;
  assign sel_975978 = array_index_975625 == array_index_949015 ? add_975977 : sel_975974;
  assign add_975981 = sel_975978 + 8'h01;
  assign sel_975982 = array_index_975625 == array_index_949021 ? add_975981 : sel_975978;
  assign add_975985 = sel_975982 + 8'h01;
  assign sel_975986 = array_index_975625 == array_index_949027 ? add_975985 : sel_975982;
  assign add_975989 = sel_975986 + 8'h01;
  assign sel_975990 = array_index_975625 == array_index_949033 ? add_975989 : sel_975986;
  assign add_975993 = sel_975990 + 8'h01;
  assign sel_975994 = array_index_975625 == array_index_949039 ? add_975993 : sel_975990;
  assign add_975997 = sel_975994 + 8'h01;
  assign sel_975998 = array_index_975625 == array_index_949045 ? add_975997 : sel_975994;
  assign add_976001 = sel_975998 + 8'h01;
  assign sel_976002 = array_index_975625 == array_index_949051 ? add_976001 : sel_975998;
  assign add_976005 = sel_976002 + 8'h01;
  assign sel_976006 = array_index_975625 == array_index_949057 ? add_976005 : sel_976002;
  assign add_976009 = sel_976006 + 8'h01;
  assign sel_976010 = array_index_975625 == array_index_949063 ? add_976009 : sel_976006;
  assign add_976013 = sel_976010 + 8'h01;
  assign sel_976014 = array_index_975625 == array_index_949069 ? add_976013 : sel_976010;
  assign add_976017 = sel_976014 + 8'h01;
  assign sel_976018 = array_index_975625 == array_index_949075 ? add_976017 : sel_976014;
  assign add_976021 = sel_976018 + 8'h01;
  assign sel_976022 = array_index_975625 == array_index_949081 ? add_976021 : sel_976018;
  assign add_976026 = sel_976022 + 8'h01;
  assign array_index_976027 = set1_unflattened[7'h44];
  assign sel_976028 = array_index_975625 == array_index_949087 ? add_976026 : sel_976022;
  assign add_976031 = sel_976028 + 8'h01;
  assign sel_976032 = array_index_976027 == array_index_948483 ? add_976031 : sel_976028;
  assign add_976035 = sel_976032 + 8'h01;
  assign sel_976036 = array_index_976027 == array_index_948487 ? add_976035 : sel_976032;
  assign add_976039 = sel_976036 + 8'h01;
  assign sel_976040 = array_index_976027 == array_index_948495 ? add_976039 : sel_976036;
  assign add_976043 = sel_976040 + 8'h01;
  assign sel_976044 = array_index_976027 == array_index_948503 ? add_976043 : sel_976040;
  assign add_976047 = sel_976044 + 8'h01;
  assign sel_976048 = array_index_976027 == array_index_948511 ? add_976047 : sel_976044;
  assign add_976051 = sel_976048 + 8'h01;
  assign sel_976052 = array_index_976027 == array_index_948519 ? add_976051 : sel_976048;
  assign add_976055 = sel_976052 + 8'h01;
  assign sel_976056 = array_index_976027 == array_index_948527 ? add_976055 : sel_976052;
  assign add_976059 = sel_976056 + 8'h01;
  assign sel_976060 = array_index_976027 == array_index_948535 ? add_976059 : sel_976056;
  assign add_976063 = sel_976060 + 8'h01;
  assign sel_976064 = array_index_976027 == array_index_948541 ? add_976063 : sel_976060;
  assign add_976067 = sel_976064 + 8'h01;
  assign sel_976068 = array_index_976027 == array_index_948547 ? add_976067 : sel_976064;
  assign add_976071 = sel_976068 + 8'h01;
  assign sel_976072 = array_index_976027 == array_index_948553 ? add_976071 : sel_976068;
  assign add_976075 = sel_976072 + 8'h01;
  assign sel_976076 = array_index_976027 == array_index_948559 ? add_976075 : sel_976072;
  assign add_976079 = sel_976076 + 8'h01;
  assign sel_976080 = array_index_976027 == array_index_948565 ? add_976079 : sel_976076;
  assign add_976083 = sel_976080 + 8'h01;
  assign sel_976084 = array_index_976027 == array_index_948571 ? add_976083 : sel_976080;
  assign add_976087 = sel_976084 + 8'h01;
  assign sel_976088 = array_index_976027 == array_index_948577 ? add_976087 : sel_976084;
  assign add_976091 = sel_976088 + 8'h01;
  assign sel_976092 = array_index_976027 == array_index_948583 ? add_976091 : sel_976088;
  assign add_976095 = sel_976092 + 8'h01;
  assign sel_976096 = array_index_976027 == array_index_948589 ? add_976095 : sel_976092;
  assign add_976099 = sel_976096 + 8'h01;
  assign sel_976100 = array_index_976027 == array_index_948595 ? add_976099 : sel_976096;
  assign add_976103 = sel_976100 + 8'h01;
  assign sel_976104 = array_index_976027 == array_index_948601 ? add_976103 : sel_976100;
  assign add_976107 = sel_976104 + 8'h01;
  assign sel_976108 = array_index_976027 == array_index_948607 ? add_976107 : sel_976104;
  assign add_976111 = sel_976108 + 8'h01;
  assign sel_976112 = array_index_976027 == array_index_948613 ? add_976111 : sel_976108;
  assign add_976115 = sel_976112 + 8'h01;
  assign sel_976116 = array_index_976027 == array_index_948619 ? add_976115 : sel_976112;
  assign add_976119 = sel_976116 + 8'h01;
  assign sel_976120 = array_index_976027 == array_index_948625 ? add_976119 : sel_976116;
  assign add_976123 = sel_976120 + 8'h01;
  assign sel_976124 = array_index_976027 == array_index_948631 ? add_976123 : sel_976120;
  assign add_976127 = sel_976124 + 8'h01;
  assign sel_976128 = array_index_976027 == array_index_948637 ? add_976127 : sel_976124;
  assign add_976131 = sel_976128 + 8'h01;
  assign sel_976132 = array_index_976027 == array_index_948643 ? add_976131 : sel_976128;
  assign add_976135 = sel_976132 + 8'h01;
  assign sel_976136 = array_index_976027 == array_index_948649 ? add_976135 : sel_976132;
  assign add_976139 = sel_976136 + 8'h01;
  assign sel_976140 = array_index_976027 == array_index_948655 ? add_976139 : sel_976136;
  assign add_976143 = sel_976140 + 8'h01;
  assign sel_976144 = array_index_976027 == array_index_948661 ? add_976143 : sel_976140;
  assign add_976147 = sel_976144 + 8'h01;
  assign sel_976148 = array_index_976027 == array_index_948667 ? add_976147 : sel_976144;
  assign add_976151 = sel_976148 + 8'h01;
  assign sel_976152 = array_index_976027 == array_index_948673 ? add_976151 : sel_976148;
  assign add_976155 = sel_976152 + 8'h01;
  assign sel_976156 = array_index_976027 == array_index_948679 ? add_976155 : sel_976152;
  assign add_976159 = sel_976156 + 8'h01;
  assign sel_976160 = array_index_976027 == array_index_948685 ? add_976159 : sel_976156;
  assign add_976163 = sel_976160 + 8'h01;
  assign sel_976164 = array_index_976027 == array_index_948691 ? add_976163 : sel_976160;
  assign add_976167 = sel_976164 + 8'h01;
  assign sel_976168 = array_index_976027 == array_index_948697 ? add_976167 : sel_976164;
  assign add_976171 = sel_976168 + 8'h01;
  assign sel_976172 = array_index_976027 == array_index_948703 ? add_976171 : sel_976168;
  assign add_976175 = sel_976172 + 8'h01;
  assign sel_976176 = array_index_976027 == array_index_948709 ? add_976175 : sel_976172;
  assign add_976179 = sel_976176 + 8'h01;
  assign sel_976180 = array_index_976027 == array_index_948715 ? add_976179 : sel_976176;
  assign add_976183 = sel_976180 + 8'h01;
  assign sel_976184 = array_index_976027 == array_index_948721 ? add_976183 : sel_976180;
  assign add_976187 = sel_976184 + 8'h01;
  assign sel_976188 = array_index_976027 == array_index_948727 ? add_976187 : sel_976184;
  assign add_976191 = sel_976188 + 8'h01;
  assign sel_976192 = array_index_976027 == array_index_948733 ? add_976191 : sel_976188;
  assign add_976195 = sel_976192 + 8'h01;
  assign sel_976196 = array_index_976027 == array_index_948739 ? add_976195 : sel_976192;
  assign add_976199 = sel_976196 + 8'h01;
  assign sel_976200 = array_index_976027 == array_index_948745 ? add_976199 : sel_976196;
  assign add_976203 = sel_976200 + 8'h01;
  assign sel_976204 = array_index_976027 == array_index_948751 ? add_976203 : sel_976200;
  assign add_976207 = sel_976204 + 8'h01;
  assign sel_976208 = array_index_976027 == array_index_948757 ? add_976207 : sel_976204;
  assign add_976211 = sel_976208 + 8'h01;
  assign sel_976212 = array_index_976027 == array_index_948763 ? add_976211 : sel_976208;
  assign add_976215 = sel_976212 + 8'h01;
  assign sel_976216 = array_index_976027 == array_index_948769 ? add_976215 : sel_976212;
  assign add_976219 = sel_976216 + 8'h01;
  assign sel_976220 = array_index_976027 == array_index_948775 ? add_976219 : sel_976216;
  assign add_976223 = sel_976220 + 8'h01;
  assign sel_976224 = array_index_976027 == array_index_948781 ? add_976223 : sel_976220;
  assign add_976227 = sel_976224 + 8'h01;
  assign sel_976228 = array_index_976027 == array_index_948787 ? add_976227 : sel_976224;
  assign add_976231 = sel_976228 + 8'h01;
  assign sel_976232 = array_index_976027 == array_index_948793 ? add_976231 : sel_976228;
  assign add_976235 = sel_976232 + 8'h01;
  assign sel_976236 = array_index_976027 == array_index_948799 ? add_976235 : sel_976232;
  assign add_976239 = sel_976236 + 8'h01;
  assign sel_976240 = array_index_976027 == array_index_948805 ? add_976239 : sel_976236;
  assign add_976243 = sel_976240 + 8'h01;
  assign sel_976244 = array_index_976027 == array_index_948811 ? add_976243 : sel_976240;
  assign add_976247 = sel_976244 + 8'h01;
  assign sel_976248 = array_index_976027 == array_index_948817 ? add_976247 : sel_976244;
  assign add_976251 = sel_976248 + 8'h01;
  assign sel_976252 = array_index_976027 == array_index_948823 ? add_976251 : sel_976248;
  assign add_976255 = sel_976252 + 8'h01;
  assign sel_976256 = array_index_976027 == array_index_948829 ? add_976255 : sel_976252;
  assign add_976259 = sel_976256 + 8'h01;
  assign sel_976260 = array_index_976027 == array_index_948835 ? add_976259 : sel_976256;
  assign add_976263 = sel_976260 + 8'h01;
  assign sel_976264 = array_index_976027 == array_index_948841 ? add_976263 : sel_976260;
  assign add_976267 = sel_976264 + 8'h01;
  assign sel_976268 = array_index_976027 == array_index_948847 ? add_976267 : sel_976264;
  assign add_976271 = sel_976268 + 8'h01;
  assign sel_976272 = array_index_976027 == array_index_948853 ? add_976271 : sel_976268;
  assign add_976275 = sel_976272 + 8'h01;
  assign sel_976276 = array_index_976027 == array_index_948859 ? add_976275 : sel_976272;
  assign add_976279 = sel_976276 + 8'h01;
  assign sel_976280 = array_index_976027 == array_index_948865 ? add_976279 : sel_976276;
  assign add_976283 = sel_976280 + 8'h01;
  assign sel_976284 = array_index_976027 == array_index_948871 ? add_976283 : sel_976280;
  assign add_976287 = sel_976284 + 8'h01;
  assign sel_976288 = array_index_976027 == array_index_948877 ? add_976287 : sel_976284;
  assign add_976291 = sel_976288 + 8'h01;
  assign sel_976292 = array_index_976027 == array_index_948883 ? add_976291 : sel_976288;
  assign add_976295 = sel_976292 + 8'h01;
  assign sel_976296 = array_index_976027 == array_index_948889 ? add_976295 : sel_976292;
  assign add_976299 = sel_976296 + 8'h01;
  assign sel_976300 = array_index_976027 == array_index_948895 ? add_976299 : sel_976296;
  assign add_976303 = sel_976300 + 8'h01;
  assign sel_976304 = array_index_976027 == array_index_948901 ? add_976303 : sel_976300;
  assign add_976307 = sel_976304 + 8'h01;
  assign sel_976308 = array_index_976027 == array_index_948907 ? add_976307 : sel_976304;
  assign add_976311 = sel_976308 + 8'h01;
  assign sel_976312 = array_index_976027 == array_index_948913 ? add_976311 : sel_976308;
  assign add_976315 = sel_976312 + 8'h01;
  assign sel_976316 = array_index_976027 == array_index_948919 ? add_976315 : sel_976312;
  assign add_976319 = sel_976316 + 8'h01;
  assign sel_976320 = array_index_976027 == array_index_948925 ? add_976319 : sel_976316;
  assign add_976323 = sel_976320 + 8'h01;
  assign sel_976324 = array_index_976027 == array_index_948931 ? add_976323 : sel_976320;
  assign add_976327 = sel_976324 + 8'h01;
  assign sel_976328 = array_index_976027 == array_index_948937 ? add_976327 : sel_976324;
  assign add_976331 = sel_976328 + 8'h01;
  assign sel_976332 = array_index_976027 == array_index_948943 ? add_976331 : sel_976328;
  assign add_976335 = sel_976332 + 8'h01;
  assign sel_976336 = array_index_976027 == array_index_948949 ? add_976335 : sel_976332;
  assign add_976339 = sel_976336 + 8'h01;
  assign sel_976340 = array_index_976027 == array_index_948955 ? add_976339 : sel_976336;
  assign add_976343 = sel_976340 + 8'h01;
  assign sel_976344 = array_index_976027 == array_index_948961 ? add_976343 : sel_976340;
  assign add_976347 = sel_976344 + 8'h01;
  assign sel_976348 = array_index_976027 == array_index_948967 ? add_976347 : sel_976344;
  assign add_976351 = sel_976348 + 8'h01;
  assign sel_976352 = array_index_976027 == array_index_948973 ? add_976351 : sel_976348;
  assign add_976355 = sel_976352 + 8'h01;
  assign sel_976356 = array_index_976027 == array_index_948979 ? add_976355 : sel_976352;
  assign add_976359 = sel_976356 + 8'h01;
  assign sel_976360 = array_index_976027 == array_index_948985 ? add_976359 : sel_976356;
  assign add_976363 = sel_976360 + 8'h01;
  assign sel_976364 = array_index_976027 == array_index_948991 ? add_976363 : sel_976360;
  assign add_976367 = sel_976364 + 8'h01;
  assign sel_976368 = array_index_976027 == array_index_948997 ? add_976367 : sel_976364;
  assign add_976371 = sel_976368 + 8'h01;
  assign sel_976372 = array_index_976027 == array_index_949003 ? add_976371 : sel_976368;
  assign add_976375 = sel_976372 + 8'h01;
  assign sel_976376 = array_index_976027 == array_index_949009 ? add_976375 : sel_976372;
  assign add_976379 = sel_976376 + 8'h01;
  assign sel_976380 = array_index_976027 == array_index_949015 ? add_976379 : sel_976376;
  assign add_976383 = sel_976380 + 8'h01;
  assign sel_976384 = array_index_976027 == array_index_949021 ? add_976383 : sel_976380;
  assign add_976387 = sel_976384 + 8'h01;
  assign sel_976388 = array_index_976027 == array_index_949027 ? add_976387 : sel_976384;
  assign add_976391 = sel_976388 + 8'h01;
  assign sel_976392 = array_index_976027 == array_index_949033 ? add_976391 : sel_976388;
  assign add_976395 = sel_976392 + 8'h01;
  assign sel_976396 = array_index_976027 == array_index_949039 ? add_976395 : sel_976392;
  assign add_976399 = sel_976396 + 8'h01;
  assign sel_976400 = array_index_976027 == array_index_949045 ? add_976399 : sel_976396;
  assign add_976403 = sel_976400 + 8'h01;
  assign sel_976404 = array_index_976027 == array_index_949051 ? add_976403 : sel_976400;
  assign add_976407 = sel_976404 + 8'h01;
  assign sel_976408 = array_index_976027 == array_index_949057 ? add_976407 : sel_976404;
  assign add_976411 = sel_976408 + 8'h01;
  assign sel_976412 = array_index_976027 == array_index_949063 ? add_976411 : sel_976408;
  assign add_976415 = sel_976412 + 8'h01;
  assign sel_976416 = array_index_976027 == array_index_949069 ? add_976415 : sel_976412;
  assign add_976419 = sel_976416 + 8'h01;
  assign sel_976420 = array_index_976027 == array_index_949075 ? add_976419 : sel_976416;
  assign add_976423 = sel_976420 + 8'h01;
  assign sel_976424 = array_index_976027 == array_index_949081 ? add_976423 : sel_976420;
  assign add_976428 = sel_976424 + 8'h01;
  assign array_index_976429 = set1_unflattened[7'h45];
  assign sel_976430 = array_index_976027 == array_index_949087 ? add_976428 : sel_976424;
  assign add_976433 = sel_976430 + 8'h01;
  assign sel_976434 = array_index_976429 == array_index_948483 ? add_976433 : sel_976430;
  assign add_976437 = sel_976434 + 8'h01;
  assign sel_976438 = array_index_976429 == array_index_948487 ? add_976437 : sel_976434;
  assign add_976441 = sel_976438 + 8'h01;
  assign sel_976442 = array_index_976429 == array_index_948495 ? add_976441 : sel_976438;
  assign add_976445 = sel_976442 + 8'h01;
  assign sel_976446 = array_index_976429 == array_index_948503 ? add_976445 : sel_976442;
  assign add_976449 = sel_976446 + 8'h01;
  assign sel_976450 = array_index_976429 == array_index_948511 ? add_976449 : sel_976446;
  assign add_976453 = sel_976450 + 8'h01;
  assign sel_976454 = array_index_976429 == array_index_948519 ? add_976453 : sel_976450;
  assign add_976457 = sel_976454 + 8'h01;
  assign sel_976458 = array_index_976429 == array_index_948527 ? add_976457 : sel_976454;
  assign add_976461 = sel_976458 + 8'h01;
  assign sel_976462 = array_index_976429 == array_index_948535 ? add_976461 : sel_976458;
  assign add_976465 = sel_976462 + 8'h01;
  assign sel_976466 = array_index_976429 == array_index_948541 ? add_976465 : sel_976462;
  assign add_976469 = sel_976466 + 8'h01;
  assign sel_976470 = array_index_976429 == array_index_948547 ? add_976469 : sel_976466;
  assign add_976473 = sel_976470 + 8'h01;
  assign sel_976474 = array_index_976429 == array_index_948553 ? add_976473 : sel_976470;
  assign add_976477 = sel_976474 + 8'h01;
  assign sel_976478 = array_index_976429 == array_index_948559 ? add_976477 : sel_976474;
  assign add_976481 = sel_976478 + 8'h01;
  assign sel_976482 = array_index_976429 == array_index_948565 ? add_976481 : sel_976478;
  assign add_976485 = sel_976482 + 8'h01;
  assign sel_976486 = array_index_976429 == array_index_948571 ? add_976485 : sel_976482;
  assign add_976489 = sel_976486 + 8'h01;
  assign sel_976490 = array_index_976429 == array_index_948577 ? add_976489 : sel_976486;
  assign add_976493 = sel_976490 + 8'h01;
  assign sel_976494 = array_index_976429 == array_index_948583 ? add_976493 : sel_976490;
  assign add_976497 = sel_976494 + 8'h01;
  assign sel_976498 = array_index_976429 == array_index_948589 ? add_976497 : sel_976494;
  assign add_976501 = sel_976498 + 8'h01;
  assign sel_976502 = array_index_976429 == array_index_948595 ? add_976501 : sel_976498;
  assign add_976505 = sel_976502 + 8'h01;
  assign sel_976506 = array_index_976429 == array_index_948601 ? add_976505 : sel_976502;
  assign add_976509 = sel_976506 + 8'h01;
  assign sel_976510 = array_index_976429 == array_index_948607 ? add_976509 : sel_976506;
  assign add_976513 = sel_976510 + 8'h01;
  assign sel_976514 = array_index_976429 == array_index_948613 ? add_976513 : sel_976510;
  assign add_976517 = sel_976514 + 8'h01;
  assign sel_976518 = array_index_976429 == array_index_948619 ? add_976517 : sel_976514;
  assign add_976521 = sel_976518 + 8'h01;
  assign sel_976522 = array_index_976429 == array_index_948625 ? add_976521 : sel_976518;
  assign add_976525 = sel_976522 + 8'h01;
  assign sel_976526 = array_index_976429 == array_index_948631 ? add_976525 : sel_976522;
  assign add_976529 = sel_976526 + 8'h01;
  assign sel_976530 = array_index_976429 == array_index_948637 ? add_976529 : sel_976526;
  assign add_976533 = sel_976530 + 8'h01;
  assign sel_976534 = array_index_976429 == array_index_948643 ? add_976533 : sel_976530;
  assign add_976537 = sel_976534 + 8'h01;
  assign sel_976538 = array_index_976429 == array_index_948649 ? add_976537 : sel_976534;
  assign add_976541 = sel_976538 + 8'h01;
  assign sel_976542 = array_index_976429 == array_index_948655 ? add_976541 : sel_976538;
  assign add_976545 = sel_976542 + 8'h01;
  assign sel_976546 = array_index_976429 == array_index_948661 ? add_976545 : sel_976542;
  assign add_976549 = sel_976546 + 8'h01;
  assign sel_976550 = array_index_976429 == array_index_948667 ? add_976549 : sel_976546;
  assign add_976553 = sel_976550 + 8'h01;
  assign sel_976554 = array_index_976429 == array_index_948673 ? add_976553 : sel_976550;
  assign add_976557 = sel_976554 + 8'h01;
  assign sel_976558 = array_index_976429 == array_index_948679 ? add_976557 : sel_976554;
  assign add_976561 = sel_976558 + 8'h01;
  assign sel_976562 = array_index_976429 == array_index_948685 ? add_976561 : sel_976558;
  assign add_976565 = sel_976562 + 8'h01;
  assign sel_976566 = array_index_976429 == array_index_948691 ? add_976565 : sel_976562;
  assign add_976569 = sel_976566 + 8'h01;
  assign sel_976570 = array_index_976429 == array_index_948697 ? add_976569 : sel_976566;
  assign add_976573 = sel_976570 + 8'h01;
  assign sel_976574 = array_index_976429 == array_index_948703 ? add_976573 : sel_976570;
  assign add_976577 = sel_976574 + 8'h01;
  assign sel_976578 = array_index_976429 == array_index_948709 ? add_976577 : sel_976574;
  assign add_976581 = sel_976578 + 8'h01;
  assign sel_976582 = array_index_976429 == array_index_948715 ? add_976581 : sel_976578;
  assign add_976585 = sel_976582 + 8'h01;
  assign sel_976586 = array_index_976429 == array_index_948721 ? add_976585 : sel_976582;
  assign add_976589 = sel_976586 + 8'h01;
  assign sel_976590 = array_index_976429 == array_index_948727 ? add_976589 : sel_976586;
  assign add_976593 = sel_976590 + 8'h01;
  assign sel_976594 = array_index_976429 == array_index_948733 ? add_976593 : sel_976590;
  assign add_976597 = sel_976594 + 8'h01;
  assign sel_976598 = array_index_976429 == array_index_948739 ? add_976597 : sel_976594;
  assign add_976601 = sel_976598 + 8'h01;
  assign sel_976602 = array_index_976429 == array_index_948745 ? add_976601 : sel_976598;
  assign add_976605 = sel_976602 + 8'h01;
  assign sel_976606 = array_index_976429 == array_index_948751 ? add_976605 : sel_976602;
  assign add_976609 = sel_976606 + 8'h01;
  assign sel_976610 = array_index_976429 == array_index_948757 ? add_976609 : sel_976606;
  assign add_976613 = sel_976610 + 8'h01;
  assign sel_976614 = array_index_976429 == array_index_948763 ? add_976613 : sel_976610;
  assign add_976617 = sel_976614 + 8'h01;
  assign sel_976618 = array_index_976429 == array_index_948769 ? add_976617 : sel_976614;
  assign add_976621 = sel_976618 + 8'h01;
  assign sel_976622 = array_index_976429 == array_index_948775 ? add_976621 : sel_976618;
  assign add_976625 = sel_976622 + 8'h01;
  assign sel_976626 = array_index_976429 == array_index_948781 ? add_976625 : sel_976622;
  assign add_976629 = sel_976626 + 8'h01;
  assign sel_976630 = array_index_976429 == array_index_948787 ? add_976629 : sel_976626;
  assign add_976633 = sel_976630 + 8'h01;
  assign sel_976634 = array_index_976429 == array_index_948793 ? add_976633 : sel_976630;
  assign add_976637 = sel_976634 + 8'h01;
  assign sel_976638 = array_index_976429 == array_index_948799 ? add_976637 : sel_976634;
  assign add_976641 = sel_976638 + 8'h01;
  assign sel_976642 = array_index_976429 == array_index_948805 ? add_976641 : sel_976638;
  assign add_976645 = sel_976642 + 8'h01;
  assign sel_976646 = array_index_976429 == array_index_948811 ? add_976645 : sel_976642;
  assign add_976649 = sel_976646 + 8'h01;
  assign sel_976650 = array_index_976429 == array_index_948817 ? add_976649 : sel_976646;
  assign add_976653 = sel_976650 + 8'h01;
  assign sel_976654 = array_index_976429 == array_index_948823 ? add_976653 : sel_976650;
  assign add_976657 = sel_976654 + 8'h01;
  assign sel_976658 = array_index_976429 == array_index_948829 ? add_976657 : sel_976654;
  assign add_976661 = sel_976658 + 8'h01;
  assign sel_976662 = array_index_976429 == array_index_948835 ? add_976661 : sel_976658;
  assign add_976665 = sel_976662 + 8'h01;
  assign sel_976666 = array_index_976429 == array_index_948841 ? add_976665 : sel_976662;
  assign add_976669 = sel_976666 + 8'h01;
  assign sel_976670 = array_index_976429 == array_index_948847 ? add_976669 : sel_976666;
  assign add_976673 = sel_976670 + 8'h01;
  assign sel_976674 = array_index_976429 == array_index_948853 ? add_976673 : sel_976670;
  assign add_976677 = sel_976674 + 8'h01;
  assign sel_976678 = array_index_976429 == array_index_948859 ? add_976677 : sel_976674;
  assign add_976681 = sel_976678 + 8'h01;
  assign sel_976682 = array_index_976429 == array_index_948865 ? add_976681 : sel_976678;
  assign add_976685 = sel_976682 + 8'h01;
  assign sel_976686 = array_index_976429 == array_index_948871 ? add_976685 : sel_976682;
  assign add_976689 = sel_976686 + 8'h01;
  assign sel_976690 = array_index_976429 == array_index_948877 ? add_976689 : sel_976686;
  assign add_976693 = sel_976690 + 8'h01;
  assign sel_976694 = array_index_976429 == array_index_948883 ? add_976693 : sel_976690;
  assign add_976697 = sel_976694 + 8'h01;
  assign sel_976698 = array_index_976429 == array_index_948889 ? add_976697 : sel_976694;
  assign add_976701 = sel_976698 + 8'h01;
  assign sel_976702 = array_index_976429 == array_index_948895 ? add_976701 : sel_976698;
  assign add_976705 = sel_976702 + 8'h01;
  assign sel_976706 = array_index_976429 == array_index_948901 ? add_976705 : sel_976702;
  assign add_976709 = sel_976706 + 8'h01;
  assign sel_976710 = array_index_976429 == array_index_948907 ? add_976709 : sel_976706;
  assign add_976713 = sel_976710 + 8'h01;
  assign sel_976714 = array_index_976429 == array_index_948913 ? add_976713 : sel_976710;
  assign add_976717 = sel_976714 + 8'h01;
  assign sel_976718 = array_index_976429 == array_index_948919 ? add_976717 : sel_976714;
  assign add_976721 = sel_976718 + 8'h01;
  assign sel_976722 = array_index_976429 == array_index_948925 ? add_976721 : sel_976718;
  assign add_976725 = sel_976722 + 8'h01;
  assign sel_976726 = array_index_976429 == array_index_948931 ? add_976725 : sel_976722;
  assign add_976729 = sel_976726 + 8'h01;
  assign sel_976730 = array_index_976429 == array_index_948937 ? add_976729 : sel_976726;
  assign add_976733 = sel_976730 + 8'h01;
  assign sel_976734 = array_index_976429 == array_index_948943 ? add_976733 : sel_976730;
  assign add_976737 = sel_976734 + 8'h01;
  assign sel_976738 = array_index_976429 == array_index_948949 ? add_976737 : sel_976734;
  assign add_976741 = sel_976738 + 8'h01;
  assign sel_976742 = array_index_976429 == array_index_948955 ? add_976741 : sel_976738;
  assign add_976745 = sel_976742 + 8'h01;
  assign sel_976746 = array_index_976429 == array_index_948961 ? add_976745 : sel_976742;
  assign add_976749 = sel_976746 + 8'h01;
  assign sel_976750 = array_index_976429 == array_index_948967 ? add_976749 : sel_976746;
  assign add_976753 = sel_976750 + 8'h01;
  assign sel_976754 = array_index_976429 == array_index_948973 ? add_976753 : sel_976750;
  assign add_976757 = sel_976754 + 8'h01;
  assign sel_976758 = array_index_976429 == array_index_948979 ? add_976757 : sel_976754;
  assign add_976761 = sel_976758 + 8'h01;
  assign sel_976762 = array_index_976429 == array_index_948985 ? add_976761 : sel_976758;
  assign add_976765 = sel_976762 + 8'h01;
  assign sel_976766 = array_index_976429 == array_index_948991 ? add_976765 : sel_976762;
  assign add_976769 = sel_976766 + 8'h01;
  assign sel_976770 = array_index_976429 == array_index_948997 ? add_976769 : sel_976766;
  assign add_976773 = sel_976770 + 8'h01;
  assign sel_976774 = array_index_976429 == array_index_949003 ? add_976773 : sel_976770;
  assign add_976777 = sel_976774 + 8'h01;
  assign sel_976778 = array_index_976429 == array_index_949009 ? add_976777 : sel_976774;
  assign add_976781 = sel_976778 + 8'h01;
  assign sel_976782 = array_index_976429 == array_index_949015 ? add_976781 : sel_976778;
  assign add_976785 = sel_976782 + 8'h01;
  assign sel_976786 = array_index_976429 == array_index_949021 ? add_976785 : sel_976782;
  assign add_976789 = sel_976786 + 8'h01;
  assign sel_976790 = array_index_976429 == array_index_949027 ? add_976789 : sel_976786;
  assign add_976793 = sel_976790 + 8'h01;
  assign sel_976794 = array_index_976429 == array_index_949033 ? add_976793 : sel_976790;
  assign add_976797 = sel_976794 + 8'h01;
  assign sel_976798 = array_index_976429 == array_index_949039 ? add_976797 : sel_976794;
  assign add_976801 = sel_976798 + 8'h01;
  assign sel_976802 = array_index_976429 == array_index_949045 ? add_976801 : sel_976798;
  assign add_976805 = sel_976802 + 8'h01;
  assign sel_976806 = array_index_976429 == array_index_949051 ? add_976805 : sel_976802;
  assign add_976809 = sel_976806 + 8'h01;
  assign sel_976810 = array_index_976429 == array_index_949057 ? add_976809 : sel_976806;
  assign add_976813 = sel_976810 + 8'h01;
  assign sel_976814 = array_index_976429 == array_index_949063 ? add_976813 : sel_976810;
  assign add_976817 = sel_976814 + 8'h01;
  assign sel_976818 = array_index_976429 == array_index_949069 ? add_976817 : sel_976814;
  assign add_976821 = sel_976818 + 8'h01;
  assign sel_976822 = array_index_976429 == array_index_949075 ? add_976821 : sel_976818;
  assign add_976825 = sel_976822 + 8'h01;
  assign sel_976826 = array_index_976429 == array_index_949081 ? add_976825 : sel_976822;
  assign add_976830 = sel_976826 + 8'h01;
  assign array_index_976831 = set1_unflattened[7'h46];
  assign sel_976832 = array_index_976429 == array_index_949087 ? add_976830 : sel_976826;
  assign add_976835 = sel_976832 + 8'h01;
  assign sel_976836 = array_index_976831 == array_index_948483 ? add_976835 : sel_976832;
  assign add_976839 = sel_976836 + 8'h01;
  assign sel_976840 = array_index_976831 == array_index_948487 ? add_976839 : sel_976836;
  assign add_976843 = sel_976840 + 8'h01;
  assign sel_976844 = array_index_976831 == array_index_948495 ? add_976843 : sel_976840;
  assign add_976847 = sel_976844 + 8'h01;
  assign sel_976848 = array_index_976831 == array_index_948503 ? add_976847 : sel_976844;
  assign add_976851 = sel_976848 + 8'h01;
  assign sel_976852 = array_index_976831 == array_index_948511 ? add_976851 : sel_976848;
  assign add_976855 = sel_976852 + 8'h01;
  assign sel_976856 = array_index_976831 == array_index_948519 ? add_976855 : sel_976852;
  assign add_976859 = sel_976856 + 8'h01;
  assign sel_976860 = array_index_976831 == array_index_948527 ? add_976859 : sel_976856;
  assign add_976863 = sel_976860 + 8'h01;
  assign sel_976864 = array_index_976831 == array_index_948535 ? add_976863 : sel_976860;
  assign add_976867 = sel_976864 + 8'h01;
  assign sel_976868 = array_index_976831 == array_index_948541 ? add_976867 : sel_976864;
  assign add_976871 = sel_976868 + 8'h01;
  assign sel_976872 = array_index_976831 == array_index_948547 ? add_976871 : sel_976868;
  assign add_976875 = sel_976872 + 8'h01;
  assign sel_976876 = array_index_976831 == array_index_948553 ? add_976875 : sel_976872;
  assign add_976879 = sel_976876 + 8'h01;
  assign sel_976880 = array_index_976831 == array_index_948559 ? add_976879 : sel_976876;
  assign add_976883 = sel_976880 + 8'h01;
  assign sel_976884 = array_index_976831 == array_index_948565 ? add_976883 : sel_976880;
  assign add_976887 = sel_976884 + 8'h01;
  assign sel_976888 = array_index_976831 == array_index_948571 ? add_976887 : sel_976884;
  assign add_976891 = sel_976888 + 8'h01;
  assign sel_976892 = array_index_976831 == array_index_948577 ? add_976891 : sel_976888;
  assign add_976895 = sel_976892 + 8'h01;
  assign sel_976896 = array_index_976831 == array_index_948583 ? add_976895 : sel_976892;
  assign add_976899 = sel_976896 + 8'h01;
  assign sel_976900 = array_index_976831 == array_index_948589 ? add_976899 : sel_976896;
  assign add_976903 = sel_976900 + 8'h01;
  assign sel_976904 = array_index_976831 == array_index_948595 ? add_976903 : sel_976900;
  assign add_976907 = sel_976904 + 8'h01;
  assign sel_976908 = array_index_976831 == array_index_948601 ? add_976907 : sel_976904;
  assign add_976911 = sel_976908 + 8'h01;
  assign sel_976912 = array_index_976831 == array_index_948607 ? add_976911 : sel_976908;
  assign add_976915 = sel_976912 + 8'h01;
  assign sel_976916 = array_index_976831 == array_index_948613 ? add_976915 : sel_976912;
  assign add_976919 = sel_976916 + 8'h01;
  assign sel_976920 = array_index_976831 == array_index_948619 ? add_976919 : sel_976916;
  assign add_976923 = sel_976920 + 8'h01;
  assign sel_976924 = array_index_976831 == array_index_948625 ? add_976923 : sel_976920;
  assign add_976927 = sel_976924 + 8'h01;
  assign sel_976928 = array_index_976831 == array_index_948631 ? add_976927 : sel_976924;
  assign add_976931 = sel_976928 + 8'h01;
  assign sel_976932 = array_index_976831 == array_index_948637 ? add_976931 : sel_976928;
  assign add_976935 = sel_976932 + 8'h01;
  assign sel_976936 = array_index_976831 == array_index_948643 ? add_976935 : sel_976932;
  assign add_976939 = sel_976936 + 8'h01;
  assign sel_976940 = array_index_976831 == array_index_948649 ? add_976939 : sel_976936;
  assign add_976943 = sel_976940 + 8'h01;
  assign sel_976944 = array_index_976831 == array_index_948655 ? add_976943 : sel_976940;
  assign add_976947 = sel_976944 + 8'h01;
  assign sel_976948 = array_index_976831 == array_index_948661 ? add_976947 : sel_976944;
  assign add_976951 = sel_976948 + 8'h01;
  assign sel_976952 = array_index_976831 == array_index_948667 ? add_976951 : sel_976948;
  assign add_976955 = sel_976952 + 8'h01;
  assign sel_976956 = array_index_976831 == array_index_948673 ? add_976955 : sel_976952;
  assign add_976959 = sel_976956 + 8'h01;
  assign sel_976960 = array_index_976831 == array_index_948679 ? add_976959 : sel_976956;
  assign add_976963 = sel_976960 + 8'h01;
  assign sel_976964 = array_index_976831 == array_index_948685 ? add_976963 : sel_976960;
  assign add_976967 = sel_976964 + 8'h01;
  assign sel_976968 = array_index_976831 == array_index_948691 ? add_976967 : sel_976964;
  assign add_976971 = sel_976968 + 8'h01;
  assign sel_976972 = array_index_976831 == array_index_948697 ? add_976971 : sel_976968;
  assign add_976975 = sel_976972 + 8'h01;
  assign sel_976976 = array_index_976831 == array_index_948703 ? add_976975 : sel_976972;
  assign add_976979 = sel_976976 + 8'h01;
  assign sel_976980 = array_index_976831 == array_index_948709 ? add_976979 : sel_976976;
  assign add_976983 = sel_976980 + 8'h01;
  assign sel_976984 = array_index_976831 == array_index_948715 ? add_976983 : sel_976980;
  assign add_976987 = sel_976984 + 8'h01;
  assign sel_976988 = array_index_976831 == array_index_948721 ? add_976987 : sel_976984;
  assign add_976991 = sel_976988 + 8'h01;
  assign sel_976992 = array_index_976831 == array_index_948727 ? add_976991 : sel_976988;
  assign add_976995 = sel_976992 + 8'h01;
  assign sel_976996 = array_index_976831 == array_index_948733 ? add_976995 : sel_976992;
  assign add_976999 = sel_976996 + 8'h01;
  assign sel_977000 = array_index_976831 == array_index_948739 ? add_976999 : sel_976996;
  assign add_977003 = sel_977000 + 8'h01;
  assign sel_977004 = array_index_976831 == array_index_948745 ? add_977003 : sel_977000;
  assign add_977007 = sel_977004 + 8'h01;
  assign sel_977008 = array_index_976831 == array_index_948751 ? add_977007 : sel_977004;
  assign add_977011 = sel_977008 + 8'h01;
  assign sel_977012 = array_index_976831 == array_index_948757 ? add_977011 : sel_977008;
  assign add_977015 = sel_977012 + 8'h01;
  assign sel_977016 = array_index_976831 == array_index_948763 ? add_977015 : sel_977012;
  assign add_977019 = sel_977016 + 8'h01;
  assign sel_977020 = array_index_976831 == array_index_948769 ? add_977019 : sel_977016;
  assign add_977023 = sel_977020 + 8'h01;
  assign sel_977024 = array_index_976831 == array_index_948775 ? add_977023 : sel_977020;
  assign add_977027 = sel_977024 + 8'h01;
  assign sel_977028 = array_index_976831 == array_index_948781 ? add_977027 : sel_977024;
  assign add_977031 = sel_977028 + 8'h01;
  assign sel_977032 = array_index_976831 == array_index_948787 ? add_977031 : sel_977028;
  assign add_977035 = sel_977032 + 8'h01;
  assign sel_977036 = array_index_976831 == array_index_948793 ? add_977035 : sel_977032;
  assign add_977039 = sel_977036 + 8'h01;
  assign sel_977040 = array_index_976831 == array_index_948799 ? add_977039 : sel_977036;
  assign add_977043 = sel_977040 + 8'h01;
  assign sel_977044 = array_index_976831 == array_index_948805 ? add_977043 : sel_977040;
  assign add_977047 = sel_977044 + 8'h01;
  assign sel_977048 = array_index_976831 == array_index_948811 ? add_977047 : sel_977044;
  assign add_977051 = sel_977048 + 8'h01;
  assign sel_977052 = array_index_976831 == array_index_948817 ? add_977051 : sel_977048;
  assign add_977055 = sel_977052 + 8'h01;
  assign sel_977056 = array_index_976831 == array_index_948823 ? add_977055 : sel_977052;
  assign add_977059 = sel_977056 + 8'h01;
  assign sel_977060 = array_index_976831 == array_index_948829 ? add_977059 : sel_977056;
  assign add_977063 = sel_977060 + 8'h01;
  assign sel_977064 = array_index_976831 == array_index_948835 ? add_977063 : sel_977060;
  assign add_977067 = sel_977064 + 8'h01;
  assign sel_977068 = array_index_976831 == array_index_948841 ? add_977067 : sel_977064;
  assign add_977071 = sel_977068 + 8'h01;
  assign sel_977072 = array_index_976831 == array_index_948847 ? add_977071 : sel_977068;
  assign add_977075 = sel_977072 + 8'h01;
  assign sel_977076 = array_index_976831 == array_index_948853 ? add_977075 : sel_977072;
  assign add_977079 = sel_977076 + 8'h01;
  assign sel_977080 = array_index_976831 == array_index_948859 ? add_977079 : sel_977076;
  assign add_977083 = sel_977080 + 8'h01;
  assign sel_977084 = array_index_976831 == array_index_948865 ? add_977083 : sel_977080;
  assign add_977087 = sel_977084 + 8'h01;
  assign sel_977088 = array_index_976831 == array_index_948871 ? add_977087 : sel_977084;
  assign add_977091 = sel_977088 + 8'h01;
  assign sel_977092 = array_index_976831 == array_index_948877 ? add_977091 : sel_977088;
  assign add_977095 = sel_977092 + 8'h01;
  assign sel_977096 = array_index_976831 == array_index_948883 ? add_977095 : sel_977092;
  assign add_977099 = sel_977096 + 8'h01;
  assign sel_977100 = array_index_976831 == array_index_948889 ? add_977099 : sel_977096;
  assign add_977103 = sel_977100 + 8'h01;
  assign sel_977104 = array_index_976831 == array_index_948895 ? add_977103 : sel_977100;
  assign add_977107 = sel_977104 + 8'h01;
  assign sel_977108 = array_index_976831 == array_index_948901 ? add_977107 : sel_977104;
  assign add_977111 = sel_977108 + 8'h01;
  assign sel_977112 = array_index_976831 == array_index_948907 ? add_977111 : sel_977108;
  assign add_977115 = sel_977112 + 8'h01;
  assign sel_977116 = array_index_976831 == array_index_948913 ? add_977115 : sel_977112;
  assign add_977119 = sel_977116 + 8'h01;
  assign sel_977120 = array_index_976831 == array_index_948919 ? add_977119 : sel_977116;
  assign add_977123 = sel_977120 + 8'h01;
  assign sel_977124 = array_index_976831 == array_index_948925 ? add_977123 : sel_977120;
  assign add_977127 = sel_977124 + 8'h01;
  assign sel_977128 = array_index_976831 == array_index_948931 ? add_977127 : sel_977124;
  assign add_977131 = sel_977128 + 8'h01;
  assign sel_977132 = array_index_976831 == array_index_948937 ? add_977131 : sel_977128;
  assign add_977135 = sel_977132 + 8'h01;
  assign sel_977136 = array_index_976831 == array_index_948943 ? add_977135 : sel_977132;
  assign add_977139 = sel_977136 + 8'h01;
  assign sel_977140 = array_index_976831 == array_index_948949 ? add_977139 : sel_977136;
  assign add_977143 = sel_977140 + 8'h01;
  assign sel_977144 = array_index_976831 == array_index_948955 ? add_977143 : sel_977140;
  assign add_977147 = sel_977144 + 8'h01;
  assign sel_977148 = array_index_976831 == array_index_948961 ? add_977147 : sel_977144;
  assign add_977151 = sel_977148 + 8'h01;
  assign sel_977152 = array_index_976831 == array_index_948967 ? add_977151 : sel_977148;
  assign add_977155 = sel_977152 + 8'h01;
  assign sel_977156 = array_index_976831 == array_index_948973 ? add_977155 : sel_977152;
  assign add_977159 = sel_977156 + 8'h01;
  assign sel_977160 = array_index_976831 == array_index_948979 ? add_977159 : sel_977156;
  assign add_977163 = sel_977160 + 8'h01;
  assign sel_977164 = array_index_976831 == array_index_948985 ? add_977163 : sel_977160;
  assign add_977167 = sel_977164 + 8'h01;
  assign sel_977168 = array_index_976831 == array_index_948991 ? add_977167 : sel_977164;
  assign add_977171 = sel_977168 + 8'h01;
  assign sel_977172 = array_index_976831 == array_index_948997 ? add_977171 : sel_977168;
  assign add_977175 = sel_977172 + 8'h01;
  assign sel_977176 = array_index_976831 == array_index_949003 ? add_977175 : sel_977172;
  assign add_977179 = sel_977176 + 8'h01;
  assign sel_977180 = array_index_976831 == array_index_949009 ? add_977179 : sel_977176;
  assign add_977183 = sel_977180 + 8'h01;
  assign sel_977184 = array_index_976831 == array_index_949015 ? add_977183 : sel_977180;
  assign add_977187 = sel_977184 + 8'h01;
  assign sel_977188 = array_index_976831 == array_index_949021 ? add_977187 : sel_977184;
  assign add_977191 = sel_977188 + 8'h01;
  assign sel_977192 = array_index_976831 == array_index_949027 ? add_977191 : sel_977188;
  assign add_977195 = sel_977192 + 8'h01;
  assign sel_977196 = array_index_976831 == array_index_949033 ? add_977195 : sel_977192;
  assign add_977199 = sel_977196 + 8'h01;
  assign sel_977200 = array_index_976831 == array_index_949039 ? add_977199 : sel_977196;
  assign add_977203 = sel_977200 + 8'h01;
  assign sel_977204 = array_index_976831 == array_index_949045 ? add_977203 : sel_977200;
  assign add_977207 = sel_977204 + 8'h01;
  assign sel_977208 = array_index_976831 == array_index_949051 ? add_977207 : sel_977204;
  assign add_977211 = sel_977208 + 8'h01;
  assign sel_977212 = array_index_976831 == array_index_949057 ? add_977211 : sel_977208;
  assign add_977215 = sel_977212 + 8'h01;
  assign sel_977216 = array_index_976831 == array_index_949063 ? add_977215 : sel_977212;
  assign add_977219 = sel_977216 + 8'h01;
  assign sel_977220 = array_index_976831 == array_index_949069 ? add_977219 : sel_977216;
  assign add_977223 = sel_977220 + 8'h01;
  assign sel_977224 = array_index_976831 == array_index_949075 ? add_977223 : sel_977220;
  assign add_977227 = sel_977224 + 8'h01;
  assign sel_977228 = array_index_976831 == array_index_949081 ? add_977227 : sel_977224;
  assign add_977232 = sel_977228 + 8'h01;
  assign array_index_977233 = set1_unflattened[7'h47];
  assign sel_977234 = array_index_976831 == array_index_949087 ? add_977232 : sel_977228;
  assign add_977237 = sel_977234 + 8'h01;
  assign sel_977238 = array_index_977233 == array_index_948483 ? add_977237 : sel_977234;
  assign add_977241 = sel_977238 + 8'h01;
  assign sel_977242 = array_index_977233 == array_index_948487 ? add_977241 : sel_977238;
  assign add_977245 = sel_977242 + 8'h01;
  assign sel_977246 = array_index_977233 == array_index_948495 ? add_977245 : sel_977242;
  assign add_977249 = sel_977246 + 8'h01;
  assign sel_977250 = array_index_977233 == array_index_948503 ? add_977249 : sel_977246;
  assign add_977253 = sel_977250 + 8'h01;
  assign sel_977254 = array_index_977233 == array_index_948511 ? add_977253 : sel_977250;
  assign add_977257 = sel_977254 + 8'h01;
  assign sel_977258 = array_index_977233 == array_index_948519 ? add_977257 : sel_977254;
  assign add_977261 = sel_977258 + 8'h01;
  assign sel_977262 = array_index_977233 == array_index_948527 ? add_977261 : sel_977258;
  assign add_977265 = sel_977262 + 8'h01;
  assign sel_977266 = array_index_977233 == array_index_948535 ? add_977265 : sel_977262;
  assign add_977269 = sel_977266 + 8'h01;
  assign sel_977270 = array_index_977233 == array_index_948541 ? add_977269 : sel_977266;
  assign add_977273 = sel_977270 + 8'h01;
  assign sel_977274 = array_index_977233 == array_index_948547 ? add_977273 : sel_977270;
  assign add_977277 = sel_977274 + 8'h01;
  assign sel_977278 = array_index_977233 == array_index_948553 ? add_977277 : sel_977274;
  assign add_977281 = sel_977278 + 8'h01;
  assign sel_977282 = array_index_977233 == array_index_948559 ? add_977281 : sel_977278;
  assign add_977285 = sel_977282 + 8'h01;
  assign sel_977286 = array_index_977233 == array_index_948565 ? add_977285 : sel_977282;
  assign add_977289 = sel_977286 + 8'h01;
  assign sel_977290 = array_index_977233 == array_index_948571 ? add_977289 : sel_977286;
  assign add_977293 = sel_977290 + 8'h01;
  assign sel_977294 = array_index_977233 == array_index_948577 ? add_977293 : sel_977290;
  assign add_977297 = sel_977294 + 8'h01;
  assign sel_977298 = array_index_977233 == array_index_948583 ? add_977297 : sel_977294;
  assign add_977301 = sel_977298 + 8'h01;
  assign sel_977302 = array_index_977233 == array_index_948589 ? add_977301 : sel_977298;
  assign add_977305 = sel_977302 + 8'h01;
  assign sel_977306 = array_index_977233 == array_index_948595 ? add_977305 : sel_977302;
  assign add_977309 = sel_977306 + 8'h01;
  assign sel_977310 = array_index_977233 == array_index_948601 ? add_977309 : sel_977306;
  assign add_977313 = sel_977310 + 8'h01;
  assign sel_977314 = array_index_977233 == array_index_948607 ? add_977313 : sel_977310;
  assign add_977317 = sel_977314 + 8'h01;
  assign sel_977318 = array_index_977233 == array_index_948613 ? add_977317 : sel_977314;
  assign add_977321 = sel_977318 + 8'h01;
  assign sel_977322 = array_index_977233 == array_index_948619 ? add_977321 : sel_977318;
  assign add_977325 = sel_977322 + 8'h01;
  assign sel_977326 = array_index_977233 == array_index_948625 ? add_977325 : sel_977322;
  assign add_977329 = sel_977326 + 8'h01;
  assign sel_977330 = array_index_977233 == array_index_948631 ? add_977329 : sel_977326;
  assign add_977333 = sel_977330 + 8'h01;
  assign sel_977334 = array_index_977233 == array_index_948637 ? add_977333 : sel_977330;
  assign add_977337 = sel_977334 + 8'h01;
  assign sel_977338 = array_index_977233 == array_index_948643 ? add_977337 : sel_977334;
  assign add_977341 = sel_977338 + 8'h01;
  assign sel_977342 = array_index_977233 == array_index_948649 ? add_977341 : sel_977338;
  assign add_977345 = sel_977342 + 8'h01;
  assign sel_977346 = array_index_977233 == array_index_948655 ? add_977345 : sel_977342;
  assign add_977349 = sel_977346 + 8'h01;
  assign sel_977350 = array_index_977233 == array_index_948661 ? add_977349 : sel_977346;
  assign add_977353 = sel_977350 + 8'h01;
  assign sel_977354 = array_index_977233 == array_index_948667 ? add_977353 : sel_977350;
  assign add_977357 = sel_977354 + 8'h01;
  assign sel_977358 = array_index_977233 == array_index_948673 ? add_977357 : sel_977354;
  assign add_977361 = sel_977358 + 8'h01;
  assign sel_977362 = array_index_977233 == array_index_948679 ? add_977361 : sel_977358;
  assign add_977365 = sel_977362 + 8'h01;
  assign sel_977366 = array_index_977233 == array_index_948685 ? add_977365 : sel_977362;
  assign add_977369 = sel_977366 + 8'h01;
  assign sel_977370 = array_index_977233 == array_index_948691 ? add_977369 : sel_977366;
  assign add_977373 = sel_977370 + 8'h01;
  assign sel_977374 = array_index_977233 == array_index_948697 ? add_977373 : sel_977370;
  assign add_977377 = sel_977374 + 8'h01;
  assign sel_977378 = array_index_977233 == array_index_948703 ? add_977377 : sel_977374;
  assign add_977381 = sel_977378 + 8'h01;
  assign sel_977382 = array_index_977233 == array_index_948709 ? add_977381 : sel_977378;
  assign add_977385 = sel_977382 + 8'h01;
  assign sel_977386 = array_index_977233 == array_index_948715 ? add_977385 : sel_977382;
  assign add_977389 = sel_977386 + 8'h01;
  assign sel_977390 = array_index_977233 == array_index_948721 ? add_977389 : sel_977386;
  assign add_977393 = sel_977390 + 8'h01;
  assign sel_977394 = array_index_977233 == array_index_948727 ? add_977393 : sel_977390;
  assign add_977397 = sel_977394 + 8'h01;
  assign sel_977398 = array_index_977233 == array_index_948733 ? add_977397 : sel_977394;
  assign add_977401 = sel_977398 + 8'h01;
  assign sel_977402 = array_index_977233 == array_index_948739 ? add_977401 : sel_977398;
  assign add_977405 = sel_977402 + 8'h01;
  assign sel_977406 = array_index_977233 == array_index_948745 ? add_977405 : sel_977402;
  assign add_977409 = sel_977406 + 8'h01;
  assign sel_977410 = array_index_977233 == array_index_948751 ? add_977409 : sel_977406;
  assign add_977413 = sel_977410 + 8'h01;
  assign sel_977414 = array_index_977233 == array_index_948757 ? add_977413 : sel_977410;
  assign add_977417 = sel_977414 + 8'h01;
  assign sel_977418 = array_index_977233 == array_index_948763 ? add_977417 : sel_977414;
  assign add_977421 = sel_977418 + 8'h01;
  assign sel_977422 = array_index_977233 == array_index_948769 ? add_977421 : sel_977418;
  assign add_977425 = sel_977422 + 8'h01;
  assign sel_977426 = array_index_977233 == array_index_948775 ? add_977425 : sel_977422;
  assign add_977429 = sel_977426 + 8'h01;
  assign sel_977430 = array_index_977233 == array_index_948781 ? add_977429 : sel_977426;
  assign add_977433 = sel_977430 + 8'h01;
  assign sel_977434 = array_index_977233 == array_index_948787 ? add_977433 : sel_977430;
  assign add_977437 = sel_977434 + 8'h01;
  assign sel_977438 = array_index_977233 == array_index_948793 ? add_977437 : sel_977434;
  assign add_977441 = sel_977438 + 8'h01;
  assign sel_977442 = array_index_977233 == array_index_948799 ? add_977441 : sel_977438;
  assign add_977445 = sel_977442 + 8'h01;
  assign sel_977446 = array_index_977233 == array_index_948805 ? add_977445 : sel_977442;
  assign add_977449 = sel_977446 + 8'h01;
  assign sel_977450 = array_index_977233 == array_index_948811 ? add_977449 : sel_977446;
  assign add_977453 = sel_977450 + 8'h01;
  assign sel_977454 = array_index_977233 == array_index_948817 ? add_977453 : sel_977450;
  assign add_977457 = sel_977454 + 8'h01;
  assign sel_977458 = array_index_977233 == array_index_948823 ? add_977457 : sel_977454;
  assign add_977461 = sel_977458 + 8'h01;
  assign sel_977462 = array_index_977233 == array_index_948829 ? add_977461 : sel_977458;
  assign add_977465 = sel_977462 + 8'h01;
  assign sel_977466 = array_index_977233 == array_index_948835 ? add_977465 : sel_977462;
  assign add_977469 = sel_977466 + 8'h01;
  assign sel_977470 = array_index_977233 == array_index_948841 ? add_977469 : sel_977466;
  assign add_977473 = sel_977470 + 8'h01;
  assign sel_977474 = array_index_977233 == array_index_948847 ? add_977473 : sel_977470;
  assign add_977477 = sel_977474 + 8'h01;
  assign sel_977478 = array_index_977233 == array_index_948853 ? add_977477 : sel_977474;
  assign add_977481 = sel_977478 + 8'h01;
  assign sel_977482 = array_index_977233 == array_index_948859 ? add_977481 : sel_977478;
  assign add_977485 = sel_977482 + 8'h01;
  assign sel_977486 = array_index_977233 == array_index_948865 ? add_977485 : sel_977482;
  assign add_977489 = sel_977486 + 8'h01;
  assign sel_977490 = array_index_977233 == array_index_948871 ? add_977489 : sel_977486;
  assign add_977493 = sel_977490 + 8'h01;
  assign sel_977494 = array_index_977233 == array_index_948877 ? add_977493 : sel_977490;
  assign add_977497 = sel_977494 + 8'h01;
  assign sel_977498 = array_index_977233 == array_index_948883 ? add_977497 : sel_977494;
  assign add_977501 = sel_977498 + 8'h01;
  assign sel_977502 = array_index_977233 == array_index_948889 ? add_977501 : sel_977498;
  assign add_977505 = sel_977502 + 8'h01;
  assign sel_977506 = array_index_977233 == array_index_948895 ? add_977505 : sel_977502;
  assign add_977509 = sel_977506 + 8'h01;
  assign sel_977510 = array_index_977233 == array_index_948901 ? add_977509 : sel_977506;
  assign add_977513 = sel_977510 + 8'h01;
  assign sel_977514 = array_index_977233 == array_index_948907 ? add_977513 : sel_977510;
  assign add_977517 = sel_977514 + 8'h01;
  assign sel_977518 = array_index_977233 == array_index_948913 ? add_977517 : sel_977514;
  assign add_977521 = sel_977518 + 8'h01;
  assign sel_977522 = array_index_977233 == array_index_948919 ? add_977521 : sel_977518;
  assign add_977525 = sel_977522 + 8'h01;
  assign sel_977526 = array_index_977233 == array_index_948925 ? add_977525 : sel_977522;
  assign add_977529 = sel_977526 + 8'h01;
  assign sel_977530 = array_index_977233 == array_index_948931 ? add_977529 : sel_977526;
  assign add_977533 = sel_977530 + 8'h01;
  assign sel_977534 = array_index_977233 == array_index_948937 ? add_977533 : sel_977530;
  assign add_977537 = sel_977534 + 8'h01;
  assign sel_977538 = array_index_977233 == array_index_948943 ? add_977537 : sel_977534;
  assign add_977541 = sel_977538 + 8'h01;
  assign sel_977542 = array_index_977233 == array_index_948949 ? add_977541 : sel_977538;
  assign add_977545 = sel_977542 + 8'h01;
  assign sel_977546 = array_index_977233 == array_index_948955 ? add_977545 : sel_977542;
  assign add_977549 = sel_977546 + 8'h01;
  assign sel_977550 = array_index_977233 == array_index_948961 ? add_977549 : sel_977546;
  assign add_977553 = sel_977550 + 8'h01;
  assign sel_977554 = array_index_977233 == array_index_948967 ? add_977553 : sel_977550;
  assign add_977557 = sel_977554 + 8'h01;
  assign sel_977558 = array_index_977233 == array_index_948973 ? add_977557 : sel_977554;
  assign add_977561 = sel_977558 + 8'h01;
  assign sel_977562 = array_index_977233 == array_index_948979 ? add_977561 : sel_977558;
  assign add_977565 = sel_977562 + 8'h01;
  assign sel_977566 = array_index_977233 == array_index_948985 ? add_977565 : sel_977562;
  assign add_977569 = sel_977566 + 8'h01;
  assign sel_977570 = array_index_977233 == array_index_948991 ? add_977569 : sel_977566;
  assign add_977573 = sel_977570 + 8'h01;
  assign sel_977574 = array_index_977233 == array_index_948997 ? add_977573 : sel_977570;
  assign add_977577 = sel_977574 + 8'h01;
  assign sel_977578 = array_index_977233 == array_index_949003 ? add_977577 : sel_977574;
  assign add_977581 = sel_977578 + 8'h01;
  assign sel_977582 = array_index_977233 == array_index_949009 ? add_977581 : sel_977578;
  assign add_977585 = sel_977582 + 8'h01;
  assign sel_977586 = array_index_977233 == array_index_949015 ? add_977585 : sel_977582;
  assign add_977589 = sel_977586 + 8'h01;
  assign sel_977590 = array_index_977233 == array_index_949021 ? add_977589 : sel_977586;
  assign add_977593 = sel_977590 + 8'h01;
  assign sel_977594 = array_index_977233 == array_index_949027 ? add_977593 : sel_977590;
  assign add_977597 = sel_977594 + 8'h01;
  assign sel_977598 = array_index_977233 == array_index_949033 ? add_977597 : sel_977594;
  assign add_977601 = sel_977598 + 8'h01;
  assign sel_977602 = array_index_977233 == array_index_949039 ? add_977601 : sel_977598;
  assign add_977605 = sel_977602 + 8'h01;
  assign sel_977606 = array_index_977233 == array_index_949045 ? add_977605 : sel_977602;
  assign add_977609 = sel_977606 + 8'h01;
  assign sel_977610 = array_index_977233 == array_index_949051 ? add_977609 : sel_977606;
  assign add_977613 = sel_977610 + 8'h01;
  assign sel_977614 = array_index_977233 == array_index_949057 ? add_977613 : sel_977610;
  assign add_977617 = sel_977614 + 8'h01;
  assign sel_977618 = array_index_977233 == array_index_949063 ? add_977617 : sel_977614;
  assign add_977621 = sel_977618 + 8'h01;
  assign sel_977622 = array_index_977233 == array_index_949069 ? add_977621 : sel_977618;
  assign add_977625 = sel_977622 + 8'h01;
  assign sel_977626 = array_index_977233 == array_index_949075 ? add_977625 : sel_977622;
  assign add_977629 = sel_977626 + 8'h01;
  assign sel_977630 = array_index_977233 == array_index_949081 ? add_977629 : sel_977626;
  assign add_977634 = sel_977630 + 8'h01;
  assign array_index_977635 = set1_unflattened[7'h48];
  assign sel_977636 = array_index_977233 == array_index_949087 ? add_977634 : sel_977630;
  assign add_977639 = sel_977636 + 8'h01;
  assign sel_977640 = array_index_977635 == array_index_948483 ? add_977639 : sel_977636;
  assign add_977643 = sel_977640 + 8'h01;
  assign sel_977644 = array_index_977635 == array_index_948487 ? add_977643 : sel_977640;
  assign add_977647 = sel_977644 + 8'h01;
  assign sel_977648 = array_index_977635 == array_index_948495 ? add_977647 : sel_977644;
  assign add_977651 = sel_977648 + 8'h01;
  assign sel_977652 = array_index_977635 == array_index_948503 ? add_977651 : sel_977648;
  assign add_977655 = sel_977652 + 8'h01;
  assign sel_977656 = array_index_977635 == array_index_948511 ? add_977655 : sel_977652;
  assign add_977659 = sel_977656 + 8'h01;
  assign sel_977660 = array_index_977635 == array_index_948519 ? add_977659 : sel_977656;
  assign add_977663 = sel_977660 + 8'h01;
  assign sel_977664 = array_index_977635 == array_index_948527 ? add_977663 : sel_977660;
  assign add_977667 = sel_977664 + 8'h01;
  assign sel_977668 = array_index_977635 == array_index_948535 ? add_977667 : sel_977664;
  assign add_977671 = sel_977668 + 8'h01;
  assign sel_977672 = array_index_977635 == array_index_948541 ? add_977671 : sel_977668;
  assign add_977675 = sel_977672 + 8'h01;
  assign sel_977676 = array_index_977635 == array_index_948547 ? add_977675 : sel_977672;
  assign add_977679 = sel_977676 + 8'h01;
  assign sel_977680 = array_index_977635 == array_index_948553 ? add_977679 : sel_977676;
  assign add_977683 = sel_977680 + 8'h01;
  assign sel_977684 = array_index_977635 == array_index_948559 ? add_977683 : sel_977680;
  assign add_977687 = sel_977684 + 8'h01;
  assign sel_977688 = array_index_977635 == array_index_948565 ? add_977687 : sel_977684;
  assign add_977691 = sel_977688 + 8'h01;
  assign sel_977692 = array_index_977635 == array_index_948571 ? add_977691 : sel_977688;
  assign add_977695 = sel_977692 + 8'h01;
  assign sel_977696 = array_index_977635 == array_index_948577 ? add_977695 : sel_977692;
  assign add_977699 = sel_977696 + 8'h01;
  assign sel_977700 = array_index_977635 == array_index_948583 ? add_977699 : sel_977696;
  assign add_977703 = sel_977700 + 8'h01;
  assign sel_977704 = array_index_977635 == array_index_948589 ? add_977703 : sel_977700;
  assign add_977707 = sel_977704 + 8'h01;
  assign sel_977708 = array_index_977635 == array_index_948595 ? add_977707 : sel_977704;
  assign add_977711 = sel_977708 + 8'h01;
  assign sel_977712 = array_index_977635 == array_index_948601 ? add_977711 : sel_977708;
  assign add_977715 = sel_977712 + 8'h01;
  assign sel_977716 = array_index_977635 == array_index_948607 ? add_977715 : sel_977712;
  assign add_977719 = sel_977716 + 8'h01;
  assign sel_977720 = array_index_977635 == array_index_948613 ? add_977719 : sel_977716;
  assign add_977723 = sel_977720 + 8'h01;
  assign sel_977724 = array_index_977635 == array_index_948619 ? add_977723 : sel_977720;
  assign add_977727 = sel_977724 + 8'h01;
  assign sel_977728 = array_index_977635 == array_index_948625 ? add_977727 : sel_977724;
  assign add_977731 = sel_977728 + 8'h01;
  assign sel_977732 = array_index_977635 == array_index_948631 ? add_977731 : sel_977728;
  assign add_977735 = sel_977732 + 8'h01;
  assign sel_977736 = array_index_977635 == array_index_948637 ? add_977735 : sel_977732;
  assign add_977739 = sel_977736 + 8'h01;
  assign sel_977740 = array_index_977635 == array_index_948643 ? add_977739 : sel_977736;
  assign add_977743 = sel_977740 + 8'h01;
  assign sel_977744 = array_index_977635 == array_index_948649 ? add_977743 : sel_977740;
  assign add_977747 = sel_977744 + 8'h01;
  assign sel_977748 = array_index_977635 == array_index_948655 ? add_977747 : sel_977744;
  assign add_977751 = sel_977748 + 8'h01;
  assign sel_977752 = array_index_977635 == array_index_948661 ? add_977751 : sel_977748;
  assign add_977755 = sel_977752 + 8'h01;
  assign sel_977756 = array_index_977635 == array_index_948667 ? add_977755 : sel_977752;
  assign add_977759 = sel_977756 + 8'h01;
  assign sel_977760 = array_index_977635 == array_index_948673 ? add_977759 : sel_977756;
  assign add_977763 = sel_977760 + 8'h01;
  assign sel_977764 = array_index_977635 == array_index_948679 ? add_977763 : sel_977760;
  assign add_977767 = sel_977764 + 8'h01;
  assign sel_977768 = array_index_977635 == array_index_948685 ? add_977767 : sel_977764;
  assign add_977771 = sel_977768 + 8'h01;
  assign sel_977772 = array_index_977635 == array_index_948691 ? add_977771 : sel_977768;
  assign add_977775 = sel_977772 + 8'h01;
  assign sel_977776 = array_index_977635 == array_index_948697 ? add_977775 : sel_977772;
  assign add_977779 = sel_977776 + 8'h01;
  assign sel_977780 = array_index_977635 == array_index_948703 ? add_977779 : sel_977776;
  assign add_977783 = sel_977780 + 8'h01;
  assign sel_977784 = array_index_977635 == array_index_948709 ? add_977783 : sel_977780;
  assign add_977787 = sel_977784 + 8'h01;
  assign sel_977788 = array_index_977635 == array_index_948715 ? add_977787 : sel_977784;
  assign add_977791 = sel_977788 + 8'h01;
  assign sel_977792 = array_index_977635 == array_index_948721 ? add_977791 : sel_977788;
  assign add_977795 = sel_977792 + 8'h01;
  assign sel_977796 = array_index_977635 == array_index_948727 ? add_977795 : sel_977792;
  assign add_977799 = sel_977796 + 8'h01;
  assign sel_977800 = array_index_977635 == array_index_948733 ? add_977799 : sel_977796;
  assign add_977803 = sel_977800 + 8'h01;
  assign sel_977804 = array_index_977635 == array_index_948739 ? add_977803 : sel_977800;
  assign add_977807 = sel_977804 + 8'h01;
  assign sel_977808 = array_index_977635 == array_index_948745 ? add_977807 : sel_977804;
  assign add_977811 = sel_977808 + 8'h01;
  assign sel_977812 = array_index_977635 == array_index_948751 ? add_977811 : sel_977808;
  assign add_977815 = sel_977812 + 8'h01;
  assign sel_977816 = array_index_977635 == array_index_948757 ? add_977815 : sel_977812;
  assign add_977819 = sel_977816 + 8'h01;
  assign sel_977820 = array_index_977635 == array_index_948763 ? add_977819 : sel_977816;
  assign add_977823 = sel_977820 + 8'h01;
  assign sel_977824 = array_index_977635 == array_index_948769 ? add_977823 : sel_977820;
  assign add_977827 = sel_977824 + 8'h01;
  assign sel_977828 = array_index_977635 == array_index_948775 ? add_977827 : sel_977824;
  assign add_977831 = sel_977828 + 8'h01;
  assign sel_977832 = array_index_977635 == array_index_948781 ? add_977831 : sel_977828;
  assign add_977835 = sel_977832 + 8'h01;
  assign sel_977836 = array_index_977635 == array_index_948787 ? add_977835 : sel_977832;
  assign add_977839 = sel_977836 + 8'h01;
  assign sel_977840 = array_index_977635 == array_index_948793 ? add_977839 : sel_977836;
  assign add_977843 = sel_977840 + 8'h01;
  assign sel_977844 = array_index_977635 == array_index_948799 ? add_977843 : sel_977840;
  assign add_977847 = sel_977844 + 8'h01;
  assign sel_977848 = array_index_977635 == array_index_948805 ? add_977847 : sel_977844;
  assign add_977851 = sel_977848 + 8'h01;
  assign sel_977852 = array_index_977635 == array_index_948811 ? add_977851 : sel_977848;
  assign add_977855 = sel_977852 + 8'h01;
  assign sel_977856 = array_index_977635 == array_index_948817 ? add_977855 : sel_977852;
  assign add_977859 = sel_977856 + 8'h01;
  assign sel_977860 = array_index_977635 == array_index_948823 ? add_977859 : sel_977856;
  assign add_977863 = sel_977860 + 8'h01;
  assign sel_977864 = array_index_977635 == array_index_948829 ? add_977863 : sel_977860;
  assign add_977867 = sel_977864 + 8'h01;
  assign sel_977868 = array_index_977635 == array_index_948835 ? add_977867 : sel_977864;
  assign add_977871 = sel_977868 + 8'h01;
  assign sel_977872 = array_index_977635 == array_index_948841 ? add_977871 : sel_977868;
  assign add_977875 = sel_977872 + 8'h01;
  assign sel_977876 = array_index_977635 == array_index_948847 ? add_977875 : sel_977872;
  assign add_977879 = sel_977876 + 8'h01;
  assign sel_977880 = array_index_977635 == array_index_948853 ? add_977879 : sel_977876;
  assign add_977883 = sel_977880 + 8'h01;
  assign sel_977884 = array_index_977635 == array_index_948859 ? add_977883 : sel_977880;
  assign add_977887 = sel_977884 + 8'h01;
  assign sel_977888 = array_index_977635 == array_index_948865 ? add_977887 : sel_977884;
  assign add_977891 = sel_977888 + 8'h01;
  assign sel_977892 = array_index_977635 == array_index_948871 ? add_977891 : sel_977888;
  assign add_977895 = sel_977892 + 8'h01;
  assign sel_977896 = array_index_977635 == array_index_948877 ? add_977895 : sel_977892;
  assign add_977899 = sel_977896 + 8'h01;
  assign sel_977900 = array_index_977635 == array_index_948883 ? add_977899 : sel_977896;
  assign add_977903 = sel_977900 + 8'h01;
  assign sel_977904 = array_index_977635 == array_index_948889 ? add_977903 : sel_977900;
  assign add_977907 = sel_977904 + 8'h01;
  assign sel_977908 = array_index_977635 == array_index_948895 ? add_977907 : sel_977904;
  assign add_977911 = sel_977908 + 8'h01;
  assign sel_977912 = array_index_977635 == array_index_948901 ? add_977911 : sel_977908;
  assign add_977915 = sel_977912 + 8'h01;
  assign sel_977916 = array_index_977635 == array_index_948907 ? add_977915 : sel_977912;
  assign add_977919 = sel_977916 + 8'h01;
  assign sel_977920 = array_index_977635 == array_index_948913 ? add_977919 : sel_977916;
  assign add_977923 = sel_977920 + 8'h01;
  assign sel_977924 = array_index_977635 == array_index_948919 ? add_977923 : sel_977920;
  assign add_977927 = sel_977924 + 8'h01;
  assign sel_977928 = array_index_977635 == array_index_948925 ? add_977927 : sel_977924;
  assign add_977931 = sel_977928 + 8'h01;
  assign sel_977932 = array_index_977635 == array_index_948931 ? add_977931 : sel_977928;
  assign add_977935 = sel_977932 + 8'h01;
  assign sel_977936 = array_index_977635 == array_index_948937 ? add_977935 : sel_977932;
  assign add_977939 = sel_977936 + 8'h01;
  assign sel_977940 = array_index_977635 == array_index_948943 ? add_977939 : sel_977936;
  assign add_977943 = sel_977940 + 8'h01;
  assign sel_977944 = array_index_977635 == array_index_948949 ? add_977943 : sel_977940;
  assign add_977947 = sel_977944 + 8'h01;
  assign sel_977948 = array_index_977635 == array_index_948955 ? add_977947 : sel_977944;
  assign add_977951 = sel_977948 + 8'h01;
  assign sel_977952 = array_index_977635 == array_index_948961 ? add_977951 : sel_977948;
  assign add_977955 = sel_977952 + 8'h01;
  assign sel_977956 = array_index_977635 == array_index_948967 ? add_977955 : sel_977952;
  assign add_977959 = sel_977956 + 8'h01;
  assign sel_977960 = array_index_977635 == array_index_948973 ? add_977959 : sel_977956;
  assign add_977963 = sel_977960 + 8'h01;
  assign sel_977964 = array_index_977635 == array_index_948979 ? add_977963 : sel_977960;
  assign add_977967 = sel_977964 + 8'h01;
  assign sel_977968 = array_index_977635 == array_index_948985 ? add_977967 : sel_977964;
  assign add_977971 = sel_977968 + 8'h01;
  assign sel_977972 = array_index_977635 == array_index_948991 ? add_977971 : sel_977968;
  assign add_977975 = sel_977972 + 8'h01;
  assign sel_977976 = array_index_977635 == array_index_948997 ? add_977975 : sel_977972;
  assign add_977979 = sel_977976 + 8'h01;
  assign sel_977980 = array_index_977635 == array_index_949003 ? add_977979 : sel_977976;
  assign add_977983 = sel_977980 + 8'h01;
  assign sel_977984 = array_index_977635 == array_index_949009 ? add_977983 : sel_977980;
  assign add_977987 = sel_977984 + 8'h01;
  assign sel_977988 = array_index_977635 == array_index_949015 ? add_977987 : sel_977984;
  assign add_977991 = sel_977988 + 8'h01;
  assign sel_977992 = array_index_977635 == array_index_949021 ? add_977991 : sel_977988;
  assign add_977995 = sel_977992 + 8'h01;
  assign sel_977996 = array_index_977635 == array_index_949027 ? add_977995 : sel_977992;
  assign add_977999 = sel_977996 + 8'h01;
  assign sel_978000 = array_index_977635 == array_index_949033 ? add_977999 : sel_977996;
  assign add_978003 = sel_978000 + 8'h01;
  assign sel_978004 = array_index_977635 == array_index_949039 ? add_978003 : sel_978000;
  assign add_978007 = sel_978004 + 8'h01;
  assign sel_978008 = array_index_977635 == array_index_949045 ? add_978007 : sel_978004;
  assign add_978011 = sel_978008 + 8'h01;
  assign sel_978012 = array_index_977635 == array_index_949051 ? add_978011 : sel_978008;
  assign add_978015 = sel_978012 + 8'h01;
  assign sel_978016 = array_index_977635 == array_index_949057 ? add_978015 : sel_978012;
  assign add_978019 = sel_978016 + 8'h01;
  assign sel_978020 = array_index_977635 == array_index_949063 ? add_978019 : sel_978016;
  assign add_978023 = sel_978020 + 8'h01;
  assign sel_978024 = array_index_977635 == array_index_949069 ? add_978023 : sel_978020;
  assign add_978027 = sel_978024 + 8'h01;
  assign sel_978028 = array_index_977635 == array_index_949075 ? add_978027 : sel_978024;
  assign add_978031 = sel_978028 + 8'h01;
  assign sel_978032 = array_index_977635 == array_index_949081 ? add_978031 : sel_978028;
  assign add_978036 = sel_978032 + 8'h01;
  assign array_index_978037 = set1_unflattened[7'h49];
  assign sel_978038 = array_index_977635 == array_index_949087 ? add_978036 : sel_978032;
  assign add_978041 = sel_978038 + 8'h01;
  assign sel_978042 = array_index_978037 == array_index_948483 ? add_978041 : sel_978038;
  assign add_978045 = sel_978042 + 8'h01;
  assign sel_978046 = array_index_978037 == array_index_948487 ? add_978045 : sel_978042;
  assign add_978049 = sel_978046 + 8'h01;
  assign sel_978050 = array_index_978037 == array_index_948495 ? add_978049 : sel_978046;
  assign add_978053 = sel_978050 + 8'h01;
  assign sel_978054 = array_index_978037 == array_index_948503 ? add_978053 : sel_978050;
  assign add_978057 = sel_978054 + 8'h01;
  assign sel_978058 = array_index_978037 == array_index_948511 ? add_978057 : sel_978054;
  assign add_978061 = sel_978058 + 8'h01;
  assign sel_978062 = array_index_978037 == array_index_948519 ? add_978061 : sel_978058;
  assign add_978065 = sel_978062 + 8'h01;
  assign sel_978066 = array_index_978037 == array_index_948527 ? add_978065 : sel_978062;
  assign add_978069 = sel_978066 + 8'h01;
  assign sel_978070 = array_index_978037 == array_index_948535 ? add_978069 : sel_978066;
  assign add_978073 = sel_978070 + 8'h01;
  assign sel_978074 = array_index_978037 == array_index_948541 ? add_978073 : sel_978070;
  assign add_978077 = sel_978074 + 8'h01;
  assign sel_978078 = array_index_978037 == array_index_948547 ? add_978077 : sel_978074;
  assign add_978081 = sel_978078 + 8'h01;
  assign sel_978082 = array_index_978037 == array_index_948553 ? add_978081 : sel_978078;
  assign add_978085 = sel_978082 + 8'h01;
  assign sel_978086 = array_index_978037 == array_index_948559 ? add_978085 : sel_978082;
  assign add_978089 = sel_978086 + 8'h01;
  assign sel_978090 = array_index_978037 == array_index_948565 ? add_978089 : sel_978086;
  assign add_978093 = sel_978090 + 8'h01;
  assign sel_978094 = array_index_978037 == array_index_948571 ? add_978093 : sel_978090;
  assign add_978097 = sel_978094 + 8'h01;
  assign sel_978098 = array_index_978037 == array_index_948577 ? add_978097 : sel_978094;
  assign add_978101 = sel_978098 + 8'h01;
  assign sel_978102 = array_index_978037 == array_index_948583 ? add_978101 : sel_978098;
  assign add_978105 = sel_978102 + 8'h01;
  assign sel_978106 = array_index_978037 == array_index_948589 ? add_978105 : sel_978102;
  assign add_978109 = sel_978106 + 8'h01;
  assign sel_978110 = array_index_978037 == array_index_948595 ? add_978109 : sel_978106;
  assign add_978113 = sel_978110 + 8'h01;
  assign sel_978114 = array_index_978037 == array_index_948601 ? add_978113 : sel_978110;
  assign add_978117 = sel_978114 + 8'h01;
  assign sel_978118 = array_index_978037 == array_index_948607 ? add_978117 : sel_978114;
  assign add_978121 = sel_978118 + 8'h01;
  assign sel_978122 = array_index_978037 == array_index_948613 ? add_978121 : sel_978118;
  assign add_978125 = sel_978122 + 8'h01;
  assign sel_978126 = array_index_978037 == array_index_948619 ? add_978125 : sel_978122;
  assign add_978129 = sel_978126 + 8'h01;
  assign sel_978130 = array_index_978037 == array_index_948625 ? add_978129 : sel_978126;
  assign add_978133 = sel_978130 + 8'h01;
  assign sel_978134 = array_index_978037 == array_index_948631 ? add_978133 : sel_978130;
  assign add_978137 = sel_978134 + 8'h01;
  assign sel_978138 = array_index_978037 == array_index_948637 ? add_978137 : sel_978134;
  assign add_978141 = sel_978138 + 8'h01;
  assign sel_978142 = array_index_978037 == array_index_948643 ? add_978141 : sel_978138;
  assign add_978145 = sel_978142 + 8'h01;
  assign sel_978146 = array_index_978037 == array_index_948649 ? add_978145 : sel_978142;
  assign add_978149 = sel_978146 + 8'h01;
  assign sel_978150 = array_index_978037 == array_index_948655 ? add_978149 : sel_978146;
  assign add_978153 = sel_978150 + 8'h01;
  assign sel_978154 = array_index_978037 == array_index_948661 ? add_978153 : sel_978150;
  assign add_978157 = sel_978154 + 8'h01;
  assign sel_978158 = array_index_978037 == array_index_948667 ? add_978157 : sel_978154;
  assign add_978161 = sel_978158 + 8'h01;
  assign sel_978162 = array_index_978037 == array_index_948673 ? add_978161 : sel_978158;
  assign add_978165 = sel_978162 + 8'h01;
  assign sel_978166 = array_index_978037 == array_index_948679 ? add_978165 : sel_978162;
  assign add_978169 = sel_978166 + 8'h01;
  assign sel_978170 = array_index_978037 == array_index_948685 ? add_978169 : sel_978166;
  assign add_978173 = sel_978170 + 8'h01;
  assign sel_978174 = array_index_978037 == array_index_948691 ? add_978173 : sel_978170;
  assign add_978177 = sel_978174 + 8'h01;
  assign sel_978178 = array_index_978037 == array_index_948697 ? add_978177 : sel_978174;
  assign add_978181 = sel_978178 + 8'h01;
  assign sel_978182 = array_index_978037 == array_index_948703 ? add_978181 : sel_978178;
  assign add_978185 = sel_978182 + 8'h01;
  assign sel_978186 = array_index_978037 == array_index_948709 ? add_978185 : sel_978182;
  assign add_978189 = sel_978186 + 8'h01;
  assign sel_978190 = array_index_978037 == array_index_948715 ? add_978189 : sel_978186;
  assign add_978193 = sel_978190 + 8'h01;
  assign sel_978194 = array_index_978037 == array_index_948721 ? add_978193 : sel_978190;
  assign add_978197 = sel_978194 + 8'h01;
  assign sel_978198 = array_index_978037 == array_index_948727 ? add_978197 : sel_978194;
  assign add_978201 = sel_978198 + 8'h01;
  assign sel_978202 = array_index_978037 == array_index_948733 ? add_978201 : sel_978198;
  assign add_978205 = sel_978202 + 8'h01;
  assign sel_978206 = array_index_978037 == array_index_948739 ? add_978205 : sel_978202;
  assign add_978209 = sel_978206 + 8'h01;
  assign sel_978210 = array_index_978037 == array_index_948745 ? add_978209 : sel_978206;
  assign add_978213 = sel_978210 + 8'h01;
  assign sel_978214 = array_index_978037 == array_index_948751 ? add_978213 : sel_978210;
  assign add_978217 = sel_978214 + 8'h01;
  assign sel_978218 = array_index_978037 == array_index_948757 ? add_978217 : sel_978214;
  assign add_978221 = sel_978218 + 8'h01;
  assign sel_978222 = array_index_978037 == array_index_948763 ? add_978221 : sel_978218;
  assign add_978225 = sel_978222 + 8'h01;
  assign sel_978226 = array_index_978037 == array_index_948769 ? add_978225 : sel_978222;
  assign add_978229 = sel_978226 + 8'h01;
  assign sel_978230 = array_index_978037 == array_index_948775 ? add_978229 : sel_978226;
  assign add_978233 = sel_978230 + 8'h01;
  assign sel_978234 = array_index_978037 == array_index_948781 ? add_978233 : sel_978230;
  assign add_978237 = sel_978234 + 8'h01;
  assign sel_978238 = array_index_978037 == array_index_948787 ? add_978237 : sel_978234;
  assign add_978241 = sel_978238 + 8'h01;
  assign sel_978242 = array_index_978037 == array_index_948793 ? add_978241 : sel_978238;
  assign add_978245 = sel_978242 + 8'h01;
  assign sel_978246 = array_index_978037 == array_index_948799 ? add_978245 : sel_978242;
  assign add_978249 = sel_978246 + 8'h01;
  assign sel_978250 = array_index_978037 == array_index_948805 ? add_978249 : sel_978246;
  assign add_978253 = sel_978250 + 8'h01;
  assign sel_978254 = array_index_978037 == array_index_948811 ? add_978253 : sel_978250;
  assign add_978257 = sel_978254 + 8'h01;
  assign sel_978258 = array_index_978037 == array_index_948817 ? add_978257 : sel_978254;
  assign add_978261 = sel_978258 + 8'h01;
  assign sel_978262 = array_index_978037 == array_index_948823 ? add_978261 : sel_978258;
  assign add_978265 = sel_978262 + 8'h01;
  assign sel_978266 = array_index_978037 == array_index_948829 ? add_978265 : sel_978262;
  assign add_978269 = sel_978266 + 8'h01;
  assign sel_978270 = array_index_978037 == array_index_948835 ? add_978269 : sel_978266;
  assign add_978273 = sel_978270 + 8'h01;
  assign sel_978274 = array_index_978037 == array_index_948841 ? add_978273 : sel_978270;
  assign add_978277 = sel_978274 + 8'h01;
  assign sel_978278 = array_index_978037 == array_index_948847 ? add_978277 : sel_978274;
  assign add_978281 = sel_978278 + 8'h01;
  assign sel_978282 = array_index_978037 == array_index_948853 ? add_978281 : sel_978278;
  assign add_978285 = sel_978282 + 8'h01;
  assign sel_978286 = array_index_978037 == array_index_948859 ? add_978285 : sel_978282;
  assign add_978289 = sel_978286 + 8'h01;
  assign sel_978290 = array_index_978037 == array_index_948865 ? add_978289 : sel_978286;
  assign add_978293 = sel_978290 + 8'h01;
  assign sel_978294 = array_index_978037 == array_index_948871 ? add_978293 : sel_978290;
  assign add_978297 = sel_978294 + 8'h01;
  assign sel_978298 = array_index_978037 == array_index_948877 ? add_978297 : sel_978294;
  assign add_978301 = sel_978298 + 8'h01;
  assign sel_978302 = array_index_978037 == array_index_948883 ? add_978301 : sel_978298;
  assign add_978305 = sel_978302 + 8'h01;
  assign sel_978306 = array_index_978037 == array_index_948889 ? add_978305 : sel_978302;
  assign add_978309 = sel_978306 + 8'h01;
  assign sel_978310 = array_index_978037 == array_index_948895 ? add_978309 : sel_978306;
  assign add_978313 = sel_978310 + 8'h01;
  assign sel_978314 = array_index_978037 == array_index_948901 ? add_978313 : sel_978310;
  assign add_978317 = sel_978314 + 8'h01;
  assign sel_978318 = array_index_978037 == array_index_948907 ? add_978317 : sel_978314;
  assign add_978321 = sel_978318 + 8'h01;
  assign sel_978322 = array_index_978037 == array_index_948913 ? add_978321 : sel_978318;
  assign add_978325 = sel_978322 + 8'h01;
  assign sel_978326 = array_index_978037 == array_index_948919 ? add_978325 : sel_978322;
  assign add_978329 = sel_978326 + 8'h01;
  assign sel_978330 = array_index_978037 == array_index_948925 ? add_978329 : sel_978326;
  assign add_978333 = sel_978330 + 8'h01;
  assign sel_978334 = array_index_978037 == array_index_948931 ? add_978333 : sel_978330;
  assign add_978337 = sel_978334 + 8'h01;
  assign sel_978338 = array_index_978037 == array_index_948937 ? add_978337 : sel_978334;
  assign add_978341 = sel_978338 + 8'h01;
  assign sel_978342 = array_index_978037 == array_index_948943 ? add_978341 : sel_978338;
  assign add_978345 = sel_978342 + 8'h01;
  assign sel_978346 = array_index_978037 == array_index_948949 ? add_978345 : sel_978342;
  assign add_978349 = sel_978346 + 8'h01;
  assign sel_978350 = array_index_978037 == array_index_948955 ? add_978349 : sel_978346;
  assign add_978353 = sel_978350 + 8'h01;
  assign sel_978354 = array_index_978037 == array_index_948961 ? add_978353 : sel_978350;
  assign add_978357 = sel_978354 + 8'h01;
  assign sel_978358 = array_index_978037 == array_index_948967 ? add_978357 : sel_978354;
  assign add_978361 = sel_978358 + 8'h01;
  assign sel_978362 = array_index_978037 == array_index_948973 ? add_978361 : sel_978358;
  assign add_978365 = sel_978362 + 8'h01;
  assign sel_978366 = array_index_978037 == array_index_948979 ? add_978365 : sel_978362;
  assign add_978369 = sel_978366 + 8'h01;
  assign sel_978370 = array_index_978037 == array_index_948985 ? add_978369 : sel_978366;
  assign add_978373 = sel_978370 + 8'h01;
  assign sel_978374 = array_index_978037 == array_index_948991 ? add_978373 : sel_978370;
  assign add_978377 = sel_978374 + 8'h01;
  assign sel_978378 = array_index_978037 == array_index_948997 ? add_978377 : sel_978374;
  assign add_978381 = sel_978378 + 8'h01;
  assign sel_978382 = array_index_978037 == array_index_949003 ? add_978381 : sel_978378;
  assign add_978385 = sel_978382 + 8'h01;
  assign sel_978386 = array_index_978037 == array_index_949009 ? add_978385 : sel_978382;
  assign add_978389 = sel_978386 + 8'h01;
  assign sel_978390 = array_index_978037 == array_index_949015 ? add_978389 : sel_978386;
  assign add_978393 = sel_978390 + 8'h01;
  assign sel_978394 = array_index_978037 == array_index_949021 ? add_978393 : sel_978390;
  assign add_978397 = sel_978394 + 8'h01;
  assign sel_978398 = array_index_978037 == array_index_949027 ? add_978397 : sel_978394;
  assign add_978401 = sel_978398 + 8'h01;
  assign sel_978402 = array_index_978037 == array_index_949033 ? add_978401 : sel_978398;
  assign add_978405 = sel_978402 + 8'h01;
  assign sel_978406 = array_index_978037 == array_index_949039 ? add_978405 : sel_978402;
  assign add_978409 = sel_978406 + 8'h01;
  assign sel_978410 = array_index_978037 == array_index_949045 ? add_978409 : sel_978406;
  assign add_978413 = sel_978410 + 8'h01;
  assign sel_978414 = array_index_978037 == array_index_949051 ? add_978413 : sel_978410;
  assign add_978417 = sel_978414 + 8'h01;
  assign sel_978418 = array_index_978037 == array_index_949057 ? add_978417 : sel_978414;
  assign add_978421 = sel_978418 + 8'h01;
  assign sel_978422 = array_index_978037 == array_index_949063 ? add_978421 : sel_978418;
  assign add_978425 = sel_978422 + 8'h01;
  assign sel_978426 = array_index_978037 == array_index_949069 ? add_978425 : sel_978422;
  assign add_978429 = sel_978426 + 8'h01;
  assign sel_978430 = array_index_978037 == array_index_949075 ? add_978429 : sel_978426;
  assign add_978433 = sel_978430 + 8'h01;
  assign sel_978434 = array_index_978037 == array_index_949081 ? add_978433 : sel_978430;
  assign add_978438 = sel_978434 + 8'h01;
  assign array_index_978439 = set1_unflattened[7'h4a];
  assign sel_978440 = array_index_978037 == array_index_949087 ? add_978438 : sel_978434;
  assign add_978443 = sel_978440 + 8'h01;
  assign sel_978444 = array_index_978439 == array_index_948483 ? add_978443 : sel_978440;
  assign add_978447 = sel_978444 + 8'h01;
  assign sel_978448 = array_index_978439 == array_index_948487 ? add_978447 : sel_978444;
  assign add_978451 = sel_978448 + 8'h01;
  assign sel_978452 = array_index_978439 == array_index_948495 ? add_978451 : sel_978448;
  assign add_978455 = sel_978452 + 8'h01;
  assign sel_978456 = array_index_978439 == array_index_948503 ? add_978455 : sel_978452;
  assign add_978459 = sel_978456 + 8'h01;
  assign sel_978460 = array_index_978439 == array_index_948511 ? add_978459 : sel_978456;
  assign add_978463 = sel_978460 + 8'h01;
  assign sel_978464 = array_index_978439 == array_index_948519 ? add_978463 : sel_978460;
  assign add_978467 = sel_978464 + 8'h01;
  assign sel_978468 = array_index_978439 == array_index_948527 ? add_978467 : sel_978464;
  assign add_978471 = sel_978468 + 8'h01;
  assign sel_978472 = array_index_978439 == array_index_948535 ? add_978471 : sel_978468;
  assign add_978475 = sel_978472 + 8'h01;
  assign sel_978476 = array_index_978439 == array_index_948541 ? add_978475 : sel_978472;
  assign add_978479 = sel_978476 + 8'h01;
  assign sel_978480 = array_index_978439 == array_index_948547 ? add_978479 : sel_978476;
  assign add_978483 = sel_978480 + 8'h01;
  assign sel_978484 = array_index_978439 == array_index_948553 ? add_978483 : sel_978480;
  assign add_978487 = sel_978484 + 8'h01;
  assign sel_978488 = array_index_978439 == array_index_948559 ? add_978487 : sel_978484;
  assign add_978491 = sel_978488 + 8'h01;
  assign sel_978492 = array_index_978439 == array_index_948565 ? add_978491 : sel_978488;
  assign add_978495 = sel_978492 + 8'h01;
  assign sel_978496 = array_index_978439 == array_index_948571 ? add_978495 : sel_978492;
  assign add_978499 = sel_978496 + 8'h01;
  assign sel_978500 = array_index_978439 == array_index_948577 ? add_978499 : sel_978496;
  assign add_978503 = sel_978500 + 8'h01;
  assign sel_978504 = array_index_978439 == array_index_948583 ? add_978503 : sel_978500;
  assign add_978507 = sel_978504 + 8'h01;
  assign sel_978508 = array_index_978439 == array_index_948589 ? add_978507 : sel_978504;
  assign add_978511 = sel_978508 + 8'h01;
  assign sel_978512 = array_index_978439 == array_index_948595 ? add_978511 : sel_978508;
  assign add_978515 = sel_978512 + 8'h01;
  assign sel_978516 = array_index_978439 == array_index_948601 ? add_978515 : sel_978512;
  assign add_978519 = sel_978516 + 8'h01;
  assign sel_978520 = array_index_978439 == array_index_948607 ? add_978519 : sel_978516;
  assign add_978523 = sel_978520 + 8'h01;
  assign sel_978524 = array_index_978439 == array_index_948613 ? add_978523 : sel_978520;
  assign add_978527 = sel_978524 + 8'h01;
  assign sel_978528 = array_index_978439 == array_index_948619 ? add_978527 : sel_978524;
  assign add_978531 = sel_978528 + 8'h01;
  assign sel_978532 = array_index_978439 == array_index_948625 ? add_978531 : sel_978528;
  assign add_978535 = sel_978532 + 8'h01;
  assign sel_978536 = array_index_978439 == array_index_948631 ? add_978535 : sel_978532;
  assign add_978539 = sel_978536 + 8'h01;
  assign sel_978540 = array_index_978439 == array_index_948637 ? add_978539 : sel_978536;
  assign add_978543 = sel_978540 + 8'h01;
  assign sel_978544 = array_index_978439 == array_index_948643 ? add_978543 : sel_978540;
  assign add_978547 = sel_978544 + 8'h01;
  assign sel_978548 = array_index_978439 == array_index_948649 ? add_978547 : sel_978544;
  assign add_978551 = sel_978548 + 8'h01;
  assign sel_978552 = array_index_978439 == array_index_948655 ? add_978551 : sel_978548;
  assign add_978555 = sel_978552 + 8'h01;
  assign sel_978556 = array_index_978439 == array_index_948661 ? add_978555 : sel_978552;
  assign add_978559 = sel_978556 + 8'h01;
  assign sel_978560 = array_index_978439 == array_index_948667 ? add_978559 : sel_978556;
  assign add_978563 = sel_978560 + 8'h01;
  assign sel_978564 = array_index_978439 == array_index_948673 ? add_978563 : sel_978560;
  assign add_978567 = sel_978564 + 8'h01;
  assign sel_978568 = array_index_978439 == array_index_948679 ? add_978567 : sel_978564;
  assign add_978571 = sel_978568 + 8'h01;
  assign sel_978572 = array_index_978439 == array_index_948685 ? add_978571 : sel_978568;
  assign add_978575 = sel_978572 + 8'h01;
  assign sel_978576 = array_index_978439 == array_index_948691 ? add_978575 : sel_978572;
  assign add_978579 = sel_978576 + 8'h01;
  assign sel_978580 = array_index_978439 == array_index_948697 ? add_978579 : sel_978576;
  assign add_978583 = sel_978580 + 8'h01;
  assign sel_978584 = array_index_978439 == array_index_948703 ? add_978583 : sel_978580;
  assign add_978587 = sel_978584 + 8'h01;
  assign sel_978588 = array_index_978439 == array_index_948709 ? add_978587 : sel_978584;
  assign add_978591 = sel_978588 + 8'h01;
  assign sel_978592 = array_index_978439 == array_index_948715 ? add_978591 : sel_978588;
  assign add_978595 = sel_978592 + 8'h01;
  assign sel_978596 = array_index_978439 == array_index_948721 ? add_978595 : sel_978592;
  assign add_978599 = sel_978596 + 8'h01;
  assign sel_978600 = array_index_978439 == array_index_948727 ? add_978599 : sel_978596;
  assign add_978603 = sel_978600 + 8'h01;
  assign sel_978604 = array_index_978439 == array_index_948733 ? add_978603 : sel_978600;
  assign add_978607 = sel_978604 + 8'h01;
  assign sel_978608 = array_index_978439 == array_index_948739 ? add_978607 : sel_978604;
  assign add_978611 = sel_978608 + 8'h01;
  assign sel_978612 = array_index_978439 == array_index_948745 ? add_978611 : sel_978608;
  assign add_978615 = sel_978612 + 8'h01;
  assign sel_978616 = array_index_978439 == array_index_948751 ? add_978615 : sel_978612;
  assign add_978619 = sel_978616 + 8'h01;
  assign sel_978620 = array_index_978439 == array_index_948757 ? add_978619 : sel_978616;
  assign add_978623 = sel_978620 + 8'h01;
  assign sel_978624 = array_index_978439 == array_index_948763 ? add_978623 : sel_978620;
  assign add_978627 = sel_978624 + 8'h01;
  assign sel_978628 = array_index_978439 == array_index_948769 ? add_978627 : sel_978624;
  assign add_978631 = sel_978628 + 8'h01;
  assign sel_978632 = array_index_978439 == array_index_948775 ? add_978631 : sel_978628;
  assign add_978635 = sel_978632 + 8'h01;
  assign sel_978636 = array_index_978439 == array_index_948781 ? add_978635 : sel_978632;
  assign add_978639 = sel_978636 + 8'h01;
  assign sel_978640 = array_index_978439 == array_index_948787 ? add_978639 : sel_978636;
  assign add_978643 = sel_978640 + 8'h01;
  assign sel_978644 = array_index_978439 == array_index_948793 ? add_978643 : sel_978640;
  assign add_978647 = sel_978644 + 8'h01;
  assign sel_978648 = array_index_978439 == array_index_948799 ? add_978647 : sel_978644;
  assign add_978651 = sel_978648 + 8'h01;
  assign sel_978652 = array_index_978439 == array_index_948805 ? add_978651 : sel_978648;
  assign add_978655 = sel_978652 + 8'h01;
  assign sel_978656 = array_index_978439 == array_index_948811 ? add_978655 : sel_978652;
  assign add_978659 = sel_978656 + 8'h01;
  assign sel_978660 = array_index_978439 == array_index_948817 ? add_978659 : sel_978656;
  assign add_978663 = sel_978660 + 8'h01;
  assign sel_978664 = array_index_978439 == array_index_948823 ? add_978663 : sel_978660;
  assign add_978667 = sel_978664 + 8'h01;
  assign sel_978668 = array_index_978439 == array_index_948829 ? add_978667 : sel_978664;
  assign add_978671 = sel_978668 + 8'h01;
  assign sel_978672 = array_index_978439 == array_index_948835 ? add_978671 : sel_978668;
  assign add_978675 = sel_978672 + 8'h01;
  assign sel_978676 = array_index_978439 == array_index_948841 ? add_978675 : sel_978672;
  assign add_978679 = sel_978676 + 8'h01;
  assign sel_978680 = array_index_978439 == array_index_948847 ? add_978679 : sel_978676;
  assign add_978683 = sel_978680 + 8'h01;
  assign sel_978684 = array_index_978439 == array_index_948853 ? add_978683 : sel_978680;
  assign add_978687 = sel_978684 + 8'h01;
  assign sel_978688 = array_index_978439 == array_index_948859 ? add_978687 : sel_978684;
  assign add_978691 = sel_978688 + 8'h01;
  assign sel_978692 = array_index_978439 == array_index_948865 ? add_978691 : sel_978688;
  assign add_978695 = sel_978692 + 8'h01;
  assign sel_978696 = array_index_978439 == array_index_948871 ? add_978695 : sel_978692;
  assign add_978699 = sel_978696 + 8'h01;
  assign sel_978700 = array_index_978439 == array_index_948877 ? add_978699 : sel_978696;
  assign add_978703 = sel_978700 + 8'h01;
  assign sel_978704 = array_index_978439 == array_index_948883 ? add_978703 : sel_978700;
  assign add_978707 = sel_978704 + 8'h01;
  assign sel_978708 = array_index_978439 == array_index_948889 ? add_978707 : sel_978704;
  assign add_978711 = sel_978708 + 8'h01;
  assign sel_978712 = array_index_978439 == array_index_948895 ? add_978711 : sel_978708;
  assign add_978715 = sel_978712 + 8'h01;
  assign sel_978716 = array_index_978439 == array_index_948901 ? add_978715 : sel_978712;
  assign add_978719 = sel_978716 + 8'h01;
  assign sel_978720 = array_index_978439 == array_index_948907 ? add_978719 : sel_978716;
  assign add_978723 = sel_978720 + 8'h01;
  assign sel_978724 = array_index_978439 == array_index_948913 ? add_978723 : sel_978720;
  assign add_978727 = sel_978724 + 8'h01;
  assign sel_978728 = array_index_978439 == array_index_948919 ? add_978727 : sel_978724;
  assign add_978731 = sel_978728 + 8'h01;
  assign sel_978732 = array_index_978439 == array_index_948925 ? add_978731 : sel_978728;
  assign add_978735 = sel_978732 + 8'h01;
  assign sel_978736 = array_index_978439 == array_index_948931 ? add_978735 : sel_978732;
  assign add_978739 = sel_978736 + 8'h01;
  assign sel_978740 = array_index_978439 == array_index_948937 ? add_978739 : sel_978736;
  assign add_978743 = sel_978740 + 8'h01;
  assign sel_978744 = array_index_978439 == array_index_948943 ? add_978743 : sel_978740;
  assign add_978747 = sel_978744 + 8'h01;
  assign sel_978748 = array_index_978439 == array_index_948949 ? add_978747 : sel_978744;
  assign add_978751 = sel_978748 + 8'h01;
  assign sel_978752 = array_index_978439 == array_index_948955 ? add_978751 : sel_978748;
  assign add_978755 = sel_978752 + 8'h01;
  assign sel_978756 = array_index_978439 == array_index_948961 ? add_978755 : sel_978752;
  assign add_978759 = sel_978756 + 8'h01;
  assign sel_978760 = array_index_978439 == array_index_948967 ? add_978759 : sel_978756;
  assign add_978763 = sel_978760 + 8'h01;
  assign sel_978764 = array_index_978439 == array_index_948973 ? add_978763 : sel_978760;
  assign add_978767 = sel_978764 + 8'h01;
  assign sel_978768 = array_index_978439 == array_index_948979 ? add_978767 : sel_978764;
  assign add_978771 = sel_978768 + 8'h01;
  assign sel_978772 = array_index_978439 == array_index_948985 ? add_978771 : sel_978768;
  assign add_978775 = sel_978772 + 8'h01;
  assign sel_978776 = array_index_978439 == array_index_948991 ? add_978775 : sel_978772;
  assign add_978779 = sel_978776 + 8'h01;
  assign sel_978780 = array_index_978439 == array_index_948997 ? add_978779 : sel_978776;
  assign add_978783 = sel_978780 + 8'h01;
  assign sel_978784 = array_index_978439 == array_index_949003 ? add_978783 : sel_978780;
  assign add_978787 = sel_978784 + 8'h01;
  assign sel_978788 = array_index_978439 == array_index_949009 ? add_978787 : sel_978784;
  assign add_978791 = sel_978788 + 8'h01;
  assign sel_978792 = array_index_978439 == array_index_949015 ? add_978791 : sel_978788;
  assign add_978795 = sel_978792 + 8'h01;
  assign sel_978796 = array_index_978439 == array_index_949021 ? add_978795 : sel_978792;
  assign add_978799 = sel_978796 + 8'h01;
  assign sel_978800 = array_index_978439 == array_index_949027 ? add_978799 : sel_978796;
  assign add_978803 = sel_978800 + 8'h01;
  assign sel_978804 = array_index_978439 == array_index_949033 ? add_978803 : sel_978800;
  assign add_978807 = sel_978804 + 8'h01;
  assign sel_978808 = array_index_978439 == array_index_949039 ? add_978807 : sel_978804;
  assign add_978811 = sel_978808 + 8'h01;
  assign sel_978812 = array_index_978439 == array_index_949045 ? add_978811 : sel_978808;
  assign add_978815 = sel_978812 + 8'h01;
  assign sel_978816 = array_index_978439 == array_index_949051 ? add_978815 : sel_978812;
  assign add_978819 = sel_978816 + 8'h01;
  assign sel_978820 = array_index_978439 == array_index_949057 ? add_978819 : sel_978816;
  assign add_978823 = sel_978820 + 8'h01;
  assign sel_978824 = array_index_978439 == array_index_949063 ? add_978823 : sel_978820;
  assign add_978827 = sel_978824 + 8'h01;
  assign sel_978828 = array_index_978439 == array_index_949069 ? add_978827 : sel_978824;
  assign add_978831 = sel_978828 + 8'h01;
  assign sel_978832 = array_index_978439 == array_index_949075 ? add_978831 : sel_978828;
  assign add_978835 = sel_978832 + 8'h01;
  assign sel_978836 = array_index_978439 == array_index_949081 ? add_978835 : sel_978832;
  assign add_978840 = sel_978836 + 8'h01;
  assign array_index_978841 = set1_unflattened[7'h4b];
  assign sel_978842 = array_index_978439 == array_index_949087 ? add_978840 : sel_978836;
  assign add_978845 = sel_978842 + 8'h01;
  assign sel_978846 = array_index_978841 == array_index_948483 ? add_978845 : sel_978842;
  assign add_978849 = sel_978846 + 8'h01;
  assign sel_978850 = array_index_978841 == array_index_948487 ? add_978849 : sel_978846;
  assign add_978853 = sel_978850 + 8'h01;
  assign sel_978854 = array_index_978841 == array_index_948495 ? add_978853 : sel_978850;
  assign add_978857 = sel_978854 + 8'h01;
  assign sel_978858 = array_index_978841 == array_index_948503 ? add_978857 : sel_978854;
  assign add_978861 = sel_978858 + 8'h01;
  assign sel_978862 = array_index_978841 == array_index_948511 ? add_978861 : sel_978858;
  assign add_978865 = sel_978862 + 8'h01;
  assign sel_978866 = array_index_978841 == array_index_948519 ? add_978865 : sel_978862;
  assign add_978869 = sel_978866 + 8'h01;
  assign sel_978870 = array_index_978841 == array_index_948527 ? add_978869 : sel_978866;
  assign add_978873 = sel_978870 + 8'h01;
  assign sel_978874 = array_index_978841 == array_index_948535 ? add_978873 : sel_978870;
  assign add_978877 = sel_978874 + 8'h01;
  assign sel_978878 = array_index_978841 == array_index_948541 ? add_978877 : sel_978874;
  assign add_978881 = sel_978878 + 8'h01;
  assign sel_978882 = array_index_978841 == array_index_948547 ? add_978881 : sel_978878;
  assign add_978885 = sel_978882 + 8'h01;
  assign sel_978886 = array_index_978841 == array_index_948553 ? add_978885 : sel_978882;
  assign add_978889 = sel_978886 + 8'h01;
  assign sel_978890 = array_index_978841 == array_index_948559 ? add_978889 : sel_978886;
  assign add_978893 = sel_978890 + 8'h01;
  assign sel_978894 = array_index_978841 == array_index_948565 ? add_978893 : sel_978890;
  assign add_978897 = sel_978894 + 8'h01;
  assign sel_978898 = array_index_978841 == array_index_948571 ? add_978897 : sel_978894;
  assign add_978901 = sel_978898 + 8'h01;
  assign sel_978902 = array_index_978841 == array_index_948577 ? add_978901 : sel_978898;
  assign add_978905 = sel_978902 + 8'h01;
  assign sel_978906 = array_index_978841 == array_index_948583 ? add_978905 : sel_978902;
  assign add_978909 = sel_978906 + 8'h01;
  assign sel_978910 = array_index_978841 == array_index_948589 ? add_978909 : sel_978906;
  assign add_978913 = sel_978910 + 8'h01;
  assign sel_978914 = array_index_978841 == array_index_948595 ? add_978913 : sel_978910;
  assign add_978917 = sel_978914 + 8'h01;
  assign sel_978918 = array_index_978841 == array_index_948601 ? add_978917 : sel_978914;
  assign add_978921 = sel_978918 + 8'h01;
  assign sel_978922 = array_index_978841 == array_index_948607 ? add_978921 : sel_978918;
  assign add_978925 = sel_978922 + 8'h01;
  assign sel_978926 = array_index_978841 == array_index_948613 ? add_978925 : sel_978922;
  assign add_978929 = sel_978926 + 8'h01;
  assign sel_978930 = array_index_978841 == array_index_948619 ? add_978929 : sel_978926;
  assign add_978933 = sel_978930 + 8'h01;
  assign sel_978934 = array_index_978841 == array_index_948625 ? add_978933 : sel_978930;
  assign add_978937 = sel_978934 + 8'h01;
  assign sel_978938 = array_index_978841 == array_index_948631 ? add_978937 : sel_978934;
  assign add_978941 = sel_978938 + 8'h01;
  assign sel_978942 = array_index_978841 == array_index_948637 ? add_978941 : sel_978938;
  assign add_978945 = sel_978942 + 8'h01;
  assign sel_978946 = array_index_978841 == array_index_948643 ? add_978945 : sel_978942;
  assign add_978949 = sel_978946 + 8'h01;
  assign sel_978950 = array_index_978841 == array_index_948649 ? add_978949 : sel_978946;
  assign add_978953 = sel_978950 + 8'h01;
  assign sel_978954 = array_index_978841 == array_index_948655 ? add_978953 : sel_978950;
  assign add_978957 = sel_978954 + 8'h01;
  assign sel_978958 = array_index_978841 == array_index_948661 ? add_978957 : sel_978954;
  assign add_978961 = sel_978958 + 8'h01;
  assign sel_978962 = array_index_978841 == array_index_948667 ? add_978961 : sel_978958;
  assign add_978965 = sel_978962 + 8'h01;
  assign sel_978966 = array_index_978841 == array_index_948673 ? add_978965 : sel_978962;
  assign add_978969 = sel_978966 + 8'h01;
  assign sel_978970 = array_index_978841 == array_index_948679 ? add_978969 : sel_978966;
  assign add_978973 = sel_978970 + 8'h01;
  assign sel_978974 = array_index_978841 == array_index_948685 ? add_978973 : sel_978970;
  assign add_978977 = sel_978974 + 8'h01;
  assign sel_978978 = array_index_978841 == array_index_948691 ? add_978977 : sel_978974;
  assign add_978981 = sel_978978 + 8'h01;
  assign sel_978982 = array_index_978841 == array_index_948697 ? add_978981 : sel_978978;
  assign add_978985 = sel_978982 + 8'h01;
  assign sel_978986 = array_index_978841 == array_index_948703 ? add_978985 : sel_978982;
  assign add_978989 = sel_978986 + 8'h01;
  assign sel_978990 = array_index_978841 == array_index_948709 ? add_978989 : sel_978986;
  assign add_978993 = sel_978990 + 8'h01;
  assign sel_978994 = array_index_978841 == array_index_948715 ? add_978993 : sel_978990;
  assign add_978997 = sel_978994 + 8'h01;
  assign sel_978998 = array_index_978841 == array_index_948721 ? add_978997 : sel_978994;
  assign add_979001 = sel_978998 + 8'h01;
  assign sel_979002 = array_index_978841 == array_index_948727 ? add_979001 : sel_978998;
  assign add_979005 = sel_979002 + 8'h01;
  assign sel_979006 = array_index_978841 == array_index_948733 ? add_979005 : sel_979002;
  assign add_979009 = sel_979006 + 8'h01;
  assign sel_979010 = array_index_978841 == array_index_948739 ? add_979009 : sel_979006;
  assign add_979013 = sel_979010 + 8'h01;
  assign sel_979014 = array_index_978841 == array_index_948745 ? add_979013 : sel_979010;
  assign add_979017 = sel_979014 + 8'h01;
  assign sel_979018 = array_index_978841 == array_index_948751 ? add_979017 : sel_979014;
  assign add_979021 = sel_979018 + 8'h01;
  assign sel_979022 = array_index_978841 == array_index_948757 ? add_979021 : sel_979018;
  assign add_979025 = sel_979022 + 8'h01;
  assign sel_979026 = array_index_978841 == array_index_948763 ? add_979025 : sel_979022;
  assign add_979029 = sel_979026 + 8'h01;
  assign sel_979030 = array_index_978841 == array_index_948769 ? add_979029 : sel_979026;
  assign add_979033 = sel_979030 + 8'h01;
  assign sel_979034 = array_index_978841 == array_index_948775 ? add_979033 : sel_979030;
  assign add_979037 = sel_979034 + 8'h01;
  assign sel_979038 = array_index_978841 == array_index_948781 ? add_979037 : sel_979034;
  assign add_979041 = sel_979038 + 8'h01;
  assign sel_979042 = array_index_978841 == array_index_948787 ? add_979041 : sel_979038;
  assign add_979045 = sel_979042 + 8'h01;
  assign sel_979046 = array_index_978841 == array_index_948793 ? add_979045 : sel_979042;
  assign add_979049 = sel_979046 + 8'h01;
  assign sel_979050 = array_index_978841 == array_index_948799 ? add_979049 : sel_979046;
  assign add_979053 = sel_979050 + 8'h01;
  assign sel_979054 = array_index_978841 == array_index_948805 ? add_979053 : sel_979050;
  assign add_979057 = sel_979054 + 8'h01;
  assign sel_979058 = array_index_978841 == array_index_948811 ? add_979057 : sel_979054;
  assign add_979061 = sel_979058 + 8'h01;
  assign sel_979062 = array_index_978841 == array_index_948817 ? add_979061 : sel_979058;
  assign add_979065 = sel_979062 + 8'h01;
  assign sel_979066 = array_index_978841 == array_index_948823 ? add_979065 : sel_979062;
  assign add_979069 = sel_979066 + 8'h01;
  assign sel_979070 = array_index_978841 == array_index_948829 ? add_979069 : sel_979066;
  assign add_979073 = sel_979070 + 8'h01;
  assign sel_979074 = array_index_978841 == array_index_948835 ? add_979073 : sel_979070;
  assign add_979077 = sel_979074 + 8'h01;
  assign sel_979078 = array_index_978841 == array_index_948841 ? add_979077 : sel_979074;
  assign add_979081 = sel_979078 + 8'h01;
  assign sel_979082 = array_index_978841 == array_index_948847 ? add_979081 : sel_979078;
  assign add_979085 = sel_979082 + 8'h01;
  assign sel_979086 = array_index_978841 == array_index_948853 ? add_979085 : sel_979082;
  assign add_979089 = sel_979086 + 8'h01;
  assign sel_979090 = array_index_978841 == array_index_948859 ? add_979089 : sel_979086;
  assign add_979093 = sel_979090 + 8'h01;
  assign sel_979094 = array_index_978841 == array_index_948865 ? add_979093 : sel_979090;
  assign add_979097 = sel_979094 + 8'h01;
  assign sel_979098 = array_index_978841 == array_index_948871 ? add_979097 : sel_979094;
  assign add_979101 = sel_979098 + 8'h01;
  assign sel_979102 = array_index_978841 == array_index_948877 ? add_979101 : sel_979098;
  assign add_979105 = sel_979102 + 8'h01;
  assign sel_979106 = array_index_978841 == array_index_948883 ? add_979105 : sel_979102;
  assign add_979109 = sel_979106 + 8'h01;
  assign sel_979110 = array_index_978841 == array_index_948889 ? add_979109 : sel_979106;
  assign add_979113 = sel_979110 + 8'h01;
  assign sel_979114 = array_index_978841 == array_index_948895 ? add_979113 : sel_979110;
  assign add_979117 = sel_979114 + 8'h01;
  assign sel_979118 = array_index_978841 == array_index_948901 ? add_979117 : sel_979114;
  assign add_979121 = sel_979118 + 8'h01;
  assign sel_979122 = array_index_978841 == array_index_948907 ? add_979121 : sel_979118;
  assign add_979125 = sel_979122 + 8'h01;
  assign sel_979126 = array_index_978841 == array_index_948913 ? add_979125 : sel_979122;
  assign add_979129 = sel_979126 + 8'h01;
  assign sel_979130 = array_index_978841 == array_index_948919 ? add_979129 : sel_979126;
  assign add_979133 = sel_979130 + 8'h01;
  assign sel_979134 = array_index_978841 == array_index_948925 ? add_979133 : sel_979130;
  assign add_979137 = sel_979134 + 8'h01;
  assign sel_979138 = array_index_978841 == array_index_948931 ? add_979137 : sel_979134;
  assign add_979141 = sel_979138 + 8'h01;
  assign sel_979142 = array_index_978841 == array_index_948937 ? add_979141 : sel_979138;
  assign add_979145 = sel_979142 + 8'h01;
  assign sel_979146 = array_index_978841 == array_index_948943 ? add_979145 : sel_979142;
  assign add_979149 = sel_979146 + 8'h01;
  assign sel_979150 = array_index_978841 == array_index_948949 ? add_979149 : sel_979146;
  assign add_979153 = sel_979150 + 8'h01;
  assign sel_979154 = array_index_978841 == array_index_948955 ? add_979153 : sel_979150;
  assign add_979157 = sel_979154 + 8'h01;
  assign sel_979158 = array_index_978841 == array_index_948961 ? add_979157 : sel_979154;
  assign add_979161 = sel_979158 + 8'h01;
  assign sel_979162 = array_index_978841 == array_index_948967 ? add_979161 : sel_979158;
  assign add_979165 = sel_979162 + 8'h01;
  assign sel_979166 = array_index_978841 == array_index_948973 ? add_979165 : sel_979162;
  assign add_979169 = sel_979166 + 8'h01;
  assign sel_979170 = array_index_978841 == array_index_948979 ? add_979169 : sel_979166;
  assign add_979173 = sel_979170 + 8'h01;
  assign sel_979174 = array_index_978841 == array_index_948985 ? add_979173 : sel_979170;
  assign add_979177 = sel_979174 + 8'h01;
  assign sel_979178 = array_index_978841 == array_index_948991 ? add_979177 : sel_979174;
  assign add_979181 = sel_979178 + 8'h01;
  assign sel_979182 = array_index_978841 == array_index_948997 ? add_979181 : sel_979178;
  assign add_979185 = sel_979182 + 8'h01;
  assign sel_979186 = array_index_978841 == array_index_949003 ? add_979185 : sel_979182;
  assign add_979189 = sel_979186 + 8'h01;
  assign sel_979190 = array_index_978841 == array_index_949009 ? add_979189 : sel_979186;
  assign add_979193 = sel_979190 + 8'h01;
  assign sel_979194 = array_index_978841 == array_index_949015 ? add_979193 : sel_979190;
  assign add_979197 = sel_979194 + 8'h01;
  assign sel_979198 = array_index_978841 == array_index_949021 ? add_979197 : sel_979194;
  assign add_979201 = sel_979198 + 8'h01;
  assign sel_979202 = array_index_978841 == array_index_949027 ? add_979201 : sel_979198;
  assign add_979205 = sel_979202 + 8'h01;
  assign sel_979206 = array_index_978841 == array_index_949033 ? add_979205 : sel_979202;
  assign add_979209 = sel_979206 + 8'h01;
  assign sel_979210 = array_index_978841 == array_index_949039 ? add_979209 : sel_979206;
  assign add_979213 = sel_979210 + 8'h01;
  assign sel_979214 = array_index_978841 == array_index_949045 ? add_979213 : sel_979210;
  assign add_979217 = sel_979214 + 8'h01;
  assign sel_979218 = array_index_978841 == array_index_949051 ? add_979217 : sel_979214;
  assign add_979221 = sel_979218 + 8'h01;
  assign sel_979222 = array_index_978841 == array_index_949057 ? add_979221 : sel_979218;
  assign add_979225 = sel_979222 + 8'h01;
  assign sel_979226 = array_index_978841 == array_index_949063 ? add_979225 : sel_979222;
  assign add_979229 = sel_979226 + 8'h01;
  assign sel_979230 = array_index_978841 == array_index_949069 ? add_979229 : sel_979226;
  assign add_979233 = sel_979230 + 8'h01;
  assign sel_979234 = array_index_978841 == array_index_949075 ? add_979233 : sel_979230;
  assign add_979237 = sel_979234 + 8'h01;
  assign sel_979238 = array_index_978841 == array_index_949081 ? add_979237 : sel_979234;
  assign add_979242 = sel_979238 + 8'h01;
  assign array_index_979243 = set1_unflattened[7'h4c];
  assign sel_979244 = array_index_978841 == array_index_949087 ? add_979242 : sel_979238;
  assign add_979247 = sel_979244 + 8'h01;
  assign sel_979248 = array_index_979243 == array_index_948483 ? add_979247 : sel_979244;
  assign add_979251 = sel_979248 + 8'h01;
  assign sel_979252 = array_index_979243 == array_index_948487 ? add_979251 : sel_979248;
  assign add_979255 = sel_979252 + 8'h01;
  assign sel_979256 = array_index_979243 == array_index_948495 ? add_979255 : sel_979252;
  assign add_979259 = sel_979256 + 8'h01;
  assign sel_979260 = array_index_979243 == array_index_948503 ? add_979259 : sel_979256;
  assign add_979263 = sel_979260 + 8'h01;
  assign sel_979264 = array_index_979243 == array_index_948511 ? add_979263 : sel_979260;
  assign add_979267 = sel_979264 + 8'h01;
  assign sel_979268 = array_index_979243 == array_index_948519 ? add_979267 : sel_979264;
  assign add_979271 = sel_979268 + 8'h01;
  assign sel_979272 = array_index_979243 == array_index_948527 ? add_979271 : sel_979268;
  assign add_979275 = sel_979272 + 8'h01;
  assign sel_979276 = array_index_979243 == array_index_948535 ? add_979275 : sel_979272;
  assign add_979279 = sel_979276 + 8'h01;
  assign sel_979280 = array_index_979243 == array_index_948541 ? add_979279 : sel_979276;
  assign add_979283 = sel_979280 + 8'h01;
  assign sel_979284 = array_index_979243 == array_index_948547 ? add_979283 : sel_979280;
  assign add_979287 = sel_979284 + 8'h01;
  assign sel_979288 = array_index_979243 == array_index_948553 ? add_979287 : sel_979284;
  assign add_979291 = sel_979288 + 8'h01;
  assign sel_979292 = array_index_979243 == array_index_948559 ? add_979291 : sel_979288;
  assign add_979295 = sel_979292 + 8'h01;
  assign sel_979296 = array_index_979243 == array_index_948565 ? add_979295 : sel_979292;
  assign add_979299 = sel_979296 + 8'h01;
  assign sel_979300 = array_index_979243 == array_index_948571 ? add_979299 : sel_979296;
  assign add_979303 = sel_979300 + 8'h01;
  assign sel_979304 = array_index_979243 == array_index_948577 ? add_979303 : sel_979300;
  assign add_979307 = sel_979304 + 8'h01;
  assign sel_979308 = array_index_979243 == array_index_948583 ? add_979307 : sel_979304;
  assign add_979311 = sel_979308 + 8'h01;
  assign sel_979312 = array_index_979243 == array_index_948589 ? add_979311 : sel_979308;
  assign add_979315 = sel_979312 + 8'h01;
  assign sel_979316 = array_index_979243 == array_index_948595 ? add_979315 : sel_979312;
  assign add_979319 = sel_979316 + 8'h01;
  assign sel_979320 = array_index_979243 == array_index_948601 ? add_979319 : sel_979316;
  assign add_979323 = sel_979320 + 8'h01;
  assign sel_979324 = array_index_979243 == array_index_948607 ? add_979323 : sel_979320;
  assign add_979327 = sel_979324 + 8'h01;
  assign sel_979328 = array_index_979243 == array_index_948613 ? add_979327 : sel_979324;
  assign add_979331 = sel_979328 + 8'h01;
  assign sel_979332 = array_index_979243 == array_index_948619 ? add_979331 : sel_979328;
  assign add_979335 = sel_979332 + 8'h01;
  assign sel_979336 = array_index_979243 == array_index_948625 ? add_979335 : sel_979332;
  assign add_979339 = sel_979336 + 8'h01;
  assign sel_979340 = array_index_979243 == array_index_948631 ? add_979339 : sel_979336;
  assign add_979343 = sel_979340 + 8'h01;
  assign sel_979344 = array_index_979243 == array_index_948637 ? add_979343 : sel_979340;
  assign add_979347 = sel_979344 + 8'h01;
  assign sel_979348 = array_index_979243 == array_index_948643 ? add_979347 : sel_979344;
  assign add_979351 = sel_979348 + 8'h01;
  assign sel_979352 = array_index_979243 == array_index_948649 ? add_979351 : sel_979348;
  assign add_979355 = sel_979352 + 8'h01;
  assign sel_979356 = array_index_979243 == array_index_948655 ? add_979355 : sel_979352;
  assign add_979359 = sel_979356 + 8'h01;
  assign sel_979360 = array_index_979243 == array_index_948661 ? add_979359 : sel_979356;
  assign add_979363 = sel_979360 + 8'h01;
  assign sel_979364 = array_index_979243 == array_index_948667 ? add_979363 : sel_979360;
  assign add_979367 = sel_979364 + 8'h01;
  assign sel_979368 = array_index_979243 == array_index_948673 ? add_979367 : sel_979364;
  assign add_979371 = sel_979368 + 8'h01;
  assign sel_979372 = array_index_979243 == array_index_948679 ? add_979371 : sel_979368;
  assign add_979375 = sel_979372 + 8'h01;
  assign sel_979376 = array_index_979243 == array_index_948685 ? add_979375 : sel_979372;
  assign add_979379 = sel_979376 + 8'h01;
  assign sel_979380 = array_index_979243 == array_index_948691 ? add_979379 : sel_979376;
  assign add_979383 = sel_979380 + 8'h01;
  assign sel_979384 = array_index_979243 == array_index_948697 ? add_979383 : sel_979380;
  assign add_979387 = sel_979384 + 8'h01;
  assign sel_979388 = array_index_979243 == array_index_948703 ? add_979387 : sel_979384;
  assign add_979391 = sel_979388 + 8'h01;
  assign sel_979392 = array_index_979243 == array_index_948709 ? add_979391 : sel_979388;
  assign add_979395 = sel_979392 + 8'h01;
  assign sel_979396 = array_index_979243 == array_index_948715 ? add_979395 : sel_979392;
  assign add_979399 = sel_979396 + 8'h01;
  assign sel_979400 = array_index_979243 == array_index_948721 ? add_979399 : sel_979396;
  assign add_979403 = sel_979400 + 8'h01;
  assign sel_979404 = array_index_979243 == array_index_948727 ? add_979403 : sel_979400;
  assign add_979407 = sel_979404 + 8'h01;
  assign sel_979408 = array_index_979243 == array_index_948733 ? add_979407 : sel_979404;
  assign add_979411 = sel_979408 + 8'h01;
  assign sel_979412 = array_index_979243 == array_index_948739 ? add_979411 : sel_979408;
  assign add_979415 = sel_979412 + 8'h01;
  assign sel_979416 = array_index_979243 == array_index_948745 ? add_979415 : sel_979412;
  assign add_979419 = sel_979416 + 8'h01;
  assign sel_979420 = array_index_979243 == array_index_948751 ? add_979419 : sel_979416;
  assign add_979423 = sel_979420 + 8'h01;
  assign sel_979424 = array_index_979243 == array_index_948757 ? add_979423 : sel_979420;
  assign add_979427 = sel_979424 + 8'h01;
  assign sel_979428 = array_index_979243 == array_index_948763 ? add_979427 : sel_979424;
  assign add_979431 = sel_979428 + 8'h01;
  assign sel_979432 = array_index_979243 == array_index_948769 ? add_979431 : sel_979428;
  assign add_979435 = sel_979432 + 8'h01;
  assign sel_979436 = array_index_979243 == array_index_948775 ? add_979435 : sel_979432;
  assign add_979439 = sel_979436 + 8'h01;
  assign sel_979440 = array_index_979243 == array_index_948781 ? add_979439 : sel_979436;
  assign add_979443 = sel_979440 + 8'h01;
  assign sel_979444 = array_index_979243 == array_index_948787 ? add_979443 : sel_979440;
  assign add_979447 = sel_979444 + 8'h01;
  assign sel_979448 = array_index_979243 == array_index_948793 ? add_979447 : sel_979444;
  assign add_979451 = sel_979448 + 8'h01;
  assign sel_979452 = array_index_979243 == array_index_948799 ? add_979451 : sel_979448;
  assign add_979455 = sel_979452 + 8'h01;
  assign sel_979456 = array_index_979243 == array_index_948805 ? add_979455 : sel_979452;
  assign add_979459 = sel_979456 + 8'h01;
  assign sel_979460 = array_index_979243 == array_index_948811 ? add_979459 : sel_979456;
  assign add_979463 = sel_979460 + 8'h01;
  assign sel_979464 = array_index_979243 == array_index_948817 ? add_979463 : sel_979460;
  assign add_979467 = sel_979464 + 8'h01;
  assign sel_979468 = array_index_979243 == array_index_948823 ? add_979467 : sel_979464;
  assign add_979471 = sel_979468 + 8'h01;
  assign sel_979472 = array_index_979243 == array_index_948829 ? add_979471 : sel_979468;
  assign add_979475 = sel_979472 + 8'h01;
  assign sel_979476 = array_index_979243 == array_index_948835 ? add_979475 : sel_979472;
  assign add_979479 = sel_979476 + 8'h01;
  assign sel_979480 = array_index_979243 == array_index_948841 ? add_979479 : sel_979476;
  assign add_979483 = sel_979480 + 8'h01;
  assign sel_979484 = array_index_979243 == array_index_948847 ? add_979483 : sel_979480;
  assign add_979487 = sel_979484 + 8'h01;
  assign sel_979488 = array_index_979243 == array_index_948853 ? add_979487 : sel_979484;
  assign add_979491 = sel_979488 + 8'h01;
  assign sel_979492 = array_index_979243 == array_index_948859 ? add_979491 : sel_979488;
  assign add_979495 = sel_979492 + 8'h01;
  assign sel_979496 = array_index_979243 == array_index_948865 ? add_979495 : sel_979492;
  assign add_979499 = sel_979496 + 8'h01;
  assign sel_979500 = array_index_979243 == array_index_948871 ? add_979499 : sel_979496;
  assign add_979503 = sel_979500 + 8'h01;
  assign sel_979504 = array_index_979243 == array_index_948877 ? add_979503 : sel_979500;
  assign add_979507 = sel_979504 + 8'h01;
  assign sel_979508 = array_index_979243 == array_index_948883 ? add_979507 : sel_979504;
  assign add_979511 = sel_979508 + 8'h01;
  assign sel_979512 = array_index_979243 == array_index_948889 ? add_979511 : sel_979508;
  assign add_979515 = sel_979512 + 8'h01;
  assign sel_979516 = array_index_979243 == array_index_948895 ? add_979515 : sel_979512;
  assign add_979519 = sel_979516 + 8'h01;
  assign sel_979520 = array_index_979243 == array_index_948901 ? add_979519 : sel_979516;
  assign add_979523 = sel_979520 + 8'h01;
  assign sel_979524 = array_index_979243 == array_index_948907 ? add_979523 : sel_979520;
  assign add_979527 = sel_979524 + 8'h01;
  assign sel_979528 = array_index_979243 == array_index_948913 ? add_979527 : sel_979524;
  assign add_979531 = sel_979528 + 8'h01;
  assign sel_979532 = array_index_979243 == array_index_948919 ? add_979531 : sel_979528;
  assign add_979535 = sel_979532 + 8'h01;
  assign sel_979536 = array_index_979243 == array_index_948925 ? add_979535 : sel_979532;
  assign add_979539 = sel_979536 + 8'h01;
  assign sel_979540 = array_index_979243 == array_index_948931 ? add_979539 : sel_979536;
  assign add_979543 = sel_979540 + 8'h01;
  assign sel_979544 = array_index_979243 == array_index_948937 ? add_979543 : sel_979540;
  assign add_979547 = sel_979544 + 8'h01;
  assign sel_979548 = array_index_979243 == array_index_948943 ? add_979547 : sel_979544;
  assign add_979551 = sel_979548 + 8'h01;
  assign sel_979552 = array_index_979243 == array_index_948949 ? add_979551 : sel_979548;
  assign add_979555 = sel_979552 + 8'h01;
  assign sel_979556 = array_index_979243 == array_index_948955 ? add_979555 : sel_979552;
  assign add_979559 = sel_979556 + 8'h01;
  assign sel_979560 = array_index_979243 == array_index_948961 ? add_979559 : sel_979556;
  assign add_979563 = sel_979560 + 8'h01;
  assign sel_979564 = array_index_979243 == array_index_948967 ? add_979563 : sel_979560;
  assign add_979567 = sel_979564 + 8'h01;
  assign sel_979568 = array_index_979243 == array_index_948973 ? add_979567 : sel_979564;
  assign add_979571 = sel_979568 + 8'h01;
  assign sel_979572 = array_index_979243 == array_index_948979 ? add_979571 : sel_979568;
  assign add_979575 = sel_979572 + 8'h01;
  assign sel_979576 = array_index_979243 == array_index_948985 ? add_979575 : sel_979572;
  assign add_979579 = sel_979576 + 8'h01;
  assign sel_979580 = array_index_979243 == array_index_948991 ? add_979579 : sel_979576;
  assign add_979583 = sel_979580 + 8'h01;
  assign sel_979584 = array_index_979243 == array_index_948997 ? add_979583 : sel_979580;
  assign add_979587 = sel_979584 + 8'h01;
  assign sel_979588 = array_index_979243 == array_index_949003 ? add_979587 : sel_979584;
  assign add_979591 = sel_979588 + 8'h01;
  assign sel_979592 = array_index_979243 == array_index_949009 ? add_979591 : sel_979588;
  assign add_979595 = sel_979592 + 8'h01;
  assign sel_979596 = array_index_979243 == array_index_949015 ? add_979595 : sel_979592;
  assign add_979599 = sel_979596 + 8'h01;
  assign sel_979600 = array_index_979243 == array_index_949021 ? add_979599 : sel_979596;
  assign add_979603 = sel_979600 + 8'h01;
  assign sel_979604 = array_index_979243 == array_index_949027 ? add_979603 : sel_979600;
  assign add_979607 = sel_979604 + 8'h01;
  assign sel_979608 = array_index_979243 == array_index_949033 ? add_979607 : sel_979604;
  assign add_979611 = sel_979608 + 8'h01;
  assign sel_979612 = array_index_979243 == array_index_949039 ? add_979611 : sel_979608;
  assign add_979615 = sel_979612 + 8'h01;
  assign sel_979616 = array_index_979243 == array_index_949045 ? add_979615 : sel_979612;
  assign add_979619 = sel_979616 + 8'h01;
  assign sel_979620 = array_index_979243 == array_index_949051 ? add_979619 : sel_979616;
  assign add_979623 = sel_979620 + 8'h01;
  assign sel_979624 = array_index_979243 == array_index_949057 ? add_979623 : sel_979620;
  assign add_979627 = sel_979624 + 8'h01;
  assign sel_979628 = array_index_979243 == array_index_949063 ? add_979627 : sel_979624;
  assign add_979631 = sel_979628 + 8'h01;
  assign sel_979632 = array_index_979243 == array_index_949069 ? add_979631 : sel_979628;
  assign add_979635 = sel_979632 + 8'h01;
  assign sel_979636 = array_index_979243 == array_index_949075 ? add_979635 : sel_979632;
  assign add_979639 = sel_979636 + 8'h01;
  assign sel_979640 = array_index_979243 == array_index_949081 ? add_979639 : sel_979636;
  assign add_979644 = sel_979640 + 8'h01;
  assign array_index_979645 = set1_unflattened[7'h4d];
  assign sel_979646 = array_index_979243 == array_index_949087 ? add_979644 : sel_979640;
  assign add_979649 = sel_979646 + 8'h01;
  assign sel_979650 = array_index_979645 == array_index_948483 ? add_979649 : sel_979646;
  assign add_979653 = sel_979650 + 8'h01;
  assign sel_979654 = array_index_979645 == array_index_948487 ? add_979653 : sel_979650;
  assign add_979657 = sel_979654 + 8'h01;
  assign sel_979658 = array_index_979645 == array_index_948495 ? add_979657 : sel_979654;
  assign add_979661 = sel_979658 + 8'h01;
  assign sel_979662 = array_index_979645 == array_index_948503 ? add_979661 : sel_979658;
  assign add_979665 = sel_979662 + 8'h01;
  assign sel_979666 = array_index_979645 == array_index_948511 ? add_979665 : sel_979662;
  assign add_979669 = sel_979666 + 8'h01;
  assign sel_979670 = array_index_979645 == array_index_948519 ? add_979669 : sel_979666;
  assign add_979673 = sel_979670 + 8'h01;
  assign sel_979674 = array_index_979645 == array_index_948527 ? add_979673 : sel_979670;
  assign add_979677 = sel_979674 + 8'h01;
  assign sel_979678 = array_index_979645 == array_index_948535 ? add_979677 : sel_979674;
  assign add_979681 = sel_979678 + 8'h01;
  assign sel_979682 = array_index_979645 == array_index_948541 ? add_979681 : sel_979678;
  assign add_979685 = sel_979682 + 8'h01;
  assign sel_979686 = array_index_979645 == array_index_948547 ? add_979685 : sel_979682;
  assign add_979689 = sel_979686 + 8'h01;
  assign sel_979690 = array_index_979645 == array_index_948553 ? add_979689 : sel_979686;
  assign add_979693 = sel_979690 + 8'h01;
  assign sel_979694 = array_index_979645 == array_index_948559 ? add_979693 : sel_979690;
  assign add_979697 = sel_979694 + 8'h01;
  assign sel_979698 = array_index_979645 == array_index_948565 ? add_979697 : sel_979694;
  assign add_979701 = sel_979698 + 8'h01;
  assign sel_979702 = array_index_979645 == array_index_948571 ? add_979701 : sel_979698;
  assign add_979705 = sel_979702 + 8'h01;
  assign sel_979706 = array_index_979645 == array_index_948577 ? add_979705 : sel_979702;
  assign add_979709 = sel_979706 + 8'h01;
  assign sel_979710 = array_index_979645 == array_index_948583 ? add_979709 : sel_979706;
  assign add_979713 = sel_979710 + 8'h01;
  assign sel_979714 = array_index_979645 == array_index_948589 ? add_979713 : sel_979710;
  assign add_979717 = sel_979714 + 8'h01;
  assign sel_979718 = array_index_979645 == array_index_948595 ? add_979717 : sel_979714;
  assign add_979721 = sel_979718 + 8'h01;
  assign sel_979722 = array_index_979645 == array_index_948601 ? add_979721 : sel_979718;
  assign add_979725 = sel_979722 + 8'h01;
  assign sel_979726 = array_index_979645 == array_index_948607 ? add_979725 : sel_979722;
  assign add_979729 = sel_979726 + 8'h01;
  assign sel_979730 = array_index_979645 == array_index_948613 ? add_979729 : sel_979726;
  assign add_979733 = sel_979730 + 8'h01;
  assign sel_979734 = array_index_979645 == array_index_948619 ? add_979733 : sel_979730;
  assign add_979737 = sel_979734 + 8'h01;
  assign sel_979738 = array_index_979645 == array_index_948625 ? add_979737 : sel_979734;
  assign add_979741 = sel_979738 + 8'h01;
  assign sel_979742 = array_index_979645 == array_index_948631 ? add_979741 : sel_979738;
  assign add_979745 = sel_979742 + 8'h01;
  assign sel_979746 = array_index_979645 == array_index_948637 ? add_979745 : sel_979742;
  assign add_979749 = sel_979746 + 8'h01;
  assign sel_979750 = array_index_979645 == array_index_948643 ? add_979749 : sel_979746;
  assign add_979753 = sel_979750 + 8'h01;
  assign sel_979754 = array_index_979645 == array_index_948649 ? add_979753 : sel_979750;
  assign add_979757 = sel_979754 + 8'h01;
  assign sel_979758 = array_index_979645 == array_index_948655 ? add_979757 : sel_979754;
  assign add_979761 = sel_979758 + 8'h01;
  assign sel_979762 = array_index_979645 == array_index_948661 ? add_979761 : sel_979758;
  assign add_979765 = sel_979762 + 8'h01;
  assign sel_979766 = array_index_979645 == array_index_948667 ? add_979765 : sel_979762;
  assign add_979769 = sel_979766 + 8'h01;
  assign sel_979770 = array_index_979645 == array_index_948673 ? add_979769 : sel_979766;
  assign add_979773 = sel_979770 + 8'h01;
  assign sel_979774 = array_index_979645 == array_index_948679 ? add_979773 : sel_979770;
  assign add_979777 = sel_979774 + 8'h01;
  assign sel_979778 = array_index_979645 == array_index_948685 ? add_979777 : sel_979774;
  assign add_979781 = sel_979778 + 8'h01;
  assign sel_979782 = array_index_979645 == array_index_948691 ? add_979781 : sel_979778;
  assign add_979785 = sel_979782 + 8'h01;
  assign sel_979786 = array_index_979645 == array_index_948697 ? add_979785 : sel_979782;
  assign add_979789 = sel_979786 + 8'h01;
  assign sel_979790 = array_index_979645 == array_index_948703 ? add_979789 : sel_979786;
  assign add_979793 = sel_979790 + 8'h01;
  assign sel_979794 = array_index_979645 == array_index_948709 ? add_979793 : sel_979790;
  assign add_979797 = sel_979794 + 8'h01;
  assign sel_979798 = array_index_979645 == array_index_948715 ? add_979797 : sel_979794;
  assign add_979801 = sel_979798 + 8'h01;
  assign sel_979802 = array_index_979645 == array_index_948721 ? add_979801 : sel_979798;
  assign add_979805 = sel_979802 + 8'h01;
  assign sel_979806 = array_index_979645 == array_index_948727 ? add_979805 : sel_979802;
  assign add_979809 = sel_979806 + 8'h01;
  assign sel_979810 = array_index_979645 == array_index_948733 ? add_979809 : sel_979806;
  assign add_979813 = sel_979810 + 8'h01;
  assign sel_979814 = array_index_979645 == array_index_948739 ? add_979813 : sel_979810;
  assign add_979817 = sel_979814 + 8'h01;
  assign sel_979818 = array_index_979645 == array_index_948745 ? add_979817 : sel_979814;
  assign add_979821 = sel_979818 + 8'h01;
  assign sel_979822 = array_index_979645 == array_index_948751 ? add_979821 : sel_979818;
  assign add_979825 = sel_979822 + 8'h01;
  assign sel_979826 = array_index_979645 == array_index_948757 ? add_979825 : sel_979822;
  assign add_979829 = sel_979826 + 8'h01;
  assign sel_979830 = array_index_979645 == array_index_948763 ? add_979829 : sel_979826;
  assign add_979833 = sel_979830 + 8'h01;
  assign sel_979834 = array_index_979645 == array_index_948769 ? add_979833 : sel_979830;
  assign add_979837 = sel_979834 + 8'h01;
  assign sel_979838 = array_index_979645 == array_index_948775 ? add_979837 : sel_979834;
  assign add_979841 = sel_979838 + 8'h01;
  assign sel_979842 = array_index_979645 == array_index_948781 ? add_979841 : sel_979838;
  assign add_979845 = sel_979842 + 8'h01;
  assign sel_979846 = array_index_979645 == array_index_948787 ? add_979845 : sel_979842;
  assign add_979849 = sel_979846 + 8'h01;
  assign sel_979850 = array_index_979645 == array_index_948793 ? add_979849 : sel_979846;
  assign add_979853 = sel_979850 + 8'h01;
  assign sel_979854 = array_index_979645 == array_index_948799 ? add_979853 : sel_979850;
  assign add_979857 = sel_979854 + 8'h01;
  assign sel_979858 = array_index_979645 == array_index_948805 ? add_979857 : sel_979854;
  assign add_979861 = sel_979858 + 8'h01;
  assign sel_979862 = array_index_979645 == array_index_948811 ? add_979861 : sel_979858;
  assign add_979865 = sel_979862 + 8'h01;
  assign sel_979866 = array_index_979645 == array_index_948817 ? add_979865 : sel_979862;
  assign add_979869 = sel_979866 + 8'h01;
  assign sel_979870 = array_index_979645 == array_index_948823 ? add_979869 : sel_979866;
  assign add_979873 = sel_979870 + 8'h01;
  assign sel_979874 = array_index_979645 == array_index_948829 ? add_979873 : sel_979870;
  assign add_979877 = sel_979874 + 8'h01;
  assign sel_979878 = array_index_979645 == array_index_948835 ? add_979877 : sel_979874;
  assign add_979881 = sel_979878 + 8'h01;
  assign sel_979882 = array_index_979645 == array_index_948841 ? add_979881 : sel_979878;
  assign add_979885 = sel_979882 + 8'h01;
  assign sel_979886 = array_index_979645 == array_index_948847 ? add_979885 : sel_979882;
  assign add_979889 = sel_979886 + 8'h01;
  assign sel_979890 = array_index_979645 == array_index_948853 ? add_979889 : sel_979886;
  assign add_979893 = sel_979890 + 8'h01;
  assign sel_979894 = array_index_979645 == array_index_948859 ? add_979893 : sel_979890;
  assign add_979897 = sel_979894 + 8'h01;
  assign sel_979898 = array_index_979645 == array_index_948865 ? add_979897 : sel_979894;
  assign add_979901 = sel_979898 + 8'h01;
  assign sel_979902 = array_index_979645 == array_index_948871 ? add_979901 : sel_979898;
  assign add_979905 = sel_979902 + 8'h01;
  assign sel_979906 = array_index_979645 == array_index_948877 ? add_979905 : sel_979902;
  assign add_979909 = sel_979906 + 8'h01;
  assign sel_979910 = array_index_979645 == array_index_948883 ? add_979909 : sel_979906;
  assign add_979913 = sel_979910 + 8'h01;
  assign sel_979914 = array_index_979645 == array_index_948889 ? add_979913 : sel_979910;
  assign add_979917 = sel_979914 + 8'h01;
  assign sel_979918 = array_index_979645 == array_index_948895 ? add_979917 : sel_979914;
  assign add_979921 = sel_979918 + 8'h01;
  assign sel_979922 = array_index_979645 == array_index_948901 ? add_979921 : sel_979918;
  assign add_979925 = sel_979922 + 8'h01;
  assign sel_979926 = array_index_979645 == array_index_948907 ? add_979925 : sel_979922;
  assign add_979929 = sel_979926 + 8'h01;
  assign sel_979930 = array_index_979645 == array_index_948913 ? add_979929 : sel_979926;
  assign add_979933 = sel_979930 + 8'h01;
  assign sel_979934 = array_index_979645 == array_index_948919 ? add_979933 : sel_979930;
  assign add_979937 = sel_979934 + 8'h01;
  assign sel_979938 = array_index_979645 == array_index_948925 ? add_979937 : sel_979934;
  assign add_979941 = sel_979938 + 8'h01;
  assign sel_979942 = array_index_979645 == array_index_948931 ? add_979941 : sel_979938;
  assign add_979945 = sel_979942 + 8'h01;
  assign sel_979946 = array_index_979645 == array_index_948937 ? add_979945 : sel_979942;
  assign add_979949 = sel_979946 + 8'h01;
  assign sel_979950 = array_index_979645 == array_index_948943 ? add_979949 : sel_979946;
  assign add_979953 = sel_979950 + 8'h01;
  assign sel_979954 = array_index_979645 == array_index_948949 ? add_979953 : sel_979950;
  assign add_979957 = sel_979954 + 8'h01;
  assign sel_979958 = array_index_979645 == array_index_948955 ? add_979957 : sel_979954;
  assign add_979961 = sel_979958 + 8'h01;
  assign sel_979962 = array_index_979645 == array_index_948961 ? add_979961 : sel_979958;
  assign add_979965 = sel_979962 + 8'h01;
  assign sel_979966 = array_index_979645 == array_index_948967 ? add_979965 : sel_979962;
  assign add_979969 = sel_979966 + 8'h01;
  assign sel_979970 = array_index_979645 == array_index_948973 ? add_979969 : sel_979966;
  assign add_979973 = sel_979970 + 8'h01;
  assign sel_979974 = array_index_979645 == array_index_948979 ? add_979973 : sel_979970;
  assign add_979977 = sel_979974 + 8'h01;
  assign sel_979978 = array_index_979645 == array_index_948985 ? add_979977 : sel_979974;
  assign add_979981 = sel_979978 + 8'h01;
  assign sel_979982 = array_index_979645 == array_index_948991 ? add_979981 : sel_979978;
  assign add_979985 = sel_979982 + 8'h01;
  assign sel_979986 = array_index_979645 == array_index_948997 ? add_979985 : sel_979982;
  assign add_979989 = sel_979986 + 8'h01;
  assign sel_979990 = array_index_979645 == array_index_949003 ? add_979989 : sel_979986;
  assign add_979993 = sel_979990 + 8'h01;
  assign sel_979994 = array_index_979645 == array_index_949009 ? add_979993 : sel_979990;
  assign add_979997 = sel_979994 + 8'h01;
  assign sel_979998 = array_index_979645 == array_index_949015 ? add_979997 : sel_979994;
  assign add_980001 = sel_979998 + 8'h01;
  assign sel_980002 = array_index_979645 == array_index_949021 ? add_980001 : sel_979998;
  assign add_980005 = sel_980002 + 8'h01;
  assign sel_980006 = array_index_979645 == array_index_949027 ? add_980005 : sel_980002;
  assign add_980009 = sel_980006 + 8'h01;
  assign sel_980010 = array_index_979645 == array_index_949033 ? add_980009 : sel_980006;
  assign add_980013 = sel_980010 + 8'h01;
  assign sel_980014 = array_index_979645 == array_index_949039 ? add_980013 : sel_980010;
  assign add_980017 = sel_980014 + 8'h01;
  assign sel_980018 = array_index_979645 == array_index_949045 ? add_980017 : sel_980014;
  assign add_980021 = sel_980018 + 8'h01;
  assign sel_980022 = array_index_979645 == array_index_949051 ? add_980021 : sel_980018;
  assign add_980025 = sel_980022 + 8'h01;
  assign sel_980026 = array_index_979645 == array_index_949057 ? add_980025 : sel_980022;
  assign add_980029 = sel_980026 + 8'h01;
  assign sel_980030 = array_index_979645 == array_index_949063 ? add_980029 : sel_980026;
  assign add_980033 = sel_980030 + 8'h01;
  assign sel_980034 = array_index_979645 == array_index_949069 ? add_980033 : sel_980030;
  assign add_980037 = sel_980034 + 8'h01;
  assign sel_980038 = array_index_979645 == array_index_949075 ? add_980037 : sel_980034;
  assign add_980041 = sel_980038 + 8'h01;
  assign sel_980042 = array_index_979645 == array_index_949081 ? add_980041 : sel_980038;
  assign add_980046 = sel_980042 + 8'h01;
  assign array_index_980047 = set1_unflattened[7'h4e];
  assign sel_980048 = array_index_979645 == array_index_949087 ? add_980046 : sel_980042;
  assign add_980051 = sel_980048 + 8'h01;
  assign sel_980052 = array_index_980047 == array_index_948483 ? add_980051 : sel_980048;
  assign add_980055 = sel_980052 + 8'h01;
  assign sel_980056 = array_index_980047 == array_index_948487 ? add_980055 : sel_980052;
  assign add_980059 = sel_980056 + 8'h01;
  assign sel_980060 = array_index_980047 == array_index_948495 ? add_980059 : sel_980056;
  assign add_980063 = sel_980060 + 8'h01;
  assign sel_980064 = array_index_980047 == array_index_948503 ? add_980063 : sel_980060;
  assign add_980067 = sel_980064 + 8'h01;
  assign sel_980068 = array_index_980047 == array_index_948511 ? add_980067 : sel_980064;
  assign add_980071 = sel_980068 + 8'h01;
  assign sel_980072 = array_index_980047 == array_index_948519 ? add_980071 : sel_980068;
  assign add_980075 = sel_980072 + 8'h01;
  assign sel_980076 = array_index_980047 == array_index_948527 ? add_980075 : sel_980072;
  assign add_980079 = sel_980076 + 8'h01;
  assign sel_980080 = array_index_980047 == array_index_948535 ? add_980079 : sel_980076;
  assign add_980083 = sel_980080 + 8'h01;
  assign sel_980084 = array_index_980047 == array_index_948541 ? add_980083 : sel_980080;
  assign add_980087 = sel_980084 + 8'h01;
  assign sel_980088 = array_index_980047 == array_index_948547 ? add_980087 : sel_980084;
  assign add_980091 = sel_980088 + 8'h01;
  assign sel_980092 = array_index_980047 == array_index_948553 ? add_980091 : sel_980088;
  assign add_980095 = sel_980092 + 8'h01;
  assign sel_980096 = array_index_980047 == array_index_948559 ? add_980095 : sel_980092;
  assign add_980099 = sel_980096 + 8'h01;
  assign sel_980100 = array_index_980047 == array_index_948565 ? add_980099 : sel_980096;
  assign add_980103 = sel_980100 + 8'h01;
  assign sel_980104 = array_index_980047 == array_index_948571 ? add_980103 : sel_980100;
  assign add_980107 = sel_980104 + 8'h01;
  assign sel_980108 = array_index_980047 == array_index_948577 ? add_980107 : sel_980104;
  assign add_980111 = sel_980108 + 8'h01;
  assign sel_980112 = array_index_980047 == array_index_948583 ? add_980111 : sel_980108;
  assign add_980115 = sel_980112 + 8'h01;
  assign sel_980116 = array_index_980047 == array_index_948589 ? add_980115 : sel_980112;
  assign add_980119 = sel_980116 + 8'h01;
  assign sel_980120 = array_index_980047 == array_index_948595 ? add_980119 : sel_980116;
  assign add_980123 = sel_980120 + 8'h01;
  assign sel_980124 = array_index_980047 == array_index_948601 ? add_980123 : sel_980120;
  assign add_980127 = sel_980124 + 8'h01;
  assign sel_980128 = array_index_980047 == array_index_948607 ? add_980127 : sel_980124;
  assign add_980131 = sel_980128 + 8'h01;
  assign sel_980132 = array_index_980047 == array_index_948613 ? add_980131 : sel_980128;
  assign add_980135 = sel_980132 + 8'h01;
  assign sel_980136 = array_index_980047 == array_index_948619 ? add_980135 : sel_980132;
  assign add_980139 = sel_980136 + 8'h01;
  assign sel_980140 = array_index_980047 == array_index_948625 ? add_980139 : sel_980136;
  assign add_980143 = sel_980140 + 8'h01;
  assign sel_980144 = array_index_980047 == array_index_948631 ? add_980143 : sel_980140;
  assign add_980147 = sel_980144 + 8'h01;
  assign sel_980148 = array_index_980047 == array_index_948637 ? add_980147 : sel_980144;
  assign add_980151 = sel_980148 + 8'h01;
  assign sel_980152 = array_index_980047 == array_index_948643 ? add_980151 : sel_980148;
  assign add_980155 = sel_980152 + 8'h01;
  assign sel_980156 = array_index_980047 == array_index_948649 ? add_980155 : sel_980152;
  assign add_980159 = sel_980156 + 8'h01;
  assign sel_980160 = array_index_980047 == array_index_948655 ? add_980159 : sel_980156;
  assign add_980163 = sel_980160 + 8'h01;
  assign sel_980164 = array_index_980047 == array_index_948661 ? add_980163 : sel_980160;
  assign add_980167 = sel_980164 + 8'h01;
  assign sel_980168 = array_index_980047 == array_index_948667 ? add_980167 : sel_980164;
  assign add_980171 = sel_980168 + 8'h01;
  assign sel_980172 = array_index_980047 == array_index_948673 ? add_980171 : sel_980168;
  assign add_980175 = sel_980172 + 8'h01;
  assign sel_980176 = array_index_980047 == array_index_948679 ? add_980175 : sel_980172;
  assign add_980179 = sel_980176 + 8'h01;
  assign sel_980180 = array_index_980047 == array_index_948685 ? add_980179 : sel_980176;
  assign add_980183 = sel_980180 + 8'h01;
  assign sel_980184 = array_index_980047 == array_index_948691 ? add_980183 : sel_980180;
  assign add_980187 = sel_980184 + 8'h01;
  assign sel_980188 = array_index_980047 == array_index_948697 ? add_980187 : sel_980184;
  assign add_980191 = sel_980188 + 8'h01;
  assign sel_980192 = array_index_980047 == array_index_948703 ? add_980191 : sel_980188;
  assign add_980195 = sel_980192 + 8'h01;
  assign sel_980196 = array_index_980047 == array_index_948709 ? add_980195 : sel_980192;
  assign add_980199 = sel_980196 + 8'h01;
  assign sel_980200 = array_index_980047 == array_index_948715 ? add_980199 : sel_980196;
  assign add_980203 = sel_980200 + 8'h01;
  assign sel_980204 = array_index_980047 == array_index_948721 ? add_980203 : sel_980200;
  assign add_980207 = sel_980204 + 8'h01;
  assign sel_980208 = array_index_980047 == array_index_948727 ? add_980207 : sel_980204;
  assign add_980211 = sel_980208 + 8'h01;
  assign sel_980212 = array_index_980047 == array_index_948733 ? add_980211 : sel_980208;
  assign add_980215 = sel_980212 + 8'h01;
  assign sel_980216 = array_index_980047 == array_index_948739 ? add_980215 : sel_980212;
  assign add_980219 = sel_980216 + 8'h01;
  assign sel_980220 = array_index_980047 == array_index_948745 ? add_980219 : sel_980216;
  assign add_980223 = sel_980220 + 8'h01;
  assign sel_980224 = array_index_980047 == array_index_948751 ? add_980223 : sel_980220;
  assign add_980227 = sel_980224 + 8'h01;
  assign sel_980228 = array_index_980047 == array_index_948757 ? add_980227 : sel_980224;
  assign add_980231 = sel_980228 + 8'h01;
  assign sel_980232 = array_index_980047 == array_index_948763 ? add_980231 : sel_980228;
  assign add_980235 = sel_980232 + 8'h01;
  assign sel_980236 = array_index_980047 == array_index_948769 ? add_980235 : sel_980232;
  assign add_980239 = sel_980236 + 8'h01;
  assign sel_980240 = array_index_980047 == array_index_948775 ? add_980239 : sel_980236;
  assign add_980243 = sel_980240 + 8'h01;
  assign sel_980244 = array_index_980047 == array_index_948781 ? add_980243 : sel_980240;
  assign add_980247 = sel_980244 + 8'h01;
  assign sel_980248 = array_index_980047 == array_index_948787 ? add_980247 : sel_980244;
  assign add_980251 = sel_980248 + 8'h01;
  assign sel_980252 = array_index_980047 == array_index_948793 ? add_980251 : sel_980248;
  assign add_980255 = sel_980252 + 8'h01;
  assign sel_980256 = array_index_980047 == array_index_948799 ? add_980255 : sel_980252;
  assign add_980259 = sel_980256 + 8'h01;
  assign sel_980260 = array_index_980047 == array_index_948805 ? add_980259 : sel_980256;
  assign add_980263 = sel_980260 + 8'h01;
  assign sel_980264 = array_index_980047 == array_index_948811 ? add_980263 : sel_980260;
  assign add_980267 = sel_980264 + 8'h01;
  assign sel_980268 = array_index_980047 == array_index_948817 ? add_980267 : sel_980264;
  assign add_980271 = sel_980268 + 8'h01;
  assign sel_980272 = array_index_980047 == array_index_948823 ? add_980271 : sel_980268;
  assign add_980275 = sel_980272 + 8'h01;
  assign sel_980276 = array_index_980047 == array_index_948829 ? add_980275 : sel_980272;
  assign add_980279 = sel_980276 + 8'h01;
  assign sel_980280 = array_index_980047 == array_index_948835 ? add_980279 : sel_980276;
  assign add_980283 = sel_980280 + 8'h01;
  assign sel_980284 = array_index_980047 == array_index_948841 ? add_980283 : sel_980280;
  assign add_980287 = sel_980284 + 8'h01;
  assign sel_980288 = array_index_980047 == array_index_948847 ? add_980287 : sel_980284;
  assign add_980291 = sel_980288 + 8'h01;
  assign sel_980292 = array_index_980047 == array_index_948853 ? add_980291 : sel_980288;
  assign add_980295 = sel_980292 + 8'h01;
  assign sel_980296 = array_index_980047 == array_index_948859 ? add_980295 : sel_980292;
  assign add_980299 = sel_980296 + 8'h01;
  assign sel_980300 = array_index_980047 == array_index_948865 ? add_980299 : sel_980296;
  assign add_980303 = sel_980300 + 8'h01;
  assign sel_980304 = array_index_980047 == array_index_948871 ? add_980303 : sel_980300;
  assign add_980307 = sel_980304 + 8'h01;
  assign sel_980308 = array_index_980047 == array_index_948877 ? add_980307 : sel_980304;
  assign add_980311 = sel_980308 + 8'h01;
  assign sel_980312 = array_index_980047 == array_index_948883 ? add_980311 : sel_980308;
  assign add_980315 = sel_980312 + 8'h01;
  assign sel_980316 = array_index_980047 == array_index_948889 ? add_980315 : sel_980312;
  assign add_980319 = sel_980316 + 8'h01;
  assign sel_980320 = array_index_980047 == array_index_948895 ? add_980319 : sel_980316;
  assign add_980323 = sel_980320 + 8'h01;
  assign sel_980324 = array_index_980047 == array_index_948901 ? add_980323 : sel_980320;
  assign add_980327 = sel_980324 + 8'h01;
  assign sel_980328 = array_index_980047 == array_index_948907 ? add_980327 : sel_980324;
  assign add_980331 = sel_980328 + 8'h01;
  assign sel_980332 = array_index_980047 == array_index_948913 ? add_980331 : sel_980328;
  assign add_980335 = sel_980332 + 8'h01;
  assign sel_980336 = array_index_980047 == array_index_948919 ? add_980335 : sel_980332;
  assign add_980339 = sel_980336 + 8'h01;
  assign sel_980340 = array_index_980047 == array_index_948925 ? add_980339 : sel_980336;
  assign add_980343 = sel_980340 + 8'h01;
  assign sel_980344 = array_index_980047 == array_index_948931 ? add_980343 : sel_980340;
  assign add_980347 = sel_980344 + 8'h01;
  assign sel_980348 = array_index_980047 == array_index_948937 ? add_980347 : sel_980344;
  assign add_980351 = sel_980348 + 8'h01;
  assign sel_980352 = array_index_980047 == array_index_948943 ? add_980351 : sel_980348;
  assign add_980355 = sel_980352 + 8'h01;
  assign sel_980356 = array_index_980047 == array_index_948949 ? add_980355 : sel_980352;
  assign add_980359 = sel_980356 + 8'h01;
  assign sel_980360 = array_index_980047 == array_index_948955 ? add_980359 : sel_980356;
  assign add_980363 = sel_980360 + 8'h01;
  assign sel_980364 = array_index_980047 == array_index_948961 ? add_980363 : sel_980360;
  assign add_980367 = sel_980364 + 8'h01;
  assign sel_980368 = array_index_980047 == array_index_948967 ? add_980367 : sel_980364;
  assign add_980371 = sel_980368 + 8'h01;
  assign sel_980372 = array_index_980047 == array_index_948973 ? add_980371 : sel_980368;
  assign add_980375 = sel_980372 + 8'h01;
  assign sel_980376 = array_index_980047 == array_index_948979 ? add_980375 : sel_980372;
  assign add_980379 = sel_980376 + 8'h01;
  assign sel_980380 = array_index_980047 == array_index_948985 ? add_980379 : sel_980376;
  assign add_980383 = sel_980380 + 8'h01;
  assign sel_980384 = array_index_980047 == array_index_948991 ? add_980383 : sel_980380;
  assign add_980387 = sel_980384 + 8'h01;
  assign sel_980388 = array_index_980047 == array_index_948997 ? add_980387 : sel_980384;
  assign add_980391 = sel_980388 + 8'h01;
  assign sel_980392 = array_index_980047 == array_index_949003 ? add_980391 : sel_980388;
  assign add_980395 = sel_980392 + 8'h01;
  assign sel_980396 = array_index_980047 == array_index_949009 ? add_980395 : sel_980392;
  assign add_980399 = sel_980396 + 8'h01;
  assign sel_980400 = array_index_980047 == array_index_949015 ? add_980399 : sel_980396;
  assign add_980403 = sel_980400 + 8'h01;
  assign sel_980404 = array_index_980047 == array_index_949021 ? add_980403 : sel_980400;
  assign add_980407 = sel_980404 + 8'h01;
  assign sel_980408 = array_index_980047 == array_index_949027 ? add_980407 : sel_980404;
  assign add_980411 = sel_980408 + 8'h01;
  assign sel_980412 = array_index_980047 == array_index_949033 ? add_980411 : sel_980408;
  assign add_980415 = sel_980412 + 8'h01;
  assign sel_980416 = array_index_980047 == array_index_949039 ? add_980415 : sel_980412;
  assign add_980419 = sel_980416 + 8'h01;
  assign sel_980420 = array_index_980047 == array_index_949045 ? add_980419 : sel_980416;
  assign add_980423 = sel_980420 + 8'h01;
  assign sel_980424 = array_index_980047 == array_index_949051 ? add_980423 : sel_980420;
  assign add_980427 = sel_980424 + 8'h01;
  assign sel_980428 = array_index_980047 == array_index_949057 ? add_980427 : sel_980424;
  assign add_980431 = sel_980428 + 8'h01;
  assign sel_980432 = array_index_980047 == array_index_949063 ? add_980431 : sel_980428;
  assign add_980435 = sel_980432 + 8'h01;
  assign sel_980436 = array_index_980047 == array_index_949069 ? add_980435 : sel_980432;
  assign add_980439 = sel_980436 + 8'h01;
  assign sel_980440 = array_index_980047 == array_index_949075 ? add_980439 : sel_980436;
  assign add_980443 = sel_980440 + 8'h01;
  assign sel_980444 = array_index_980047 == array_index_949081 ? add_980443 : sel_980440;
  assign add_980448 = sel_980444 + 8'h01;
  assign array_index_980449 = set1_unflattened[7'h4f];
  assign sel_980450 = array_index_980047 == array_index_949087 ? add_980448 : sel_980444;
  assign add_980453 = sel_980450 + 8'h01;
  assign sel_980454 = array_index_980449 == array_index_948483 ? add_980453 : sel_980450;
  assign add_980457 = sel_980454 + 8'h01;
  assign sel_980458 = array_index_980449 == array_index_948487 ? add_980457 : sel_980454;
  assign add_980461 = sel_980458 + 8'h01;
  assign sel_980462 = array_index_980449 == array_index_948495 ? add_980461 : sel_980458;
  assign add_980465 = sel_980462 + 8'h01;
  assign sel_980466 = array_index_980449 == array_index_948503 ? add_980465 : sel_980462;
  assign add_980469 = sel_980466 + 8'h01;
  assign sel_980470 = array_index_980449 == array_index_948511 ? add_980469 : sel_980466;
  assign add_980473 = sel_980470 + 8'h01;
  assign sel_980474 = array_index_980449 == array_index_948519 ? add_980473 : sel_980470;
  assign add_980477 = sel_980474 + 8'h01;
  assign sel_980478 = array_index_980449 == array_index_948527 ? add_980477 : sel_980474;
  assign add_980481 = sel_980478 + 8'h01;
  assign sel_980482 = array_index_980449 == array_index_948535 ? add_980481 : sel_980478;
  assign add_980485 = sel_980482 + 8'h01;
  assign sel_980486 = array_index_980449 == array_index_948541 ? add_980485 : sel_980482;
  assign add_980489 = sel_980486 + 8'h01;
  assign sel_980490 = array_index_980449 == array_index_948547 ? add_980489 : sel_980486;
  assign add_980493 = sel_980490 + 8'h01;
  assign sel_980494 = array_index_980449 == array_index_948553 ? add_980493 : sel_980490;
  assign add_980497 = sel_980494 + 8'h01;
  assign sel_980498 = array_index_980449 == array_index_948559 ? add_980497 : sel_980494;
  assign add_980501 = sel_980498 + 8'h01;
  assign sel_980502 = array_index_980449 == array_index_948565 ? add_980501 : sel_980498;
  assign add_980505 = sel_980502 + 8'h01;
  assign sel_980506 = array_index_980449 == array_index_948571 ? add_980505 : sel_980502;
  assign add_980509 = sel_980506 + 8'h01;
  assign sel_980510 = array_index_980449 == array_index_948577 ? add_980509 : sel_980506;
  assign add_980513 = sel_980510 + 8'h01;
  assign sel_980514 = array_index_980449 == array_index_948583 ? add_980513 : sel_980510;
  assign add_980517 = sel_980514 + 8'h01;
  assign sel_980518 = array_index_980449 == array_index_948589 ? add_980517 : sel_980514;
  assign add_980521 = sel_980518 + 8'h01;
  assign sel_980522 = array_index_980449 == array_index_948595 ? add_980521 : sel_980518;
  assign add_980525 = sel_980522 + 8'h01;
  assign sel_980526 = array_index_980449 == array_index_948601 ? add_980525 : sel_980522;
  assign add_980529 = sel_980526 + 8'h01;
  assign sel_980530 = array_index_980449 == array_index_948607 ? add_980529 : sel_980526;
  assign add_980533 = sel_980530 + 8'h01;
  assign sel_980534 = array_index_980449 == array_index_948613 ? add_980533 : sel_980530;
  assign add_980537 = sel_980534 + 8'h01;
  assign sel_980538 = array_index_980449 == array_index_948619 ? add_980537 : sel_980534;
  assign add_980541 = sel_980538 + 8'h01;
  assign sel_980542 = array_index_980449 == array_index_948625 ? add_980541 : sel_980538;
  assign add_980545 = sel_980542 + 8'h01;
  assign sel_980546 = array_index_980449 == array_index_948631 ? add_980545 : sel_980542;
  assign add_980549 = sel_980546 + 8'h01;
  assign sel_980550 = array_index_980449 == array_index_948637 ? add_980549 : sel_980546;
  assign add_980553 = sel_980550 + 8'h01;
  assign sel_980554 = array_index_980449 == array_index_948643 ? add_980553 : sel_980550;
  assign add_980557 = sel_980554 + 8'h01;
  assign sel_980558 = array_index_980449 == array_index_948649 ? add_980557 : sel_980554;
  assign add_980561 = sel_980558 + 8'h01;
  assign sel_980562 = array_index_980449 == array_index_948655 ? add_980561 : sel_980558;
  assign add_980565 = sel_980562 + 8'h01;
  assign sel_980566 = array_index_980449 == array_index_948661 ? add_980565 : sel_980562;
  assign add_980569 = sel_980566 + 8'h01;
  assign sel_980570 = array_index_980449 == array_index_948667 ? add_980569 : sel_980566;
  assign add_980573 = sel_980570 + 8'h01;
  assign sel_980574 = array_index_980449 == array_index_948673 ? add_980573 : sel_980570;
  assign add_980577 = sel_980574 + 8'h01;
  assign sel_980578 = array_index_980449 == array_index_948679 ? add_980577 : sel_980574;
  assign add_980581 = sel_980578 + 8'h01;
  assign sel_980582 = array_index_980449 == array_index_948685 ? add_980581 : sel_980578;
  assign add_980585 = sel_980582 + 8'h01;
  assign sel_980586 = array_index_980449 == array_index_948691 ? add_980585 : sel_980582;
  assign add_980589 = sel_980586 + 8'h01;
  assign sel_980590 = array_index_980449 == array_index_948697 ? add_980589 : sel_980586;
  assign add_980593 = sel_980590 + 8'h01;
  assign sel_980594 = array_index_980449 == array_index_948703 ? add_980593 : sel_980590;
  assign add_980597 = sel_980594 + 8'h01;
  assign sel_980598 = array_index_980449 == array_index_948709 ? add_980597 : sel_980594;
  assign add_980601 = sel_980598 + 8'h01;
  assign sel_980602 = array_index_980449 == array_index_948715 ? add_980601 : sel_980598;
  assign add_980605 = sel_980602 + 8'h01;
  assign sel_980606 = array_index_980449 == array_index_948721 ? add_980605 : sel_980602;
  assign add_980609 = sel_980606 + 8'h01;
  assign sel_980610 = array_index_980449 == array_index_948727 ? add_980609 : sel_980606;
  assign add_980613 = sel_980610 + 8'h01;
  assign sel_980614 = array_index_980449 == array_index_948733 ? add_980613 : sel_980610;
  assign add_980617 = sel_980614 + 8'h01;
  assign sel_980618 = array_index_980449 == array_index_948739 ? add_980617 : sel_980614;
  assign add_980621 = sel_980618 + 8'h01;
  assign sel_980622 = array_index_980449 == array_index_948745 ? add_980621 : sel_980618;
  assign add_980625 = sel_980622 + 8'h01;
  assign sel_980626 = array_index_980449 == array_index_948751 ? add_980625 : sel_980622;
  assign add_980629 = sel_980626 + 8'h01;
  assign sel_980630 = array_index_980449 == array_index_948757 ? add_980629 : sel_980626;
  assign add_980633 = sel_980630 + 8'h01;
  assign sel_980634 = array_index_980449 == array_index_948763 ? add_980633 : sel_980630;
  assign add_980637 = sel_980634 + 8'h01;
  assign sel_980638 = array_index_980449 == array_index_948769 ? add_980637 : sel_980634;
  assign add_980641 = sel_980638 + 8'h01;
  assign sel_980642 = array_index_980449 == array_index_948775 ? add_980641 : sel_980638;
  assign add_980645 = sel_980642 + 8'h01;
  assign sel_980646 = array_index_980449 == array_index_948781 ? add_980645 : sel_980642;
  assign add_980649 = sel_980646 + 8'h01;
  assign sel_980650 = array_index_980449 == array_index_948787 ? add_980649 : sel_980646;
  assign add_980653 = sel_980650 + 8'h01;
  assign sel_980654 = array_index_980449 == array_index_948793 ? add_980653 : sel_980650;
  assign add_980657 = sel_980654 + 8'h01;
  assign sel_980658 = array_index_980449 == array_index_948799 ? add_980657 : sel_980654;
  assign add_980661 = sel_980658 + 8'h01;
  assign sel_980662 = array_index_980449 == array_index_948805 ? add_980661 : sel_980658;
  assign add_980665 = sel_980662 + 8'h01;
  assign sel_980666 = array_index_980449 == array_index_948811 ? add_980665 : sel_980662;
  assign add_980669 = sel_980666 + 8'h01;
  assign sel_980670 = array_index_980449 == array_index_948817 ? add_980669 : sel_980666;
  assign add_980673 = sel_980670 + 8'h01;
  assign sel_980674 = array_index_980449 == array_index_948823 ? add_980673 : sel_980670;
  assign add_980677 = sel_980674 + 8'h01;
  assign sel_980678 = array_index_980449 == array_index_948829 ? add_980677 : sel_980674;
  assign add_980681 = sel_980678 + 8'h01;
  assign sel_980682 = array_index_980449 == array_index_948835 ? add_980681 : sel_980678;
  assign add_980685 = sel_980682 + 8'h01;
  assign sel_980686 = array_index_980449 == array_index_948841 ? add_980685 : sel_980682;
  assign add_980689 = sel_980686 + 8'h01;
  assign sel_980690 = array_index_980449 == array_index_948847 ? add_980689 : sel_980686;
  assign add_980693 = sel_980690 + 8'h01;
  assign sel_980694 = array_index_980449 == array_index_948853 ? add_980693 : sel_980690;
  assign add_980697 = sel_980694 + 8'h01;
  assign sel_980698 = array_index_980449 == array_index_948859 ? add_980697 : sel_980694;
  assign add_980701 = sel_980698 + 8'h01;
  assign sel_980702 = array_index_980449 == array_index_948865 ? add_980701 : sel_980698;
  assign add_980705 = sel_980702 + 8'h01;
  assign sel_980706 = array_index_980449 == array_index_948871 ? add_980705 : sel_980702;
  assign add_980709 = sel_980706 + 8'h01;
  assign sel_980710 = array_index_980449 == array_index_948877 ? add_980709 : sel_980706;
  assign add_980713 = sel_980710 + 8'h01;
  assign sel_980714 = array_index_980449 == array_index_948883 ? add_980713 : sel_980710;
  assign add_980717 = sel_980714 + 8'h01;
  assign sel_980718 = array_index_980449 == array_index_948889 ? add_980717 : sel_980714;
  assign add_980721 = sel_980718 + 8'h01;
  assign sel_980722 = array_index_980449 == array_index_948895 ? add_980721 : sel_980718;
  assign add_980725 = sel_980722 + 8'h01;
  assign sel_980726 = array_index_980449 == array_index_948901 ? add_980725 : sel_980722;
  assign add_980729 = sel_980726 + 8'h01;
  assign sel_980730 = array_index_980449 == array_index_948907 ? add_980729 : sel_980726;
  assign add_980733 = sel_980730 + 8'h01;
  assign sel_980734 = array_index_980449 == array_index_948913 ? add_980733 : sel_980730;
  assign add_980737 = sel_980734 + 8'h01;
  assign sel_980738 = array_index_980449 == array_index_948919 ? add_980737 : sel_980734;
  assign add_980741 = sel_980738 + 8'h01;
  assign sel_980742 = array_index_980449 == array_index_948925 ? add_980741 : sel_980738;
  assign add_980745 = sel_980742 + 8'h01;
  assign sel_980746 = array_index_980449 == array_index_948931 ? add_980745 : sel_980742;
  assign add_980749 = sel_980746 + 8'h01;
  assign sel_980750 = array_index_980449 == array_index_948937 ? add_980749 : sel_980746;
  assign add_980753 = sel_980750 + 8'h01;
  assign sel_980754 = array_index_980449 == array_index_948943 ? add_980753 : sel_980750;
  assign add_980757 = sel_980754 + 8'h01;
  assign sel_980758 = array_index_980449 == array_index_948949 ? add_980757 : sel_980754;
  assign add_980761 = sel_980758 + 8'h01;
  assign sel_980762 = array_index_980449 == array_index_948955 ? add_980761 : sel_980758;
  assign add_980765 = sel_980762 + 8'h01;
  assign sel_980766 = array_index_980449 == array_index_948961 ? add_980765 : sel_980762;
  assign add_980769 = sel_980766 + 8'h01;
  assign sel_980770 = array_index_980449 == array_index_948967 ? add_980769 : sel_980766;
  assign add_980773 = sel_980770 + 8'h01;
  assign sel_980774 = array_index_980449 == array_index_948973 ? add_980773 : sel_980770;
  assign add_980777 = sel_980774 + 8'h01;
  assign sel_980778 = array_index_980449 == array_index_948979 ? add_980777 : sel_980774;
  assign add_980781 = sel_980778 + 8'h01;
  assign sel_980782 = array_index_980449 == array_index_948985 ? add_980781 : sel_980778;
  assign add_980785 = sel_980782 + 8'h01;
  assign sel_980786 = array_index_980449 == array_index_948991 ? add_980785 : sel_980782;
  assign add_980789 = sel_980786 + 8'h01;
  assign sel_980790 = array_index_980449 == array_index_948997 ? add_980789 : sel_980786;
  assign add_980793 = sel_980790 + 8'h01;
  assign sel_980794 = array_index_980449 == array_index_949003 ? add_980793 : sel_980790;
  assign add_980797 = sel_980794 + 8'h01;
  assign sel_980798 = array_index_980449 == array_index_949009 ? add_980797 : sel_980794;
  assign add_980801 = sel_980798 + 8'h01;
  assign sel_980802 = array_index_980449 == array_index_949015 ? add_980801 : sel_980798;
  assign add_980805 = sel_980802 + 8'h01;
  assign sel_980806 = array_index_980449 == array_index_949021 ? add_980805 : sel_980802;
  assign add_980809 = sel_980806 + 8'h01;
  assign sel_980810 = array_index_980449 == array_index_949027 ? add_980809 : sel_980806;
  assign add_980813 = sel_980810 + 8'h01;
  assign sel_980814 = array_index_980449 == array_index_949033 ? add_980813 : sel_980810;
  assign add_980817 = sel_980814 + 8'h01;
  assign sel_980818 = array_index_980449 == array_index_949039 ? add_980817 : sel_980814;
  assign add_980821 = sel_980818 + 8'h01;
  assign sel_980822 = array_index_980449 == array_index_949045 ? add_980821 : sel_980818;
  assign add_980825 = sel_980822 + 8'h01;
  assign sel_980826 = array_index_980449 == array_index_949051 ? add_980825 : sel_980822;
  assign add_980829 = sel_980826 + 8'h01;
  assign sel_980830 = array_index_980449 == array_index_949057 ? add_980829 : sel_980826;
  assign add_980833 = sel_980830 + 8'h01;
  assign sel_980834 = array_index_980449 == array_index_949063 ? add_980833 : sel_980830;
  assign add_980837 = sel_980834 + 8'h01;
  assign sel_980838 = array_index_980449 == array_index_949069 ? add_980837 : sel_980834;
  assign add_980841 = sel_980838 + 8'h01;
  assign sel_980842 = array_index_980449 == array_index_949075 ? add_980841 : sel_980838;
  assign add_980845 = sel_980842 + 8'h01;
  assign sel_980846 = array_index_980449 == array_index_949081 ? add_980845 : sel_980842;
  assign add_980850 = sel_980846 + 8'h01;
  assign array_index_980851 = set1_unflattened[7'h50];
  assign sel_980852 = array_index_980449 == array_index_949087 ? add_980850 : sel_980846;
  assign add_980855 = sel_980852 + 8'h01;
  assign sel_980856 = array_index_980851 == array_index_948483 ? add_980855 : sel_980852;
  assign add_980859 = sel_980856 + 8'h01;
  assign sel_980860 = array_index_980851 == array_index_948487 ? add_980859 : sel_980856;
  assign add_980863 = sel_980860 + 8'h01;
  assign sel_980864 = array_index_980851 == array_index_948495 ? add_980863 : sel_980860;
  assign add_980867 = sel_980864 + 8'h01;
  assign sel_980868 = array_index_980851 == array_index_948503 ? add_980867 : sel_980864;
  assign add_980871 = sel_980868 + 8'h01;
  assign sel_980872 = array_index_980851 == array_index_948511 ? add_980871 : sel_980868;
  assign add_980875 = sel_980872 + 8'h01;
  assign sel_980876 = array_index_980851 == array_index_948519 ? add_980875 : sel_980872;
  assign add_980879 = sel_980876 + 8'h01;
  assign sel_980880 = array_index_980851 == array_index_948527 ? add_980879 : sel_980876;
  assign add_980883 = sel_980880 + 8'h01;
  assign sel_980884 = array_index_980851 == array_index_948535 ? add_980883 : sel_980880;
  assign add_980887 = sel_980884 + 8'h01;
  assign sel_980888 = array_index_980851 == array_index_948541 ? add_980887 : sel_980884;
  assign add_980891 = sel_980888 + 8'h01;
  assign sel_980892 = array_index_980851 == array_index_948547 ? add_980891 : sel_980888;
  assign add_980895 = sel_980892 + 8'h01;
  assign sel_980896 = array_index_980851 == array_index_948553 ? add_980895 : sel_980892;
  assign add_980899 = sel_980896 + 8'h01;
  assign sel_980900 = array_index_980851 == array_index_948559 ? add_980899 : sel_980896;
  assign add_980903 = sel_980900 + 8'h01;
  assign sel_980904 = array_index_980851 == array_index_948565 ? add_980903 : sel_980900;
  assign add_980907 = sel_980904 + 8'h01;
  assign sel_980908 = array_index_980851 == array_index_948571 ? add_980907 : sel_980904;
  assign add_980911 = sel_980908 + 8'h01;
  assign sel_980912 = array_index_980851 == array_index_948577 ? add_980911 : sel_980908;
  assign add_980915 = sel_980912 + 8'h01;
  assign sel_980916 = array_index_980851 == array_index_948583 ? add_980915 : sel_980912;
  assign add_980919 = sel_980916 + 8'h01;
  assign sel_980920 = array_index_980851 == array_index_948589 ? add_980919 : sel_980916;
  assign add_980923 = sel_980920 + 8'h01;
  assign sel_980924 = array_index_980851 == array_index_948595 ? add_980923 : sel_980920;
  assign add_980927 = sel_980924 + 8'h01;
  assign sel_980928 = array_index_980851 == array_index_948601 ? add_980927 : sel_980924;
  assign add_980931 = sel_980928 + 8'h01;
  assign sel_980932 = array_index_980851 == array_index_948607 ? add_980931 : sel_980928;
  assign add_980935 = sel_980932 + 8'h01;
  assign sel_980936 = array_index_980851 == array_index_948613 ? add_980935 : sel_980932;
  assign add_980939 = sel_980936 + 8'h01;
  assign sel_980940 = array_index_980851 == array_index_948619 ? add_980939 : sel_980936;
  assign add_980943 = sel_980940 + 8'h01;
  assign sel_980944 = array_index_980851 == array_index_948625 ? add_980943 : sel_980940;
  assign add_980947 = sel_980944 + 8'h01;
  assign sel_980948 = array_index_980851 == array_index_948631 ? add_980947 : sel_980944;
  assign add_980951 = sel_980948 + 8'h01;
  assign sel_980952 = array_index_980851 == array_index_948637 ? add_980951 : sel_980948;
  assign add_980955 = sel_980952 + 8'h01;
  assign sel_980956 = array_index_980851 == array_index_948643 ? add_980955 : sel_980952;
  assign add_980959 = sel_980956 + 8'h01;
  assign sel_980960 = array_index_980851 == array_index_948649 ? add_980959 : sel_980956;
  assign add_980963 = sel_980960 + 8'h01;
  assign sel_980964 = array_index_980851 == array_index_948655 ? add_980963 : sel_980960;
  assign add_980967 = sel_980964 + 8'h01;
  assign sel_980968 = array_index_980851 == array_index_948661 ? add_980967 : sel_980964;
  assign add_980971 = sel_980968 + 8'h01;
  assign sel_980972 = array_index_980851 == array_index_948667 ? add_980971 : sel_980968;
  assign add_980975 = sel_980972 + 8'h01;
  assign sel_980976 = array_index_980851 == array_index_948673 ? add_980975 : sel_980972;
  assign add_980979 = sel_980976 + 8'h01;
  assign sel_980980 = array_index_980851 == array_index_948679 ? add_980979 : sel_980976;
  assign add_980983 = sel_980980 + 8'h01;
  assign sel_980984 = array_index_980851 == array_index_948685 ? add_980983 : sel_980980;
  assign add_980987 = sel_980984 + 8'h01;
  assign sel_980988 = array_index_980851 == array_index_948691 ? add_980987 : sel_980984;
  assign add_980991 = sel_980988 + 8'h01;
  assign sel_980992 = array_index_980851 == array_index_948697 ? add_980991 : sel_980988;
  assign add_980995 = sel_980992 + 8'h01;
  assign sel_980996 = array_index_980851 == array_index_948703 ? add_980995 : sel_980992;
  assign add_980999 = sel_980996 + 8'h01;
  assign sel_981000 = array_index_980851 == array_index_948709 ? add_980999 : sel_980996;
  assign add_981003 = sel_981000 + 8'h01;
  assign sel_981004 = array_index_980851 == array_index_948715 ? add_981003 : sel_981000;
  assign add_981007 = sel_981004 + 8'h01;
  assign sel_981008 = array_index_980851 == array_index_948721 ? add_981007 : sel_981004;
  assign add_981011 = sel_981008 + 8'h01;
  assign sel_981012 = array_index_980851 == array_index_948727 ? add_981011 : sel_981008;
  assign add_981015 = sel_981012 + 8'h01;
  assign sel_981016 = array_index_980851 == array_index_948733 ? add_981015 : sel_981012;
  assign add_981019 = sel_981016 + 8'h01;
  assign sel_981020 = array_index_980851 == array_index_948739 ? add_981019 : sel_981016;
  assign add_981023 = sel_981020 + 8'h01;
  assign sel_981024 = array_index_980851 == array_index_948745 ? add_981023 : sel_981020;
  assign add_981027 = sel_981024 + 8'h01;
  assign sel_981028 = array_index_980851 == array_index_948751 ? add_981027 : sel_981024;
  assign add_981031 = sel_981028 + 8'h01;
  assign sel_981032 = array_index_980851 == array_index_948757 ? add_981031 : sel_981028;
  assign add_981035 = sel_981032 + 8'h01;
  assign sel_981036 = array_index_980851 == array_index_948763 ? add_981035 : sel_981032;
  assign add_981039 = sel_981036 + 8'h01;
  assign sel_981040 = array_index_980851 == array_index_948769 ? add_981039 : sel_981036;
  assign add_981043 = sel_981040 + 8'h01;
  assign sel_981044 = array_index_980851 == array_index_948775 ? add_981043 : sel_981040;
  assign add_981047 = sel_981044 + 8'h01;
  assign sel_981048 = array_index_980851 == array_index_948781 ? add_981047 : sel_981044;
  assign add_981051 = sel_981048 + 8'h01;
  assign sel_981052 = array_index_980851 == array_index_948787 ? add_981051 : sel_981048;
  assign add_981055 = sel_981052 + 8'h01;
  assign sel_981056 = array_index_980851 == array_index_948793 ? add_981055 : sel_981052;
  assign add_981059 = sel_981056 + 8'h01;
  assign sel_981060 = array_index_980851 == array_index_948799 ? add_981059 : sel_981056;
  assign add_981063 = sel_981060 + 8'h01;
  assign sel_981064 = array_index_980851 == array_index_948805 ? add_981063 : sel_981060;
  assign add_981067 = sel_981064 + 8'h01;
  assign sel_981068 = array_index_980851 == array_index_948811 ? add_981067 : sel_981064;
  assign add_981071 = sel_981068 + 8'h01;
  assign sel_981072 = array_index_980851 == array_index_948817 ? add_981071 : sel_981068;
  assign add_981075 = sel_981072 + 8'h01;
  assign sel_981076 = array_index_980851 == array_index_948823 ? add_981075 : sel_981072;
  assign add_981079 = sel_981076 + 8'h01;
  assign sel_981080 = array_index_980851 == array_index_948829 ? add_981079 : sel_981076;
  assign add_981083 = sel_981080 + 8'h01;
  assign sel_981084 = array_index_980851 == array_index_948835 ? add_981083 : sel_981080;
  assign add_981087 = sel_981084 + 8'h01;
  assign sel_981088 = array_index_980851 == array_index_948841 ? add_981087 : sel_981084;
  assign add_981091 = sel_981088 + 8'h01;
  assign sel_981092 = array_index_980851 == array_index_948847 ? add_981091 : sel_981088;
  assign add_981095 = sel_981092 + 8'h01;
  assign sel_981096 = array_index_980851 == array_index_948853 ? add_981095 : sel_981092;
  assign add_981099 = sel_981096 + 8'h01;
  assign sel_981100 = array_index_980851 == array_index_948859 ? add_981099 : sel_981096;
  assign add_981103 = sel_981100 + 8'h01;
  assign sel_981104 = array_index_980851 == array_index_948865 ? add_981103 : sel_981100;
  assign add_981107 = sel_981104 + 8'h01;
  assign sel_981108 = array_index_980851 == array_index_948871 ? add_981107 : sel_981104;
  assign add_981111 = sel_981108 + 8'h01;
  assign sel_981112 = array_index_980851 == array_index_948877 ? add_981111 : sel_981108;
  assign add_981115 = sel_981112 + 8'h01;
  assign sel_981116 = array_index_980851 == array_index_948883 ? add_981115 : sel_981112;
  assign add_981119 = sel_981116 + 8'h01;
  assign sel_981120 = array_index_980851 == array_index_948889 ? add_981119 : sel_981116;
  assign add_981123 = sel_981120 + 8'h01;
  assign sel_981124 = array_index_980851 == array_index_948895 ? add_981123 : sel_981120;
  assign add_981127 = sel_981124 + 8'h01;
  assign sel_981128 = array_index_980851 == array_index_948901 ? add_981127 : sel_981124;
  assign add_981131 = sel_981128 + 8'h01;
  assign sel_981132 = array_index_980851 == array_index_948907 ? add_981131 : sel_981128;
  assign add_981135 = sel_981132 + 8'h01;
  assign sel_981136 = array_index_980851 == array_index_948913 ? add_981135 : sel_981132;
  assign add_981139 = sel_981136 + 8'h01;
  assign sel_981140 = array_index_980851 == array_index_948919 ? add_981139 : sel_981136;
  assign add_981143 = sel_981140 + 8'h01;
  assign sel_981144 = array_index_980851 == array_index_948925 ? add_981143 : sel_981140;
  assign add_981147 = sel_981144 + 8'h01;
  assign sel_981148 = array_index_980851 == array_index_948931 ? add_981147 : sel_981144;
  assign add_981151 = sel_981148 + 8'h01;
  assign sel_981152 = array_index_980851 == array_index_948937 ? add_981151 : sel_981148;
  assign add_981155 = sel_981152 + 8'h01;
  assign sel_981156 = array_index_980851 == array_index_948943 ? add_981155 : sel_981152;
  assign add_981159 = sel_981156 + 8'h01;
  assign sel_981160 = array_index_980851 == array_index_948949 ? add_981159 : sel_981156;
  assign add_981163 = sel_981160 + 8'h01;
  assign sel_981164 = array_index_980851 == array_index_948955 ? add_981163 : sel_981160;
  assign add_981167 = sel_981164 + 8'h01;
  assign sel_981168 = array_index_980851 == array_index_948961 ? add_981167 : sel_981164;
  assign add_981171 = sel_981168 + 8'h01;
  assign sel_981172 = array_index_980851 == array_index_948967 ? add_981171 : sel_981168;
  assign add_981175 = sel_981172 + 8'h01;
  assign sel_981176 = array_index_980851 == array_index_948973 ? add_981175 : sel_981172;
  assign add_981179 = sel_981176 + 8'h01;
  assign sel_981180 = array_index_980851 == array_index_948979 ? add_981179 : sel_981176;
  assign add_981183 = sel_981180 + 8'h01;
  assign sel_981184 = array_index_980851 == array_index_948985 ? add_981183 : sel_981180;
  assign add_981187 = sel_981184 + 8'h01;
  assign sel_981188 = array_index_980851 == array_index_948991 ? add_981187 : sel_981184;
  assign add_981191 = sel_981188 + 8'h01;
  assign sel_981192 = array_index_980851 == array_index_948997 ? add_981191 : sel_981188;
  assign add_981195 = sel_981192 + 8'h01;
  assign sel_981196 = array_index_980851 == array_index_949003 ? add_981195 : sel_981192;
  assign add_981199 = sel_981196 + 8'h01;
  assign sel_981200 = array_index_980851 == array_index_949009 ? add_981199 : sel_981196;
  assign add_981203 = sel_981200 + 8'h01;
  assign sel_981204 = array_index_980851 == array_index_949015 ? add_981203 : sel_981200;
  assign add_981207 = sel_981204 + 8'h01;
  assign sel_981208 = array_index_980851 == array_index_949021 ? add_981207 : sel_981204;
  assign add_981211 = sel_981208 + 8'h01;
  assign sel_981212 = array_index_980851 == array_index_949027 ? add_981211 : sel_981208;
  assign add_981215 = sel_981212 + 8'h01;
  assign sel_981216 = array_index_980851 == array_index_949033 ? add_981215 : sel_981212;
  assign add_981219 = sel_981216 + 8'h01;
  assign sel_981220 = array_index_980851 == array_index_949039 ? add_981219 : sel_981216;
  assign add_981223 = sel_981220 + 8'h01;
  assign sel_981224 = array_index_980851 == array_index_949045 ? add_981223 : sel_981220;
  assign add_981227 = sel_981224 + 8'h01;
  assign sel_981228 = array_index_980851 == array_index_949051 ? add_981227 : sel_981224;
  assign add_981231 = sel_981228 + 8'h01;
  assign sel_981232 = array_index_980851 == array_index_949057 ? add_981231 : sel_981228;
  assign add_981235 = sel_981232 + 8'h01;
  assign sel_981236 = array_index_980851 == array_index_949063 ? add_981235 : sel_981232;
  assign add_981239 = sel_981236 + 8'h01;
  assign sel_981240 = array_index_980851 == array_index_949069 ? add_981239 : sel_981236;
  assign add_981243 = sel_981240 + 8'h01;
  assign sel_981244 = array_index_980851 == array_index_949075 ? add_981243 : sel_981240;
  assign add_981247 = sel_981244 + 8'h01;
  assign sel_981248 = array_index_980851 == array_index_949081 ? add_981247 : sel_981244;
  assign add_981252 = sel_981248 + 8'h01;
  assign array_index_981253 = set1_unflattened[7'h51];
  assign sel_981254 = array_index_980851 == array_index_949087 ? add_981252 : sel_981248;
  assign add_981257 = sel_981254 + 8'h01;
  assign sel_981258 = array_index_981253 == array_index_948483 ? add_981257 : sel_981254;
  assign add_981261 = sel_981258 + 8'h01;
  assign sel_981262 = array_index_981253 == array_index_948487 ? add_981261 : sel_981258;
  assign add_981265 = sel_981262 + 8'h01;
  assign sel_981266 = array_index_981253 == array_index_948495 ? add_981265 : sel_981262;
  assign add_981269 = sel_981266 + 8'h01;
  assign sel_981270 = array_index_981253 == array_index_948503 ? add_981269 : sel_981266;
  assign add_981273 = sel_981270 + 8'h01;
  assign sel_981274 = array_index_981253 == array_index_948511 ? add_981273 : sel_981270;
  assign add_981277 = sel_981274 + 8'h01;
  assign sel_981278 = array_index_981253 == array_index_948519 ? add_981277 : sel_981274;
  assign add_981281 = sel_981278 + 8'h01;
  assign sel_981282 = array_index_981253 == array_index_948527 ? add_981281 : sel_981278;
  assign add_981285 = sel_981282 + 8'h01;
  assign sel_981286 = array_index_981253 == array_index_948535 ? add_981285 : sel_981282;
  assign add_981289 = sel_981286 + 8'h01;
  assign sel_981290 = array_index_981253 == array_index_948541 ? add_981289 : sel_981286;
  assign add_981293 = sel_981290 + 8'h01;
  assign sel_981294 = array_index_981253 == array_index_948547 ? add_981293 : sel_981290;
  assign add_981297 = sel_981294 + 8'h01;
  assign sel_981298 = array_index_981253 == array_index_948553 ? add_981297 : sel_981294;
  assign add_981301 = sel_981298 + 8'h01;
  assign sel_981302 = array_index_981253 == array_index_948559 ? add_981301 : sel_981298;
  assign add_981305 = sel_981302 + 8'h01;
  assign sel_981306 = array_index_981253 == array_index_948565 ? add_981305 : sel_981302;
  assign add_981309 = sel_981306 + 8'h01;
  assign sel_981310 = array_index_981253 == array_index_948571 ? add_981309 : sel_981306;
  assign add_981313 = sel_981310 + 8'h01;
  assign sel_981314 = array_index_981253 == array_index_948577 ? add_981313 : sel_981310;
  assign add_981317 = sel_981314 + 8'h01;
  assign sel_981318 = array_index_981253 == array_index_948583 ? add_981317 : sel_981314;
  assign add_981321 = sel_981318 + 8'h01;
  assign sel_981322 = array_index_981253 == array_index_948589 ? add_981321 : sel_981318;
  assign add_981325 = sel_981322 + 8'h01;
  assign sel_981326 = array_index_981253 == array_index_948595 ? add_981325 : sel_981322;
  assign add_981329 = sel_981326 + 8'h01;
  assign sel_981330 = array_index_981253 == array_index_948601 ? add_981329 : sel_981326;
  assign add_981333 = sel_981330 + 8'h01;
  assign sel_981334 = array_index_981253 == array_index_948607 ? add_981333 : sel_981330;
  assign add_981337 = sel_981334 + 8'h01;
  assign sel_981338 = array_index_981253 == array_index_948613 ? add_981337 : sel_981334;
  assign add_981341 = sel_981338 + 8'h01;
  assign sel_981342 = array_index_981253 == array_index_948619 ? add_981341 : sel_981338;
  assign add_981345 = sel_981342 + 8'h01;
  assign sel_981346 = array_index_981253 == array_index_948625 ? add_981345 : sel_981342;
  assign add_981349 = sel_981346 + 8'h01;
  assign sel_981350 = array_index_981253 == array_index_948631 ? add_981349 : sel_981346;
  assign add_981353 = sel_981350 + 8'h01;
  assign sel_981354 = array_index_981253 == array_index_948637 ? add_981353 : sel_981350;
  assign add_981357 = sel_981354 + 8'h01;
  assign sel_981358 = array_index_981253 == array_index_948643 ? add_981357 : sel_981354;
  assign add_981361 = sel_981358 + 8'h01;
  assign sel_981362 = array_index_981253 == array_index_948649 ? add_981361 : sel_981358;
  assign add_981365 = sel_981362 + 8'h01;
  assign sel_981366 = array_index_981253 == array_index_948655 ? add_981365 : sel_981362;
  assign add_981369 = sel_981366 + 8'h01;
  assign sel_981370 = array_index_981253 == array_index_948661 ? add_981369 : sel_981366;
  assign add_981373 = sel_981370 + 8'h01;
  assign sel_981374 = array_index_981253 == array_index_948667 ? add_981373 : sel_981370;
  assign add_981377 = sel_981374 + 8'h01;
  assign sel_981378 = array_index_981253 == array_index_948673 ? add_981377 : sel_981374;
  assign add_981381 = sel_981378 + 8'h01;
  assign sel_981382 = array_index_981253 == array_index_948679 ? add_981381 : sel_981378;
  assign add_981385 = sel_981382 + 8'h01;
  assign sel_981386 = array_index_981253 == array_index_948685 ? add_981385 : sel_981382;
  assign add_981389 = sel_981386 + 8'h01;
  assign sel_981390 = array_index_981253 == array_index_948691 ? add_981389 : sel_981386;
  assign add_981393 = sel_981390 + 8'h01;
  assign sel_981394 = array_index_981253 == array_index_948697 ? add_981393 : sel_981390;
  assign add_981397 = sel_981394 + 8'h01;
  assign sel_981398 = array_index_981253 == array_index_948703 ? add_981397 : sel_981394;
  assign add_981401 = sel_981398 + 8'h01;
  assign sel_981402 = array_index_981253 == array_index_948709 ? add_981401 : sel_981398;
  assign add_981405 = sel_981402 + 8'h01;
  assign sel_981406 = array_index_981253 == array_index_948715 ? add_981405 : sel_981402;
  assign add_981409 = sel_981406 + 8'h01;
  assign sel_981410 = array_index_981253 == array_index_948721 ? add_981409 : sel_981406;
  assign add_981413 = sel_981410 + 8'h01;
  assign sel_981414 = array_index_981253 == array_index_948727 ? add_981413 : sel_981410;
  assign add_981417 = sel_981414 + 8'h01;
  assign sel_981418 = array_index_981253 == array_index_948733 ? add_981417 : sel_981414;
  assign add_981421 = sel_981418 + 8'h01;
  assign sel_981422 = array_index_981253 == array_index_948739 ? add_981421 : sel_981418;
  assign add_981425 = sel_981422 + 8'h01;
  assign sel_981426 = array_index_981253 == array_index_948745 ? add_981425 : sel_981422;
  assign add_981429 = sel_981426 + 8'h01;
  assign sel_981430 = array_index_981253 == array_index_948751 ? add_981429 : sel_981426;
  assign add_981433 = sel_981430 + 8'h01;
  assign sel_981434 = array_index_981253 == array_index_948757 ? add_981433 : sel_981430;
  assign add_981437 = sel_981434 + 8'h01;
  assign sel_981438 = array_index_981253 == array_index_948763 ? add_981437 : sel_981434;
  assign add_981441 = sel_981438 + 8'h01;
  assign sel_981442 = array_index_981253 == array_index_948769 ? add_981441 : sel_981438;
  assign add_981445 = sel_981442 + 8'h01;
  assign sel_981446 = array_index_981253 == array_index_948775 ? add_981445 : sel_981442;
  assign add_981449 = sel_981446 + 8'h01;
  assign sel_981450 = array_index_981253 == array_index_948781 ? add_981449 : sel_981446;
  assign add_981453 = sel_981450 + 8'h01;
  assign sel_981454 = array_index_981253 == array_index_948787 ? add_981453 : sel_981450;
  assign add_981457 = sel_981454 + 8'h01;
  assign sel_981458 = array_index_981253 == array_index_948793 ? add_981457 : sel_981454;
  assign add_981461 = sel_981458 + 8'h01;
  assign sel_981462 = array_index_981253 == array_index_948799 ? add_981461 : sel_981458;
  assign add_981465 = sel_981462 + 8'h01;
  assign sel_981466 = array_index_981253 == array_index_948805 ? add_981465 : sel_981462;
  assign add_981469 = sel_981466 + 8'h01;
  assign sel_981470 = array_index_981253 == array_index_948811 ? add_981469 : sel_981466;
  assign add_981473 = sel_981470 + 8'h01;
  assign sel_981474 = array_index_981253 == array_index_948817 ? add_981473 : sel_981470;
  assign add_981477 = sel_981474 + 8'h01;
  assign sel_981478 = array_index_981253 == array_index_948823 ? add_981477 : sel_981474;
  assign add_981481 = sel_981478 + 8'h01;
  assign sel_981482 = array_index_981253 == array_index_948829 ? add_981481 : sel_981478;
  assign add_981485 = sel_981482 + 8'h01;
  assign sel_981486 = array_index_981253 == array_index_948835 ? add_981485 : sel_981482;
  assign add_981489 = sel_981486 + 8'h01;
  assign sel_981490 = array_index_981253 == array_index_948841 ? add_981489 : sel_981486;
  assign add_981493 = sel_981490 + 8'h01;
  assign sel_981494 = array_index_981253 == array_index_948847 ? add_981493 : sel_981490;
  assign add_981497 = sel_981494 + 8'h01;
  assign sel_981498 = array_index_981253 == array_index_948853 ? add_981497 : sel_981494;
  assign add_981501 = sel_981498 + 8'h01;
  assign sel_981502 = array_index_981253 == array_index_948859 ? add_981501 : sel_981498;
  assign add_981505 = sel_981502 + 8'h01;
  assign sel_981506 = array_index_981253 == array_index_948865 ? add_981505 : sel_981502;
  assign add_981509 = sel_981506 + 8'h01;
  assign sel_981510 = array_index_981253 == array_index_948871 ? add_981509 : sel_981506;
  assign add_981513 = sel_981510 + 8'h01;
  assign sel_981514 = array_index_981253 == array_index_948877 ? add_981513 : sel_981510;
  assign add_981517 = sel_981514 + 8'h01;
  assign sel_981518 = array_index_981253 == array_index_948883 ? add_981517 : sel_981514;
  assign add_981521 = sel_981518 + 8'h01;
  assign sel_981522 = array_index_981253 == array_index_948889 ? add_981521 : sel_981518;
  assign add_981525 = sel_981522 + 8'h01;
  assign sel_981526 = array_index_981253 == array_index_948895 ? add_981525 : sel_981522;
  assign add_981529 = sel_981526 + 8'h01;
  assign sel_981530 = array_index_981253 == array_index_948901 ? add_981529 : sel_981526;
  assign add_981533 = sel_981530 + 8'h01;
  assign sel_981534 = array_index_981253 == array_index_948907 ? add_981533 : sel_981530;
  assign add_981537 = sel_981534 + 8'h01;
  assign sel_981538 = array_index_981253 == array_index_948913 ? add_981537 : sel_981534;
  assign add_981541 = sel_981538 + 8'h01;
  assign sel_981542 = array_index_981253 == array_index_948919 ? add_981541 : sel_981538;
  assign add_981545 = sel_981542 + 8'h01;
  assign sel_981546 = array_index_981253 == array_index_948925 ? add_981545 : sel_981542;
  assign add_981549 = sel_981546 + 8'h01;
  assign sel_981550 = array_index_981253 == array_index_948931 ? add_981549 : sel_981546;
  assign add_981553 = sel_981550 + 8'h01;
  assign sel_981554 = array_index_981253 == array_index_948937 ? add_981553 : sel_981550;
  assign add_981557 = sel_981554 + 8'h01;
  assign sel_981558 = array_index_981253 == array_index_948943 ? add_981557 : sel_981554;
  assign add_981561 = sel_981558 + 8'h01;
  assign sel_981562 = array_index_981253 == array_index_948949 ? add_981561 : sel_981558;
  assign add_981565 = sel_981562 + 8'h01;
  assign sel_981566 = array_index_981253 == array_index_948955 ? add_981565 : sel_981562;
  assign add_981569 = sel_981566 + 8'h01;
  assign sel_981570 = array_index_981253 == array_index_948961 ? add_981569 : sel_981566;
  assign add_981573 = sel_981570 + 8'h01;
  assign sel_981574 = array_index_981253 == array_index_948967 ? add_981573 : sel_981570;
  assign add_981577 = sel_981574 + 8'h01;
  assign sel_981578 = array_index_981253 == array_index_948973 ? add_981577 : sel_981574;
  assign add_981581 = sel_981578 + 8'h01;
  assign sel_981582 = array_index_981253 == array_index_948979 ? add_981581 : sel_981578;
  assign add_981585 = sel_981582 + 8'h01;
  assign sel_981586 = array_index_981253 == array_index_948985 ? add_981585 : sel_981582;
  assign add_981589 = sel_981586 + 8'h01;
  assign sel_981590 = array_index_981253 == array_index_948991 ? add_981589 : sel_981586;
  assign add_981593 = sel_981590 + 8'h01;
  assign sel_981594 = array_index_981253 == array_index_948997 ? add_981593 : sel_981590;
  assign add_981597 = sel_981594 + 8'h01;
  assign sel_981598 = array_index_981253 == array_index_949003 ? add_981597 : sel_981594;
  assign add_981601 = sel_981598 + 8'h01;
  assign sel_981602 = array_index_981253 == array_index_949009 ? add_981601 : sel_981598;
  assign add_981605 = sel_981602 + 8'h01;
  assign sel_981606 = array_index_981253 == array_index_949015 ? add_981605 : sel_981602;
  assign add_981609 = sel_981606 + 8'h01;
  assign sel_981610 = array_index_981253 == array_index_949021 ? add_981609 : sel_981606;
  assign add_981613 = sel_981610 + 8'h01;
  assign sel_981614 = array_index_981253 == array_index_949027 ? add_981613 : sel_981610;
  assign add_981617 = sel_981614 + 8'h01;
  assign sel_981618 = array_index_981253 == array_index_949033 ? add_981617 : sel_981614;
  assign add_981621 = sel_981618 + 8'h01;
  assign sel_981622 = array_index_981253 == array_index_949039 ? add_981621 : sel_981618;
  assign add_981625 = sel_981622 + 8'h01;
  assign sel_981626 = array_index_981253 == array_index_949045 ? add_981625 : sel_981622;
  assign add_981629 = sel_981626 + 8'h01;
  assign sel_981630 = array_index_981253 == array_index_949051 ? add_981629 : sel_981626;
  assign add_981633 = sel_981630 + 8'h01;
  assign sel_981634 = array_index_981253 == array_index_949057 ? add_981633 : sel_981630;
  assign add_981637 = sel_981634 + 8'h01;
  assign sel_981638 = array_index_981253 == array_index_949063 ? add_981637 : sel_981634;
  assign add_981641 = sel_981638 + 8'h01;
  assign sel_981642 = array_index_981253 == array_index_949069 ? add_981641 : sel_981638;
  assign add_981645 = sel_981642 + 8'h01;
  assign sel_981646 = array_index_981253 == array_index_949075 ? add_981645 : sel_981642;
  assign add_981649 = sel_981646 + 8'h01;
  assign sel_981650 = array_index_981253 == array_index_949081 ? add_981649 : sel_981646;
  assign add_981654 = sel_981650 + 8'h01;
  assign array_index_981655 = set1_unflattened[7'h52];
  assign sel_981656 = array_index_981253 == array_index_949087 ? add_981654 : sel_981650;
  assign add_981659 = sel_981656 + 8'h01;
  assign sel_981660 = array_index_981655 == array_index_948483 ? add_981659 : sel_981656;
  assign add_981663 = sel_981660 + 8'h01;
  assign sel_981664 = array_index_981655 == array_index_948487 ? add_981663 : sel_981660;
  assign add_981667 = sel_981664 + 8'h01;
  assign sel_981668 = array_index_981655 == array_index_948495 ? add_981667 : sel_981664;
  assign add_981671 = sel_981668 + 8'h01;
  assign sel_981672 = array_index_981655 == array_index_948503 ? add_981671 : sel_981668;
  assign add_981675 = sel_981672 + 8'h01;
  assign sel_981676 = array_index_981655 == array_index_948511 ? add_981675 : sel_981672;
  assign add_981679 = sel_981676 + 8'h01;
  assign sel_981680 = array_index_981655 == array_index_948519 ? add_981679 : sel_981676;
  assign add_981683 = sel_981680 + 8'h01;
  assign sel_981684 = array_index_981655 == array_index_948527 ? add_981683 : sel_981680;
  assign add_981687 = sel_981684 + 8'h01;
  assign sel_981688 = array_index_981655 == array_index_948535 ? add_981687 : sel_981684;
  assign add_981691 = sel_981688 + 8'h01;
  assign sel_981692 = array_index_981655 == array_index_948541 ? add_981691 : sel_981688;
  assign add_981695 = sel_981692 + 8'h01;
  assign sel_981696 = array_index_981655 == array_index_948547 ? add_981695 : sel_981692;
  assign add_981699 = sel_981696 + 8'h01;
  assign sel_981700 = array_index_981655 == array_index_948553 ? add_981699 : sel_981696;
  assign add_981703 = sel_981700 + 8'h01;
  assign sel_981704 = array_index_981655 == array_index_948559 ? add_981703 : sel_981700;
  assign add_981707 = sel_981704 + 8'h01;
  assign sel_981708 = array_index_981655 == array_index_948565 ? add_981707 : sel_981704;
  assign add_981711 = sel_981708 + 8'h01;
  assign sel_981712 = array_index_981655 == array_index_948571 ? add_981711 : sel_981708;
  assign add_981715 = sel_981712 + 8'h01;
  assign sel_981716 = array_index_981655 == array_index_948577 ? add_981715 : sel_981712;
  assign add_981719 = sel_981716 + 8'h01;
  assign sel_981720 = array_index_981655 == array_index_948583 ? add_981719 : sel_981716;
  assign add_981723 = sel_981720 + 8'h01;
  assign sel_981724 = array_index_981655 == array_index_948589 ? add_981723 : sel_981720;
  assign add_981727 = sel_981724 + 8'h01;
  assign sel_981728 = array_index_981655 == array_index_948595 ? add_981727 : sel_981724;
  assign add_981731 = sel_981728 + 8'h01;
  assign sel_981732 = array_index_981655 == array_index_948601 ? add_981731 : sel_981728;
  assign add_981735 = sel_981732 + 8'h01;
  assign sel_981736 = array_index_981655 == array_index_948607 ? add_981735 : sel_981732;
  assign add_981739 = sel_981736 + 8'h01;
  assign sel_981740 = array_index_981655 == array_index_948613 ? add_981739 : sel_981736;
  assign add_981743 = sel_981740 + 8'h01;
  assign sel_981744 = array_index_981655 == array_index_948619 ? add_981743 : sel_981740;
  assign add_981747 = sel_981744 + 8'h01;
  assign sel_981748 = array_index_981655 == array_index_948625 ? add_981747 : sel_981744;
  assign add_981751 = sel_981748 + 8'h01;
  assign sel_981752 = array_index_981655 == array_index_948631 ? add_981751 : sel_981748;
  assign add_981755 = sel_981752 + 8'h01;
  assign sel_981756 = array_index_981655 == array_index_948637 ? add_981755 : sel_981752;
  assign add_981759 = sel_981756 + 8'h01;
  assign sel_981760 = array_index_981655 == array_index_948643 ? add_981759 : sel_981756;
  assign add_981763 = sel_981760 + 8'h01;
  assign sel_981764 = array_index_981655 == array_index_948649 ? add_981763 : sel_981760;
  assign add_981767 = sel_981764 + 8'h01;
  assign sel_981768 = array_index_981655 == array_index_948655 ? add_981767 : sel_981764;
  assign add_981771 = sel_981768 + 8'h01;
  assign sel_981772 = array_index_981655 == array_index_948661 ? add_981771 : sel_981768;
  assign add_981775 = sel_981772 + 8'h01;
  assign sel_981776 = array_index_981655 == array_index_948667 ? add_981775 : sel_981772;
  assign add_981779 = sel_981776 + 8'h01;
  assign sel_981780 = array_index_981655 == array_index_948673 ? add_981779 : sel_981776;
  assign add_981783 = sel_981780 + 8'h01;
  assign sel_981784 = array_index_981655 == array_index_948679 ? add_981783 : sel_981780;
  assign add_981787 = sel_981784 + 8'h01;
  assign sel_981788 = array_index_981655 == array_index_948685 ? add_981787 : sel_981784;
  assign add_981791 = sel_981788 + 8'h01;
  assign sel_981792 = array_index_981655 == array_index_948691 ? add_981791 : sel_981788;
  assign add_981795 = sel_981792 + 8'h01;
  assign sel_981796 = array_index_981655 == array_index_948697 ? add_981795 : sel_981792;
  assign add_981799 = sel_981796 + 8'h01;
  assign sel_981800 = array_index_981655 == array_index_948703 ? add_981799 : sel_981796;
  assign add_981803 = sel_981800 + 8'h01;
  assign sel_981804 = array_index_981655 == array_index_948709 ? add_981803 : sel_981800;
  assign add_981807 = sel_981804 + 8'h01;
  assign sel_981808 = array_index_981655 == array_index_948715 ? add_981807 : sel_981804;
  assign add_981811 = sel_981808 + 8'h01;
  assign sel_981812 = array_index_981655 == array_index_948721 ? add_981811 : sel_981808;
  assign add_981815 = sel_981812 + 8'h01;
  assign sel_981816 = array_index_981655 == array_index_948727 ? add_981815 : sel_981812;
  assign add_981819 = sel_981816 + 8'h01;
  assign sel_981820 = array_index_981655 == array_index_948733 ? add_981819 : sel_981816;
  assign add_981823 = sel_981820 + 8'h01;
  assign sel_981824 = array_index_981655 == array_index_948739 ? add_981823 : sel_981820;
  assign add_981827 = sel_981824 + 8'h01;
  assign sel_981828 = array_index_981655 == array_index_948745 ? add_981827 : sel_981824;
  assign add_981831 = sel_981828 + 8'h01;
  assign sel_981832 = array_index_981655 == array_index_948751 ? add_981831 : sel_981828;
  assign add_981835 = sel_981832 + 8'h01;
  assign sel_981836 = array_index_981655 == array_index_948757 ? add_981835 : sel_981832;
  assign add_981839 = sel_981836 + 8'h01;
  assign sel_981840 = array_index_981655 == array_index_948763 ? add_981839 : sel_981836;
  assign add_981843 = sel_981840 + 8'h01;
  assign sel_981844 = array_index_981655 == array_index_948769 ? add_981843 : sel_981840;
  assign add_981847 = sel_981844 + 8'h01;
  assign sel_981848 = array_index_981655 == array_index_948775 ? add_981847 : sel_981844;
  assign add_981851 = sel_981848 + 8'h01;
  assign sel_981852 = array_index_981655 == array_index_948781 ? add_981851 : sel_981848;
  assign add_981855 = sel_981852 + 8'h01;
  assign sel_981856 = array_index_981655 == array_index_948787 ? add_981855 : sel_981852;
  assign add_981859 = sel_981856 + 8'h01;
  assign sel_981860 = array_index_981655 == array_index_948793 ? add_981859 : sel_981856;
  assign add_981863 = sel_981860 + 8'h01;
  assign sel_981864 = array_index_981655 == array_index_948799 ? add_981863 : sel_981860;
  assign add_981867 = sel_981864 + 8'h01;
  assign sel_981868 = array_index_981655 == array_index_948805 ? add_981867 : sel_981864;
  assign add_981871 = sel_981868 + 8'h01;
  assign sel_981872 = array_index_981655 == array_index_948811 ? add_981871 : sel_981868;
  assign add_981875 = sel_981872 + 8'h01;
  assign sel_981876 = array_index_981655 == array_index_948817 ? add_981875 : sel_981872;
  assign add_981879 = sel_981876 + 8'h01;
  assign sel_981880 = array_index_981655 == array_index_948823 ? add_981879 : sel_981876;
  assign add_981883 = sel_981880 + 8'h01;
  assign sel_981884 = array_index_981655 == array_index_948829 ? add_981883 : sel_981880;
  assign add_981887 = sel_981884 + 8'h01;
  assign sel_981888 = array_index_981655 == array_index_948835 ? add_981887 : sel_981884;
  assign add_981891 = sel_981888 + 8'h01;
  assign sel_981892 = array_index_981655 == array_index_948841 ? add_981891 : sel_981888;
  assign add_981895 = sel_981892 + 8'h01;
  assign sel_981896 = array_index_981655 == array_index_948847 ? add_981895 : sel_981892;
  assign add_981899 = sel_981896 + 8'h01;
  assign sel_981900 = array_index_981655 == array_index_948853 ? add_981899 : sel_981896;
  assign add_981903 = sel_981900 + 8'h01;
  assign sel_981904 = array_index_981655 == array_index_948859 ? add_981903 : sel_981900;
  assign add_981907 = sel_981904 + 8'h01;
  assign sel_981908 = array_index_981655 == array_index_948865 ? add_981907 : sel_981904;
  assign add_981911 = sel_981908 + 8'h01;
  assign sel_981912 = array_index_981655 == array_index_948871 ? add_981911 : sel_981908;
  assign add_981915 = sel_981912 + 8'h01;
  assign sel_981916 = array_index_981655 == array_index_948877 ? add_981915 : sel_981912;
  assign add_981919 = sel_981916 + 8'h01;
  assign sel_981920 = array_index_981655 == array_index_948883 ? add_981919 : sel_981916;
  assign add_981923 = sel_981920 + 8'h01;
  assign sel_981924 = array_index_981655 == array_index_948889 ? add_981923 : sel_981920;
  assign add_981927 = sel_981924 + 8'h01;
  assign sel_981928 = array_index_981655 == array_index_948895 ? add_981927 : sel_981924;
  assign add_981931 = sel_981928 + 8'h01;
  assign sel_981932 = array_index_981655 == array_index_948901 ? add_981931 : sel_981928;
  assign add_981935 = sel_981932 + 8'h01;
  assign sel_981936 = array_index_981655 == array_index_948907 ? add_981935 : sel_981932;
  assign add_981939 = sel_981936 + 8'h01;
  assign sel_981940 = array_index_981655 == array_index_948913 ? add_981939 : sel_981936;
  assign add_981943 = sel_981940 + 8'h01;
  assign sel_981944 = array_index_981655 == array_index_948919 ? add_981943 : sel_981940;
  assign add_981947 = sel_981944 + 8'h01;
  assign sel_981948 = array_index_981655 == array_index_948925 ? add_981947 : sel_981944;
  assign add_981951 = sel_981948 + 8'h01;
  assign sel_981952 = array_index_981655 == array_index_948931 ? add_981951 : sel_981948;
  assign add_981955 = sel_981952 + 8'h01;
  assign sel_981956 = array_index_981655 == array_index_948937 ? add_981955 : sel_981952;
  assign add_981959 = sel_981956 + 8'h01;
  assign sel_981960 = array_index_981655 == array_index_948943 ? add_981959 : sel_981956;
  assign add_981963 = sel_981960 + 8'h01;
  assign sel_981964 = array_index_981655 == array_index_948949 ? add_981963 : sel_981960;
  assign add_981967 = sel_981964 + 8'h01;
  assign sel_981968 = array_index_981655 == array_index_948955 ? add_981967 : sel_981964;
  assign add_981971 = sel_981968 + 8'h01;
  assign sel_981972 = array_index_981655 == array_index_948961 ? add_981971 : sel_981968;
  assign add_981975 = sel_981972 + 8'h01;
  assign sel_981976 = array_index_981655 == array_index_948967 ? add_981975 : sel_981972;
  assign add_981979 = sel_981976 + 8'h01;
  assign sel_981980 = array_index_981655 == array_index_948973 ? add_981979 : sel_981976;
  assign add_981983 = sel_981980 + 8'h01;
  assign sel_981984 = array_index_981655 == array_index_948979 ? add_981983 : sel_981980;
  assign add_981987 = sel_981984 + 8'h01;
  assign sel_981988 = array_index_981655 == array_index_948985 ? add_981987 : sel_981984;
  assign add_981991 = sel_981988 + 8'h01;
  assign sel_981992 = array_index_981655 == array_index_948991 ? add_981991 : sel_981988;
  assign add_981995 = sel_981992 + 8'h01;
  assign sel_981996 = array_index_981655 == array_index_948997 ? add_981995 : sel_981992;
  assign add_981999 = sel_981996 + 8'h01;
  assign sel_982000 = array_index_981655 == array_index_949003 ? add_981999 : sel_981996;
  assign add_982003 = sel_982000 + 8'h01;
  assign sel_982004 = array_index_981655 == array_index_949009 ? add_982003 : sel_982000;
  assign add_982007 = sel_982004 + 8'h01;
  assign sel_982008 = array_index_981655 == array_index_949015 ? add_982007 : sel_982004;
  assign add_982011 = sel_982008 + 8'h01;
  assign sel_982012 = array_index_981655 == array_index_949021 ? add_982011 : sel_982008;
  assign add_982015 = sel_982012 + 8'h01;
  assign sel_982016 = array_index_981655 == array_index_949027 ? add_982015 : sel_982012;
  assign add_982019 = sel_982016 + 8'h01;
  assign sel_982020 = array_index_981655 == array_index_949033 ? add_982019 : sel_982016;
  assign add_982023 = sel_982020 + 8'h01;
  assign sel_982024 = array_index_981655 == array_index_949039 ? add_982023 : sel_982020;
  assign add_982027 = sel_982024 + 8'h01;
  assign sel_982028 = array_index_981655 == array_index_949045 ? add_982027 : sel_982024;
  assign add_982031 = sel_982028 + 8'h01;
  assign sel_982032 = array_index_981655 == array_index_949051 ? add_982031 : sel_982028;
  assign add_982035 = sel_982032 + 8'h01;
  assign sel_982036 = array_index_981655 == array_index_949057 ? add_982035 : sel_982032;
  assign add_982039 = sel_982036 + 8'h01;
  assign sel_982040 = array_index_981655 == array_index_949063 ? add_982039 : sel_982036;
  assign add_982043 = sel_982040 + 8'h01;
  assign sel_982044 = array_index_981655 == array_index_949069 ? add_982043 : sel_982040;
  assign add_982047 = sel_982044 + 8'h01;
  assign sel_982048 = array_index_981655 == array_index_949075 ? add_982047 : sel_982044;
  assign add_982051 = sel_982048 + 8'h01;
  assign sel_982052 = array_index_981655 == array_index_949081 ? add_982051 : sel_982048;
  assign add_982056 = sel_982052 + 8'h01;
  assign array_index_982057 = set1_unflattened[7'h53];
  assign sel_982058 = array_index_981655 == array_index_949087 ? add_982056 : sel_982052;
  assign add_982061 = sel_982058 + 8'h01;
  assign sel_982062 = array_index_982057 == array_index_948483 ? add_982061 : sel_982058;
  assign add_982065 = sel_982062 + 8'h01;
  assign sel_982066 = array_index_982057 == array_index_948487 ? add_982065 : sel_982062;
  assign add_982069 = sel_982066 + 8'h01;
  assign sel_982070 = array_index_982057 == array_index_948495 ? add_982069 : sel_982066;
  assign add_982073 = sel_982070 + 8'h01;
  assign sel_982074 = array_index_982057 == array_index_948503 ? add_982073 : sel_982070;
  assign add_982077 = sel_982074 + 8'h01;
  assign sel_982078 = array_index_982057 == array_index_948511 ? add_982077 : sel_982074;
  assign add_982081 = sel_982078 + 8'h01;
  assign sel_982082 = array_index_982057 == array_index_948519 ? add_982081 : sel_982078;
  assign add_982085 = sel_982082 + 8'h01;
  assign sel_982086 = array_index_982057 == array_index_948527 ? add_982085 : sel_982082;
  assign add_982089 = sel_982086 + 8'h01;
  assign sel_982090 = array_index_982057 == array_index_948535 ? add_982089 : sel_982086;
  assign add_982093 = sel_982090 + 8'h01;
  assign sel_982094 = array_index_982057 == array_index_948541 ? add_982093 : sel_982090;
  assign add_982097 = sel_982094 + 8'h01;
  assign sel_982098 = array_index_982057 == array_index_948547 ? add_982097 : sel_982094;
  assign add_982101 = sel_982098 + 8'h01;
  assign sel_982102 = array_index_982057 == array_index_948553 ? add_982101 : sel_982098;
  assign add_982105 = sel_982102 + 8'h01;
  assign sel_982106 = array_index_982057 == array_index_948559 ? add_982105 : sel_982102;
  assign add_982109 = sel_982106 + 8'h01;
  assign sel_982110 = array_index_982057 == array_index_948565 ? add_982109 : sel_982106;
  assign add_982113 = sel_982110 + 8'h01;
  assign sel_982114 = array_index_982057 == array_index_948571 ? add_982113 : sel_982110;
  assign add_982117 = sel_982114 + 8'h01;
  assign sel_982118 = array_index_982057 == array_index_948577 ? add_982117 : sel_982114;
  assign add_982121 = sel_982118 + 8'h01;
  assign sel_982122 = array_index_982057 == array_index_948583 ? add_982121 : sel_982118;
  assign add_982125 = sel_982122 + 8'h01;
  assign sel_982126 = array_index_982057 == array_index_948589 ? add_982125 : sel_982122;
  assign add_982129 = sel_982126 + 8'h01;
  assign sel_982130 = array_index_982057 == array_index_948595 ? add_982129 : sel_982126;
  assign add_982133 = sel_982130 + 8'h01;
  assign sel_982134 = array_index_982057 == array_index_948601 ? add_982133 : sel_982130;
  assign add_982137 = sel_982134 + 8'h01;
  assign sel_982138 = array_index_982057 == array_index_948607 ? add_982137 : sel_982134;
  assign add_982141 = sel_982138 + 8'h01;
  assign sel_982142 = array_index_982057 == array_index_948613 ? add_982141 : sel_982138;
  assign add_982145 = sel_982142 + 8'h01;
  assign sel_982146 = array_index_982057 == array_index_948619 ? add_982145 : sel_982142;
  assign add_982149 = sel_982146 + 8'h01;
  assign sel_982150 = array_index_982057 == array_index_948625 ? add_982149 : sel_982146;
  assign add_982153 = sel_982150 + 8'h01;
  assign sel_982154 = array_index_982057 == array_index_948631 ? add_982153 : sel_982150;
  assign add_982157 = sel_982154 + 8'h01;
  assign sel_982158 = array_index_982057 == array_index_948637 ? add_982157 : sel_982154;
  assign add_982161 = sel_982158 + 8'h01;
  assign sel_982162 = array_index_982057 == array_index_948643 ? add_982161 : sel_982158;
  assign add_982165 = sel_982162 + 8'h01;
  assign sel_982166 = array_index_982057 == array_index_948649 ? add_982165 : sel_982162;
  assign add_982169 = sel_982166 + 8'h01;
  assign sel_982170 = array_index_982057 == array_index_948655 ? add_982169 : sel_982166;
  assign add_982173 = sel_982170 + 8'h01;
  assign sel_982174 = array_index_982057 == array_index_948661 ? add_982173 : sel_982170;
  assign add_982177 = sel_982174 + 8'h01;
  assign sel_982178 = array_index_982057 == array_index_948667 ? add_982177 : sel_982174;
  assign add_982181 = sel_982178 + 8'h01;
  assign sel_982182 = array_index_982057 == array_index_948673 ? add_982181 : sel_982178;
  assign add_982185 = sel_982182 + 8'h01;
  assign sel_982186 = array_index_982057 == array_index_948679 ? add_982185 : sel_982182;
  assign add_982189 = sel_982186 + 8'h01;
  assign sel_982190 = array_index_982057 == array_index_948685 ? add_982189 : sel_982186;
  assign add_982193 = sel_982190 + 8'h01;
  assign sel_982194 = array_index_982057 == array_index_948691 ? add_982193 : sel_982190;
  assign add_982197 = sel_982194 + 8'h01;
  assign sel_982198 = array_index_982057 == array_index_948697 ? add_982197 : sel_982194;
  assign add_982201 = sel_982198 + 8'h01;
  assign sel_982202 = array_index_982057 == array_index_948703 ? add_982201 : sel_982198;
  assign add_982205 = sel_982202 + 8'h01;
  assign sel_982206 = array_index_982057 == array_index_948709 ? add_982205 : sel_982202;
  assign add_982209 = sel_982206 + 8'h01;
  assign sel_982210 = array_index_982057 == array_index_948715 ? add_982209 : sel_982206;
  assign add_982213 = sel_982210 + 8'h01;
  assign sel_982214 = array_index_982057 == array_index_948721 ? add_982213 : sel_982210;
  assign add_982217 = sel_982214 + 8'h01;
  assign sel_982218 = array_index_982057 == array_index_948727 ? add_982217 : sel_982214;
  assign add_982221 = sel_982218 + 8'h01;
  assign sel_982222 = array_index_982057 == array_index_948733 ? add_982221 : sel_982218;
  assign add_982225 = sel_982222 + 8'h01;
  assign sel_982226 = array_index_982057 == array_index_948739 ? add_982225 : sel_982222;
  assign add_982229 = sel_982226 + 8'h01;
  assign sel_982230 = array_index_982057 == array_index_948745 ? add_982229 : sel_982226;
  assign add_982233 = sel_982230 + 8'h01;
  assign sel_982234 = array_index_982057 == array_index_948751 ? add_982233 : sel_982230;
  assign add_982237 = sel_982234 + 8'h01;
  assign sel_982238 = array_index_982057 == array_index_948757 ? add_982237 : sel_982234;
  assign add_982241 = sel_982238 + 8'h01;
  assign sel_982242 = array_index_982057 == array_index_948763 ? add_982241 : sel_982238;
  assign add_982245 = sel_982242 + 8'h01;
  assign sel_982246 = array_index_982057 == array_index_948769 ? add_982245 : sel_982242;
  assign add_982249 = sel_982246 + 8'h01;
  assign sel_982250 = array_index_982057 == array_index_948775 ? add_982249 : sel_982246;
  assign add_982253 = sel_982250 + 8'h01;
  assign sel_982254 = array_index_982057 == array_index_948781 ? add_982253 : sel_982250;
  assign add_982257 = sel_982254 + 8'h01;
  assign sel_982258 = array_index_982057 == array_index_948787 ? add_982257 : sel_982254;
  assign add_982261 = sel_982258 + 8'h01;
  assign sel_982262 = array_index_982057 == array_index_948793 ? add_982261 : sel_982258;
  assign add_982265 = sel_982262 + 8'h01;
  assign sel_982266 = array_index_982057 == array_index_948799 ? add_982265 : sel_982262;
  assign add_982269 = sel_982266 + 8'h01;
  assign sel_982270 = array_index_982057 == array_index_948805 ? add_982269 : sel_982266;
  assign add_982273 = sel_982270 + 8'h01;
  assign sel_982274 = array_index_982057 == array_index_948811 ? add_982273 : sel_982270;
  assign add_982277 = sel_982274 + 8'h01;
  assign sel_982278 = array_index_982057 == array_index_948817 ? add_982277 : sel_982274;
  assign add_982281 = sel_982278 + 8'h01;
  assign sel_982282 = array_index_982057 == array_index_948823 ? add_982281 : sel_982278;
  assign add_982285 = sel_982282 + 8'h01;
  assign sel_982286 = array_index_982057 == array_index_948829 ? add_982285 : sel_982282;
  assign add_982289 = sel_982286 + 8'h01;
  assign sel_982290 = array_index_982057 == array_index_948835 ? add_982289 : sel_982286;
  assign add_982293 = sel_982290 + 8'h01;
  assign sel_982294 = array_index_982057 == array_index_948841 ? add_982293 : sel_982290;
  assign add_982297 = sel_982294 + 8'h01;
  assign sel_982298 = array_index_982057 == array_index_948847 ? add_982297 : sel_982294;
  assign add_982301 = sel_982298 + 8'h01;
  assign sel_982302 = array_index_982057 == array_index_948853 ? add_982301 : sel_982298;
  assign add_982305 = sel_982302 + 8'h01;
  assign sel_982306 = array_index_982057 == array_index_948859 ? add_982305 : sel_982302;
  assign add_982309 = sel_982306 + 8'h01;
  assign sel_982310 = array_index_982057 == array_index_948865 ? add_982309 : sel_982306;
  assign add_982313 = sel_982310 + 8'h01;
  assign sel_982314 = array_index_982057 == array_index_948871 ? add_982313 : sel_982310;
  assign add_982317 = sel_982314 + 8'h01;
  assign sel_982318 = array_index_982057 == array_index_948877 ? add_982317 : sel_982314;
  assign add_982321 = sel_982318 + 8'h01;
  assign sel_982322 = array_index_982057 == array_index_948883 ? add_982321 : sel_982318;
  assign add_982325 = sel_982322 + 8'h01;
  assign sel_982326 = array_index_982057 == array_index_948889 ? add_982325 : sel_982322;
  assign add_982329 = sel_982326 + 8'h01;
  assign sel_982330 = array_index_982057 == array_index_948895 ? add_982329 : sel_982326;
  assign add_982333 = sel_982330 + 8'h01;
  assign sel_982334 = array_index_982057 == array_index_948901 ? add_982333 : sel_982330;
  assign add_982337 = sel_982334 + 8'h01;
  assign sel_982338 = array_index_982057 == array_index_948907 ? add_982337 : sel_982334;
  assign add_982341 = sel_982338 + 8'h01;
  assign sel_982342 = array_index_982057 == array_index_948913 ? add_982341 : sel_982338;
  assign add_982345 = sel_982342 + 8'h01;
  assign sel_982346 = array_index_982057 == array_index_948919 ? add_982345 : sel_982342;
  assign add_982349 = sel_982346 + 8'h01;
  assign sel_982350 = array_index_982057 == array_index_948925 ? add_982349 : sel_982346;
  assign add_982353 = sel_982350 + 8'h01;
  assign sel_982354 = array_index_982057 == array_index_948931 ? add_982353 : sel_982350;
  assign add_982357 = sel_982354 + 8'h01;
  assign sel_982358 = array_index_982057 == array_index_948937 ? add_982357 : sel_982354;
  assign add_982361 = sel_982358 + 8'h01;
  assign sel_982362 = array_index_982057 == array_index_948943 ? add_982361 : sel_982358;
  assign add_982365 = sel_982362 + 8'h01;
  assign sel_982366 = array_index_982057 == array_index_948949 ? add_982365 : sel_982362;
  assign add_982369 = sel_982366 + 8'h01;
  assign sel_982370 = array_index_982057 == array_index_948955 ? add_982369 : sel_982366;
  assign add_982373 = sel_982370 + 8'h01;
  assign sel_982374 = array_index_982057 == array_index_948961 ? add_982373 : sel_982370;
  assign add_982377 = sel_982374 + 8'h01;
  assign sel_982378 = array_index_982057 == array_index_948967 ? add_982377 : sel_982374;
  assign add_982381 = sel_982378 + 8'h01;
  assign sel_982382 = array_index_982057 == array_index_948973 ? add_982381 : sel_982378;
  assign add_982385 = sel_982382 + 8'h01;
  assign sel_982386 = array_index_982057 == array_index_948979 ? add_982385 : sel_982382;
  assign add_982389 = sel_982386 + 8'h01;
  assign sel_982390 = array_index_982057 == array_index_948985 ? add_982389 : sel_982386;
  assign add_982393 = sel_982390 + 8'h01;
  assign sel_982394 = array_index_982057 == array_index_948991 ? add_982393 : sel_982390;
  assign add_982397 = sel_982394 + 8'h01;
  assign sel_982398 = array_index_982057 == array_index_948997 ? add_982397 : sel_982394;
  assign add_982401 = sel_982398 + 8'h01;
  assign sel_982402 = array_index_982057 == array_index_949003 ? add_982401 : sel_982398;
  assign add_982405 = sel_982402 + 8'h01;
  assign sel_982406 = array_index_982057 == array_index_949009 ? add_982405 : sel_982402;
  assign add_982409 = sel_982406 + 8'h01;
  assign sel_982410 = array_index_982057 == array_index_949015 ? add_982409 : sel_982406;
  assign add_982413 = sel_982410 + 8'h01;
  assign sel_982414 = array_index_982057 == array_index_949021 ? add_982413 : sel_982410;
  assign add_982417 = sel_982414 + 8'h01;
  assign sel_982418 = array_index_982057 == array_index_949027 ? add_982417 : sel_982414;
  assign add_982421 = sel_982418 + 8'h01;
  assign sel_982422 = array_index_982057 == array_index_949033 ? add_982421 : sel_982418;
  assign add_982425 = sel_982422 + 8'h01;
  assign sel_982426 = array_index_982057 == array_index_949039 ? add_982425 : sel_982422;
  assign add_982429 = sel_982426 + 8'h01;
  assign sel_982430 = array_index_982057 == array_index_949045 ? add_982429 : sel_982426;
  assign add_982433 = sel_982430 + 8'h01;
  assign sel_982434 = array_index_982057 == array_index_949051 ? add_982433 : sel_982430;
  assign add_982437 = sel_982434 + 8'h01;
  assign sel_982438 = array_index_982057 == array_index_949057 ? add_982437 : sel_982434;
  assign add_982441 = sel_982438 + 8'h01;
  assign sel_982442 = array_index_982057 == array_index_949063 ? add_982441 : sel_982438;
  assign add_982445 = sel_982442 + 8'h01;
  assign sel_982446 = array_index_982057 == array_index_949069 ? add_982445 : sel_982442;
  assign add_982449 = sel_982446 + 8'h01;
  assign sel_982450 = array_index_982057 == array_index_949075 ? add_982449 : sel_982446;
  assign add_982453 = sel_982450 + 8'h01;
  assign sel_982454 = array_index_982057 == array_index_949081 ? add_982453 : sel_982450;
  assign add_982458 = sel_982454 + 8'h01;
  assign array_index_982459 = set1_unflattened[7'h54];
  assign sel_982460 = array_index_982057 == array_index_949087 ? add_982458 : sel_982454;
  assign add_982463 = sel_982460 + 8'h01;
  assign sel_982464 = array_index_982459 == array_index_948483 ? add_982463 : sel_982460;
  assign add_982467 = sel_982464 + 8'h01;
  assign sel_982468 = array_index_982459 == array_index_948487 ? add_982467 : sel_982464;
  assign add_982471 = sel_982468 + 8'h01;
  assign sel_982472 = array_index_982459 == array_index_948495 ? add_982471 : sel_982468;
  assign add_982475 = sel_982472 + 8'h01;
  assign sel_982476 = array_index_982459 == array_index_948503 ? add_982475 : sel_982472;
  assign add_982479 = sel_982476 + 8'h01;
  assign sel_982480 = array_index_982459 == array_index_948511 ? add_982479 : sel_982476;
  assign add_982483 = sel_982480 + 8'h01;
  assign sel_982484 = array_index_982459 == array_index_948519 ? add_982483 : sel_982480;
  assign add_982487 = sel_982484 + 8'h01;
  assign sel_982488 = array_index_982459 == array_index_948527 ? add_982487 : sel_982484;
  assign add_982491 = sel_982488 + 8'h01;
  assign sel_982492 = array_index_982459 == array_index_948535 ? add_982491 : sel_982488;
  assign add_982495 = sel_982492 + 8'h01;
  assign sel_982496 = array_index_982459 == array_index_948541 ? add_982495 : sel_982492;
  assign add_982499 = sel_982496 + 8'h01;
  assign sel_982500 = array_index_982459 == array_index_948547 ? add_982499 : sel_982496;
  assign add_982503 = sel_982500 + 8'h01;
  assign sel_982504 = array_index_982459 == array_index_948553 ? add_982503 : sel_982500;
  assign add_982507 = sel_982504 + 8'h01;
  assign sel_982508 = array_index_982459 == array_index_948559 ? add_982507 : sel_982504;
  assign add_982511 = sel_982508 + 8'h01;
  assign sel_982512 = array_index_982459 == array_index_948565 ? add_982511 : sel_982508;
  assign add_982515 = sel_982512 + 8'h01;
  assign sel_982516 = array_index_982459 == array_index_948571 ? add_982515 : sel_982512;
  assign add_982519 = sel_982516 + 8'h01;
  assign sel_982520 = array_index_982459 == array_index_948577 ? add_982519 : sel_982516;
  assign add_982523 = sel_982520 + 8'h01;
  assign sel_982524 = array_index_982459 == array_index_948583 ? add_982523 : sel_982520;
  assign add_982527 = sel_982524 + 8'h01;
  assign sel_982528 = array_index_982459 == array_index_948589 ? add_982527 : sel_982524;
  assign add_982531 = sel_982528 + 8'h01;
  assign sel_982532 = array_index_982459 == array_index_948595 ? add_982531 : sel_982528;
  assign add_982535 = sel_982532 + 8'h01;
  assign sel_982536 = array_index_982459 == array_index_948601 ? add_982535 : sel_982532;
  assign add_982539 = sel_982536 + 8'h01;
  assign sel_982540 = array_index_982459 == array_index_948607 ? add_982539 : sel_982536;
  assign add_982543 = sel_982540 + 8'h01;
  assign sel_982544 = array_index_982459 == array_index_948613 ? add_982543 : sel_982540;
  assign add_982547 = sel_982544 + 8'h01;
  assign sel_982548 = array_index_982459 == array_index_948619 ? add_982547 : sel_982544;
  assign add_982551 = sel_982548 + 8'h01;
  assign sel_982552 = array_index_982459 == array_index_948625 ? add_982551 : sel_982548;
  assign add_982555 = sel_982552 + 8'h01;
  assign sel_982556 = array_index_982459 == array_index_948631 ? add_982555 : sel_982552;
  assign add_982559 = sel_982556 + 8'h01;
  assign sel_982560 = array_index_982459 == array_index_948637 ? add_982559 : sel_982556;
  assign add_982563 = sel_982560 + 8'h01;
  assign sel_982564 = array_index_982459 == array_index_948643 ? add_982563 : sel_982560;
  assign add_982567 = sel_982564 + 8'h01;
  assign sel_982568 = array_index_982459 == array_index_948649 ? add_982567 : sel_982564;
  assign add_982571 = sel_982568 + 8'h01;
  assign sel_982572 = array_index_982459 == array_index_948655 ? add_982571 : sel_982568;
  assign add_982575 = sel_982572 + 8'h01;
  assign sel_982576 = array_index_982459 == array_index_948661 ? add_982575 : sel_982572;
  assign add_982579 = sel_982576 + 8'h01;
  assign sel_982580 = array_index_982459 == array_index_948667 ? add_982579 : sel_982576;
  assign add_982583 = sel_982580 + 8'h01;
  assign sel_982584 = array_index_982459 == array_index_948673 ? add_982583 : sel_982580;
  assign add_982587 = sel_982584 + 8'h01;
  assign sel_982588 = array_index_982459 == array_index_948679 ? add_982587 : sel_982584;
  assign add_982591 = sel_982588 + 8'h01;
  assign sel_982592 = array_index_982459 == array_index_948685 ? add_982591 : sel_982588;
  assign add_982595 = sel_982592 + 8'h01;
  assign sel_982596 = array_index_982459 == array_index_948691 ? add_982595 : sel_982592;
  assign add_982599 = sel_982596 + 8'h01;
  assign sel_982600 = array_index_982459 == array_index_948697 ? add_982599 : sel_982596;
  assign add_982603 = sel_982600 + 8'h01;
  assign sel_982604 = array_index_982459 == array_index_948703 ? add_982603 : sel_982600;
  assign add_982607 = sel_982604 + 8'h01;
  assign sel_982608 = array_index_982459 == array_index_948709 ? add_982607 : sel_982604;
  assign add_982611 = sel_982608 + 8'h01;
  assign sel_982612 = array_index_982459 == array_index_948715 ? add_982611 : sel_982608;
  assign add_982615 = sel_982612 + 8'h01;
  assign sel_982616 = array_index_982459 == array_index_948721 ? add_982615 : sel_982612;
  assign add_982619 = sel_982616 + 8'h01;
  assign sel_982620 = array_index_982459 == array_index_948727 ? add_982619 : sel_982616;
  assign add_982623 = sel_982620 + 8'h01;
  assign sel_982624 = array_index_982459 == array_index_948733 ? add_982623 : sel_982620;
  assign add_982627 = sel_982624 + 8'h01;
  assign sel_982628 = array_index_982459 == array_index_948739 ? add_982627 : sel_982624;
  assign add_982631 = sel_982628 + 8'h01;
  assign sel_982632 = array_index_982459 == array_index_948745 ? add_982631 : sel_982628;
  assign add_982635 = sel_982632 + 8'h01;
  assign sel_982636 = array_index_982459 == array_index_948751 ? add_982635 : sel_982632;
  assign add_982639 = sel_982636 + 8'h01;
  assign sel_982640 = array_index_982459 == array_index_948757 ? add_982639 : sel_982636;
  assign add_982643 = sel_982640 + 8'h01;
  assign sel_982644 = array_index_982459 == array_index_948763 ? add_982643 : sel_982640;
  assign add_982647 = sel_982644 + 8'h01;
  assign sel_982648 = array_index_982459 == array_index_948769 ? add_982647 : sel_982644;
  assign add_982651 = sel_982648 + 8'h01;
  assign sel_982652 = array_index_982459 == array_index_948775 ? add_982651 : sel_982648;
  assign add_982655 = sel_982652 + 8'h01;
  assign sel_982656 = array_index_982459 == array_index_948781 ? add_982655 : sel_982652;
  assign add_982659 = sel_982656 + 8'h01;
  assign sel_982660 = array_index_982459 == array_index_948787 ? add_982659 : sel_982656;
  assign add_982663 = sel_982660 + 8'h01;
  assign sel_982664 = array_index_982459 == array_index_948793 ? add_982663 : sel_982660;
  assign add_982667 = sel_982664 + 8'h01;
  assign sel_982668 = array_index_982459 == array_index_948799 ? add_982667 : sel_982664;
  assign add_982671 = sel_982668 + 8'h01;
  assign sel_982672 = array_index_982459 == array_index_948805 ? add_982671 : sel_982668;
  assign add_982675 = sel_982672 + 8'h01;
  assign sel_982676 = array_index_982459 == array_index_948811 ? add_982675 : sel_982672;
  assign add_982679 = sel_982676 + 8'h01;
  assign sel_982680 = array_index_982459 == array_index_948817 ? add_982679 : sel_982676;
  assign add_982683 = sel_982680 + 8'h01;
  assign sel_982684 = array_index_982459 == array_index_948823 ? add_982683 : sel_982680;
  assign add_982687 = sel_982684 + 8'h01;
  assign sel_982688 = array_index_982459 == array_index_948829 ? add_982687 : sel_982684;
  assign add_982691 = sel_982688 + 8'h01;
  assign sel_982692 = array_index_982459 == array_index_948835 ? add_982691 : sel_982688;
  assign add_982695 = sel_982692 + 8'h01;
  assign sel_982696 = array_index_982459 == array_index_948841 ? add_982695 : sel_982692;
  assign add_982699 = sel_982696 + 8'h01;
  assign sel_982700 = array_index_982459 == array_index_948847 ? add_982699 : sel_982696;
  assign add_982703 = sel_982700 + 8'h01;
  assign sel_982704 = array_index_982459 == array_index_948853 ? add_982703 : sel_982700;
  assign add_982707 = sel_982704 + 8'h01;
  assign sel_982708 = array_index_982459 == array_index_948859 ? add_982707 : sel_982704;
  assign add_982711 = sel_982708 + 8'h01;
  assign sel_982712 = array_index_982459 == array_index_948865 ? add_982711 : sel_982708;
  assign add_982715 = sel_982712 + 8'h01;
  assign sel_982716 = array_index_982459 == array_index_948871 ? add_982715 : sel_982712;
  assign add_982719 = sel_982716 + 8'h01;
  assign sel_982720 = array_index_982459 == array_index_948877 ? add_982719 : sel_982716;
  assign add_982723 = sel_982720 + 8'h01;
  assign sel_982724 = array_index_982459 == array_index_948883 ? add_982723 : sel_982720;
  assign add_982727 = sel_982724 + 8'h01;
  assign sel_982728 = array_index_982459 == array_index_948889 ? add_982727 : sel_982724;
  assign add_982731 = sel_982728 + 8'h01;
  assign sel_982732 = array_index_982459 == array_index_948895 ? add_982731 : sel_982728;
  assign add_982735 = sel_982732 + 8'h01;
  assign sel_982736 = array_index_982459 == array_index_948901 ? add_982735 : sel_982732;
  assign add_982739 = sel_982736 + 8'h01;
  assign sel_982740 = array_index_982459 == array_index_948907 ? add_982739 : sel_982736;
  assign add_982743 = sel_982740 + 8'h01;
  assign sel_982744 = array_index_982459 == array_index_948913 ? add_982743 : sel_982740;
  assign add_982747 = sel_982744 + 8'h01;
  assign sel_982748 = array_index_982459 == array_index_948919 ? add_982747 : sel_982744;
  assign add_982751 = sel_982748 + 8'h01;
  assign sel_982752 = array_index_982459 == array_index_948925 ? add_982751 : sel_982748;
  assign add_982755 = sel_982752 + 8'h01;
  assign sel_982756 = array_index_982459 == array_index_948931 ? add_982755 : sel_982752;
  assign add_982759 = sel_982756 + 8'h01;
  assign sel_982760 = array_index_982459 == array_index_948937 ? add_982759 : sel_982756;
  assign add_982763 = sel_982760 + 8'h01;
  assign sel_982764 = array_index_982459 == array_index_948943 ? add_982763 : sel_982760;
  assign add_982767 = sel_982764 + 8'h01;
  assign sel_982768 = array_index_982459 == array_index_948949 ? add_982767 : sel_982764;
  assign add_982771 = sel_982768 + 8'h01;
  assign sel_982772 = array_index_982459 == array_index_948955 ? add_982771 : sel_982768;
  assign add_982775 = sel_982772 + 8'h01;
  assign sel_982776 = array_index_982459 == array_index_948961 ? add_982775 : sel_982772;
  assign add_982779 = sel_982776 + 8'h01;
  assign sel_982780 = array_index_982459 == array_index_948967 ? add_982779 : sel_982776;
  assign add_982783 = sel_982780 + 8'h01;
  assign sel_982784 = array_index_982459 == array_index_948973 ? add_982783 : sel_982780;
  assign add_982787 = sel_982784 + 8'h01;
  assign sel_982788 = array_index_982459 == array_index_948979 ? add_982787 : sel_982784;
  assign add_982791 = sel_982788 + 8'h01;
  assign sel_982792 = array_index_982459 == array_index_948985 ? add_982791 : sel_982788;
  assign add_982795 = sel_982792 + 8'h01;
  assign sel_982796 = array_index_982459 == array_index_948991 ? add_982795 : sel_982792;
  assign add_982799 = sel_982796 + 8'h01;
  assign sel_982800 = array_index_982459 == array_index_948997 ? add_982799 : sel_982796;
  assign add_982803 = sel_982800 + 8'h01;
  assign sel_982804 = array_index_982459 == array_index_949003 ? add_982803 : sel_982800;
  assign add_982807 = sel_982804 + 8'h01;
  assign sel_982808 = array_index_982459 == array_index_949009 ? add_982807 : sel_982804;
  assign add_982811 = sel_982808 + 8'h01;
  assign sel_982812 = array_index_982459 == array_index_949015 ? add_982811 : sel_982808;
  assign add_982815 = sel_982812 + 8'h01;
  assign sel_982816 = array_index_982459 == array_index_949021 ? add_982815 : sel_982812;
  assign add_982819 = sel_982816 + 8'h01;
  assign sel_982820 = array_index_982459 == array_index_949027 ? add_982819 : sel_982816;
  assign add_982823 = sel_982820 + 8'h01;
  assign sel_982824 = array_index_982459 == array_index_949033 ? add_982823 : sel_982820;
  assign add_982827 = sel_982824 + 8'h01;
  assign sel_982828 = array_index_982459 == array_index_949039 ? add_982827 : sel_982824;
  assign add_982831 = sel_982828 + 8'h01;
  assign sel_982832 = array_index_982459 == array_index_949045 ? add_982831 : sel_982828;
  assign add_982835 = sel_982832 + 8'h01;
  assign sel_982836 = array_index_982459 == array_index_949051 ? add_982835 : sel_982832;
  assign add_982839 = sel_982836 + 8'h01;
  assign sel_982840 = array_index_982459 == array_index_949057 ? add_982839 : sel_982836;
  assign add_982843 = sel_982840 + 8'h01;
  assign sel_982844 = array_index_982459 == array_index_949063 ? add_982843 : sel_982840;
  assign add_982847 = sel_982844 + 8'h01;
  assign sel_982848 = array_index_982459 == array_index_949069 ? add_982847 : sel_982844;
  assign add_982851 = sel_982848 + 8'h01;
  assign sel_982852 = array_index_982459 == array_index_949075 ? add_982851 : sel_982848;
  assign add_982855 = sel_982852 + 8'h01;
  assign sel_982856 = array_index_982459 == array_index_949081 ? add_982855 : sel_982852;
  assign add_982860 = sel_982856 + 8'h01;
  assign array_index_982861 = set1_unflattened[7'h55];
  assign sel_982862 = array_index_982459 == array_index_949087 ? add_982860 : sel_982856;
  assign add_982865 = sel_982862 + 8'h01;
  assign sel_982866 = array_index_982861 == array_index_948483 ? add_982865 : sel_982862;
  assign add_982869 = sel_982866 + 8'h01;
  assign sel_982870 = array_index_982861 == array_index_948487 ? add_982869 : sel_982866;
  assign add_982873 = sel_982870 + 8'h01;
  assign sel_982874 = array_index_982861 == array_index_948495 ? add_982873 : sel_982870;
  assign add_982877 = sel_982874 + 8'h01;
  assign sel_982878 = array_index_982861 == array_index_948503 ? add_982877 : sel_982874;
  assign add_982881 = sel_982878 + 8'h01;
  assign sel_982882 = array_index_982861 == array_index_948511 ? add_982881 : sel_982878;
  assign add_982885 = sel_982882 + 8'h01;
  assign sel_982886 = array_index_982861 == array_index_948519 ? add_982885 : sel_982882;
  assign add_982889 = sel_982886 + 8'h01;
  assign sel_982890 = array_index_982861 == array_index_948527 ? add_982889 : sel_982886;
  assign add_982893 = sel_982890 + 8'h01;
  assign sel_982894 = array_index_982861 == array_index_948535 ? add_982893 : sel_982890;
  assign add_982897 = sel_982894 + 8'h01;
  assign sel_982898 = array_index_982861 == array_index_948541 ? add_982897 : sel_982894;
  assign add_982901 = sel_982898 + 8'h01;
  assign sel_982902 = array_index_982861 == array_index_948547 ? add_982901 : sel_982898;
  assign add_982905 = sel_982902 + 8'h01;
  assign sel_982906 = array_index_982861 == array_index_948553 ? add_982905 : sel_982902;
  assign add_982909 = sel_982906 + 8'h01;
  assign sel_982910 = array_index_982861 == array_index_948559 ? add_982909 : sel_982906;
  assign add_982913 = sel_982910 + 8'h01;
  assign sel_982914 = array_index_982861 == array_index_948565 ? add_982913 : sel_982910;
  assign add_982917 = sel_982914 + 8'h01;
  assign sel_982918 = array_index_982861 == array_index_948571 ? add_982917 : sel_982914;
  assign add_982921 = sel_982918 + 8'h01;
  assign sel_982922 = array_index_982861 == array_index_948577 ? add_982921 : sel_982918;
  assign add_982925 = sel_982922 + 8'h01;
  assign sel_982926 = array_index_982861 == array_index_948583 ? add_982925 : sel_982922;
  assign add_982929 = sel_982926 + 8'h01;
  assign sel_982930 = array_index_982861 == array_index_948589 ? add_982929 : sel_982926;
  assign add_982933 = sel_982930 + 8'h01;
  assign sel_982934 = array_index_982861 == array_index_948595 ? add_982933 : sel_982930;
  assign add_982937 = sel_982934 + 8'h01;
  assign sel_982938 = array_index_982861 == array_index_948601 ? add_982937 : sel_982934;
  assign add_982941 = sel_982938 + 8'h01;
  assign sel_982942 = array_index_982861 == array_index_948607 ? add_982941 : sel_982938;
  assign add_982945 = sel_982942 + 8'h01;
  assign sel_982946 = array_index_982861 == array_index_948613 ? add_982945 : sel_982942;
  assign add_982949 = sel_982946 + 8'h01;
  assign sel_982950 = array_index_982861 == array_index_948619 ? add_982949 : sel_982946;
  assign add_982953 = sel_982950 + 8'h01;
  assign sel_982954 = array_index_982861 == array_index_948625 ? add_982953 : sel_982950;
  assign add_982957 = sel_982954 + 8'h01;
  assign sel_982958 = array_index_982861 == array_index_948631 ? add_982957 : sel_982954;
  assign add_982961 = sel_982958 + 8'h01;
  assign sel_982962 = array_index_982861 == array_index_948637 ? add_982961 : sel_982958;
  assign add_982965 = sel_982962 + 8'h01;
  assign sel_982966 = array_index_982861 == array_index_948643 ? add_982965 : sel_982962;
  assign add_982969 = sel_982966 + 8'h01;
  assign sel_982970 = array_index_982861 == array_index_948649 ? add_982969 : sel_982966;
  assign add_982973 = sel_982970 + 8'h01;
  assign sel_982974 = array_index_982861 == array_index_948655 ? add_982973 : sel_982970;
  assign add_982977 = sel_982974 + 8'h01;
  assign sel_982978 = array_index_982861 == array_index_948661 ? add_982977 : sel_982974;
  assign add_982981 = sel_982978 + 8'h01;
  assign sel_982982 = array_index_982861 == array_index_948667 ? add_982981 : sel_982978;
  assign add_982985 = sel_982982 + 8'h01;
  assign sel_982986 = array_index_982861 == array_index_948673 ? add_982985 : sel_982982;
  assign add_982989 = sel_982986 + 8'h01;
  assign sel_982990 = array_index_982861 == array_index_948679 ? add_982989 : sel_982986;
  assign add_982993 = sel_982990 + 8'h01;
  assign sel_982994 = array_index_982861 == array_index_948685 ? add_982993 : sel_982990;
  assign add_982997 = sel_982994 + 8'h01;
  assign sel_982998 = array_index_982861 == array_index_948691 ? add_982997 : sel_982994;
  assign add_983001 = sel_982998 + 8'h01;
  assign sel_983002 = array_index_982861 == array_index_948697 ? add_983001 : sel_982998;
  assign add_983005 = sel_983002 + 8'h01;
  assign sel_983006 = array_index_982861 == array_index_948703 ? add_983005 : sel_983002;
  assign add_983009 = sel_983006 + 8'h01;
  assign sel_983010 = array_index_982861 == array_index_948709 ? add_983009 : sel_983006;
  assign add_983013 = sel_983010 + 8'h01;
  assign sel_983014 = array_index_982861 == array_index_948715 ? add_983013 : sel_983010;
  assign add_983017 = sel_983014 + 8'h01;
  assign sel_983018 = array_index_982861 == array_index_948721 ? add_983017 : sel_983014;
  assign add_983021 = sel_983018 + 8'h01;
  assign sel_983022 = array_index_982861 == array_index_948727 ? add_983021 : sel_983018;
  assign add_983025 = sel_983022 + 8'h01;
  assign sel_983026 = array_index_982861 == array_index_948733 ? add_983025 : sel_983022;
  assign add_983029 = sel_983026 + 8'h01;
  assign sel_983030 = array_index_982861 == array_index_948739 ? add_983029 : sel_983026;
  assign add_983033 = sel_983030 + 8'h01;
  assign sel_983034 = array_index_982861 == array_index_948745 ? add_983033 : sel_983030;
  assign add_983037 = sel_983034 + 8'h01;
  assign sel_983038 = array_index_982861 == array_index_948751 ? add_983037 : sel_983034;
  assign add_983041 = sel_983038 + 8'h01;
  assign sel_983042 = array_index_982861 == array_index_948757 ? add_983041 : sel_983038;
  assign add_983045 = sel_983042 + 8'h01;
  assign sel_983046 = array_index_982861 == array_index_948763 ? add_983045 : sel_983042;
  assign add_983049 = sel_983046 + 8'h01;
  assign sel_983050 = array_index_982861 == array_index_948769 ? add_983049 : sel_983046;
  assign add_983053 = sel_983050 + 8'h01;
  assign sel_983054 = array_index_982861 == array_index_948775 ? add_983053 : sel_983050;
  assign add_983057 = sel_983054 + 8'h01;
  assign sel_983058 = array_index_982861 == array_index_948781 ? add_983057 : sel_983054;
  assign add_983061 = sel_983058 + 8'h01;
  assign sel_983062 = array_index_982861 == array_index_948787 ? add_983061 : sel_983058;
  assign add_983065 = sel_983062 + 8'h01;
  assign sel_983066 = array_index_982861 == array_index_948793 ? add_983065 : sel_983062;
  assign add_983069 = sel_983066 + 8'h01;
  assign sel_983070 = array_index_982861 == array_index_948799 ? add_983069 : sel_983066;
  assign add_983073 = sel_983070 + 8'h01;
  assign sel_983074 = array_index_982861 == array_index_948805 ? add_983073 : sel_983070;
  assign add_983077 = sel_983074 + 8'h01;
  assign sel_983078 = array_index_982861 == array_index_948811 ? add_983077 : sel_983074;
  assign add_983081 = sel_983078 + 8'h01;
  assign sel_983082 = array_index_982861 == array_index_948817 ? add_983081 : sel_983078;
  assign add_983085 = sel_983082 + 8'h01;
  assign sel_983086 = array_index_982861 == array_index_948823 ? add_983085 : sel_983082;
  assign add_983089 = sel_983086 + 8'h01;
  assign sel_983090 = array_index_982861 == array_index_948829 ? add_983089 : sel_983086;
  assign add_983093 = sel_983090 + 8'h01;
  assign sel_983094 = array_index_982861 == array_index_948835 ? add_983093 : sel_983090;
  assign add_983097 = sel_983094 + 8'h01;
  assign sel_983098 = array_index_982861 == array_index_948841 ? add_983097 : sel_983094;
  assign add_983101 = sel_983098 + 8'h01;
  assign sel_983102 = array_index_982861 == array_index_948847 ? add_983101 : sel_983098;
  assign add_983105 = sel_983102 + 8'h01;
  assign sel_983106 = array_index_982861 == array_index_948853 ? add_983105 : sel_983102;
  assign add_983109 = sel_983106 + 8'h01;
  assign sel_983110 = array_index_982861 == array_index_948859 ? add_983109 : sel_983106;
  assign add_983113 = sel_983110 + 8'h01;
  assign sel_983114 = array_index_982861 == array_index_948865 ? add_983113 : sel_983110;
  assign add_983117 = sel_983114 + 8'h01;
  assign sel_983118 = array_index_982861 == array_index_948871 ? add_983117 : sel_983114;
  assign add_983121 = sel_983118 + 8'h01;
  assign sel_983122 = array_index_982861 == array_index_948877 ? add_983121 : sel_983118;
  assign add_983125 = sel_983122 + 8'h01;
  assign sel_983126 = array_index_982861 == array_index_948883 ? add_983125 : sel_983122;
  assign add_983129 = sel_983126 + 8'h01;
  assign sel_983130 = array_index_982861 == array_index_948889 ? add_983129 : sel_983126;
  assign add_983133 = sel_983130 + 8'h01;
  assign sel_983134 = array_index_982861 == array_index_948895 ? add_983133 : sel_983130;
  assign add_983137 = sel_983134 + 8'h01;
  assign sel_983138 = array_index_982861 == array_index_948901 ? add_983137 : sel_983134;
  assign add_983141 = sel_983138 + 8'h01;
  assign sel_983142 = array_index_982861 == array_index_948907 ? add_983141 : sel_983138;
  assign add_983145 = sel_983142 + 8'h01;
  assign sel_983146 = array_index_982861 == array_index_948913 ? add_983145 : sel_983142;
  assign add_983149 = sel_983146 + 8'h01;
  assign sel_983150 = array_index_982861 == array_index_948919 ? add_983149 : sel_983146;
  assign add_983153 = sel_983150 + 8'h01;
  assign sel_983154 = array_index_982861 == array_index_948925 ? add_983153 : sel_983150;
  assign add_983157 = sel_983154 + 8'h01;
  assign sel_983158 = array_index_982861 == array_index_948931 ? add_983157 : sel_983154;
  assign add_983161 = sel_983158 + 8'h01;
  assign sel_983162 = array_index_982861 == array_index_948937 ? add_983161 : sel_983158;
  assign add_983165 = sel_983162 + 8'h01;
  assign sel_983166 = array_index_982861 == array_index_948943 ? add_983165 : sel_983162;
  assign add_983169 = sel_983166 + 8'h01;
  assign sel_983170 = array_index_982861 == array_index_948949 ? add_983169 : sel_983166;
  assign add_983173 = sel_983170 + 8'h01;
  assign sel_983174 = array_index_982861 == array_index_948955 ? add_983173 : sel_983170;
  assign add_983177 = sel_983174 + 8'h01;
  assign sel_983178 = array_index_982861 == array_index_948961 ? add_983177 : sel_983174;
  assign add_983181 = sel_983178 + 8'h01;
  assign sel_983182 = array_index_982861 == array_index_948967 ? add_983181 : sel_983178;
  assign add_983185 = sel_983182 + 8'h01;
  assign sel_983186 = array_index_982861 == array_index_948973 ? add_983185 : sel_983182;
  assign add_983189 = sel_983186 + 8'h01;
  assign sel_983190 = array_index_982861 == array_index_948979 ? add_983189 : sel_983186;
  assign add_983193 = sel_983190 + 8'h01;
  assign sel_983194 = array_index_982861 == array_index_948985 ? add_983193 : sel_983190;
  assign add_983197 = sel_983194 + 8'h01;
  assign sel_983198 = array_index_982861 == array_index_948991 ? add_983197 : sel_983194;
  assign add_983201 = sel_983198 + 8'h01;
  assign sel_983202 = array_index_982861 == array_index_948997 ? add_983201 : sel_983198;
  assign add_983205 = sel_983202 + 8'h01;
  assign sel_983206 = array_index_982861 == array_index_949003 ? add_983205 : sel_983202;
  assign add_983209 = sel_983206 + 8'h01;
  assign sel_983210 = array_index_982861 == array_index_949009 ? add_983209 : sel_983206;
  assign add_983213 = sel_983210 + 8'h01;
  assign sel_983214 = array_index_982861 == array_index_949015 ? add_983213 : sel_983210;
  assign add_983217 = sel_983214 + 8'h01;
  assign sel_983218 = array_index_982861 == array_index_949021 ? add_983217 : sel_983214;
  assign add_983221 = sel_983218 + 8'h01;
  assign sel_983222 = array_index_982861 == array_index_949027 ? add_983221 : sel_983218;
  assign add_983225 = sel_983222 + 8'h01;
  assign sel_983226 = array_index_982861 == array_index_949033 ? add_983225 : sel_983222;
  assign add_983229 = sel_983226 + 8'h01;
  assign sel_983230 = array_index_982861 == array_index_949039 ? add_983229 : sel_983226;
  assign add_983233 = sel_983230 + 8'h01;
  assign sel_983234 = array_index_982861 == array_index_949045 ? add_983233 : sel_983230;
  assign add_983237 = sel_983234 + 8'h01;
  assign sel_983238 = array_index_982861 == array_index_949051 ? add_983237 : sel_983234;
  assign add_983241 = sel_983238 + 8'h01;
  assign sel_983242 = array_index_982861 == array_index_949057 ? add_983241 : sel_983238;
  assign add_983245 = sel_983242 + 8'h01;
  assign sel_983246 = array_index_982861 == array_index_949063 ? add_983245 : sel_983242;
  assign add_983249 = sel_983246 + 8'h01;
  assign sel_983250 = array_index_982861 == array_index_949069 ? add_983249 : sel_983246;
  assign add_983253 = sel_983250 + 8'h01;
  assign sel_983254 = array_index_982861 == array_index_949075 ? add_983253 : sel_983250;
  assign add_983257 = sel_983254 + 8'h01;
  assign sel_983258 = array_index_982861 == array_index_949081 ? add_983257 : sel_983254;
  assign add_983262 = sel_983258 + 8'h01;
  assign array_index_983263 = set1_unflattened[7'h56];
  assign sel_983264 = array_index_982861 == array_index_949087 ? add_983262 : sel_983258;
  assign add_983267 = sel_983264 + 8'h01;
  assign sel_983268 = array_index_983263 == array_index_948483 ? add_983267 : sel_983264;
  assign add_983271 = sel_983268 + 8'h01;
  assign sel_983272 = array_index_983263 == array_index_948487 ? add_983271 : sel_983268;
  assign add_983275 = sel_983272 + 8'h01;
  assign sel_983276 = array_index_983263 == array_index_948495 ? add_983275 : sel_983272;
  assign add_983279 = sel_983276 + 8'h01;
  assign sel_983280 = array_index_983263 == array_index_948503 ? add_983279 : sel_983276;
  assign add_983283 = sel_983280 + 8'h01;
  assign sel_983284 = array_index_983263 == array_index_948511 ? add_983283 : sel_983280;
  assign add_983287 = sel_983284 + 8'h01;
  assign sel_983288 = array_index_983263 == array_index_948519 ? add_983287 : sel_983284;
  assign add_983291 = sel_983288 + 8'h01;
  assign sel_983292 = array_index_983263 == array_index_948527 ? add_983291 : sel_983288;
  assign add_983295 = sel_983292 + 8'h01;
  assign sel_983296 = array_index_983263 == array_index_948535 ? add_983295 : sel_983292;
  assign add_983299 = sel_983296 + 8'h01;
  assign sel_983300 = array_index_983263 == array_index_948541 ? add_983299 : sel_983296;
  assign add_983303 = sel_983300 + 8'h01;
  assign sel_983304 = array_index_983263 == array_index_948547 ? add_983303 : sel_983300;
  assign add_983307 = sel_983304 + 8'h01;
  assign sel_983308 = array_index_983263 == array_index_948553 ? add_983307 : sel_983304;
  assign add_983311 = sel_983308 + 8'h01;
  assign sel_983312 = array_index_983263 == array_index_948559 ? add_983311 : sel_983308;
  assign add_983315 = sel_983312 + 8'h01;
  assign sel_983316 = array_index_983263 == array_index_948565 ? add_983315 : sel_983312;
  assign add_983319 = sel_983316 + 8'h01;
  assign sel_983320 = array_index_983263 == array_index_948571 ? add_983319 : sel_983316;
  assign add_983323 = sel_983320 + 8'h01;
  assign sel_983324 = array_index_983263 == array_index_948577 ? add_983323 : sel_983320;
  assign add_983327 = sel_983324 + 8'h01;
  assign sel_983328 = array_index_983263 == array_index_948583 ? add_983327 : sel_983324;
  assign add_983331 = sel_983328 + 8'h01;
  assign sel_983332 = array_index_983263 == array_index_948589 ? add_983331 : sel_983328;
  assign add_983335 = sel_983332 + 8'h01;
  assign sel_983336 = array_index_983263 == array_index_948595 ? add_983335 : sel_983332;
  assign add_983339 = sel_983336 + 8'h01;
  assign sel_983340 = array_index_983263 == array_index_948601 ? add_983339 : sel_983336;
  assign add_983343 = sel_983340 + 8'h01;
  assign sel_983344 = array_index_983263 == array_index_948607 ? add_983343 : sel_983340;
  assign add_983347 = sel_983344 + 8'h01;
  assign sel_983348 = array_index_983263 == array_index_948613 ? add_983347 : sel_983344;
  assign add_983351 = sel_983348 + 8'h01;
  assign sel_983352 = array_index_983263 == array_index_948619 ? add_983351 : sel_983348;
  assign add_983355 = sel_983352 + 8'h01;
  assign sel_983356 = array_index_983263 == array_index_948625 ? add_983355 : sel_983352;
  assign add_983359 = sel_983356 + 8'h01;
  assign sel_983360 = array_index_983263 == array_index_948631 ? add_983359 : sel_983356;
  assign add_983363 = sel_983360 + 8'h01;
  assign sel_983364 = array_index_983263 == array_index_948637 ? add_983363 : sel_983360;
  assign add_983367 = sel_983364 + 8'h01;
  assign sel_983368 = array_index_983263 == array_index_948643 ? add_983367 : sel_983364;
  assign add_983371 = sel_983368 + 8'h01;
  assign sel_983372 = array_index_983263 == array_index_948649 ? add_983371 : sel_983368;
  assign add_983375 = sel_983372 + 8'h01;
  assign sel_983376 = array_index_983263 == array_index_948655 ? add_983375 : sel_983372;
  assign add_983379 = sel_983376 + 8'h01;
  assign sel_983380 = array_index_983263 == array_index_948661 ? add_983379 : sel_983376;
  assign add_983383 = sel_983380 + 8'h01;
  assign sel_983384 = array_index_983263 == array_index_948667 ? add_983383 : sel_983380;
  assign add_983387 = sel_983384 + 8'h01;
  assign sel_983388 = array_index_983263 == array_index_948673 ? add_983387 : sel_983384;
  assign add_983391 = sel_983388 + 8'h01;
  assign sel_983392 = array_index_983263 == array_index_948679 ? add_983391 : sel_983388;
  assign add_983395 = sel_983392 + 8'h01;
  assign sel_983396 = array_index_983263 == array_index_948685 ? add_983395 : sel_983392;
  assign add_983399 = sel_983396 + 8'h01;
  assign sel_983400 = array_index_983263 == array_index_948691 ? add_983399 : sel_983396;
  assign add_983403 = sel_983400 + 8'h01;
  assign sel_983404 = array_index_983263 == array_index_948697 ? add_983403 : sel_983400;
  assign add_983407 = sel_983404 + 8'h01;
  assign sel_983408 = array_index_983263 == array_index_948703 ? add_983407 : sel_983404;
  assign add_983411 = sel_983408 + 8'h01;
  assign sel_983412 = array_index_983263 == array_index_948709 ? add_983411 : sel_983408;
  assign add_983415 = sel_983412 + 8'h01;
  assign sel_983416 = array_index_983263 == array_index_948715 ? add_983415 : sel_983412;
  assign add_983419 = sel_983416 + 8'h01;
  assign sel_983420 = array_index_983263 == array_index_948721 ? add_983419 : sel_983416;
  assign add_983423 = sel_983420 + 8'h01;
  assign sel_983424 = array_index_983263 == array_index_948727 ? add_983423 : sel_983420;
  assign add_983427 = sel_983424 + 8'h01;
  assign sel_983428 = array_index_983263 == array_index_948733 ? add_983427 : sel_983424;
  assign add_983431 = sel_983428 + 8'h01;
  assign sel_983432 = array_index_983263 == array_index_948739 ? add_983431 : sel_983428;
  assign add_983435 = sel_983432 + 8'h01;
  assign sel_983436 = array_index_983263 == array_index_948745 ? add_983435 : sel_983432;
  assign add_983439 = sel_983436 + 8'h01;
  assign sel_983440 = array_index_983263 == array_index_948751 ? add_983439 : sel_983436;
  assign add_983443 = sel_983440 + 8'h01;
  assign sel_983444 = array_index_983263 == array_index_948757 ? add_983443 : sel_983440;
  assign add_983447 = sel_983444 + 8'h01;
  assign sel_983448 = array_index_983263 == array_index_948763 ? add_983447 : sel_983444;
  assign add_983451 = sel_983448 + 8'h01;
  assign sel_983452 = array_index_983263 == array_index_948769 ? add_983451 : sel_983448;
  assign add_983455 = sel_983452 + 8'h01;
  assign sel_983456 = array_index_983263 == array_index_948775 ? add_983455 : sel_983452;
  assign add_983459 = sel_983456 + 8'h01;
  assign sel_983460 = array_index_983263 == array_index_948781 ? add_983459 : sel_983456;
  assign add_983463 = sel_983460 + 8'h01;
  assign sel_983464 = array_index_983263 == array_index_948787 ? add_983463 : sel_983460;
  assign add_983467 = sel_983464 + 8'h01;
  assign sel_983468 = array_index_983263 == array_index_948793 ? add_983467 : sel_983464;
  assign add_983471 = sel_983468 + 8'h01;
  assign sel_983472 = array_index_983263 == array_index_948799 ? add_983471 : sel_983468;
  assign add_983475 = sel_983472 + 8'h01;
  assign sel_983476 = array_index_983263 == array_index_948805 ? add_983475 : sel_983472;
  assign add_983479 = sel_983476 + 8'h01;
  assign sel_983480 = array_index_983263 == array_index_948811 ? add_983479 : sel_983476;
  assign add_983483 = sel_983480 + 8'h01;
  assign sel_983484 = array_index_983263 == array_index_948817 ? add_983483 : sel_983480;
  assign add_983487 = sel_983484 + 8'h01;
  assign sel_983488 = array_index_983263 == array_index_948823 ? add_983487 : sel_983484;
  assign add_983491 = sel_983488 + 8'h01;
  assign sel_983492 = array_index_983263 == array_index_948829 ? add_983491 : sel_983488;
  assign add_983495 = sel_983492 + 8'h01;
  assign sel_983496 = array_index_983263 == array_index_948835 ? add_983495 : sel_983492;
  assign add_983499 = sel_983496 + 8'h01;
  assign sel_983500 = array_index_983263 == array_index_948841 ? add_983499 : sel_983496;
  assign add_983503 = sel_983500 + 8'h01;
  assign sel_983504 = array_index_983263 == array_index_948847 ? add_983503 : sel_983500;
  assign add_983507 = sel_983504 + 8'h01;
  assign sel_983508 = array_index_983263 == array_index_948853 ? add_983507 : sel_983504;
  assign add_983511 = sel_983508 + 8'h01;
  assign sel_983512 = array_index_983263 == array_index_948859 ? add_983511 : sel_983508;
  assign add_983515 = sel_983512 + 8'h01;
  assign sel_983516 = array_index_983263 == array_index_948865 ? add_983515 : sel_983512;
  assign add_983519 = sel_983516 + 8'h01;
  assign sel_983520 = array_index_983263 == array_index_948871 ? add_983519 : sel_983516;
  assign add_983523 = sel_983520 + 8'h01;
  assign sel_983524 = array_index_983263 == array_index_948877 ? add_983523 : sel_983520;
  assign add_983527 = sel_983524 + 8'h01;
  assign sel_983528 = array_index_983263 == array_index_948883 ? add_983527 : sel_983524;
  assign add_983531 = sel_983528 + 8'h01;
  assign sel_983532 = array_index_983263 == array_index_948889 ? add_983531 : sel_983528;
  assign add_983535 = sel_983532 + 8'h01;
  assign sel_983536 = array_index_983263 == array_index_948895 ? add_983535 : sel_983532;
  assign add_983539 = sel_983536 + 8'h01;
  assign sel_983540 = array_index_983263 == array_index_948901 ? add_983539 : sel_983536;
  assign add_983543 = sel_983540 + 8'h01;
  assign sel_983544 = array_index_983263 == array_index_948907 ? add_983543 : sel_983540;
  assign add_983547 = sel_983544 + 8'h01;
  assign sel_983548 = array_index_983263 == array_index_948913 ? add_983547 : sel_983544;
  assign add_983551 = sel_983548 + 8'h01;
  assign sel_983552 = array_index_983263 == array_index_948919 ? add_983551 : sel_983548;
  assign add_983555 = sel_983552 + 8'h01;
  assign sel_983556 = array_index_983263 == array_index_948925 ? add_983555 : sel_983552;
  assign add_983559 = sel_983556 + 8'h01;
  assign sel_983560 = array_index_983263 == array_index_948931 ? add_983559 : sel_983556;
  assign add_983563 = sel_983560 + 8'h01;
  assign sel_983564 = array_index_983263 == array_index_948937 ? add_983563 : sel_983560;
  assign add_983567 = sel_983564 + 8'h01;
  assign sel_983568 = array_index_983263 == array_index_948943 ? add_983567 : sel_983564;
  assign add_983571 = sel_983568 + 8'h01;
  assign sel_983572 = array_index_983263 == array_index_948949 ? add_983571 : sel_983568;
  assign add_983575 = sel_983572 + 8'h01;
  assign sel_983576 = array_index_983263 == array_index_948955 ? add_983575 : sel_983572;
  assign add_983579 = sel_983576 + 8'h01;
  assign sel_983580 = array_index_983263 == array_index_948961 ? add_983579 : sel_983576;
  assign add_983583 = sel_983580 + 8'h01;
  assign sel_983584 = array_index_983263 == array_index_948967 ? add_983583 : sel_983580;
  assign add_983587 = sel_983584 + 8'h01;
  assign sel_983588 = array_index_983263 == array_index_948973 ? add_983587 : sel_983584;
  assign add_983591 = sel_983588 + 8'h01;
  assign sel_983592 = array_index_983263 == array_index_948979 ? add_983591 : sel_983588;
  assign add_983595 = sel_983592 + 8'h01;
  assign sel_983596 = array_index_983263 == array_index_948985 ? add_983595 : sel_983592;
  assign add_983599 = sel_983596 + 8'h01;
  assign sel_983600 = array_index_983263 == array_index_948991 ? add_983599 : sel_983596;
  assign add_983603 = sel_983600 + 8'h01;
  assign sel_983604 = array_index_983263 == array_index_948997 ? add_983603 : sel_983600;
  assign add_983607 = sel_983604 + 8'h01;
  assign sel_983608 = array_index_983263 == array_index_949003 ? add_983607 : sel_983604;
  assign add_983611 = sel_983608 + 8'h01;
  assign sel_983612 = array_index_983263 == array_index_949009 ? add_983611 : sel_983608;
  assign add_983615 = sel_983612 + 8'h01;
  assign sel_983616 = array_index_983263 == array_index_949015 ? add_983615 : sel_983612;
  assign add_983619 = sel_983616 + 8'h01;
  assign sel_983620 = array_index_983263 == array_index_949021 ? add_983619 : sel_983616;
  assign add_983623 = sel_983620 + 8'h01;
  assign sel_983624 = array_index_983263 == array_index_949027 ? add_983623 : sel_983620;
  assign add_983627 = sel_983624 + 8'h01;
  assign sel_983628 = array_index_983263 == array_index_949033 ? add_983627 : sel_983624;
  assign add_983631 = sel_983628 + 8'h01;
  assign sel_983632 = array_index_983263 == array_index_949039 ? add_983631 : sel_983628;
  assign add_983635 = sel_983632 + 8'h01;
  assign sel_983636 = array_index_983263 == array_index_949045 ? add_983635 : sel_983632;
  assign add_983639 = sel_983636 + 8'h01;
  assign sel_983640 = array_index_983263 == array_index_949051 ? add_983639 : sel_983636;
  assign add_983643 = sel_983640 + 8'h01;
  assign sel_983644 = array_index_983263 == array_index_949057 ? add_983643 : sel_983640;
  assign add_983647 = sel_983644 + 8'h01;
  assign sel_983648 = array_index_983263 == array_index_949063 ? add_983647 : sel_983644;
  assign add_983651 = sel_983648 + 8'h01;
  assign sel_983652 = array_index_983263 == array_index_949069 ? add_983651 : sel_983648;
  assign add_983655 = sel_983652 + 8'h01;
  assign sel_983656 = array_index_983263 == array_index_949075 ? add_983655 : sel_983652;
  assign add_983659 = sel_983656 + 8'h01;
  assign sel_983660 = array_index_983263 == array_index_949081 ? add_983659 : sel_983656;
  assign add_983664 = sel_983660 + 8'h01;
  assign array_index_983665 = set1_unflattened[7'h57];
  assign sel_983666 = array_index_983263 == array_index_949087 ? add_983664 : sel_983660;
  assign add_983669 = sel_983666 + 8'h01;
  assign sel_983670 = array_index_983665 == array_index_948483 ? add_983669 : sel_983666;
  assign add_983673 = sel_983670 + 8'h01;
  assign sel_983674 = array_index_983665 == array_index_948487 ? add_983673 : sel_983670;
  assign add_983677 = sel_983674 + 8'h01;
  assign sel_983678 = array_index_983665 == array_index_948495 ? add_983677 : sel_983674;
  assign add_983681 = sel_983678 + 8'h01;
  assign sel_983682 = array_index_983665 == array_index_948503 ? add_983681 : sel_983678;
  assign add_983685 = sel_983682 + 8'h01;
  assign sel_983686 = array_index_983665 == array_index_948511 ? add_983685 : sel_983682;
  assign add_983689 = sel_983686 + 8'h01;
  assign sel_983690 = array_index_983665 == array_index_948519 ? add_983689 : sel_983686;
  assign add_983693 = sel_983690 + 8'h01;
  assign sel_983694 = array_index_983665 == array_index_948527 ? add_983693 : sel_983690;
  assign add_983697 = sel_983694 + 8'h01;
  assign sel_983698 = array_index_983665 == array_index_948535 ? add_983697 : sel_983694;
  assign add_983701 = sel_983698 + 8'h01;
  assign sel_983702 = array_index_983665 == array_index_948541 ? add_983701 : sel_983698;
  assign add_983705 = sel_983702 + 8'h01;
  assign sel_983706 = array_index_983665 == array_index_948547 ? add_983705 : sel_983702;
  assign add_983709 = sel_983706 + 8'h01;
  assign sel_983710 = array_index_983665 == array_index_948553 ? add_983709 : sel_983706;
  assign add_983713 = sel_983710 + 8'h01;
  assign sel_983714 = array_index_983665 == array_index_948559 ? add_983713 : sel_983710;
  assign add_983717 = sel_983714 + 8'h01;
  assign sel_983718 = array_index_983665 == array_index_948565 ? add_983717 : sel_983714;
  assign add_983721 = sel_983718 + 8'h01;
  assign sel_983722 = array_index_983665 == array_index_948571 ? add_983721 : sel_983718;
  assign add_983725 = sel_983722 + 8'h01;
  assign sel_983726 = array_index_983665 == array_index_948577 ? add_983725 : sel_983722;
  assign add_983729 = sel_983726 + 8'h01;
  assign sel_983730 = array_index_983665 == array_index_948583 ? add_983729 : sel_983726;
  assign add_983733 = sel_983730 + 8'h01;
  assign sel_983734 = array_index_983665 == array_index_948589 ? add_983733 : sel_983730;
  assign add_983737 = sel_983734 + 8'h01;
  assign sel_983738 = array_index_983665 == array_index_948595 ? add_983737 : sel_983734;
  assign add_983741 = sel_983738 + 8'h01;
  assign sel_983742 = array_index_983665 == array_index_948601 ? add_983741 : sel_983738;
  assign add_983745 = sel_983742 + 8'h01;
  assign sel_983746 = array_index_983665 == array_index_948607 ? add_983745 : sel_983742;
  assign add_983749 = sel_983746 + 8'h01;
  assign sel_983750 = array_index_983665 == array_index_948613 ? add_983749 : sel_983746;
  assign add_983753 = sel_983750 + 8'h01;
  assign sel_983754 = array_index_983665 == array_index_948619 ? add_983753 : sel_983750;
  assign add_983757 = sel_983754 + 8'h01;
  assign sel_983758 = array_index_983665 == array_index_948625 ? add_983757 : sel_983754;
  assign add_983761 = sel_983758 + 8'h01;
  assign sel_983762 = array_index_983665 == array_index_948631 ? add_983761 : sel_983758;
  assign add_983765 = sel_983762 + 8'h01;
  assign sel_983766 = array_index_983665 == array_index_948637 ? add_983765 : sel_983762;
  assign add_983769 = sel_983766 + 8'h01;
  assign sel_983770 = array_index_983665 == array_index_948643 ? add_983769 : sel_983766;
  assign add_983773 = sel_983770 + 8'h01;
  assign sel_983774 = array_index_983665 == array_index_948649 ? add_983773 : sel_983770;
  assign add_983777 = sel_983774 + 8'h01;
  assign sel_983778 = array_index_983665 == array_index_948655 ? add_983777 : sel_983774;
  assign add_983781 = sel_983778 + 8'h01;
  assign sel_983782 = array_index_983665 == array_index_948661 ? add_983781 : sel_983778;
  assign add_983785 = sel_983782 + 8'h01;
  assign sel_983786 = array_index_983665 == array_index_948667 ? add_983785 : sel_983782;
  assign add_983789 = sel_983786 + 8'h01;
  assign sel_983790 = array_index_983665 == array_index_948673 ? add_983789 : sel_983786;
  assign add_983793 = sel_983790 + 8'h01;
  assign sel_983794 = array_index_983665 == array_index_948679 ? add_983793 : sel_983790;
  assign add_983797 = sel_983794 + 8'h01;
  assign sel_983798 = array_index_983665 == array_index_948685 ? add_983797 : sel_983794;
  assign add_983801 = sel_983798 + 8'h01;
  assign sel_983802 = array_index_983665 == array_index_948691 ? add_983801 : sel_983798;
  assign add_983805 = sel_983802 + 8'h01;
  assign sel_983806 = array_index_983665 == array_index_948697 ? add_983805 : sel_983802;
  assign add_983809 = sel_983806 + 8'h01;
  assign sel_983810 = array_index_983665 == array_index_948703 ? add_983809 : sel_983806;
  assign add_983813 = sel_983810 + 8'h01;
  assign sel_983814 = array_index_983665 == array_index_948709 ? add_983813 : sel_983810;
  assign add_983817 = sel_983814 + 8'h01;
  assign sel_983818 = array_index_983665 == array_index_948715 ? add_983817 : sel_983814;
  assign add_983821 = sel_983818 + 8'h01;
  assign sel_983822 = array_index_983665 == array_index_948721 ? add_983821 : sel_983818;
  assign add_983825 = sel_983822 + 8'h01;
  assign sel_983826 = array_index_983665 == array_index_948727 ? add_983825 : sel_983822;
  assign add_983829 = sel_983826 + 8'h01;
  assign sel_983830 = array_index_983665 == array_index_948733 ? add_983829 : sel_983826;
  assign add_983833 = sel_983830 + 8'h01;
  assign sel_983834 = array_index_983665 == array_index_948739 ? add_983833 : sel_983830;
  assign add_983837 = sel_983834 + 8'h01;
  assign sel_983838 = array_index_983665 == array_index_948745 ? add_983837 : sel_983834;
  assign add_983841 = sel_983838 + 8'h01;
  assign sel_983842 = array_index_983665 == array_index_948751 ? add_983841 : sel_983838;
  assign add_983845 = sel_983842 + 8'h01;
  assign sel_983846 = array_index_983665 == array_index_948757 ? add_983845 : sel_983842;
  assign add_983849 = sel_983846 + 8'h01;
  assign sel_983850 = array_index_983665 == array_index_948763 ? add_983849 : sel_983846;
  assign add_983853 = sel_983850 + 8'h01;
  assign sel_983854 = array_index_983665 == array_index_948769 ? add_983853 : sel_983850;
  assign add_983857 = sel_983854 + 8'h01;
  assign sel_983858 = array_index_983665 == array_index_948775 ? add_983857 : sel_983854;
  assign add_983861 = sel_983858 + 8'h01;
  assign sel_983862 = array_index_983665 == array_index_948781 ? add_983861 : sel_983858;
  assign add_983865 = sel_983862 + 8'h01;
  assign sel_983866 = array_index_983665 == array_index_948787 ? add_983865 : sel_983862;
  assign add_983869 = sel_983866 + 8'h01;
  assign sel_983870 = array_index_983665 == array_index_948793 ? add_983869 : sel_983866;
  assign add_983873 = sel_983870 + 8'h01;
  assign sel_983874 = array_index_983665 == array_index_948799 ? add_983873 : sel_983870;
  assign add_983877 = sel_983874 + 8'h01;
  assign sel_983878 = array_index_983665 == array_index_948805 ? add_983877 : sel_983874;
  assign add_983881 = sel_983878 + 8'h01;
  assign sel_983882 = array_index_983665 == array_index_948811 ? add_983881 : sel_983878;
  assign add_983885 = sel_983882 + 8'h01;
  assign sel_983886 = array_index_983665 == array_index_948817 ? add_983885 : sel_983882;
  assign add_983889 = sel_983886 + 8'h01;
  assign sel_983890 = array_index_983665 == array_index_948823 ? add_983889 : sel_983886;
  assign add_983893 = sel_983890 + 8'h01;
  assign sel_983894 = array_index_983665 == array_index_948829 ? add_983893 : sel_983890;
  assign add_983897 = sel_983894 + 8'h01;
  assign sel_983898 = array_index_983665 == array_index_948835 ? add_983897 : sel_983894;
  assign add_983901 = sel_983898 + 8'h01;
  assign sel_983902 = array_index_983665 == array_index_948841 ? add_983901 : sel_983898;
  assign add_983905 = sel_983902 + 8'h01;
  assign sel_983906 = array_index_983665 == array_index_948847 ? add_983905 : sel_983902;
  assign add_983909 = sel_983906 + 8'h01;
  assign sel_983910 = array_index_983665 == array_index_948853 ? add_983909 : sel_983906;
  assign add_983913 = sel_983910 + 8'h01;
  assign sel_983914 = array_index_983665 == array_index_948859 ? add_983913 : sel_983910;
  assign add_983917 = sel_983914 + 8'h01;
  assign sel_983918 = array_index_983665 == array_index_948865 ? add_983917 : sel_983914;
  assign add_983921 = sel_983918 + 8'h01;
  assign sel_983922 = array_index_983665 == array_index_948871 ? add_983921 : sel_983918;
  assign add_983925 = sel_983922 + 8'h01;
  assign sel_983926 = array_index_983665 == array_index_948877 ? add_983925 : sel_983922;
  assign add_983929 = sel_983926 + 8'h01;
  assign sel_983930 = array_index_983665 == array_index_948883 ? add_983929 : sel_983926;
  assign add_983933 = sel_983930 + 8'h01;
  assign sel_983934 = array_index_983665 == array_index_948889 ? add_983933 : sel_983930;
  assign add_983937 = sel_983934 + 8'h01;
  assign sel_983938 = array_index_983665 == array_index_948895 ? add_983937 : sel_983934;
  assign add_983941 = sel_983938 + 8'h01;
  assign sel_983942 = array_index_983665 == array_index_948901 ? add_983941 : sel_983938;
  assign add_983945 = sel_983942 + 8'h01;
  assign sel_983946 = array_index_983665 == array_index_948907 ? add_983945 : sel_983942;
  assign add_983949 = sel_983946 + 8'h01;
  assign sel_983950 = array_index_983665 == array_index_948913 ? add_983949 : sel_983946;
  assign add_983953 = sel_983950 + 8'h01;
  assign sel_983954 = array_index_983665 == array_index_948919 ? add_983953 : sel_983950;
  assign add_983957 = sel_983954 + 8'h01;
  assign sel_983958 = array_index_983665 == array_index_948925 ? add_983957 : sel_983954;
  assign add_983961 = sel_983958 + 8'h01;
  assign sel_983962 = array_index_983665 == array_index_948931 ? add_983961 : sel_983958;
  assign add_983965 = sel_983962 + 8'h01;
  assign sel_983966 = array_index_983665 == array_index_948937 ? add_983965 : sel_983962;
  assign add_983969 = sel_983966 + 8'h01;
  assign sel_983970 = array_index_983665 == array_index_948943 ? add_983969 : sel_983966;
  assign add_983973 = sel_983970 + 8'h01;
  assign sel_983974 = array_index_983665 == array_index_948949 ? add_983973 : sel_983970;
  assign add_983977 = sel_983974 + 8'h01;
  assign sel_983978 = array_index_983665 == array_index_948955 ? add_983977 : sel_983974;
  assign add_983981 = sel_983978 + 8'h01;
  assign sel_983982 = array_index_983665 == array_index_948961 ? add_983981 : sel_983978;
  assign add_983985 = sel_983982 + 8'h01;
  assign sel_983986 = array_index_983665 == array_index_948967 ? add_983985 : sel_983982;
  assign add_983989 = sel_983986 + 8'h01;
  assign sel_983990 = array_index_983665 == array_index_948973 ? add_983989 : sel_983986;
  assign add_983993 = sel_983990 + 8'h01;
  assign sel_983994 = array_index_983665 == array_index_948979 ? add_983993 : sel_983990;
  assign add_983997 = sel_983994 + 8'h01;
  assign sel_983998 = array_index_983665 == array_index_948985 ? add_983997 : sel_983994;
  assign add_984001 = sel_983998 + 8'h01;
  assign sel_984002 = array_index_983665 == array_index_948991 ? add_984001 : sel_983998;
  assign add_984005 = sel_984002 + 8'h01;
  assign sel_984006 = array_index_983665 == array_index_948997 ? add_984005 : sel_984002;
  assign add_984009 = sel_984006 + 8'h01;
  assign sel_984010 = array_index_983665 == array_index_949003 ? add_984009 : sel_984006;
  assign add_984013 = sel_984010 + 8'h01;
  assign sel_984014 = array_index_983665 == array_index_949009 ? add_984013 : sel_984010;
  assign add_984017 = sel_984014 + 8'h01;
  assign sel_984018 = array_index_983665 == array_index_949015 ? add_984017 : sel_984014;
  assign add_984021 = sel_984018 + 8'h01;
  assign sel_984022 = array_index_983665 == array_index_949021 ? add_984021 : sel_984018;
  assign add_984025 = sel_984022 + 8'h01;
  assign sel_984026 = array_index_983665 == array_index_949027 ? add_984025 : sel_984022;
  assign add_984029 = sel_984026 + 8'h01;
  assign sel_984030 = array_index_983665 == array_index_949033 ? add_984029 : sel_984026;
  assign add_984033 = sel_984030 + 8'h01;
  assign sel_984034 = array_index_983665 == array_index_949039 ? add_984033 : sel_984030;
  assign add_984037 = sel_984034 + 8'h01;
  assign sel_984038 = array_index_983665 == array_index_949045 ? add_984037 : sel_984034;
  assign add_984041 = sel_984038 + 8'h01;
  assign sel_984042 = array_index_983665 == array_index_949051 ? add_984041 : sel_984038;
  assign add_984045 = sel_984042 + 8'h01;
  assign sel_984046 = array_index_983665 == array_index_949057 ? add_984045 : sel_984042;
  assign add_984049 = sel_984046 + 8'h01;
  assign sel_984050 = array_index_983665 == array_index_949063 ? add_984049 : sel_984046;
  assign add_984053 = sel_984050 + 8'h01;
  assign sel_984054 = array_index_983665 == array_index_949069 ? add_984053 : sel_984050;
  assign add_984057 = sel_984054 + 8'h01;
  assign sel_984058 = array_index_983665 == array_index_949075 ? add_984057 : sel_984054;
  assign add_984061 = sel_984058 + 8'h01;
  assign sel_984062 = array_index_983665 == array_index_949081 ? add_984061 : sel_984058;
  assign add_984066 = sel_984062 + 8'h01;
  assign array_index_984067 = set1_unflattened[7'h58];
  assign sel_984068 = array_index_983665 == array_index_949087 ? add_984066 : sel_984062;
  assign add_984071 = sel_984068 + 8'h01;
  assign sel_984072 = array_index_984067 == array_index_948483 ? add_984071 : sel_984068;
  assign add_984075 = sel_984072 + 8'h01;
  assign sel_984076 = array_index_984067 == array_index_948487 ? add_984075 : sel_984072;
  assign add_984079 = sel_984076 + 8'h01;
  assign sel_984080 = array_index_984067 == array_index_948495 ? add_984079 : sel_984076;
  assign add_984083 = sel_984080 + 8'h01;
  assign sel_984084 = array_index_984067 == array_index_948503 ? add_984083 : sel_984080;
  assign add_984087 = sel_984084 + 8'h01;
  assign sel_984088 = array_index_984067 == array_index_948511 ? add_984087 : sel_984084;
  assign add_984091 = sel_984088 + 8'h01;
  assign sel_984092 = array_index_984067 == array_index_948519 ? add_984091 : sel_984088;
  assign add_984095 = sel_984092 + 8'h01;
  assign sel_984096 = array_index_984067 == array_index_948527 ? add_984095 : sel_984092;
  assign add_984099 = sel_984096 + 8'h01;
  assign sel_984100 = array_index_984067 == array_index_948535 ? add_984099 : sel_984096;
  assign add_984103 = sel_984100 + 8'h01;
  assign sel_984104 = array_index_984067 == array_index_948541 ? add_984103 : sel_984100;
  assign add_984107 = sel_984104 + 8'h01;
  assign sel_984108 = array_index_984067 == array_index_948547 ? add_984107 : sel_984104;
  assign add_984111 = sel_984108 + 8'h01;
  assign sel_984112 = array_index_984067 == array_index_948553 ? add_984111 : sel_984108;
  assign add_984115 = sel_984112 + 8'h01;
  assign sel_984116 = array_index_984067 == array_index_948559 ? add_984115 : sel_984112;
  assign add_984119 = sel_984116 + 8'h01;
  assign sel_984120 = array_index_984067 == array_index_948565 ? add_984119 : sel_984116;
  assign add_984123 = sel_984120 + 8'h01;
  assign sel_984124 = array_index_984067 == array_index_948571 ? add_984123 : sel_984120;
  assign add_984127 = sel_984124 + 8'h01;
  assign sel_984128 = array_index_984067 == array_index_948577 ? add_984127 : sel_984124;
  assign add_984131 = sel_984128 + 8'h01;
  assign sel_984132 = array_index_984067 == array_index_948583 ? add_984131 : sel_984128;
  assign add_984135 = sel_984132 + 8'h01;
  assign sel_984136 = array_index_984067 == array_index_948589 ? add_984135 : sel_984132;
  assign add_984139 = sel_984136 + 8'h01;
  assign sel_984140 = array_index_984067 == array_index_948595 ? add_984139 : sel_984136;
  assign add_984143 = sel_984140 + 8'h01;
  assign sel_984144 = array_index_984067 == array_index_948601 ? add_984143 : sel_984140;
  assign add_984147 = sel_984144 + 8'h01;
  assign sel_984148 = array_index_984067 == array_index_948607 ? add_984147 : sel_984144;
  assign add_984151 = sel_984148 + 8'h01;
  assign sel_984152 = array_index_984067 == array_index_948613 ? add_984151 : sel_984148;
  assign add_984155 = sel_984152 + 8'h01;
  assign sel_984156 = array_index_984067 == array_index_948619 ? add_984155 : sel_984152;
  assign add_984159 = sel_984156 + 8'h01;
  assign sel_984160 = array_index_984067 == array_index_948625 ? add_984159 : sel_984156;
  assign add_984163 = sel_984160 + 8'h01;
  assign sel_984164 = array_index_984067 == array_index_948631 ? add_984163 : sel_984160;
  assign add_984167 = sel_984164 + 8'h01;
  assign sel_984168 = array_index_984067 == array_index_948637 ? add_984167 : sel_984164;
  assign add_984171 = sel_984168 + 8'h01;
  assign sel_984172 = array_index_984067 == array_index_948643 ? add_984171 : sel_984168;
  assign add_984175 = sel_984172 + 8'h01;
  assign sel_984176 = array_index_984067 == array_index_948649 ? add_984175 : sel_984172;
  assign add_984179 = sel_984176 + 8'h01;
  assign sel_984180 = array_index_984067 == array_index_948655 ? add_984179 : sel_984176;
  assign add_984183 = sel_984180 + 8'h01;
  assign sel_984184 = array_index_984067 == array_index_948661 ? add_984183 : sel_984180;
  assign add_984187 = sel_984184 + 8'h01;
  assign sel_984188 = array_index_984067 == array_index_948667 ? add_984187 : sel_984184;
  assign add_984191 = sel_984188 + 8'h01;
  assign sel_984192 = array_index_984067 == array_index_948673 ? add_984191 : sel_984188;
  assign add_984195 = sel_984192 + 8'h01;
  assign sel_984196 = array_index_984067 == array_index_948679 ? add_984195 : sel_984192;
  assign add_984199 = sel_984196 + 8'h01;
  assign sel_984200 = array_index_984067 == array_index_948685 ? add_984199 : sel_984196;
  assign add_984203 = sel_984200 + 8'h01;
  assign sel_984204 = array_index_984067 == array_index_948691 ? add_984203 : sel_984200;
  assign add_984207 = sel_984204 + 8'h01;
  assign sel_984208 = array_index_984067 == array_index_948697 ? add_984207 : sel_984204;
  assign add_984211 = sel_984208 + 8'h01;
  assign sel_984212 = array_index_984067 == array_index_948703 ? add_984211 : sel_984208;
  assign add_984215 = sel_984212 + 8'h01;
  assign sel_984216 = array_index_984067 == array_index_948709 ? add_984215 : sel_984212;
  assign add_984219 = sel_984216 + 8'h01;
  assign sel_984220 = array_index_984067 == array_index_948715 ? add_984219 : sel_984216;
  assign add_984223 = sel_984220 + 8'h01;
  assign sel_984224 = array_index_984067 == array_index_948721 ? add_984223 : sel_984220;
  assign add_984227 = sel_984224 + 8'h01;
  assign sel_984228 = array_index_984067 == array_index_948727 ? add_984227 : sel_984224;
  assign add_984231 = sel_984228 + 8'h01;
  assign sel_984232 = array_index_984067 == array_index_948733 ? add_984231 : sel_984228;
  assign add_984235 = sel_984232 + 8'h01;
  assign sel_984236 = array_index_984067 == array_index_948739 ? add_984235 : sel_984232;
  assign add_984239 = sel_984236 + 8'h01;
  assign sel_984240 = array_index_984067 == array_index_948745 ? add_984239 : sel_984236;
  assign add_984243 = sel_984240 + 8'h01;
  assign sel_984244 = array_index_984067 == array_index_948751 ? add_984243 : sel_984240;
  assign add_984247 = sel_984244 + 8'h01;
  assign sel_984248 = array_index_984067 == array_index_948757 ? add_984247 : sel_984244;
  assign add_984251 = sel_984248 + 8'h01;
  assign sel_984252 = array_index_984067 == array_index_948763 ? add_984251 : sel_984248;
  assign add_984255 = sel_984252 + 8'h01;
  assign sel_984256 = array_index_984067 == array_index_948769 ? add_984255 : sel_984252;
  assign add_984259 = sel_984256 + 8'h01;
  assign sel_984260 = array_index_984067 == array_index_948775 ? add_984259 : sel_984256;
  assign add_984263 = sel_984260 + 8'h01;
  assign sel_984264 = array_index_984067 == array_index_948781 ? add_984263 : sel_984260;
  assign add_984267 = sel_984264 + 8'h01;
  assign sel_984268 = array_index_984067 == array_index_948787 ? add_984267 : sel_984264;
  assign add_984271 = sel_984268 + 8'h01;
  assign sel_984272 = array_index_984067 == array_index_948793 ? add_984271 : sel_984268;
  assign add_984275 = sel_984272 + 8'h01;
  assign sel_984276 = array_index_984067 == array_index_948799 ? add_984275 : sel_984272;
  assign add_984279 = sel_984276 + 8'h01;
  assign sel_984280 = array_index_984067 == array_index_948805 ? add_984279 : sel_984276;
  assign add_984283 = sel_984280 + 8'h01;
  assign sel_984284 = array_index_984067 == array_index_948811 ? add_984283 : sel_984280;
  assign add_984287 = sel_984284 + 8'h01;
  assign sel_984288 = array_index_984067 == array_index_948817 ? add_984287 : sel_984284;
  assign add_984291 = sel_984288 + 8'h01;
  assign sel_984292 = array_index_984067 == array_index_948823 ? add_984291 : sel_984288;
  assign add_984295 = sel_984292 + 8'h01;
  assign sel_984296 = array_index_984067 == array_index_948829 ? add_984295 : sel_984292;
  assign add_984299 = sel_984296 + 8'h01;
  assign sel_984300 = array_index_984067 == array_index_948835 ? add_984299 : sel_984296;
  assign add_984303 = sel_984300 + 8'h01;
  assign sel_984304 = array_index_984067 == array_index_948841 ? add_984303 : sel_984300;
  assign add_984307 = sel_984304 + 8'h01;
  assign sel_984308 = array_index_984067 == array_index_948847 ? add_984307 : sel_984304;
  assign add_984311 = sel_984308 + 8'h01;
  assign sel_984312 = array_index_984067 == array_index_948853 ? add_984311 : sel_984308;
  assign add_984315 = sel_984312 + 8'h01;
  assign sel_984316 = array_index_984067 == array_index_948859 ? add_984315 : sel_984312;
  assign add_984319 = sel_984316 + 8'h01;
  assign sel_984320 = array_index_984067 == array_index_948865 ? add_984319 : sel_984316;
  assign add_984323 = sel_984320 + 8'h01;
  assign sel_984324 = array_index_984067 == array_index_948871 ? add_984323 : sel_984320;
  assign add_984327 = sel_984324 + 8'h01;
  assign sel_984328 = array_index_984067 == array_index_948877 ? add_984327 : sel_984324;
  assign add_984331 = sel_984328 + 8'h01;
  assign sel_984332 = array_index_984067 == array_index_948883 ? add_984331 : sel_984328;
  assign add_984335 = sel_984332 + 8'h01;
  assign sel_984336 = array_index_984067 == array_index_948889 ? add_984335 : sel_984332;
  assign add_984339 = sel_984336 + 8'h01;
  assign sel_984340 = array_index_984067 == array_index_948895 ? add_984339 : sel_984336;
  assign add_984343 = sel_984340 + 8'h01;
  assign sel_984344 = array_index_984067 == array_index_948901 ? add_984343 : sel_984340;
  assign add_984347 = sel_984344 + 8'h01;
  assign sel_984348 = array_index_984067 == array_index_948907 ? add_984347 : sel_984344;
  assign add_984351 = sel_984348 + 8'h01;
  assign sel_984352 = array_index_984067 == array_index_948913 ? add_984351 : sel_984348;
  assign add_984355 = sel_984352 + 8'h01;
  assign sel_984356 = array_index_984067 == array_index_948919 ? add_984355 : sel_984352;
  assign add_984359 = sel_984356 + 8'h01;
  assign sel_984360 = array_index_984067 == array_index_948925 ? add_984359 : sel_984356;
  assign add_984363 = sel_984360 + 8'h01;
  assign sel_984364 = array_index_984067 == array_index_948931 ? add_984363 : sel_984360;
  assign add_984367 = sel_984364 + 8'h01;
  assign sel_984368 = array_index_984067 == array_index_948937 ? add_984367 : sel_984364;
  assign add_984371 = sel_984368 + 8'h01;
  assign sel_984372 = array_index_984067 == array_index_948943 ? add_984371 : sel_984368;
  assign add_984375 = sel_984372 + 8'h01;
  assign sel_984376 = array_index_984067 == array_index_948949 ? add_984375 : sel_984372;
  assign add_984379 = sel_984376 + 8'h01;
  assign sel_984380 = array_index_984067 == array_index_948955 ? add_984379 : sel_984376;
  assign add_984383 = sel_984380 + 8'h01;
  assign sel_984384 = array_index_984067 == array_index_948961 ? add_984383 : sel_984380;
  assign add_984387 = sel_984384 + 8'h01;
  assign sel_984388 = array_index_984067 == array_index_948967 ? add_984387 : sel_984384;
  assign add_984391 = sel_984388 + 8'h01;
  assign sel_984392 = array_index_984067 == array_index_948973 ? add_984391 : sel_984388;
  assign add_984395 = sel_984392 + 8'h01;
  assign sel_984396 = array_index_984067 == array_index_948979 ? add_984395 : sel_984392;
  assign add_984399 = sel_984396 + 8'h01;
  assign sel_984400 = array_index_984067 == array_index_948985 ? add_984399 : sel_984396;
  assign add_984403 = sel_984400 + 8'h01;
  assign sel_984404 = array_index_984067 == array_index_948991 ? add_984403 : sel_984400;
  assign add_984407 = sel_984404 + 8'h01;
  assign sel_984408 = array_index_984067 == array_index_948997 ? add_984407 : sel_984404;
  assign add_984411 = sel_984408 + 8'h01;
  assign sel_984412 = array_index_984067 == array_index_949003 ? add_984411 : sel_984408;
  assign add_984415 = sel_984412 + 8'h01;
  assign sel_984416 = array_index_984067 == array_index_949009 ? add_984415 : sel_984412;
  assign add_984419 = sel_984416 + 8'h01;
  assign sel_984420 = array_index_984067 == array_index_949015 ? add_984419 : sel_984416;
  assign add_984423 = sel_984420 + 8'h01;
  assign sel_984424 = array_index_984067 == array_index_949021 ? add_984423 : sel_984420;
  assign add_984427 = sel_984424 + 8'h01;
  assign sel_984428 = array_index_984067 == array_index_949027 ? add_984427 : sel_984424;
  assign add_984431 = sel_984428 + 8'h01;
  assign sel_984432 = array_index_984067 == array_index_949033 ? add_984431 : sel_984428;
  assign add_984435 = sel_984432 + 8'h01;
  assign sel_984436 = array_index_984067 == array_index_949039 ? add_984435 : sel_984432;
  assign add_984439 = sel_984436 + 8'h01;
  assign sel_984440 = array_index_984067 == array_index_949045 ? add_984439 : sel_984436;
  assign add_984443 = sel_984440 + 8'h01;
  assign sel_984444 = array_index_984067 == array_index_949051 ? add_984443 : sel_984440;
  assign add_984447 = sel_984444 + 8'h01;
  assign sel_984448 = array_index_984067 == array_index_949057 ? add_984447 : sel_984444;
  assign add_984451 = sel_984448 + 8'h01;
  assign sel_984452 = array_index_984067 == array_index_949063 ? add_984451 : sel_984448;
  assign add_984455 = sel_984452 + 8'h01;
  assign sel_984456 = array_index_984067 == array_index_949069 ? add_984455 : sel_984452;
  assign add_984459 = sel_984456 + 8'h01;
  assign sel_984460 = array_index_984067 == array_index_949075 ? add_984459 : sel_984456;
  assign add_984463 = sel_984460 + 8'h01;
  assign sel_984464 = array_index_984067 == array_index_949081 ? add_984463 : sel_984460;
  assign add_984468 = sel_984464 + 8'h01;
  assign array_index_984469 = set1_unflattened[7'h59];
  assign sel_984470 = array_index_984067 == array_index_949087 ? add_984468 : sel_984464;
  assign add_984473 = sel_984470 + 8'h01;
  assign sel_984474 = array_index_984469 == array_index_948483 ? add_984473 : sel_984470;
  assign add_984477 = sel_984474 + 8'h01;
  assign sel_984478 = array_index_984469 == array_index_948487 ? add_984477 : sel_984474;
  assign add_984481 = sel_984478 + 8'h01;
  assign sel_984482 = array_index_984469 == array_index_948495 ? add_984481 : sel_984478;
  assign add_984485 = sel_984482 + 8'h01;
  assign sel_984486 = array_index_984469 == array_index_948503 ? add_984485 : sel_984482;
  assign add_984489 = sel_984486 + 8'h01;
  assign sel_984490 = array_index_984469 == array_index_948511 ? add_984489 : sel_984486;
  assign add_984493 = sel_984490 + 8'h01;
  assign sel_984494 = array_index_984469 == array_index_948519 ? add_984493 : sel_984490;
  assign add_984497 = sel_984494 + 8'h01;
  assign sel_984498 = array_index_984469 == array_index_948527 ? add_984497 : sel_984494;
  assign add_984501 = sel_984498 + 8'h01;
  assign sel_984502 = array_index_984469 == array_index_948535 ? add_984501 : sel_984498;
  assign add_984505 = sel_984502 + 8'h01;
  assign sel_984506 = array_index_984469 == array_index_948541 ? add_984505 : sel_984502;
  assign add_984509 = sel_984506 + 8'h01;
  assign sel_984510 = array_index_984469 == array_index_948547 ? add_984509 : sel_984506;
  assign add_984513 = sel_984510 + 8'h01;
  assign sel_984514 = array_index_984469 == array_index_948553 ? add_984513 : sel_984510;
  assign add_984517 = sel_984514 + 8'h01;
  assign sel_984518 = array_index_984469 == array_index_948559 ? add_984517 : sel_984514;
  assign add_984521 = sel_984518 + 8'h01;
  assign sel_984522 = array_index_984469 == array_index_948565 ? add_984521 : sel_984518;
  assign add_984525 = sel_984522 + 8'h01;
  assign sel_984526 = array_index_984469 == array_index_948571 ? add_984525 : sel_984522;
  assign add_984529 = sel_984526 + 8'h01;
  assign sel_984530 = array_index_984469 == array_index_948577 ? add_984529 : sel_984526;
  assign add_984533 = sel_984530 + 8'h01;
  assign sel_984534 = array_index_984469 == array_index_948583 ? add_984533 : sel_984530;
  assign add_984537 = sel_984534 + 8'h01;
  assign sel_984538 = array_index_984469 == array_index_948589 ? add_984537 : sel_984534;
  assign add_984541 = sel_984538 + 8'h01;
  assign sel_984542 = array_index_984469 == array_index_948595 ? add_984541 : sel_984538;
  assign add_984545 = sel_984542 + 8'h01;
  assign sel_984546 = array_index_984469 == array_index_948601 ? add_984545 : sel_984542;
  assign add_984549 = sel_984546 + 8'h01;
  assign sel_984550 = array_index_984469 == array_index_948607 ? add_984549 : sel_984546;
  assign add_984553 = sel_984550 + 8'h01;
  assign sel_984554 = array_index_984469 == array_index_948613 ? add_984553 : sel_984550;
  assign add_984557 = sel_984554 + 8'h01;
  assign sel_984558 = array_index_984469 == array_index_948619 ? add_984557 : sel_984554;
  assign add_984561 = sel_984558 + 8'h01;
  assign sel_984562 = array_index_984469 == array_index_948625 ? add_984561 : sel_984558;
  assign add_984565 = sel_984562 + 8'h01;
  assign sel_984566 = array_index_984469 == array_index_948631 ? add_984565 : sel_984562;
  assign add_984569 = sel_984566 + 8'h01;
  assign sel_984570 = array_index_984469 == array_index_948637 ? add_984569 : sel_984566;
  assign add_984573 = sel_984570 + 8'h01;
  assign sel_984574 = array_index_984469 == array_index_948643 ? add_984573 : sel_984570;
  assign add_984577 = sel_984574 + 8'h01;
  assign sel_984578 = array_index_984469 == array_index_948649 ? add_984577 : sel_984574;
  assign add_984581 = sel_984578 + 8'h01;
  assign sel_984582 = array_index_984469 == array_index_948655 ? add_984581 : sel_984578;
  assign add_984585 = sel_984582 + 8'h01;
  assign sel_984586 = array_index_984469 == array_index_948661 ? add_984585 : sel_984582;
  assign add_984589 = sel_984586 + 8'h01;
  assign sel_984590 = array_index_984469 == array_index_948667 ? add_984589 : sel_984586;
  assign add_984593 = sel_984590 + 8'h01;
  assign sel_984594 = array_index_984469 == array_index_948673 ? add_984593 : sel_984590;
  assign add_984597 = sel_984594 + 8'h01;
  assign sel_984598 = array_index_984469 == array_index_948679 ? add_984597 : sel_984594;
  assign add_984601 = sel_984598 + 8'h01;
  assign sel_984602 = array_index_984469 == array_index_948685 ? add_984601 : sel_984598;
  assign add_984605 = sel_984602 + 8'h01;
  assign sel_984606 = array_index_984469 == array_index_948691 ? add_984605 : sel_984602;
  assign add_984609 = sel_984606 + 8'h01;
  assign sel_984610 = array_index_984469 == array_index_948697 ? add_984609 : sel_984606;
  assign add_984613 = sel_984610 + 8'h01;
  assign sel_984614 = array_index_984469 == array_index_948703 ? add_984613 : sel_984610;
  assign add_984617 = sel_984614 + 8'h01;
  assign sel_984618 = array_index_984469 == array_index_948709 ? add_984617 : sel_984614;
  assign add_984621 = sel_984618 + 8'h01;
  assign sel_984622 = array_index_984469 == array_index_948715 ? add_984621 : sel_984618;
  assign add_984625 = sel_984622 + 8'h01;
  assign sel_984626 = array_index_984469 == array_index_948721 ? add_984625 : sel_984622;
  assign add_984629 = sel_984626 + 8'h01;
  assign sel_984630 = array_index_984469 == array_index_948727 ? add_984629 : sel_984626;
  assign add_984633 = sel_984630 + 8'h01;
  assign sel_984634 = array_index_984469 == array_index_948733 ? add_984633 : sel_984630;
  assign add_984637 = sel_984634 + 8'h01;
  assign sel_984638 = array_index_984469 == array_index_948739 ? add_984637 : sel_984634;
  assign add_984641 = sel_984638 + 8'h01;
  assign sel_984642 = array_index_984469 == array_index_948745 ? add_984641 : sel_984638;
  assign add_984645 = sel_984642 + 8'h01;
  assign sel_984646 = array_index_984469 == array_index_948751 ? add_984645 : sel_984642;
  assign add_984649 = sel_984646 + 8'h01;
  assign sel_984650 = array_index_984469 == array_index_948757 ? add_984649 : sel_984646;
  assign add_984653 = sel_984650 + 8'h01;
  assign sel_984654 = array_index_984469 == array_index_948763 ? add_984653 : sel_984650;
  assign add_984657 = sel_984654 + 8'h01;
  assign sel_984658 = array_index_984469 == array_index_948769 ? add_984657 : sel_984654;
  assign add_984661 = sel_984658 + 8'h01;
  assign sel_984662 = array_index_984469 == array_index_948775 ? add_984661 : sel_984658;
  assign add_984665 = sel_984662 + 8'h01;
  assign sel_984666 = array_index_984469 == array_index_948781 ? add_984665 : sel_984662;
  assign add_984669 = sel_984666 + 8'h01;
  assign sel_984670 = array_index_984469 == array_index_948787 ? add_984669 : sel_984666;
  assign add_984673 = sel_984670 + 8'h01;
  assign sel_984674 = array_index_984469 == array_index_948793 ? add_984673 : sel_984670;
  assign add_984677 = sel_984674 + 8'h01;
  assign sel_984678 = array_index_984469 == array_index_948799 ? add_984677 : sel_984674;
  assign add_984681 = sel_984678 + 8'h01;
  assign sel_984682 = array_index_984469 == array_index_948805 ? add_984681 : sel_984678;
  assign add_984685 = sel_984682 + 8'h01;
  assign sel_984686 = array_index_984469 == array_index_948811 ? add_984685 : sel_984682;
  assign add_984689 = sel_984686 + 8'h01;
  assign sel_984690 = array_index_984469 == array_index_948817 ? add_984689 : sel_984686;
  assign add_984693 = sel_984690 + 8'h01;
  assign sel_984694 = array_index_984469 == array_index_948823 ? add_984693 : sel_984690;
  assign add_984697 = sel_984694 + 8'h01;
  assign sel_984698 = array_index_984469 == array_index_948829 ? add_984697 : sel_984694;
  assign add_984701 = sel_984698 + 8'h01;
  assign sel_984702 = array_index_984469 == array_index_948835 ? add_984701 : sel_984698;
  assign add_984705 = sel_984702 + 8'h01;
  assign sel_984706 = array_index_984469 == array_index_948841 ? add_984705 : sel_984702;
  assign add_984709 = sel_984706 + 8'h01;
  assign sel_984710 = array_index_984469 == array_index_948847 ? add_984709 : sel_984706;
  assign add_984713 = sel_984710 + 8'h01;
  assign sel_984714 = array_index_984469 == array_index_948853 ? add_984713 : sel_984710;
  assign add_984717 = sel_984714 + 8'h01;
  assign sel_984718 = array_index_984469 == array_index_948859 ? add_984717 : sel_984714;
  assign add_984721 = sel_984718 + 8'h01;
  assign sel_984722 = array_index_984469 == array_index_948865 ? add_984721 : sel_984718;
  assign add_984725 = sel_984722 + 8'h01;
  assign sel_984726 = array_index_984469 == array_index_948871 ? add_984725 : sel_984722;
  assign add_984729 = sel_984726 + 8'h01;
  assign sel_984730 = array_index_984469 == array_index_948877 ? add_984729 : sel_984726;
  assign add_984733 = sel_984730 + 8'h01;
  assign sel_984734 = array_index_984469 == array_index_948883 ? add_984733 : sel_984730;
  assign add_984737 = sel_984734 + 8'h01;
  assign sel_984738 = array_index_984469 == array_index_948889 ? add_984737 : sel_984734;
  assign add_984741 = sel_984738 + 8'h01;
  assign sel_984742 = array_index_984469 == array_index_948895 ? add_984741 : sel_984738;
  assign add_984745 = sel_984742 + 8'h01;
  assign sel_984746 = array_index_984469 == array_index_948901 ? add_984745 : sel_984742;
  assign add_984749 = sel_984746 + 8'h01;
  assign sel_984750 = array_index_984469 == array_index_948907 ? add_984749 : sel_984746;
  assign add_984753 = sel_984750 + 8'h01;
  assign sel_984754 = array_index_984469 == array_index_948913 ? add_984753 : sel_984750;
  assign add_984757 = sel_984754 + 8'h01;
  assign sel_984758 = array_index_984469 == array_index_948919 ? add_984757 : sel_984754;
  assign add_984761 = sel_984758 + 8'h01;
  assign sel_984762 = array_index_984469 == array_index_948925 ? add_984761 : sel_984758;
  assign add_984765 = sel_984762 + 8'h01;
  assign sel_984766 = array_index_984469 == array_index_948931 ? add_984765 : sel_984762;
  assign add_984769 = sel_984766 + 8'h01;
  assign sel_984770 = array_index_984469 == array_index_948937 ? add_984769 : sel_984766;
  assign add_984773 = sel_984770 + 8'h01;
  assign sel_984774 = array_index_984469 == array_index_948943 ? add_984773 : sel_984770;
  assign add_984777 = sel_984774 + 8'h01;
  assign sel_984778 = array_index_984469 == array_index_948949 ? add_984777 : sel_984774;
  assign add_984781 = sel_984778 + 8'h01;
  assign sel_984782 = array_index_984469 == array_index_948955 ? add_984781 : sel_984778;
  assign add_984785 = sel_984782 + 8'h01;
  assign sel_984786 = array_index_984469 == array_index_948961 ? add_984785 : sel_984782;
  assign add_984789 = sel_984786 + 8'h01;
  assign sel_984790 = array_index_984469 == array_index_948967 ? add_984789 : sel_984786;
  assign add_984793 = sel_984790 + 8'h01;
  assign sel_984794 = array_index_984469 == array_index_948973 ? add_984793 : sel_984790;
  assign add_984797 = sel_984794 + 8'h01;
  assign sel_984798 = array_index_984469 == array_index_948979 ? add_984797 : sel_984794;
  assign add_984801 = sel_984798 + 8'h01;
  assign sel_984802 = array_index_984469 == array_index_948985 ? add_984801 : sel_984798;
  assign add_984805 = sel_984802 + 8'h01;
  assign sel_984806 = array_index_984469 == array_index_948991 ? add_984805 : sel_984802;
  assign add_984809 = sel_984806 + 8'h01;
  assign sel_984810 = array_index_984469 == array_index_948997 ? add_984809 : sel_984806;
  assign add_984813 = sel_984810 + 8'h01;
  assign sel_984814 = array_index_984469 == array_index_949003 ? add_984813 : sel_984810;
  assign add_984817 = sel_984814 + 8'h01;
  assign sel_984818 = array_index_984469 == array_index_949009 ? add_984817 : sel_984814;
  assign add_984821 = sel_984818 + 8'h01;
  assign sel_984822 = array_index_984469 == array_index_949015 ? add_984821 : sel_984818;
  assign add_984825 = sel_984822 + 8'h01;
  assign sel_984826 = array_index_984469 == array_index_949021 ? add_984825 : sel_984822;
  assign add_984829 = sel_984826 + 8'h01;
  assign sel_984830 = array_index_984469 == array_index_949027 ? add_984829 : sel_984826;
  assign add_984833 = sel_984830 + 8'h01;
  assign sel_984834 = array_index_984469 == array_index_949033 ? add_984833 : sel_984830;
  assign add_984837 = sel_984834 + 8'h01;
  assign sel_984838 = array_index_984469 == array_index_949039 ? add_984837 : sel_984834;
  assign add_984841 = sel_984838 + 8'h01;
  assign sel_984842 = array_index_984469 == array_index_949045 ? add_984841 : sel_984838;
  assign add_984845 = sel_984842 + 8'h01;
  assign sel_984846 = array_index_984469 == array_index_949051 ? add_984845 : sel_984842;
  assign add_984849 = sel_984846 + 8'h01;
  assign sel_984850 = array_index_984469 == array_index_949057 ? add_984849 : sel_984846;
  assign add_984853 = sel_984850 + 8'h01;
  assign sel_984854 = array_index_984469 == array_index_949063 ? add_984853 : sel_984850;
  assign add_984857 = sel_984854 + 8'h01;
  assign sel_984858 = array_index_984469 == array_index_949069 ? add_984857 : sel_984854;
  assign add_984861 = sel_984858 + 8'h01;
  assign sel_984862 = array_index_984469 == array_index_949075 ? add_984861 : sel_984858;
  assign add_984865 = sel_984862 + 8'h01;
  assign sel_984866 = array_index_984469 == array_index_949081 ? add_984865 : sel_984862;
  assign add_984870 = sel_984866 + 8'h01;
  assign array_index_984871 = set1_unflattened[7'h5a];
  assign sel_984872 = array_index_984469 == array_index_949087 ? add_984870 : sel_984866;
  assign add_984875 = sel_984872 + 8'h01;
  assign sel_984876 = array_index_984871 == array_index_948483 ? add_984875 : sel_984872;
  assign add_984879 = sel_984876 + 8'h01;
  assign sel_984880 = array_index_984871 == array_index_948487 ? add_984879 : sel_984876;
  assign add_984883 = sel_984880 + 8'h01;
  assign sel_984884 = array_index_984871 == array_index_948495 ? add_984883 : sel_984880;
  assign add_984887 = sel_984884 + 8'h01;
  assign sel_984888 = array_index_984871 == array_index_948503 ? add_984887 : sel_984884;
  assign add_984891 = sel_984888 + 8'h01;
  assign sel_984892 = array_index_984871 == array_index_948511 ? add_984891 : sel_984888;
  assign add_984895 = sel_984892 + 8'h01;
  assign sel_984896 = array_index_984871 == array_index_948519 ? add_984895 : sel_984892;
  assign add_984899 = sel_984896 + 8'h01;
  assign sel_984900 = array_index_984871 == array_index_948527 ? add_984899 : sel_984896;
  assign add_984903 = sel_984900 + 8'h01;
  assign sel_984904 = array_index_984871 == array_index_948535 ? add_984903 : sel_984900;
  assign add_984907 = sel_984904 + 8'h01;
  assign sel_984908 = array_index_984871 == array_index_948541 ? add_984907 : sel_984904;
  assign add_984911 = sel_984908 + 8'h01;
  assign sel_984912 = array_index_984871 == array_index_948547 ? add_984911 : sel_984908;
  assign add_984915 = sel_984912 + 8'h01;
  assign sel_984916 = array_index_984871 == array_index_948553 ? add_984915 : sel_984912;
  assign add_984919 = sel_984916 + 8'h01;
  assign sel_984920 = array_index_984871 == array_index_948559 ? add_984919 : sel_984916;
  assign add_984923 = sel_984920 + 8'h01;
  assign sel_984924 = array_index_984871 == array_index_948565 ? add_984923 : sel_984920;
  assign add_984927 = sel_984924 + 8'h01;
  assign sel_984928 = array_index_984871 == array_index_948571 ? add_984927 : sel_984924;
  assign add_984931 = sel_984928 + 8'h01;
  assign sel_984932 = array_index_984871 == array_index_948577 ? add_984931 : sel_984928;
  assign add_984935 = sel_984932 + 8'h01;
  assign sel_984936 = array_index_984871 == array_index_948583 ? add_984935 : sel_984932;
  assign add_984939 = sel_984936 + 8'h01;
  assign sel_984940 = array_index_984871 == array_index_948589 ? add_984939 : sel_984936;
  assign add_984943 = sel_984940 + 8'h01;
  assign sel_984944 = array_index_984871 == array_index_948595 ? add_984943 : sel_984940;
  assign add_984947 = sel_984944 + 8'h01;
  assign sel_984948 = array_index_984871 == array_index_948601 ? add_984947 : sel_984944;
  assign add_984951 = sel_984948 + 8'h01;
  assign sel_984952 = array_index_984871 == array_index_948607 ? add_984951 : sel_984948;
  assign add_984955 = sel_984952 + 8'h01;
  assign sel_984956 = array_index_984871 == array_index_948613 ? add_984955 : sel_984952;
  assign add_984959 = sel_984956 + 8'h01;
  assign sel_984960 = array_index_984871 == array_index_948619 ? add_984959 : sel_984956;
  assign add_984963 = sel_984960 + 8'h01;
  assign sel_984964 = array_index_984871 == array_index_948625 ? add_984963 : sel_984960;
  assign add_984967 = sel_984964 + 8'h01;
  assign sel_984968 = array_index_984871 == array_index_948631 ? add_984967 : sel_984964;
  assign add_984971 = sel_984968 + 8'h01;
  assign sel_984972 = array_index_984871 == array_index_948637 ? add_984971 : sel_984968;
  assign add_984975 = sel_984972 + 8'h01;
  assign sel_984976 = array_index_984871 == array_index_948643 ? add_984975 : sel_984972;
  assign add_984979 = sel_984976 + 8'h01;
  assign sel_984980 = array_index_984871 == array_index_948649 ? add_984979 : sel_984976;
  assign add_984983 = sel_984980 + 8'h01;
  assign sel_984984 = array_index_984871 == array_index_948655 ? add_984983 : sel_984980;
  assign add_984987 = sel_984984 + 8'h01;
  assign sel_984988 = array_index_984871 == array_index_948661 ? add_984987 : sel_984984;
  assign add_984991 = sel_984988 + 8'h01;
  assign sel_984992 = array_index_984871 == array_index_948667 ? add_984991 : sel_984988;
  assign add_984995 = sel_984992 + 8'h01;
  assign sel_984996 = array_index_984871 == array_index_948673 ? add_984995 : sel_984992;
  assign add_984999 = sel_984996 + 8'h01;
  assign sel_985000 = array_index_984871 == array_index_948679 ? add_984999 : sel_984996;
  assign add_985003 = sel_985000 + 8'h01;
  assign sel_985004 = array_index_984871 == array_index_948685 ? add_985003 : sel_985000;
  assign add_985007 = sel_985004 + 8'h01;
  assign sel_985008 = array_index_984871 == array_index_948691 ? add_985007 : sel_985004;
  assign add_985011 = sel_985008 + 8'h01;
  assign sel_985012 = array_index_984871 == array_index_948697 ? add_985011 : sel_985008;
  assign add_985015 = sel_985012 + 8'h01;
  assign sel_985016 = array_index_984871 == array_index_948703 ? add_985015 : sel_985012;
  assign add_985019 = sel_985016 + 8'h01;
  assign sel_985020 = array_index_984871 == array_index_948709 ? add_985019 : sel_985016;
  assign add_985023 = sel_985020 + 8'h01;
  assign sel_985024 = array_index_984871 == array_index_948715 ? add_985023 : sel_985020;
  assign add_985027 = sel_985024 + 8'h01;
  assign sel_985028 = array_index_984871 == array_index_948721 ? add_985027 : sel_985024;
  assign add_985031 = sel_985028 + 8'h01;
  assign sel_985032 = array_index_984871 == array_index_948727 ? add_985031 : sel_985028;
  assign add_985035 = sel_985032 + 8'h01;
  assign sel_985036 = array_index_984871 == array_index_948733 ? add_985035 : sel_985032;
  assign add_985039 = sel_985036 + 8'h01;
  assign sel_985040 = array_index_984871 == array_index_948739 ? add_985039 : sel_985036;
  assign add_985043 = sel_985040 + 8'h01;
  assign sel_985044 = array_index_984871 == array_index_948745 ? add_985043 : sel_985040;
  assign add_985047 = sel_985044 + 8'h01;
  assign sel_985048 = array_index_984871 == array_index_948751 ? add_985047 : sel_985044;
  assign add_985051 = sel_985048 + 8'h01;
  assign sel_985052 = array_index_984871 == array_index_948757 ? add_985051 : sel_985048;
  assign add_985055 = sel_985052 + 8'h01;
  assign sel_985056 = array_index_984871 == array_index_948763 ? add_985055 : sel_985052;
  assign add_985059 = sel_985056 + 8'h01;
  assign sel_985060 = array_index_984871 == array_index_948769 ? add_985059 : sel_985056;
  assign add_985063 = sel_985060 + 8'h01;
  assign sel_985064 = array_index_984871 == array_index_948775 ? add_985063 : sel_985060;
  assign add_985067 = sel_985064 + 8'h01;
  assign sel_985068 = array_index_984871 == array_index_948781 ? add_985067 : sel_985064;
  assign add_985071 = sel_985068 + 8'h01;
  assign sel_985072 = array_index_984871 == array_index_948787 ? add_985071 : sel_985068;
  assign add_985075 = sel_985072 + 8'h01;
  assign sel_985076 = array_index_984871 == array_index_948793 ? add_985075 : sel_985072;
  assign add_985079 = sel_985076 + 8'h01;
  assign sel_985080 = array_index_984871 == array_index_948799 ? add_985079 : sel_985076;
  assign add_985083 = sel_985080 + 8'h01;
  assign sel_985084 = array_index_984871 == array_index_948805 ? add_985083 : sel_985080;
  assign add_985087 = sel_985084 + 8'h01;
  assign sel_985088 = array_index_984871 == array_index_948811 ? add_985087 : sel_985084;
  assign add_985091 = sel_985088 + 8'h01;
  assign sel_985092 = array_index_984871 == array_index_948817 ? add_985091 : sel_985088;
  assign add_985095 = sel_985092 + 8'h01;
  assign sel_985096 = array_index_984871 == array_index_948823 ? add_985095 : sel_985092;
  assign add_985099 = sel_985096 + 8'h01;
  assign sel_985100 = array_index_984871 == array_index_948829 ? add_985099 : sel_985096;
  assign add_985103 = sel_985100 + 8'h01;
  assign sel_985104 = array_index_984871 == array_index_948835 ? add_985103 : sel_985100;
  assign add_985107 = sel_985104 + 8'h01;
  assign sel_985108 = array_index_984871 == array_index_948841 ? add_985107 : sel_985104;
  assign add_985111 = sel_985108 + 8'h01;
  assign sel_985112 = array_index_984871 == array_index_948847 ? add_985111 : sel_985108;
  assign add_985115 = sel_985112 + 8'h01;
  assign sel_985116 = array_index_984871 == array_index_948853 ? add_985115 : sel_985112;
  assign add_985119 = sel_985116 + 8'h01;
  assign sel_985120 = array_index_984871 == array_index_948859 ? add_985119 : sel_985116;
  assign add_985123 = sel_985120 + 8'h01;
  assign sel_985124 = array_index_984871 == array_index_948865 ? add_985123 : sel_985120;
  assign add_985127 = sel_985124 + 8'h01;
  assign sel_985128 = array_index_984871 == array_index_948871 ? add_985127 : sel_985124;
  assign add_985131 = sel_985128 + 8'h01;
  assign sel_985132 = array_index_984871 == array_index_948877 ? add_985131 : sel_985128;
  assign add_985135 = sel_985132 + 8'h01;
  assign sel_985136 = array_index_984871 == array_index_948883 ? add_985135 : sel_985132;
  assign add_985139 = sel_985136 + 8'h01;
  assign sel_985140 = array_index_984871 == array_index_948889 ? add_985139 : sel_985136;
  assign add_985143 = sel_985140 + 8'h01;
  assign sel_985144 = array_index_984871 == array_index_948895 ? add_985143 : sel_985140;
  assign add_985147 = sel_985144 + 8'h01;
  assign sel_985148 = array_index_984871 == array_index_948901 ? add_985147 : sel_985144;
  assign add_985151 = sel_985148 + 8'h01;
  assign sel_985152 = array_index_984871 == array_index_948907 ? add_985151 : sel_985148;
  assign add_985155 = sel_985152 + 8'h01;
  assign sel_985156 = array_index_984871 == array_index_948913 ? add_985155 : sel_985152;
  assign add_985159 = sel_985156 + 8'h01;
  assign sel_985160 = array_index_984871 == array_index_948919 ? add_985159 : sel_985156;
  assign add_985163 = sel_985160 + 8'h01;
  assign sel_985164 = array_index_984871 == array_index_948925 ? add_985163 : sel_985160;
  assign add_985167 = sel_985164 + 8'h01;
  assign sel_985168 = array_index_984871 == array_index_948931 ? add_985167 : sel_985164;
  assign add_985171 = sel_985168 + 8'h01;
  assign sel_985172 = array_index_984871 == array_index_948937 ? add_985171 : sel_985168;
  assign add_985175 = sel_985172 + 8'h01;
  assign sel_985176 = array_index_984871 == array_index_948943 ? add_985175 : sel_985172;
  assign add_985179 = sel_985176 + 8'h01;
  assign sel_985180 = array_index_984871 == array_index_948949 ? add_985179 : sel_985176;
  assign add_985183 = sel_985180 + 8'h01;
  assign sel_985184 = array_index_984871 == array_index_948955 ? add_985183 : sel_985180;
  assign add_985187 = sel_985184 + 8'h01;
  assign sel_985188 = array_index_984871 == array_index_948961 ? add_985187 : sel_985184;
  assign add_985191 = sel_985188 + 8'h01;
  assign sel_985192 = array_index_984871 == array_index_948967 ? add_985191 : sel_985188;
  assign add_985195 = sel_985192 + 8'h01;
  assign sel_985196 = array_index_984871 == array_index_948973 ? add_985195 : sel_985192;
  assign add_985199 = sel_985196 + 8'h01;
  assign sel_985200 = array_index_984871 == array_index_948979 ? add_985199 : sel_985196;
  assign add_985203 = sel_985200 + 8'h01;
  assign sel_985204 = array_index_984871 == array_index_948985 ? add_985203 : sel_985200;
  assign add_985207 = sel_985204 + 8'h01;
  assign sel_985208 = array_index_984871 == array_index_948991 ? add_985207 : sel_985204;
  assign add_985211 = sel_985208 + 8'h01;
  assign sel_985212 = array_index_984871 == array_index_948997 ? add_985211 : sel_985208;
  assign add_985215 = sel_985212 + 8'h01;
  assign sel_985216 = array_index_984871 == array_index_949003 ? add_985215 : sel_985212;
  assign add_985219 = sel_985216 + 8'h01;
  assign sel_985220 = array_index_984871 == array_index_949009 ? add_985219 : sel_985216;
  assign add_985223 = sel_985220 + 8'h01;
  assign sel_985224 = array_index_984871 == array_index_949015 ? add_985223 : sel_985220;
  assign add_985227 = sel_985224 + 8'h01;
  assign sel_985228 = array_index_984871 == array_index_949021 ? add_985227 : sel_985224;
  assign add_985231 = sel_985228 + 8'h01;
  assign sel_985232 = array_index_984871 == array_index_949027 ? add_985231 : sel_985228;
  assign add_985235 = sel_985232 + 8'h01;
  assign sel_985236 = array_index_984871 == array_index_949033 ? add_985235 : sel_985232;
  assign add_985239 = sel_985236 + 8'h01;
  assign sel_985240 = array_index_984871 == array_index_949039 ? add_985239 : sel_985236;
  assign add_985243 = sel_985240 + 8'h01;
  assign sel_985244 = array_index_984871 == array_index_949045 ? add_985243 : sel_985240;
  assign add_985247 = sel_985244 + 8'h01;
  assign sel_985248 = array_index_984871 == array_index_949051 ? add_985247 : sel_985244;
  assign add_985251 = sel_985248 + 8'h01;
  assign sel_985252 = array_index_984871 == array_index_949057 ? add_985251 : sel_985248;
  assign add_985255 = sel_985252 + 8'h01;
  assign sel_985256 = array_index_984871 == array_index_949063 ? add_985255 : sel_985252;
  assign add_985259 = sel_985256 + 8'h01;
  assign sel_985260 = array_index_984871 == array_index_949069 ? add_985259 : sel_985256;
  assign add_985263 = sel_985260 + 8'h01;
  assign sel_985264 = array_index_984871 == array_index_949075 ? add_985263 : sel_985260;
  assign add_985267 = sel_985264 + 8'h01;
  assign sel_985268 = array_index_984871 == array_index_949081 ? add_985267 : sel_985264;
  assign add_985272 = sel_985268 + 8'h01;
  assign array_index_985273 = set1_unflattened[7'h5b];
  assign sel_985274 = array_index_984871 == array_index_949087 ? add_985272 : sel_985268;
  assign add_985277 = sel_985274 + 8'h01;
  assign sel_985278 = array_index_985273 == array_index_948483 ? add_985277 : sel_985274;
  assign add_985281 = sel_985278 + 8'h01;
  assign sel_985282 = array_index_985273 == array_index_948487 ? add_985281 : sel_985278;
  assign add_985285 = sel_985282 + 8'h01;
  assign sel_985286 = array_index_985273 == array_index_948495 ? add_985285 : sel_985282;
  assign add_985289 = sel_985286 + 8'h01;
  assign sel_985290 = array_index_985273 == array_index_948503 ? add_985289 : sel_985286;
  assign add_985293 = sel_985290 + 8'h01;
  assign sel_985294 = array_index_985273 == array_index_948511 ? add_985293 : sel_985290;
  assign add_985297 = sel_985294 + 8'h01;
  assign sel_985298 = array_index_985273 == array_index_948519 ? add_985297 : sel_985294;
  assign add_985301 = sel_985298 + 8'h01;
  assign sel_985302 = array_index_985273 == array_index_948527 ? add_985301 : sel_985298;
  assign add_985305 = sel_985302 + 8'h01;
  assign sel_985306 = array_index_985273 == array_index_948535 ? add_985305 : sel_985302;
  assign add_985309 = sel_985306 + 8'h01;
  assign sel_985310 = array_index_985273 == array_index_948541 ? add_985309 : sel_985306;
  assign add_985313 = sel_985310 + 8'h01;
  assign sel_985314 = array_index_985273 == array_index_948547 ? add_985313 : sel_985310;
  assign add_985317 = sel_985314 + 8'h01;
  assign sel_985318 = array_index_985273 == array_index_948553 ? add_985317 : sel_985314;
  assign add_985321 = sel_985318 + 8'h01;
  assign sel_985322 = array_index_985273 == array_index_948559 ? add_985321 : sel_985318;
  assign add_985325 = sel_985322 + 8'h01;
  assign sel_985326 = array_index_985273 == array_index_948565 ? add_985325 : sel_985322;
  assign add_985329 = sel_985326 + 8'h01;
  assign sel_985330 = array_index_985273 == array_index_948571 ? add_985329 : sel_985326;
  assign add_985333 = sel_985330 + 8'h01;
  assign sel_985334 = array_index_985273 == array_index_948577 ? add_985333 : sel_985330;
  assign add_985337 = sel_985334 + 8'h01;
  assign sel_985338 = array_index_985273 == array_index_948583 ? add_985337 : sel_985334;
  assign add_985341 = sel_985338 + 8'h01;
  assign sel_985342 = array_index_985273 == array_index_948589 ? add_985341 : sel_985338;
  assign add_985345 = sel_985342 + 8'h01;
  assign sel_985346 = array_index_985273 == array_index_948595 ? add_985345 : sel_985342;
  assign add_985349 = sel_985346 + 8'h01;
  assign sel_985350 = array_index_985273 == array_index_948601 ? add_985349 : sel_985346;
  assign add_985353 = sel_985350 + 8'h01;
  assign sel_985354 = array_index_985273 == array_index_948607 ? add_985353 : sel_985350;
  assign add_985357 = sel_985354 + 8'h01;
  assign sel_985358 = array_index_985273 == array_index_948613 ? add_985357 : sel_985354;
  assign add_985361 = sel_985358 + 8'h01;
  assign sel_985362 = array_index_985273 == array_index_948619 ? add_985361 : sel_985358;
  assign add_985365 = sel_985362 + 8'h01;
  assign sel_985366 = array_index_985273 == array_index_948625 ? add_985365 : sel_985362;
  assign add_985369 = sel_985366 + 8'h01;
  assign sel_985370 = array_index_985273 == array_index_948631 ? add_985369 : sel_985366;
  assign add_985373 = sel_985370 + 8'h01;
  assign sel_985374 = array_index_985273 == array_index_948637 ? add_985373 : sel_985370;
  assign add_985377 = sel_985374 + 8'h01;
  assign sel_985378 = array_index_985273 == array_index_948643 ? add_985377 : sel_985374;
  assign add_985381 = sel_985378 + 8'h01;
  assign sel_985382 = array_index_985273 == array_index_948649 ? add_985381 : sel_985378;
  assign add_985385 = sel_985382 + 8'h01;
  assign sel_985386 = array_index_985273 == array_index_948655 ? add_985385 : sel_985382;
  assign add_985389 = sel_985386 + 8'h01;
  assign sel_985390 = array_index_985273 == array_index_948661 ? add_985389 : sel_985386;
  assign add_985393 = sel_985390 + 8'h01;
  assign sel_985394 = array_index_985273 == array_index_948667 ? add_985393 : sel_985390;
  assign add_985397 = sel_985394 + 8'h01;
  assign sel_985398 = array_index_985273 == array_index_948673 ? add_985397 : sel_985394;
  assign add_985401 = sel_985398 + 8'h01;
  assign sel_985402 = array_index_985273 == array_index_948679 ? add_985401 : sel_985398;
  assign add_985405 = sel_985402 + 8'h01;
  assign sel_985406 = array_index_985273 == array_index_948685 ? add_985405 : sel_985402;
  assign add_985409 = sel_985406 + 8'h01;
  assign sel_985410 = array_index_985273 == array_index_948691 ? add_985409 : sel_985406;
  assign add_985413 = sel_985410 + 8'h01;
  assign sel_985414 = array_index_985273 == array_index_948697 ? add_985413 : sel_985410;
  assign add_985417 = sel_985414 + 8'h01;
  assign sel_985418 = array_index_985273 == array_index_948703 ? add_985417 : sel_985414;
  assign add_985421 = sel_985418 + 8'h01;
  assign sel_985422 = array_index_985273 == array_index_948709 ? add_985421 : sel_985418;
  assign add_985425 = sel_985422 + 8'h01;
  assign sel_985426 = array_index_985273 == array_index_948715 ? add_985425 : sel_985422;
  assign add_985429 = sel_985426 + 8'h01;
  assign sel_985430 = array_index_985273 == array_index_948721 ? add_985429 : sel_985426;
  assign add_985433 = sel_985430 + 8'h01;
  assign sel_985434 = array_index_985273 == array_index_948727 ? add_985433 : sel_985430;
  assign add_985437 = sel_985434 + 8'h01;
  assign sel_985438 = array_index_985273 == array_index_948733 ? add_985437 : sel_985434;
  assign add_985441 = sel_985438 + 8'h01;
  assign sel_985442 = array_index_985273 == array_index_948739 ? add_985441 : sel_985438;
  assign add_985445 = sel_985442 + 8'h01;
  assign sel_985446 = array_index_985273 == array_index_948745 ? add_985445 : sel_985442;
  assign add_985449 = sel_985446 + 8'h01;
  assign sel_985450 = array_index_985273 == array_index_948751 ? add_985449 : sel_985446;
  assign add_985453 = sel_985450 + 8'h01;
  assign sel_985454 = array_index_985273 == array_index_948757 ? add_985453 : sel_985450;
  assign add_985457 = sel_985454 + 8'h01;
  assign sel_985458 = array_index_985273 == array_index_948763 ? add_985457 : sel_985454;
  assign add_985461 = sel_985458 + 8'h01;
  assign sel_985462 = array_index_985273 == array_index_948769 ? add_985461 : sel_985458;
  assign add_985465 = sel_985462 + 8'h01;
  assign sel_985466 = array_index_985273 == array_index_948775 ? add_985465 : sel_985462;
  assign add_985469 = sel_985466 + 8'h01;
  assign sel_985470 = array_index_985273 == array_index_948781 ? add_985469 : sel_985466;
  assign add_985473 = sel_985470 + 8'h01;
  assign sel_985474 = array_index_985273 == array_index_948787 ? add_985473 : sel_985470;
  assign add_985477 = sel_985474 + 8'h01;
  assign sel_985478 = array_index_985273 == array_index_948793 ? add_985477 : sel_985474;
  assign add_985481 = sel_985478 + 8'h01;
  assign sel_985482 = array_index_985273 == array_index_948799 ? add_985481 : sel_985478;
  assign add_985485 = sel_985482 + 8'h01;
  assign sel_985486 = array_index_985273 == array_index_948805 ? add_985485 : sel_985482;
  assign add_985489 = sel_985486 + 8'h01;
  assign sel_985490 = array_index_985273 == array_index_948811 ? add_985489 : sel_985486;
  assign add_985493 = sel_985490 + 8'h01;
  assign sel_985494 = array_index_985273 == array_index_948817 ? add_985493 : sel_985490;
  assign add_985497 = sel_985494 + 8'h01;
  assign sel_985498 = array_index_985273 == array_index_948823 ? add_985497 : sel_985494;
  assign add_985501 = sel_985498 + 8'h01;
  assign sel_985502 = array_index_985273 == array_index_948829 ? add_985501 : sel_985498;
  assign add_985505 = sel_985502 + 8'h01;
  assign sel_985506 = array_index_985273 == array_index_948835 ? add_985505 : sel_985502;
  assign add_985509 = sel_985506 + 8'h01;
  assign sel_985510 = array_index_985273 == array_index_948841 ? add_985509 : sel_985506;
  assign add_985513 = sel_985510 + 8'h01;
  assign sel_985514 = array_index_985273 == array_index_948847 ? add_985513 : sel_985510;
  assign add_985517 = sel_985514 + 8'h01;
  assign sel_985518 = array_index_985273 == array_index_948853 ? add_985517 : sel_985514;
  assign add_985521 = sel_985518 + 8'h01;
  assign sel_985522 = array_index_985273 == array_index_948859 ? add_985521 : sel_985518;
  assign add_985525 = sel_985522 + 8'h01;
  assign sel_985526 = array_index_985273 == array_index_948865 ? add_985525 : sel_985522;
  assign add_985529 = sel_985526 + 8'h01;
  assign sel_985530 = array_index_985273 == array_index_948871 ? add_985529 : sel_985526;
  assign add_985533 = sel_985530 + 8'h01;
  assign sel_985534 = array_index_985273 == array_index_948877 ? add_985533 : sel_985530;
  assign add_985537 = sel_985534 + 8'h01;
  assign sel_985538 = array_index_985273 == array_index_948883 ? add_985537 : sel_985534;
  assign add_985541 = sel_985538 + 8'h01;
  assign sel_985542 = array_index_985273 == array_index_948889 ? add_985541 : sel_985538;
  assign add_985545 = sel_985542 + 8'h01;
  assign sel_985546 = array_index_985273 == array_index_948895 ? add_985545 : sel_985542;
  assign add_985549 = sel_985546 + 8'h01;
  assign sel_985550 = array_index_985273 == array_index_948901 ? add_985549 : sel_985546;
  assign add_985553 = sel_985550 + 8'h01;
  assign sel_985554 = array_index_985273 == array_index_948907 ? add_985553 : sel_985550;
  assign add_985557 = sel_985554 + 8'h01;
  assign sel_985558 = array_index_985273 == array_index_948913 ? add_985557 : sel_985554;
  assign add_985561 = sel_985558 + 8'h01;
  assign sel_985562 = array_index_985273 == array_index_948919 ? add_985561 : sel_985558;
  assign add_985565 = sel_985562 + 8'h01;
  assign sel_985566 = array_index_985273 == array_index_948925 ? add_985565 : sel_985562;
  assign add_985569 = sel_985566 + 8'h01;
  assign sel_985570 = array_index_985273 == array_index_948931 ? add_985569 : sel_985566;
  assign add_985573 = sel_985570 + 8'h01;
  assign sel_985574 = array_index_985273 == array_index_948937 ? add_985573 : sel_985570;
  assign add_985577 = sel_985574 + 8'h01;
  assign sel_985578 = array_index_985273 == array_index_948943 ? add_985577 : sel_985574;
  assign add_985581 = sel_985578 + 8'h01;
  assign sel_985582 = array_index_985273 == array_index_948949 ? add_985581 : sel_985578;
  assign add_985585 = sel_985582 + 8'h01;
  assign sel_985586 = array_index_985273 == array_index_948955 ? add_985585 : sel_985582;
  assign add_985589 = sel_985586 + 8'h01;
  assign sel_985590 = array_index_985273 == array_index_948961 ? add_985589 : sel_985586;
  assign add_985593 = sel_985590 + 8'h01;
  assign sel_985594 = array_index_985273 == array_index_948967 ? add_985593 : sel_985590;
  assign add_985597 = sel_985594 + 8'h01;
  assign sel_985598 = array_index_985273 == array_index_948973 ? add_985597 : sel_985594;
  assign add_985601 = sel_985598 + 8'h01;
  assign sel_985602 = array_index_985273 == array_index_948979 ? add_985601 : sel_985598;
  assign add_985605 = sel_985602 + 8'h01;
  assign sel_985606 = array_index_985273 == array_index_948985 ? add_985605 : sel_985602;
  assign add_985609 = sel_985606 + 8'h01;
  assign sel_985610 = array_index_985273 == array_index_948991 ? add_985609 : sel_985606;
  assign add_985613 = sel_985610 + 8'h01;
  assign sel_985614 = array_index_985273 == array_index_948997 ? add_985613 : sel_985610;
  assign add_985617 = sel_985614 + 8'h01;
  assign sel_985618 = array_index_985273 == array_index_949003 ? add_985617 : sel_985614;
  assign add_985621 = sel_985618 + 8'h01;
  assign sel_985622 = array_index_985273 == array_index_949009 ? add_985621 : sel_985618;
  assign add_985625 = sel_985622 + 8'h01;
  assign sel_985626 = array_index_985273 == array_index_949015 ? add_985625 : sel_985622;
  assign add_985629 = sel_985626 + 8'h01;
  assign sel_985630 = array_index_985273 == array_index_949021 ? add_985629 : sel_985626;
  assign add_985633 = sel_985630 + 8'h01;
  assign sel_985634 = array_index_985273 == array_index_949027 ? add_985633 : sel_985630;
  assign add_985637 = sel_985634 + 8'h01;
  assign sel_985638 = array_index_985273 == array_index_949033 ? add_985637 : sel_985634;
  assign add_985641 = sel_985638 + 8'h01;
  assign sel_985642 = array_index_985273 == array_index_949039 ? add_985641 : sel_985638;
  assign add_985645 = sel_985642 + 8'h01;
  assign sel_985646 = array_index_985273 == array_index_949045 ? add_985645 : sel_985642;
  assign add_985649 = sel_985646 + 8'h01;
  assign sel_985650 = array_index_985273 == array_index_949051 ? add_985649 : sel_985646;
  assign add_985653 = sel_985650 + 8'h01;
  assign sel_985654 = array_index_985273 == array_index_949057 ? add_985653 : sel_985650;
  assign add_985657 = sel_985654 + 8'h01;
  assign sel_985658 = array_index_985273 == array_index_949063 ? add_985657 : sel_985654;
  assign add_985661 = sel_985658 + 8'h01;
  assign sel_985662 = array_index_985273 == array_index_949069 ? add_985661 : sel_985658;
  assign add_985665 = sel_985662 + 8'h01;
  assign sel_985666 = array_index_985273 == array_index_949075 ? add_985665 : sel_985662;
  assign add_985669 = sel_985666 + 8'h01;
  assign sel_985670 = array_index_985273 == array_index_949081 ? add_985669 : sel_985666;
  assign add_985674 = sel_985670 + 8'h01;
  assign array_index_985675 = set1_unflattened[7'h5c];
  assign sel_985676 = array_index_985273 == array_index_949087 ? add_985674 : sel_985670;
  assign add_985679 = sel_985676 + 8'h01;
  assign sel_985680 = array_index_985675 == array_index_948483 ? add_985679 : sel_985676;
  assign add_985683 = sel_985680 + 8'h01;
  assign sel_985684 = array_index_985675 == array_index_948487 ? add_985683 : sel_985680;
  assign add_985687 = sel_985684 + 8'h01;
  assign sel_985688 = array_index_985675 == array_index_948495 ? add_985687 : sel_985684;
  assign add_985691 = sel_985688 + 8'h01;
  assign sel_985692 = array_index_985675 == array_index_948503 ? add_985691 : sel_985688;
  assign add_985695 = sel_985692 + 8'h01;
  assign sel_985696 = array_index_985675 == array_index_948511 ? add_985695 : sel_985692;
  assign add_985699 = sel_985696 + 8'h01;
  assign sel_985700 = array_index_985675 == array_index_948519 ? add_985699 : sel_985696;
  assign add_985703 = sel_985700 + 8'h01;
  assign sel_985704 = array_index_985675 == array_index_948527 ? add_985703 : sel_985700;
  assign add_985707 = sel_985704 + 8'h01;
  assign sel_985708 = array_index_985675 == array_index_948535 ? add_985707 : sel_985704;
  assign add_985711 = sel_985708 + 8'h01;
  assign sel_985712 = array_index_985675 == array_index_948541 ? add_985711 : sel_985708;
  assign add_985715 = sel_985712 + 8'h01;
  assign sel_985716 = array_index_985675 == array_index_948547 ? add_985715 : sel_985712;
  assign add_985719 = sel_985716 + 8'h01;
  assign sel_985720 = array_index_985675 == array_index_948553 ? add_985719 : sel_985716;
  assign add_985723 = sel_985720 + 8'h01;
  assign sel_985724 = array_index_985675 == array_index_948559 ? add_985723 : sel_985720;
  assign add_985727 = sel_985724 + 8'h01;
  assign sel_985728 = array_index_985675 == array_index_948565 ? add_985727 : sel_985724;
  assign add_985731 = sel_985728 + 8'h01;
  assign sel_985732 = array_index_985675 == array_index_948571 ? add_985731 : sel_985728;
  assign add_985735 = sel_985732 + 8'h01;
  assign sel_985736 = array_index_985675 == array_index_948577 ? add_985735 : sel_985732;
  assign add_985739 = sel_985736 + 8'h01;
  assign sel_985740 = array_index_985675 == array_index_948583 ? add_985739 : sel_985736;
  assign add_985743 = sel_985740 + 8'h01;
  assign sel_985744 = array_index_985675 == array_index_948589 ? add_985743 : sel_985740;
  assign add_985747 = sel_985744 + 8'h01;
  assign sel_985748 = array_index_985675 == array_index_948595 ? add_985747 : sel_985744;
  assign add_985751 = sel_985748 + 8'h01;
  assign sel_985752 = array_index_985675 == array_index_948601 ? add_985751 : sel_985748;
  assign add_985755 = sel_985752 + 8'h01;
  assign sel_985756 = array_index_985675 == array_index_948607 ? add_985755 : sel_985752;
  assign add_985759 = sel_985756 + 8'h01;
  assign sel_985760 = array_index_985675 == array_index_948613 ? add_985759 : sel_985756;
  assign add_985763 = sel_985760 + 8'h01;
  assign sel_985764 = array_index_985675 == array_index_948619 ? add_985763 : sel_985760;
  assign add_985767 = sel_985764 + 8'h01;
  assign sel_985768 = array_index_985675 == array_index_948625 ? add_985767 : sel_985764;
  assign add_985771 = sel_985768 + 8'h01;
  assign sel_985772 = array_index_985675 == array_index_948631 ? add_985771 : sel_985768;
  assign add_985775 = sel_985772 + 8'h01;
  assign sel_985776 = array_index_985675 == array_index_948637 ? add_985775 : sel_985772;
  assign add_985779 = sel_985776 + 8'h01;
  assign sel_985780 = array_index_985675 == array_index_948643 ? add_985779 : sel_985776;
  assign add_985783 = sel_985780 + 8'h01;
  assign sel_985784 = array_index_985675 == array_index_948649 ? add_985783 : sel_985780;
  assign add_985787 = sel_985784 + 8'h01;
  assign sel_985788 = array_index_985675 == array_index_948655 ? add_985787 : sel_985784;
  assign add_985791 = sel_985788 + 8'h01;
  assign sel_985792 = array_index_985675 == array_index_948661 ? add_985791 : sel_985788;
  assign add_985795 = sel_985792 + 8'h01;
  assign sel_985796 = array_index_985675 == array_index_948667 ? add_985795 : sel_985792;
  assign add_985799 = sel_985796 + 8'h01;
  assign sel_985800 = array_index_985675 == array_index_948673 ? add_985799 : sel_985796;
  assign add_985803 = sel_985800 + 8'h01;
  assign sel_985804 = array_index_985675 == array_index_948679 ? add_985803 : sel_985800;
  assign add_985807 = sel_985804 + 8'h01;
  assign sel_985808 = array_index_985675 == array_index_948685 ? add_985807 : sel_985804;
  assign add_985811 = sel_985808 + 8'h01;
  assign sel_985812 = array_index_985675 == array_index_948691 ? add_985811 : sel_985808;
  assign add_985815 = sel_985812 + 8'h01;
  assign sel_985816 = array_index_985675 == array_index_948697 ? add_985815 : sel_985812;
  assign add_985819 = sel_985816 + 8'h01;
  assign sel_985820 = array_index_985675 == array_index_948703 ? add_985819 : sel_985816;
  assign add_985823 = sel_985820 + 8'h01;
  assign sel_985824 = array_index_985675 == array_index_948709 ? add_985823 : sel_985820;
  assign add_985827 = sel_985824 + 8'h01;
  assign sel_985828 = array_index_985675 == array_index_948715 ? add_985827 : sel_985824;
  assign add_985831 = sel_985828 + 8'h01;
  assign sel_985832 = array_index_985675 == array_index_948721 ? add_985831 : sel_985828;
  assign add_985835 = sel_985832 + 8'h01;
  assign sel_985836 = array_index_985675 == array_index_948727 ? add_985835 : sel_985832;
  assign add_985839 = sel_985836 + 8'h01;
  assign sel_985840 = array_index_985675 == array_index_948733 ? add_985839 : sel_985836;
  assign add_985843 = sel_985840 + 8'h01;
  assign sel_985844 = array_index_985675 == array_index_948739 ? add_985843 : sel_985840;
  assign add_985847 = sel_985844 + 8'h01;
  assign sel_985848 = array_index_985675 == array_index_948745 ? add_985847 : sel_985844;
  assign add_985851 = sel_985848 + 8'h01;
  assign sel_985852 = array_index_985675 == array_index_948751 ? add_985851 : sel_985848;
  assign add_985855 = sel_985852 + 8'h01;
  assign sel_985856 = array_index_985675 == array_index_948757 ? add_985855 : sel_985852;
  assign add_985859 = sel_985856 + 8'h01;
  assign sel_985860 = array_index_985675 == array_index_948763 ? add_985859 : sel_985856;
  assign add_985863 = sel_985860 + 8'h01;
  assign sel_985864 = array_index_985675 == array_index_948769 ? add_985863 : sel_985860;
  assign add_985867 = sel_985864 + 8'h01;
  assign sel_985868 = array_index_985675 == array_index_948775 ? add_985867 : sel_985864;
  assign add_985871 = sel_985868 + 8'h01;
  assign sel_985872 = array_index_985675 == array_index_948781 ? add_985871 : sel_985868;
  assign add_985875 = sel_985872 + 8'h01;
  assign sel_985876 = array_index_985675 == array_index_948787 ? add_985875 : sel_985872;
  assign add_985879 = sel_985876 + 8'h01;
  assign sel_985880 = array_index_985675 == array_index_948793 ? add_985879 : sel_985876;
  assign add_985883 = sel_985880 + 8'h01;
  assign sel_985884 = array_index_985675 == array_index_948799 ? add_985883 : sel_985880;
  assign add_985887 = sel_985884 + 8'h01;
  assign sel_985888 = array_index_985675 == array_index_948805 ? add_985887 : sel_985884;
  assign add_985891 = sel_985888 + 8'h01;
  assign sel_985892 = array_index_985675 == array_index_948811 ? add_985891 : sel_985888;
  assign add_985895 = sel_985892 + 8'h01;
  assign sel_985896 = array_index_985675 == array_index_948817 ? add_985895 : sel_985892;
  assign add_985899 = sel_985896 + 8'h01;
  assign sel_985900 = array_index_985675 == array_index_948823 ? add_985899 : sel_985896;
  assign add_985903 = sel_985900 + 8'h01;
  assign sel_985904 = array_index_985675 == array_index_948829 ? add_985903 : sel_985900;
  assign add_985907 = sel_985904 + 8'h01;
  assign sel_985908 = array_index_985675 == array_index_948835 ? add_985907 : sel_985904;
  assign add_985911 = sel_985908 + 8'h01;
  assign sel_985912 = array_index_985675 == array_index_948841 ? add_985911 : sel_985908;
  assign add_985915 = sel_985912 + 8'h01;
  assign sel_985916 = array_index_985675 == array_index_948847 ? add_985915 : sel_985912;
  assign add_985919 = sel_985916 + 8'h01;
  assign sel_985920 = array_index_985675 == array_index_948853 ? add_985919 : sel_985916;
  assign add_985923 = sel_985920 + 8'h01;
  assign sel_985924 = array_index_985675 == array_index_948859 ? add_985923 : sel_985920;
  assign add_985927 = sel_985924 + 8'h01;
  assign sel_985928 = array_index_985675 == array_index_948865 ? add_985927 : sel_985924;
  assign add_985931 = sel_985928 + 8'h01;
  assign sel_985932 = array_index_985675 == array_index_948871 ? add_985931 : sel_985928;
  assign add_985935 = sel_985932 + 8'h01;
  assign sel_985936 = array_index_985675 == array_index_948877 ? add_985935 : sel_985932;
  assign add_985939 = sel_985936 + 8'h01;
  assign sel_985940 = array_index_985675 == array_index_948883 ? add_985939 : sel_985936;
  assign add_985943 = sel_985940 + 8'h01;
  assign sel_985944 = array_index_985675 == array_index_948889 ? add_985943 : sel_985940;
  assign add_985947 = sel_985944 + 8'h01;
  assign sel_985948 = array_index_985675 == array_index_948895 ? add_985947 : sel_985944;
  assign add_985951 = sel_985948 + 8'h01;
  assign sel_985952 = array_index_985675 == array_index_948901 ? add_985951 : sel_985948;
  assign add_985955 = sel_985952 + 8'h01;
  assign sel_985956 = array_index_985675 == array_index_948907 ? add_985955 : sel_985952;
  assign add_985959 = sel_985956 + 8'h01;
  assign sel_985960 = array_index_985675 == array_index_948913 ? add_985959 : sel_985956;
  assign add_985963 = sel_985960 + 8'h01;
  assign sel_985964 = array_index_985675 == array_index_948919 ? add_985963 : sel_985960;
  assign add_985967 = sel_985964 + 8'h01;
  assign sel_985968 = array_index_985675 == array_index_948925 ? add_985967 : sel_985964;
  assign add_985971 = sel_985968 + 8'h01;
  assign sel_985972 = array_index_985675 == array_index_948931 ? add_985971 : sel_985968;
  assign add_985975 = sel_985972 + 8'h01;
  assign sel_985976 = array_index_985675 == array_index_948937 ? add_985975 : sel_985972;
  assign add_985979 = sel_985976 + 8'h01;
  assign sel_985980 = array_index_985675 == array_index_948943 ? add_985979 : sel_985976;
  assign add_985983 = sel_985980 + 8'h01;
  assign sel_985984 = array_index_985675 == array_index_948949 ? add_985983 : sel_985980;
  assign add_985987 = sel_985984 + 8'h01;
  assign sel_985988 = array_index_985675 == array_index_948955 ? add_985987 : sel_985984;
  assign add_985991 = sel_985988 + 8'h01;
  assign sel_985992 = array_index_985675 == array_index_948961 ? add_985991 : sel_985988;
  assign add_985995 = sel_985992 + 8'h01;
  assign sel_985996 = array_index_985675 == array_index_948967 ? add_985995 : sel_985992;
  assign add_985999 = sel_985996 + 8'h01;
  assign sel_986000 = array_index_985675 == array_index_948973 ? add_985999 : sel_985996;
  assign add_986003 = sel_986000 + 8'h01;
  assign sel_986004 = array_index_985675 == array_index_948979 ? add_986003 : sel_986000;
  assign add_986007 = sel_986004 + 8'h01;
  assign sel_986008 = array_index_985675 == array_index_948985 ? add_986007 : sel_986004;
  assign add_986011 = sel_986008 + 8'h01;
  assign sel_986012 = array_index_985675 == array_index_948991 ? add_986011 : sel_986008;
  assign add_986015 = sel_986012 + 8'h01;
  assign sel_986016 = array_index_985675 == array_index_948997 ? add_986015 : sel_986012;
  assign add_986019 = sel_986016 + 8'h01;
  assign sel_986020 = array_index_985675 == array_index_949003 ? add_986019 : sel_986016;
  assign add_986023 = sel_986020 + 8'h01;
  assign sel_986024 = array_index_985675 == array_index_949009 ? add_986023 : sel_986020;
  assign add_986027 = sel_986024 + 8'h01;
  assign sel_986028 = array_index_985675 == array_index_949015 ? add_986027 : sel_986024;
  assign add_986031 = sel_986028 + 8'h01;
  assign sel_986032 = array_index_985675 == array_index_949021 ? add_986031 : sel_986028;
  assign add_986035 = sel_986032 + 8'h01;
  assign sel_986036 = array_index_985675 == array_index_949027 ? add_986035 : sel_986032;
  assign add_986039 = sel_986036 + 8'h01;
  assign sel_986040 = array_index_985675 == array_index_949033 ? add_986039 : sel_986036;
  assign add_986043 = sel_986040 + 8'h01;
  assign sel_986044 = array_index_985675 == array_index_949039 ? add_986043 : sel_986040;
  assign add_986047 = sel_986044 + 8'h01;
  assign sel_986048 = array_index_985675 == array_index_949045 ? add_986047 : sel_986044;
  assign add_986051 = sel_986048 + 8'h01;
  assign sel_986052 = array_index_985675 == array_index_949051 ? add_986051 : sel_986048;
  assign add_986055 = sel_986052 + 8'h01;
  assign sel_986056 = array_index_985675 == array_index_949057 ? add_986055 : sel_986052;
  assign add_986059 = sel_986056 + 8'h01;
  assign sel_986060 = array_index_985675 == array_index_949063 ? add_986059 : sel_986056;
  assign add_986063 = sel_986060 + 8'h01;
  assign sel_986064 = array_index_985675 == array_index_949069 ? add_986063 : sel_986060;
  assign add_986067 = sel_986064 + 8'h01;
  assign sel_986068 = array_index_985675 == array_index_949075 ? add_986067 : sel_986064;
  assign add_986071 = sel_986068 + 8'h01;
  assign sel_986072 = array_index_985675 == array_index_949081 ? add_986071 : sel_986068;
  assign add_986076 = sel_986072 + 8'h01;
  assign array_index_986077 = set1_unflattened[7'h5d];
  assign sel_986078 = array_index_985675 == array_index_949087 ? add_986076 : sel_986072;
  assign add_986081 = sel_986078 + 8'h01;
  assign sel_986082 = array_index_986077 == array_index_948483 ? add_986081 : sel_986078;
  assign add_986085 = sel_986082 + 8'h01;
  assign sel_986086 = array_index_986077 == array_index_948487 ? add_986085 : sel_986082;
  assign add_986089 = sel_986086 + 8'h01;
  assign sel_986090 = array_index_986077 == array_index_948495 ? add_986089 : sel_986086;
  assign add_986093 = sel_986090 + 8'h01;
  assign sel_986094 = array_index_986077 == array_index_948503 ? add_986093 : sel_986090;
  assign add_986097 = sel_986094 + 8'h01;
  assign sel_986098 = array_index_986077 == array_index_948511 ? add_986097 : sel_986094;
  assign add_986101 = sel_986098 + 8'h01;
  assign sel_986102 = array_index_986077 == array_index_948519 ? add_986101 : sel_986098;
  assign add_986105 = sel_986102 + 8'h01;
  assign sel_986106 = array_index_986077 == array_index_948527 ? add_986105 : sel_986102;
  assign add_986109 = sel_986106 + 8'h01;
  assign sel_986110 = array_index_986077 == array_index_948535 ? add_986109 : sel_986106;
  assign add_986113 = sel_986110 + 8'h01;
  assign sel_986114 = array_index_986077 == array_index_948541 ? add_986113 : sel_986110;
  assign add_986117 = sel_986114 + 8'h01;
  assign sel_986118 = array_index_986077 == array_index_948547 ? add_986117 : sel_986114;
  assign add_986121 = sel_986118 + 8'h01;
  assign sel_986122 = array_index_986077 == array_index_948553 ? add_986121 : sel_986118;
  assign add_986125 = sel_986122 + 8'h01;
  assign sel_986126 = array_index_986077 == array_index_948559 ? add_986125 : sel_986122;
  assign add_986129 = sel_986126 + 8'h01;
  assign sel_986130 = array_index_986077 == array_index_948565 ? add_986129 : sel_986126;
  assign add_986133 = sel_986130 + 8'h01;
  assign sel_986134 = array_index_986077 == array_index_948571 ? add_986133 : sel_986130;
  assign add_986137 = sel_986134 + 8'h01;
  assign sel_986138 = array_index_986077 == array_index_948577 ? add_986137 : sel_986134;
  assign add_986141 = sel_986138 + 8'h01;
  assign sel_986142 = array_index_986077 == array_index_948583 ? add_986141 : sel_986138;
  assign add_986145 = sel_986142 + 8'h01;
  assign sel_986146 = array_index_986077 == array_index_948589 ? add_986145 : sel_986142;
  assign add_986149 = sel_986146 + 8'h01;
  assign sel_986150 = array_index_986077 == array_index_948595 ? add_986149 : sel_986146;
  assign add_986153 = sel_986150 + 8'h01;
  assign sel_986154 = array_index_986077 == array_index_948601 ? add_986153 : sel_986150;
  assign add_986157 = sel_986154 + 8'h01;
  assign sel_986158 = array_index_986077 == array_index_948607 ? add_986157 : sel_986154;
  assign add_986161 = sel_986158 + 8'h01;
  assign sel_986162 = array_index_986077 == array_index_948613 ? add_986161 : sel_986158;
  assign add_986165 = sel_986162 + 8'h01;
  assign sel_986166 = array_index_986077 == array_index_948619 ? add_986165 : sel_986162;
  assign add_986169 = sel_986166 + 8'h01;
  assign sel_986170 = array_index_986077 == array_index_948625 ? add_986169 : sel_986166;
  assign add_986173 = sel_986170 + 8'h01;
  assign sel_986174 = array_index_986077 == array_index_948631 ? add_986173 : sel_986170;
  assign add_986177 = sel_986174 + 8'h01;
  assign sel_986178 = array_index_986077 == array_index_948637 ? add_986177 : sel_986174;
  assign add_986181 = sel_986178 + 8'h01;
  assign sel_986182 = array_index_986077 == array_index_948643 ? add_986181 : sel_986178;
  assign add_986185 = sel_986182 + 8'h01;
  assign sel_986186 = array_index_986077 == array_index_948649 ? add_986185 : sel_986182;
  assign add_986189 = sel_986186 + 8'h01;
  assign sel_986190 = array_index_986077 == array_index_948655 ? add_986189 : sel_986186;
  assign add_986193 = sel_986190 + 8'h01;
  assign sel_986194 = array_index_986077 == array_index_948661 ? add_986193 : sel_986190;
  assign add_986197 = sel_986194 + 8'h01;
  assign sel_986198 = array_index_986077 == array_index_948667 ? add_986197 : sel_986194;
  assign add_986201 = sel_986198 + 8'h01;
  assign sel_986202 = array_index_986077 == array_index_948673 ? add_986201 : sel_986198;
  assign add_986205 = sel_986202 + 8'h01;
  assign sel_986206 = array_index_986077 == array_index_948679 ? add_986205 : sel_986202;
  assign add_986209 = sel_986206 + 8'h01;
  assign sel_986210 = array_index_986077 == array_index_948685 ? add_986209 : sel_986206;
  assign add_986213 = sel_986210 + 8'h01;
  assign sel_986214 = array_index_986077 == array_index_948691 ? add_986213 : sel_986210;
  assign add_986217 = sel_986214 + 8'h01;
  assign sel_986218 = array_index_986077 == array_index_948697 ? add_986217 : sel_986214;
  assign add_986221 = sel_986218 + 8'h01;
  assign sel_986222 = array_index_986077 == array_index_948703 ? add_986221 : sel_986218;
  assign add_986225 = sel_986222 + 8'h01;
  assign sel_986226 = array_index_986077 == array_index_948709 ? add_986225 : sel_986222;
  assign add_986229 = sel_986226 + 8'h01;
  assign sel_986230 = array_index_986077 == array_index_948715 ? add_986229 : sel_986226;
  assign add_986233 = sel_986230 + 8'h01;
  assign sel_986234 = array_index_986077 == array_index_948721 ? add_986233 : sel_986230;
  assign add_986237 = sel_986234 + 8'h01;
  assign sel_986238 = array_index_986077 == array_index_948727 ? add_986237 : sel_986234;
  assign add_986241 = sel_986238 + 8'h01;
  assign sel_986242 = array_index_986077 == array_index_948733 ? add_986241 : sel_986238;
  assign add_986245 = sel_986242 + 8'h01;
  assign sel_986246 = array_index_986077 == array_index_948739 ? add_986245 : sel_986242;
  assign add_986249 = sel_986246 + 8'h01;
  assign sel_986250 = array_index_986077 == array_index_948745 ? add_986249 : sel_986246;
  assign add_986253 = sel_986250 + 8'h01;
  assign sel_986254 = array_index_986077 == array_index_948751 ? add_986253 : sel_986250;
  assign add_986257 = sel_986254 + 8'h01;
  assign sel_986258 = array_index_986077 == array_index_948757 ? add_986257 : sel_986254;
  assign add_986261 = sel_986258 + 8'h01;
  assign sel_986262 = array_index_986077 == array_index_948763 ? add_986261 : sel_986258;
  assign add_986265 = sel_986262 + 8'h01;
  assign sel_986266 = array_index_986077 == array_index_948769 ? add_986265 : sel_986262;
  assign add_986269 = sel_986266 + 8'h01;
  assign sel_986270 = array_index_986077 == array_index_948775 ? add_986269 : sel_986266;
  assign add_986273 = sel_986270 + 8'h01;
  assign sel_986274 = array_index_986077 == array_index_948781 ? add_986273 : sel_986270;
  assign add_986277 = sel_986274 + 8'h01;
  assign sel_986278 = array_index_986077 == array_index_948787 ? add_986277 : sel_986274;
  assign add_986281 = sel_986278 + 8'h01;
  assign sel_986282 = array_index_986077 == array_index_948793 ? add_986281 : sel_986278;
  assign add_986285 = sel_986282 + 8'h01;
  assign sel_986286 = array_index_986077 == array_index_948799 ? add_986285 : sel_986282;
  assign add_986289 = sel_986286 + 8'h01;
  assign sel_986290 = array_index_986077 == array_index_948805 ? add_986289 : sel_986286;
  assign add_986293 = sel_986290 + 8'h01;
  assign sel_986294 = array_index_986077 == array_index_948811 ? add_986293 : sel_986290;
  assign add_986297 = sel_986294 + 8'h01;
  assign sel_986298 = array_index_986077 == array_index_948817 ? add_986297 : sel_986294;
  assign add_986301 = sel_986298 + 8'h01;
  assign sel_986302 = array_index_986077 == array_index_948823 ? add_986301 : sel_986298;
  assign add_986305 = sel_986302 + 8'h01;
  assign sel_986306 = array_index_986077 == array_index_948829 ? add_986305 : sel_986302;
  assign add_986309 = sel_986306 + 8'h01;
  assign sel_986310 = array_index_986077 == array_index_948835 ? add_986309 : sel_986306;
  assign add_986313 = sel_986310 + 8'h01;
  assign sel_986314 = array_index_986077 == array_index_948841 ? add_986313 : sel_986310;
  assign add_986317 = sel_986314 + 8'h01;
  assign sel_986318 = array_index_986077 == array_index_948847 ? add_986317 : sel_986314;
  assign add_986321 = sel_986318 + 8'h01;
  assign sel_986322 = array_index_986077 == array_index_948853 ? add_986321 : sel_986318;
  assign add_986325 = sel_986322 + 8'h01;
  assign sel_986326 = array_index_986077 == array_index_948859 ? add_986325 : sel_986322;
  assign add_986329 = sel_986326 + 8'h01;
  assign sel_986330 = array_index_986077 == array_index_948865 ? add_986329 : sel_986326;
  assign add_986333 = sel_986330 + 8'h01;
  assign sel_986334 = array_index_986077 == array_index_948871 ? add_986333 : sel_986330;
  assign add_986337 = sel_986334 + 8'h01;
  assign sel_986338 = array_index_986077 == array_index_948877 ? add_986337 : sel_986334;
  assign add_986341 = sel_986338 + 8'h01;
  assign sel_986342 = array_index_986077 == array_index_948883 ? add_986341 : sel_986338;
  assign add_986345 = sel_986342 + 8'h01;
  assign sel_986346 = array_index_986077 == array_index_948889 ? add_986345 : sel_986342;
  assign add_986349 = sel_986346 + 8'h01;
  assign sel_986350 = array_index_986077 == array_index_948895 ? add_986349 : sel_986346;
  assign add_986353 = sel_986350 + 8'h01;
  assign sel_986354 = array_index_986077 == array_index_948901 ? add_986353 : sel_986350;
  assign add_986357 = sel_986354 + 8'h01;
  assign sel_986358 = array_index_986077 == array_index_948907 ? add_986357 : sel_986354;
  assign add_986361 = sel_986358 + 8'h01;
  assign sel_986362 = array_index_986077 == array_index_948913 ? add_986361 : sel_986358;
  assign add_986365 = sel_986362 + 8'h01;
  assign sel_986366 = array_index_986077 == array_index_948919 ? add_986365 : sel_986362;
  assign add_986369 = sel_986366 + 8'h01;
  assign sel_986370 = array_index_986077 == array_index_948925 ? add_986369 : sel_986366;
  assign add_986373 = sel_986370 + 8'h01;
  assign sel_986374 = array_index_986077 == array_index_948931 ? add_986373 : sel_986370;
  assign add_986377 = sel_986374 + 8'h01;
  assign sel_986378 = array_index_986077 == array_index_948937 ? add_986377 : sel_986374;
  assign add_986381 = sel_986378 + 8'h01;
  assign sel_986382 = array_index_986077 == array_index_948943 ? add_986381 : sel_986378;
  assign add_986385 = sel_986382 + 8'h01;
  assign sel_986386 = array_index_986077 == array_index_948949 ? add_986385 : sel_986382;
  assign add_986389 = sel_986386 + 8'h01;
  assign sel_986390 = array_index_986077 == array_index_948955 ? add_986389 : sel_986386;
  assign add_986393 = sel_986390 + 8'h01;
  assign sel_986394 = array_index_986077 == array_index_948961 ? add_986393 : sel_986390;
  assign add_986397 = sel_986394 + 8'h01;
  assign sel_986398 = array_index_986077 == array_index_948967 ? add_986397 : sel_986394;
  assign add_986401 = sel_986398 + 8'h01;
  assign sel_986402 = array_index_986077 == array_index_948973 ? add_986401 : sel_986398;
  assign add_986405 = sel_986402 + 8'h01;
  assign sel_986406 = array_index_986077 == array_index_948979 ? add_986405 : sel_986402;
  assign add_986409 = sel_986406 + 8'h01;
  assign sel_986410 = array_index_986077 == array_index_948985 ? add_986409 : sel_986406;
  assign add_986413 = sel_986410 + 8'h01;
  assign sel_986414 = array_index_986077 == array_index_948991 ? add_986413 : sel_986410;
  assign add_986417 = sel_986414 + 8'h01;
  assign sel_986418 = array_index_986077 == array_index_948997 ? add_986417 : sel_986414;
  assign add_986421 = sel_986418 + 8'h01;
  assign sel_986422 = array_index_986077 == array_index_949003 ? add_986421 : sel_986418;
  assign add_986425 = sel_986422 + 8'h01;
  assign sel_986426 = array_index_986077 == array_index_949009 ? add_986425 : sel_986422;
  assign add_986429 = sel_986426 + 8'h01;
  assign sel_986430 = array_index_986077 == array_index_949015 ? add_986429 : sel_986426;
  assign add_986433 = sel_986430 + 8'h01;
  assign sel_986434 = array_index_986077 == array_index_949021 ? add_986433 : sel_986430;
  assign add_986437 = sel_986434 + 8'h01;
  assign sel_986438 = array_index_986077 == array_index_949027 ? add_986437 : sel_986434;
  assign add_986441 = sel_986438 + 8'h01;
  assign sel_986442 = array_index_986077 == array_index_949033 ? add_986441 : sel_986438;
  assign add_986445 = sel_986442 + 8'h01;
  assign sel_986446 = array_index_986077 == array_index_949039 ? add_986445 : sel_986442;
  assign add_986449 = sel_986446 + 8'h01;
  assign sel_986450 = array_index_986077 == array_index_949045 ? add_986449 : sel_986446;
  assign add_986453 = sel_986450 + 8'h01;
  assign sel_986454 = array_index_986077 == array_index_949051 ? add_986453 : sel_986450;
  assign add_986457 = sel_986454 + 8'h01;
  assign sel_986458 = array_index_986077 == array_index_949057 ? add_986457 : sel_986454;
  assign add_986461 = sel_986458 + 8'h01;
  assign sel_986462 = array_index_986077 == array_index_949063 ? add_986461 : sel_986458;
  assign add_986465 = sel_986462 + 8'h01;
  assign sel_986466 = array_index_986077 == array_index_949069 ? add_986465 : sel_986462;
  assign add_986469 = sel_986466 + 8'h01;
  assign sel_986470 = array_index_986077 == array_index_949075 ? add_986469 : sel_986466;
  assign add_986473 = sel_986470 + 8'h01;
  assign sel_986474 = array_index_986077 == array_index_949081 ? add_986473 : sel_986470;
  assign add_986478 = sel_986474 + 8'h01;
  assign array_index_986479 = set1_unflattened[7'h5e];
  assign sel_986480 = array_index_986077 == array_index_949087 ? add_986478 : sel_986474;
  assign add_986483 = sel_986480 + 8'h01;
  assign sel_986484 = array_index_986479 == array_index_948483 ? add_986483 : sel_986480;
  assign add_986487 = sel_986484 + 8'h01;
  assign sel_986488 = array_index_986479 == array_index_948487 ? add_986487 : sel_986484;
  assign add_986491 = sel_986488 + 8'h01;
  assign sel_986492 = array_index_986479 == array_index_948495 ? add_986491 : sel_986488;
  assign add_986495 = sel_986492 + 8'h01;
  assign sel_986496 = array_index_986479 == array_index_948503 ? add_986495 : sel_986492;
  assign add_986499 = sel_986496 + 8'h01;
  assign sel_986500 = array_index_986479 == array_index_948511 ? add_986499 : sel_986496;
  assign add_986503 = sel_986500 + 8'h01;
  assign sel_986504 = array_index_986479 == array_index_948519 ? add_986503 : sel_986500;
  assign add_986507 = sel_986504 + 8'h01;
  assign sel_986508 = array_index_986479 == array_index_948527 ? add_986507 : sel_986504;
  assign add_986511 = sel_986508 + 8'h01;
  assign sel_986512 = array_index_986479 == array_index_948535 ? add_986511 : sel_986508;
  assign add_986515 = sel_986512 + 8'h01;
  assign sel_986516 = array_index_986479 == array_index_948541 ? add_986515 : sel_986512;
  assign add_986519 = sel_986516 + 8'h01;
  assign sel_986520 = array_index_986479 == array_index_948547 ? add_986519 : sel_986516;
  assign add_986523 = sel_986520 + 8'h01;
  assign sel_986524 = array_index_986479 == array_index_948553 ? add_986523 : sel_986520;
  assign add_986527 = sel_986524 + 8'h01;
  assign sel_986528 = array_index_986479 == array_index_948559 ? add_986527 : sel_986524;
  assign add_986531 = sel_986528 + 8'h01;
  assign sel_986532 = array_index_986479 == array_index_948565 ? add_986531 : sel_986528;
  assign add_986535 = sel_986532 + 8'h01;
  assign sel_986536 = array_index_986479 == array_index_948571 ? add_986535 : sel_986532;
  assign add_986539 = sel_986536 + 8'h01;
  assign sel_986540 = array_index_986479 == array_index_948577 ? add_986539 : sel_986536;
  assign add_986543 = sel_986540 + 8'h01;
  assign sel_986544 = array_index_986479 == array_index_948583 ? add_986543 : sel_986540;
  assign add_986547 = sel_986544 + 8'h01;
  assign sel_986548 = array_index_986479 == array_index_948589 ? add_986547 : sel_986544;
  assign add_986551 = sel_986548 + 8'h01;
  assign sel_986552 = array_index_986479 == array_index_948595 ? add_986551 : sel_986548;
  assign add_986555 = sel_986552 + 8'h01;
  assign sel_986556 = array_index_986479 == array_index_948601 ? add_986555 : sel_986552;
  assign add_986559 = sel_986556 + 8'h01;
  assign sel_986560 = array_index_986479 == array_index_948607 ? add_986559 : sel_986556;
  assign add_986563 = sel_986560 + 8'h01;
  assign sel_986564 = array_index_986479 == array_index_948613 ? add_986563 : sel_986560;
  assign add_986567 = sel_986564 + 8'h01;
  assign sel_986568 = array_index_986479 == array_index_948619 ? add_986567 : sel_986564;
  assign add_986571 = sel_986568 + 8'h01;
  assign sel_986572 = array_index_986479 == array_index_948625 ? add_986571 : sel_986568;
  assign add_986575 = sel_986572 + 8'h01;
  assign sel_986576 = array_index_986479 == array_index_948631 ? add_986575 : sel_986572;
  assign add_986579 = sel_986576 + 8'h01;
  assign sel_986580 = array_index_986479 == array_index_948637 ? add_986579 : sel_986576;
  assign add_986583 = sel_986580 + 8'h01;
  assign sel_986584 = array_index_986479 == array_index_948643 ? add_986583 : sel_986580;
  assign add_986587 = sel_986584 + 8'h01;
  assign sel_986588 = array_index_986479 == array_index_948649 ? add_986587 : sel_986584;
  assign add_986591 = sel_986588 + 8'h01;
  assign sel_986592 = array_index_986479 == array_index_948655 ? add_986591 : sel_986588;
  assign add_986595 = sel_986592 + 8'h01;
  assign sel_986596 = array_index_986479 == array_index_948661 ? add_986595 : sel_986592;
  assign add_986599 = sel_986596 + 8'h01;
  assign sel_986600 = array_index_986479 == array_index_948667 ? add_986599 : sel_986596;
  assign add_986603 = sel_986600 + 8'h01;
  assign sel_986604 = array_index_986479 == array_index_948673 ? add_986603 : sel_986600;
  assign add_986607 = sel_986604 + 8'h01;
  assign sel_986608 = array_index_986479 == array_index_948679 ? add_986607 : sel_986604;
  assign add_986611 = sel_986608 + 8'h01;
  assign sel_986612 = array_index_986479 == array_index_948685 ? add_986611 : sel_986608;
  assign add_986615 = sel_986612 + 8'h01;
  assign sel_986616 = array_index_986479 == array_index_948691 ? add_986615 : sel_986612;
  assign add_986619 = sel_986616 + 8'h01;
  assign sel_986620 = array_index_986479 == array_index_948697 ? add_986619 : sel_986616;
  assign add_986623 = sel_986620 + 8'h01;
  assign sel_986624 = array_index_986479 == array_index_948703 ? add_986623 : sel_986620;
  assign add_986627 = sel_986624 + 8'h01;
  assign sel_986628 = array_index_986479 == array_index_948709 ? add_986627 : sel_986624;
  assign add_986631 = sel_986628 + 8'h01;
  assign sel_986632 = array_index_986479 == array_index_948715 ? add_986631 : sel_986628;
  assign add_986635 = sel_986632 + 8'h01;
  assign sel_986636 = array_index_986479 == array_index_948721 ? add_986635 : sel_986632;
  assign add_986639 = sel_986636 + 8'h01;
  assign sel_986640 = array_index_986479 == array_index_948727 ? add_986639 : sel_986636;
  assign add_986643 = sel_986640 + 8'h01;
  assign sel_986644 = array_index_986479 == array_index_948733 ? add_986643 : sel_986640;
  assign add_986647 = sel_986644 + 8'h01;
  assign sel_986648 = array_index_986479 == array_index_948739 ? add_986647 : sel_986644;
  assign add_986651 = sel_986648 + 8'h01;
  assign sel_986652 = array_index_986479 == array_index_948745 ? add_986651 : sel_986648;
  assign add_986655 = sel_986652 + 8'h01;
  assign sel_986656 = array_index_986479 == array_index_948751 ? add_986655 : sel_986652;
  assign add_986659 = sel_986656 + 8'h01;
  assign sel_986660 = array_index_986479 == array_index_948757 ? add_986659 : sel_986656;
  assign add_986663 = sel_986660 + 8'h01;
  assign sel_986664 = array_index_986479 == array_index_948763 ? add_986663 : sel_986660;
  assign add_986667 = sel_986664 + 8'h01;
  assign sel_986668 = array_index_986479 == array_index_948769 ? add_986667 : sel_986664;
  assign add_986671 = sel_986668 + 8'h01;
  assign sel_986672 = array_index_986479 == array_index_948775 ? add_986671 : sel_986668;
  assign add_986675 = sel_986672 + 8'h01;
  assign sel_986676 = array_index_986479 == array_index_948781 ? add_986675 : sel_986672;
  assign add_986679 = sel_986676 + 8'h01;
  assign sel_986680 = array_index_986479 == array_index_948787 ? add_986679 : sel_986676;
  assign add_986683 = sel_986680 + 8'h01;
  assign sel_986684 = array_index_986479 == array_index_948793 ? add_986683 : sel_986680;
  assign add_986687 = sel_986684 + 8'h01;
  assign sel_986688 = array_index_986479 == array_index_948799 ? add_986687 : sel_986684;
  assign add_986691 = sel_986688 + 8'h01;
  assign sel_986692 = array_index_986479 == array_index_948805 ? add_986691 : sel_986688;
  assign add_986695 = sel_986692 + 8'h01;
  assign sel_986696 = array_index_986479 == array_index_948811 ? add_986695 : sel_986692;
  assign add_986699 = sel_986696 + 8'h01;
  assign sel_986700 = array_index_986479 == array_index_948817 ? add_986699 : sel_986696;
  assign add_986703 = sel_986700 + 8'h01;
  assign sel_986704 = array_index_986479 == array_index_948823 ? add_986703 : sel_986700;
  assign add_986707 = sel_986704 + 8'h01;
  assign sel_986708 = array_index_986479 == array_index_948829 ? add_986707 : sel_986704;
  assign add_986711 = sel_986708 + 8'h01;
  assign sel_986712 = array_index_986479 == array_index_948835 ? add_986711 : sel_986708;
  assign add_986715 = sel_986712 + 8'h01;
  assign sel_986716 = array_index_986479 == array_index_948841 ? add_986715 : sel_986712;
  assign add_986719 = sel_986716 + 8'h01;
  assign sel_986720 = array_index_986479 == array_index_948847 ? add_986719 : sel_986716;
  assign add_986723 = sel_986720 + 8'h01;
  assign sel_986724 = array_index_986479 == array_index_948853 ? add_986723 : sel_986720;
  assign add_986727 = sel_986724 + 8'h01;
  assign sel_986728 = array_index_986479 == array_index_948859 ? add_986727 : sel_986724;
  assign add_986731 = sel_986728 + 8'h01;
  assign sel_986732 = array_index_986479 == array_index_948865 ? add_986731 : sel_986728;
  assign add_986735 = sel_986732 + 8'h01;
  assign sel_986736 = array_index_986479 == array_index_948871 ? add_986735 : sel_986732;
  assign add_986739 = sel_986736 + 8'h01;
  assign sel_986740 = array_index_986479 == array_index_948877 ? add_986739 : sel_986736;
  assign add_986743 = sel_986740 + 8'h01;
  assign sel_986744 = array_index_986479 == array_index_948883 ? add_986743 : sel_986740;
  assign add_986747 = sel_986744 + 8'h01;
  assign sel_986748 = array_index_986479 == array_index_948889 ? add_986747 : sel_986744;
  assign add_986751 = sel_986748 + 8'h01;
  assign sel_986752 = array_index_986479 == array_index_948895 ? add_986751 : sel_986748;
  assign add_986755 = sel_986752 + 8'h01;
  assign sel_986756 = array_index_986479 == array_index_948901 ? add_986755 : sel_986752;
  assign add_986759 = sel_986756 + 8'h01;
  assign sel_986760 = array_index_986479 == array_index_948907 ? add_986759 : sel_986756;
  assign add_986763 = sel_986760 + 8'h01;
  assign sel_986764 = array_index_986479 == array_index_948913 ? add_986763 : sel_986760;
  assign add_986767 = sel_986764 + 8'h01;
  assign sel_986768 = array_index_986479 == array_index_948919 ? add_986767 : sel_986764;
  assign add_986771 = sel_986768 + 8'h01;
  assign sel_986772 = array_index_986479 == array_index_948925 ? add_986771 : sel_986768;
  assign add_986775 = sel_986772 + 8'h01;
  assign sel_986776 = array_index_986479 == array_index_948931 ? add_986775 : sel_986772;
  assign add_986779 = sel_986776 + 8'h01;
  assign sel_986780 = array_index_986479 == array_index_948937 ? add_986779 : sel_986776;
  assign add_986783 = sel_986780 + 8'h01;
  assign sel_986784 = array_index_986479 == array_index_948943 ? add_986783 : sel_986780;
  assign add_986787 = sel_986784 + 8'h01;
  assign sel_986788 = array_index_986479 == array_index_948949 ? add_986787 : sel_986784;
  assign add_986791 = sel_986788 + 8'h01;
  assign sel_986792 = array_index_986479 == array_index_948955 ? add_986791 : sel_986788;
  assign add_986795 = sel_986792 + 8'h01;
  assign sel_986796 = array_index_986479 == array_index_948961 ? add_986795 : sel_986792;
  assign add_986799 = sel_986796 + 8'h01;
  assign sel_986800 = array_index_986479 == array_index_948967 ? add_986799 : sel_986796;
  assign add_986803 = sel_986800 + 8'h01;
  assign sel_986804 = array_index_986479 == array_index_948973 ? add_986803 : sel_986800;
  assign add_986807 = sel_986804 + 8'h01;
  assign sel_986808 = array_index_986479 == array_index_948979 ? add_986807 : sel_986804;
  assign add_986811 = sel_986808 + 8'h01;
  assign sel_986812 = array_index_986479 == array_index_948985 ? add_986811 : sel_986808;
  assign add_986815 = sel_986812 + 8'h01;
  assign sel_986816 = array_index_986479 == array_index_948991 ? add_986815 : sel_986812;
  assign add_986819 = sel_986816 + 8'h01;
  assign sel_986820 = array_index_986479 == array_index_948997 ? add_986819 : sel_986816;
  assign add_986823 = sel_986820 + 8'h01;
  assign sel_986824 = array_index_986479 == array_index_949003 ? add_986823 : sel_986820;
  assign add_986827 = sel_986824 + 8'h01;
  assign sel_986828 = array_index_986479 == array_index_949009 ? add_986827 : sel_986824;
  assign add_986831 = sel_986828 + 8'h01;
  assign sel_986832 = array_index_986479 == array_index_949015 ? add_986831 : sel_986828;
  assign add_986835 = sel_986832 + 8'h01;
  assign sel_986836 = array_index_986479 == array_index_949021 ? add_986835 : sel_986832;
  assign add_986839 = sel_986836 + 8'h01;
  assign sel_986840 = array_index_986479 == array_index_949027 ? add_986839 : sel_986836;
  assign add_986843 = sel_986840 + 8'h01;
  assign sel_986844 = array_index_986479 == array_index_949033 ? add_986843 : sel_986840;
  assign add_986847 = sel_986844 + 8'h01;
  assign sel_986848 = array_index_986479 == array_index_949039 ? add_986847 : sel_986844;
  assign add_986851 = sel_986848 + 8'h01;
  assign sel_986852 = array_index_986479 == array_index_949045 ? add_986851 : sel_986848;
  assign add_986855 = sel_986852 + 8'h01;
  assign sel_986856 = array_index_986479 == array_index_949051 ? add_986855 : sel_986852;
  assign add_986859 = sel_986856 + 8'h01;
  assign sel_986860 = array_index_986479 == array_index_949057 ? add_986859 : sel_986856;
  assign add_986863 = sel_986860 + 8'h01;
  assign sel_986864 = array_index_986479 == array_index_949063 ? add_986863 : sel_986860;
  assign add_986867 = sel_986864 + 8'h01;
  assign sel_986868 = array_index_986479 == array_index_949069 ? add_986867 : sel_986864;
  assign add_986871 = sel_986868 + 8'h01;
  assign sel_986872 = array_index_986479 == array_index_949075 ? add_986871 : sel_986868;
  assign add_986875 = sel_986872 + 8'h01;
  assign sel_986876 = array_index_986479 == array_index_949081 ? add_986875 : sel_986872;
  assign add_986880 = sel_986876 + 8'h01;
  assign array_index_986881 = set1_unflattened[7'h5f];
  assign sel_986882 = array_index_986479 == array_index_949087 ? add_986880 : sel_986876;
  assign add_986885 = sel_986882 + 8'h01;
  assign sel_986886 = array_index_986881 == array_index_948483 ? add_986885 : sel_986882;
  assign add_986889 = sel_986886 + 8'h01;
  assign sel_986890 = array_index_986881 == array_index_948487 ? add_986889 : sel_986886;
  assign add_986893 = sel_986890 + 8'h01;
  assign sel_986894 = array_index_986881 == array_index_948495 ? add_986893 : sel_986890;
  assign add_986897 = sel_986894 + 8'h01;
  assign sel_986898 = array_index_986881 == array_index_948503 ? add_986897 : sel_986894;
  assign add_986901 = sel_986898 + 8'h01;
  assign sel_986902 = array_index_986881 == array_index_948511 ? add_986901 : sel_986898;
  assign add_986905 = sel_986902 + 8'h01;
  assign sel_986906 = array_index_986881 == array_index_948519 ? add_986905 : sel_986902;
  assign add_986909 = sel_986906 + 8'h01;
  assign sel_986910 = array_index_986881 == array_index_948527 ? add_986909 : sel_986906;
  assign add_986913 = sel_986910 + 8'h01;
  assign sel_986914 = array_index_986881 == array_index_948535 ? add_986913 : sel_986910;
  assign add_986917 = sel_986914 + 8'h01;
  assign sel_986918 = array_index_986881 == array_index_948541 ? add_986917 : sel_986914;
  assign add_986921 = sel_986918 + 8'h01;
  assign sel_986922 = array_index_986881 == array_index_948547 ? add_986921 : sel_986918;
  assign add_986925 = sel_986922 + 8'h01;
  assign sel_986926 = array_index_986881 == array_index_948553 ? add_986925 : sel_986922;
  assign add_986929 = sel_986926 + 8'h01;
  assign sel_986930 = array_index_986881 == array_index_948559 ? add_986929 : sel_986926;
  assign add_986933 = sel_986930 + 8'h01;
  assign sel_986934 = array_index_986881 == array_index_948565 ? add_986933 : sel_986930;
  assign add_986937 = sel_986934 + 8'h01;
  assign sel_986938 = array_index_986881 == array_index_948571 ? add_986937 : sel_986934;
  assign add_986941 = sel_986938 + 8'h01;
  assign sel_986942 = array_index_986881 == array_index_948577 ? add_986941 : sel_986938;
  assign add_986945 = sel_986942 + 8'h01;
  assign sel_986946 = array_index_986881 == array_index_948583 ? add_986945 : sel_986942;
  assign add_986949 = sel_986946 + 8'h01;
  assign sel_986950 = array_index_986881 == array_index_948589 ? add_986949 : sel_986946;
  assign add_986953 = sel_986950 + 8'h01;
  assign sel_986954 = array_index_986881 == array_index_948595 ? add_986953 : sel_986950;
  assign add_986957 = sel_986954 + 8'h01;
  assign sel_986958 = array_index_986881 == array_index_948601 ? add_986957 : sel_986954;
  assign add_986961 = sel_986958 + 8'h01;
  assign sel_986962 = array_index_986881 == array_index_948607 ? add_986961 : sel_986958;
  assign add_986965 = sel_986962 + 8'h01;
  assign sel_986966 = array_index_986881 == array_index_948613 ? add_986965 : sel_986962;
  assign add_986969 = sel_986966 + 8'h01;
  assign sel_986970 = array_index_986881 == array_index_948619 ? add_986969 : sel_986966;
  assign add_986973 = sel_986970 + 8'h01;
  assign sel_986974 = array_index_986881 == array_index_948625 ? add_986973 : sel_986970;
  assign add_986977 = sel_986974 + 8'h01;
  assign sel_986978 = array_index_986881 == array_index_948631 ? add_986977 : sel_986974;
  assign add_986981 = sel_986978 + 8'h01;
  assign sel_986982 = array_index_986881 == array_index_948637 ? add_986981 : sel_986978;
  assign add_986985 = sel_986982 + 8'h01;
  assign sel_986986 = array_index_986881 == array_index_948643 ? add_986985 : sel_986982;
  assign add_986989 = sel_986986 + 8'h01;
  assign sel_986990 = array_index_986881 == array_index_948649 ? add_986989 : sel_986986;
  assign add_986993 = sel_986990 + 8'h01;
  assign sel_986994 = array_index_986881 == array_index_948655 ? add_986993 : sel_986990;
  assign add_986997 = sel_986994 + 8'h01;
  assign sel_986998 = array_index_986881 == array_index_948661 ? add_986997 : sel_986994;
  assign add_987001 = sel_986998 + 8'h01;
  assign sel_987002 = array_index_986881 == array_index_948667 ? add_987001 : sel_986998;
  assign add_987005 = sel_987002 + 8'h01;
  assign sel_987006 = array_index_986881 == array_index_948673 ? add_987005 : sel_987002;
  assign add_987009 = sel_987006 + 8'h01;
  assign sel_987010 = array_index_986881 == array_index_948679 ? add_987009 : sel_987006;
  assign add_987013 = sel_987010 + 8'h01;
  assign sel_987014 = array_index_986881 == array_index_948685 ? add_987013 : sel_987010;
  assign add_987017 = sel_987014 + 8'h01;
  assign sel_987018 = array_index_986881 == array_index_948691 ? add_987017 : sel_987014;
  assign add_987021 = sel_987018 + 8'h01;
  assign sel_987022 = array_index_986881 == array_index_948697 ? add_987021 : sel_987018;
  assign add_987025 = sel_987022 + 8'h01;
  assign sel_987026 = array_index_986881 == array_index_948703 ? add_987025 : sel_987022;
  assign add_987029 = sel_987026 + 8'h01;
  assign sel_987030 = array_index_986881 == array_index_948709 ? add_987029 : sel_987026;
  assign add_987033 = sel_987030 + 8'h01;
  assign sel_987034 = array_index_986881 == array_index_948715 ? add_987033 : sel_987030;
  assign add_987037 = sel_987034 + 8'h01;
  assign sel_987038 = array_index_986881 == array_index_948721 ? add_987037 : sel_987034;
  assign add_987041 = sel_987038 + 8'h01;
  assign sel_987042 = array_index_986881 == array_index_948727 ? add_987041 : sel_987038;
  assign add_987045 = sel_987042 + 8'h01;
  assign sel_987046 = array_index_986881 == array_index_948733 ? add_987045 : sel_987042;
  assign add_987049 = sel_987046 + 8'h01;
  assign sel_987050 = array_index_986881 == array_index_948739 ? add_987049 : sel_987046;
  assign add_987053 = sel_987050 + 8'h01;
  assign sel_987054 = array_index_986881 == array_index_948745 ? add_987053 : sel_987050;
  assign add_987057 = sel_987054 + 8'h01;
  assign sel_987058 = array_index_986881 == array_index_948751 ? add_987057 : sel_987054;
  assign add_987061 = sel_987058 + 8'h01;
  assign sel_987062 = array_index_986881 == array_index_948757 ? add_987061 : sel_987058;
  assign add_987065 = sel_987062 + 8'h01;
  assign sel_987066 = array_index_986881 == array_index_948763 ? add_987065 : sel_987062;
  assign add_987069 = sel_987066 + 8'h01;
  assign sel_987070 = array_index_986881 == array_index_948769 ? add_987069 : sel_987066;
  assign add_987073 = sel_987070 + 8'h01;
  assign sel_987074 = array_index_986881 == array_index_948775 ? add_987073 : sel_987070;
  assign add_987077 = sel_987074 + 8'h01;
  assign sel_987078 = array_index_986881 == array_index_948781 ? add_987077 : sel_987074;
  assign add_987081 = sel_987078 + 8'h01;
  assign sel_987082 = array_index_986881 == array_index_948787 ? add_987081 : sel_987078;
  assign add_987085 = sel_987082 + 8'h01;
  assign sel_987086 = array_index_986881 == array_index_948793 ? add_987085 : sel_987082;
  assign add_987089 = sel_987086 + 8'h01;
  assign sel_987090 = array_index_986881 == array_index_948799 ? add_987089 : sel_987086;
  assign add_987093 = sel_987090 + 8'h01;
  assign sel_987094 = array_index_986881 == array_index_948805 ? add_987093 : sel_987090;
  assign add_987097 = sel_987094 + 8'h01;
  assign sel_987098 = array_index_986881 == array_index_948811 ? add_987097 : sel_987094;
  assign add_987101 = sel_987098 + 8'h01;
  assign sel_987102 = array_index_986881 == array_index_948817 ? add_987101 : sel_987098;
  assign add_987105 = sel_987102 + 8'h01;
  assign sel_987106 = array_index_986881 == array_index_948823 ? add_987105 : sel_987102;
  assign add_987109 = sel_987106 + 8'h01;
  assign sel_987110 = array_index_986881 == array_index_948829 ? add_987109 : sel_987106;
  assign add_987113 = sel_987110 + 8'h01;
  assign sel_987114 = array_index_986881 == array_index_948835 ? add_987113 : sel_987110;
  assign add_987117 = sel_987114 + 8'h01;
  assign sel_987118 = array_index_986881 == array_index_948841 ? add_987117 : sel_987114;
  assign add_987121 = sel_987118 + 8'h01;
  assign sel_987122 = array_index_986881 == array_index_948847 ? add_987121 : sel_987118;
  assign add_987125 = sel_987122 + 8'h01;
  assign sel_987126 = array_index_986881 == array_index_948853 ? add_987125 : sel_987122;
  assign add_987129 = sel_987126 + 8'h01;
  assign sel_987130 = array_index_986881 == array_index_948859 ? add_987129 : sel_987126;
  assign add_987133 = sel_987130 + 8'h01;
  assign sel_987134 = array_index_986881 == array_index_948865 ? add_987133 : sel_987130;
  assign add_987137 = sel_987134 + 8'h01;
  assign sel_987138 = array_index_986881 == array_index_948871 ? add_987137 : sel_987134;
  assign add_987141 = sel_987138 + 8'h01;
  assign sel_987142 = array_index_986881 == array_index_948877 ? add_987141 : sel_987138;
  assign add_987145 = sel_987142 + 8'h01;
  assign sel_987146 = array_index_986881 == array_index_948883 ? add_987145 : sel_987142;
  assign add_987149 = sel_987146 + 8'h01;
  assign sel_987150 = array_index_986881 == array_index_948889 ? add_987149 : sel_987146;
  assign add_987153 = sel_987150 + 8'h01;
  assign sel_987154 = array_index_986881 == array_index_948895 ? add_987153 : sel_987150;
  assign add_987157 = sel_987154 + 8'h01;
  assign sel_987158 = array_index_986881 == array_index_948901 ? add_987157 : sel_987154;
  assign add_987161 = sel_987158 + 8'h01;
  assign sel_987162 = array_index_986881 == array_index_948907 ? add_987161 : sel_987158;
  assign add_987165 = sel_987162 + 8'h01;
  assign sel_987166 = array_index_986881 == array_index_948913 ? add_987165 : sel_987162;
  assign add_987169 = sel_987166 + 8'h01;
  assign sel_987170 = array_index_986881 == array_index_948919 ? add_987169 : sel_987166;
  assign add_987173 = sel_987170 + 8'h01;
  assign sel_987174 = array_index_986881 == array_index_948925 ? add_987173 : sel_987170;
  assign add_987177 = sel_987174 + 8'h01;
  assign sel_987178 = array_index_986881 == array_index_948931 ? add_987177 : sel_987174;
  assign add_987181 = sel_987178 + 8'h01;
  assign sel_987182 = array_index_986881 == array_index_948937 ? add_987181 : sel_987178;
  assign add_987185 = sel_987182 + 8'h01;
  assign sel_987186 = array_index_986881 == array_index_948943 ? add_987185 : sel_987182;
  assign add_987189 = sel_987186 + 8'h01;
  assign sel_987190 = array_index_986881 == array_index_948949 ? add_987189 : sel_987186;
  assign add_987193 = sel_987190 + 8'h01;
  assign sel_987194 = array_index_986881 == array_index_948955 ? add_987193 : sel_987190;
  assign add_987197 = sel_987194 + 8'h01;
  assign sel_987198 = array_index_986881 == array_index_948961 ? add_987197 : sel_987194;
  assign add_987201 = sel_987198 + 8'h01;
  assign sel_987202 = array_index_986881 == array_index_948967 ? add_987201 : sel_987198;
  assign add_987205 = sel_987202 + 8'h01;
  assign sel_987206 = array_index_986881 == array_index_948973 ? add_987205 : sel_987202;
  assign add_987209 = sel_987206 + 8'h01;
  assign sel_987210 = array_index_986881 == array_index_948979 ? add_987209 : sel_987206;
  assign add_987213 = sel_987210 + 8'h01;
  assign sel_987214 = array_index_986881 == array_index_948985 ? add_987213 : sel_987210;
  assign add_987217 = sel_987214 + 8'h01;
  assign sel_987218 = array_index_986881 == array_index_948991 ? add_987217 : sel_987214;
  assign add_987221 = sel_987218 + 8'h01;
  assign sel_987222 = array_index_986881 == array_index_948997 ? add_987221 : sel_987218;
  assign add_987225 = sel_987222 + 8'h01;
  assign sel_987226 = array_index_986881 == array_index_949003 ? add_987225 : sel_987222;
  assign add_987229 = sel_987226 + 8'h01;
  assign sel_987230 = array_index_986881 == array_index_949009 ? add_987229 : sel_987226;
  assign add_987233 = sel_987230 + 8'h01;
  assign sel_987234 = array_index_986881 == array_index_949015 ? add_987233 : sel_987230;
  assign add_987237 = sel_987234 + 8'h01;
  assign sel_987238 = array_index_986881 == array_index_949021 ? add_987237 : sel_987234;
  assign add_987241 = sel_987238 + 8'h01;
  assign sel_987242 = array_index_986881 == array_index_949027 ? add_987241 : sel_987238;
  assign add_987245 = sel_987242 + 8'h01;
  assign sel_987246 = array_index_986881 == array_index_949033 ? add_987245 : sel_987242;
  assign add_987249 = sel_987246 + 8'h01;
  assign sel_987250 = array_index_986881 == array_index_949039 ? add_987249 : sel_987246;
  assign add_987253 = sel_987250 + 8'h01;
  assign sel_987254 = array_index_986881 == array_index_949045 ? add_987253 : sel_987250;
  assign add_987257 = sel_987254 + 8'h01;
  assign sel_987258 = array_index_986881 == array_index_949051 ? add_987257 : sel_987254;
  assign add_987261 = sel_987258 + 8'h01;
  assign sel_987262 = array_index_986881 == array_index_949057 ? add_987261 : sel_987258;
  assign add_987265 = sel_987262 + 8'h01;
  assign sel_987266 = array_index_986881 == array_index_949063 ? add_987265 : sel_987262;
  assign add_987269 = sel_987266 + 8'h01;
  assign sel_987270 = array_index_986881 == array_index_949069 ? add_987269 : sel_987266;
  assign add_987273 = sel_987270 + 8'h01;
  assign sel_987274 = array_index_986881 == array_index_949075 ? add_987273 : sel_987270;
  assign add_987277 = sel_987274 + 8'h01;
  assign sel_987278 = array_index_986881 == array_index_949081 ? add_987277 : sel_987274;
  assign add_987282 = sel_987278 + 8'h01;
  assign array_index_987283 = set1_unflattened[7'h60];
  assign sel_987284 = array_index_986881 == array_index_949087 ? add_987282 : sel_987278;
  assign add_987287 = sel_987284 + 8'h01;
  assign sel_987288 = array_index_987283 == array_index_948483 ? add_987287 : sel_987284;
  assign add_987291 = sel_987288 + 8'h01;
  assign sel_987292 = array_index_987283 == array_index_948487 ? add_987291 : sel_987288;
  assign add_987295 = sel_987292 + 8'h01;
  assign sel_987296 = array_index_987283 == array_index_948495 ? add_987295 : sel_987292;
  assign add_987299 = sel_987296 + 8'h01;
  assign sel_987300 = array_index_987283 == array_index_948503 ? add_987299 : sel_987296;
  assign add_987303 = sel_987300 + 8'h01;
  assign sel_987304 = array_index_987283 == array_index_948511 ? add_987303 : sel_987300;
  assign add_987307 = sel_987304 + 8'h01;
  assign sel_987308 = array_index_987283 == array_index_948519 ? add_987307 : sel_987304;
  assign add_987311 = sel_987308 + 8'h01;
  assign sel_987312 = array_index_987283 == array_index_948527 ? add_987311 : sel_987308;
  assign add_987315 = sel_987312 + 8'h01;
  assign sel_987316 = array_index_987283 == array_index_948535 ? add_987315 : sel_987312;
  assign add_987319 = sel_987316 + 8'h01;
  assign sel_987320 = array_index_987283 == array_index_948541 ? add_987319 : sel_987316;
  assign add_987323 = sel_987320 + 8'h01;
  assign sel_987324 = array_index_987283 == array_index_948547 ? add_987323 : sel_987320;
  assign add_987327 = sel_987324 + 8'h01;
  assign sel_987328 = array_index_987283 == array_index_948553 ? add_987327 : sel_987324;
  assign add_987331 = sel_987328 + 8'h01;
  assign sel_987332 = array_index_987283 == array_index_948559 ? add_987331 : sel_987328;
  assign add_987335 = sel_987332 + 8'h01;
  assign sel_987336 = array_index_987283 == array_index_948565 ? add_987335 : sel_987332;
  assign add_987339 = sel_987336 + 8'h01;
  assign sel_987340 = array_index_987283 == array_index_948571 ? add_987339 : sel_987336;
  assign add_987343 = sel_987340 + 8'h01;
  assign sel_987344 = array_index_987283 == array_index_948577 ? add_987343 : sel_987340;
  assign add_987347 = sel_987344 + 8'h01;
  assign sel_987348 = array_index_987283 == array_index_948583 ? add_987347 : sel_987344;
  assign add_987351 = sel_987348 + 8'h01;
  assign sel_987352 = array_index_987283 == array_index_948589 ? add_987351 : sel_987348;
  assign add_987355 = sel_987352 + 8'h01;
  assign sel_987356 = array_index_987283 == array_index_948595 ? add_987355 : sel_987352;
  assign add_987359 = sel_987356 + 8'h01;
  assign sel_987360 = array_index_987283 == array_index_948601 ? add_987359 : sel_987356;
  assign add_987363 = sel_987360 + 8'h01;
  assign sel_987364 = array_index_987283 == array_index_948607 ? add_987363 : sel_987360;
  assign add_987367 = sel_987364 + 8'h01;
  assign sel_987368 = array_index_987283 == array_index_948613 ? add_987367 : sel_987364;
  assign add_987371 = sel_987368 + 8'h01;
  assign sel_987372 = array_index_987283 == array_index_948619 ? add_987371 : sel_987368;
  assign add_987375 = sel_987372 + 8'h01;
  assign sel_987376 = array_index_987283 == array_index_948625 ? add_987375 : sel_987372;
  assign add_987379 = sel_987376 + 8'h01;
  assign sel_987380 = array_index_987283 == array_index_948631 ? add_987379 : sel_987376;
  assign add_987383 = sel_987380 + 8'h01;
  assign sel_987384 = array_index_987283 == array_index_948637 ? add_987383 : sel_987380;
  assign add_987387 = sel_987384 + 8'h01;
  assign sel_987388 = array_index_987283 == array_index_948643 ? add_987387 : sel_987384;
  assign add_987391 = sel_987388 + 8'h01;
  assign sel_987392 = array_index_987283 == array_index_948649 ? add_987391 : sel_987388;
  assign add_987395 = sel_987392 + 8'h01;
  assign sel_987396 = array_index_987283 == array_index_948655 ? add_987395 : sel_987392;
  assign add_987399 = sel_987396 + 8'h01;
  assign sel_987400 = array_index_987283 == array_index_948661 ? add_987399 : sel_987396;
  assign add_987403 = sel_987400 + 8'h01;
  assign sel_987404 = array_index_987283 == array_index_948667 ? add_987403 : sel_987400;
  assign add_987407 = sel_987404 + 8'h01;
  assign sel_987408 = array_index_987283 == array_index_948673 ? add_987407 : sel_987404;
  assign add_987411 = sel_987408 + 8'h01;
  assign sel_987412 = array_index_987283 == array_index_948679 ? add_987411 : sel_987408;
  assign add_987415 = sel_987412 + 8'h01;
  assign sel_987416 = array_index_987283 == array_index_948685 ? add_987415 : sel_987412;
  assign add_987419 = sel_987416 + 8'h01;
  assign sel_987420 = array_index_987283 == array_index_948691 ? add_987419 : sel_987416;
  assign add_987423 = sel_987420 + 8'h01;
  assign sel_987424 = array_index_987283 == array_index_948697 ? add_987423 : sel_987420;
  assign add_987427 = sel_987424 + 8'h01;
  assign sel_987428 = array_index_987283 == array_index_948703 ? add_987427 : sel_987424;
  assign add_987431 = sel_987428 + 8'h01;
  assign sel_987432 = array_index_987283 == array_index_948709 ? add_987431 : sel_987428;
  assign add_987435 = sel_987432 + 8'h01;
  assign sel_987436 = array_index_987283 == array_index_948715 ? add_987435 : sel_987432;
  assign add_987439 = sel_987436 + 8'h01;
  assign sel_987440 = array_index_987283 == array_index_948721 ? add_987439 : sel_987436;
  assign add_987443 = sel_987440 + 8'h01;
  assign sel_987444 = array_index_987283 == array_index_948727 ? add_987443 : sel_987440;
  assign add_987447 = sel_987444 + 8'h01;
  assign sel_987448 = array_index_987283 == array_index_948733 ? add_987447 : sel_987444;
  assign add_987451 = sel_987448 + 8'h01;
  assign sel_987452 = array_index_987283 == array_index_948739 ? add_987451 : sel_987448;
  assign add_987455 = sel_987452 + 8'h01;
  assign sel_987456 = array_index_987283 == array_index_948745 ? add_987455 : sel_987452;
  assign add_987459 = sel_987456 + 8'h01;
  assign sel_987460 = array_index_987283 == array_index_948751 ? add_987459 : sel_987456;
  assign add_987463 = sel_987460 + 8'h01;
  assign sel_987464 = array_index_987283 == array_index_948757 ? add_987463 : sel_987460;
  assign add_987467 = sel_987464 + 8'h01;
  assign sel_987468 = array_index_987283 == array_index_948763 ? add_987467 : sel_987464;
  assign add_987471 = sel_987468 + 8'h01;
  assign sel_987472 = array_index_987283 == array_index_948769 ? add_987471 : sel_987468;
  assign add_987475 = sel_987472 + 8'h01;
  assign sel_987476 = array_index_987283 == array_index_948775 ? add_987475 : sel_987472;
  assign add_987479 = sel_987476 + 8'h01;
  assign sel_987480 = array_index_987283 == array_index_948781 ? add_987479 : sel_987476;
  assign add_987483 = sel_987480 + 8'h01;
  assign sel_987484 = array_index_987283 == array_index_948787 ? add_987483 : sel_987480;
  assign add_987487 = sel_987484 + 8'h01;
  assign sel_987488 = array_index_987283 == array_index_948793 ? add_987487 : sel_987484;
  assign add_987491 = sel_987488 + 8'h01;
  assign sel_987492 = array_index_987283 == array_index_948799 ? add_987491 : sel_987488;
  assign add_987495 = sel_987492 + 8'h01;
  assign sel_987496 = array_index_987283 == array_index_948805 ? add_987495 : sel_987492;
  assign add_987499 = sel_987496 + 8'h01;
  assign sel_987500 = array_index_987283 == array_index_948811 ? add_987499 : sel_987496;
  assign add_987503 = sel_987500 + 8'h01;
  assign sel_987504 = array_index_987283 == array_index_948817 ? add_987503 : sel_987500;
  assign add_987507 = sel_987504 + 8'h01;
  assign sel_987508 = array_index_987283 == array_index_948823 ? add_987507 : sel_987504;
  assign add_987511 = sel_987508 + 8'h01;
  assign sel_987512 = array_index_987283 == array_index_948829 ? add_987511 : sel_987508;
  assign add_987515 = sel_987512 + 8'h01;
  assign sel_987516 = array_index_987283 == array_index_948835 ? add_987515 : sel_987512;
  assign add_987519 = sel_987516 + 8'h01;
  assign sel_987520 = array_index_987283 == array_index_948841 ? add_987519 : sel_987516;
  assign add_987523 = sel_987520 + 8'h01;
  assign sel_987524 = array_index_987283 == array_index_948847 ? add_987523 : sel_987520;
  assign add_987527 = sel_987524 + 8'h01;
  assign sel_987528 = array_index_987283 == array_index_948853 ? add_987527 : sel_987524;
  assign add_987531 = sel_987528 + 8'h01;
  assign sel_987532 = array_index_987283 == array_index_948859 ? add_987531 : sel_987528;
  assign add_987535 = sel_987532 + 8'h01;
  assign sel_987536 = array_index_987283 == array_index_948865 ? add_987535 : sel_987532;
  assign add_987539 = sel_987536 + 8'h01;
  assign sel_987540 = array_index_987283 == array_index_948871 ? add_987539 : sel_987536;
  assign add_987543 = sel_987540 + 8'h01;
  assign sel_987544 = array_index_987283 == array_index_948877 ? add_987543 : sel_987540;
  assign add_987547 = sel_987544 + 8'h01;
  assign sel_987548 = array_index_987283 == array_index_948883 ? add_987547 : sel_987544;
  assign add_987551 = sel_987548 + 8'h01;
  assign sel_987552 = array_index_987283 == array_index_948889 ? add_987551 : sel_987548;
  assign add_987555 = sel_987552 + 8'h01;
  assign sel_987556 = array_index_987283 == array_index_948895 ? add_987555 : sel_987552;
  assign add_987559 = sel_987556 + 8'h01;
  assign sel_987560 = array_index_987283 == array_index_948901 ? add_987559 : sel_987556;
  assign add_987563 = sel_987560 + 8'h01;
  assign sel_987564 = array_index_987283 == array_index_948907 ? add_987563 : sel_987560;
  assign add_987567 = sel_987564 + 8'h01;
  assign sel_987568 = array_index_987283 == array_index_948913 ? add_987567 : sel_987564;
  assign add_987571 = sel_987568 + 8'h01;
  assign sel_987572 = array_index_987283 == array_index_948919 ? add_987571 : sel_987568;
  assign add_987575 = sel_987572 + 8'h01;
  assign sel_987576 = array_index_987283 == array_index_948925 ? add_987575 : sel_987572;
  assign add_987579 = sel_987576 + 8'h01;
  assign sel_987580 = array_index_987283 == array_index_948931 ? add_987579 : sel_987576;
  assign add_987583 = sel_987580 + 8'h01;
  assign sel_987584 = array_index_987283 == array_index_948937 ? add_987583 : sel_987580;
  assign add_987587 = sel_987584 + 8'h01;
  assign sel_987588 = array_index_987283 == array_index_948943 ? add_987587 : sel_987584;
  assign add_987591 = sel_987588 + 8'h01;
  assign sel_987592 = array_index_987283 == array_index_948949 ? add_987591 : sel_987588;
  assign add_987595 = sel_987592 + 8'h01;
  assign sel_987596 = array_index_987283 == array_index_948955 ? add_987595 : sel_987592;
  assign add_987599 = sel_987596 + 8'h01;
  assign sel_987600 = array_index_987283 == array_index_948961 ? add_987599 : sel_987596;
  assign add_987603 = sel_987600 + 8'h01;
  assign sel_987604 = array_index_987283 == array_index_948967 ? add_987603 : sel_987600;
  assign add_987607 = sel_987604 + 8'h01;
  assign sel_987608 = array_index_987283 == array_index_948973 ? add_987607 : sel_987604;
  assign add_987611 = sel_987608 + 8'h01;
  assign sel_987612 = array_index_987283 == array_index_948979 ? add_987611 : sel_987608;
  assign add_987615 = sel_987612 + 8'h01;
  assign sel_987616 = array_index_987283 == array_index_948985 ? add_987615 : sel_987612;
  assign add_987619 = sel_987616 + 8'h01;
  assign sel_987620 = array_index_987283 == array_index_948991 ? add_987619 : sel_987616;
  assign add_987623 = sel_987620 + 8'h01;
  assign sel_987624 = array_index_987283 == array_index_948997 ? add_987623 : sel_987620;
  assign add_987627 = sel_987624 + 8'h01;
  assign sel_987628 = array_index_987283 == array_index_949003 ? add_987627 : sel_987624;
  assign add_987631 = sel_987628 + 8'h01;
  assign sel_987632 = array_index_987283 == array_index_949009 ? add_987631 : sel_987628;
  assign add_987635 = sel_987632 + 8'h01;
  assign sel_987636 = array_index_987283 == array_index_949015 ? add_987635 : sel_987632;
  assign add_987639 = sel_987636 + 8'h01;
  assign sel_987640 = array_index_987283 == array_index_949021 ? add_987639 : sel_987636;
  assign add_987643 = sel_987640 + 8'h01;
  assign sel_987644 = array_index_987283 == array_index_949027 ? add_987643 : sel_987640;
  assign add_987647 = sel_987644 + 8'h01;
  assign sel_987648 = array_index_987283 == array_index_949033 ? add_987647 : sel_987644;
  assign add_987651 = sel_987648 + 8'h01;
  assign sel_987652 = array_index_987283 == array_index_949039 ? add_987651 : sel_987648;
  assign add_987655 = sel_987652 + 8'h01;
  assign sel_987656 = array_index_987283 == array_index_949045 ? add_987655 : sel_987652;
  assign add_987659 = sel_987656 + 8'h01;
  assign sel_987660 = array_index_987283 == array_index_949051 ? add_987659 : sel_987656;
  assign add_987663 = sel_987660 + 8'h01;
  assign sel_987664 = array_index_987283 == array_index_949057 ? add_987663 : sel_987660;
  assign add_987667 = sel_987664 + 8'h01;
  assign sel_987668 = array_index_987283 == array_index_949063 ? add_987667 : sel_987664;
  assign add_987671 = sel_987668 + 8'h01;
  assign sel_987672 = array_index_987283 == array_index_949069 ? add_987671 : sel_987668;
  assign add_987675 = sel_987672 + 8'h01;
  assign sel_987676 = array_index_987283 == array_index_949075 ? add_987675 : sel_987672;
  assign add_987679 = sel_987676 + 8'h01;
  assign sel_987680 = array_index_987283 == array_index_949081 ? add_987679 : sel_987676;
  assign add_987684 = sel_987680 + 8'h01;
  assign array_index_987685 = set1_unflattened[7'h61];
  assign sel_987686 = array_index_987283 == array_index_949087 ? add_987684 : sel_987680;
  assign add_987689 = sel_987686 + 8'h01;
  assign sel_987690 = array_index_987685 == array_index_948483 ? add_987689 : sel_987686;
  assign add_987693 = sel_987690 + 8'h01;
  assign sel_987694 = array_index_987685 == array_index_948487 ? add_987693 : sel_987690;
  assign add_987697 = sel_987694 + 8'h01;
  assign sel_987698 = array_index_987685 == array_index_948495 ? add_987697 : sel_987694;
  assign add_987701 = sel_987698 + 8'h01;
  assign sel_987702 = array_index_987685 == array_index_948503 ? add_987701 : sel_987698;
  assign add_987705 = sel_987702 + 8'h01;
  assign sel_987706 = array_index_987685 == array_index_948511 ? add_987705 : sel_987702;
  assign add_987709 = sel_987706 + 8'h01;
  assign sel_987710 = array_index_987685 == array_index_948519 ? add_987709 : sel_987706;
  assign add_987713 = sel_987710 + 8'h01;
  assign sel_987714 = array_index_987685 == array_index_948527 ? add_987713 : sel_987710;
  assign add_987717 = sel_987714 + 8'h01;
  assign sel_987718 = array_index_987685 == array_index_948535 ? add_987717 : sel_987714;
  assign add_987721 = sel_987718 + 8'h01;
  assign sel_987722 = array_index_987685 == array_index_948541 ? add_987721 : sel_987718;
  assign add_987725 = sel_987722 + 8'h01;
  assign sel_987726 = array_index_987685 == array_index_948547 ? add_987725 : sel_987722;
  assign add_987729 = sel_987726 + 8'h01;
  assign sel_987730 = array_index_987685 == array_index_948553 ? add_987729 : sel_987726;
  assign add_987733 = sel_987730 + 8'h01;
  assign sel_987734 = array_index_987685 == array_index_948559 ? add_987733 : sel_987730;
  assign add_987737 = sel_987734 + 8'h01;
  assign sel_987738 = array_index_987685 == array_index_948565 ? add_987737 : sel_987734;
  assign add_987741 = sel_987738 + 8'h01;
  assign sel_987742 = array_index_987685 == array_index_948571 ? add_987741 : sel_987738;
  assign add_987745 = sel_987742 + 8'h01;
  assign sel_987746 = array_index_987685 == array_index_948577 ? add_987745 : sel_987742;
  assign add_987749 = sel_987746 + 8'h01;
  assign sel_987750 = array_index_987685 == array_index_948583 ? add_987749 : sel_987746;
  assign add_987753 = sel_987750 + 8'h01;
  assign sel_987754 = array_index_987685 == array_index_948589 ? add_987753 : sel_987750;
  assign add_987757 = sel_987754 + 8'h01;
  assign sel_987758 = array_index_987685 == array_index_948595 ? add_987757 : sel_987754;
  assign add_987761 = sel_987758 + 8'h01;
  assign sel_987762 = array_index_987685 == array_index_948601 ? add_987761 : sel_987758;
  assign add_987765 = sel_987762 + 8'h01;
  assign sel_987766 = array_index_987685 == array_index_948607 ? add_987765 : sel_987762;
  assign add_987769 = sel_987766 + 8'h01;
  assign sel_987770 = array_index_987685 == array_index_948613 ? add_987769 : sel_987766;
  assign add_987773 = sel_987770 + 8'h01;
  assign sel_987774 = array_index_987685 == array_index_948619 ? add_987773 : sel_987770;
  assign add_987777 = sel_987774 + 8'h01;
  assign sel_987778 = array_index_987685 == array_index_948625 ? add_987777 : sel_987774;
  assign add_987781 = sel_987778 + 8'h01;
  assign sel_987782 = array_index_987685 == array_index_948631 ? add_987781 : sel_987778;
  assign add_987785 = sel_987782 + 8'h01;
  assign sel_987786 = array_index_987685 == array_index_948637 ? add_987785 : sel_987782;
  assign add_987789 = sel_987786 + 8'h01;
  assign sel_987790 = array_index_987685 == array_index_948643 ? add_987789 : sel_987786;
  assign add_987793 = sel_987790 + 8'h01;
  assign sel_987794 = array_index_987685 == array_index_948649 ? add_987793 : sel_987790;
  assign add_987797 = sel_987794 + 8'h01;
  assign sel_987798 = array_index_987685 == array_index_948655 ? add_987797 : sel_987794;
  assign add_987801 = sel_987798 + 8'h01;
  assign sel_987802 = array_index_987685 == array_index_948661 ? add_987801 : sel_987798;
  assign add_987805 = sel_987802 + 8'h01;
  assign sel_987806 = array_index_987685 == array_index_948667 ? add_987805 : sel_987802;
  assign add_987809 = sel_987806 + 8'h01;
  assign sel_987810 = array_index_987685 == array_index_948673 ? add_987809 : sel_987806;
  assign add_987813 = sel_987810 + 8'h01;
  assign sel_987814 = array_index_987685 == array_index_948679 ? add_987813 : sel_987810;
  assign add_987817 = sel_987814 + 8'h01;
  assign sel_987818 = array_index_987685 == array_index_948685 ? add_987817 : sel_987814;
  assign add_987821 = sel_987818 + 8'h01;
  assign sel_987822 = array_index_987685 == array_index_948691 ? add_987821 : sel_987818;
  assign add_987825 = sel_987822 + 8'h01;
  assign sel_987826 = array_index_987685 == array_index_948697 ? add_987825 : sel_987822;
  assign add_987829 = sel_987826 + 8'h01;
  assign sel_987830 = array_index_987685 == array_index_948703 ? add_987829 : sel_987826;
  assign add_987833 = sel_987830 + 8'h01;
  assign sel_987834 = array_index_987685 == array_index_948709 ? add_987833 : sel_987830;
  assign add_987837 = sel_987834 + 8'h01;
  assign sel_987838 = array_index_987685 == array_index_948715 ? add_987837 : sel_987834;
  assign add_987841 = sel_987838 + 8'h01;
  assign sel_987842 = array_index_987685 == array_index_948721 ? add_987841 : sel_987838;
  assign add_987845 = sel_987842 + 8'h01;
  assign sel_987846 = array_index_987685 == array_index_948727 ? add_987845 : sel_987842;
  assign add_987849 = sel_987846 + 8'h01;
  assign sel_987850 = array_index_987685 == array_index_948733 ? add_987849 : sel_987846;
  assign add_987853 = sel_987850 + 8'h01;
  assign sel_987854 = array_index_987685 == array_index_948739 ? add_987853 : sel_987850;
  assign add_987857 = sel_987854 + 8'h01;
  assign sel_987858 = array_index_987685 == array_index_948745 ? add_987857 : sel_987854;
  assign add_987861 = sel_987858 + 8'h01;
  assign sel_987862 = array_index_987685 == array_index_948751 ? add_987861 : sel_987858;
  assign add_987865 = sel_987862 + 8'h01;
  assign sel_987866 = array_index_987685 == array_index_948757 ? add_987865 : sel_987862;
  assign add_987869 = sel_987866 + 8'h01;
  assign sel_987870 = array_index_987685 == array_index_948763 ? add_987869 : sel_987866;
  assign add_987873 = sel_987870 + 8'h01;
  assign sel_987874 = array_index_987685 == array_index_948769 ? add_987873 : sel_987870;
  assign add_987877 = sel_987874 + 8'h01;
  assign sel_987878 = array_index_987685 == array_index_948775 ? add_987877 : sel_987874;
  assign add_987881 = sel_987878 + 8'h01;
  assign sel_987882 = array_index_987685 == array_index_948781 ? add_987881 : sel_987878;
  assign add_987885 = sel_987882 + 8'h01;
  assign sel_987886 = array_index_987685 == array_index_948787 ? add_987885 : sel_987882;
  assign add_987889 = sel_987886 + 8'h01;
  assign sel_987890 = array_index_987685 == array_index_948793 ? add_987889 : sel_987886;
  assign add_987893 = sel_987890 + 8'h01;
  assign sel_987894 = array_index_987685 == array_index_948799 ? add_987893 : sel_987890;
  assign add_987897 = sel_987894 + 8'h01;
  assign sel_987898 = array_index_987685 == array_index_948805 ? add_987897 : sel_987894;
  assign add_987901 = sel_987898 + 8'h01;
  assign sel_987902 = array_index_987685 == array_index_948811 ? add_987901 : sel_987898;
  assign add_987905 = sel_987902 + 8'h01;
  assign sel_987906 = array_index_987685 == array_index_948817 ? add_987905 : sel_987902;
  assign add_987909 = sel_987906 + 8'h01;
  assign sel_987910 = array_index_987685 == array_index_948823 ? add_987909 : sel_987906;
  assign add_987913 = sel_987910 + 8'h01;
  assign sel_987914 = array_index_987685 == array_index_948829 ? add_987913 : sel_987910;
  assign add_987917 = sel_987914 + 8'h01;
  assign sel_987918 = array_index_987685 == array_index_948835 ? add_987917 : sel_987914;
  assign add_987921 = sel_987918 + 8'h01;
  assign sel_987922 = array_index_987685 == array_index_948841 ? add_987921 : sel_987918;
  assign add_987925 = sel_987922 + 8'h01;
  assign sel_987926 = array_index_987685 == array_index_948847 ? add_987925 : sel_987922;
  assign add_987929 = sel_987926 + 8'h01;
  assign sel_987930 = array_index_987685 == array_index_948853 ? add_987929 : sel_987926;
  assign add_987933 = sel_987930 + 8'h01;
  assign sel_987934 = array_index_987685 == array_index_948859 ? add_987933 : sel_987930;
  assign add_987937 = sel_987934 + 8'h01;
  assign sel_987938 = array_index_987685 == array_index_948865 ? add_987937 : sel_987934;
  assign add_987941 = sel_987938 + 8'h01;
  assign sel_987942 = array_index_987685 == array_index_948871 ? add_987941 : sel_987938;
  assign add_987945 = sel_987942 + 8'h01;
  assign sel_987946 = array_index_987685 == array_index_948877 ? add_987945 : sel_987942;
  assign add_987949 = sel_987946 + 8'h01;
  assign sel_987950 = array_index_987685 == array_index_948883 ? add_987949 : sel_987946;
  assign add_987953 = sel_987950 + 8'h01;
  assign sel_987954 = array_index_987685 == array_index_948889 ? add_987953 : sel_987950;
  assign add_987957 = sel_987954 + 8'h01;
  assign sel_987958 = array_index_987685 == array_index_948895 ? add_987957 : sel_987954;
  assign add_987961 = sel_987958 + 8'h01;
  assign sel_987962 = array_index_987685 == array_index_948901 ? add_987961 : sel_987958;
  assign add_987965 = sel_987962 + 8'h01;
  assign sel_987966 = array_index_987685 == array_index_948907 ? add_987965 : sel_987962;
  assign add_987969 = sel_987966 + 8'h01;
  assign sel_987970 = array_index_987685 == array_index_948913 ? add_987969 : sel_987966;
  assign add_987973 = sel_987970 + 8'h01;
  assign sel_987974 = array_index_987685 == array_index_948919 ? add_987973 : sel_987970;
  assign add_987977 = sel_987974 + 8'h01;
  assign sel_987978 = array_index_987685 == array_index_948925 ? add_987977 : sel_987974;
  assign add_987981 = sel_987978 + 8'h01;
  assign sel_987982 = array_index_987685 == array_index_948931 ? add_987981 : sel_987978;
  assign add_987985 = sel_987982 + 8'h01;
  assign sel_987986 = array_index_987685 == array_index_948937 ? add_987985 : sel_987982;
  assign add_987989 = sel_987986 + 8'h01;
  assign sel_987990 = array_index_987685 == array_index_948943 ? add_987989 : sel_987986;
  assign add_987993 = sel_987990 + 8'h01;
  assign sel_987994 = array_index_987685 == array_index_948949 ? add_987993 : sel_987990;
  assign add_987997 = sel_987994 + 8'h01;
  assign sel_987998 = array_index_987685 == array_index_948955 ? add_987997 : sel_987994;
  assign add_988001 = sel_987998 + 8'h01;
  assign sel_988002 = array_index_987685 == array_index_948961 ? add_988001 : sel_987998;
  assign add_988005 = sel_988002 + 8'h01;
  assign sel_988006 = array_index_987685 == array_index_948967 ? add_988005 : sel_988002;
  assign add_988009 = sel_988006 + 8'h01;
  assign sel_988010 = array_index_987685 == array_index_948973 ? add_988009 : sel_988006;
  assign add_988013 = sel_988010 + 8'h01;
  assign sel_988014 = array_index_987685 == array_index_948979 ? add_988013 : sel_988010;
  assign add_988017 = sel_988014 + 8'h01;
  assign sel_988018 = array_index_987685 == array_index_948985 ? add_988017 : sel_988014;
  assign add_988021 = sel_988018 + 8'h01;
  assign sel_988022 = array_index_987685 == array_index_948991 ? add_988021 : sel_988018;
  assign add_988025 = sel_988022 + 8'h01;
  assign sel_988026 = array_index_987685 == array_index_948997 ? add_988025 : sel_988022;
  assign add_988029 = sel_988026 + 8'h01;
  assign sel_988030 = array_index_987685 == array_index_949003 ? add_988029 : sel_988026;
  assign add_988033 = sel_988030 + 8'h01;
  assign sel_988034 = array_index_987685 == array_index_949009 ? add_988033 : sel_988030;
  assign add_988037 = sel_988034 + 8'h01;
  assign sel_988038 = array_index_987685 == array_index_949015 ? add_988037 : sel_988034;
  assign add_988041 = sel_988038 + 8'h01;
  assign sel_988042 = array_index_987685 == array_index_949021 ? add_988041 : sel_988038;
  assign add_988045 = sel_988042 + 8'h01;
  assign sel_988046 = array_index_987685 == array_index_949027 ? add_988045 : sel_988042;
  assign add_988049 = sel_988046 + 8'h01;
  assign sel_988050 = array_index_987685 == array_index_949033 ? add_988049 : sel_988046;
  assign add_988053 = sel_988050 + 8'h01;
  assign sel_988054 = array_index_987685 == array_index_949039 ? add_988053 : sel_988050;
  assign add_988057 = sel_988054 + 8'h01;
  assign sel_988058 = array_index_987685 == array_index_949045 ? add_988057 : sel_988054;
  assign add_988061 = sel_988058 + 8'h01;
  assign sel_988062 = array_index_987685 == array_index_949051 ? add_988061 : sel_988058;
  assign add_988065 = sel_988062 + 8'h01;
  assign sel_988066 = array_index_987685 == array_index_949057 ? add_988065 : sel_988062;
  assign add_988069 = sel_988066 + 8'h01;
  assign sel_988070 = array_index_987685 == array_index_949063 ? add_988069 : sel_988066;
  assign add_988073 = sel_988070 + 8'h01;
  assign sel_988074 = array_index_987685 == array_index_949069 ? add_988073 : sel_988070;
  assign add_988077 = sel_988074 + 8'h01;
  assign sel_988078 = array_index_987685 == array_index_949075 ? add_988077 : sel_988074;
  assign add_988081 = sel_988078 + 8'h01;
  assign sel_988082 = array_index_987685 == array_index_949081 ? add_988081 : sel_988078;
  assign add_988086 = sel_988082 + 8'h01;
  assign array_index_988087 = set1_unflattened[7'h62];
  assign sel_988088 = array_index_987685 == array_index_949087 ? add_988086 : sel_988082;
  assign add_988091 = sel_988088 + 8'h01;
  assign sel_988092 = array_index_988087 == array_index_948483 ? add_988091 : sel_988088;
  assign add_988095 = sel_988092 + 8'h01;
  assign sel_988096 = array_index_988087 == array_index_948487 ? add_988095 : sel_988092;
  assign add_988099 = sel_988096 + 8'h01;
  assign sel_988100 = array_index_988087 == array_index_948495 ? add_988099 : sel_988096;
  assign add_988103 = sel_988100 + 8'h01;
  assign sel_988104 = array_index_988087 == array_index_948503 ? add_988103 : sel_988100;
  assign add_988107 = sel_988104 + 8'h01;
  assign sel_988108 = array_index_988087 == array_index_948511 ? add_988107 : sel_988104;
  assign add_988111 = sel_988108 + 8'h01;
  assign sel_988112 = array_index_988087 == array_index_948519 ? add_988111 : sel_988108;
  assign add_988115 = sel_988112 + 8'h01;
  assign sel_988116 = array_index_988087 == array_index_948527 ? add_988115 : sel_988112;
  assign add_988119 = sel_988116 + 8'h01;
  assign sel_988120 = array_index_988087 == array_index_948535 ? add_988119 : sel_988116;
  assign add_988123 = sel_988120 + 8'h01;
  assign sel_988124 = array_index_988087 == array_index_948541 ? add_988123 : sel_988120;
  assign add_988127 = sel_988124 + 8'h01;
  assign sel_988128 = array_index_988087 == array_index_948547 ? add_988127 : sel_988124;
  assign add_988131 = sel_988128 + 8'h01;
  assign sel_988132 = array_index_988087 == array_index_948553 ? add_988131 : sel_988128;
  assign add_988135 = sel_988132 + 8'h01;
  assign sel_988136 = array_index_988087 == array_index_948559 ? add_988135 : sel_988132;
  assign add_988139 = sel_988136 + 8'h01;
  assign sel_988140 = array_index_988087 == array_index_948565 ? add_988139 : sel_988136;
  assign add_988143 = sel_988140 + 8'h01;
  assign sel_988144 = array_index_988087 == array_index_948571 ? add_988143 : sel_988140;
  assign add_988147 = sel_988144 + 8'h01;
  assign sel_988148 = array_index_988087 == array_index_948577 ? add_988147 : sel_988144;
  assign add_988151 = sel_988148 + 8'h01;
  assign sel_988152 = array_index_988087 == array_index_948583 ? add_988151 : sel_988148;
  assign add_988155 = sel_988152 + 8'h01;
  assign sel_988156 = array_index_988087 == array_index_948589 ? add_988155 : sel_988152;
  assign add_988159 = sel_988156 + 8'h01;
  assign sel_988160 = array_index_988087 == array_index_948595 ? add_988159 : sel_988156;
  assign add_988163 = sel_988160 + 8'h01;
  assign sel_988164 = array_index_988087 == array_index_948601 ? add_988163 : sel_988160;
  assign add_988167 = sel_988164 + 8'h01;
  assign sel_988168 = array_index_988087 == array_index_948607 ? add_988167 : sel_988164;
  assign add_988171 = sel_988168 + 8'h01;
  assign sel_988172 = array_index_988087 == array_index_948613 ? add_988171 : sel_988168;
  assign add_988175 = sel_988172 + 8'h01;
  assign sel_988176 = array_index_988087 == array_index_948619 ? add_988175 : sel_988172;
  assign add_988179 = sel_988176 + 8'h01;
  assign sel_988180 = array_index_988087 == array_index_948625 ? add_988179 : sel_988176;
  assign add_988183 = sel_988180 + 8'h01;
  assign sel_988184 = array_index_988087 == array_index_948631 ? add_988183 : sel_988180;
  assign add_988187 = sel_988184 + 8'h01;
  assign sel_988188 = array_index_988087 == array_index_948637 ? add_988187 : sel_988184;
  assign add_988191 = sel_988188 + 8'h01;
  assign sel_988192 = array_index_988087 == array_index_948643 ? add_988191 : sel_988188;
  assign add_988195 = sel_988192 + 8'h01;
  assign sel_988196 = array_index_988087 == array_index_948649 ? add_988195 : sel_988192;
  assign add_988199 = sel_988196 + 8'h01;
  assign sel_988200 = array_index_988087 == array_index_948655 ? add_988199 : sel_988196;
  assign add_988203 = sel_988200 + 8'h01;
  assign sel_988204 = array_index_988087 == array_index_948661 ? add_988203 : sel_988200;
  assign add_988207 = sel_988204 + 8'h01;
  assign sel_988208 = array_index_988087 == array_index_948667 ? add_988207 : sel_988204;
  assign add_988211 = sel_988208 + 8'h01;
  assign sel_988212 = array_index_988087 == array_index_948673 ? add_988211 : sel_988208;
  assign add_988215 = sel_988212 + 8'h01;
  assign sel_988216 = array_index_988087 == array_index_948679 ? add_988215 : sel_988212;
  assign add_988219 = sel_988216 + 8'h01;
  assign sel_988220 = array_index_988087 == array_index_948685 ? add_988219 : sel_988216;
  assign add_988223 = sel_988220 + 8'h01;
  assign sel_988224 = array_index_988087 == array_index_948691 ? add_988223 : sel_988220;
  assign add_988227 = sel_988224 + 8'h01;
  assign sel_988228 = array_index_988087 == array_index_948697 ? add_988227 : sel_988224;
  assign add_988231 = sel_988228 + 8'h01;
  assign sel_988232 = array_index_988087 == array_index_948703 ? add_988231 : sel_988228;
  assign add_988235 = sel_988232 + 8'h01;
  assign sel_988236 = array_index_988087 == array_index_948709 ? add_988235 : sel_988232;
  assign add_988239 = sel_988236 + 8'h01;
  assign sel_988240 = array_index_988087 == array_index_948715 ? add_988239 : sel_988236;
  assign add_988243 = sel_988240 + 8'h01;
  assign sel_988244 = array_index_988087 == array_index_948721 ? add_988243 : sel_988240;
  assign add_988247 = sel_988244 + 8'h01;
  assign sel_988248 = array_index_988087 == array_index_948727 ? add_988247 : sel_988244;
  assign add_988251 = sel_988248 + 8'h01;
  assign sel_988252 = array_index_988087 == array_index_948733 ? add_988251 : sel_988248;
  assign add_988255 = sel_988252 + 8'h01;
  assign sel_988256 = array_index_988087 == array_index_948739 ? add_988255 : sel_988252;
  assign add_988259 = sel_988256 + 8'h01;
  assign sel_988260 = array_index_988087 == array_index_948745 ? add_988259 : sel_988256;
  assign add_988263 = sel_988260 + 8'h01;
  assign sel_988264 = array_index_988087 == array_index_948751 ? add_988263 : sel_988260;
  assign add_988267 = sel_988264 + 8'h01;
  assign sel_988268 = array_index_988087 == array_index_948757 ? add_988267 : sel_988264;
  assign add_988271 = sel_988268 + 8'h01;
  assign sel_988272 = array_index_988087 == array_index_948763 ? add_988271 : sel_988268;
  assign add_988275 = sel_988272 + 8'h01;
  assign sel_988276 = array_index_988087 == array_index_948769 ? add_988275 : sel_988272;
  assign add_988279 = sel_988276 + 8'h01;
  assign sel_988280 = array_index_988087 == array_index_948775 ? add_988279 : sel_988276;
  assign add_988283 = sel_988280 + 8'h01;
  assign sel_988284 = array_index_988087 == array_index_948781 ? add_988283 : sel_988280;
  assign add_988287 = sel_988284 + 8'h01;
  assign sel_988288 = array_index_988087 == array_index_948787 ? add_988287 : sel_988284;
  assign add_988291 = sel_988288 + 8'h01;
  assign sel_988292 = array_index_988087 == array_index_948793 ? add_988291 : sel_988288;
  assign add_988295 = sel_988292 + 8'h01;
  assign sel_988296 = array_index_988087 == array_index_948799 ? add_988295 : sel_988292;
  assign add_988299 = sel_988296 + 8'h01;
  assign sel_988300 = array_index_988087 == array_index_948805 ? add_988299 : sel_988296;
  assign add_988303 = sel_988300 + 8'h01;
  assign sel_988304 = array_index_988087 == array_index_948811 ? add_988303 : sel_988300;
  assign add_988307 = sel_988304 + 8'h01;
  assign sel_988308 = array_index_988087 == array_index_948817 ? add_988307 : sel_988304;
  assign add_988311 = sel_988308 + 8'h01;
  assign sel_988312 = array_index_988087 == array_index_948823 ? add_988311 : sel_988308;
  assign add_988315 = sel_988312 + 8'h01;
  assign sel_988316 = array_index_988087 == array_index_948829 ? add_988315 : sel_988312;
  assign add_988319 = sel_988316 + 8'h01;
  assign sel_988320 = array_index_988087 == array_index_948835 ? add_988319 : sel_988316;
  assign add_988323 = sel_988320 + 8'h01;
  assign sel_988324 = array_index_988087 == array_index_948841 ? add_988323 : sel_988320;
  assign add_988327 = sel_988324 + 8'h01;
  assign sel_988328 = array_index_988087 == array_index_948847 ? add_988327 : sel_988324;
  assign add_988331 = sel_988328 + 8'h01;
  assign sel_988332 = array_index_988087 == array_index_948853 ? add_988331 : sel_988328;
  assign add_988335 = sel_988332 + 8'h01;
  assign sel_988336 = array_index_988087 == array_index_948859 ? add_988335 : sel_988332;
  assign add_988339 = sel_988336 + 8'h01;
  assign sel_988340 = array_index_988087 == array_index_948865 ? add_988339 : sel_988336;
  assign add_988343 = sel_988340 + 8'h01;
  assign sel_988344 = array_index_988087 == array_index_948871 ? add_988343 : sel_988340;
  assign add_988347 = sel_988344 + 8'h01;
  assign sel_988348 = array_index_988087 == array_index_948877 ? add_988347 : sel_988344;
  assign add_988351 = sel_988348 + 8'h01;
  assign sel_988352 = array_index_988087 == array_index_948883 ? add_988351 : sel_988348;
  assign add_988355 = sel_988352 + 8'h01;
  assign sel_988356 = array_index_988087 == array_index_948889 ? add_988355 : sel_988352;
  assign add_988359 = sel_988356 + 8'h01;
  assign sel_988360 = array_index_988087 == array_index_948895 ? add_988359 : sel_988356;
  assign add_988363 = sel_988360 + 8'h01;
  assign sel_988364 = array_index_988087 == array_index_948901 ? add_988363 : sel_988360;
  assign add_988367 = sel_988364 + 8'h01;
  assign sel_988368 = array_index_988087 == array_index_948907 ? add_988367 : sel_988364;
  assign add_988371 = sel_988368 + 8'h01;
  assign sel_988372 = array_index_988087 == array_index_948913 ? add_988371 : sel_988368;
  assign add_988375 = sel_988372 + 8'h01;
  assign sel_988376 = array_index_988087 == array_index_948919 ? add_988375 : sel_988372;
  assign add_988379 = sel_988376 + 8'h01;
  assign sel_988380 = array_index_988087 == array_index_948925 ? add_988379 : sel_988376;
  assign add_988383 = sel_988380 + 8'h01;
  assign sel_988384 = array_index_988087 == array_index_948931 ? add_988383 : sel_988380;
  assign add_988387 = sel_988384 + 8'h01;
  assign sel_988388 = array_index_988087 == array_index_948937 ? add_988387 : sel_988384;
  assign add_988391 = sel_988388 + 8'h01;
  assign sel_988392 = array_index_988087 == array_index_948943 ? add_988391 : sel_988388;
  assign add_988395 = sel_988392 + 8'h01;
  assign sel_988396 = array_index_988087 == array_index_948949 ? add_988395 : sel_988392;
  assign add_988399 = sel_988396 + 8'h01;
  assign sel_988400 = array_index_988087 == array_index_948955 ? add_988399 : sel_988396;
  assign add_988403 = sel_988400 + 8'h01;
  assign sel_988404 = array_index_988087 == array_index_948961 ? add_988403 : sel_988400;
  assign add_988407 = sel_988404 + 8'h01;
  assign sel_988408 = array_index_988087 == array_index_948967 ? add_988407 : sel_988404;
  assign add_988411 = sel_988408 + 8'h01;
  assign sel_988412 = array_index_988087 == array_index_948973 ? add_988411 : sel_988408;
  assign add_988415 = sel_988412 + 8'h01;
  assign sel_988416 = array_index_988087 == array_index_948979 ? add_988415 : sel_988412;
  assign add_988419 = sel_988416 + 8'h01;
  assign sel_988420 = array_index_988087 == array_index_948985 ? add_988419 : sel_988416;
  assign add_988423 = sel_988420 + 8'h01;
  assign sel_988424 = array_index_988087 == array_index_948991 ? add_988423 : sel_988420;
  assign add_988427 = sel_988424 + 8'h01;
  assign sel_988428 = array_index_988087 == array_index_948997 ? add_988427 : sel_988424;
  assign add_988431 = sel_988428 + 8'h01;
  assign sel_988432 = array_index_988087 == array_index_949003 ? add_988431 : sel_988428;
  assign add_988435 = sel_988432 + 8'h01;
  assign sel_988436 = array_index_988087 == array_index_949009 ? add_988435 : sel_988432;
  assign add_988439 = sel_988436 + 8'h01;
  assign sel_988440 = array_index_988087 == array_index_949015 ? add_988439 : sel_988436;
  assign add_988443 = sel_988440 + 8'h01;
  assign sel_988444 = array_index_988087 == array_index_949021 ? add_988443 : sel_988440;
  assign add_988447 = sel_988444 + 8'h01;
  assign sel_988448 = array_index_988087 == array_index_949027 ? add_988447 : sel_988444;
  assign add_988451 = sel_988448 + 8'h01;
  assign sel_988452 = array_index_988087 == array_index_949033 ? add_988451 : sel_988448;
  assign add_988455 = sel_988452 + 8'h01;
  assign sel_988456 = array_index_988087 == array_index_949039 ? add_988455 : sel_988452;
  assign add_988459 = sel_988456 + 8'h01;
  assign sel_988460 = array_index_988087 == array_index_949045 ? add_988459 : sel_988456;
  assign add_988463 = sel_988460 + 8'h01;
  assign sel_988464 = array_index_988087 == array_index_949051 ? add_988463 : sel_988460;
  assign add_988467 = sel_988464 + 8'h01;
  assign sel_988468 = array_index_988087 == array_index_949057 ? add_988467 : sel_988464;
  assign add_988471 = sel_988468 + 8'h01;
  assign sel_988472 = array_index_988087 == array_index_949063 ? add_988471 : sel_988468;
  assign add_988475 = sel_988472 + 8'h01;
  assign sel_988476 = array_index_988087 == array_index_949069 ? add_988475 : sel_988472;
  assign add_988479 = sel_988476 + 8'h01;
  assign sel_988480 = array_index_988087 == array_index_949075 ? add_988479 : sel_988476;
  assign add_988483 = sel_988480 + 8'h01;
  assign sel_988484 = array_index_988087 == array_index_949081 ? add_988483 : sel_988480;
  assign add_988488 = sel_988484 + 8'h01;
  assign array_index_988489 = set1_unflattened[7'h63];
  assign sel_988490 = array_index_988087 == array_index_949087 ? add_988488 : sel_988484;
  assign add_988493 = sel_988490 + 8'h01;
  assign sel_988494 = array_index_988489 == array_index_948483 ? add_988493 : sel_988490;
  assign add_988497 = sel_988494 + 8'h01;
  assign sel_988498 = array_index_988489 == array_index_948487 ? add_988497 : sel_988494;
  assign add_988501 = sel_988498 + 8'h01;
  assign sel_988502 = array_index_988489 == array_index_948495 ? add_988501 : sel_988498;
  assign add_988505 = sel_988502 + 8'h01;
  assign sel_988506 = array_index_988489 == array_index_948503 ? add_988505 : sel_988502;
  assign add_988509 = sel_988506 + 8'h01;
  assign sel_988510 = array_index_988489 == array_index_948511 ? add_988509 : sel_988506;
  assign add_988513 = sel_988510 + 8'h01;
  assign sel_988514 = array_index_988489 == array_index_948519 ? add_988513 : sel_988510;
  assign add_988517 = sel_988514 + 8'h01;
  assign sel_988518 = array_index_988489 == array_index_948527 ? add_988517 : sel_988514;
  assign add_988521 = sel_988518 + 8'h01;
  assign sel_988522 = array_index_988489 == array_index_948535 ? add_988521 : sel_988518;
  assign add_988525 = sel_988522 + 8'h01;
  assign sel_988526 = array_index_988489 == array_index_948541 ? add_988525 : sel_988522;
  assign add_988529 = sel_988526 + 8'h01;
  assign sel_988530 = array_index_988489 == array_index_948547 ? add_988529 : sel_988526;
  assign add_988533 = sel_988530 + 8'h01;
  assign sel_988534 = array_index_988489 == array_index_948553 ? add_988533 : sel_988530;
  assign add_988537 = sel_988534 + 8'h01;
  assign sel_988538 = array_index_988489 == array_index_948559 ? add_988537 : sel_988534;
  assign add_988541 = sel_988538 + 8'h01;
  assign sel_988542 = array_index_988489 == array_index_948565 ? add_988541 : sel_988538;
  assign add_988545 = sel_988542 + 8'h01;
  assign sel_988546 = array_index_988489 == array_index_948571 ? add_988545 : sel_988542;
  assign add_988549 = sel_988546 + 8'h01;
  assign sel_988550 = array_index_988489 == array_index_948577 ? add_988549 : sel_988546;
  assign add_988553 = sel_988550 + 8'h01;
  assign sel_988554 = array_index_988489 == array_index_948583 ? add_988553 : sel_988550;
  assign add_988557 = sel_988554 + 8'h01;
  assign sel_988558 = array_index_988489 == array_index_948589 ? add_988557 : sel_988554;
  assign add_988561 = sel_988558 + 8'h01;
  assign sel_988562 = array_index_988489 == array_index_948595 ? add_988561 : sel_988558;
  assign add_988565 = sel_988562 + 8'h01;
  assign sel_988566 = array_index_988489 == array_index_948601 ? add_988565 : sel_988562;
  assign add_988569 = sel_988566 + 8'h01;
  assign sel_988570 = array_index_988489 == array_index_948607 ? add_988569 : sel_988566;
  assign add_988573 = sel_988570 + 8'h01;
  assign sel_988574 = array_index_988489 == array_index_948613 ? add_988573 : sel_988570;
  assign add_988577 = sel_988574 + 8'h01;
  assign sel_988578 = array_index_988489 == array_index_948619 ? add_988577 : sel_988574;
  assign add_988581 = sel_988578 + 8'h01;
  assign sel_988582 = array_index_988489 == array_index_948625 ? add_988581 : sel_988578;
  assign add_988585 = sel_988582 + 8'h01;
  assign sel_988586 = array_index_988489 == array_index_948631 ? add_988585 : sel_988582;
  assign add_988589 = sel_988586 + 8'h01;
  assign sel_988590 = array_index_988489 == array_index_948637 ? add_988589 : sel_988586;
  assign add_988593 = sel_988590 + 8'h01;
  assign sel_988594 = array_index_988489 == array_index_948643 ? add_988593 : sel_988590;
  assign add_988597 = sel_988594 + 8'h01;
  assign sel_988598 = array_index_988489 == array_index_948649 ? add_988597 : sel_988594;
  assign add_988601 = sel_988598 + 8'h01;
  assign sel_988602 = array_index_988489 == array_index_948655 ? add_988601 : sel_988598;
  assign add_988605 = sel_988602 + 8'h01;
  assign sel_988606 = array_index_988489 == array_index_948661 ? add_988605 : sel_988602;
  assign add_988609 = sel_988606 + 8'h01;
  assign sel_988610 = array_index_988489 == array_index_948667 ? add_988609 : sel_988606;
  assign add_988613 = sel_988610 + 8'h01;
  assign sel_988614 = array_index_988489 == array_index_948673 ? add_988613 : sel_988610;
  assign add_988617 = sel_988614 + 8'h01;
  assign sel_988618 = array_index_988489 == array_index_948679 ? add_988617 : sel_988614;
  assign add_988621 = sel_988618 + 8'h01;
  assign sel_988622 = array_index_988489 == array_index_948685 ? add_988621 : sel_988618;
  assign add_988625 = sel_988622 + 8'h01;
  assign sel_988626 = array_index_988489 == array_index_948691 ? add_988625 : sel_988622;
  assign add_988629 = sel_988626 + 8'h01;
  assign sel_988630 = array_index_988489 == array_index_948697 ? add_988629 : sel_988626;
  assign add_988633 = sel_988630 + 8'h01;
  assign sel_988634 = array_index_988489 == array_index_948703 ? add_988633 : sel_988630;
  assign add_988637 = sel_988634 + 8'h01;
  assign sel_988638 = array_index_988489 == array_index_948709 ? add_988637 : sel_988634;
  assign add_988641 = sel_988638 + 8'h01;
  assign sel_988642 = array_index_988489 == array_index_948715 ? add_988641 : sel_988638;
  assign add_988645 = sel_988642 + 8'h01;
  assign sel_988646 = array_index_988489 == array_index_948721 ? add_988645 : sel_988642;
  assign add_988649 = sel_988646 + 8'h01;
  assign sel_988650 = array_index_988489 == array_index_948727 ? add_988649 : sel_988646;
  assign add_988653 = sel_988650 + 8'h01;
  assign sel_988654 = array_index_988489 == array_index_948733 ? add_988653 : sel_988650;
  assign add_988657 = sel_988654 + 8'h01;
  assign sel_988658 = array_index_988489 == array_index_948739 ? add_988657 : sel_988654;
  assign add_988661 = sel_988658 + 8'h01;
  assign sel_988662 = array_index_988489 == array_index_948745 ? add_988661 : sel_988658;
  assign add_988665 = sel_988662 + 8'h01;
  assign sel_988666 = array_index_988489 == array_index_948751 ? add_988665 : sel_988662;
  assign add_988669 = sel_988666 + 8'h01;
  assign sel_988670 = array_index_988489 == array_index_948757 ? add_988669 : sel_988666;
  assign add_988673 = sel_988670 + 8'h01;
  assign sel_988674 = array_index_988489 == array_index_948763 ? add_988673 : sel_988670;
  assign add_988677 = sel_988674 + 8'h01;
  assign sel_988678 = array_index_988489 == array_index_948769 ? add_988677 : sel_988674;
  assign add_988681 = sel_988678 + 8'h01;
  assign sel_988682 = array_index_988489 == array_index_948775 ? add_988681 : sel_988678;
  assign add_988685 = sel_988682 + 8'h01;
  assign sel_988686 = array_index_988489 == array_index_948781 ? add_988685 : sel_988682;
  assign add_988689 = sel_988686 + 8'h01;
  assign sel_988690 = array_index_988489 == array_index_948787 ? add_988689 : sel_988686;
  assign add_988693 = sel_988690 + 8'h01;
  assign sel_988694 = array_index_988489 == array_index_948793 ? add_988693 : sel_988690;
  assign add_988697 = sel_988694 + 8'h01;
  assign sel_988698 = array_index_988489 == array_index_948799 ? add_988697 : sel_988694;
  assign add_988701 = sel_988698 + 8'h01;
  assign sel_988702 = array_index_988489 == array_index_948805 ? add_988701 : sel_988698;
  assign add_988705 = sel_988702 + 8'h01;
  assign sel_988706 = array_index_988489 == array_index_948811 ? add_988705 : sel_988702;
  assign add_988709 = sel_988706 + 8'h01;
  assign sel_988710 = array_index_988489 == array_index_948817 ? add_988709 : sel_988706;
  assign add_988713 = sel_988710 + 8'h01;
  assign sel_988714 = array_index_988489 == array_index_948823 ? add_988713 : sel_988710;
  assign add_988717 = sel_988714 + 8'h01;
  assign sel_988718 = array_index_988489 == array_index_948829 ? add_988717 : sel_988714;
  assign add_988721 = sel_988718 + 8'h01;
  assign sel_988722 = array_index_988489 == array_index_948835 ? add_988721 : sel_988718;
  assign add_988725 = sel_988722 + 8'h01;
  assign sel_988726 = array_index_988489 == array_index_948841 ? add_988725 : sel_988722;
  assign add_988729 = sel_988726 + 8'h01;
  assign sel_988730 = array_index_988489 == array_index_948847 ? add_988729 : sel_988726;
  assign add_988733 = sel_988730 + 8'h01;
  assign sel_988734 = array_index_988489 == array_index_948853 ? add_988733 : sel_988730;
  assign add_988737 = sel_988734 + 8'h01;
  assign sel_988738 = array_index_988489 == array_index_948859 ? add_988737 : sel_988734;
  assign add_988741 = sel_988738 + 8'h01;
  assign sel_988742 = array_index_988489 == array_index_948865 ? add_988741 : sel_988738;
  assign add_988745 = sel_988742 + 8'h01;
  assign sel_988746 = array_index_988489 == array_index_948871 ? add_988745 : sel_988742;
  assign add_988749 = sel_988746 + 8'h01;
  assign sel_988750 = array_index_988489 == array_index_948877 ? add_988749 : sel_988746;
  assign add_988753 = sel_988750 + 8'h01;
  assign sel_988754 = array_index_988489 == array_index_948883 ? add_988753 : sel_988750;
  assign add_988757 = sel_988754 + 8'h01;
  assign sel_988758 = array_index_988489 == array_index_948889 ? add_988757 : sel_988754;
  assign add_988761 = sel_988758 + 8'h01;
  assign sel_988762 = array_index_988489 == array_index_948895 ? add_988761 : sel_988758;
  assign add_988765 = sel_988762 + 8'h01;
  assign sel_988766 = array_index_988489 == array_index_948901 ? add_988765 : sel_988762;
  assign add_988769 = sel_988766 + 8'h01;
  assign sel_988770 = array_index_988489 == array_index_948907 ? add_988769 : sel_988766;
  assign add_988773 = sel_988770 + 8'h01;
  assign sel_988774 = array_index_988489 == array_index_948913 ? add_988773 : sel_988770;
  assign add_988777 = sel_988774 + 8'h01;
  assign sel_988778 = array_index_988489 == array_index_948919 ? add_988777 : sel_988774;
  assign add_988781 = sel_988778 + 8'h01;
  assign sel_988782 = array_index_988489 == array_index_948925 ? add_988781 : sel_988778;
  assign add_988785 = sel_988782 + 8'h01;
  assign sel_988786 = array_index_988489 == array_index_948931 ? add_988785 : sel_988782;
  assign add_988789 = sel_988786 + 8'h01;
  assign sel_988790 = array_index_988489 == array_index_948937 ? add_988789 : sel_988786;
  assign add_988793 = sel_988790 + 8'h01;
  assign sel_988794 = array_index_988489 == array_index_948943 ? add_988793 : sel_988790;
  assign add_988797 = sel_988794 + 8'h01;
  assign sel_988798 = array_index_988489 == array_index_948949 ? add_988797 : sel_988794;
  assign add_988801 = sel_988798 + 8'h01;
  assign sel_988802 = array_index_988489 == array_index_948955 ? add_988801 : sel_988798;
  assign add_988805 = sel_988802 + 8'h01;
  assign sel_988806 = array_index_988489 == array_index_948961 ? add_988805 : sel_988802;
  assign add_988809 = sel_988806 + 8'h01;
  assign sel_988810 = array_index_988489 == array_index_948967 ? add_988809 : sel_988806;
  assign add_988813 = sel_988810 + 8'h01;
  assign sel_988814 = array_index_988489 == array_index_948973 ? add_988813 : sel_988810;
  assign add_988817 = sel_988814 + 8'h01;
  assign sel_988818 = array_index_988489 == array_index_948979 ? add_988817 : sel_988814;
  assign add_988821 = sel_988818 + 8'h01;
  assign sel_988822 = array_index_988489 == array_index_948985 ? add_988821 : sel_988818;
  assign add_988825 = sel_988822 + 8'h01;
  assign sel_988826 = array_index_988489 == array_index_948991 ? add_988825 : sel_988822;
  assign add_988829 = sel_988826 + 8'h01;
  assign sel_988830 = array_index_988489 == array_index_948997 ? add_988829 : sel_988826;
  assign add_988833 = sel_988830 + 8'h01;
  assign sel_988834 = array_index_988489 == array_index_949003 ? add_988833 : sel_988830;
  assign add_988837 = sel_988834 + 8'h01;
  assign sel_988838 = array_index_988489 == array_index_949009 ? add_988837 : sel_988834;
  assign add_988841 = sel_988838 + 8'h01;
  assign sel_988842 = array_index_988489 == array_index_949015 ? add_988841 : sel_988838;
  assign add_988845 = sel_988842 + 8'h01;
  assign sel_988846 = array_index_988489 == array_index_949021 ? add_988845 : sel_988842;
  assign add_988849 = sel_988846 + 8'h01;
  assign sel_988850 = array_index_988489 == array_index_949027 ? add_988849 : sel_988846;
  assign add_988853 = sel_988850 + 8'h01;
  assign sel_988854 = array_index_988489 == array_index_949033 ? add_988853 : sel_988850;
  assign add_988857 = sel_988854 + 8'h01;
  assign sel_988858 = array_index_988489 == array_index_949039 ? add_988857 : sel_988854;
  assign add_988861 = sel_988858 + 8'h01;
  assign sel_988862 = array_index_988489 == array_index_949045 ? add_988861 : sel_988858;
  assign add_988865 = sel_988862 + 8'h01;
  assign sel_988866 = array_index_988489 == array_index_949051 ? add_988865 : sel_988862;
  assign add_988869 = sel_988866 + 8'h01;
  assign sel_988870 = array_index_988489 == array_index_949057 ? add_988869 : sel_988866;
  assign add_988873 = sel_988870 + 8'h01;
  assign sel_988874 = array_index_988489 == array_index_949063 ? add_988873 : sel_988870;
  assign add_988877 = sel_988874 + 8'h01;
  assign sel_988878 = array_index_988489 == array_index_949069 ? add_988877 : sel_988874;
  assign add_988881 = sel_988878 + 8'h01;
  assign sel_988882 = array_index_988489 == array_index_949075 ? add_988881 : sel_988878;
  assign add_988885 = sel_988882 + 8'h01;
  assign sel_988886 = array_index_988489 == array_index_949081 ? add_988885 : sel_988882;
  assign add_988889 = sel_988886 + 8'h01;
  assign out = {array_index_988489 == array_index_949087 ? add_988889 : sel_988886, {set1_unflattened[99], set1_unflattened[98], set1_unflattened[97], set1_unflattened[96], set1_unflattened[95], set1_unflattened[94], set1_unflattened[93], set1_unflattened[92], set1_unflattened[91], set1_unflattened[90], set1_unflattened[89], set1_unflattened[88], set1_unflattened[87], set1_unflattened[86], set1_unflattened[85], set1_unflattened[84], set1_unflattened[83], set1_unflattened[82], set1_unflattened[81], set1_unflattened[80], set1_unflattened[79], set1_unflattened[78], set1_unflattened[77], set1_unflattened[76], set1_unflattened[75], set1_unflattened[74], set1_unflattened[73], set1_unflattened[72], set1_unflattened[71], set1_unflattened[70], set1_unflattened[69], set1_unflattened[68], set1_unflattened[67], set1_unflattened[66], set1_unflattened[65], set1_unflattened[64], set1_unflattened[63], set1_unflattened[62], set1_unflattened[61], set1_unflattened[60], set1_unflattened[59], set1_unflattened[58], set1_unflattened[57], set1_unflattened[56], set1_unflattened[55], set1_unflattened[54], set1_unflattened[53], set1_unflattened[52], set1_unflattened[51], set1_unflattened[50], set1_unflattened[49], set1_unflattened[48], set1_unflattened[47], set1_unflattened[46], set1_unflattened[45], set1_unflattened[44], set1_unflattened[43], set1_unflattened[42], set1_unflattened[41], set1_unflattened[40], set1_unflattened[39], set1_unflattened[38], set1_unflattened[37], set1_unflattened[36], set1_unflattened[35], set1_unflattened[34], set1_unflattened[33], set1_unflattened[32], set1_unflattened[31], set1_unflattened[30], set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[99], set2_unflattened[98], set2_unflattened[97], set2_unflattened[96], set2_unflattened[95], set2_unflattened[94], set2_unflattened[93], set2_unflattened[92], set2_unflattened[91], set2_unflattened[90], set2_unflattened[89], set2_unflattened[88], set2_unflattened[87], set2_unflattened[86], set2_unflattened[85], set2_unflattened[84], set2_unflattened[83], set2_unflattened[82], set2_unflattened[81], set2_unflattened[80], set2_unflattened[79], set2_unflattened[78], set2_unflattened[77], set2_unflattened[76], set2_unflattened[75], set2_unflattened[74], set2_unflattened[73], set2_unflattened[72], set2_unflattened[71], set2_unflattened[70], set2_unflattened[69], set2_unflattened[68], set2_unflattened[67], set2_unflattened[66], set2_unflattened[65], set2_unflattened[64], set2_unflattened[63], set2_unflattened[62], set2_unflattened[61], set2_unflattened[60], set2_unflattened[59], set2_unflattened[58], set2_unflattened[57], set2_unflattened[56], set2_unflattened[55], set2_unflattened[54], set2_unflattened[53], set2_unflattened[52], set2_unflattened[51], set2_unflattened[50], set2_unflattened[49], set2_unflattened[48], set2_unflattened[47], set2_unflattened[46], set2_unflattened[45], set2_unflattened[44], set2_unflattened[43], set2_unflattened[42], set2_unflattened[41], set2_unflattened[40], set2_unflattened[39], set2_unflattened[38], set2_unflattened[37], set2_unflattened[36], set2_unflattened[35], set2_unflattened[34], set2_unflattened[33], set2_unflattened[32], set2_unflattened[31], set2_unflattened[30], set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
