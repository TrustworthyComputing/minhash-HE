module min_hash(
  input wire [1199:0] set1,
  input wire [1199:0] set2,
  output wire [2407:0] out
);
  wire [15:0] set1_unflattened[75];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  assign set1_unflattened[30] = set1[495:480];
  assign set1_unflattened[31] = set1[511:496];
  assign set1_unflattened[32] = set1[527:512];
  assign set1_unflattened[33] = set1[543:528];
  assign set1_unflattened[34] = set1[559:544];
  assign set1_unflattened[35] = set1[575:560];
  assign set1_unflattened[36] = set1[591:576];
  assign set1_unflattened[37] = set1[607:592];
  assign set1_unflattened[38] = set1[623:608];
  assign set1_unflattened[39] = set1[639:624];
  assign set1_unflattened[40] = set1[655:640];
  assign set1_unflattened[41] = set1[671:656];
  assign set1_unflattened[42] = set1[687:672];
  assign set1_unflattened[43] = set1[703:688];
  assign set1_unflattened[44] = set1[719:704];
  assign set1_unflattened[45] = set1[735:720];
  assign set1_unflattened[46] = set1[751:736];
  assign set1_unflattened[47] = set1[767:752];
  assign set1_unflattened[48] = set1[783:768];
  assign set1_unflattened[49] = set1[799:784];
  assign set1_unflattened[50] = set1[815:800];
  assign set1_unflattened[51] = set1[831:816];
  assign set1_unflattened[52] = set1[847:832];
  assign set1_unflattened[53] = set1[863:848];
  assign set1_unflattened[54] = set1[879:864];
  assign set1_unflattened[55] = set1[895:880];
  assign set1_unflattened[56] = set1[911:896];
  assign set1_unflattened[57] = set1[927:912];
  assign set1_unflattened[58] = set1[943:928];
  assign set1_unflattened[59] = set1[959:944];
  assign set1_unflattened[60] = set1[975:960];
  assign set1_unflattened[61] = set1[991:976];
  assign set1_unflattened[62] = set1[1007:992];
  assign set1_unflattened[63] = set1[1023:1008];
  assign set1_unflattened[64] = set1[1039:1024];
  assign set1_unflattened[65] = set1[1055:1040];
  assign set1_unflattened[66] = set1[1071:1056];
  assign set1_unflattened[67] = set1[1087:1072];
  assign set1_unflattened[68] = set1[1103:1088];
  assign set1_unflattened[69] = set1[1119:1104];
  assign set1_unflattened[70] = set1[1135:1120];
  assign set1_unflattened[71] = set1[1151:1136];
  assign set1_unflattened[72] = set1[1167:1152];
  assign set1_unflattened[73] = set1[1183:1168];
  assign set1_unflattened[74] = set1[1199:1184];
  wire [15:0] set2_unflattened[75];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  assign set2_unflattened[30] = set2[495:480];
  assign set2_unflattened[31] = set2[511:496];
  assign set2_unflattened[32] = set2[527:512];
  assign set2_unflattened[33] = set2[543:528];
  assign set2_unflattened[34] = set2[559:544];
  assign set2_unflattened[35] = set2[575:560];
  assign set2_unflattened[36] = set2[591:576];
  assign set2_unflattened[37] = set2[607:592];
  assign set2_unflattened[38] = set2[623:608];
  assign set2_unflattened[39] = set2[639:624];
  assign set2_unflattened[40] = set2[655:640];
  assign set2_unflattened[41] = set2[671:656];
  assign set2_unflattened[42] = set2[687:672];
  assign set2_unflattened[43] = set2[703:688];
  assign set2_unflattened[44] = set2[719:704];
  assign set2_unflattened[45] = set2[735:720];
  assign set2_unflattened[46] = set2[751:736];
  assign set2_unflattened[47] = set2[767:752];
  assign set2_unflattened[48] = set2[783:768];
  assign set2_unflattened[49] = set2[799:784];
  assign set2_unflattened[50] = set2[815:800];
  assign set2_unflattened[51] = set2[831:816];
  assign set2_unflattened[52] = set2[847:832];
  assign set2_unflattened[53] = set2[863:848];
  assign set2_unflattened[54] = set2[879:864];
  assign set2_unflattened[55] = set2[895:880];
  assign set2_unflattened[56] = set2[911:896];
  assign set2_unflattened[57] = set2[927:912];
  assign set2_unflattened[58] = set2[943:928];
  assign set2_unflattened[59] = set2[959:944];
  assign set2_unflattened[60] = set2[975:960];
  assign set2_unflattened[61] = set2[991:976];
  assign set2_unflattened[62] = set2[1007:992];
  assign set2_unflattened[63] = set2[1023:1008];
  assign set2_unflattened[64] = set2[1039:1024];
  assign set2_unflattened[65] = set2[1055:1040];
  assign set2_unflattened[66] = set2[1071:1056];
  assign set2_unflattened[67] = set2[1087:1072];
  assign set2_unflattened[68] = set2[1103:1088];
  assign set2_unflattened[69] = set2[1119:1104];
  assign set2_unflattened[70] = set2[1135:1120];
  assign set2_unflattened[71] = set2[1151:1136];
  assign set2_unflattened[72] = set2[1167:1152];
  assign set2_unflattened[73] = set2[1183:1168];
  assign set2_unflattened[74] = set2[1199:1184];
  wire [15:0] array_index_537011;
  wire [15:0] array_index_537012;
  wire [15:0] array_index_537016;
  wire [1:0] concat_537017;
  wire [1:0] add_537020;
  wire [15:0] array_index_537024;
  wire [2:0] concat_537025;
  wire [2:0] add_537028;
  wire [15:0] array_index_537032;
  wire [3:0] concat_537033;
  wire [3:0] add_537036;
  wire [15:0] array_index_537040;
  wire [4:0] concat_537041;
  wire [4:0] add_537044;
  wire [15:0] array_index_537048;
  wire [5:0] concat_537049;
  wire [5:0] add_537052;
  wire [15:0] array_index_537056;
  wire [6:0] concat_537057;
  wire [6:0] add_537060;
  wire [15:0] array_index_537064;
  wire [7:0] concat_537065;
  wire [7:0] add_537069;
  wire [15:0] array_index_537070;
  wire [7:0] sel_537071;
  wire [7:0] add_537075;
  wire [15:0] array_index_537076;
  wire [7:0] sel_537077;
  wire [7:0] add_537081;
  wire [15:0] array_index_537082;
  wire [7:0] sel_537083;
  wire [7:0] add_537087;
  wire [15:0] array_index_537088;
  wire [7:0] sel_537089;
  wire [7:0] add_537093;
  wire [15:0] array_index_537094;
  wire [7:0] sel_537095;
  wire [7:0] add_537099;
  wire [15:0] array_index_537100;
  wire [7:0] sel_537101;
  wire [7:0] add_537105;
  wire [15:0] array_index_537106;
  wire [7:0] sel_537107;
  wire [7:0] add_537111;
  wire [15:0] array_index_537112;
  wire [7:0] sel_537113;
  wire [7:0] add_537117;
  wire [15:0] array_index_537118;
  wire [7:0] sel_537119;
  wire [7:0] add_537123;
  wire [15:0] array_index_537124;
  wire [7:0] sel_537125;
  wire [7:0] add_537129;
  wire [15:0] array_index_537130;
  wire [7:0] sel_537131;
  wire [7:0] add_537135;
  wire [15:0] array_index_537136;
  wire [7:0] sel_537137;
  wire [7:0] add_537141;
  wire [15:0] array_index_537142;
  wire [7:0] sel_537143;
  wire [7:0] add_537147;
  wire [15:0] array_index_537148;
  wire [7:0] sel_537149;
  wire [7:0] add_537153;
  wire [15:0] array_index_537154;
  wire [7:0] sel_537155;
  wire [7:0] add_537159;
  wire [15:0] array_index_537160;
  wire [7:0] sel_537161;
  wire [7:0] add_537165;
  wire [15:0] array_index_537166;
  wire [7:0] sel_537167;
  wire [7:0] add_537171;
  wire [15:0] array_index_537172;
  wire [7:0] sel_537173;
  wire [7:0] add_537177;
  wire [15:0] array_index_537178;
  wire [7:0] sel_537179;
  wire [7:0] add_537183;
  wire [15:0] array_index_537184;
  wire [7:0] sel_537185;
  wire [7:0] add_537189;
  wire [15:0] array_index_537190;
  wire [7:0] sel_537191;
  wire [7:0] add_537195;
  wire [15:0] array_index_537196;
  wire [7:0] sel_537197;
  wire [7:0] add_537201;
  wire [15:0] array_index_537202;
  wire [7:0] sel_537203;
  wire [7:0] add_537207;
  wire [15:0] array_index_537208;
  wire [7:0] sel_537209;
  wire [7:0] add_537213;
  wire [15:0] array_index_537214;
  wire [7:0] sel_537215;
  wire [7:0] add_537219;
  wire [15:0] array_index_537220;
  wire [7:0] sel_537221;
  wire [7:0] add_537225;
  wire [15:0] array_index_537226;
  wire [7:0] sel_537227;
  wire [7:0] add_537231;
  wire [15:0] array_index_537232;
  wire [7:0] sel_537233;
  wire [7:0] add_537237;
  wire [15:0] array_index_537238;
  wire [7:0] sel_537239;
  wire [7:0] add_537243;
  wire [15:0] array_index_537244;
  wire [7:0] sel_537245;
  wire [7:0] add_537249;
  wire [15:0] array_index_537250;
  wire [7:0] sel_537251;
  wire [7:0] add_537255;
  wire [15:0] array_index_537256;
  wire [7:0] sel_537257;
  wire [7:0] add_537261;
  wire [15:0] array_index_537262;
  wire [7:0] sel_537263;
  wire [7:0] add_537267;
  wire [15:0] array_index_537268;
  wire [7:0] sel_537269;
  wire [7:0] add_537273;
  wire [15:0] array_index_537274;
  wire [7:0] sel_537275;
  wire [7:0] add_537279;
  wire [15:0] array_index_537280;
  wire [7:0] sel_537281;
  wire [7:0] add_537285;
  wire [15:0] array_index_537286;
  wire [7:0] sel_537287;
  wire [7:0] add_537291;
  wire [15:0] array_index_537292;
  wire [7:0] sel_537293;
  wire [7:0] add_537297;
  wire [15:0] array_index_537298;
  wire [7:0] sel_537299;
  wire [7:0] add_537303;
  wire [15:0] array_index_537304;
  wire [7:0] sel_537305;
  wire [7:0] add_537309;
  wire [15:0] array_index_537310;
  wire [7:0] sel_537311;
  wire [7:0] add_537315;
  wire [15:0] array_index_537316;
  wire [7:0] sel_537317;
  wire [7:0] add_537321;
  wire [15:0] array_index_537322;
  wire [7:0] sel_537323;
  wire [7:0] add_537327;
  wire [15:0] array_index_537328;
  wire [7:0] sel_537329;
  wire [7:0] add_537333;
  wire [15:0] array_index_537334;
  wire [7:0] sel_537335;
  wire [7:0] add_537339;
  wire [15:0] array_index_537340;
  wire [7:0] sel_537341;
  wire [7:0] add_537345;
  wire [15:0] array_index_537346;
  wire [7:0] sel_537347;
  wire [7:0] add_537351;
  wire [15:0] array_index_537352;
  wire [7:0] sel_537353;
  wire [7:0] add_537357;
  wire [15:0] array_index_537358;
  wire [7:0] sel_537359;
  wire [7:0] add_537363;
  wire [15:0] array_index_537364;
  wire [7:0] sel_537365;
  wire [7:0] add_537369;
  wire [15:0] array_index_537370;
  wire [7:0] sel_537371;
  wire [7:0] add_537375;
  wire [15:0] array_index_537376;
  wire [7:0] sel_537377;
  wire [7:0] add_537381;
  wire [15:0] array_index_537382;
  wire [7:0] sel_537383;
  wire [7:0] add_537387;
  wire [15:0] array_index_537388;
  wire [7:0] sel_537389;
  wire [7:0] add_537393;
  wire [15:0] array_index_537394;
  wire [7:0] sel_537395;
  wire [7:0] add_537399;
  wire [15:0] array_index_537400;
  wire [7:0] sel_537401;
  wire [7:0] add_537405;
  wire [15:0] array_index_537406;
  wire [7:0] sel_537407;
  wire [7:0] add_537411;
  wire [15:0] array_index_537412;
  wire [7:0] sel_537413;
  wire [7:0] add_537417;
  wire [15:0] array_index_537418;
  wire [7:0] sel_537419;
  wire [7:0] add_537423;
  wire [15:0] array_index_537424;
  wire [7:0] sel_537425;
  wire [7:0] add_537429;
  wire [15:0] array_index_537430;
  wire [7:0] sel_537431;
  wire [7:0] add_537435;
  wire [15:0] array_index_537436;
  wire [7:0] sel_537437;
  wire [7:0] add_537441;
  wire [15:0] array_index_537442;
  wire [7:0] sel_537443;
  wire [7:0] add_537447;
  wire [15:0] array_index_537448;
  wire [7:0] sel_537449;
  wire [7:0] add_537453;
  wire [15:0] array_index_537454;
  wire [7:0] sel_537455;
  wire [7:0] add_537459;
  wire [15:0] array_index_537460;
  wire [7:0] sel_537461;
  wire [7:0] add_537465;
  wire [15:0] array_index_537466;
  wire [7:0] sel_537467;
  wire [7:0] add_537471;
  wire [15:0] array_index_537472;
  wire [7:0] sel_537473;
  wire [7:0] add_537476;
  wire [7:0] sel_537477;
  wire [7:0] add_537480;
  wire [7:0] sel_537481;
  wire [7:0] add_537484;
  wire [7:0] sel_537485;
  wire [7:0] add_537488;
  wire [7:0] sel_537489;
  wire [7:0] add_537492;
  wire [7:0] sel_537493;
  wire [7:0] add_537496;
  wire [7:0] sel_537497;
  wire [7:0] add_537500;
  wire [7:0] sel_537501;
  wire [7:0] add_537504;
  wire [7:0] sel_537505;
  wire [7:0] add_537508;
  wire [7:0] sel_537509;
  wire [7:0] add_537512;
  wire [7:0] sel_537513;
  wire [7:0] add_537516;
  wire [7:0] sel_537517;
  wire [7:0] add_537520;
  wire [7:0] sel_537521;
  wire [7:0] add_537524;
  wire [7:0] sel_537525;
  wire [7:0] add_537528;
  wire [7:0] sel_537529;
  wire [7:0] add_537532;
  wire [7:0] sel_537533;
  wire [7:0] add_537536;
  wire [7:0] sel_537537;
  wire [7:0] add_537540;
  wire [7:0] sel_537541;
  wire [7:0] add_537544;
  wire [7:0] sel_537545;
  wire [7:0] add_537548;
  wire [7:0] sel_537549;
  wire [7:0] add_537552;
  wire [7:0] sel_537553;
  wire [7:0] add_537556;
  wire [7:0] sel_537557;
  wire [7:0] add_537560;
  wire [7:0] sel_537561;
  wire [7:0] add_537564;
  wire [7:0] sel_537565;
  wire [7:0] add_537568;
  wire [7:0] sel_537569;
  wire [7:0] add_537572;
  wire [7:0] sel_537573;
  wire [7:0] add_537576;
  wire [7:0] sel_537577;
  wire [7:0] add_537580;
  wire [7:0] sel_537581;
  wire [7:0] add_537584;
  wire [7:0] sel_537585;
  wire [7:0] add_537588;
  wire [7:0] sel_537589;
  wire [7:0] add_537592;
  wire [7:0] sel_537593;
  wire [7:0] add_537596;
  wire [7:0] sel_537597;
  wire [7:0] add_537600;
  wire [7:0] sel_537601;
  wire [7:0] add_537604;
  wire [7:0] sel_537605;
  wire [7:0] add_537608;
  wire [7:0] sel_537609;
  wire [7:0] add_537612;
  wire [7:0] sel_537613;
  wire [7:0] add_537616;
  wire [7:0] sel_537617;
  wire [7:0] add_537620;
  wire [7:0] sel_537621;
  wire [7:0] add_537624;
  wire [7:0] sel_537625;
  wire [7:0] add_537628;
  wire [7:0] sel_537629;
  wire [7:0] add_537632;
  wire [7:0] sel_537633;
  wire [7:0] add_537636;
  wire [7:0] sel_537637;
  wire [7:0] add_537640;
  wire [7:0] sel_537641;
  wire [7:0] add_537644;
  wire [7:0] sel_537645;
  wire [7:0] add_537648;
  wire [7:0] sel_537649;
  wire [7:0] add_537652;
  wire [7:0] sel_537653;
  wire [7:0] add_537656;
  wire [7:0] sel_537657;
  wire [7:0] add_537660;
  wire [7:0] sel_537661;
  wire [7:0] add_537664;
  wire [7:0] sel_537665;
  wire [7:0] add_537668;
  wire [7:0] sel_537669;
  wire [7:0] add_537672;
  wire [7:0] sel_537673;
  wire [7:0] add_537676;
  wire [7:0] sel_537677;
  wire [7:0] add_537680;
  wire [7:0] sel_537681;
  wire [7:0] add_537684;
  wire [7:0] sel_537685;
  wire [7:0] add_537688;
  wire [7:0] sel_537689;
  wire [7:0] add_537692;
  wire [7:0] sel_537693;
  wire [7:0] add_537696;
  wire [7:0] sel_537697;
  wire [7:0] add_537700;
  wire [7:0] sel_537701;
  wire [7:0] add_537704;
  wire [7:0] sel_537705;
  wire [7:0] add_537708;
  wire [7:0] sel_537709;
  wire [7:0] add_537712;
  wire [7:0] sel_537713;
  wire [7:0] add_537716;
  wire [7:0] sel_537717;
  wire [7:0] add_537720;
  wire [7:0] sel_537721;
  wire [7:0] add_537724;
  wire [7:0] sel_537725;
  wire [7:0] add_537728;
  wire [7:0] sel_537729;
  wire [7:0] add_537732;
  wire [7:0] sel_537733;
  wire [7:0] add_537736;
  wire [7:0] sel_537737;
  wire [7:0] add_537740;
  wire [7:0] sel_537741;
  wire [7:0] add_537744;
  wire [7:0] sel_537745;
  wire [7:0] add_537748;
  wire [7:0] sel_537749;
  wire [7:0] add_537752;
  wire [7:0] sel_537753;
  wire [7:0] add_537756;
  wire [7:0] sel_537757;
  wire [7:0] add_537760;
  wire [7:0] sel_537761;
  wire [7:0] add_537764;
  wire [7:0] sel_537765;
  wire [7:0] add_537768;
  wire [7:0] sel_537769;
  wire [7:0] add_537773;
  wire [15:0] array_index_537774;
  wire [7:0] sel_537775;
  wire [7:0] add_537778;
  wire [7:0] sel_537779;
  wire [7:0] add_537782;
  wire [7:0] sel_537783;
  wire [7:0] add_537786;
  wire [7:0] sel_537787;
  wire [7:0] add_537790;
  wire [7:0] sel_537791;
  wire [7:0] add_537794;
  wire [7:0] sel_537795;
  wire [7:0] add_537798;
  wire [7:0] sel_537799;
  wire [7:0] add_537802;
  wire [7:0] sel_537803;
  wire [7:0] add_537806;
  wire [7:0] sel_537807;
  wire [7:0] add_537810;
  wire [7:0] sel_537811;
  wire [7:0] add_537814;
  wire [7:0] sel_537815;
  wire [7:0] add_537818;
  wire [7:0] sel_537819;
  wire [7:0] add_537822;
  wire [7:0] sel_537823;
  wire [7:0] add_537826;
  wire [7:0] sel_537827;
  wire [7:0] add_537830;
  wire [7:0] sel_537831;
  wire [7:0] add_537834;
  wire [7:0] sel_537835;
  wire [7:0] add_537838;
  wire [7:0] sel_537839;
  wire [7:0] add_537842;
  wire [7:0] sel_537843;
  wire [7:0] add_537846;
  wire [7:0] sel_537847;
  wire [7:0] add_537850;
  wire [7:0] sel_537851;
  wire [7:0] add_537854;
  wire [7:0] sel_537855;
  wire [7:0] add_537858;
  wire [7:0] sel_537859;
  wire [7:0] add_537862;
  wire [7:0] sel_537863;
  wire [7:0] add_537866;
  wire [7:0] sel_537867;
  wire [7:0] add_537870;
  wire [7:0] sel_537871;
  wire [7:0] add_537874;
  wire [7:0] sel_537875;
  wire [7:0] add_537878;
  wire [7:0] sel_537879;
  wire [7:0] add_537882;
  wire [7:0] sel_537883;
  wire [7:0] add_537886;
  wire [7:0] sel_537887;
  wire [7:0] add_537890;
  wire [7:0] sel_537891;
  wire [7:0] add_537894;
  wire [7:0] sel_537895;
  wire [7:0] add_537898;
  wire [7:0] sel_537899;
  wire [7:0] add_537902;
  wire [7:0] sel_537903;
  wire [7:0] add_537906;
  wire [7:0] sel_537907;
  wire [7:0] add_537910;
  wire [7:0] sel_537911;
  wire [7:0] add_537914;
  wire [7:0] sel_537915;
  wire [7:0] add_537918;
  wire [7:0] sel_537919;
  wire [7:0] add_537922;
  wire [7:0] sel_537923;
  wire [7:0] add_537926;
  wire [7:0] sel_537927;
  wire [7:0] add_537930;
  wire [7:0] sel_537931;
  wire [7:0] add_537934;
  wire [7:0] sel_537935;
  wire [7:0] add_537938;
  wire [7:0] sel_537939;
  wire [7:0] add_537942;
  wire [7:0] sel_537943;
  wire [7:0] add_537946;
  wire [7:0] sel_537947;
  wire [7:0] add_537950;
  wire [7:0] sel_537951;
  wire [7:0] add_537954;
  wire [7:0] sel_537955;
  wire [7:0] add_537958;
  wire [7:0] sel_537959;
  wire [7:0] add_537962;
  wire [7:0] sel_537963;
  wire [7:0] add_537966;
  wire [7:0] sel_537967;
  wire [7:0] add_537970;
  wire [7:0] sel_537971;
  wire [7:0] add_537974;
  wire [7:0] sel_537975;
  wire [7:0] add_537978;
  wire [7:0] sel_537979;
  wire [7:0] add_537982;
  wire [7:0] sel_537983;
  wire [7:0] add_537986;
  wire [7:0] sel_537987;
  wire [7:0] add_537990;
  wire [7:0] sel_537991;
  wire [7:0] add_537994;
  wire [7:0] sel_537995;
  wire [7:0] add_537998;
  wire [7:0] sel_537999;
  wire [7:0] add_538002;
  wire [7:0] sel_538003;
  wire [7:0] add_538006;
  wire [7:0] sel_538007;
  wire [7:0] add_538010;
  wire [7:0] sel_538011;
  wire [7:0] add_538014;
  wire [7:0] sel_538015;
  wire [7:0] add_538018;
  wire [7:0] sel_538019;
  wire [7:0] add_538022;
  wire [7:0] sel_538023;
  wire [7:0] add_538026;
  wire [7:0] sel_538027;
  wire [7:0] add_538030;
  wire [7:0] sel_538031;
  wire [7:0] add_538034;
  wire [7:0] sel_538035;
  wire [7:0] add_538038;
  wire [7:0] sel_538039;
  wire [7:0] add_538042;
  wire [7:0] sel_538043;
  wire [7:0] add_538046;
  wire [7:0] sel_538047;
  wire [7:0] add_538050;
  wire [7:0] sel_538051;
  wire [7:0] add_538054;
  wire [7:0] sel_538055;
  wire [7:0] add_538058;
  wire [7:0] sel_538059;
  wire [7:0] add_538062;
  wire [7:0] sel_538063;
  wire [7:0] add_538066;
  wire [7:0] sel_538067;
  wire [7:0] add_538070;
  wire [7:0] sel_538071;
  wire [7:0] add_538075;
  wire [15:0] array_index_538076;
  wire [7:0] sel_538077;
  wire [7:0] add_538080;
  wire [7:0] sel_538081;
  wire [7:0] add_538084;
  wire [7:0] sel_538085;
  wire [7:0] add_538088;
  wire [7:0] sel_538089;
  wire [7:0] add_538092;
  wire [7:0] sel_538093;
  wire [7:0] add_538096;
  wire [7:0] sel_538097;
  wire [7:0] add_538100;
  wire [7:0] sel_538101;
  wire [7:0] add_538104;
  wire [7:0] sel_538105;
  wire [7:0] add_538108;
  wire [7:0] sel_538109;
  wire [7:0] add_538112;
  wire [7:0] sel_538113;
  wire [7:0] add_538116;
  wire [7:0] sel_538117;
  wire [7:0] add_538120;
  wire [7:0] sel_538121;
  wire [7:0] add_538124;
  wire [7:0] sel_538125;
  wire [7:0] add_538128;
  wire [7:0] sel_538129;
  wire [7:0] add_538132;
  wire [7:0] sel_538133;
  wire [7:0] add_538136;
  wire [7:0] sel_538137;
  wire [7:0] add_538140;
  wire [7:0] sel_538141;
  wire [7:0] add_538144;
  wire [7:0] sel_538145;
  wire [7:0] add_538148;
  wire [7:0] sel_538149;
  wire [7:0] add_538152;
  wire [7:0] sel_538153;
  wire [7:0] add_538156;
  wire [7:0] sel_538157;
  wire [7:0] add_538160;
  wire [7:0] sel_538161;
  wire [7:0] add_538164;
  wire [7:0] sel_538165;
  wire [7:0] add_538168;
  wire [7:0] sel_538169;
  wire [7:0] add_538172;
  wire [7:0] sel_538173;
  wire [7:0] add_538176;
  wire [7:0] sel_538177;
  wire [7:0] add_538180;
  wire [7:0] sel_538181;
  wire [7:0] add_538184;
  wire [7:0] sel_538185;
  wire [7:0] add_538188;
  wire [7:0] sel_538189;
  wire [7:0] add_538192;
  wire [7:0] sel_538193;
  wire [7:0] add_538196;
  wire [7:0] sel_538197;
  wire [7:0] add_538200;
  wire [7:0] sel_538201;
  wire [7:0] add_538204;
  wire [7:0] sel_538205;
  wire [7:0] add_538208;
  wire [7:0] sel_538209;
  wire [7:0] add_538212;
  wire [7:0] sel_538213;
  wire [7:0] add_538216;
  wire [7:0] sel_538217;
  wire [7:0] add_538220;
  wire [7:0] sel_538221;
  wire [7:0] add_538224;
  wire [7:0] sel_538225;
  wire [7:0] add_538228;
  wire [7:0] sel_538229;
  wire [7:0] add_538232;
  wire [7:0] sel_538233;
  wire [7:0] add_538236;
  wire [7:0] sel_538237;
  wire [7:0] add_538240;
  wire [7:0] sel_538241;
  wire [7:0] add_538244;
  wire [7:0] sel_538245;
  wire [7:0] add_538248;
  wire [7:0] sel_538249;
  wire [7:0] add_538252;
  wire [7:0] sel_538253;
  wire [7:0] add_538256;
  wire [7:0] sel_538257;
  wire [7:0] add_538260;
  wire [7:0] sel_538261;
  wire [7:0] add_538264;
  wire [7:0] sel_538265;
  wire [7:0] add_538268;
  wire [7:0] sel_538269;
  wire [7:0] add_538272;
  wire [7:0] sel_538273;
  wire [7:0] add_538276;
  wire [7:0] sel_538277;
  wire [7:0] add_538280;
  wire [7:0] sel_538281;
  wire [7:0] add_538284;
  wire [7:0] sel_538285;
  wire [7:0] add_538288;
  wire [7:0] sel_538289;
  wire [7:0] add_538292;
  wire [7:0] sel_538293;
  wire [7:0] add_538296;
  wire [7:0] sel_538297;
  wire [7:0] add_538300;
  wire [7:0] sel_538301;
  wire [7:0] add_538304;
  wire [7:0] sel_538305;
  wire [7:0] add_538308;
  wire [7:0] sel_538309;
  wire [7:0] add_538312;
  wire [7:0] sel_538313;
  wire [7:0] add_538316;
  wire [7:0] sel_538317;
  wire [7:0] add_538320;
  wire [7:0] sel_538321;
  wire [7:0] add_538324;
  wire [7:0] sel_538325;
  wire [7:0] add_538328;
  wire [7:0] sel_538329;
  wire [7:0] add_538332;
  wire [7:0] sel_538333;
  wire [7:0] add_538336;
  wire [7:0] sel_538337;
  wire [7:0] add_538340;
  wire [7:0] sel_538341;
  wire [7:0] add_538344;
  wire [7:0] sel_538345;
  wire [7:0] add_538348;
  wire [7:0] sel_538349;
  wire [7:0] add_538352;
  wire [7:0] sel_538353;
  wire [7:0] add_538356;
  wire [7:0] sel_538357;
  wire [7:0] add_538360;
  wire [7:0] sel_538361;
  wire [7:0] add_538364;
  wire [7:0] sel_538365;
  wire [7:0] add_538368;
  wire [7:0] sel_538369;
  wire [7:0] add_538372;
  wire [7:0] sel_538373;
  wire [7:0] add_538377;
  wire [15:0] array_index_538378;
  wire [7:0] sel_538379;
  wire [7:0] add_538382;
  wire [7:0] sel_538383;
  wire [7:0] add_538386;
  wire [7:0] sel_538387;
  wire [7:0] add_538390;
  wire [7:0] sel_538391;
  wire [7:0] add_538394;
  wire [7:0] sel_538395;
  wire [7:0] add_538398;
  wire [7:0] sel_538399;
  wire [7:0] add_538402;
  wire [7:0] sel_538403;
  wire [7:0] add_538406;
  wire [7:0] sel_538407;
  wire [7:0] add_538410;
  wire [7:0] sel_538411;
  wire [7:0] add_538414;
  wire [7:0] sel_538415;
  wire [7:0] add_538418;
  wire [7:0] sel_538419;
  wire [7:0] add_538422;
  wire [7:0] sel_538423;
  wire [7:0] add_538426;
  wire [7:0] sel_538427;
  wire [7:0] add_538430;
  wire [7:0] sel_538431;
  wire [7:0] add_538434;
  wire [7:0] sel_538435;
  wire [7:0] add_538438;
  wire [7:0] sel_538439;
  wire [7:0] add_538442;
  wire [7:0] sel_538443;
  wire [7:0] add_538446;
  wire [7:0] sel_538447;
  wire [7:0] add_538450;
  wire [7:0] sel_538451;
  wire [7:0] add_538454;
  wire [7:0] sel_538455;
  wire [7:0] add_538458;
  wire [7:0] sel_538459;
  wire [7:0] add_538462;
  wire [7:0] sel_538463;
  wire [7:0] add_538466;
  wire [7:0] sel_538467;
  wire [7:0] add_538470;
  wire [7:0] sel_538471;
  wire [7:0] add_538474;
  wire [7:0] sel_538475;
  wire [7:0] add_538478;
  wire [7:0] sel_538479;
  wire [7:0] add_538482;
  wire [7:0] sel_538483;
  wire [7:0] add_538486;
  wire [7:0] sel_538487;
  wire [7:0] add_538490;
  wire [7:0] sel_538491;
  wire [7:0] add_538494;
  wire [7:0] sel_538495;
  wire [7:0] add_538498;
  wire [7:0] sel_538499;
  wire [7:0] add_538502;
  wire [7:0] sel_538503;
  wire [7:0] add_538506;
  wire [7:0] sel_538507;
  wire [7:0] add_538510;
  wire [7:0] sel_538511;
  wire [7:0] add_538514;
  wire [7:0] sel_538515;
  wire [7:0] add_538518;
  wire [7:0] sel_538519;
  wire [7:0] add_538522;
  wire [7:0] sel_538523;
  wire [7:0] add_538526;
  wire [7:0] sel_538527;
  wire [7:0] add_538530;
  wire [7:0] sel_538531;
  wire [7:0] add_538534;
  wire [7:0] sel_538535;
  wire [7:0] add_538538;
  wire [7:0] sel_538539;
  wire [7:0] add_538542;
  wire [7:0] sel_538543;
  wire [7:0] add_538546;
  wire [7:0] sel_538547;
  wire [7:0] add_538550;
  wire [7:0] sel_538551;
  wire [7:0] add_538554;
  wire [7:0] sel_538555;
  wire [7:0] add_538558;
  wire [7:0] sel_538559;
  wire [7:0] add_538562;
  wire [7:0] sel_538563;
  wire [7:0] add_538566;
  wire [7:0] sel_538567;
  wire [7:0] add_538570;
  wire [7:0] sel_538571;
  wire [7:0] add_538574;
  wire [7:0] sel_538575;
  wire [7:0] add_538578;
  wire [7:0] sel_538579;
  wire [7:0] add_538582;
  wire [7:0] sel_538583;
  wire [7:0] add_538586;
  wire [7:0] sel_538587;
  wire [7:0] add_538590;
  wire [7:0] sel_538591;
  wire [7:0] add_538594;
  wire [7:0] sel_538595;
  wire [7:0] add_538598;
  wire [7:0] sel_538599;
  wire [7:0] add_538602;
  wire [7:0] sel_538603;
  wire [7:0] add_538606;
  wire [7:0] sel_538607;
  wire [7:0] add_538610;
  wire [7:0] sel_538611;
  wire [7:0] add_538614;
  wire [7:0] sel_538615;
  wire [7:0] add_538618;
  wire [7:0] sel_538619;
  wire [7:0] add_538622;
  wire [7:0] sel_538623;
  wire [7:0] add_538626;
  wire [7:0] sel_538627;
  wire [7:0] add_538630;
  wire [7:0] sel_538631;
  wire [7:0] add_538634;
  wire [7:0] sel_538635;
  wire [7:0] add_538638;
  wire [7:0] sel_538639;
  wire [7:0] add_538642;
  wire [7:0] sel_538643;
  wire [7:0] add_538646;
  wire [7:0] sel_538647;
  wire [7:0] add_538650;
  wire [7:0] sel_538651;
  wire [7:0] add_538654;
  wire [7:0] sel_538655;
  wire [7:0] add_538658;
  wire [7:0] sel_538659;
  wire [7:0] add_538662;
  wire [7:0] sel_538663;
  wire [7:0] add_538666;
  wire [7:0] sel_538667;
  wire [7:0] add_538670;
  wire [7:0] sel_538671;
  wire [7:0] add_538674;
  wire [7:0] sel_538675;
  wire [7:0] add_538679;
  wire [15:0] array_index_538680;
  wire [7:0] sel_538681;
  wire [7:0] add_538684;
  wire [7:0] sel_538685;
  wire [7:0] add_538688;
  wire [7:0] sel_538689;
  wire [7:0] add_538692;
  wire [7:0] sel_538693;
  wire [7:0] add_538696;
  wire [7:0] sel_538697;
  wire [7:0] add_538700;
  wire [7:0] sel_538701;
  wire [7:0] add_538704;
  wire [7:0] sel_538705;
  wire [7:0] add_538708;
  wire [7:0] sel_538709;
  wire [7:0] add_538712;
  wire [7:0] sel_538713;
  wire [7:0] add_538716;
  wire [7:0] sel_538717;
  wire [7:0] add_538720;
  wire [7:0] sel_538721;
  wire [7:0] add_538724;
  wire [7:0] sel_538725;
  wire [7:0] add_538728;
  wire [7:0] sel_538729;
  wire [7:0] add_538732;
  wire [7:0] sel_538733;
  wire [7:0] add_538736;
  wire [7:0] sel_538737;
  wire [7:0] add_538740;
  wire [7:0] sel_538741;
  wire [7:0] add_538744;
  wire [7:0] sel_538745;
  wire [7:0] add_538748;
  wire [7:0] sel_538749;
  wire [7:0] add_538752;
  wire [7:0] sel_538753;
  wire [7:0] add_538756;
  wire [7:0] sel_538757;
  wire [7:0] add_538760;
  wire [7:0] sel_538761;
  wire [7:0] add_538764;
  wire [7:0] sel_538765;
  wire [7:0] add_538768;
  wire [7:0] sel_538769;
  wire [7:0] add_538772;
  wire [7:0] sel_538773;
  wire [7:0] add_538776;
  wire [7:0] sel_538777;
  wire [7:0] add_538780;
  wire [7:0] sel_538781;
  wire [7:0] add_538784;
  wire [7:0] sel_538785;
  wire [7:0] add_538788;
  wire [7:0] sel_538789;
  wire [7:0] add_538792;
  wire [7:0] sel_538793;
  wire [7:0] add_538796;
  wire [7:0] sel_538797;
  wire [7:0] add_538800;
  wire [7:0] sel_538801;
  wire [7:0] add_538804;
  wire [7:0] sel_538805;
  wire [7:0] add_538808;
  wire [7:0] sel_538809;
  wire [7:0] add_538812;
  wire [7:0] sel_538813;
  wire [7:0] add_538816;
  wire [7:0] sel_538817;
  wire [7:0] add_538820;
  wire [7:0] sel_538821;
  wire [7:0] add_538824;
  wire [7:0] sel_538825;
  wire [7:0] add_538828;
  wire [7:0] sel_538829;
  wire [7:0] add_538832;
  wire [7:0] sel_538833;
  wire [7:0] add_538836;
  wire [7:0] sel_538837;
  wire [7:0] add_538840;
  wire [7:0] sel_538841;
  wire [7:0] add_538844;
  wire [7:0] sel_538845;
  wire [7:0] add_538848;
  wire [7:0] sel_538849;
  wire [7:0] add_538852;
  wire [7:0] sel_538853;
  wire [7:0] add_538856;
  wire [7:0] sel_538857;
  wire [7:0] add_538860;
  wire [7:0] sel_538861;
  wire [7:0] add_538864;
  wire [7:0] sel_538865;
  wire [7:0] add_538868;
  wire [7:0] sel_538869;
  wire [7:0] add_538872;
  wire [7:0] sel_538873;
  wire [7:0] add_538876;
  wire [7:0] sel_538877;
  wire [7:0] add_538880;
  wire [7:0] sel_538881;
  wire [7:0] add_538884;
  wire [7:0] sel_538885;
  wire [7:0] add_538888;
  wire [7:0] sel_538889;
  wire [7:0] add_538892;
  wire [7:0] sel_538893;
  wire [7:0] add_538896;
  wire [7:0] sel_538897;
  wire [7:0] add_538900;
  wire [7:0] sel_538901;
  wire [7:0] add_538904;
  wire [7:0] sel_538905;
  wire [7:0] add_538908;
  wire [7:0] sel_538909;
  wire [7:0] add_538912;
  wire [7:0] sel_538913;
  wire [7:0] add_538916;
  wire [7:0] sel_538917;
  wire [7:0] add_538920;
  wire [7:0] sel_538921;
  wire [7:0] add_538924;
  wire [7:0] sel_538925;
  wire [7:0] add_538928;
  wire [7:0] sel_538929;
  wire [7:0] add_538932;
  wire [7:0] sel_538933;
  wire [7:0] add_538936;
  wire [7:0] sel_538937;
  wire [7:0] add_538940;
  wire [7:0] sel_538941;
  wire [7:0] add_538944;
  wire [7:0] sel_538945;
  wire [7:0] add_538948;
  wire [7:0] sel_538949;
  wire [7:0] add_538952;
  wire [7:0] sel_538953;
  wire [7:0] add_538956;
  wire [7:0] sel_538957;
  wire [7:0] add_538960;
  wire [7:0] sel_538961;
  wire [7:0] add_538964;
  wire [7:0] sel_538965;
  wire [7:0] add_538968;
  wire [7:0] sel_538969;
  wire [7:0] add_538972;
  wire [7:0] sel_538973;
  wire [7:0] add_538976;
  wire [7:0] sel_538977;
  wire [7:0] add_538981;
  wire [15:0] array_index_538982;
  wire [7:0] sel_538983;
  wire [7:0] add_538986;
  wire [7:0] sel_538987;
  wire [7:0] add_538990;
  wire [7:0] sel_538991;
  wire [7:0] add_538994;
  wire [7:0] sel_538995;
  wire [7:0] add_538998;
  wire [7:0] sel_538999;
  wire [7:0] add_539002;
  wire [7:0] sel_539003;
  wire [7:0] add_539006;
  wire [7:0] sel_539007;
  wire [7:0] add_539010;
  wire [7:0] sel_539011;
  wire [7:0] add_539014;
  wire [7:0] sel_539015;
  wire [7:0] add_539018;
  wire [7:0] sel_539019;
  wire [7:0] add_539022;
  wire [7:0] sel_539023;
  wire [7:0] add_539026;
  wire [7:0] sel_539027;
  wire [7:0] add_539030;
  wire [7:0] sel_539031;
  wire [7:0] add_539034;
  wire [7:0] sel_539035;
  wire [7:0] add_539038;
  wire [7:0] sel_539039;
  wire [7:0] add_539042;
  wire [7:0] sel_539043;
  wire [7:0] add_539046;
  wire [7:0] sel_539047;
  wire [7:0] add_539050;
  wire [7:0] sel_539051;
  wire [7:0] add_539054;
  wire [7:0] sel_539055;
  wire [7:0] add_539058;
  wire [7:0] sel_539059;
  wire [7:0] add_539062;
  wire [7:0] sel_539063;
  wire [7:0] add_539066;
  wire [7:0] sel_539067;
  wire [7:0] add_539070;
  wire [7:0] sel_539071;
  wire [7:0] add_539074;
  wire [7:0] sel_539075;
  wire [7:0] add_539078;
  wire [7:0] sel_539079;
  wire [7:0] add_539082;
  wire [7:0] sel_539083;
  wire [7:0] add_539086;
  wire [7:0] sel_539087;
  wire [7:0] add_539090;
  wire [7:0] sel_539091;
  wire [7:0] add_539094;
  wire [7:0] sel_539095;
  wire [7:0] add_539098;
  wire [7:0] sel_539099;
  wire [7:0] add_539102;
  wire [7:0] sel_539103;
  wire [7:0] add_539106;
  wire [7:0] sel_539107;
  wire [7:0] add_539110;
  wire [7:0] sel_539111;
  wire [7:0] add_539114;
  wire [7:0] sel_539115;
  wire [7:0] add_539118;
  wire [7:0] sel_539119;
  wire [7:0] add_539122;
  wire [7:0] sel_539123;
  wire [7:0] add_539126;
  wire [7:0] sel_539127;
  wire [7:0] add_539130;
  wire [7:0] sel_539131;
  wire [7:0] add_539134;
  wire [7:0] sel_539135;
  wire [7:0] add_539138;
  wire [7:0] sel_539139;
  wire [7:0] add_539142;
  wire [7:0] sel_539143;
  wire [7:0] add_539146;
  wire [7:0] sel_539147;
  wire [7:0] add_539150;
  wire [7:0] sel_539151;
  wire [7:0] add_539154;
  wire [7:0] sel_539155;
  wire [7:0] add_539158;
  wire [7:0] sel_539159;
  wire [7:0] add_539162;
  wire [7:0] sel_539163;
  wire [7:0] add_539166;
  wire [7:0] sel_539167;
  wire [7:0] add_539170;
  wire [7:0] sel_539171;
  wire [7:0] add_539174;
  wire [7:0] sel_539175;
  wire [7:0] add_539178;
  wire [7:0] sel_539179;
  wire [7:0] add_539182;
  wire [7:0] sel_539183;
  wire [7:0] add_539186;
  wire [7:0] sel_539187;
  wire [7:0] add_539190;
  wire [7:0] sel_539191;
  wire [7:0] add_539194;
  wire [7:0] sel_539195;
  wire [7:0] add_539198;
  wire [7:0] sel_539199;
  wire [7:0] add_539202;
  wire [7:0] sel_539203;
  wire [7:0] add_539206;
  wire [7:0] sel_539207;
  wire [7:0] add_539210;
  wire [7:0] sel_539211;
  wire [7:0] add_539214;
  wire [7:0] sel_539215;
  wire [7:0] add_539218;
  wire [7:0] sel_539219;
  wire [7:0] add_539222;
  wire [7:0] sel_539223;
  wire [7:0] add_539226;
  wire [7:0] sel_539227;
  wire [7:0] add_539230;
  wire [7:0] sel_539231;
  wire [7:0] add_539234;
  wire [7:0] sel_539235;
  wire [7:0] add_539238;
  wire [7:0] sel_539239;
  wire [7:0] add_539242;
  wire [7:0] sel_539243;
  wire [7:0] add_539246;
  wire [7:0] sel_539247;
  wire [7:0] add_539250;
  wire [7:0] sel_539251;
  wire [7:0] add_539254;
  wire [7:0] sel_539255;
  wire [7:0] add_539258;
  wire [7:0] sel_539259;
  wire [7:0] add_539262;
  wire [7:0] sel_539263;
  wire [7:0] add_539266;
  wire [7:0] sel_539267;
  wire [7:0] add_539270;
  wire [7:0] sel_539271;
  wire [7:0] add_539274;
  wire [7:0] sel_539275;
  wire [7:0] add_539278;
  wire [7:0] sel_539279;
  wire [7:0] add_539283;
  wire [15:0] array_index_539284;
  wire [7:0] sel_539285;
  wire [7:0] add_539288;
  wire [7:0] sel_539289;
  wire [7:0] add_539292;
  wire [7:0] sel_539293;
  wire [7:0] add_539296;
  wire [7:0] sel_539297;
  wire [7:0] add_539300;
  wire [7:0] sel_539301;
  wire [7:0] add_539304;
  wire [7:0] sel_539305;
  wire [7:0] add_539308;
  wire [7:0] sel_539309;
  wire [7:0] add_539312;
  wire [7:0] sel_539313;
  wire [7:0] add_539316;
  wire [7:0] sel_539317;
  wire [7:0] add_539320;
  wire [7:0] sel_539321;
  wire [7:0] add_539324;
  wire [7:0] sel_539325;
  wire [7:0] add_539328;
  wire [7:0] sel_539329;
  wire [7:0] add_539332;
  wire [7:0] sel_539333;
  wire [7:0] add_539336;
  wire [7:0] sel_539337;
  wire [7:0] add_539340;
  wire [7:0] sel_539341;
  wire [7:0] add_539344;
  wire [7:0] sel_539345;
  wire [7:0] add_539348;
  wire [7:0] sel_539349;
  wire [7:0] add_539352;
  wire [7:0] sel_539353;
  wire [7:0] add_539356;
  wire [7:0] sel_539357;
  wire [7:0] add_539360;
  wire [7:0] sel_539361;
  wire [7:0] add_539364;
  wire [7:0] sel_539365;
  wire [7:0] add_539368;
  wire [7:0] sel_539369;
  wire [7:0] add_539372;
  wire [7:0] sel_539373;
  wire [7:0] add_539376;
  wire [7:0] sel_539377;
  wire [7:0] add_539380;
  wire [7:0] sel_539381;
  wire [7:0] add_539384;
  wire [7:0] sel_539385;
  wire [7:0] add_539388;
  wire [7:0] sel_539389;
  wire [7:0] add_539392;
  wire [7:0] sel_539393;
  wire [7:0] add_539396;
  wire [7:0] sel_539397;
  wire [7:0] add_539400;
  wire [7:0] sel_539401;
  wire [7:0] add_539404;
  wire [7:0] sel_539405;
  wire [7:0] add_539408;
  wire [7:0] sel_539409;
  wire [7:0] add_539412;
  wire [7:0] sel_539413;
  wire [7:0] add_539416;
  wire [7:0] sel_539417;
  wire [7:0] add_539420;
  wire [7:0] sel_539421;
  wire [7:0] add_539424;
  wire [7:0] sel_539425;
  wire [7:0] add_539428;
  wire [7:0] sel_539429;
  wire [7:0] add_539432;
  wire [7:0] sel_539433;
  wire [7:0] add_539436;
  wire [7:0] sel_539437;
  wire [7:0] add_539440;
  wire [7:0] sel_539441;
  wire [7:0] add_539444;
  wire [7:0] sel_539445;
  wire [7:0] add_539448;
  wire [7:0] sel_539449;
  wire [7:0] add_539452;
  wire [7:0] sel_539453;
  wire [7:0] add_539456;
  wire [7:0] sel_539457;
  wire [7:0] add_539460;
  wire [7:0] sel_539461;
  wire [7:0] add_539464;
  wire [7:0] sel_539465;
  wire [7:0] add_539468;
  wire [7:0] sel_539469;
  wire [7:0] add_539472;
  wire [7:0] sel_539473;
  wire [7:0] add_539476;
  wire [7:0] sel_539477;
  wire [7:0] add_539480;
  wire [7:0] sel_539481;
  wire [7:0] add_539484;
  wire [7:0] sel_539485;
  wire [7:0] add_539488;
  wire [7:0] sel_539489;
  wire [7:0] add_539492;
  wire [7:0] sel_539493;
  wire [7:0] add_539496;
  wire [7:0] sel_539497;
  wire [7:0] add_539500;
  wire [7:0] sel_539501;
  wire [7:0] add_539504;
  wire [7:0] sel_539505;
  wire [7:0] add_539508;
  wire [7:0] sel_539509;
  wire [7:0] add_539512;
  wire [7:0] sel_539513;
  wire [7:0] add_539516;
  wire [7:0] sel_539517;
  wire [7:0] add_539520;
  wire [7:0] sel_539521;
  wire [7:0] add_539524;
  wire [7:0] sel_539525;
  wire [7:0] add_539528;
  wire [7:0] sel_539529;
  wire [7:0] add_539532;
  wire [7:0] sel_539533;
  wire [7:0] add_539536;
  wire [7:0] sel_539537;
  wire [7:0] add_539540;
  wire [7:0] sel_539541;
  wire [7:0] add_539544;
  wire [7:0] sel_539545;
  wire [7:0] add_539548;
  wire [7:0] sel_539549;
  wire [7:0] add_539552;
  wire [7:0] sel_539553;
  wire [7:0] add_539556;
  wire [7:0] sel_539557;
  wire [7:0] add_539560;
  wire [7:0] sel_539561;
  wire [7:0] add_539564;
  wire [7:0] sel_539565;
  wire [7:0] add_539568;
  wire [7:0] sel_539569;
  wire [7:0] add_539572;
  wire [7:0] sel_539573;
  wire [7:0] add_539576;
  wire [7:0] sel_539577;
  wire [7:0] add_539580;
  wire [7:0] sel_539581;
  wire [7:0] add_539585;
  wire [15:0] array_index_539586;
  wire [7:0] sel_539587;
  wire [7:0] add_539590;
  wire [7:0] sel_539591;
  wire [7:0] add_539594;
  wire [7:0] sel_539595;
  wire [7:0] add_539598;
  wire [7:0] sel_539599;
  wire [7:0] add_539602;
  wire [7:0] sel_539603;
  wire [7:0] add_539606;
  wire [7:0] sel_539607;
  wire [7:0] add_539610;
  wire [7:0] sel_539611;
  wire [7:0] add_539614;
  wire [7:0] sel_539615;
  wire [7:0] add_539618;
  wire [7:0] sel_539619;
  wire [7:0] add_539622;
  wire [7:0] sel_539623;
  wire [7:0] add_539626;
  wire [7:0] sel_539627;
  wire [7:0] add_539630;
  wire [7:0] sel_539631;
  wire [7:0] add_539634;
  wire [7:0] sel_539635;
  wire [7:0] add_539638;
  wire [7:0] sel_539639;
  wire [7:0] add_539642;
  wire [7:0] sel_539643;
  wire [7:0] add_539646;
  wire [7:0] sel_539647;
  wire [7:0] add_539650;
  wire [7:0] sel_539651;
  wire [7:0] add_539654;
  wire [7:0] sel_539655;
  wire [7:0] add_539658;
  wire [7:0] sel_539659;
  wire [7:0] add_539662;
  wire [7:0] sel_539663;
  wire [7:0] add_539666;
  wire [7:0] sel_539667;
  wire [7:0] add_539670;
  wire [7:0] sel_539671;
  wire [7:0] add_539674;
  wire [7:0] sel_539675;
  wire [7:0] add_539678;
  wire [7:0] sel_539679;
  wire [7:0] add_539682;
  wire [7:0] sel_539683;
  wire [7:0] add_539686;
  wire [7:0] sel_539687;
  wire [7:0] add_539690;
  wire [7:0] sel_539691;
  wire [7:0] add_539694;
  wire [7:0] sel_539695;
  wire [7:0] add_539698;
  wire [7:0] sel_539699;
  wire [7:0] add_539702;
  wire [7:0] sel_539703;
  wire [7:0] add_539706;
  wire [7:0] sel_539707;
  wire [7:0] add_539710;
  wire [7:0] sel_539711;
  wire [7:0] add_539714;
  wire [7:0] sel_539715;
  wire [7:0] add_539718;
  wire [7:0] sel_539719;
  wire [7:0] add_539722;
  wire [7:0] sel_539723;
  wire [7:0] add_539726;
  wire [7:0] sel_539727;
  wire [7:0] add_539730;
  wire [7:0] sel_539731;
  wire [7:0] add_539734;
  wire [7:0] sel_539735;
  wire [7:0] add_539738;
  wire [7:0] sel_539739;
  wire [7:0] add_539742;
  wire [7:0] sel_539743;
  wire [7:0] add_539746;
  wire [7:0] sel_539747;
  wire [7:0] add_539750;
  wire [7:0] sel_539751;
  wire [7:0] add_539754;
  wire [7:0] sel_539755;
  wire [7:0] add_539758;
  wire [7:0] sel_539759;
  wire [7:0] add_539762;
  wire [7:0] sel_539763;
  wire [7:0] add_539766;
  wire [7:0] sel_539767;
  wire [7:0] add_539770;
  wire [7:0] sel_539771;
  wire [7:0] add_539774;
  wire [7:0] sel_539775;
  wire [7:0] add_539778;
  wire [7:0] sel_539779;
  wire [7:0] add_539782;
  wire [7:0] sel_539783;
  wire [7:0] add_539786;
  wire [7:0] sel_539787;
  wire [7:0] add_539790;
  wire [7:0] sel_539791;
  wire [7:0] add_539794;
  wire [7:0] sel_539795;
  wire [7:0] add_539798;
  wire [7:0] sel_539799;
  wire [7:0] add_539802;
  wire [7:0] sel_539803;
  wire [7:0] add_539806;
  wire [7:0] sel_539807;
  wire [7:0] add_539810;
  wire [7:0] sel_539811;
  wire [7:0] add_539814;
  wire [7:0] sel_539815;
  wire [7:0] add_539818;
  wire [7:0] sel_539819;
  wire [7:0] add_539822;
  wire [7:0] sel_539823;
  wire [7:0] add_539826;
  wire [7:0] sel_539827;
  wire [7:0] add_539830;
  wire [7:0] sel_539831;
  wire [7:0] add_539834;
  wire [7:0] sel_539835;
  wire [7:0] add_539838;
  wire [7:0] sel_539839;
  wire [7:0] add_539842;
  wire [7:0] sel_539843;
  wire [7:0] add_539846;
  wire [7:0] sel_539847;
  wire [7:0] add_539850;
  wire [7:0] sel_539851;
  wire [7:0] add_539854;
  wire [7:0] sel_539855;
  wire [7:0] add_539858;
  wire [7:0] sel_539859;
  wire [7:0] add_539862;
  wire [7:0] sel_539863;
  wire [7:0] add_539866;
  wire [7:0] sel_539867;
  wire [7:0] add_539870;
  wire [7:0] sel_539871;
  wire [7:0] add_539874;
  wire [7:0] sel_539875;
  wire [7:0] add_539878;
  wire [7:0] sel_539879;
  wire [7:0] add_539882;
  wire [7:0] sel_539883;
  wire [7:0] add_539887;
  wire [15:0] array_index_539888;
  wire [7:0] sel_539889;
  wire [7:0] add_539892;
  wire [7:0] sel_539893;
  wire [7:0] add_539896;
  wire [7:0] sel_539897;
  wire [7:0] add_539900;
  wire [7:0] sel_539901;
  wire [7:0] add_539904;
  wire [7:0] sel_539905;
  wire [7:0] add_539908;
  wire [7:0] sel_539909;
  wire [7:0] add_539912;
  wire [7:0] sel_539913;
  wire [7:0] add_539916;
  wire [7:0] sel_539917;
  wire [7:0] add_539920;
  wire [7:0] sel_539921;
  wire [7:0] add_539924;
  wire [7:0] sel_539925;
  wire [7:0] add_539928;
  wire [7:0] sel_539929;
  wire [7:0] add_539932;
  wire [7:0] sel_539933;
  wire [7:0] add_539936;
  wire [7:0] sel_539937;
  wire [7:0] add_539940;
  wire [7:0] sel_539941;
  wire [7:0] add_539944;
  wire [7:0] sel_539945;
  wire [7:0] add_539948;
  wire [7:0] sel_539949;
  wire [7:0] add_539952;
  wire [7:0] sel_539953;
  wire [7:0] add_539956;
  wire [7:0] sel_539957;
  wire [7:0] add_539960;
  wire [7:0] sel_539961;
  wire [7:0] add_539964;
  wire [7:0] sel_539965;
  wire [7:0] add_539968;
  wire [7:0] sel_539969;
  wire [7:0] add_539972;
  wire [7:0] sel_539973;
  wire [7:0] add_539976;
  wire [7:0] sel_539977;
  wire [7:0] add_539980;
  wire [7:0] sel_539981;
  wire [7:0] add_539984;
  wire [7:0] sel_539985;
  wire [7:0] add_539988;
  wire [7:0] sel_539989;
  wire [7:0] add_539992;
  wire [7:0] sel_539993;
  wire [7:0] add_539996;
  wire [7:0] sel_539997;
  wire [7:0] add_540000;
  wire [7:0] sel_540001;
  wire [7:0] add_540004;
  wire [7:0] sel_540005;
  wire [7:0] add_540008;
  wire [7:0] sel_540009;
  wire [7:0] add_540012;
  wire [7:0] sel_540013;
  wire [7:0] add_540016;
  wire [7:0] sel_540017;
  wire [7:0] add_540020;
  wire [7:0] sel_540021;
  wire [7:0] add_540024;
  wire [7:0] sel_540025;
  wire [7:0] add_540028;
  wire [7:0] sel_540029;
  wire [7:0] add_540032;
  wire [7:0] sel_540033;
  wire [7:0] add_540036;
  wire [7:0] sel_540037;
  wire [7:0] add_540040;
  wire [7:0] sel_540041;
  wire [7:0] add_540044;
  wire [7:0] sel_540045;
  wire [7:0] add_540048;
  wire [7:0] sel_540049;
  wire [7:0] add_540052;
  wire [7:0] sel_540053;
  wire [7:0] add_540056;
  wire [7:0] sel_540057;
  wire [7:0] add_540060;
  wire [7:0] sel_540061;
  wire [7:0] add_540064;
  wire [7:0] sel_540065;
  wire [7:0] add_540068;
  wire [7:0] sel_540069;
  wire [7:0] add_540072;
  wire [7:0] sel_540073;
  wire [7:0] add_540076;
  wire [7:0] sel_540077;
  wire [7:0] add_540080;
  wire [7:0] sel_540081;
  wire [7:0] add_540084;
  wire [7:0] sel_540085;
  wire [7:0] add_540088;
  wire [7:0] sel_540089;
  wire [7:0] add_540092;
  wire [7:0] sel_540093;
  wire [7:0] add_540096;
  wire [7:0] sel_540097;
  wire [7:0] add_540100;
  wire [7:0] sel_540101;
  wire [7:0] add_540104;
  wire [7:0] sel_540105;
  wire [7:0] add_540108;
  wire [7:0] sel_540109;
  wire [7:0] add_540112;
  wire [7:0] sel_540113;
  wire [7:0] add_540116;
  wire [7:0] sel_540117;
  wire [7:0] add_540120;
  wire [7:0] sel_540121;
  wire [7:0] add_540124;
  wire [7:0] sel_540125;
  wire [7:0] add_540128;
  wire [7:0] sel_540129;
  wire [7:0] add_540132;
  wire [7:0] sel_540133;
  wire [7:0] add_540136;
  wire [7:0] sel_540137;
  wire [7:0] add_540140;
  wire [7:0] sel_540141;
  wire [7:0] add_540144;
  wire [7:0] sel_540145;
  wire [7:0] add_540148;
  wire [7:0] sel_540149;
  wire [7:0] add_540152;
  wire [7:0] sel_540153;
  wire [7:0] add_540156;
  wire [7:0] sel_540157;
  wire [7:0] add_540160;
  wire [7:0] sel_540161;
  wire [7:0] add_540164;
  wire [7:0] sel_540165;
  wire [7:0] add_540168;
  wire [7:0] sel_540169;
  wire [7:0] add_540172;
  wire [7:0] sel_540173;
  wire [7:0] add_540176;
  wire [7:0] sel_540177;
  wire [7:0] add_540180;
  wire [7:0] sel_540181;
  wire [7:0] add_540184;
  wire [7:0] sel_540185;
  wire [7:0] add_540189;
  wire [15:0] array_index_540190;
  wire [7:0] sel_540191;
  wire [7:0] add_540194;
  wire [7:0] sel_540195;
  wire [7:0] add_540198;
  wire [7:0] sel_540199;
  wire [7:0] add_540202;
  wire [7:0] sel_540203;
  wire [7:0] add_540206;
  wire [7:0] sel_540207;
  wire [7:0] add_540210;
  wire [7:0] sel_540211;
  wire [7:0] add_540214;
  wire [7:0] sel_540215;
  wire [7:0] add_540218;
  wire [7:0] sel_540219;
  wire [7:0] add_540222;
  wire [7:0] sel_540223;
  wire [7:0] add_540226;
  wire [7:0] sel_540227;
  wire [7:0] add_540230;
  wire [7:0] sel_540231;
  wire [7:0] add_540234;
  wire [7:0] sel_540235;
  wire [7:0] add_540238;
  wire [7:0] sel_540239;
  wire [7:0] add_540242;
  wire [7:0] sel_540243;
  wire [7:0] add_540246;
  wire [7:0] sel_540247;
  wire [7:0] add_540250;
  wire [7:0] sel_540251;
  wire [7:0] add_540254;
  wire [7:0] sel_540255;
  wire [7:0] add_540258;
  wire [7:0] sel_540259;
  wire [7:0] add_540262;
  wire [7:0] sel_540263;
  wire [7:0] add_540266;
  wire [7:0] sel_540267;
  wire [7:0] add_540270;
  wire [7:0] sel_540271;
  wire [7:0] add_540274;
  wire [7:0] sel_540275;
  wire [7:0] add_540278;
  wire [7:0] sel_540279;
  wire [7:0] add_540282;
  wire [7:0] sel_540283;
  wire [7:0] add_540286;
  wire [7:0] sel_540287;
  wire [7:0] add_540290;
  wire [7:0] sel_540291;
  wire [7:0] add_540294;
  wire [7:0] sel_540295;
  wire [7:0] add_540298;
  wire [7:0] sel_540299;
  wire [7:0] add_540302;
  wire [7:0] sel_540303;
  wire [7:0] add_540306;
  wire [7:0] sel_540307;
  wire [7:0] add_540310;
  wire [7:0] sel_540311;
  wire [7:0] add_540314;
  wire [7:0] sel_540315;
  wire [7:0] add_540318;
  wire [7:0] sel_540319;
  wire [7:0] add_540322;
  wire [7:0] sel_540323;
  wire [7:0] add_540326;
  wire [7:0] sel_540327;
  wire [7:0] add_540330;
  wire [7:0] sel_540331;
  wire [7:0] add_540334;
  wire [7:0] sel_540335;
  wire [7:0] add_540338;
  wire [7:0] sel_540339;
  wire [7:0] add_540342;
  wire [7:0] sel_540343;
  wire [7:0] add_540346;
  wire [7:0] sel_540347;
  wire [7:0] add_540350;
  wire [7:0] sel_540351;
  wire [7:0] add_540354;
  wire [7:0] sel_540355;
  wire [7:0] add_540358;
  wire [7:0] sel_540359;
  wire [7:0] add_540362;
  wire [7:0] sel_540363;
  wire [7:0] add_540366;
  wire [7:0] sel_540367;
  wire [7:0] add_540370;
  wire [7:0] sel_540371;
  wire [7:0] add_540374;
  wire [7:0] sel_540375;
  wire [7:0] add_540378;
  wire [7:0] sel_540379;
  wire [7:0] add_540382;
  wire [7:0] sel_540383;
  wire [7:0] add_540386;
  wire [7:0] sel_540387;
  wire [7:0] add_540390;
  wire [7:0] sel_540391;
  wire [7:0] add_540394;
  wire [7:0] sel_540395;
  wire [7:0] add_540398;
  wire [7:0] sel_540399;
  wire [7:0] add_540402;
  wire [7:0] sel_540403;
  wire [7:0] add_540406;
  wire [7:0] sel_540407;
  wire [7:0] add_540410;
  wire [7:0] sel_540411;
  wire [7:0] add_540414;
  wire [7:0] sel_540415;
  wire [7:0] add_540418;
  wire [7:0] sel_540419;
  wire [7:0] add_540422;
  wire [7:0] sel_540423;
  wire [7:0] add_540426;
  wire [7:0] sel_540427;
  wire [7:0] add_540430;
  wire [7:0] sel_540431;
  wire [7:0] add_540434;
  wire [7:0] sel_540435;
  wire [7:0] add_540438;
  wire [7:0] sel_540439;
  wire [7:0] add_540442;
  wire [7:0] sel_540443;
  wire [7:0] add_540446;
  wire [7:0] sel_540447;
  wire [7:0] add_540450;
  wire [7:0] sel_540451;
  wire [7:0] add_540454;
  wire [7:0] sel_540455;
  wire [7:0] add_540458;
  wire [7:0] sel_540459;
  wire [7:0] add_540462;
  wire [7:0] sel_540463;
  wire [7:0] add_540466;
  wire [7:0] sel_540467;
  wire [7:0] add_540470;
  wire [7:0] sel_540471;
  wire [7:0] add_540474;
  wire [7:0] sel_540475;
  wire [7:0] add_540478;
  wire [7:0] sel_540479;
  wire [7:0] add_540482;
  wire [7:0] sel_540483;
  wire [7:0] add_540486;
  wire [7:0] sel_540487;
  wire [7:0] add_540491;
  wire [15:0] array_index_540492;
  wire [7:0] sel_540493;
  wire [7:0] add_540496;
  wire [7:0] sel_540497;
  wire [7:0] add_540500;
  wire [7:0] sel_540501;
  wire [7:0] add_540504;
  wire [7:0] sel_540505;
  wire [7:0] add_540508;
  wire [7:0] sel_540509;
  wire [7:0] add_540512;
  wire [7:0] sel_540513;
  wire [7:0] add_540516;
  wire [7:0] sel_540517;
  wire [7:0] add_540520;
  wire [7:0] sel_540521;
  wire [7:0] add_540524;
  wire [7:0] sel_540525;
  wire [7:0] add_540528;
  wire [7:0] sel_540529;
  wire [7:0] add_540532;
  wire [7:0] sel_540533;
  wire [7:0] add_540536;
  wire [7:0] sel_540537;
  wire [7:0] add_540540;
  wire [7:0] sel_540541;
  wire [7:0] add_540544;
  wire [7:0] sel_540545;
  wire [7:0] add_540548;
  wire [7:0] sel_540549;
  wire [7:0] add_540552;
  wire [7:0] sel_540553;
  wire [7:0] add_540556;
  wire [7:0] sel_540557;
  wire [7:0] add_540560;
  wire [7:0] sel_540561;
  wire [7:0] add_540564;
  wire [7:0] sel_540565;
  wire [7:0] add_540568;
  wire [7:0] sel_540569;
  wire [7:0] add_540572;
  wire [7:0] sel_540573;
  wire [7:0] add_540576;
  wire [7:0] sel_540577;
  wire [7:0] add_540580;
  wire [7:0] sel_540581;
  wire [7:0] add_540584;
  wire [7:0] sel_540585;
  wire [7:0] add_540588;
  wire [7:0] sel_540589;
  wire [7:0] add_540592;
  wire [7:0] sel_540593;
  wire [7:0] add_540596;
  wire [7:0] sel_540597;
  wire [7:0] add_540600;
  wire [7:0] sel_540601;
  wire [7:0] add_540604;
  wire [7:0] sel_540605;
  wire [7:0] add_540608;
  wire [7:0] sel_540609;
  wire [7:0] add_540612;
  wire [7:0] sel_540613;
  wire [7:0] add_540616;
  wire [7:0] sel_540617;
  wire [7:0] add_540620;
  wire [7:0] sel_540621;
  wire [7:0] add_540624;
  wire [7:0] sel_540625;
  wire [7:0] add_540628;
  wire [7:0] sel_540629;
  wire [7:0] add_540632;
  wire [7:0] sel_540633;
  wire [7:0] add_540636;
  wire [7:0] sel_540637;
  wire [7:0] add_540640;
  wire [7:0] sel_540641;
  wire [7:0] add_540644;
  wire [7:0] sel_540645;
  wire [7:0] add_540648;
  wire [7:0] sel_540649;
  wire [7:0] add_540652;
  wire [7:0] sel_540653;
  wire [7:0] add_540656;
  wire [7:0] sel_540657;
  wire [7:0] add_540660;
  wire [7:0] sel_540661;
  wire [7:0] add_540664;
  wire [7:0] sel_540665;
  wire [7:0] add_540668;
  wire [7:0] sel_540669;
  wire [7:0] add_540672;
  wire [7:0] sel_540673;
  wire [7:0] add_540676;
  wire [7:0] sel_540677;
  wire [7:0] add_540680;
  wire [7:0] sel_540681;
  wire [7:0] add_540684;
  wire [7:0] sel_540685;
  wire [7:0] add_540688;
  wire [7:0] sel_540689;
  wire [7:0] add_540692;
  wire [7:0] sel_540693;
  wire [7:0] add_540696;
  wire [7:0] sel_540697;
  wire [7:0] add_540700;
  wire [7:0] sel_540701;
  wire [7:0] add_540704;
  wire [7:0] sel_540705;
  wire [7:0] add_540708;
  wire [7:0] sel_540709;
  wire [7:0] add_540712;
  wire [7:0] sel_540713;
  wire [7:0] add_540716;
  wire [7:0] sel_540717;
  wire [7:0] add_540720;
  wire [7:0] sel_540721;
  wire [7:0] add_540724;
  wire [7:0] sel_540725;
  wire [7:0] add_540728;
  wire [7:0] sel_540729;
  wire [7:0] add_540732;
  wire [7:0] sel_540733;
  wire [7:0] add_540736;
  wire [7:0] sel_540737;
  wire [7:0] add_540740;
  wire [7:0] sel_540741;
  wire [7:0] add_540744;
  wire [7:0] sel_540745;
  wire [7:0] add_540748;
  wire [7:0] sel_540749;
  wire [7:0] add_540752;
  wire [7:0] sel_540753;
  wire [7:0] add_540756;
  wire [7:0] sel_540757;
  wire [7:0] add_540760;
  wire [7:0] sel_540761;
  wire [7:0] add_540764;
  wire [7:0] sel_540765;
  wire [7:0] add_540768;
  wire [7:0] sel_540769;
  wire [7:0] add_540772;
  wire [7:0] sel_540773;
  wire [7:0] add_540776;
  wire [7:0] sel_540777;
  wire [7:0] add_540780;
  wire [7:0] sel_540781;
  wire [7:0] add_540784;
  wire [7:0] sel_540785;
  wire [7:0] add_540788;
  wire [7:0] sel_540789;
  wire [7:0] add_540793;
  wire [15:0] array_index_540794;
  wire [7:0] sel_540795;
  wire [7:0] add_540798;
  wire [7:0] sel_540799;
  wire [7:0] add_540802;
  wire [7:0] sel_540803;
  wire [7:0] add_540806;
  wire [7:0] sel_540807;
  wire [7:0] add_540810;
  wire [7:0] sel_540811;
  wire [7:0] add_540814;
  wire [7:0] sel_540815;
  wire [7:0] add_540818;
  wire [7:0] sel_540819;
  wire [7:0] add_540822;
  wire [7:0] sel_540823;
  wire [7:0] add_540826;
  wire [7:0] sel_540827;
  wire [7:0] add_540830;
  wire [7:0] sel_540831;
  wire [7:0] add_540834;
  wire [7:0] sel_540835;
  wire [7:0] add_540838;
  wire [7:0] sel_540839;
  wire [7:0] add_540842;
  wire [7:0] sel_540843;
  wire [7:0] add_540846;
  wire [7:0] sel_540847;
  wire [7:0] add_540850;
  wire [7:0] sel_540851;
  wire [7:0] add_540854;
  wire [7:0] sel_540855;
  wire [7:0] add_540858;
  wire [7:0] sel_540859;
  wire [7:0] add_540862;
  wire [7:0] sel_540863;
  wire [7:0] add_540866;
  wire [7:0] sel_540867;
  wire [7:0] add_540870;
  wire [7:0] sel_540871;
  wire [7:0] add_540874;
  wire [7:0] sel_540875;
  wire [7:0] add_540878;
  wire [7:0] sel_540879;
  wire [7:0] add_540882;
  wire [7:0] sel_540883;
  wire [7:0] add_540886;
  wire [7:0] sel_540887;
  wire [7:0] add_540890;
  wire [7:0] sel_540891;
  wire [7:0] add_540894;
  wire [7:0] sel_540895;
  wire [7:0] add_540898;
  wire [7:0] sel_540899;
  wire [7:0] add_540902;
  wire [7:0] sel_540903;
  wire [7:0] add_540906;
  wire [7:0] sel_540907;
  wire [7:0] add_540910;
  wire [7:0] sel_540911;
  wire [7:0] add_540914;
  wire [7:0] sel_540915;
  wire [7:0] add_540918;
  wire [7:0] sel_540919;
  wire [7:0] add_540922;
  wire [7:0] sel_540923;
  wire [7:0] add_540926;
  wire [7:0] sel_540927;
  wire [7:0] add_540930;
  wire [7:0] sel_540931;
  wire [7:0] add_540934;
  wire [7:0] sel_540935;
  wire [7:0] add_540938;
  wire [7:0] sel_540939;
  wire [7:0] add_540942;
  wire [7:0] sel_540943;
  wire [7:0] add_540946;
  wire [7:0] sel_540947;
  wire [7:0] add_540950;
  wire [7:0] sel_540951;
  wire [7:0] add_540954;
  wire [7:0] sel_540955;
  wire [7:0] add_540958;
  wire [7:0] sel_540959;
  wire [7:0] add_540962;
  wire [7:0] sel_540963;
  wire [7:0] add_540966;
  wire [7:0] sel_540967;
  wire [7:0] add_540970;
  wire [7:0] sel_540971;
  wire [7:0] add_540974;
  wire [7:0] sel_540975;
  wire [7:0] add_540978;
  wire [7:0] sel_540979;
  wire [7:0] add_540982;
  wire [7:0] sel_540983;
  wire [7:0] add_540986;
  wire [7:0] sel_540987;
  wire [7:0] add_540990;
  wire [7:0] sel_540991;
  wire [7:0] add_540994;
  wire [7:0] sel_540995;
  wire [7:0] add_540998;
  wire [7:0] sel_540999;
  wire [7:0] add_541002;
  wire [7:0] sel_541003;
  wire [7:0] add_541006;
  wire [7:0] sel_541007;
  wire [7:0] add_541010;
  wire [7:0] sel_541011;
  wire [7:0] add_541014;
  wire [7:0] sel_541015;
  wire [7:0] add_541018;
  wire [7:0] sel_541019;
  wire [7:0] add_541022;
  wire [7:0] sel_541023;
  wire [7:0] add_541026;
  wire [7:0] sel_541027;
  wire [7:0] add_541030;
  wire [7:0] sel_541031;
  wire [7:0] add_541034;
  wire [7:0] sel_541035;
  wire [7:0] add_541038;
  wire [7:0] sel_541039;
  wire [7:0] add_541042;
  wire [7:0] sel_541043;
  wire [7:0] add_541046;
  wire [7:0] sel_541047;
  wire [7:0] add_541050;
  wire [7:0] sel_541051;
  wire [7:0] add_541054;
  wire [7:0] sel_541055;
  wire [7:0] add_541058;
  wire [7:0] sel_541059;
  wire [7:0] add_541062;
  wire [7:0] sel_541063;
  wire [7:0] add_541066;
  wire [7:0] sel_541067;
  wire [7:0] add_541070;
  wire [7:0] sel_541071;
  wire [7:0] add_541074;
  wire [7:0] sel_541075;
  wire [7:0] add_541078;
  wire [7:0] sel_541079;
  wire [7:0] add_541082;
  wire [7:0] sel_541083;
  wire [7:0] add_541086;
  wire [7:0] sel_541087;
  wire [7:0] add_541090;
  wire [7:0] sel_541091;
  wire [7:0] add_541095;
  wire [15:0] array_index_541096;
  wire [7:0] sel_541097;
  wire [7:0] add_541100;
  wire [7:0] sel_541101;
  wire [7:0] add_541104;
  wire [7:0] sel_541105;
  wire [7:0] add_541108;
  wire [7:0] sel_541109;
  wire [7:0] add_541112;
  wire [7:0] sel_541113;
  wire [7:0] add_541116;
  wire [7:0] sel_541117;
  wire [7:0] add_541120;
  wire [7:0] sel_541121;
  wire [7:0] add_541124;
  wire [7:0] sel_541125;
  wire [7:0] add_541128;
  wire [7:0] sel_541129;
  wire [7:0] add_541132;
  wire [7:0] sel_541133;
  wire [7:0] add_541136;
  wire [7:0] sel_541137;
  wire [7:0] add_541140;
  wire [7:0] sel_541141;
  wire [7:0] add_541144;
  wire [7:0] sel_541145;
  wire [7:0] add_541148;
  wire [7:0] sel_541149;
  wire [7:0] add_541152;
  wire [7:0] sel_541153;
  wire [7:0] add_541156;
  wire [7:0] sel_541157;
  wire [7:0] add_541160;
  wire [7:0] sel_541161;
  wire [7:0] add_541164;
  wire [7:0] sel_541165;
  wire [7:0] add_541168;
  wire [7:0] sel_541169;
  wire [7:0] add_541172;
  wire [7:0] sel_541173;
  wire [7:0] add_541176;
  wire [7:0] sel_541177;
  wire [7:0] add_541180;
  wire [7:0] sel_541181;
  wire [7:0] add_541184;
  wire [7:0] sel_541185;
  wire [7:0] add_541188;
  wire [7:0] sel_541189;
  wire [7:0] add_541192;
  wire [7:0] sel_541193;
  wire [7:0] add_541196;
  wire [7:0] sel_541197;
  wire [7:0] add_541200;
  wire [7:0] sel_541201;
  wire [7:0] add_541204;
  wire [7:0] sel_541205;
  wire [7:0] add_541208;
  wire [7:0] sel_541209;
  wire [7:0] add_541212;
  wire [7:0] sel_541213;
  wire [7:0] add_541216;
  wire [7:0] sel_541217;
  wire [7:0] add_541220;
  wire [7:0] sel_541221;
  wire [7:0] add_541224;
  wire [7:0] sel_541225;
  wire [7:0] add_541228;
  wire [7:0] sel_541229;
  wire [7:0] add_541232;
  wire [7:0] sel_541233;
  wire [7:0] add_541236;
  wire [7:0] sel_541237;
  wire [7:0] add_541240;
  wire [7:0] sel_541241;
  wire [7:0] add_541244;
  wire [7:0] sel_541245;
  wire [7:0] add_541248;
  wire [7:0] sel_541249;
  wire [7:0] add_541252;
  wire [7:0] sel_541253;
  wire [7:0] add_541256;
  wire [7:0] sel_541257;
  wire [7:0] add_541260;
  wire [7:0] sel_541261;
  wire [7:0] add_541264;
  wire [7:0] sel_541265;
  wire [7:0] add_541268;
  wire [7:0] sel_541269;
  wire [7:0] add_541272;
  wire [7:0] sel_541273;
  wire [7:0] add_541276;
  wire [7:0] sel_541277;
  wire [7:0] add_541280;
  wire [7:0] sel_541281;
  wire [7:0] add_541284;
  wire [7:0] sel_541285;
  wire [7:0] add_541288;
  wire [7:0] sel_541289;
  wire [7:0] add_541292;
  wire [7:0] sel_541293;
  wire [7:0] add_541296;
  wire [7:0] sel_541297;
  wire [7:0] add_541300;
  wire [7:0] sel_541301;
  wire [7:0] add_541304;
  wire [7:0] sel_541305;
  wire [7:0] add_541308;
  wire [7:0] sel_541309;
  wire [7:0] add_541312;
  wire [7:0] sel_541313;
  wire [7:0] add_541316;
  wire [7:0] sel_541317;
  wire [7:0] add_541320;
  wire [7:0] sel_541321;
  wire [7:0] add_541324;
  wire [7:0] sel_541325;
  wire [7:0] add_541328;
  wire [7:0] sel_541329;
  wire [7:0] add_541332;
  wire [7:0] sel_541333;
  wire [7:0] add_541336;
  wire [7:0] sel_541337;
  wire [7:0] add_541340;
  wire [7:0] sel_541341;
  wire [7:0] add_541344;
  wire [7:0] sel_541345;
  wire [7:0] add_541348;
  wire [7:0] sel_541349;
  wire [7:0] add_541352;
  wire [7:0] sel_541353;
  wire [7:0] add_541356;
  wire [7:0] sel_541357;
  wire [7:0] add_541360;
  wire [7:0] sel_541361;
  wire [7:0] add_541364;
  wire [7:0] sel_541365;
  wire [7:0] add_541368;
  wire [7:0] sel_541369;
  wire [7:0] add_541372;
  wire [7:0] sel_541373;
  wire [7:0] add_541376;
  wire [7:0] sel_541377;
  wire [7:0] add_541380;
  wire [7:0] sel_541381;
  wire [7:0] add_541384;
  wire [7:0] sel_541385;
  wire [7:0] add_541388;
  wire [7:0] sel_541389;
  wire [7:0] add_541392;
  wire [7:0] sel_541393;
  wire [7:0] add_541397;
  wire [15:0] array_index_541398;
  wire [7:0] sel_541399;
  wire [7:0] add_541402;
  wire [7:0] sel_541403;
  wire [7:0] add_541406;
  wire [7:0] sel_541407;
  wire [7:0] add_541410;
  wire [7:0] sel_541411;
  wire [7:0] add_541414;
  wire [7:0] sel_541415;
  wire [7:0] add_541418;
  wire [7:0] sel_541419;
  wire [7:0] add_541422;
  wire [7:0] sel_541423;
  wire [7:0] add_541426;
  wire [7:0] sel_541427;
  wire [7:0] add_541430;
  wire [7:0] sel_541431;
  wire [7:0] add_541434;
  wire [7:0] sel_541435;
  wire [7:0] add_541438;
  wire [7:0] sel_541439;
  wire [7:0] add_541442;
  wire [7:0] sel_541443;
  wire [7:0] add_541446;
  wire [7:0] sel_541447;
  wire [7:0] add_541450;
  wire [7:0] sel_541451;
  wire [7:0] add_541454;
  wire [7:0] sel_541455;
  wire [7:0] add_541458;
  wire [7:0] sel_541459;
  wire [7:0] add_541462;
  wire [7:0] sel_541463;
  wire [7:0] add_541466;
  wire [7:0] sel_541467;
  wire [7:0] add_541470;
  wire [7:0] sel_541471;
  wire [7:0] add_541474;
  wire [7:0] sel_541475;
  wire [7:0] add_541478;
  wire [7:0] sel_541479;
  wire [7:0] add_541482;
  wire [7:0] sel_541483;
  wire [7:0] add_541486;
  wire [7:0] sel_541487;
  wire [7:0] add_541490;
  wire [7:0] sel_541491;
  wire [7:0] add_541494;
  wire [7:0] sel_541495;
  wire [7:0] add_541498;
  wire [7:0] sel_541499;
  wire [7:0] add_541502;
  wire [7:0] sel_541503;
  wire [7:0] add_541506;
  wire [7:0] sel_541507;
  wire [7:0] add_541510;
  wire [7:0] sel_541511;
  wire [7:0] add_541514;
  wire [7:0] sel_541515;
  wire [7:0] add_541518;
  wire [7:0] sel_541519;
  wire [7:0] add_541522;
  wire [7:0] sel_541523;
  wire [7:0] add_541526;
  wire [7:0] sel_541527;
  wire [7:0] add_541530;
  wire [7:0] sel_541531;
  wire [7:0] add_541534;
  wire [7:0] sel_541535;
  wire [7:0] add_541538;
  wire [7:0] sel_541539;
  wire [7:0] add_541542;
  wire [7:0] sel_541543;
  wire [7:0] add_541546;
  wire [7:0] sel_541547;
  wire [7:0] add_541550;
  wire [7:0] sel_541551;
  wire [7:0] add_541554;
  wire [7:0] sel_541555;
  wire [7:0] add_541558;
  wire [7:0] sel_541559;
  wire [7:0] add_541562;
  wire [7:0] sel_541563;
  wire [7:0] add_541566;
  wire [7:0] sel_541567;
  wire [7:0] add_541570;
  wire [7:0] sel_541571;
  wire [7:0] add_541574;
  wire [7:0] sel_541575;
  wire [7:0] add_541578;
  wire [7:0] sel_541579;
  wire [7:0] add_541582;
  wire [7:0] sel_541583;
  wire [7:0] add_541586;
  wire [7:0] sel_541587;
  wire [7:0] add_541590;
  wire [7:0] sel_541591;
  wire [7:0] add_541594;
  wire [7:0] sel_541595;
  wire [7:0] add_541598;
  wire [7:0] sel_541599;
  wire [7:0] add_541602;
  wire [7:0] sel_541603;
  wire [7:0] add_541606;
  wire [7:0] sel_541607;
  wire [7:0] add_541610;
  wire [7:0] sel_541611;
  wire [7:0] add_541614;
  wire [7:0] sel_541615;
  wire [7:0] add_541618;
  wire [7:0] sel_541619;
  wire [7:0] add_541622;
  wire [7:0] sel_541623;
  wire [7:0] add_541626;
  wire [7:0] sel_541627;
  wire [7:0] add_541630;
  wire [7:0] sel_541631;
  wire [7:0] add_541634;
  wire [7:0] sel_541635;
  wire [7:0] add_541638;
  wire [7:0] sel_541639;
  wire [7:0] add_541642;
  wire [7:0] sel_541643;
  wire [7:0] add_541646;
  wire [7:0] sel_541647;
  wire [7:0] add_541650;
  wire [7:0] sel_541651;
  wire [7:0] add_541654;
  wire [7:0] sel_541655;
  wire [7:0] add_541658;
  wire [7:0] sel_541659;
  wire [7:0] add_541662;
  wire [7:0] sel_541663;
  wire [7:0] add_541666;
  wire [7:0] sel_541667;
  wire [7:0] add_541670;
  wire [7:0] sel_541671;
  wire [7:0] add_541674;
  wire [7:0] sel_541675;
  wire [7:0] add_541678;
  wire [7:0] sel_541679;
  wire [7:0] add_541682;
  wire [7:0] sel_541683;
  wire [7:0] add_541686;
  wire [7:0] sel_541687;
  wire [7:0] add_541690;
  wire [7:0] sel_541691;
  wire [7:0] add_541694;
  wire [7:0] sel_541695;
  wire [7:0] add_541699;
  wire [15:0] array_index_541700;
  wire [7:0] sel_541701;
  wire [7:0] add_541704;
  wire [7:0] sel_541705;
  wire [7:0] add_541708;
  wire [7:0] sel_541709;
  wire [7:0] add_541712;
  wire [7:0] sel_541713;
  wire [7:0] add_541716;
  wire [7:0] sel_541717;
  wire [7:0] add_541720;
  wire [7:0] sel_541721;
  wire [7:0] add_541724;
  wire [7:0] sel_541725;
  wire [7:0] add_541728;
  wire [7:0] sel_541729;
  wire [7:0] add_541732;
  wire [7:0] sel_541733;
  wire [7:0] add_541736;
  wire [7:0] sel_541737;
  wire [7:0] add_541740;
  wire [7:0] sel_541741;
  wire [7:0] add_541744;
  wire [7:0] sel_541745;
  wire [7:0] add_541748;
  wire [7:0] sel_541749;
  wire [7:0] add_541752;
  wire [7:0] sel_541753;
  wire [7:0] add_541756;
  wire [7:0] sel_541757;
  wire [7:0] add_541760;
  wire [7:0] sel_541761;
  wire [7:0] add_541764;
  wire [7:0] sel_541765;
  wire [7:0] add_541768;
  wire [7:0] sel_541769;
  wire [7:0] add_541772;
  wire [7:0] sel_541773;
  wire [7:0] add_541776;
  wire [7:0] sel_541777;
  wire [7:0] add_541780;
  wire [7:0] sel_541781;
  wire [7:0] add_541784;
  wire [7:0] sel_541785;
  wire [7:0] add_541788;
  wire [7:0] sel_541789;
  wire [7:0] add_541792;
  wire [7:0] sel_541793;
  wire [7:0] add_541796;
  wire [7:0] sel_541797;
  wire [7:0] add_541800;
  wire [7:0] sel_541801;
  wire [7:0] add_541804;
  wire [7:0] sel_541805;
  wire [7:0] add_541808;
  wire [7:0] sel_541809;
  wire [7:0] add_541812;
  wire [7:0] sel_541813;
  wire [7:0] add_541816;
  wire [7:0] sel_541817;
  wire [7:0] add_541820;
  wire [7:0] sel_541821;
  wire [7:0] add_541824;
  wire [7:0] sel_541825;
  wire [7:0] add_541828;
  wire [7:0] sel_541829;
  wire [7:0] add_541832;
  wire [7:0] sel_541833;
  wire [7:0] add_541836;
  wire [7:0] sel_541837;
  wire [7:0] add_541840;
  wire [7:0] sel_541841;
  wire [7:0] add_541844;
  wire [7:0] sel_541845;
  wire [7:0] add_541848;
  wire [7:0] sel_541849;
  wire [7:0] add_541852;
  wire [7:0] sel_541853;
  wire [7:0] add_541856;
  wire [7:0] sel_541857;
  wire [7:0] add_541860;
  wire [7:0] sel_541861;
  wire [7:0] add_541864;
  wire [7:0] sel_541865;
  wire [7:0] add_541868;
  wire [7:0] sel_541869;
  wire [7:0] add_541872;
  wire [7:0] sel_541873;
  wire [7:0] add_541876;
  wire [7:0] sel_541877;
  wire [7:0] add_541880;
  wire [7:0] sel_541881;
  wire [7:0] add_541884;
  wire [7:0] sel_541885;
  wire [7:0] add_541888;
  wire [7:0] sel_541889;
  wire [7:0] add_541892;
  wire [7:0] sel_541893;
  wire [7:0] add_541896;
  wire [7:0] sel_541897;
  wire [7:0] add_541900;
  wire [7:0] sel_541901;
  wire [7:0] add_541904;
  wire [7:0] sel_541905;
  wire [7:0] add_541908;
  wire [7:0] sel_541909;
  wire [7:0] add_541912;
  wire [7:0] sel_541913;
  wire [7:0] add_541916;
  wire [7:0] sel_541917;
  wire [7:0] add_541920;
  wire [7:0] sel_541921;
  wire [7:0] add_541924;
  wire [7:0] sel_541925;
  wire [7:0] add_541928;
  wire [7:0] sel_541929;
  wire [7:0] add_541932;
  wire [7:0] sel_541933;
  wire [7:0] add_541936;
  wire [7:0] sel_541937;
  wire [7:0] add_541940;
  wire [7:0] sel_541941;
  wire [7:0] add_541944;
  wire [7:0] sel_541945;
  wire [7:0] add_541948;
  wire [7:0] sel_541949;
  wire [7:0] add_541952;
  wire [7:0] sel_541953;
  wire [7:0] add_541956;
  wire [7:0] sel_541957;
  wire [7:0] add_541960;
  wire [7:0] sel_541961;
  wire [7:0] add_541964;
  wire [7:0] sel_541965;
  wire [7:0] add_541968;
  wire [7:0] sel_541969;
  wire [7:0] add_541972;
  wire [7:0] sel_541973;
  wire [7:0] add_541976;
  wire [7:0] sel_541977;
  wire [7:0] add_541980;
  wire [7:0] sel_541981;
  wire [7:0] add_541984;
  wire [7:0] sel_541985;
  wire [7:0] add_541988;
  wire [7:0] sel_541989;
  wire [7:0] add_541992;
  wire [7:0] sel_541993;
  wire [7:0] add_541996;
  wire [7:0] sel_541997;
  wire [7:0] add_542001;
  wire [15:0] array_index_542002;
  wire [7:0] sel_542003;
  wire [7:0] add_542006;
  wire [7:0] sel_542007;
  wire [7:0] add_542010;
  wire [7:0] sel_542011;
  wire [7:0] add_542014;
  wire [7:0] sel_542015;
  wire [7:0] add_542018;
  wire [7:0] sel_542019;
  wire [7:0] add_542022;
  wire [7:0] sel_542023;
  wire [7:0] add_542026;
  wire [7:0] sel_542027;
  wire [7:0] add_542030;
  wire [7:0] sel_542031;
  wire [7:0] add_542034;
  wire [7:0] sel_542035;
  wire [7:0] add_542038;
  wire [7:0] sel_542039;
  wire [7:0] add_542042;
  wire [7:0] sel_542043;
  wire [7:0] add_542046;
  wire [7:0] sel_542047;
  wire [7:0] add_542050;
  wire [7:0] sel_542051;
  wire [7:0] add_542054;
  wire [7:0] sel_542055;
  wire [7:0] add_542058;
  wire [7:0] sel_542059;
  wire [7:0] add_542062;
  wire [7:0] sel_542063;
  wire [7:0] add_542066;
  wire [7:0] sel_542067;
  wire [7:0] add_542070;
  wire [7:0] sel_542071;
  wire [7:0] add_542074;
  wire [7:0] sel_542075;
  wire [7:0] add_542078;
  wire [7:0] sel_542079;
  wire [7:0] add_542082;
  wire [7:0] sel_542083;
  wire [7:0] add_542086;
  wire [7:0] sel_542087;
  wire [7:0] add_542090;
  wire [7:0] sel_542091;
  wire [7:0] add_542094;
  wire [7:0] sel_542095;
  wire [7:0] add_542098;
  wire [7:0] sel_542099;
  wire [7:0] add_542102;
  wire [7:0] sel_542103;
  wire [7:0] add_542106;
  wire [7:0] sel_542107;
  wire [7:0] add_542110;
  wire [7:0] sel_542111;
  wire [7:0] add_542114;
  wire [7:0] sel_542115;
  wire [7:0] add_542118;
  wire [7:0] sel_542119;
  wire [7:0] add_542122;
  wire [7:0] sel_542123;
  wire [7:0] add_542126;
  wire [7:0] sel_542127;
  wire [7:0] add_542130;
  wire [7:0] sel_542131;
  wire [7:0] add_542134;
  wire [7:0] sel_542135;
  wire [7:0] add_542138;
  wire [7:0] sel_542139;
  wire [7:0] add_542142;
  wire [7:0] sel_542143;
  wire [7:0] add_542146;
  wire [7:0] sel_542147;
  wire [7:0] add_542150;
  wire [7:0] sel_542151;
  wire [7:0] add_542154;
  wire [7:0] sel_542155;
  wire [7:0] add_542158;
  wire [7:0] sel_542159;
  wire [7:0] add_542162;
  wire [7:0] sel_542163;
  wire [7:0] add_542166;
  wire [7:0] sel_542167;
  wire [7:0] add_542170;
  wire [7:0] sel_542171;
  wire [7:0] add_542174;
  wire [7:0] sel_542175;
  wire [7:0] add_542178;
  wire [7:0] sel_542179;
  wire [7:0] add_542182;
  wire [7:0] sel_542183;
  wire [7:0] add_542186;
  wire [7:0] sel_542187;
  wire [7:0] add_542190;
  wire [7:0] sel_542191;
  wire [7:0] add_542194;
  wire [7:0] sel_542195;
  wire [7:0] add_542198;
  wire [7:0] sel_542199;
  wire [7:0] add_542202;
  wire [7:0] sel_542203;
  wire [7:0] add_542206;
  wire [7:0] sel_542207;
  wire [7:0] add_542210;
  wire [7:0] sel_542211;
  wire [7:0] add_542214;
  wire [7:0] sel_542215;
  wire [7:0] add_542218;
  wire [7:0] sel_542219;
  wire [7:0] add_542222;
  wire [7:0] sel_542223;
  wire [7:0] add_542226;
  wire [7:0] sel_542227;
  wire [7:0] add_542230;
  wire [7:0] sel_542231;
  wire [7:0] add_542234;
  wire [7:0] sel_542235;
  wire [7:0] add_542238;
  wire [7:0] sel_542239;
  wire [7:0] add_542242;
  wire [7:0] sel_542243;
  wire [7:0] add_542246;
  wire [7:0] sel_542247;
  wire [7:0] add_542250;
  wire [7:0] sel_542251;
  wire [7:0] add_542254;
  wire [7:0] sel_542255;
  wire [7:0] add_542258;
  wire [7:0] sel_542259;
  wire [7:0] add_542262;
  wire [7:0] sel_542263;
  wire [7:0] add_542266;
  wire [7:0] sel_542267;
  wire [7:0] add_542270;
  wire [7:0] sel_542271;
  wire [7:0] add_542274;
  wire [7:0] sel_542275;
  wire [7:0] add_542278;
  wire [7:0] sel_542279;
  wire [7:0] add_542282;
  wire [7:0] sel_542283;
  wire [7:0] add_542286;
  wire [7:0] sel_542287;
  wire [7:0] add_542290;
  wire [7:0] sel_542291;
  wire [7:0] add_542294;
  wire [7:0] sel_542295;
  wire [7:0] add_542298;
  wire [7:0] sel_542299;
  wire [7:0] add_542303;
  wire [15:0] array_index_542304;
  wire [7:0] sel_542305;
  wire [7:0] add_542308;
  wire [7:0] sel_542309;
  wire [7:0] add_542312;
  wire [7:0] sel_542313;
  wire [7:0] add_542316;
  wire [7:0] sel_542317;
  wire [7:0] add_542320;
  wire [7:0] sel_542321;
  wire [7:0] add_542324;
  wire [7:0] sel_542325;
  wire [7:0] add_542328;
  wire [7:0] sel_542329;
  wire [7:0] add_542332;
  wire [7:0] sel_542333;
  wire [7:0] add_542336;
  wire [7:0] sel_542337;
  wire [7:0] add_542340;
  wire [7:0] sel_542341;
  wire [7:0] add_542344;
  wire [7:0] sel_542345;
  wire [7:0] add_542348;
  wire [7:0] sel_542349;
  wire [7:0] add_542352;
  wire [7:0] sel_542353;
  wire [7:0] add_542356;
  wire [7:0] sel_542357;
  wire [7:0] add_542360;
  wire [7:0] sel_542361;
  wire [7:0] add_542364;
  wire [7:0] sel_542365;
  wire [7:0] add_542368;
  wire [7:0] sel_542369;
  wire [7:0] add_542372;
  wire [7:0] sel_542373;
  wire [7:0] add_542376;
  wire [7:0] sel_542377;
  wire [7:0] add_542380;
  wire [7:0] sel_542381;
  wire [7:0] add_542384;
  wire [7:0] sel_542385;
  wire [7:0] add_542388;
  wire [7:0] sel_542389;
  wire [7:0] add_542392;
  wire [7:0] sel_542393;
  wire [7:0] add_542396;
  wire [7:0] sel_542397;
  wire [7:0] add_542400;
  wire [7:0] sel_542401;
  wire [7:0] add_542404;
  wire [7:0] sel_542405;
  wire [7:0] add_542408;
  wire [7:0] sel_542409;
  wire [7:0] add_542412;
  wire [7:0] sel_542413;
  wire [7:0] add_542416;
  wire [7:0] sel_542417;
  wire [7:0] add_542420;
  wire [7:0] sel_542421;
  wire [7:0] add_542424;
  wire [7:0] sel_542425;
  wire [7:0] add_542428;
  wire [7:0] sel_542429;
  wire [7:0] add_542432;
  wire [7:0] sel_542433;
  wire [7:0] add_542436;
  wire [7:0] sel_542437;
  wire [7:0] add_542440;
  wire [7:0] sel_542441;
  wire [7:0] add_542444;
  wire [7:0] sel_542445;
  wire [7:0] add_542448;
  wire [7:0] sel_542449;
  wire [7:0] add_542452;
  wire [7:0] sel_542453;
  wire [7:0] add_542456;
  wire [7:0] sel_542457;
  wire [7:0] add_542460;
  wire [7:0] sel_542461;
  wire [7:0] add_542464;
  wire [7:0] sel_542465;
  wire [7:0] add_542468;
  wire [7:0] sel_542469;
  wire [7:0] add_542472;
  wire [7:0] sel_542473;
  wire [7:0] add_542476;
  wire [7:0] sel_542477;
  wire [7:0] add_542480;
  wire [7:0] sel_542481;
  wire [7:0] add_542484;
  wire [7:0] sel_542485;
  wire [7:0] add_542488;
  wire [7:0] sel_542489;
  wire [7:0] add_542492;
  wire [7:0] sel_542493;
  wire [7:0] add_542496;
  wire [7:0] sel_542497;
  wire [7:0] add_542500;
  wire [7:0] sel_542501;
  wire [7:0] add_542504;
  wire [7:0] sel_542505;
  wire [7:0] add_542508;
  wire [7:0] sel_542509;
  wire [7:0] add_542512;
  wire [7:0] sel_542513;
  wire [7:0] add_542516;
  wire [7:0] sel_542517;
  wire [7:0] add_542520;
  wire [7:0] sel_542521;
  wire [7:0] add_542524;
  wire [7:0] sel_542525;
  wire [7:0] add_542528;
  wire [7:0] sel_542529;
  wire [7:0] add_542532;
  wire [7:0] sel_542533;
  wire [7:0] add_542536;
  wire [7:0] sel_542537;
  wire [7:0] add_542540;
  wire [7:0] sel_542541;
  wire [7:0] add_542544;
  wire [7:0] sel_542545;
  wire [7:0] add_542548;
  wire [7:0] sel_542549;
  wire [7:0] add_542552;
  wire [7:0] sel_542553;
  wire [7:0] add_542556;
  wire [7:0] sel_542557;
  wire [7:0] add_542560;
  wire [7:0] sel_542561;
  wire [7:0] add_542564;
  wire [7:0] sel_542565;
  wire [7:0] add_542568;
  wire [7:0] sel_542569;
  wire [7:0] add_542572;
  wire [7:0] sel_542573;
  wire [7:0] add_542576;
  wire [7:0] sel_542577;
  wire [7:0] add_542580;
  wire [7:0] sel_542581;
  wire [7:0] add_542584;
  wire [7:0] sel_542585;
  wire [7:0] add_542588;
  wire [7:0] sel_542589;
  wire [7:0] add_542592;
  wire [7:0] sel_542593;
  wire [7:0] add_542596;
  wire [7:0] sel_542597;
  wire [7:0] add_542600;
  wire [7:0] sel_542601;
  wire [7:0] add_542605;
  wire [15:0] array_index_542606;
  wire [7:0] sel_542607;
  wire [7:0] add_542610;
  wire [7:0] sel_542611;
  wire [7:0] add_542614;
  wire [7:0] sel_542615;
  wire [7:0] add_542618;
  wire [7:0] sel_542619;
  wire [7:0] add_542622;
  wire [7:0] sel_542623;
  wire [7:0] add_542626;
  wire [7:0] sel_542627;
  wire [7:0] add_542630;
  wire [7:0] sel_542631;
  wire [7:0] add_542634;
  wire [7:0] sel_542635;
  wire [7:0] add_542638;
  wire [7:0] sel_542639;
  wire [7:0] add_542642;
  wire [7:0] sel_542643;
  wire [7:0] add_542646;
  wire [7:0] sel_542647;
  wire [7:0] add_542650;
  wire [7:0] sel_542651;
  wire [7:0] add_542654;
  wire [7:0] sel_542655;
  wire [7:0] add_542658;
  wire [7:0] sel_542659;
  wire [7:0] add_542662;
  wire [7:0] sel_542663;
  wire [7:0] add_542666;
  wire [7:0] sel_542667;
  wire [7:0] add_542670;
  wire [7:0] sel_542671;
  wire [7:0] add_542674;
  wire [7:0] sel_542675;
  wire [7:0] add_542678;
  wire [7:0] sel_542679;
  wire [7:0] add_542682;
  wire [7:0] sel_542683;
  wire [7:0] add_542686;
  wire [7:0] sel_542687;
  wire [7:0] add_542690;
  wire [7:0] sel_542691;
  wire [7:0] add_542694;
  wire [7:0] sel_542695;
  wire [7:0] add_542698;
  wire [7:0] sel_542699;
  wire [7:0] add_542702;
  wire [7:0] sel_542703;
  wire [7:0] add_542706;
  wire [7:0] sel_542707;
  wire [7:0] add_542710;
  wire [7:0] sel_542711;
  wire [7:0] add_542714;
  wire [7:0] sel_542715;
  wire [7:0] add_542718;
  wire [7:0] sel_542719;
  wire [7:0] add_542722;
  wire [7:0] sel_542723;
  wire [7:0] add_542726;
  wire [7:0] sel_542727;
  wire [7:0] add_542730;
  wire [7:0] sel_542731;
  wire [7:0] add_542734;
  wire [7:0] sel_542735;
  wire [7:0] add_542738;
  wire [7:0] sel_542739;
  wire [7:0] add_542742;
  wire [7:0] sel_542743;
  wire [7:0] add_542746;
  wire [7:0] sel_542747;
  wire [7:0] add_542750;
  wire [7:0] sel_542751;
  wire [7:0] add_542754;
  wire [7:0] sel_542755;
  wire [7:0] add_542758;
  wire [7:0] sel_542759;
  wire [7:0] add_542762;
  wire [7:0] sel_542763;
  wire [7:0] add_542766;
  wire [7:0] sel_542767;
  wire [7:0] add_542770;
  wire [7:0] sel_542771;
  wire [7:0] add_542774;
  wire [7:0] sel_542775;
  wire [7:0] add_542778;
  wire [7:0] sel_542779;
  wire [7:0] add_542782;
  wire [7:0] sel_542783;
  wire [7:0] add_542786;
  wire [7:0] sel_542787;
  wire [7:0] add_542790;
  wire [7:0] sel_542791;
  wire [7:0] add_542794;
  wire [7:0] sel_542795;
  wire [7:0] add_542798;
  wire [7:0] sel_542799;
  wire [7:0] add_542802;
  wire [7:0] sel_542803;
  wire [7:0] add_542806;
  wire [7:0] sel_542807;
  wire [7:0] add_542810;
  wire [7:0] sel_542811;
  wire [7:0] add_542814;
  wire [7:0] sel_542815;
  wire [7:0] add_542818;
  wire [7:0] sel_542819;
  wire [7:0] add_542822;
  wire [7:0] sel_542823;
  wire [7:0] add_542826;
  wire [7:0] sel_542827;
  wire [7:0] add_542830;
  wire [7:0] sel_542831;
  wire [7:0] add_542834;
  wire [7:0] sel_542835;
  wire [7:0] add_542838;
  wire [7:0] sel_542839;
  wire [7:0] add_542842;
  wire [7:0] sel_542843;
  wire [7:0] add_542846;
  wire [7:0] sel_542847;
  wire [7:0] add_542850;
  wire [7:0] sel_542851;
  wire [7:0] add_542854;
  wire [7:0] sel_542855;
  wire [7:0] add_542858;
  wire [7:0] sel_542859;
  wire [7:0] add_542862;
  wire [7:0] sel_542863;
  wire [7:0] add_542866;
  wire [7:0] sel_542867;
  wire [7:0] add_542870;
  wire [7:0] sel_542871;
  wire [7:0] add_542874;
  wire [7:0] sel_542875;
  wire [7:0] add_542878;
  wire [7:0] sel_542879;
  wire [7:0] add_542882;
  wire [7:0] sel_542883;
  wire [7:0] add_542886;
  wire [7:0] sel_542887;
  wire [7:0] add_542890;
  wire [7:0] sel_542891;
  wire [7:0] add_542894;
  wire [7:0] sel_542895;
  wire [7:0] add_542898;
  wire [7:0] sel_542899;
  wire [7:0] add_542902;
  wire [7:0] sel_542903;
  wire [7:0] add_542907;
  wire [15:0] array_index_542908;
  wire [7:0] sel_542909;
  wire [7:0] add_542912;
  wire [7:0] sel_542913;
  wire [7:0] add_542916;
  wire [7:0] sel_542917;
  wire [7:0] add_542920;
  wire [7:0] sel_542921;
  wire [7:0] add_542924;
  wire [7:0] sel_542925;
  wire [7:0] add_542928;
  wire [7:0] sel_542929;
  wire [7:0] add_542932;
  wire [7:0] sel_542933;
  wire [7:0] add_542936;
  wire [7:0] sel_542937;
  wire [7:0] add_542940;
  wire [7:0] sel_542941;
  wire [7:0] add_542944;
  wire [7:0] sel_542945;
  wire [7:0] add_542948;
  wire [7:0] sel_542949;
  wire [7:0] add_542952;
  wire [7:0] sel_542953;
  wire [7:0] add_542956;
  wire [7:0] sel_542957;
  wire [7:0] add_542960;
  wire [7:0] sel_542961;
  wire [7:0] add_542964;
  wire [7:0] sel_542965;
  wire [7:0] add_542968;
  wire [7:0] sel_542969;
  wire [7:0] add_542972;
  wire [7:0] sel_542973;
  wire [7:0] add_542976;
  wire [7:0] sel_542977;
  wire [7:0] add_542980;
  wire [7:0] sel_542981;
  wire [7:0] add_542984;
  wire [7:0] sel_542985;
  wire [7:0] add_542988;
  wire [7:0] sel_542989;
  wire [7:0] add_542992;
  wire [7:0] sel_542993;
  wire [7:0] add_542996;
  wire [7:0] sel_542997;
  wire [7:0] add_543000;
  wire [7:0] sel_543001;
  wire [7:0] add_543004;
  wire [7:0] sel_543005;
  wire [7:0] add_543008;
  wire [7:0] sel_543009;
  wire [7:0] add_543012;
  wire [7:0] sel_543013;
  wire [7:0] add_543016;
  wire [7:0] sel_543017;
  wire [7:0] add_543020;
  wire [7:0] sel_543021;
  wire [7:0] add_543024;
  wire [7:0] sel_543025;
  wire [7:0] add_543028;
  wire [7:0] sel_543029;
  wire [7:0] add_543032;
  wire [7:0] sel_543033;
  wire [7:0] add_543036;
  wire [7:0] sel_543037;
  wire [7:0] add_543040;
  wire [7:0] sel_543041;
  wire [7:0] add_543044;
  wire [7:0] sel_543045;
  wire [7:0] add_543048;
  wire [7:0] sel_543049;
  wire [7:0] add_543052;
  wire [7:0] sel_543053;
  wire [7:0] add_543056;
  wire [7:0] sel_543057;
  wire [7:0] add_543060;
  wire [7:0] sel_543061;
  wire [7:0] add_543064;
  wire [7:0] sel_543065;
  wire [7:0] add_543068;
  wire [7:0] sel_543069;
  wire [7:0] add_543072;
  wire [7:0] sel_543073;
  wire [7:0] add_543076;
  wire [7:0] sel_543077;
  wire [7:0] add_543080;
  wire [7:0] sel_543081;
  wire [7:0] add_543084;
  wire [7:0] sel_543085;
  wire [7:0] add_543088;
  wire [7:0] sel_543089;
  wire [7:0] add_543092;
  wire [7:0] sel_543093;
  wire [7:0] add_543096;
  wire [7:0] sel_543097;
  wire [7:0] add_543100;
  wire [7:0] sel_543101;
  wire [7:0] add_543104;
  wire [7:0] sel_543105;
  wire [7:0] add_543108;
  wire [7:0] sel_543109;
  wire [7:0] add_543112;
  wire [7:0] sel_543113;
  wire [7:0] add_543116;
  wire [7:0] sel_543117;
  wire [7:0] add_543120;
  wire [7:0] sel_543121;
  wire [7:0] add_543124;
  wire [7:0] sel_543125;
  wire [7:0] add_543128;
  wire [7:0] sel_543129;
  wire [7:0] add_543132;
  wire [7:0] sel_543133;
  wire [7:0] add_543136;
  wire [7:0] sel_543137;
  wire [7:0] add_543140;
  wire [7:0] sel_543141;
  wire [7:0] add_543144;
  wire [7:0] sel_543145;
  wire [7:0] add_543148;
  wire [7:0] sel_543149;
  wire [7:0] add_543152;
  wire [7:0] sel_543153;
  wire [7:0] add_543156;
  wire [7:0] sel_543157;
  wire [7:0] add_543160;
  wire [7:0] sel_543161;
  wire [7:0] add_543164;
  wire [7:0] sel_543165;
  wire [7:0] add_543168;
  wire [7:0] sel_543169;
  wire [7:0] add_543172;
  wire [7:0] sel_543173;
  wire [7:0] add_543176;
  wire [7:0] sel_543177;
  wire [7:0] add_543180;
  wire [7:0] sel_543181;
  wire [7:0] add_543184;
  wire [7:0] sel_543185;
  wire [7:0] add_543188;
  wire [7:0] sel_543189;
  wire [7:0] add_543192;
  wire [7:0] sel_543193;
  wire [7:0] add_543196;
  wire [7:0] sel_543197;
  wire [7:0] add_543200;
  wire [7:0] sel_543201;
  wire [7:0] add_543204;
  wire [7:0] sel_543205;
  wire [7:0] add_543209;
  wire [15:0] array_index_543210;
  wire [7:0] sel_543211;
  wire [7:0] add_543214;
  wire [7:0] sel_543215;
  wire [7:0] add_543218;
  wire [7:0] sel_543219;
  wire [7:0] add_543222;
  wire [7:0] sel_543223;
  wire [7:0] add_543226;
  wire [7:0] sel_543227;
  wire [7:0] add_543230;
  wire [7:0] sel_543231;
  wire [7:0] add_543234;
  wire [7:0] sel_543235;
  wire [7:0] add_543238;
  wire [7:0] sel_543239;
  wire [7:0] add_543242;
  wire [7:0] sel_543243;
  wire [7:0] add_543246;
  wire [7:0] sel_543247;
  wire [7:0] add_543250;
  wire [7:0] sel_543251;
  wire [7:0] add_543254;
  wire [7:0] sel_543255;
  wire [7:0] add_543258;
  wire [7:0] sel_543259;
  wire [7:0] add_543262;
  wire [7:0] sel_543263;
  wire [7:0] add_543266;
  wire [7:0] sel_543267;
  wire [7:0] add_543270;
  wire [7:0] sel_543271;
  wire [7:0] add_543274;
  wire [7:0] sel_543275;
  wire [7:0] add_543278;
  wire [7:0] sel_543279;
  wire [7:0] add_543282;
  wire [7:0] sel_543283;
  wire [7:0] add_543286;
  wire [7:0] sel_543287;
  wire [7:0] add_543290;
  wire [7:0] sel_543291;
  wire [7:0] add_543294;
  wire [7:0] sel_543295;
  wire [7:0] add_543298;
  wire [7:0] sel_543299;
  wire [7:0] add_543302;
  wire [7:0] sel_543303;
  wire [7:0] add_543306;
  wire [7:0] sel_543307;
  wire [7:0] add_543310;
  wire [7:0] sel_543311;
  wire [7:0] add_543314;
  wire [7:0] sel_543315;
  wire [7:0] add_543318;
  wire [7:0] sel_543319;
  wire [7:0] add_543322;
  wire [7:0] sel_543323;
  wire [7:0] add_543326;
  wire [7:0] sel_543327;
  wire [7:0] add_543330;
  wire [7:0] sel_543331;
  wire [7:0] add_543334;
  wire [7:0] sel_543335;
  wire [7:0] add_543338;
  wire [7:0] sel_543339;
  wire [7:0] add_543342;
  wire [7:0] sel_543343;
  wire [7:0] add_543346;
  wire [7:0] sel_543347;
  wire [7:0] add_543350;
  wire [7:0] sel_543351;
  wire [7:0] add_543354;
  wire [7:0] sel_543355;
  wire [7:0] add_543358;
  wire [7:0] sel_543359;
  wire [7:0] add_543362;
  wire [7:0] sel_543363;
  wire [7:0] add_543366;
  wire [7:0] sel_543367;
  wire [7:0] add_543370;
  wire [7:0] sel_543371;
  wire [7:0] add_543374;
  wire [7:0] sel_543375;
  wire [7:0] add_543378;
  wire [7:0] sel_543379;
  wire [7:0] add_543382;
  wire [7:0] sel_543383;
  wire [7:0] add_543386;
  wire [7:0] sel_543387;
  wire [7:0] add_543390;
  wire [7:0] sel_543391;
  wire [7:0] add_543394;
  wire [7:0] sel_543395;
  wire [7:0] add_543398;
  wire [7:0] sel_543399;
  wire [7:0] add_543402;
  wire [7:0] sel_543403;
  wire [7:0] add_543406;
  wire [7:0] sel_543407;
  wire [7:0] add_543410;
  wire [7:0] sel_543411;
  wire [7:0] add_543414;
  wire [7:0] sel_543415;
  wire [7:0] add_543418;
  wire [7:0] sel_543419;
  wire [7:0] add_543422;
  wire [7:0] sel_543423;
  wire [7:0] add_543426;
  wire [7:0] sel_543427;
  wire [7:0] add_543430;
  wire [7:0] sel_543431;
  wire [7:0] add_543434;
  wire [7:0] sel_543435;
  wire [7:0] add_543438;
  wire [7:0] sel_543439;
  wire [7:0] add_543442;
  wire [7:0] sel_543443;
  wire [7:0] add_543446;
  wire [7:0] sel_543447;
  wire [7:0] add_543450;
  wire [7:0] sel_543451;
  wire [7:0] add_543454;
  wire [7:0] sel_543455;
  wire [7:0] add_543458;
  wire [7:0] sel_543459;
  wire [7:0] add_543462;
  wire [7:0] sel_543463;
  wire [7:0] add_543466;
  wire [7:0] sel_543467;
  wire [7:0] add_543470;
  wire [7:0] sel_543471;
  wire [7:0] add_543474;
  wire [7:0] sel_543475;
  wire [7:0] add_543478;
  wire [7:0] sel_543479;
  wire [7:0] add_543482;
  wire [7:0] sel_543483;
  wire [7:0] add_543486;
  wire [7:0] sel_543487;
  wire [7:0] add_543490;
  wire [7:0] sel_543491;
  wire [7:0] add_543494;
  wire [7:0] sel_543495;
  wire [7:0] add_543498;
  wire [7:0] sel_543499;
  wire [7:0] add_543502;
  wire [7:0] sel_543503;
  wire [7:0] add_543506;
  wire [7:0] sel_543507;
  wire [7:0] add_543511;
  wire [15:0] array_index_543512;
  wire [7:0] sel_543513;
  wire [7:0] add_543516;
  wire [7:0] sel_543517;
  wire [7:0] add_543520;
  wire [7:0] sel_543521;
  wire [7:0] add_543524;
  wire [7:0] sel_543525;
  wire [7:0] add_543528;
  wire [7:0] sel_543529;
  wire [7:0] add_543532;
  wire [7:0] sel_543533;
  wire [7:0] add_543536;
  wire [7:0] sel_543537;
  wire [7:0] add_543540;
  wire [7:0] sel_543541;
  wire [7:0] add_543544;
  wire [7:0] sel_543545;
  wire [7:0] add_543548;
  wire [7:0] sel_543549;
  wire [7:0] add_543552;
  wire [7:0] sel_543553;
  wire [7:0] add_543556;
  wire [7:0] sel_543557;
  wire [7:0] add_543560;
  wire [7:0] sel_543561;
  wire [7:0] add_543564;
  wire [7:0] sel_543565;
  wire [7:0] add_543568;
  wire [7:0] sel_543569;
  wire [7:0] add_543572;
  wire [7:0] sel_543573;
  wire [7:0] add_543576;
  wire [7:0] sel_543577;
  wire [7:0] add_543580;
  wire [7:0] sel_543581;
  wire [7:0] add_543584;
  wire [7:0] sel_543585;
  wire [7:0] add_543588;
  wire [7:0] sel_543589;
  wire [7:0] add_543592;
  wire [7:0] sel_543593;
  wire [7:0] add_543596;
  wire [7:0] sel_543597;
  wire [7:0] add_543600;
  wire [7:0] sel_543601;
  wire [7:0] add_543604;
  wire [7:0] sel_543605;
  wire [7:0] add_543608;
  wire [7:0] sel_543609;
  wire [7:0] add_543612;
  wire [7:0] sel_543613;
  wire [7:0] add_543616;
  wire [7:0] sel_543617;
  wire [7:0] add_543620;
  wire [7:0] sel_543621;
  wire [7:0] add_543624;
  wire [7:0] sel_543625;
  wire [7:0] add_543628;
  wire [7:0] sel_543629;
  wire [7:0] add_543632;
  wire [7:0] sel_543633;
  wire [7:0] add_543636;
  wire [7:0] sel_543637;
  wire [7:0] add_543640;
  wire [7:0] sel_543641;
  wire [7:0] add_543644;
  wire [7:0] sel_543645;
  wire [7:0] add_543648;
  wire [7:0] sel_543649;
  wire [7:0] add_543652;
  wire [7:0] sel_543653;
  wire [7:0] add_543656;
  wire [7:0] sel_543657;
  wire [7:0] add_543660;
  wire [7:0] sel_543661;
  wire [7:0] add_543664;
  wire [7:0] sel_543665;
  wire [7:0] add_543668;
  wire [7:0] sel_543669;
  wire [7:0] add_543672;
  wire [7:0] sel_543673;
  wire [7:0] add_543676;
  wire [7:0] sel_543677;
  wire [7:0] add_543680;
  wire [7:0] sel_543681;
  wire [7:0] add_543684;
  wire [7:0] sel_543685;
  wire [7:0] add_543688;
  wire [7:0] sel_543689;
  wire [7:0] add_543692;
  wire [7:0] sel_543693;
  wire [7:0] add_543696;
  wire [7:0] sel_543697;
  wire [7:0] add_543700;
  wire [7:0] sel_543701;
  wire [7:0] add_543704;
  wire [7:0] sel_543705;
  wire [7:0] add_543708;
  wire [7:0] sel_543709;
  wire [7:0] add_543712;
  wire [7:0] sel_543713;
  wire [7:0] add_543716;
  wire [7:0] sel_543717;
  wire [7:0] add_543720;
  wire [7:0] sel_543721;
  wire [7:0] add_543724;
  wire [7:0] sel_543725;
  wire [7:0] add_543728;
  wire [7:0] sel_543729;
  wire [7:0] add_543732;
  wire [7:0] sel_543733;
  wire [7:0] add_543736;
  wire [7:0] sel_543737;
  wire [7:0] add_543740;
  wire [7:0] sel_543741;
  wire [7:0] add_543744;
  wire [7:0] sel_543745;
  wire [7:0] add_543748;
  wire [7:0] sel_543749;
  wire [7:0] add_543752;
  wire [7:0] sel_543753;
  wire [7:0] add_543756;
  wire [7:0] sel_543757;
  wire [7:0] add_543760;
  wire [7:0] sel_543761;
  wire [7:0] add_543764;
  wire [7:0] sel_543765;
  wire [7:0] add_543768;
  wire [7:0] sel_543769;
  wire [7:0] add_543772;
  wire [7:0] sel_543773;
  wire [7:0] add_543776;
  wire [7:0] sel_543777;
  wire [7:0] add_543780;
  wire [7:0] sel_543781;
  wire [7:0] add_543784;
  wire [7:0] sel_543785;
  wire [7:0] add_543788;
  wire [7:0] sel_543789;
  wire [7:0] add_543792;
  wire [7:0] sel_543793;
  wire [7:0] add_543796;
  wire [7:0] sel_543797;
  wire [7:0] add_543800;
  wire [7:0] sel_543801;
  wire [7:0] add_543804;
  wire [7:0] sel_543805;
  wire [7:0] add_543808;
  wire [7:0] sel_543809;
  wire [7:0] add_543813;
  wire [15:0] array_index_543814;
  wire [7:0] sel_543815;
  wire [7:0] add_543818;
  wire [7:0] sel_543819;
  wire [7:0] add_543822;
  wire [7:0] sel_543823;
  wire [7:0] add_543826;
  wire [7:0] sel_543827;
  wire [7:0] add_543830;
  wire [7:0] sel_543831;
  wire [7:0] add_543834;
  wire [7:0] sel_543835;
  wire [7:0] add_543838;
  wire [7:0] sel_543839;
  wire [7:0] add_543842;
  wire [7:0] sel_543843;
  wire [7:0] add_543846;
  wire [7:0] sel_543847;
  wire [7:0] add_543850;
  wire [7:0] sel_543851;
  wire [7:0] add_543854;
  wire [7:0] sel_543855;
  wire [7:0] add_543858;
  wire [7:0] sel_543859;
  wire [7:0] add_543862;
  wire [7:0] sel_543863;
  wire [7:0] add_543866;
  wire [7:0] sel_543867;
  wire [7:0] add_543870;
  wire [7:0] sel_543871;
  wire [7:0] add_543874;
  wire [7:0] sel_543875;
  wire [7:0] add_543878;
  wire [7:0] sel_543879;
  wire [7:0] add_543882;
  wire [7:0] sel_543883;
  wire [7:0] add_543886;
  wire [7:0] sel_543887;
  wire [7:0] add_543890;
  wire [7:0] sel_543891;
  wire [7:0] add_543894;
  wire [7:0] sel_543895;
  wire [7:0] add_543898;
  wire [7:0] sel_543899;
  wire [7:0] add_543902;
  wire [7:0] sel_543903;
  wire [7:0] add_543906;
  wire [7:0] sel_543907;
  wire [7:0] add_543910;
  wire [7:0] sel_543911;
  wire [7:0] add_543914;
  wire [7:0] sel_543915;
  wire [7:0] add_543918;
  wire [7:0] sel_543919;
  wire [7:0] add_543922;
  wire [7:0] sel_543923;
  wire [7:0] add_543926;
  wire [7:0] sel_543927;
  wire [7:0] add_543930;
  wire [7:0] sel_543931;
  wire [7:0] add_543934;
  wire [7:0] sel_543935;
  wire [7:0] add_543938;
  wire [7:0] sel_543939;
  wire [7:0] add_543942;
  wire [7:0] sel_543943;
  wire [7:0] add_543946;
  wire [7:0] sel_543947;
  wire [7:0] add_543950;
  wire [7:0] sel_543951;
  wire [7:0] add_543954;
  wire [7:0] sel_543955;
  wire [7:0] add_543958;
  wire [7:0] sel_543959;
  wire [7:0] add_543962;
  wire [7:0] sel_543963;
  wire [7:0] add_543966;
  wire [7:0] sel_543967;
  wire [7:0] add_543970;
  wire [7:0] sel_543971;
  wire [7:0] add_543974;
  wire [7:0] sel_543975;
  wire [7:0] add_543978;
  wire [7:0] sel_543979;
  wire [7:0] add_543982;
  wire [7:0] sel_543983;
  wire [7:0] add_543986;
  wire [7:0] sel_543987;
  wire [7:0] add_543990;
  wire [7:0] sel_543991;
  wire [7:0] add_543994;
  wire [7:0] sel_543995;
  wire [7:0] add_543998;
  wire [7:0] sel_543999;
  wire [7:0] add_544002;
  wire [7:0] sel_544003;
  wire [7:0] add_544006;
  wire [7:0] sel_544007;
  wire [7:0] add_544010;
  wire [7:0] sel_544011;
  wire [7:0] add_544014;
  wire [7:0] sel_544015;
  wire [7:0] add_544018;
  wire [7:0] sel_544019;
  wire [7:0] add_544022;
  wire [7:0] sel_544023;
  wire [7:0] add_544026;
  wire [7:0] sel_544027;
  wire [7:0] add_544030;
  wire [7:0] sel_544031;
  wire [7:0] add_544034;
  wire [7:0] sel_544035;
  wire [7:0] add_544038;
  wire [7:0] sel_544039;
  wire [7:0] add_544042;
  wire [7:0] sel_544043;
  wire [7:0] add_544046;
  wire [7:0] sel_544047;
  wire [7:0] add_544050;
  wire [7:0] sel_544051;
  wire [7:0] add_544054;
  wire [7:0] sel_544055;
  wire [7:0] add_544058;
  wire [7:0] sel_544059;
  wire [7:0] add_544062;
  wire [7:0] sel_544063;
  wire [7:0] add_544066;
  wire [7:0] sel_544067;
  wire [7:0] add_544070;
  wire [7:0] sel_544071;
  wire [7:0] add_544074;
  wire [7:0] sel_544075;
  wire [7:0] add_544078;
  wire [7:0] sel_544079;
  wire [7:0] add_544082;
  wire [7:0] sel_544083;
  wire [7:0] add_544086;
  wire [7:0] sel_544087;
  wire [7:0] add_544090;
  wire [7:0] sel_544091;
  wire [7:0] add_544094;
  wire [7:0] sel_544095;
  wire [7:0] add_544098;
  wire [7:0] sel_544099;
  wire [7:0] add_544102;
  wire [7:0] sel_544103;
  wire [7:0] add_544106;
  wire [7:0] sel_544107;
  wire [7:0] add_544110;
  wire [7:0] sel_544111;
  wire [7:0] add_544115;
  wire [15:0] array_index_544116;
  wire [7:0] sel_544117;
  wire [7:0] add_544120;
  wire [7:0] sel_544121;
  wire [7:0] add_544124;
  wire [7:0] sel_544125;
  wire [7:0] add_544128;
  wire [7:0] sel_544129;
  wire [7:0] add_544132;
  wire [7:0] sel_544133;
  wire [7:0] add_544136;
  wire [7:0] sel_544137;
  wire [7:0] add_544140;
  wire [7:0] sel_544141;
  wire [7:0] add_544144;
  wire [7:0] sel_544145;
  wire [7:0] add_544148;
  wire [7:0] sel_544149;
  wire [7:0] add_544152;
  wire [7:0] sel_544153;
  wire [7:0] add_544156;
  wire [7:0] sel_544157;
  wire [7:0] add_544160;
  wire [7:0] sel_544161;
  wire [7:0] add_544164;
  wire [7:0] sel_544165;
  wire [7:0] add_544168;
  wire [7:0] sel_544169;
  wire [7:0] add_544172;
  wire [7:0] sel_544173;
  wire [7:0] add_544176;
  wire [7:0] sel_544177;
  wire [7:0] add_544180;
  wire [7:0] sel_544181;
  wire [7:0] add_544184;
  wire [7:0] sel_544185;
  wire [7:0] add_544188;
  wire [7:0] sel_544189;
  wire [7:0] add_544192;
  wire [7:0] sel_544193;
  wire [7:0] add_544196;
  wire [7:0] sel_544197;
  wire [7:0] add_544200;
  wire [7:0] sel_544201;
  wire [7:0] add_544204;
  wire [7:0] sel_544205;
  wire [7:0] add_544208;
  wire [7:0] sel_544209;
  wire [7:0] add_544212;
  wire [7:0] sel_544213;
  wire [7:0] add_544216;
  wire [7:0] sel_544217;
  wire [7:0] add_544220;
  wire [7:0] sel_544221;
  wire [7:0] add_544224;
  wire [7:0] sel_544225;
  wire [7:0] add_544228;
  wire [7:0] sel_544229;
  wire [7:0] add_544232;
  wire [7:0] sel_544233;
  wire [7:0] add_544236;
  wire [7:0] sel_544237;
  wire [7:0] add_544240;
  wire [7:0] sel_544241;
  wire [7:0] add_544244;
  wire [7:0] sel_544245;
  wire [7:0] add_544248;
  wire [7:0] sel_544249;
  wire [7:0] add_544252;
  wire [7:0] sel_544253;
  wire [7:0] add_544256;
  wire [7:0] sel_544257;
  wire [7:0] add_544260;
  wire [7:0] sel_544261;
  wire [7:0] add_544264;
  wire [7:0] sel_544265;
  wire [7:0] add_544268;
  wire [7:0] sel_544269;
  wire [7:0] add_544272;
  wire [7:0] sel_544273;
  wire [7:0] add_544276;
  wire [7:0] sel_544277;
  wire [7:0] add_544280;
  wire [7:0] sel_544281;
  wire [7:0] add_544284;
  wire [7:0] sel_544285;
  wire [7:0] add_544288;
  wire [7:0] sel_544289;
  wire [7:0] add_544292;
  wire [7:0] sel_544293;
  wire [7:0] add_544296;
  wire [7:0] sel_544297;
  wire [7:0] add_544300;
  wire [7:0] sel_544301;
  wire [7:0] add_544304;
  wire [7:0] sel_544305;
  wire [7:0] add_544308;
  wire [7:0] sel_544309;
  wire [7:0] add_544312;
  wire [7:0] sel_544313;
  wire [7:0] add_544316;
  wire [7:0] sel_544317;
  wire [7:0] add_544320;
  wire [7:0] sel_544321;
  wire [7:0] add_544324;
  wire [7:0] sel_544325;
  wire [7:0] add_544328;
  wire [7:0] sel_544329;
  wire [7:0] add_544332;
  wire [7:0] sel_544333;
  wire [7:0] add_544336;
  wire [7:0] sel_544337;
  wire [7:0] add_544340;
  wire [7:0] sel_544341;
  wire [7:0] add_544344;
  wire [7:0] sel_544345;
  wire [7:0] add_544348;
  wire [7:0] sel_544349;
  wire [7:0] add_544352;
  wire [7:0] sel_544353;
  wire [7:0] add_544356;
  wire [7:0] sel_544357;
  wire [7:0] add_544360;
  wire [7:0] sel_544361;
  wire [7:0] add_544364;
  wire [7:0] sel_544365;
  wire [7:0] add_544368;
  wire [7:0] sel_544369;
  wire [7:0] add_544372;
  wire [7:0] sel_544373;
  wire [7:0] add_544376;
  wire [7:0] sel_544377;
  wire [7:0] add_544380;
  wire [7:0] sel_544381;
  wire [7:0] add_544384;
  wire [7:0] sel_544385;
  wire [7:0] add_544388;
  wire [7:0] sel_544389;
  wire [7:0] add_544392;
  wire [7:0] sel_544393;
  wire [7:0] add_544396;
  wire [7:0] sel_544397;
  wire [7:0] add_544400;
  wire [7:0] sel_544401;
  wire [7:0] add_544404;
  wire [7:0] sel_544405;
  wire [7:0] add_544408;
  wire [7:0] sel_544409;
  wire [7:0] add_544412;
  wire [7:0] sel_544413;
  wire [7:0] add_544417;
  wire [15:0] array_index_544418;
  wire [7:0] sel_544419;
  wire [7:0] add_544422;
  wire [7:0] sel_544423;
  wire [7:0] add_544426;
  wire [7:0] sel_544427;
  wire [7:0] add_544430;
  wire [7:0] sel_544431;
  wire [7:0] add_544434;
  wire [7:0] sel_544435;
  wire [7:0] add_544438;
  wire [7:0] sel_544439;
  wire [7:0] add_544442;
  wire [7:0] sel_544443;
  wire [7:0] add_544446;
  wire [7:0] sel_544447;
  wire [7:0] add_544450;
  wire [7:0] sel_544451;
  wire [7:0] add_544454;
  wire [7:0] sel_544455;
  wire [7:0] add_544458;
  wire [7:0] sel_544459;
  wire [7:0] add_544462;
  wire [7:0] sel_544463;
  wire [7:0] add_544466;
  wire [7:0] sel_544467;
  wire [7:0] add_544470;
  wire [7:0] sel_544471;
  wire [7:0] add_544474;
  wire [7:0] sel_544475;
  wire [7:0] add_544478;
  wire [7:0] sel_544479;
  wire [7:0] add_544482;
  wire [7:0] sel_544483;
  wire [7:0] add_544486;
  wire [7:0] sel_544487;
  wire [7:0] add_544490;
  wire [7:0] sel_544491;
  wire [7:0] add_544494;
  wire [7:0] sel_544495;
  wire [7:0] add_544498;
  wire [7:0] sel_544499;
  wire [7:0] add_544502;
  wire [7:0] sel_544503;
  wire [7:0] add_544506;
  wire [7:0] sel_544507;
  wire [7:0] add_544510;
  wire [7:0] sel_544511;
  wire [7:0] add_544514;
  wire [7:0] sel_544515;
  wire [7:0] add_544518;
  wire [7:0] sel_544519;
  wire [7:0] add_544522;
  wire [7:0] sel_544523;
  wire [7:0] add_544526;
  wire [7:0] sel_544527;
  wire [7:0] add_544530;
  wire [7:0] sel_544531;
  wire [7:0] add_544534;
  wire [7:0] sel_544535;
  wire [7:0] add_544538;
  wire [7:0] sel_544539;
  wire [7:0] add_544542;
  wire [7:0] sel_544543;
  wire [7:0] add_544546;
  wire [7:0] sel_544547;
  wire [7:0] add_544550;
  wire [7:0] sel_544551;
  wire [7:0] add_544554;
  wire [7:0] sel_544555;
  wire [7:0] add_544558;
  wire [7:0] sel_544559;
  wire [7:0] add_544562;
  wire [7:0] sel_544563;
  wire [7:0] add_544566;
  wire [7:0] sel_544567;
  wire [7:0] add_544570;
  wire [7:0] sel_544571;
  wire [7:0] add_544574;
  wire [7:0] sel_544575;
  wire [7:0] add_544578;
  wire [7:0] sel_544579;
  wire [7:0] add_544582;
  wire [7:0] sel_544583;
  wire [7:0] add_544586;
  wire [7:0] sel_544587;
  wire [7:0] add_544590;
  wire [7:0] sel_544591;
  wire [7:0] add_544594;
  wire [7:0] sel_544595;
  wire [7:0] add_544598;
  wire [7:0] sel_544599;
  wire [7:0] add_544602;
  wire [7:0] sel_544603;
  wire [7:0] add_544606;
  wire [7:0] sel_544607;
  wire [7:0] add_544610;
  wire [7:0] sel_544611;
  wire [7:0] add_544614;
  wire [7:0] sel_544615;
  wire [7:0] add_544618;
  wire [7:0] sel_544619;
  wire [7:0] add_544622;
  wire [7:0] sel_544623;
  wire [7:0] add_544626;
  wire [7:0] sel_544627;
  wire [7:0] add_544630;
  wire [7:0] sel_544631;
  wire [7:0] add_544634;
  wire [7:0] sel_544635;
  wire [7:0] add_544638;
  wire [7:0] sel_544639;
  wire [7:0] add_544642;
  wire [7:0] sel_544643;
  wire [7:0] add_544646;
  wire [7:0] sel_544647;
  wire [7:0] add_544650;
  wire [7:0] sel_544651;
  wire [7:0] add_544654;
  wire [7:0] sel_544655;
  wire [7:0] add_544658;
  wire [7:0] sel_544659;
  wire [7:0] add_544662;
  wire [7:0] sel_544663;
  wire [7:0] add_544666;
  wire [7:0] sel_544667;
  wire [7:0] add_544670;
  wire [7:0] sel_544671;
  wire [7:0] add_544674;
  wire [7:0] sel_544675;
  wire [7:0] add_544678;
  wire [7:0] sel_544679;
  wire [7:0] add_544682;
  wire [7:0] sel_544683;
  wire [7:0] add_544686;
  wire [7:0] sel_544687;
  wire [7:0] add_544690;
  wire [7:0] sel_544691;
  wire [7:0] add_544694;
  wire [7:0] sel_544695;
  wire [7:0] add_544698;
  wire [7:0] sel_544699;
  wire [7:0] add_544702;
  wire [7:0] sel_544703;
  wire [7:0] add_544706;
  wire [7:0] sel_544707;
  wire [7:0] add_544710;
  wire [7:0] sel_544711;
  wire [7:0] add_544714;
  wire [7:0] sel_544715;
  wire [7:0] add_544719;
  wire [15:0] array_index_544720;
  wire [7:0] sel_544721;
  wire [7:0] add_544724;
  wire [7:0] sel_544725;
  wire [7:0] add_544728;
  wire [7:0] sel_544729;
  wire [7:0] add_544732;
  wire [7:0] sel_544733;
  wire [7:0] add_544736;
  wire [7:0] sel_544737;
  wire [7:0] add_544740;
  wire [7:0] sel_544741;
  wire [7:0] add_544744;
  wire [7:0] sel_544745;
  wire [7:0] add_544748;
  wire [7:0] sel_544749;
  wire [7:0] add_544752;
  wire [7:0] sel_544753;
  wire [7:0] add_544756;
  wire [7:0] sel_544757;
  wire [7:0] add_544760;
  wire [7:0] sel_544761;
  wire [7:0] add_544764;
  wire [7:0] sel_544765;
  wire [7:0] add_544768;
  wire [7:0] sel_544769;
  wire [7:0] add_544772;
  wire [7:0] sel_544773;
  wire [7:0] add_544776;
  wire [7:0] sel_544777;
  wire [7:0] add_544780;
  wire [7:0] sel_544781;
  wire [7:0] add_544784;
  wire [7:0] sel_544785;
  wire [7:0] add_544788;
  wire [7:0] sel_544789;
  wire [7:0] add_544792;
  wire [7:0] sel_544793;
  wire [7:0] add_544796;
  wire [7:0] sel_544797;
  wire [7:0] add_544800;
  wire [7:0] sel_544801;
  wire [7:0] add_544804;
  wire [7:0] sel_544805;
  wire [7:0] add_544808;
  wire [7:0] sel_544809;
  wire [7:0] add_544812;
  wire [7:0] sel_544813;
  wire [7:0] add_544816;
  wire [7:0] sel_544817;
  wire [7:0] add_544820;
  wire [7:0] sel_544821;
  wire [7:0] add_544824;
  wire [7:0] sel_544825;
  wire [7:0] add_544828;
  wire [7:0] sel_544829;
  wire [7:0] add_544832;
  wire [7:0] sel_544833;
  wire [7:0] add_544836;
  wire [7:0] sel_544837;
  wire [7:0] add_544840;
  wire [7:0] sel_544841;
  wire [7:0] add_544844;
  wire [7:0] sel_544845;
  wire [7:0] add_544848;
  wire [7:0] sel_544849;
  wire [7:0] add_544852;
  wire [7:0] sel_544853;
  wire [7:0] add_544856;
  wire [7:0] sel_544857;
  wire [7:0] add_544860;
  wire [7:0] sel_544861;
  wire [7:0] add_544864;
  wire [7:0] sel_544865;
  wire [7:0] add_544868;
  wire [7:0] sel_544869;
  wire [7:0] add_544872;
  wire [7:0] sel_544873;
  wire [7:0] add_544876;
  wire [7:0] sel_544877;
  wire [7:0] add_544880;
  wire [7:0] sel_544881;
  wire [7:0] add_544884;
  wire [7:0] sel_544885;
  wire [7:0] add_544888;
  wire [7:0] sel_544889;
  wire [7:0] add_544892;
  wire [7:0] sel_544893;
  wire [7:0] add_544896;
  wire [7:0] sel_544897;
  wire [7:0] add_544900;
  wire [7:0] sel_544901;
  wire [7:0] add_544904;
  wire [7:0] sel_544905;
  wire [7:0] add_544908;
  wire [7:0] sel_544909;
  wire [7:0] add_544912;
  wire [7:0] sel_544913;
  wire [7:0] add_544916;
  wire [7:0] sel_544917;
  wire [7:0] add_544920;
  wire [7:0] sel_544921;
  wire [7:0] add_544924;
  wire [7:0] sel_544925;
  wire [7:0] add_544928;
  wire [7:0] sel_544929;
  wire [7:0] add_544932;
  wire [7:0] sel_544933;
  wire [7:0] add_544936;
  wire [7:0] sel_544937;
  wire [7:0] add_544940;
  wire [7:0] sel_544941;
  wire [7:0] add_544944;
  wire [7:0] sel_544945;
  wire [7:0] add_544948;
  wire [7:0] sel_544949;
  wire [7:0] add_544952;
  wire [7:0] sel_544953;
  wire [7:0] add_544956;
  wire [7:0] sel_544957;
  wire [7:0] add_544960;
  wire [7:0] sel_544961;
  wire [7:0] add_544964;
  wire [7:0] sel_544965;
  wire [7:0] add_544968;
  wire [7:0] sel_544969;
  wire [7:0] add_544972;
  wire [7:0] sel_544973;
  wire [7:0] add_544976;
  wire [7:0] sel_544977;
  wire [7:0] add_544980;
  wire [7:0] sel_544981;
  wire [7:0] add_544984;
  wire [7:0] sel_544985;
  wire [7:0] add_544988;
  wire [7:0] sel_544989;
  wire [7:0] add_544992;
  wire [7:0] sel_544993;
  wire [7:0] add_544996;
  wire [7:0] sel_544997;
  wire [7:0] add_545000;
  wire [7:0] sel_545001;
  wire [7:0] add_545004;
  wire [7:0] sel_545005;
  wire [7:0] add_545008;
  wire [7:0] sel_545009;
  wire [7:0] add_545012;
  wire [7:0] sel_545013;
  wire [7:0] add_545016;
  wire [7:0] sel_545017;
  wire [7:0] add_545021;
  wire [15:0] array_index_545022;
  wire [7:0] sel_545023;
  wire [7:0] add_545026;
  wire [7:0] sel_545027;
  wire [7:0] add_545030;
  wire [7:0] sel_545031;
  wire [7:0] add_545034;
  wire [7:0] sel_545035;
  wire [7:0] add_545038;
  wire [7:0] sel_545039;
  wire [7:0] add_545042;
  wire [7:0] sel_545043;
  wire [7:0] add_545046;
  wire [7:0] sel_545047;
  wire [7:0] add_545050;
  wire [7:0] sel_545051;
  wire [7:0] add_545054;
  wire [7:0] sel_545055;
  wire [7:0] add_545058;
  wire [7:0] sel_545059;
  wire [7:0] add_545062;
  wire [7:0] sel_545063;
  wire [7:0] add_545066;
  wire [7:0] sel_545067;
  wire [7:0] add_545070;
  wire [7:0] sel_545071;
  wire [7:0] add_545074;
  wire [7:0] sel_545075;
  wire [7:0] add_545078;
  wire [7:0] sel_545079;
  wire [7:0] add_545082;
  wire [7:0] sel_545083;
  wire [7:0] add_545086;
  wire [7:0] sel_545087;
  wire [7:0] add_545090;
  wire [7:0] sel_545091;
  wire [7:0] add_545094;
  wire [7:0] sel_545095;
  wire [7:0] add_545098;
  wire [7:0] sel_545099;
  wire [7:0] add_545102;
  wire [7:0] sel_545103;
  wire [7:0] add_545106;
  wire [7:0] sel_545107;
  wire [7:0] add_545110;
  wire [7:0] sel_545111;
  wire [7:0] add_545114;
  wire [7:0] sel_545115;
  wire [7:0] add_545118;
  wire [7:0] sel_545119;
  wire [7:0] add_545122;
  wire [7:0] sel_545123;
  wire [7:0] add_545126;
  wire [7:0] sel_545127;
  wire [7:0] add_545130;
  wire [7:0] sel_545131;
  wire [7:0] add_545134;
  wire [7:0] sel_545135;
  wire [7:0] add_545138;
  wire [7:0] sel_545139;
  wire [7:0] add_545142;
  wire [7:0] sel_545143;
  wire [7:0] add_545146;
  wire [7:0] sel_545147;
  wire [7:0] add_545150;
  wire [7:0] sel_545151;
  wire [7:0] add_545154;
  wire [7:0] sel_545155;
  wire [7:0] add_545158;
  wire [7:0] sel_545159;
  wire [7:0] add_545162;
  wire [7:0] sel_545163;
  wire [7:0] add_545166;
  wire [7:0] sel_545167;
  wire [7:0] add_545170;
  wire [7:0] sel_545171;
  wire [7:0] add_545174;
  wire [7:0] sel_545175;
  wire [7:0] add_545178;
  wire [7:0] sel_545179;
  wire [7:0] add_545182;
  wire [7:0] sel_545183;
  wire [7:0] add_545186;
  wire [7:0] sel_545187;
  wire [7:0] add_545190;
  wire [7:0] sel_545191;
  wire [7:0] add_545194;
  wire [7:0] sel_545195;
  wire [7:0] add_545198;
  wire [7:0] sel_545199;
  wire [7:0] add_545202;
  wire [7:0] sel_545203;
  wire [7:0] add_545206;
  wire [7:0] sel_545207;
  wire [7:0] add_545210;
  wire [7:0] sel_545211;
  wire [7:0] add_545214;
  wire [7:0] sel_545215;
  wire [7:0] add_545218;
  wire [7:0] sel_545219;
  wire [7:0] add_545222;
  wire [7:0] sel_545223;
  wire [7:0] add_545226;
  wire [7:0] sel_545227;
  wire [7:0] add_545230;
  wire [7:0] sel_545231;
  wire [7:0] add_545234;
  wire [7:0] sel_545235;
  wire [7:0] add_545238;
  wire [7:0] sel_545239;
  wire [7:0] add_545242;
  wire [7:0] sel_545243;
  wire [7:0] add_545246;
  wire [7:0] sel_545247;
  wire [7:0] add_545250;
  wire [7:0] sel_545251;
  wire [7:0] add_545254;
  wire [7:0] sel_545255;
  wire [7:0] add_545258;
  wire [7:0] sel_545259;
  wire [7:0] add_545262;
  wire [7:0] sel_545263;
  wire [7:0] add_545266;
  wire [7:0] sel_545267;
  wire [7:0] add_545270;
  wire [7:0] sel_545271;
  wire [7:0] add_545274;
  wire [7:0] sel_545275;
  wire [7:0] add_545278;
  wire [7:0] sel_545279;
  wire [7:0] add_545282;
  wire [7:0] sel_545283;
  wire [7:0] add_545286;
  wire [7:0] sel_545287;
  wire [7:0] add_545290;
  wire [7:0] sel_545291;
  wire [7:0] add_545294;
  wire [7:0] sel_545295;
  wire [7:0] add_545298;
  wire [7:0] sel_545299;
  wire [7:0] add_545302;
  wire [7:0] sel_545303;
  wire [7:0] add_545306;
  wire [7:0] sel_545307;
  wire [7:0] add_545310;
  wire [7:0] sel_545311;
  wire [7:0] add_545314;
  wire [7:0] sel_545315;
  wire [7:0] add_545318;
  wire [7:0] sel_545319;
  wire [7:0] add_545323;
  wire [15:0] array_index_545324;
  wire [7:0] sel_545325;
  wire [7:0] add_545328;
  wire [7:0] sel_545329;
  wire [7:0] add_545332;
  wire [7:0] sel_545333;
  wire [7:0] add_545336;
  wire [7:0] sel_545337;
  wire [7:0] add_545340;
  wire [7:0] sel_545341;
  wire [7:0] add_545344;
  wire [7:0] sel_545345;
  wire [7:0] add_545348;
  wire [7:0] sel_545349;
  wire [7:0] add_545352;
  wire [7:0] sel_545353;
  wire [7:0] add_545356;
  wire [7:0] sel_545357;
  wire [7:0] add_545360;
  wire [7:0] sel_545361;
  wire [7:0] add_545364;
  wire [7:0] sel_545365;
  wire [7:0] add_545368;
  wire [7:0] sel_545369;
  wire [7:0] add_545372;
  wire [7:0] sel_545373;
  wire [7:0] add_545376;
  wire [7:0] sel_545377;
  wire [7:0] add_545380;
  wire [7:0] sel_545381;
  wire [7:0] add_545384;
  wire [7:0] sel_545385;
  wire [7:0] add_545388;
  wire [7:0] sel_545389;
  wire [7:0] add_545392;
  wire [7:0] sel_545393;
  wire [7:0] add_545396;
  wire [7:0] sel_545397;
  wire [7:0] add_545400;
  wire [7:0] sel_545401;
  wire [7:0] add_545404;
  wire [7:0] sel_545405;
  wire [7:0] add_545408;
  wire [7:0] sel_545409;
  wire [7:0] add_545412;
  wire [7:0] sel_545413;
  wire [7:0] add_545416;
  wire [7:0] sel_545417;
  wire [7:0] add_545420;
  wire [7:0] sel_545421;
  wire [7:0] add_545424;
  wire [7:0] sel_545425;
  wire [7:0] add_545428;
  wire [7:0] sel_545429;
  wire [7:0] add_545432;
  wire [7:0] sel_545433;
  wire [7:0] add_545436;
  wire [7:0] sel_545437;
  wire [7:0] add_545440;
  wire [7:0] sel_545441;
  wire [7:0] add_545444;
  wire [7:0] sel_545445;
  wire [7:0] add_545448;
  wire [7:0] sel_545449;
  wire [7:0] add_545452;
  wire [7:0] sel_545453;
  wire [7:0] add_545456;
  wire [7:0] sel_545457;
  wire [7:0] add_545460;
  wire [7:0] sel_545461;
  wire [7:0] add_545464;
  wire [7:0] sel_545465;
  wire [7:0] add_545468;
  wire [7:0] sel_545469;
  wire [7:0] add_545472;
  wire [7:0] sel_545473;
  wire [7:0] add_545476;
  wire [7:0] sel_545477;
  wire [7:0] add_545480;
  wire [7:0] sel_545481;
  wire [7:0] add_545484;
  wire [7:0] sel_545485;
  wire [7:0] add_545488;
  wire [7:0] sel_545489;
  wire [7:0] add_545492;
  wire [7:0] sel_545493;
  wire [7:0] add_545496;
  wire [7:0] sel_545497;
  wire [7:0] add_545500;
  wire [7:0] sel_545501;
  wire [7:0] add_545504;
  wire [7:0] sel_545505;
  wire [7:0] add_545508;
  wire [7:0] sel_545509;
  wire [7:0] add_545512;
  wire [7:0] sel_545513;
  wire [7:0] add_545516;
  wire [7:0] sel_545517;
  wire [7:0] add_545520;
  wire [7:0] sel_545521;
  wire [7:0] add_545524;
  wire [7:0] sel_545525;
  wire [7:0] add_545528;
  wire [7:0] sel_545529;
  wire [7:0] add_545532;
  wire [7:0] sel_545533;
  wire [7:0] add_545536;
  wire [7:0] sel_545537;
  wire [7:0] add_545540;
  wire [7:0] sel_545541;
  wire [7:0] add_545544;
  wire [7:0] sel_545545;
  wire [7:0] add_545548;
  wire [7:0] sel_545549;
  wire [7:0] add_545552;
  wire [7:0] sel_545553;
  wire [7:0] add_545556;
  wire [7:0] sel_545557;
  wire [7:0] add_545560;
  wire [7:0] sel_545561;
  wire [7:0] add_545564;
  wire [7:0] sel_545565;
  wire [7:0] add_545568;
  wire [7:0] sel_545569;
  wire [7:0] add_545572;
  wire [7:0] sel_545573;
  wire [7:0] add_545576;
  wire [7:0] sel_545577;
  wire [7:0] add_545580;
  wire [7:0] sel_545581;
  wire [7:0] add_545584;
  wire [7:0] sel_545585;
  wire [7:0] add_545588;
  wire [7:0] sel_545589;
  wire [7:0] add_545592;
  wire [7:0] sel_545593;
  wire [7:0] add_545596;
  wire [7:0] sel_545597;
  wire [7:0] add_545600;
  wire [7:0] sel_545601;
  wire [7:0] add_545604;
  wire [7:0] sel_545605;
  wire [7:0] add_545608;
  wire [7:0] sel_545609;
  wire [7:0] add_545612;
  wire [7:0] sel_545613;
  wire [7:0] add_545616;
  wire [7:0] sel_545617;
  wire [7:0] add_545620;
  wire [7:0] sel_545621;
  wire [7:0] add_545625;
  wire [15:0] array_index_545626;
  wire [7:0] sel_545627;
  wire [7:0] add_545630;
  wire [7:0] sel_545631;
  wire [7:0] add_545634;
  wire [7:0] sel_545635;
  wire [7:0] add_545638;
  wire [7:0] sel_545639;
  wire [7:0] add_545642;
  wire [7:0] sel_545643;
  wire [7:0] add_545646;
  wire [7:0] sel_545647;
  wire [7:0] add_545650;
  wire [7:0] sel_545651;
  wire [7:0] add_545654;
  wire [7:0] sel_545655;
  wire [7:0] add_545658;
  wire [7:0] sel_545659;
  wire [7:0] add_545662;
  wire [7:0] sel_545663;
  wire [7:0] add_545666;
  wire [7:0] sel_545667;
  wire [7:0] add_545670;
  wire [7:0] sel_545671;
  wire [7:0] add_545674;
  wire [7:0] sel_545675;
  wire [7:0] add_545678;
  wire [7:0] sel_545679;
  wire [7:0] add_545682;
  wire [7:0] sel_545683;
  wire [7:0] add_545686;
  wire [7:0] sel_545687;
  wire [7:0] add_545690;
  wire [7:0] sel_545691;
  wire [7:0] add_545694;
  wire [7:0] sel_545695;
  wire [7:0] add_545698;
  wire [7:0] sel_545699;
  wire [7:0] add_545702;
  wire [7:0] sel_545703;
  wire [7:0] add_545706;
  wire [7:0] sel_545707;
  wire [7:0] add_545710;
  wire [7:0] sel_545711;
  wire [7:0] add_545714;
  wire [7:0] sel_545715;
  wire [7:0] add_545718;
  wire [7:0] sel_545719;
  wire [7:0] add_545722;
  wire [7:0] sel_545723;
  wire [7:0] add_545726;
  wire [7:0] sel_545727;
  wire [7:0] add_545730;
  wire [7:0] sel_545731;
  wire [7:0] add_545734;
  wire [7:0] sel_545735;
  wire [7:0] add_545738;
  wire [7:0] sel_545739;
  wire [7:0] add_545742;
  wire [7:0] sel_545743;
  wire [7:0] add_545746;
  wire [7:0] sel_545747;
  wire [7:0] add_545750;
  wire [7:0] sel_545751;
  wire [7:0] add_545754;
  wire [7:0] sel_545755;
  wire [7:0] add_545758;
  wire [7:0] sel_545759;
  wire [7:0] add_545762;
  wire [7:0] sel_545763;
  wire [7:0] add_545766;
  wire [7:0] sel_545767;
  wire [7:0] add_545770;
  wire [7:0] sel_545771;
  wire [7:0] add_545774;
  wire [7:0] sel_545775;
  wire [7:0] add_545778;
  wire [7:0] sel_545779;
  wire [7:0] add_545782;
  wire [7:0] sel_545783;
  wire [7:0] add_545786;
  wire [7:0] sel_545787;
  wire [7:0] add_545790;
  wire [7:0] sel_545791;
  wire [7:0] add_545794;
  wire [7:0] sel_545795;
  wire [7:0] add_545798;
  wire [7:0] sel_545799;
  wire [7:0] add_545802;
  wire [7:0] sel_545803;
  wire [7:0] add_545806;
  wire [7:0] sel_545807;
  wire [7:0] add_545810;
  wire [7:0] sel_545811;
  wire [7:0] add_545814;
  wire [7:0] sel_545815;
  wire [7:0] add_545818;
  wire [7:0] sel_545819;
  wire [7:0] add_545822;
  wire [7:0] sel_545823;
  wire [7:0] add_545826;
  wire [7:0] sel_545827;
  wire [7:0] add_545830;
  wire [7:0] sel_545831;
  wire [7:0] add_545834;
  wire [7:0] sel_545835;
  wire [7:0] add_545838;
  wire [7:0] sel_545839;
  wire [7:0] add_545842;
  wire [7:0] sel_545843;
  wire [7:0] add_545846;
  wire [7:0] sel_545847;
  wire [7:0] add_545850;
  wire [7:0] sel_545851;
  wire [7:0] add_545854;
  wire [7:0] sel_545855;
  wire [7:0] add_545858;
  wire [7:0] sel_545859;
  wire [7:0] add_545862;
  wire [7:0] sel_545863;
  wire [7:0] add_545866;
  wire [7:0] sel_545867;
  wire [7:0] add_545870;
  wire [7:0] sel_545871;
  wire [7:0] add_545874;
  wire [7:0] sel_545875;
  wire [7:0] add_545878;
  wire [7:0] sel_545879;
  wire [7:0] add_545882;
  wire [7:0] sel_545883;
  wire [7:0] add_545886;
  wire [7:0] sel_545887;
  wire [7:0] add_545890;
  wire [7:0] sel_545891;
  wire [7:0] add_545894;
  wire [7:0] sel_545895;
  wire [7:0] add_545898;
  wire [7:0] sel_545899;
  wire [7:0] add_545902;
  wire [7:0] sel_545903;
  wire [7:0] add_545906;
  wire [7:0] sel_545907;
  wire [7:0] add_545910;
  wire [7:0] sel_545911;
  wire [7:0] add_545914;
  wire [7:0] sel_545915;
  wire [7:0] add_545918;
  wire [7:0] sel_545919;
  wire [7:0] add_545922;
  wire [7:0] sel_545923;
  wire [7:0] add_545927;
  wire [15:0] array_index_545928;
  wire [7:0] sel_545929;
  wire [7:0] add_545932;
  wire [7:0] sel_545933;
  wire [7:0] add_545936;
  wire [7:0] sel_545937;
  wire [7:0] add_545940;
  wire [7:0] sel_545941;
  wire [7:0] add_545944;
  wire [7:0] sel_545945;
  wire [7:0] add_545948;
  wire [7:0] sel_545949;
  wire [7:0] add_545952;
  wire [7:0] sel_545953;
  wire [7:0] add_545956;
  wire [7:0] sel_545957;
  wire [7:0] add_545960;
  wire [7:0] sel_545961;
  wire [7:0] add_545964;
  wire [7:0] sel_545965;
  wire [7:0] add_545968;
  wire [7:0] sel_545969;
  wire [7:0] add_545972;
  wire [7:0] sel_545973;
  wire [7:0] add_545976;
  wire [7:0] sel_545977;
  wire [7:0] add_545980;
  wire [7:0] sel_545981;
  wire [7:0] add_545984;
  wire [7:0] sel_545985;
  wire [7:0] add_545988;
  wire [7:0] sel_545989;
  wire [7:0] add_545992;
  wire [7:0] sel_545993;
  wire [7:0] add_545996;
  wire [7:0] sel_545997;
  wire [7:0] add_546000;
  wire [7:0] sel_546001;
  wire [7:0] add_546004;
  wire [7:0] sel_546005;
  wire [7:0] add_546008;
  wire [7:0] sel_546009;
  wire [7:0] add_546012;
  wire [7:0] sel_546013;
  wire [7:0] add_546016;
  wire [7:0] sel_546017;
  wire [7:0] add_546020;
  wire [7:0] sel_546021;
  wire [7:0] add_546024;
  wire [7:0] sel_546025;
  wire [7:0] add_546028;
  wire [7:0] sel_546029;
  wire [7:0] add_546032;
  wire [7:0] sel_546033;
  wire [7:0] add_546036;
  wire [7:0] sel_546037;
  wire [7:0] add_546040;
  wire [7:0] sel_546041;
  wire [7:0] add_546044;
  wire [7:0] sel_546045;
  wire [7:0] add_546048;
  wire [7:0] sel_546049;
  wire [7:0] add_546052;
  wire [7:0] sel_546053;
  wire [7:0] add_546056;
  wire [7:0] sel_546057;
  wire [7:0] add_546060;
  wire [7:0] sel_546061;
  wire [7:0] add_546064;
  wire [7:0] sel_546065;
  wire [7:0] add_546068;
  wire [7:0] sel_546069;
  wire [7:0] add_546072;
  wire [7:0] sel_546073;
  wire [7:0] add_546076;
  wire [7:0] sel_546077;
  wire [7:0] add_546080;
  wire [7:0] sel_546081;
  wire [7:0] add_546084;
  wire [7:0] sel_546085;
  wire [7:0] add_546088;
  wire [7:0] sel_546089;
  wire [7:0] add_546092;
  wire [7:0] sel_546093;
  wire [7:0] add_546096;
  wire [7:0] sel_546097;
  wire [7:0] add_546100;
  wire [7:0] sel_546101;
  wire [7:0] add_546104;
  wire [7:0] sel_546105;
  wire [7:0] add_546108;
  wire [7:0] sel_546109;
  wire [7:0] add_546112;
  wire [7:0] sel_546113;
  wire [7:0] add_546116;
  wire [7:0] sel_546117;
  wire [7:0] add_546120;
  wire [7:0] sel_546121;
  wire [7:0] add_546124;
  wire [7:0] sel_546125;
  wire [7:0] add_546128;
  wire [7:0] sel_546129;
  wire [7:0] add_546132;
  wire [7:0] sel_546133;
  wire [7:0] add_546136;
  wire [7:0] sel_546137;
  wire [7:0] add_546140;
  wire [7:0] sel_546141;
  wire [7:0] add_546144;
  wire [7:0] sel_546145;
  wire [7:0] add_546148;
  wire [7:0] sel_546149;
  wire [7:0] add_546152;
  wire [7:0] sel_546153;
  wire [7:0] add_546156;
  wire [7:0] sel_546157;
  wire [7:0] add_546160;
  wire [7:0] sel_546161;
  wire [7:0] add_546164;
  wire [7:0] sel_546165;
  wire [7:0] add_546168;
  wire [7:0] sel_546169;
  wire [7:0] add_546172;
  wire [7:0] sel_546173;
  wire [7:0] add_546176;
  wire [7:0] sel_546177;
  wire [7:0] add_546180;
  wire [7:0] sel_546181;
  wire [7:0] add_546184;
  wire [7:0] sel_546185;
  wire [7:0] add_546188;
  wire [7:0] sel_546189;
  wire [7:0] add_546192;
  wire [7:0] sel_546193;
  wire [7:0] add_546196;
  wire [7:0] sel_546197;
  wire [7:0] add_546200;
  wire [7:0] sel_546201;
  wire [7:0] add_546204;
  wire [7:0] sel_546205;
  wire [7:0] add_546208;
  wire [7:0] sel_546209;
  wire [7:0] add_546212;
  wire [7:0] sel_546213;
  wire [7:0] add_546216;
  wire [7:0] sel_546217;
  wire [7:0] add_546220;
  wire [7:0] sel_546221;
  wire [7:0] add_546224;
  wire [7:0] sel_546225;
  wire [7:0] add_546229;
  wire [15:0] array_index_546230;
  wire [7:0] sel_546231;
  wire [7:0] add_546234;
  wire [7:0] sel_546235;
  wire [7:0] add_546238;
  wire [7:0] sel_546239;
  wire [7:0] add_546242;
  wire [7:0] sel_546243;
  wire [7:0] add_546246;
  wire [7:0] sel_546247;
  wire [7:0] add_546250;
  wire [7:0] sel_546251;
  wire [7:0] add_546254;
  wire [7:0] sel_546255;
  wire [7:0] add_546258;
  wire [7:0] sel_546259;
  wire [7:0] add_546262;
  wire [7:0] sel_546263;
  wire [7:0] add_546266;
  wire [7:0] sel_546267;
  wire [7:0] add_546270;
  wire [7:0] sel_546271;
  wire [7:0] add_546274;
  wire [7:0] sel_546275;
  wire [7:0] add_546278;
  wire [7:0] sel_546279;
  wire [7:0] add_546282;
  wire [7:0] sel_546283;
  wire [7:0] add_546286;
  wire [7:0] sel_546287;
  wire [7:0] add_546290;
  wire [7:0] sel_546291;
  wire [7:0] add_546294;
  wire [7:0] sel_546295;
  wire [7:0] add_546298;
  wire [7:0] sel_546299;
  wire [7:0] add_546302;
  wire [7:0] sel_546303;
  wire [7:0] add_546306;
  wire [7:0] sel_546307;
  wire [7:0] add_546310;
  wire [7:0] sel_546311;
  wire [7:0] add_546314;
  wire [7:0] sel_546315;
  wire [7:0] add_546318;
  wire [7:0] sel_546319;
  wire [7:0] add_546322;
  wire [7:0] sel_546323;
  wire [7:0] add_546326;
  wire [7:0] sel_546327;
  wire [7:0] add_546330;
  wire [7:0] sel_546331;
  wire [7:0] add_546334;
  wire [7:0] sel_546335;
  wire [7:0] add_546338;
  wire [7:0] sel_546339;
  wire [7:0] add_546342;
  wire [7:0] sel_546343;
  wire [7:0] add_546346;
  wire [7:0] sel_546347;
  wire [7:0] add_546350;
  wire [7:0] sel_546351;
  wire [7:0] add_546354;
  wire [7:0] sel_546355;
  wire [7:0] add_546358;
  wire [7:0] sel_546359;
  wire [7:0] add_546362;
  wire [7:0] sel_546363;
  wire [7:0] add_546366;
  wire [7:0] sel_546367;
  wire [7:0] add_546370;
  wire [7:0] sel_546371;
  wire [7:0] add_546374;
  wire [7:0] sel_546375;
  wire [7:0] add_546378;
  wire [7:0] sel_546379;
  wire [7:0] add_546382;
  wire [7:0] sel_546383;
  wire [7:0] add_546386;
  wire [7:0] sel_546387;
  wire [7:0] add_546390;
  wire [7:0] sel_546391;
  wire [7:0] add_546394;
  wire [7:0] sel_546395;
  wire [7:0] add_546398;
  wire [7:0] sel_546399;
  wire [7:0] add_546402;
  wire [7:0] sel_546403;
  wire [7:0] add_546406;
  wire [7:0] sel_546407;
  wire [7:0] add_546410;
  wire [7:0] sel_546411;
  wire [7:0] add_546414;
  wire [7:0] sel_546415;
  wire [7:0] add_546418;
  wire [7:0] sel_546419;
  wire [7:0] add_546422;
  wire [7:0] sel_546423;
  wire [7:0] add_546426;
  wire [7:0] sel_546427;
  wire [7:0] add_546430;
  wire [7:0] sel_546431;
  wire [7:0] add_546434;
  wire [7:0] sel_546435;
  wire [7:0] add_546438;
  wire [7:0] sel_546439;
  wire [7:0] add_546442;
  wire [7:0] sel_546443;
  wire [7:0] add_546446;
  wire [7:0] sel_546447;
  wire [7:0] add_546450;
  wire [7:0] sel_546451;
  wire [7:0] add_546454;
  wire [7:0] sel_546455;
  wire [7:0] add_546458;
  wire [7:0] sel_546459;
  wire [7:0] add_546462;
  wire [7:0] sel_546463;
  wire [7:0] add_546466;
  wire [7:0] sel_546467;
  wire [7:0] add_546470;
  wire [7:0] sel_546471;
  wire [7:0] add_546474;
  wire [7:0] sel_546475;
  wire [7:0] add_546478;
  wire [7:0] sel_546479;
  wire [7:0] add_546482;
  wire [7:0] sel_546483;
  wire [7:0] add_546486;
  wire [7:0] sel_546487;
  wire [7:0] add_546490;
  wire [7:0] sel_546491;
  wire [7:0] add_546494;
  wire [7:0] sel_546495;
  wire [7:0] add_546498;
  wire [7:0] sel_546499;
  wire [7:0] add_546502;
  wire [7:0] sel_546503;
  wire [7:0] add_546506;
  wire [7:0] sel_546507;
  wire [7:0] add_546510;
  wire [7:0] sel_546511;
  wire [7:0] add_546514;
  wire [7:0] sel_546515;
  wire [7:0] add_546518;
  wire [7:0] sel_546519;
  wire [7:0] add_546522;
  wire [7:0] sel_546523;
  wire [7:0] add_546526;
  wire [7:0] sel_546527;
  wire [7:0] add_546531;
  wire [15:0] array_index_546532;
  wire [7:0] sel_546533;
  wire [7:0] add_546536;
  wire [7:0] sel_546537;
  wire [7:0] add_546540;
  wire [7:0] sel_546541;
  wire [7:0] add_546544;
  wire [7:0] sel_546545;
  wire [7:0] add_546548;
  wire [7:0] sel_546549;
  wire [7:0] add_546552;
  wire [7:0] sel_546553;
  wire [7:0] add_546556;
  wire [7:0] sel_546557;
  wire [7:0] add_546560;
  wire [7:0] sel_546561;
  wire [7:0] add_546564;
  wire [7:0] sel_546565;
  wire [7:0] add_546568;
  wire [7:0] sel_546569;
  wire [7:0] add_546572;
  wire [7:0] sel_546573;
  wire [7:0] add_546576;
  wire [7:0] sel_546577;
  wire [7:0] add_546580;
  wire [7:0] sel_546581;
  wire [7:0] add_546584;
  wire [7:0] sel_546585;
  wire [7:0] add_546588;
  wire [7:0] sel_546589;
  wire [7:0] add_546592;
  wire [7:0] sel_546593;
  wire [7:0] add_546596;
  wire [7:0] sel_546597;
  wire [7:0] add_546600;
  wire [7:0] sel_546601;
  wire [7:0] add_546604;
  wire [7:0] sel_546605;
  wire [7:0] add_546608;
  wire [7:0] sel_546609;
  wire [7:0] add_546612;
  wire [7:0] sel_546613;
  wire [7:0] add_546616;
  wire [7:0] sel_546617;
  wire [7:0] add_546620;
  wire [7:0] sel_546621;
  wire [7:0] add_546624;
  wire [7:0] sel_546625;
  wire [7:0] add_546628;
  wire [7:0] sel_546629;
  wire [7:0] add_546632;
  wire [7:0] sel_546633;
  wire [7:0] add_546636;
  wire [7:0] sel_546637;
  wire [7:0] add_546640;
  wire [7:0] sel_546641;
  wire [7:0] add_546644;
  wire [7:0] sel_546645;
  wire [7:0] add_546648;
  wire [7:0] sel_546649;
  wire [7:0] add_546652;
  wire [7:0] sel_546653;
  wire [7:0] add_546656;
  wire [7:0] sel_546657;
  wire [7:0] add_546660;
  wire [7:0] sel_546661;
  wire [7:0] add_546664;
  wire [7:0] sel_546665;
  wire [7:0] add_546668;
  wire [7:0] sel_546669;
  wire [7:0] add_546672;
  wire [7:0] sel_546673;
  wire [7:0] add_546676;
  wire [7:0] sel_546677;
  wire [7:0] add_546680;
  wire [7:0] sel_546681;
  wire [7:0] add_546684;
  wire [7:0] sel_546685;
  wire [7:0] add_546688;
  wire [7:0] sel_546689;
  wire [7:0] add_546692;
  wire [7:0] sel_546693;
  wire [7:0] add_546696;
  wire [7:0] sel_546697;
  wire [7:0] add_546700;
  wire [7:0] sel_546701;
  wire [7:0] add_546704;
  wire [7:0] sel_546705;
  wire [7:0] add_546708;
  wire [7:0] sel_546709;
  wire [7:0] add_546712;
  wire [7:0] sel_546713;
  wire [7:0] add_546716;
  wire [7:0] sel_546717;
  wire [7:0] add_546720;
  wire [7:0] sel_546721;
  wire [7:0] add_546724;
  wire [7:0] sel_546725;
  wire [7:0] add_546728;
  wire [7:0] sel_546729;
  wire [7:0] add_546732;
  wire [7:0] sel_546733;
  wire [7:0] add_546736;
  wire [7:0] sel_546737;
  wire [7:0] add_546740;
  wire [7:0] sel_546741;
  wire [7:0] add_546744;
  wire [7:0] sel_546745;
  wire [7:0] add_546748;
  wire [7:0] sel_546749;
  wire [7:0] add_546752;
  wire [7:0] sel_546753;
  wire [7:0] add_546756;
  wire [7:0] sel_546757;
  wire [7:0] add_546760;
  wire [7:0] sel_546761;
  wire [7:0] add_546764;
  wire [7:0] sel_546765;
  wire [7:0] add_546768;
  wire [7:0] sel_546769;
  wire [7:0] add_546772;
  wire [7:0] sel_546773;
  wire [7:0] add_546776;
  wire [7:0] sel_546777;
  wire [7:0] add_546780;
  wire [7:0] sel_546781;
  wire [7:0] add_546784;
  wire [7:0] sel_546785;
  wire [7:0] add_546788;
  wire [7:0] sel_546789;
  wire [7:0] add_546792;
  wire [7:0] sel_546793;
  wire [7:0] add_546796;
  wire [7:0] sel_546797;
  wire [7:0] add_546800;
  wire [7:0] sel_546801;
  wire [7:0] add_546804;
  wire [7:0] sel_546805;
  wire [7:0] add_546808;
  wire [7:0] sel_546809;
  wire [7:0] add_546812;
  wire [7:0] sel_546813;
  wire [7:0] add_546816;
  wire [7:0] sel_546817;
  wire [7:0] add_546820;
  wire [7:0] sel_546821;
  wire [7:0] add_546824;
  wire [7:0] sel_546825;
  wire [7:0] add_546828;
  wire [7:0] sel_546829;
  wire [7:0] add_546833;
  wire [15:0] array_index_546834;
  wire [7:0] sel_546835;
  wire [7:0] add_546838;
  wire [7:0] sel_546839;
  wire [7:0] add_546842;
  wire [7:0] sel_546843;
  wire [7:0] add_546846;
  wire [7:0] sel_546847;
  wire [7:0] add_546850;
  wire [7:0] sel_546851;
  wire [7:0] add_546854;
  wire [7:0] sel_546855;
  wire [7:0] add_546858;
  wire [7:0] sel_546859;
  wire [7:0] add_546862;
  wire [7:0] sel_546863;
  wire [7:0] add_546866;
  wire [7:0] sel_546867;
  wire [7:0] add_546870;
  wire [7:0] sel_546871;
  wire [7:0] add_546874;
  wire [7:0] sel_546875;
  wire [7:0] add_546878;
  wire [7:0] sel_546879;
  wire [7:0] add_546882;
  wire [7:0] sel_546883;
  wire [7:0] add_546886;
  wire [7:0] sel_546887;
  wire [7:0] add_546890;
  wire [7:0] sel_546891;
  wire [7:0] add_546894;
  wire [7:0] sel_546895;
  wire [7:0] add_546898;
  wire [7:0] sel_546899;
  wire [7:0] add_546902;
  wire [7:0] sel_546903;
  wire [7:0] add_546906;
  wire [7:0] sel_546907;
  wire [7:0] add_546910;
  wire [7:0] sel_546911;
  wire [7:0] add_546914;
  wire [7:0] sel_546915;
  wire [7:0] add_546918;
  wire [7:0] sel_546919;
  wire [7:0] add_546922;
  wire [7:0] sel_546923;
  wire [7:0] add_546926;
  wire [7:0] sel_546927;
  wire [7:0] add_546930;
  wire [7:0] sel_546931;
  wire [7:0] add_546934;
  wire [7:0] sel_546935;
  wire [7:0] add_546938;
  wire [7:0] sel_546939;
  wire [7:0] add_546942;
  wire [7:0] sel_546943;
  wire [7:0] add_546946;
  wire [7:0] sel_546947;
  wire [7:0] add_546950;
  wire [7:0] sel_546951;
  wire [7:0] add_546954;
  wire [7:0] sel_546955;
  wire [7:0] add_546958;
  wire [7:0] sel_546959;
  wire [7:0] add_546962;
  wire [7:0] sel_546963;
  wire [7:0] add_546966;
  wire [7:0] sel_546967;
  wire [7:0] add_546970;
  wire [7:0] sel_546971;
  wire [7:0] add_546974;
  wire [7:0] sel_546975;
  wire [7:0] add_546978;
  wire [7:0] sel_546979;
  wire [7:0] add_546982;
  wire [7:0] sel_546983;
  wire [7:0] add_546986;
  wire [7:0] sel_546987;
  wire [7:0] add_546990;
  wire [7:0] sel_546991;
  wire [7:0] add_546994;
  wire [7:0] sel_546995;
  wire [7:0] add_546998;
  wire [7:0] sel_546999;
  wire [7:0] add_547002;
  wire [7:0] sel_547003;
  wire [7:0] add_547006;
  wire [7:0] sel_547007;
  wire [7:0] add_547010;
  wire [7:0] sel_547011;
  wire [7:0] add_547014;
  wire [7:0] sel_547015;
  wire [7:0] add_547018;
  wire [7:0] sel_547019;
  wire [7:0] add_547022;
  wire [7:0] sel_547023;
  wire [7:0] add_547026;
  wire [7:0] sel_547027;
  wire [7:0] add_547030;
  wire [7:0] sel_547031;
  wire [7:0] add_547034;
  wire [7:0] sel_547035;
  wire [7:0] add_547038;
  wire [7:0] sel_547039;
  wire [7:0] add_547042;
  wire [7:0] sel_547043;
  wire [7:0] add_547046;
  wire [7:0] sel_547047;
  wire [7:0] add_547050;
  wire [7:0] sel_547051;
  wire [7:0] add_547054;
  wire [7:0] sel_547055;
  wire [7:0] add_547058;
  wire [7:0] sel_547059;
  wire [7:0] add_547062;
  wire [7:0] sel_547063;
  wire [7:0] add_547066;
  wire [7:0] sel_547067;
  wire [7:0] add_547070;
  wire [7:0] sel_547071;
  wire [7:0] add_547074;
  wire [7:0] sel_547075;
  wire [7:0] add_547078;
  wire [7:0] sel_547079;
  wire [7:0] add_547082;
  wire [7:0] sel_547083;
  wire [7:0] add_547086;
  wire [7:0] sel_547087;
  wire [7:0] add_547090;
  wire [7:0] sel_547091;
  wire [7:0] add_547094;
  wire [7:0] sel_547095;
  wire [7:0] add_547098;
  wire [7:0] sel_547099;
  wire [7:0] add_547102;
  wire [7:0] sel_547103;
  wire [7:0] add_547106;
  wire [7:0] sel_547107;
  wire [7:0] add_547110;
  wire [7:0] sel_547111;
  wire [7:0] add_547114;
  wire [7:0] sel_547115;
  wire [7:0] add_547118;
  wire [7:0] sel_547119;
  wire [7:0] add_547122;
  wire [7:0] sel_547123;
  wire [7:0] add_547126;
  wire [7:0] sel_547127;
  wire [7:0] add_547130;
  wire [7:0] sel_547131;
  wire [7:0] add_547135;
  wire [15:0] array_index_547136;
  wire [7:0] sel_547137;
  wire [7:0] add_547140;
  wire [7:0] sel_547141;
  wire [7:0] add_547144;
  wire [7:0] sel_547145;
  wire [7:0] add_547148;
  wire [7:0] sel_547149;
  wire [7:0] add_547152;
  wire [7:0] sel_547153;
  wire [7:0] add_547156;
  wire [7:0] sel_547157;
  wire [7:0] add_547160;
  wire [7:0] sel_547161;
  wire [7:0] add_547164;
  wire [7:0] sel_547165;
  wire [7:0] add_547168;
  wire [7:0] sel_547169;
  wire [7:0] add_547172;
  wire [7:0] sel_547173;
  wire [7:0] add_547176;
  wire [7:0] sel_547177;
  wire [7:0] add_547180;
  wire [7:0] sel_547181;
  wire [7:0] add_547184;
  wire [7:0] sel_547185;
  wire [7:0] add_547188;
  wire [7:0] sel_547189;
  wire [7:0] add_547192;
  wire [7:0] sel_547193;
  wire [7:0] add_547196;
  wire [7:0] sel_547197;
  wire [7:0] add_547200;
  wire [7:0] sel_547201;
  wire [7:0] add_547204;
  wire [7:0] sel_547205;
  wire [7:0] add_547208;
  wire [7:0] sel_547209;
  wire [7:0] add_547212;
  wire [7:0] sel_547213;
  wire [7:0] add_547216;
  wire [7:0] sel_547217;
  wire [7:0] add_547220;
  wire [7:0] sel_547221;
  wire [7:0] add_547224;
  wire [7:0] sel_547225;
  wire [7:0] add_547228;
  wire [7:0] sel_547229;
  wire [7:0] add_547232;
  wire [7:0] sel_547233;
  wire [7:0] add_547236;
  wire [7:0] sel_547237;
  wire [7:0] add_547240;
  wire [7:0] sel_547241;
  wire [7:0] add_547244;
  wire [7:0] sel_547245;
  wire [7:0] add_547248;
  wire [7:0] sel_547249;
  wire [7:0] add_547252;
  wire [7:0] sel_547253;
  wire [7:0] add_547256;
  wire [7:0] sel_547257;
  wire [7:0] add_547260;
  wire [7:0] sel_547261;
  wire [7:0] add_547264;
  wire [7:0] sel_547265;
  wire [7:0] add_547268;
  wire [7:0] sel_547269;
  wire [7:0] add_547272;
  wire [7:0] sel_547273;
  wire [7:0] add_547276;
  wire [7:0] sel_547277;
  wire [7:0] add_547280;
  wire [7:0] sel_547281;
  wire [7:0] add_547284;
  wire [7:0] sel_547285;
  wire [7:0] add_547288;
  wire [7:0] sel_547289;
  wire [7:0] add_547292;
  wire [7:0] sel_547293;
  wire [7:0] add_547296;
  wire [7:0] sel_547297;
  wire [7:0] add_547300;
  wire [7:0] sel_547301;
  wire [7:0] add_547304;
  wire [7:0] sel_547305;
  wire [7:0] add_547308;
  wire [7:0] sel_547309;
  wire [7:0] add_547312;
  wire [7:0] sel_547313;
  wire [7:0] add_547316;
  wire [7:0] sel_547317;
  wire [7:0] add_547320;
  wire [7:0] sel_547321;
  wire [7:0] add_547324;
  wire [7:0] sel_547325;
  wire [7:0] add_547328;
  wire [7:0] sel_547329;
  wire [7:0] add_547332;
  wire [7:0] sel_547333;
  wire [7:0] add_547336;
  wire [7:0] sel_547337;
  wire [7:0] add_547340;
  wire [7:0] sel_547341;
  wire [7:0] add_547344;
  wire [7:0] sel_547345;
  wire [7:0] add_547348;
  wire [7:0] sel_547349;
  wire [7:0] add_547352;
  wire [7:0] sel_547353;
  wire [7:0] add_547356;
  wire [7:0] sel_547357;
  wire [7:0] add_547360;
  wire [7:0] sel_547361;
  wire [7:0] add_547364;
  wire [7:0] sel_547365;
  wire [7:0] add_547368;
  wire [7:0] sel_547369;
  wire [7:0] add_547372;
  wire [7:0] sel_547373;
  wire [7:0] add_547376;
  wire [7:0] sel_547377;
  wire [7:0] add_547380;
  wire [7:0] sel_547381;
  wire [7:0] add_547384;
  wire [7:0] sel_547385;
  wire [7:0] add_547388;
  wire [7:0] sel_547389;
  wire [7:0] add_547392;
  wire [7:0] sel_547393;
  wire [7:0] add_547396;
  wire [7:0] sel_547397;
  wire [7:0] add_547400;
  wire [7:0] sel_547401;
  wire [7:0] add_547404;
  wire [7:0] sel_547405;
  wire [7:0] add_547408;
  wire [7:0] sel_547409;
  wire [7:0] add_547412;
  wire [7:0] sel_547413;
  wire [7:0] add_547416;
  wire [7:0] sel_547417;
  wire [7:0] add_547420;
  wire [7:0] sel_547421;
  wire [7:0] add_547424;
  wire [7:0] sel_547425;
  wire [7:0] add_547428;
  wire [7:0] sel_547429;
  wire [7:0] add_547432;
  wire [7:0] sel_547433;
  wire [7:0] add_547437;
  wire [15:0] array_index_547438;
  wire [7:0] sel_547439;
  wire [7:0] add_547442;
  wire [7:0] sel_547443;
  wire [7:0] add_547446;
  wire [7:0] sel_547447;
  wire [7:0] add_547450;
  wire [7:0] sel_547451;
  wire [7:0] add_547454;
  wire [7:0] sel_547455;
  wire [7:0] add_547458;
  wire [7:0] sel_547459;
  wire [7:0] add_547462;
  wire [7:0] sel_547463;
  wire [7:0] add_547466;
  wire [7:0] sel_547467;
  wire [7:0] add_547470;
  wire [7:0] sel_547471;
  wire [7:0] add_547474;
  wire [7:0] sel_547475;
  wire [7:0] add_547478;
  wire [7:0] sel_547479;
  wire [7:0] add_547482;
  wire [7:0] sel_547483;
  wire [7:0] add_547486;
  wire [7:0] sel_547487;
  wire [7:0] add_547490;
  wire [7:0] sel_547491;
  wire [7:0] add_547494;
  wire [7:0] sel_547495;
  wire [7:0] add_547498;
  wire [7:0] sel_547499;
  wire [7:0] add_547502;
  wire [7:0] sel_547503;
  wire [7:0] add_547506;
  wire [7:0] sel_547507;
  wire [7:0] add_547510;
  wire [7:0] sel_547511;
  wire [7:0] add_547514;
  wire [7:0] sel_547515;
  wire [7:0] add_547518;
  wire [7:0] sel_547519;
  wire [7:0] add_547522;
  wire [7:0] sel_547523;
  wire [7:0] add_547526;
  wire [7:0] sel_547527;
  wire [7:0] add_547530;
  wire [7:0] sel_547531;
  wire [7:0] add_547534;
  wire [7:0] sel_547535;
  wire [7:0] add_547538;
  wire [7:0] sel_547539;
  wire [7:0] add_547542;
  wire [7:0] sel_547543;
  wire [7:0] add_547546;
  wire [7:0] sel_547547;
  wire [7:0] add_547550;
  wire [7:0] sel_547551;
  wire [7:0] add_547554;
  wire [7:0] sel_547555;
  wire [7:0] add_547558;
  wire [7:0] sel_547559;
  wire [7:0] add_547562;
  wire [7:0] sel_547563;
  wire [7:0] add_547566;
  wire [7:0] sel_547567;
  wire [7:0] add_547570;
  wire [7:0] sel_547571;
  wire [7:0] add_547574;
  wire [7:0] sel_547575;
  wire [7:0] add_547578;
  wire [7:0] sel_547579;
  wire [7:0] add_547582;
  wire [7:0] sel_547583;
  wire [7:0] add_547586;
  wire [7:0] sel_547587;
  wire [7:0] add_547590;
  wire [7:0] sel_547591;
  wire [7:0] add_547594;
  wire [7:0] sel_547595;
  wire [7:0] add_547598;
  wire [7:0] sel_547599;
  wire [7:0] add_547602;
  wire [7:0] sel_547603;
  wire [7:0] add_547606;
  wire [7:0] sel_547607;
  wire [7:0] add_547610;
  wire [7:0] sel_547611;
  wire [7:0] add_547614;
  wire [7:0] sel_547615;
  wire [7:0] add_547618;
  wire [7:0] sel_547619;
  wire [7:0] add_547622;
  wire [7:0] sel_547623;
  wire [7:0] add_547626;
  wire [7:0] sel_547627;
  wire [7:0] add_547630;
  wire [7:0] sel_547631;
  wire [7:0] add_547634;
  wire [7:0] sel_547635;
  wire [7:0] add_547638;
  wire [7:0] sel_547639;
  wire [7:0] add_547642;
  wire [7:0] sel_547643;
  wire [7:0] add_547646;
  wire [7:0] sel_547647;
  wire [7:0] add_547650;
  wire [7:0] sel_547651;
  wire [7:0] add_547654;
  wire [7:0] sel_547655;
  wire [7:0] add_547658;
  wire [7:0] sel_547659;
  wire [7:0] add_547662;
  wire [7:0] sel_547663;
  wire [7:0] add_547666;
  wire [7:0] sel_547667;
  wire [7:0] add_547670;
  wire [7:0] sel_547671;
  wire [7:0] add_547674;
  wire [7:0] sel_547675;
  wire [7:0] add_547678;
  wire [7:0] sel_547679;
  wire [7:0] add_547682;
  wire [7:0] sel_547683;
  wire [7:0] add_547686;
  wire [7:0] sel_547687;
  wire [7:0] add_547690;
  wire [7:0] sel_547691;
  wire [7:0] add_547694;
  wire [7:0] sel_547695;
  wire [7:0] add_547698;
  wire [7:0] sel_547699;
  wire [7:0] add_547702;
  wire [7:0] sel_547703;
  wire [7:0] add_547706;
  wire [7:0] sel_547707;
  wire [7:0] add_547710;
  wire [7:0] sel_547711;
  wire [7:0] add_547714;
  wire [7:0] sel_547715;
  wire [7:0] add_547718;
  wire [7:0] sel_547719;
  wire [7:0] add_547722;
  wire [7:0] sel_547723;
  wire [7:0] add_547726;
  wire [7:0] sel_547727;
  wire [7:0] add_547730;
  wire [7:0] sel_547731;
  wire [7:0] add_547734;
  wire [7:0] sel_547735;
  wire [7:0] add_547739;
  wire [15:0] array_index_547740;
  wire [7:0] sel_547741;
  wire [7:0] add_547744;
  wire [7:0] sel_547745;
  wire [7:0] add_547748;
  wire [7:0] sel_547749;
  wire [7:0] add_547752;
  wire [7:0] sel_547753;
  wire [7:0] add_547756;
  wire [7:0] sel_547757;
  wire [7:0] add_547760;
  wire [7:0] sel_547761;
  wire [7:0] add_547764;
  wire [7:0] sel_547765;
  wire [7:0] add_547768;
  wire [7:0] sel_547769;
  wire [7:0] add_547772;
  wire [7:0] sel_547773;
  wire [7:0] add_547776;
  wire [7:0] sel_547777;
  wire [7:0] add_547780;
  wire [7:0] sel_547781;
  wire [7:0] add_547784;
  wire [7:0] sel_547785;
  wire [7:0] add_547788;
  wire [7:0] sel_547789;
  wire [7:0] add_547792;
  wire [7:0] sel_547793;
  wire [7:0] add_547796;
  wire [7:0] sel_547797;
  wire [7:0] add_547800;
  wire [7:0] sel_547801;
  wire [7:0] add_547804;
  wire [7:0] sel_547805;
  wire [7:0] add_547808;
  wire [7:0] sel_547809;
  wire [7:0] add_547812;
  wire [7:0] sel_547813;
  wire [7:0] add_547816;
  wire [7:0] sel_547817;
  wire [7:0] add_547820;
  wire [7:0] sel_547821;
  wire [7:0] add_547824;
  wire [7:0] sel_547825;
  wire [7:0] add_547828;
  wire [7:0] sel_547829;
  wire [7:0] add_547832;
  wire [7:0] sel_547833;
  wire [7:0] add_547836;
  wire [7:0] sel_547837;
  wire [7:0] add_547840;
  wire [7:0] sel_547841;
  wire [7:0] add_547844;
  wire [7:0] sel_547845;
  wire [7:0] add_547848;
  wire [7:0] sel_547849;
  wire [7:0] add_547852;
  wire [7:0] sel_547853;
  wire [7:0] add_547856;
  wire [7:0] sel_547857;
  wire [7:0] add_547860;
  wire [7:0] sel_547861;
  wire [7:0] add_547864;
  wire [7:0] sel_547865;
  wire [7:0] add_547868;
  wire [7:0] sel_547869;
  wire [7:0] add_547872;
  wire [7:0] sel_547873;
  wire [7:0] add_547876;
  wire [7:0] sel_547877;
  wire [7:0] add_547880;
  wire [7:0] sel_547881;
  wire [7:0] add_547884;
  wire [7:0] sel_547885;
  wire [7:0] add_547888;
  wire [7:0] sel_547889;
  wire [7:0] add_547892;
  wire [7:0] sel_547893;
  wire [7:0] add_547896;
  wire [7:0] sel_547897;
  wire [7:0] add_547900;
  wire [7:0] sel_547901;
  wire [7:0] add_547904;
  wire [7:0] sel_547905;
  wire [7:0] add_547908;
  wire [7:0] sel_547909;
  wire [7:0] add_547912;
  wire [7:0] sel_547913;
  wire [7:0] add_547916;
  wire [7:0] sel_547917;
  wire [7:0] add_547920;
  wire [7:0] sel_547921;
  wire [7:0] add_547924;
  wire [7:0] sel_547925;
  wire [7:0] add_547928;
  wire [7:0] sel_547929;
  wire [7:0] add_547932;
  wire [7:0] sel_547933;
  wire [7:0] add_547936;
  wire [7:0] sel_547937;
  wire [7:0] add_547940;
  wire [7:0] sel_547941;
  wire [7:0] add_547944;
  wire [7:0] sel_547945;
  wire [7:0] add_547948;
  wire [7:0] sel_547949;
  wire [7:0] add_547952;
  wire [7:0] sel_547953;
  wire [7:0] add_547956;
  wire [7:0] sel_547957;
  wire [7:0] add_547960;
  wire [7:0] sel_547961;
  wire [7:0] add_547964;
  wire [7:0] sel_547965;
  wire [7:0] add_547968;
  wire [7:0] sel_547969;
  wire [7:0] add_547972;
  wire [7:0] sel_547973;
  wire [7:0] add_547976;
  wire [7:0] sel_547977;
  wire [7:0] add_547980;
  wire [7:0] sel_547981;
  wire [7:0] add_547984;
  wire [7:0] sel_547985;
  wire [7:0] add_547988;
  wire [7:0] sel_547989;
  wire [7:0] add_547992;
  wire [7:0] sel_547993;
  wire [7:0] add_547996;
  wire [7:0] sel_547997;
  wire [7:0] add_548000;
  wire [7:0] sel_548001;
  wire [7:0] add_548004;
  wire [7:0] sel_548005;
  wire [7:0] add_548008;
  wire [7:0] sel_548009;
  wire [7:0] add_548012;
  wire [7:0] sel_548013;
  wire [7:0] add_548016;
  wire [7:0] sel_548017;
  wire [7:0] add_548020;
  wire [7:0] sel_548021;
  wire [7:0] add_548024;
  wire [7:0] sel_548025;
  wire [7:0] add_548028;
  wire [7:0] sel_548029;
  wire [7:0] add_548032;
  wire [7:0] sel_548033;
  wire [7:0] add_548036;
  wire [7:0] sel_548037;
  wire [7:0] add_548041;
  wire [15:0] array_index_548042;
  wire [7:0] sel_548043;
  wire [7:0] add_548046;
  wire [7:0] sel_548047;
  wire [7:0] add_548050;
  wire [7:0] sel_548051;
  wire [7:0] add_548054;
  wire [7:0] sel_548055;
  wire [7:0] add_548058;
  wire [7:0] sel_548059;
  wire [7:0] add_548062;
  wire [7:0] sel_548063;
  wire [7:0] add_548066;
  wire [7:0] sel_548067;
  wire [7:0] add_548070;
  wire [7:0] sel_548071;
  wire [7:0] add_548074;
  wire [7:0] sel_548075;
  wire [7:0] add_548078;
  wire [7:0] sel_548079;
  wire [7:0] add_548082;
  wire [7:0] sel_548083;
  wire [7:0] add_548086;
  wire [7:0] sel_548087;
  wire [7:0] add_548090;
  wire [7:0] sel_548091;
  wire [7:0] add_548094;
  wire [7:0] sel_548095;
  wire [7:0] add_548098;
  wire [7:0] sel_548099;
  wire [7:0] add_548102;
  wire [7:0] sel_548103;
  wire [7:0] add_548106;
  wire [7:0] sel_548107;
  wire [7:0] add_548110;
  wire [7:0] sel_548111;
  wire [7:0] add_548114;
  wire [7:0] sel_548115;
  wire [7:0] add_548118;
  wire [7:0] sel_548119;
  wire [7:0] add_548122;
  wire [7:0] sel_548123;
  wire [7:0] add_548126;
  wire [7:0] sel_548127;
  wire [7:0] add_548130;
  wire [7:0] sel_548131;
  wire [7:0] add_548134;
  wire [7:0] sel_548135;
  wire [7:0] add_548138;
  wire [7:0] sel_548139;
  wire [7:0] add_548142;
  wire [7:0] sel_548143;
  wire [7:0] add_548146;
  wire [7:0] sel_548147;
  wire [7:0] add_548150;
  wire [7:0] sel_548151;
  wire [7:0] add_548154;
  wire [7:0] sel_548155;
  wire [7:0] add_548158;
  wire [7:0] sel_548159;
  wire [7:0] add_548162;
  wire [7:0] sel_548163;
  wire [7:0] add_548166;
  wire [7:0] sel_548167;
  wire [7:0] add_548170;
  wire [7:0] sel_548171;
  wire [7:0] add_548174;
  wire [7:0] sel_548175;
  wire [7:0] add_548178;
  wire [7:0] sel_548179;
  wire [7:0] add_548182;
  wire [7:0] sel_548183;
  wire [7:0] add_548186;
  wire [7:0] sel_548187;
  wire [7:0] add_548190;
  wire [7:0] sel_548191;
  wire [7:0] add_548194;
  wire [7:0] sel_548195;
  wire [7:0] add_548198;
  wire [7:0] sel_548199;
  wire [7:0] add_548202;
  wire [7:0] sel_548203;
  wire [7:0] add_548206;
  wire [7:0] sel_548207;
  wire [7:0] add_548210;
  wire [7:0] sel_548211;
  wire [7:0] add_548214;
  wire [7:0] sel_548215;
  wire [7:0] add_548218;
  wire [7:0] sel_548219;
  wire [7:0] add_548222;
  wire [7:0] sel_548223;
  wire [7:0] add_548226;
  wire [7:0] sel_548227;
  wire [7:0] add_548230;
  wire [7:0] sel_548231;
  wire [7:0] add_548234;
  wire [7:0] sel_548235;
  wire [7:0] add_548238;
  wire [7:0] sel_548239;
  wire [7:0] add_548242;
  wire [7:0] sel_548243;
  wire [7:0] add_548246;
  wire [7:0] sel_548247;
  wire [7:0] add_548250;
  wire [7:0] sel_548251;
  wire [7:0] add_548254;
  wire [7:0] sel_548255;
  wire [7:0] add_548258;
  wire [7:0] sel_548259;
  wire [7:0] add_548262;
  wire [7:0] sel_548263;
  wire [7:0] add_548266;
  wire [7:0] sel_548267;
  wire [7:0] add_548270;
  wire [7:0] sel_548271;
  wire [7:0] add_548274;
  wire [7:0] sel_548275;
  wire [7:0] add_548278;
  wire [7:0] sel_548279;
  wire [7:0] add_548282;
  wire [7:0] sel_548283;
  wire [7:0] add_548286;
  wire [7:0] sel_548287;
  wire [7:0] add_548290;
  wire [7:0] sel_548291;
  wire [7:0] add_548294;
  wire [7:0] sel_548295;
  wire [7:0] add_548298;
  wire [7:0] sel_548299;
  wire [7:0] add_548302;
  wire [7:0] sel_548303;
  wire [7:0] add_548306;
  wire [7:0] sel_548307;
  wire [7:0] add_548310;
  wire [7:0] sel_548311;
  wire [7:0] add_548314;
  wire [7:0] sel_548315;
  wire [7:0] add_548318;
  wire [7:0] sel_548319;
  wire [7:0] add_548322;
  wire [7:0] sel_548323;
  wire [7:0] add_548326;
  wire [7:0] sel_548327;
  wire [7:0] add_548330;
  wire [7:0] sel_548331;
  wire [7:0] add_548334;
  wire [7:0] sel_548335;
  wire [7:0] add_548338;
  wire [7:0] sel_548339;
  wire [7:0] add_548343;
  wire [15:0] array_index_548344;
  wire [7:0] sel_548345;
  wire [7:0] add_548348;
  wire [7:0] sel_548349;
  wire [7:0] add_548352;
  wire [7:0] sel_548353;
  wire [7:0] add_548356;
  wire [7:0] sel_548357;
  wire [7:0] add_548360;
  wire [7:0] sel_548361;
  wire [7:0] add_548364;
  wire [7:0] sel_548365;
  wire [7:0] add_548368;
  wire [7:0] sel_548369;
  wire [7:0] add_548372;
  wire [7:0] sel_548373;
  wire [7:0] add_548376;
  wire [7:0] sel_548377;
  wire [7:0] add_548380;
  wire [7:0] sel_548381;
  wire [7:0] add_548384;
  wire [7:0] sel_548385;
  wire [7:0] add_548388;
  wire [7:0] sel_548389;
  wire [7:0] add_548392;
  wire [7:0] sel_548393;
  wire [7:0] add_548396;
  wire [7:0] sel_548397;
  wire [7:0] add_548400;
  wire [7:0] sel_548401;
  wire [7:0] add_548404;
  wire [7:0] sel_548405;
  wire [7:0] add_548408;
  wire [7:0] sel_548409;
  wire [7:0] add_548412;
  wire [7:0] sel_548413;
  wire [7:0] add_548416;
  wire [7:0] sel_548417;
  wire [7:0] add_548420;
  wire [7:0] sel_548421;
  wire [7:0] add_548424;
  wire [7:0] sel_548425;
  wire [7:0] add_548428;
  wire [7:0] sel_548429;
  wire [7:0] add_548432;
  wire [7:0] sel_548433;
  wire [7:0] add_548436;
  wire [7:0] sel_548437;
  wire [7:0] add_548440;
  wire [7:0] sel_548441;
  wire [7:0] add_548444;
  wire [7:0] sel_548445;
  wire [7:0] add_548448;
  wire [7:0] sel_548449;
  wire [7:0] add_548452;
  wire [7:0] sel_548453;
  wire [7:0] add_548456;
  wire [7:0] sel_548457;
  wire [7:0] add_548460;
  wire [7:0] sel_548461;
  wire [7:0] add_548464;
  wire [7:0] sel_548465;
  wire [7:0] add_548468;
  wire [7:0] sel_548469;
  wire [7:0] add_548472;
  wire [7:0] sel_548473;
  wire [7:0] add_548476;
  wire [7:0] sel_548477;
  wire [7:0] add_548480;
  wire [7:0] sel_548481;
  wire [7:0] add_548484;
  wire [7:0] sel_548485;
  wire [7:0] add_548488;
  wire [7:0] sel_548489;
  wire [7:0] add_548492;
  wire [7:0] sel_548493;
  wire [7:0] add_548496;
  wire [7:0] sel_548497;
  wire [7:0] add_548500;
  wire [7:0] sel_548501;
  wire [7:0] add_548504;
  wire [7:0] sel_548505;
  wire [7:0] add_548508;
  wire [7:0] sel_548509;
  wire [7:0] add_548512;
  wire [7:0] sel_548513;
  wire [7:0] add_548516;
  wire [7:0] sel_548517;
  wire [7:0] add_548520;
  wire [7:0] sel_548521;
  wire [7:0] add_548524;
  wire [7:0] sel_548525;
  wire [7:0] add_548528;
  wire [7:0] sel_548529;
  wire [7:0] add_548532;
  wire [7:0] sel_548533;
  wire [7:0] add_548536;
  wire [7:0] sel_548537;
  wire [7:0] add_548540;
  wire [7:0] sel_548541;
  wire [7:0] add_548544;
  wire [7:0] sel_548545;
  wire [7:0] add_548548;
  wire [7:0] sel_548549;
  wire [7:0] add_548552;
  wire [7:0] sel_548553;
  wire [7:0] add_548556;
  wire [7:0] sel_548557;
  wire [7:0] add_548560;
  wire [7:0] sel_548561;
  wire [7:0] add_548564;
  wire [7:0] sel_548565;
  wire [7:0] add_548568;
  wire [7:0] sel_548569;
  wire [7:0] add_548572;
  wire [7:0] sel_548573;
  wire [7:0] add_548576;
  wire [7:0] sel_548577;
  wire [7:0] add_548580;
  wire [7:0] sel_548581;
  wire [7:0] add_548584;
  wire [7:0] sel_548585;
  wire [7:0] add_548588;
  wire [7:0] sel_548589;
  wire [7:0] add_548592;
  wire [7:0] sel_548593;
  wire [7:0] add_548596;
  wire [7:0] sel_548597;
  wire [7:0] add_548600;
  wire [7:0] sel_548601;
  wire [7:0] add_548604;
  wire [7:0] sel_548605;
  wire [7:0] add_548608;
  wire [7:0] sel_548609;
  wire [7:0] add_548612;
  wire [7:0] sel_548613;
  wire [7:0] add_548616;
  wire [7:0] sel_548617;
  wire [7:0] add_548620;
  wire [7:0] sel_548621;
  wire [7:0] add_548624;
  wire [7:0] sel_548625;
  wire [7:0] add_548628;
  wire [7:0] sel_548629;
  wire [7:0] add_548632;
  wire [7:0] sel_548633;
  wire [7:0] add_548636;
  wire [7:0] sel_548637;
  wire [7:0] add_548640;
  wire [7:0] sel_548641;
  wire [7:0] add_548645;
  wire [15:0] array_index_548646;
  wire [7:0] sel_548647;
  wire [7:0] add_548650;
  wire [7:0] sel_548651;
  wire [7:0] add_548654;
  wire [7:0] sel_548655;
  wire [7:0] add_548658;
  wire [7:0] sel_548659;
  wire [7:0] add_548662;
  wire [7:0] sel_548663;
  wire [7:0] add_548666;
  wire [7:0] sel_548667;
  wire [7:0] add_548670;
  wire [7:0] sel_548671;
  wire [7:0] add_548674;
  wire [7:0] sel_548675;
  wire [7:0] add_548678;
  wire [7:0] sel_548679;
  wire [7:0] add_548682;
  wire [7:0] sel_548683;
  wire [7:0] add_548686;
  wire [7:0] sel_548687;
  wire [7:0] add_548690;
  wire [7:0] sel_548691;
  wire [7:0] add_548694;
  wire [7:0] sel_548695;
  wire [7:0] add_548698;
  wire [7:0] sel_548699;
  wire [7:0] add_548702;
  wire [7:0] sel_548703;
  wire [7:0] add_548706;
  wire [7:0] sel_548707;
  wire [7:0] add_548710;
  wire [7:0] sel_548711;
  wire [7:0] add_548714;
  wire [7:0] sel_548715;
  wire [7:0] add_548718;
  wire [7:0] sel_548719;
  wire [7:0] add_548722;
  wire [7:0] sel_548723;
  wire [7:0] add_548726;
  wire [7:0] sel_548727;
  wire [7:0] add_548730;
  wire [7:0] sel_548731;
  wire [7:0] add_548734;
  wire [7:0] sel_548735;
  wire [7:0] add_548738;
  wire [7:0] sel_548739;
  wire [7:0] add_548742;
  wire [7:0] sel_548743;
  wire [7:0] add_548746;
  wire [7:0] sel_548747;
  wire [7:0] add_548750;
  wire [7:0] sel_548751;
  wire [7:0] add_548754;
  wire [7:0] sel_548755;
  wire [7:0] add_548758;
  wire [7:0] sel_548759;
  wire [7:0] add_548762;
  wire [7:0] sel_548763;
  wire [7:0] add_548766;
  wire [7:0] sel_548767;
  wire [7:0] add_548770;
  wire [7:0] sel_548771;
  wire [7:0] add_548774;
  wire [7:0] sel_548775;
  wire [7:0] add_548778;
  wire [7:0] sel_548779;
  wire [7:0] add_548782;
  wire [7:0] sel_548783;
  wire [7:0] add_548786;
  wire [7:0] sel_548787;
  wire [7:0] add_548790;
  wire [7:0] sel_548791;
  wire [7:0] add_548794;
  wire [7:0] sel_548795;
  wire [7:0] add_548798;
  wire [7:0] sel_548799;
  wire [7:0] add_548802;
  wire [7:0] sel_548803;
  wire [7:0] add_548806;
  wire [7:0] sel_548807;
  wire [7:0] add_548810;
  wire [7:0] sel_548811;
  wire [7:0] add_548814;
  wire [7:0] sel_548815;
  wire [7:0] add_548818;
  wire [7:0] sel_548819;
  wire [7:0] add_548822;
  wire [7:0] sel_548823;
  wire [7:0] add_548826;
  wire [7:0] sel_548827;
  wire [7:0] add_548830;
  wire [7:0] sel_548831;
  wire [7:0] add_548834;
  wire [7:0] sel_548835;
  wire [7:0] add_548838;
  wire [7:0] sel_548839;
  wire [7:0] add_548842;
  wire [7:0] sel_548843;
  wire [7:0] add_548846;
  wire [7:0] sel_548847;
  wire [7:0] add_548850;
  wire [7:0] sel_548851;
  wire [7:0] add_548854;
  wire [7:0] sel_548855;
  wire [7:0] add_548858;
  wire [7:0] sel_548859;
  wire [7:0] add_548862;
  wire [7:0] sel_548863;
  wire [7:0] add_548866;
  wire [7:0] sel_548867;
  wire [7:0] add_548870;
  wire [7:0] sel_548871;
  wire [7:0] add_548874;
  wire [7:0] sel_548875;
  wire [7:0] add_548878;
  wire [7:0] sel_548879;
  wire [7:0] add_548882;
  wire [7:0] sel_548883;
  wire [7:0] add_548886;
  wire [7:0] sel_548887;
  wire [7:0] add_548890;
  wire [7:0] sel_548891;
  wire [7:0] add_548894;
  wire [7:0] sel_548895;
  wire [7:0] add_548898;
  wire [7:0] sel_548899;
  wire [7:0] add_548902;
  wire [7:0] sel_548903;
  wire [7:0] add_548906;
  wire [7:0] sel_548907;
  wire [7:0] add_548910;
  wire [7:0] sel_548911;
  wire [7:0] add_548914;
  wire [7:0] sel_548915;
  wire [7:0] add_548918;
  wire [7:0] sel_548919;
  wire [7:0] add_548922;
  wire [7:0] sel_548923;
  wire [7:0] add_548926;
  wire [7:0] sel_548927;
  wire [7:0] add_548930;
  wire [7:0] sel_548931;
  wire [7:0] add_548934;
  wire [7:0] sel_548935;
  wire [7:0] add_548938;
  wire [7:0] sel_548939;
  wire [7:0] add_548942;
  wire [7:0] sel_548943;
  wire [7:0] add_548947;
  wire [15:0] array_index_548948;
  wire [7:0] sel_548949;
  wire [7:0] add_548952;
  wire [7:0] sel_548953;
  wire [7:0] add_548956;
  wire [7:0] sel_548957;
  wire [7:0] add_548960;
  wire [7:0] sel_548961;
  wire [7:0] add_548964;
  wire [7:0] sel_548965;
  wire [7:0] add_548968;
  wire [7:0] sel_548969;
  wire [7:0] add_548972;
  wire [7:0] sel_548973;
  wire [7:0] add_548976;
  wire [7:0] sel_548977;
  wire [7:0] add_548980;
  wire [7:0] sel_548981;
  wire [7:0] add_548984;
  wire [7:0] sel_548985;
  wire [7:0] add_548988;
  wire [7:0] sel_548989;
  wire [7:0] add_548992;
  wire [7:0] sel_548993;
  wire [7:0] add_548996;
  wire [7:0] sel_548997;
  wire [7:0] add_549000;
  wire [7:0] sel_549001;
  wire [7:0] add_549004;
  wire [7:0] sel_549005;
  wire [7:0] add_549008;
  wire [7:0] sel_549009;
  wire [7:0] add_549012;
  wire [7:0] sel_549013;
  wire [7:0] add_549016;
  wire [7:0] sel_549017;
  wire [7:0] add_549020;
  wire [7:0] sel_549021;
  wire [7:0] add_549024;
  wire [7:0] sel_549025;
  wire [7:0] add_549028;
  wire [7:0] sel_549029;
  wire [7:0] add_549032;
  wire [7:0] sel_549033;
  wire [7:0] add_549036;
  wire [7:0] sel_549037;
  wire [7:0] add_549040;
  wire [7:0] sel_549041;
  wire [7:0] add_549044;
  wire [7:0] sel_549045;
  wire [7:0] add_549048;
  wire [7:0] sel_549049;
  wire [7:0] add_549052;
  wire [7:0] sel_549053;
  wire [7:0] add_549056;
  wire [7:0] sel_549057;
  wire [7:0] add_549060;
  wire [7:0] sel_549061;
  wire [7:0] add_549064;
  wire [7:0] sel_549065;
  wire [7:0] add_549068;
  wire [7:0] sel_549069;
  wire [7:0] add_549072;
  wire [7:0] sel_549073;
  wire [7:0] add_549076;
  wire [7:0] sel_549077;
  wire [7:0] add_549080;
  wire [7:0] sel_549081;
  wire [7:0] add_549084;
  wire [7:0] sel_549085;
  wire [7:0] add_549088;
  wire [7:0] sel_549089;
  wire [7:0] add_549092;
  wire [7:0] sel_549093;
  wire [7:0] add_549096;
  wire [7:0] sel_549097;
  wire [7:0] add_549100;
  wire [7:0] sel_549101;
  wire [7:0] add_549104;
  wire [7:0] sel_549105;
  wire [7:0] add_549108;
  wire [7:0] sel_549109;
  wire [7:0] add_549112;
  wire [7:0] sel_549113;
  wire [7:0] add_549116;
  wire [7:0] sel_549117;
  wire [7:0] add_549120;
  wire [7:0] sel_549121;
  wire [7:0] add_549124;
  wire [7:0] sel_549125;
  wire [7:0] add_549128;
  wire [7:0] sel_549129;
  wire [7:0] add_549132;
  wire [7:0] sel_549133;
  wire [7:0] add_549136;
  wire [7:0] sel_549137;
  wire [7:0] add_549140;
  wire [7:0] sel_549141;
  wire [7:0] add_549144;
  wire [7:0] sel_549145;
  wire [7:0] add_549148;
  wire [7:0] sel_549149;
  wire [7:0] add_549152;
  wire [7:0] sel_549153;
  wire [7:0] add_549156;
  wire [7:0] sel_549157;
  wire [7:0] add_549160;
  wire [7:0] sel_549161;
  wire [7:0] add_549164;
  wire [7:0] sel_549165;
  wire [7:0] add_549168;
  wire [7:0] sel_549169;
  wire [7:0] add_549172;
  wire [7:0] sel_549173;
  wire [7:0] add_549176;
  wire [7:0] sel_549177;
  wire [7:0] add_549180;
  wire [7:0] sel_549181;
  wire [7:0] add_549184;
  wire [7:0] sel_549185;
  wire [7:0] add_549188;
  wire [7:0] sel_549189;
  wire [7:0] add_549192;
  wire [7:0] sel_549193;
  wire [7:0] add_549196;
  wire [7:0] sel_549197;
  wire [7:0] add_549200;
  wire [7:0] sel_549201;
  wire [7:0] add_549204;
  wire [7:0] sel_549205;
  wire [7:0] add_549208;
  wire [7:0] sel_549209;
  wire [7:0] add_549212;
  wire [7:0] sel_549213;
  wire [7:0] add_549216;
  wire [7:0] sel_549217;
  wire [7:0] add_549220;
  wire [7:0] sel_549221;
  wire [7:0] add_549224;
  wire [7:0] sel_549225;
  wire [7:0] add_549228;
  wire [7:0] sel_549229;
  wire [7:0] add_549232;
  wire [7:0] sel_549233;
  wire [7:0] add_549236;
  wire [7:0] sel_549237;
  wire [7:0] add_549240;
  wire [7:0] sel_549241;
  wire [7:0] add_549244;
  wire [7:0] sel_549245;
  wire [7:0] add_549249;
  wire [15:0] array_index_549250;
  wire [7:0] sel_549251;
  wire [7:0] add_549254;
  wire [7:0] sel_549255;
  wire [7:0] add_549258;
  wire [7:0] sel_549259;
  wire [7:0] add_549262;
  wire [7:0] sel_549263;
  wire [7:0] add_549266;
  wire [7:0] sel_549267;
  wire [7:0] add_549270;
  wire [7:0] sel_549271;
  wire [7:0] add_549274;
  wire [7:0] sel_549275;
  wire [7:0] add_549278;
  wire [7:0] sel_549279;
  wire [7:0] add_549282;
  wire [7:0] sel_549283;
  wire [7:0] add_549286;
  wire [7:0] sel_549287;
  wire [7:0] add_549290;
  wire [7:0] sel_549291;
  wire [7:0] add_549294;
  wire [7:0] sel_549295;
  wire [7:0] add_549298;
  wire [7:0] sel_549299;
  wire [7:0] add_549302;
  wire [7:0] sel_549303;
  wire [7:0] add_549306;
  wire [7:0] sel_549307;
  wire [7:0] add_549310;
  wire [7:0] sel_549311;
  wire [7:0] add_549314;
  wire [7:0] sel_549315;
  wire [7:0] add_549318;
  wire [7:0] sel_549319;
  wire [7:0] add_549322;
  wire [7:0] sel_549323;
  wire [7:0] add_549326;
  wire [7:0] sel_549327;
  wire [7:0] add_549330;
  wire [7:0] sel_549331;
  wire [7:0] add_549334;
  wire [7:0] sel_549335;
  wire [7:0] add_549338;
  wire [7:0] sel_549339;
  wire [7:0] add_549342;
  wire [7:0] sel_549343;
  wire [7:0] add_549346;
  wire [7:0] sel_549347;
  wire [7:0] add_549350;
  wire [7:0] sel_549351;
  wire [7:0] add_549354;
  wire [7:0] sel_549355;
  wire [7:0] add_549358;
  wire [7:0] sel_549359;
  wire [7:0] add_549362;
  wire [7:0] sel_549363;
  wire [7:0] add_549366;
  wire [7:0] sel_549367;
  wire [7:0] add_549370;
  wire [7:0] sel_549371;
  wire [7:0] add_549374;
  wire [7:0] sel_549375;
  wire [7:0] add_549378;
  wire [7:0] sel_549379;
  wire [7:0] add_549382;
  wire [7:0] sel_549383;
  wire [7:0] add_549386;
  wire [7:0] sel_549387;
  wire [7:0] add_549390;
  wire [7:0] sel_549391;
  wire [7:0] add_549394;
  wire [7:0] sel_549395;
  wire [7:0] add_549398;
  wire [7:0] sel_549399;
  wire [7:0] add_549402;
  wire [7:0] sel_549403;
  wire [7:0] add_549406;
  wire [7:0] sel_549407;
  wire [7:0] add_549410;
  wire [7:0] sel_549411;
  wire [7:0] add_549414;
  wire [7:0] sel_549415;
  wire [7:0] add_549418;
  wire [7:0] sel_549419;
  wire [7:0] add_549422;
  wire [7:0] sel_549423;
  wire [7:0] add_549426;
  wire [7:0] sel_549427;
  wire [7:0] add_549430;
  wire [7:0] sel_549431;
  wire [7:0] add_549434;
  wire [7:0] sel_549435;
  wire [7:0] add_549438;
  wire [7:0] sel_549439;
  wire [7:0] add_549442;
  wire [7:0] sel_549443;
  wire [7:0] add_549446;
  wire [7:0] sel_549447;
  wire [7:0] add_549450;
  wire [7:0] sel_549451;
  wire [7:0] add_549454;
  wire [7:0] sel_549455;
  wire [7:0] add_549458;
  wire [7:0] sel_549459;
  wire [7:0] add_549462;
  wire [7:0] sel_549463;
  wire [7:0] add_549466;
  wire [7:0] sel_549467;
  wire [7:0] add_549470;
  wire [7:0] sel_549471;
  wire [7:0] add_549474;
  wire [7:0] sel_549475;
  wire [7:0] add_549478;
  wire [7:0] sel_549479;
  wire [7:0] add_549482;
  wire [7:0] sel_549483;
  wire [7:0] add_549486;
  wire [7:0] sel_549487;
  wire [7:0] add_549490;
  wire [7:0] sel_549491;
  wire [7:0] add_549494;
  wire [7:0] sel_549495;
  wire [7:0] add_549498;
  wire [7:0] sel_549499;
  wire [7:0] add_549502;
  wire [7:0] sel_549503;
  wire [7:0] add_549506;
  wire [7:0] sel_549507;
  wire [7:0] add_549510;
  wire [7:0] sel_549511;
  wire [7:0] add_549514;
  wire [7:0] sel_549515;
  wire [7:0] add_549518;
  wire [7:0] sel_549519;
  wire [7:0] add_549522;
  wire [7:0] sel_549523;
  wire [7:0] add_549526;
  wire [7:0] sel_549527;
  wire [7:0] add_549530;
  wire [7:0] sel_549531;
  wire [7:0] add_549534;
  wire [7:0] sel_549535;
  wire [7:0] add_549538;
  wire [7:0] sel_549539;
  wire [7:0] add_549542;
  wire [7:0] sel_549543;
  wire [7:0] add_549546;
  wire [7:0] sel_549547;
  wire [7:0] add_549551;
  wire [15:0] array_index_549552;
  wire [7:0] sel_549553;
  wire [7:0] add_549556;
  wire [7:0] sel_549557;
  wire [7:0] add_549560;
  wire [7:0] sel_549561;
  wire [7:0] add_549564;
  wire [7:0] sel_549565;
  wire [7:0] add_549568;
  wire [7:0] sel_549569;
  wire [7:0] add_549572;
  wire [7:0] sel_549573;
  wire [7:0] add_549576;
  wire [7:0] sel_549577;
  wire [7:0] add_549580;
  wire [7:0] sel_549581;
  wire [7:0] add_549584;
  wire [7:0] sel_549585;
  wire [7:0] add_549588;
  wire [7:0] sel_549589;
  wire [7:0] add_549592;
  wire [7:0] sel_549593;
  wire [7:0] add_549596;
  wire [7:0] sel_549597;
  wire [7:0] add_549600;
  wire [7:0] sel_549601;
  wire [7:0] add_549604;
  wire [7:0] sel_549605;
  wire [7:0] add_549608;
  wire [7:0] sel_549609;
  wire [7:0] add_549612;
  wire [7:0] sel_549613;
  wire [7:0] add_549616;
  wire [7:0] sel_549617;
  wire [7:0] add_549620;
  wire [7:0] sel_549621;
  wire [7:0] add_549624;
  wire [7:0] sel_549625;
  wire [7:0] add_549628;
  wire [7:0] sel_549629;
  wire [7:0] add_549632;
  wire [7:0] sel_549633;
  wire [7:0] add_549636;
  wire [7:0] sel_549637;
  wire [7:0] add_549640;
  wire [7:0] sel_549641;
  wire [7:0] add_549644;
  wire [7:0] sel_549645;
  wire [7:0] add_549648;
  wire [7:0] sel_549649;
  wire [7:0] add_549652;
  wire [7:0] sel_549653;
  wire [7:0] add_549656;
  wire [7:0] sel_549657;
  wire [7:0] add_549660;
  wire [7:0] sel_549661;
  wire [7:0] add_549664;
  wire [7:0] sel_549665;
  wire [7:0] add_549668;
  wire [7:0] sel_549669;
  wire [7:0] add_549672;
  wire [7:0] sel_549673;
  wire [7:0] add_549676;
  wire [7:0] sel_549677;
  wire [7:0] add_549680;
  wire [7:0] sel_549681;
  wire [7:0] add_549684;
  wire [7:0] sel_549685;
  wire [7:0] add_549688;
  wire [7:0] sel_549689;
  wire [7:0] add_549692;
  wire [7:0] sel_549693;
  wire [7:0] add_549696;
  wire [7:0] sel_549697;
  wire [7:0] add_549700;
  wire [7:0] sel_549701;
  wire [7:0] add_549704;
  wire [7:0] sel_549705;
  wire [7:0] add_549708;
  wire [7:0] sel_549709;
  wire [7:0] add_549712;
  wire [7:0] sel_549713;
  wire [7:0] add_549716;
  wire [7:0] sel_549717;
  wire [7:0] add_549720;
  wire [7:0] sel_549721;
  wire [7:0] add_549724;
  wire [7:0] sel_549725;
  wire [7:0] add_549728;
  wire [7:0] sel_549729;
  wire [7:0] add_549732;
  wire [7:0] sel_549733;
  wire [7:0] add_549736;
  wire [7:0] sel_549737;
  wire [7:0] add_549740;
  wire [7:0] sel_549741;
  wire [7:0] add_549744;
  wire [7:0] sel_549745;
  wire [7:0] add_549748;
  wire [7:0] sel_549749;
  wire [7:0] add_549752;
  wire [7:0] sel_549753;
  wire [7:0] add_549756;
  wire [7:0] sel_549757;
  wire [7:0] add_549760;
  wire [7:0] sel_549761;
  wire [7:0] add_549764;
  wire [7:0] sel_549765;
  wire [7:0] add_549768;
  wire [7:0] sel_549769;
  wire [7:0] add_549772;
  wire [7:0] sel_549773;
  wire [7:0] add_549776;
  wire [7:0] sel_549777;
  wire [7:0] add_549780;
  wire [7:0] sel_549781;
  wire [7:0] add_549784;
  wire [7:0] sel_549785;
  wire [7:0] add_549788;
  wire [7:0] sel_549789;
  wire [7:0] add_549792;
  wire [7:0] sel_549793;
  wire [7:0] add_549796;
  wire [7:0] sel_549797;
  wire [7:0] add_549800;
  wire [7:0] sel_549801;
  wire [7:0] add_549804;
  wire [7:0] sel_549805;
  wire [7:0] add_549808;
  wire [7:0] sel_549809;
  wire [7:0] add_549812;
  wire [7:0] sel_549813;
  wire [7:0] add_549816;
  wire [7:0] sel_549817;
  wire [7:0] add_549820;
  wire [7:0] sel_549821;
  wire [7:0] add_549824;
  wire [7:0] sel_549825;
  wire [7:0] add_549828;
  wire [7:0] sel_549829;
  wire [7:0] add_549832;
  wire [7:0] sel_549833;
  wire [7:0] add_549836;
  wire [7:0] sel_549837;
  wire [7:0] add_549840;
  wire [7:0] sel_549841;
  wire [7:0] add_549844;
  wire [7:0] sel_549845;
  wire [7:0] add_549848;
  wire [7:0] sel_549849;
  wire [7:0] add_549853;
  wire [15:0] array_index_549854;
  wire [7:0] sel_549855;
  wire [7:0] add_549858;
  wire [7:0] sel_549859;
  wire [7:0] add_549862;
  wire [7:0] sel_549863;
  wire [7:0] add_549866;
  wire [7:0] sel_549867;
  wire [7:0] add_549870;
  wire [7:0] sel_549871;
  wire [7:0] add_549874;
  wire [7:0] sel_549875;
  wire [7:0] add_549878;
  wire [7:0] sel_549879;
  wire [7:0] add_549882;
  wire [7:0] sel_549883;
  wire [7:0] add_549886;
  wire [7:0] sel_549887;
  wire [7:0] add_549890;
  wire [7:0] sel_549891;
  wire [7:0] add_549894;
  wire [7:0] sel_549895;
  wire [7:0] add_549898;
  wire [7:0] sel_549899;
  wire [7:0] add_549902;
  wire [7:0] sel_549903;
  wire [7:0] add_549906;
  wire [7:0] sel_549907;
  wire [7:0] add_549910;
  wire [7:0] sel_549911;
  wire [7:0] add_549914;
  wire [7:0] sel_549915;
  wire [7:0] add_549918;
  wire [7:0] sel_549919;
  wire [7:0] add_549922;
  wire [7:0] sel_549923;
  wire [7:0] add_549926;
  wire [7:0] sel_549927;
  wire [7:0] add_549930;
  wire [7:0] sel_549931;
  wire [7:0] add_549934;
  wire [7:0] sel_549935;
  wire [7:0] add_549938;
  wire [7:0] sel_549939;
  wire [7:0] add_549942;
  wire [7:0] sel_549943;
  wire [7:0] add_549946;
  wire [7:0] sel_549947;
  wire [7:0] add_549950;
  wire [7:0] sel_549951;
  wire [7:0] add_549954;
  wire [7:0] sel_549955;
  wire [7:0] add_549958;
  wire [7:0] sel_549959;
  wire [7:0] add_549962;
  wire [7:0] sel_549963;
  wire [7:0] add_549966;
  wire [7:0] sel_549967;
  wire [7:0] add_549970;
  wire [7:0] sel_549971;
  wire [7:0] add_549974;
  wire [7:0] sel_549975;
  wire [7:0] add_549978;
  wire [7:0] sel_549979;
  wire [7:0] add_549982;
  wire [7:0] sel_549983;
  wire [7:0] add_549986;
  wire [7:0] sel_549987;
  wire [7:0] add_549990;
  wire [7:0] sel_549991;
  wire [7:0] add_549994;
  wire [7:0] sel_549995;
  wire [7:0] add_549998;
  wire [7:0] sel_549999;
  wire [7:0] add_550002;
  wire [7:0] sel_550003;
  wire [7:0] add_550006;
  wire [7:0] sel_550007;
  wire [7:0] add_550010;
  wire [7:0] sel_550011;
  wire [7:0] add_550014;
  wire [7:0] sel_550015;
  wire [7:0] add_550018;
  wire [7:0] sel_550019;
  wire [7:0] add_550022;
  wire [7:0] sel_550023;
  wire [7:0] add_550026;
  wire [7:0] sel_550027;
  wire [7:0] add_550030;
  wire [7:0] sel_550031;
  wire [7:0] add_550034;
  wire [7:0] sel_550035;
  wire [7:0] add_550038;
  wire [7:0] sel_550039;
  wire [7:0] add_550042;
  wire [7:0] sel_550043;
  wire [7:0] add_550046;
  wire [7:0] sel_550047;
  wire [7:0] add_550050;
  wire [7:0] sel_550051;
  wire [7:0] add_550054;
  wire [7:0] sel_550055;
  wire [7:0] add_550058;
  wire [7:0] sel_550059;
  wire [7:0] add_550062;
  wire [7:0] sel_550063;
  wire [7:0] add_550066;
  wire [7:0] sel_550067;
  wire [7:0] add_550070;
  wire [7:0] sel_550071;
  wire [7:0] add_550074;
  wire [7:0] sel_550075;
  wire [7:0] add_550078;
  wire [7:0] sel_550079;
  wire [7:0] add_550082;
  wire [7:0] sel_550083;
  wire [7:0] add_550086;
  wire [7:0] sel_550087;
  wire [7:0] add_550090;
  wire [7:0] sel_550091;
  wire [7:0] add_550094;
  wire [7:0] sel_550095;
  wire [7:0] add_550098;
  wire [7:0] sel_550099;
  wire [7:0] add_550102;
  wire [7:0] sel_550103;
  wire [7:0] add_550106;
  wire [7:0] sel_550107;
  wire [7:0] add_550110;
  wire [7:0] sel_550111;
  wire [7:0] add_550114;
  wire [7:0] sel_550115;
  wire [7:0] add_550118;
  wire [7:0] sel_550119;
  wire [7:0] add_550122;
  wire [7:0] sel_550123;
  wire [7:0] add_550126;
  wire [7:0] sel_550127;
  wire [7:0] add_550130;
  wire [7:0] sel_550131;
  wire [7:0] add_550134;
  wire [7:0] sel_550135;
  wire [7:0] add_550138;
  wire [7:0] sel_550139;
  wire [7:0] add_550142;
  wire [7:0] sel_550143;
  wire [7:0] add_550146;
  wire [7:0] sel_550147;
  wire [7:0] add_550150;
  wire [7:0] sel_550151;
  wire [7:0] add_550155;
  wire [15:0] array_index_550156;
  wire [7:0] sel_550157;
  wire [7:0] add_550160;
  wire [7:0] sel_550161;
  wire [7:0] add_550164;
  wire [7:0] sel_550165;
  wire [7:0] add_550168;
  wire [7:0] sel_550169;
  wire [7:0] add_550172;
  wire [7:0] sel_550173;
  wire [7:0] add_550176;
  wire [7:0] sel_550177;
  wire [7:0] add_550180;
  wire [7:0] sel_550181;
  wire [7:0] add_550184;
  wire [7:0] sel_550185;
  wire [7:0] add_550188;
  wire [7:0] sel_550189;
  wire [7:0] add_550192;
  wire [7:0] sel_550193;
  wire [7:0] add_550196;
  wire [7:0] sel_550197;
  wire [7:0] add_550200;
  wire [7:0] sel_550201;
  wire [7:0] add_550204;
  wire [7:0] sel_550205;
  wire [7:0] add_550208;
  wire [7:0] sel_550209;
  wire [7:0] add_550212;
  wire [7:0] sel_550213;
  wire [7:0] add_550216;
  wire [7:0] sel_550217;
  wire [7:0] add_550220;
  wire [7:0] sel_550221;
  wire [7:0] add_550224;
  wire [7:0] sel_550225;
  wire [7:0] add_550228;
  wire [7:0] sel_550229;
  wire [7:0] add_550232;
  wire [7:0] sel_550233;
  wire [7:0] add_550236;
  wire [7:0] sel_550237;
  wire [7:0] add_550240;
  wire [7:0] sel_550241;
  wire [7:0] add_550244;
  wire [7:0] sel_550245;
  wire [7:0] add_550248;
  wire [7:0] sel_550249;
  wire [7:0] add_550252;
  wire [7:0] sel_550253;
  wire [7:0] add_550256;
  wire [7:0] sel_550257;
  wire [7:0] add_550260;
  wire [7:0] sel_550261;
  wire [7:0] add_550264;
  wire [7:0] sel_550265;
  wire [7:0] add_550268;
  wire [7:0] sel_550269;
  wire [7:0] add_550272;
  wire [7:0] sel_550273;
  wire [7:0] add_550276;
  wire [7:0] sel_550277;
  wire [7:0] add_550280;
  wire [7:0] sel_550281;
  wire [7:0] add_550284;
  wire [7:0] sel_550285;
  wire [7:0] add_550288;
  wire [7:0] sel_550289;
  wire [7:0] add_550292;
  wire [7:0] sel_550293;
  wire [7:0] add_550296;
  wire [7:0] sel_550297;
  wire [7:0] add_550300;
  wire [7:0] sel_550301;
  wire [7:0] add_550304;
  wire [7:0] sel_550305;
  wire [7:0] add_550308;
  wire [7:0] sel_550309;
  wire [7:0] add_550312;
  wire [7:0] sel_550313;
  wire [7:0] add_550316;
  wire [7:0] sel_550317;
  wire [7:0] add_550320;
  wire [7:0] sel_550321;
  wire [7:0] add_550324;
  wire [7:0] sel_550325;
  wire [7:0] add_550328;
  wire [7:0] sel_550329;
  wire [7:0] add_550332;
  wire [7:0] sel_550333;
  wire [7:0] add_550336;
  wire [7:0] sel_550337;
  wire [7:0] add_550340;
  wire [7:0] sel_550341;
  wire [7:0] add_550344;
  wire [7:0] sel_550345;
  wire [7:0] add_550348;
  wire [7:0] sel_550349;
  wire [7:0] add_550352;
  wire [7:0] sel_550353;
  wire [7:0] add_550356;
  wire [7:0] sel_550357;
  wire [7:0] add_550360;
  wire [7:0] sel_550361;
  wire [7:0] add_550364;
  wire [7:0] sel_550365;
  wire [7:0] add_550368;
  wire [7:0] sel_550369;
  wire [7:0] add_550372;
  wire [7:0] sel_550373;
  wire [7:0] add_550376;
  wire [7:0] sel_550377;
  wire [7:0] add_550380;
  wire [7:0] sel_550381;
  wire [7:0] add_550384;
  wire [7:0] sel_550385;
  wire [7:0] add_550388;
  wire [7:0] sel_550389;
  wire [7:0] add_550392;
  wire [7:0] sel_550393;
  wire [7:0] add_550396;
  wire [7:0] sel_550397;
  wire [7:0] add_550400;
  wire [7:0] sel_550401;
  wire [7:0] add_550404;
  wire [7:0] sel_550405;
  wire [7:0] add_550408;
  wire [7:0] sel_550409;
  wire [7:0] add_550412;
  wire [7:0] sel_550413;
  wire [7:0] add_550416;
  wire [7:0] sel_550417;
  wire [7:0] add_550420;
  wire [7:0] sel_550421;
  wire [7:0] add_550424;
  wire [7:0] sel_550425;
  wire [7:0] add_550428;
  wire [7:0] sel_550429;
  wire [7:0] add_550432;
  wire [7:0] sel_550433;
  wire [7:0] add_550436;
  wire [7:0] sel_550437;
  wire [7:0] add_550440;
  wire [7:0] sel_550441;
  wire [7:0] add_550444;
  wire [7:0] sel_550445;
  wire [7:0] add_550448;
  wire [7:0] sel_550449;
  wire [7:0] add_550452;
  wire [7:0] sel_550453;
  wire [7:0] add_550457;
  wire [15:0] array_index_550458;
  wire [7:0] sel_550459;
  wire [7:0] add_550462;
  wire [7:0] sel_550463;
  wire [7:0] add_550466;
  wire [7:0] sel_550467;
  wire [7:0] add_550470;
  wire [7:0] sel_550471;
  wire [7:0] add_550474;
  wire [7:0] sel_550475;
  wire [7:0] add_550478;
  wire [7:0] sel_550479;
  wire [7:0] add_550482;
  wire [7:0] sel_550483;
  wire [7:0] add_550486;
  wire [7:0] sel_550487;
  wire [7:0] add_550490;
  wire [7:0] sel_550491;
  wire [7:0] add_550494;
  wire [7:0] sel_550495;
  wire [7:0] add_550498;
  wire [7:0] sel_550499;
  wire [7:0] add_550502;
  wire [7:0] sel_550503;
  wire [7:0] add_550506;
  wire [7:0] sel_550507;
  wire [7:0] add_550510;
  wire [7:0] sel_550511;
  wire [7:0] add_550514;
  wire [7:0] sel_550515;
  wire [7:0] add_550518;
  wire [7:0] sel_550519;
  wire [7:0] add_550522;
  wire [7:0] sel_550523;
  wire [7:0] add_550526;
  wire [7:0] sel_550527;
  wire [7:0] add_550530;
  wire [7:0] sel_550531;
  wire [7:0] add_550534;
  wire [7:0] sel_550535;
  wire [7:0] add_550538;
  wire [7:0] sel_550539;
  wire [7:0] add_550542;
  wire [7:0] sel_550543;
  wire [7:0] add_550546;
  wire [7:0] sel_550547;
  wire [7:0] add_550550;
  wire [7:0] sel_550551;
  wire [7:0] add_550554;
  wire [7:0] sel_550555;
  wire [7:0] add_550558;
  wire [7:0] sel_550559;
  wire [7:0] add_550562;
  wire [7:0] sel_550563;
  wire [7:0] add_550566;
  wire [7:0] sel_550567;
  wire [7:0] add_550570;
  wire [7:0] sel_550571;
  wire [7:0] add_550574;
  wire [7:0] sel_550575;
  wire [7:0] add_550578;
  wire [7:0] sel_550579;
  wire [7:0] add_550582;
  wire [7:0] sel_550583;
  wire [7:0] add_550586;
  wire [7:0] sel_550587;
  wire [7:0] add_550590;
  wire [7:0] sel_550591;
  wire [7:0] add_550594;
  wire [7:0] sel_550595;
  wire [7:0] add_550598;
  wire [7:0] sel_550599;
  wire [7:0] add_550602;
  wire [7:0] sel_550603;
  wire [7:0] add_550606;
  wire [7:0] sel_550607;
  wire [7:0] add_550610;
  wire [7:0] sel_550611;
  wire [7:0] add_550614;
  wire [7:0] sel_550615;
  wire [7:0] add_550618;
  wire [7:0] sel_550619;
  wire [7:0] add_550622;
  wire [7:0] sel_550623;
  wire [7:0] add_550626;
  wire [7:0] sel_550627;
  wire [7:0] add_550630;
  wire [7:0] sel_550631;
  wire [7:0] add_550634;
  wire [7:0] sel_550635;
  wire [7:0] add_550638;
  wire [7:0] sel_550639;
  wire [7:0] add_550642;
  wire [7:0] sel_550643;
  wire [7:0] add_550646;
  wire [7:0] sel_550647;
  wire [7:0] add_550650;
  wire [7:0] sel_550651;
  wire [7:0] add_550654;
  wire [7:0] sel_550655;
  wire [7:0] add_550658;
  wire [7:0] sel_550659;
  wire [7:0] add_550662;
  wire [7:0] sel_550663;
  wire [7:0] add_550666;
  wire [7:0] sel_550667;
  wire [7:0] add_550670;
  wire [7:0] sel_550671;
  wire [7:0] add_550674;
  wire [7:0] sel_550675;
  wire [7:0] add_550678;
  wire [7:0] sel_550679;
  wire [7:0] add_550682;
  wire [7:0] sel_550683;
  wire [7:0] add_550686;
  wire [7:0] sel_550687;
  wire [7:0] add_550690;
  wire [7:0] sel_550691;
  wire [7:0] add_550694;
  wire [7:0] sel_550695;
  wire [7:0] add_550698;
  wire [7:0] sel_550699;
  wire [7:0] add_550702;
  wire [7:0] sel_550703;
  wire [7:0] add_550706;
  wire [7:0] sel_550707;
  wire [7:0] add_550710;
  wire [7:0] sel_550711;
  wire [7:0] add_550714;
  wire [7:0] sel_550715;
  wire [7:0] add_550718;
  wire [7:0] sel_550719;
  wire [7:0] add_550722;
  wire [7:0] sel_550723;
  wire [7:0] add_550726;
  wire [7:0] sel_550727;
  wire [7:0] add_550730;
  wire [7:0] sel_550731;
  wire [7:0] add_550734;
  wire [7:0] sel_550735;
  wire [7:0] add_550738;
  wire [7:0] sel_550739;
  wire [7:0] add_550742;
  wire [7:0] sel_550743;
  wire [7:0] add_550746;
  wire [7:0] sel_550747;
  wire [7:0] add_550750;
  wire [7:0] sel_550751;
  wire [7:0] add_550754;
  wire [7:0] sel_550755;
  wire [7:0] add_550759;
  wire [15:0] array_index_550760;
  wire [7:0] sel_550761;
  wire [7:0] add_550764;
  wire [7:0] sel_550765;
  wire [7:0] add_550768;
  wire [7:0] sel_550769;
  wire [7:0] add_550772;
  wire [7:0] sel_550773;
  wire [7:0] add_550776;
  wire [7:0] sel_550777;
  wire [7:0] add_550780;
  wire [7:0] sel_550781;
  wire [7:0] add_550784;
  wire [7:0] sel_550785;
  wire [7:0] add_550788;
  wire [7:0] sel_550789;
  wire [7:0] add_550792;
  wire [7:0] sel_550793;
  wire [7:0] add_550796;
  wire [7:0] sel_550797;
  wire [7:0] add_550800;
  wire [7:0] sel_550801;
  wire [7:0] add_550804;
  wire [7:0] sel_550805;
  wire [7:0] add_550808;
  wire [7:0] sel_550809;
  wire [7:0] add_550812;
  wire [7:0] sel_550813;
  wire [7:0] add_550816;
  wire [7:0] sel_550817;
  wire [7:0] add_550820;
  wire [7:0] sel_550821;
  wire [7:0] add_550824;
  wire [7:0] sel_550825;
  wire [7:0] add_550828;
  wire [7:0] sel_550829;
  wire [7:0] add_550832;
  wire [7:0] sel_550833;
  wire [7:0] add_550836;
  wire [7:0] sel_550837;
  wire [7:0] add_550840;
  wire [7:0] sel_550841;
  wire [7:0] add_550844;
  wire [7:0] sel_550845;
  wire [7:0] add_550848;
  wire [7:0] sel_550849;
  wire [7:0] add_550852;
  wire [7:0] sel_550853;
  wire [7:0] add_550856;
  wire [7:0] sel_550857;
  wire [7:0] add_550860;
  wire [7:0] sel_550861;
  wire [7:0] add_550864;
  wire [7:0] sel_550865;
  wire [7:0] add_550868;
  wire [7:0] sel_550869;
  wire [7:0] add_550872;
  wire [7:0] sel_550873;
  wire [7:0] add_550876;
  wire [7:0] sel_550877;
  wire [7:0] add_550880;
  wire [7:0] sel_550881;
  wire [7:0] add_550884;
  wire [7:0] sel_550885;
  wire [7:0] add_550888;
  wire [7:0] sel_550889;
  wire [7:0] add_550892;
  wire [7:0] sel_550893;
  wire [7:0] add_550896;
  wire [7:0] sel_550897;
  wire [7:0] add_550900;
  wire [7:0] sel_550901;
  wire [7:0] add_550904;
  wire [7:0] sel_550905;
  wire [7:0] add_550908;
  wire [7:0] sel_550909;
  wire [7:0] add_550912;
  wire [7:0] sel_550913;
  wire [7:0] add_550916;
  wire [7:0] sel_550917;
  wire [7:0] add_550920;
  wire [7:0] sel_550921;
  wire [7:0] add_550924;
  wire [7:0] sel_550925;
  wire [7:0] add_550928;
  wire [7:0] sel_550929;
  wire [7:0] add_550932;
  wire [7:0] sel_550933;
  wire [7:0] add_550936;
  wire [7:0] sel_550937;
  wire [7:0] add_550940;
  wire [7:0] sel_550941;
  wire [7:0] add_550944;
  wire [7:0] sel_550945;
  wire [7:0] add_550948;
  wire [7:0] sel_550949;
  wire [7:0] add_550952;
  wire [7:0] sel_550953;
  wire [7:0] add_550956;
  wire [7:0] sel_550957;
  wire [7:0] add_550960;
  wire [7:0] sel_550961;
  wire [7:0] add_550964;
  wire [7:0] sel_550965;
  wire [7:0] add_550968;
  wire [7:0] sel_550969;
  wire [7:0] add_550972;
  wire [7:0] sel_550973;
  wire [7:0] add_550976;
  wire [7:0] sel_550977;
  wire [7:0] add_550980;
  wire [7:0] sel_550981;
  wire [7:0] add_550984;
  wire [7:0] sel_550985;
  wire [7:0] add_550988;
  wire [7:0] sel_550989;
  wire [7:0] add_550992;
  wire [7:0] sel_550993;
  wire [7:0] add_550996;
  wire [7:0] sel_550997;
  wire [7:0] add_551000;
  wire [7:0] sel_551001;
  wire [7:0] add_551004;
  wire [7:0] sel_551005;
  wire [7:0] add_551008;
  wire [7:0] sel_551009;
  wire [7:0] add_551012;
  wire [7:0] sel_551013;
  wire [7:0] add_551016;
  wire [7:0] sel_551017;
  wire [7:0] add_551020;
  wire [7:0] sel_551021;
  wire [7:0] add_551024;
  wire [7:0] sel_551025;
  wire [7:0] add_551028;
  wire [7:0] sel_551029;
  wire [7:0] add_551032;
  wire [7:0] sel_551033;
  wire [7:0] add_551036;
  wire [7:0] sel_551037;
  wire [7:0] add_551040;
  wire [7:0] sel_551041;
  wire [7:0] add_551044;
  wire [7:0] sel_551045;
  wire [7:0] add_551048;
  wire [7:0] sel_551049;
  wire [7:0] add_551052;
  wire [7:0] sel_551053;
  wire [7:0] add_551056;
  wire [7:0] sel_551057;
  wire [7:0] add_551061;
  wire [15:0] array_index_551062;
  wire [7:0] sel_551063;
  wire [7:0] add_551066;
  wire [7:0] sel_551067;
  wire [7:0] add_551070;
  wire [7:0] sel_551071;
  wire [7:0] add_551074;
  wire [7:0] sel_551075;
  wire [7:0] add_551078;
  wire [7:0] sel_551079;
  wire [7:0] add_551082;
  wire [7:0] sel_551083;
  wire [7:0] add_551086;
  wire [7:0] sel_551087;
  wire [7:0] add_551090;
  wire [7:0] sel_551091;
  wire [7:0] add_551094;
  wire [7:0] sel_551095;
  wire [7:0] add_551098;
  wire [7:0] sel_551099;
  wire [7:0] add_551102;
  wire [7:0] sel_551103;
  wire [7:0] add_551106;
  wire [7:0] sel_551107;
  wire [7:0] add_551110;
  wire [7:0] sel_551111;
  wire [7:0] add_551114;
  wire [7:0] sel_551115;
  wire [7:0] add_551118;
  wire [7:0] sel_551119;
  wire [7:0] add_551122;
  wire [7:0] sel_551123;
  wire [7:0] add_551126;
  wire [7:0] sel_551127;
  wire [7:0] add_551130;
  wire [7:0] sel_551131;
  wire [7:0] add_551134;
  wire [7:0] sel_551135;
  wire [7:0] add_551138;
  wire [7:0] sel_551139;
  wire [7:0] add_551142;
  wire [7:0] sel_551143;
  wire [7:0] add_551146;
  wire [7:0] sel_551147;
  wire [7:0] add_551150;
  wire [7:0] sel_551151;
  wire [7:0] add_551154;
  wire [7:0] sel_551155;
  wire [7:0] add_551158;
  wire [7:0] sel_551159;
  wire [7:0] add_551162;
  wire [7:0] sel_551163;
  wire [7:0] add_551166;
  wire [7:0] sel_551167;
  wire [7:0] add_551170;
  wire [7:0] sel_551171;
  wire [7:0] add_551174;
  wire [7:0] sel_551175;
  wire [7:0] add_551178;
  wire [7:0] sel_551179;
  wire [7:0] add_551182;
  wire [7:0] sel_551183;
  wire [7:0] add_551186;
  wire [7:0] sel_551187;
  wire [7:0] add_551190;
  wire [7:0] sel_551191;
  wire [7:0] add_551194;
  wire [7:0] sel_551195;
  wire [7:0] add_551198;
  wire [7:0] sel_551199;
  wire [7:0] add_551202;
  wire [7:0] sel_551203;
  wire [7:0] add_551206;
  wire [7:0] sel_551207;
  wire [7:0] add_551210;
  wire [7:0] sel_551211;
  wire [7:0] add_551214;
  wire [7:0] sel_551215;
  wire [7:0] add_551218;
  wire [7:0] sel_551219;
  wire [7:0] add_551222;
  wire [7:0] sel_551223;
  wire [7:0] add_551226;
  wire [7:0] sel_551227;
  wire [7:0] add_551230;
  wire [7:0] sel_551231;
  wire [7:0] add_551234;
  wire [7:0] sel_551235;
  wire [7:0] add_551238;
  wire [7:0] sel_551239;
  wire [7:0] add_551242;
  wire [7:0] sel_551243;
  wire [7:0] add_551246;
  wire [7:0] sel_551247;
  wire [7:0] add_551250;
  wire [7:0] sel_551251;
  wire [7:0] add_551254;
  wire [7:0] sel_551255;
  wire [7:0] add_551258;
  wire [7:0] sel_551259;
  wire [7:0] add_551262;
  wire [7:0] sel_551263;
  wire [7:0] add_551266;
  wire [7:0] sel_551267;
  wire [7:0] add_551270;
  wire [7:0] sel_551271;
  wire [7:0] add_551274;
  wire [7:0] sel_551275;
  wire [7:0] add_551278;
  wire [7:0] sel_551279;
  wire [7:0] add_551282;
  wire [7:0] sel_551283;
  wire [7:0] add_551286;
  wire [7:0] sel_551287;
  wire [7:0] add_551290;
  wire [7:0] sel_551291;
  wire [7:0] add_551294;
  wire [7:0] sel_551295;
  wire [7:0] add_551298;
  wire [7:0] sel_551299;
  wire [7:0] add_551302;
  wire [7:0] sel_551303;
  wire [7:0] add_551306;
  wire [7:0] sel_551307;
  wire [7:0] add_551310;
  wire [7:0] sel_551311;
  wire [7:0] add_551314;
  wire [7:0] sel_551315;
  wire [7:0] add_551318;
  wire [7:0] sel_551319;
  wire [7:0] add_551322;
  wire [7:0] sel_551323;
  wire [7:0] add_551326;
  wire [7:0] sel_551327;
  wire [7:0] add_551330;
  wire [7:0] sel_551331;
  wire [7:0] add_551334;
  wire [7:0] sel_551335;
  wire [7:0] add_551338;
  wire [7:0] sel_551339;
  wire [7:0] add_551342;
  wire [7:0] sel_551343;
  wire [7:0] add_551346;
  wire [7:0] sel_551347;
  wire [7:0] add_551350;
  wire [7:0] sel_551351;
  wire [7:0] add_551354;
  wire [7:0] sel_551355;
  wire [7:0] add_551358;
  wire [7:0] sel_551359;
  wire [7:0] add_551363;
  wire [15:0] array_index_551364;
  wire [7:0] sel_551365;
  wire [7:0] add_551368;
  wire [7:0] sel_551369;
  wire [7:0] add_551372;
  wire [7:0] sel_551373;
  wire [7:0] add_551376;
  wire [7:0] sel_551377;
  wire [7:0] add_551380;
  wire [7:0] sel_551381;
  wire [7:0] add_551384;
  wire [7:0] sel_551385;
  wire [7:0] add_551388;
  wire [7:0] sel_551389;
  wire [7:0] add_551392;
  wire [7:0] sel_551393;
  wire [7:0] add_551396;
  wire [7:0] sel_551397;
  wire [7:0] add_551400;
  wire [7:0] sel_551401;
  wire [7:0] add_551404;
  wire [7:0] sel_551405;
  wire [7:0] add_551408;
  wire [7:0] sel_551409;
  wire [7:0] add_551412;
  wire [7:0] sel_551413;
  wire [7:0] add_551416;
  wire [7:0] sel_551417;
  wire [7:0] add_551420;
  wire [7:0] sel_551421;
  wire [7:0] add_551424;
  wire [7:0] sel_551425;
  wire [7:0] add_551428;
  wire [7:0] sel_551429;
  wire [7:0] add_551432;
  wire [7:0] sel_551433;
  wire [7:0] add_551436;
  wire [7:0] sel_551437;
  wire [7:0] add_551440;
  wire [7:0] sel_551441;
  wire [7:0] add_551444;
  wire [7:0] sel_551445;
  wire [7:0] add_551448;
  wire [7:0] sel_551449;
  wire [7:0] add_551452;
  wire [7:0] sel_551453;
  wire [7:0] add_551456;
  wire [7:0] sel_551457;
  wire [7:0] add_551460;
  wire [7:0] sel_551461;
  wire [7:0] add_551464;
  wire [7:0] sel_551465;
  wire [7:0] add_551468;
  wire [7:0] sel_551469;
  wire [7:0] add_551472;
  wire [7:0] sel_551473;
  wire [7:0] add_551476;
  wire [7:0] sel_551477;
  wire [7:0] add_551480;
  wire [7:0] sel_551481;
  wire [7:0] add_551484;
  wire [7:0] sel_551485;
  wire [7:0] add_551488;
  wire [7:0] sel_551489;
  wire [7:0] add_551492;
  wire [7:0] sel_551493;
  wire [7:0] add_551496;
  wire [7:0] sel_551497;
  wire [7:0] add_551500;
  wire [7:0] sel_551501;
  wire [7:0] add_551504;
  wire [7:0] sel_551505;
  wire [7:0] add_551508;
  wire [7:0] sel_551509;
  wire [7:0] add_551512;
  wire [7:0] sel_551513;
  wire [7:0] add_551516;
  wire [7:0] sel_551517;
  wire [7:0] add_551520;
  wire [7:0] sel_551521;
  wire [7:0] add_551524;
  wire [7:0] sel_551525;
  wire [7:0] add_551528;
  wire [7:0] sel_551529;
  wire [7:0] add_551532;
  wire [7:0] sel_551533;
  wire [7:0] add_551536;
  wire [7:0] sel_551537;
  wire [7:0] add_551540;
  wire [7:0] sel_551541;
  wire [7:0] add_551544;
  wire [7:0] sel_551545;
  wire [7:0] add_551548;
  wire [7:0] sel_551549;
  wire [7:0] add_551552;
  wire [7:0] sel_551553;
  wire [7:0] add_551556;
  wire [7:0] sel_551557;
  wire [7:0] add_551560;
  wire [7:0] sel_551561;
  wire [7:0] add_551564;
  wire [7:0] sel_551565;
  wire [7:0] add_551568;
  wire [7:0] sel_551569;
  wire [7:0] add_551572;
  wire [7:0] sel_551573;
  wire [7:0] add_551576;
  wire [7:0] sel_551577;
  wire [7:0] add_551580;
  wire [7:0] sel_551581;
  wire [7:0] add_551584;
  wire [7:0] sel_551585;
  wire [7:0] add_551588;
  wire [7:0] sel_551589;
  wire [7:0] add_551592;
  wire [7:0] sel_551593;
  wire [7:0] add_551596;
  wire [7:0] sel_551597;
  wire [7:0] add_551600;
  wire [7:0] sel_551601;
  wire [7:0] add_551604;
  wire [7:0] sel_551605;
  wire [7:0] add_551608;
  wire [7:0] sel_551609;
  wire [7:0] add_551612;
  wire [7:0] sel_551613;
  wire [7:0] add_551616;
  wire [7:0] sel_551617;
  wire [7:0] add_551620;
  wire [7:0] sel_551621;
  wire [7:0] add_551624;
  wire [7:0] sel_551625;
  wire [7:0] add_551628;
  wire [7:0] sel_551629;
  wire [7:0] add_551632;
  wire [7:0] sel_551633;
  wire [7:0] add_551636;
  wire [7:0] sel_551637;
  wire [7:0] add_551640;
  wire [7:0] sel_551641;
  wire [7:0] add_551644;
  wire [7:0] sel_551645;
  wire [7:0] add_551648;
  wire [7:0] sel_551649;
  wire [7:0] add_551652;
  wire [7:0] sel_551653;
  wire [7:0] add_551656;
  wire [7:0] sel_551657;
  wire [7:0] add_551660;
  wire [7:0] sel_551661;
  wire [7:0] add_551665;
  wire [15:0] array_index_551666;
  wire [7:0] sel_551667;
  wire [7:0] add_551670;
  wire [7:0] sel_551671;
  wire [7:0] add_551674;
  wire [7:0] sel_551675;
  wire [7:0] add_551678;
  wire [7:0] sel_551679;
  wire [7:0] add_551682;
  wire [7:0] sel_551683;
  wire [7:0] add_551686;
  wire [7:0] sel_551687;
  wire [7:0] add_551690;
  wire [7:0] sel_551691;
  wire [7:0] add_551694;
  wire [7:0] sel_551695;
  wire [7:0] add_551698;
  wire [7:0] sel_551699;
  wire [7:0] add_551702;
  wire [7:0] sel_551703;
  wire [7:0] add_551706;
  wire [7:0] sel_551707;
  wire [7:0] add_551710;
  wire [7:0] sel_551711;
  wire [7:0] add_551714;
  wire [7:0] sel_551715;
  wire [7:0] add_551718;
  wire [7:0] sel_551719;
  wire [7:0] add_551722;
  wire [7:0] sel_551723;
  wire [7:0] add_551726;
  wire [7:0] sel_551727;
  wire [7:0] add_551730;
  wire [7:0] sel_551731;
  wire [7:0] add_551734;
  wire [7:0] sel_551735;
  wire [7:0] add_551738;
  wire [7:0] sel_551739;
  wire [7:0] add_551742;
  wire [7:0] sel_551743;
  wire [7:0] add_551746;
  wire [7:0] sel_551747;
  wire [7:0] add_551750;
  wire [7:0] sel_551751;
  wire [7:0] add_551754;
  wire [7:0] sel_551755;
  wire [7:0] add_551758;
  wire [7:0] sel_551759;
  wire [7:0] add_551762;
  wire [7:0] sel_551763;
  wire [7:0] add_551766;
  wire [7:0] sel_551767;
  wire [7:0] add_551770;
  wire [7:0] sel_551771;
  wire [7:0] add_551774;
  wire [7:0] sel_551775;
  wire [7:0] add_551778;
  wire [7:0] sel_551779;
  wire [7:0] add_551782;
  wire [7:0] sel_551783;
  wire [7:0] add_551786;
  wire [7:0] sel_551787;
  wire [7:0] add_551790;
  wire [7:0] sel_551791;
  wire [7:0] add_551794;
  wire [7:0] sel_551795;
  wire [7:0] add_551798;
  wire [7:0] sel_551799;
  wire [7:0] add_551802;
  wire [7:0] sel_551803;
  wire [7:0] add_551806;
  wire [7:0] sel_551807;
  wire [7:0] add_551810;
  wire [7:0] sel_551811;
  wire [7:0] add_551814;
  wire [7:0] sel_551815;
  wire [7:0] add_551818;
  wire [7:0] sel_551819;
  wire [7:0] add_551822;
  wire [7:0] sel_551823;
  wire [7:0] add_551826;
  wire [7:0] sel_551827;
  wire [7:0] add_551830;
  wire [7:0] sel_551831;
  wire [7:0] add_551834;
  wire [7:0] sel_551835;
  wire [7:0] add_551838;
  wire [7:0] sel_551839;
  wire [7:0] add_551842;
  wire [7:0] sel_551843;
  wire [7:0] add_551846;
  wire [7:0] sel_551847;
  wire [7:0] add_551850;
  wire [7:0] sel_551851;
  wire [7:0] add_551854;
  wire [7:0] sel_551855;
  wire [7:0] add_551858;
  wire [7:0] sel_551859;
  wire [7:0] add_551862;
  wire [7:0] sel_551863;
  wire [7:0] add_551866;
  wire [7:0] sel_551867;
  wire [7:0] add_551870;
  wire [7:0] sel_551871;
  wire [7:0] add_551874;
  wire [7:0] sel_551875;
  wire [7:0] add_551878;
  wire [7:0] sel_551879;
  wire [7:0] add_551882;
  wire [7:0] sel_551883;
  wire [7:0] add_551886;
  wire [7:0] sel_551887;
  wire [7:0] add_551890;
  wire [7:0] sel_551891;
  wire [7:0] add_551894;
  wire [7:0] sel_551895;
  wire [7:0] add_551898;
  wire [7:0] sel_551899;
  wire [7:0] add_551902;
  wire [7:0] sel_551903;
  wire [7:0] add_551906;
  wire [7:0] sel_551907;
  wire [7:0] add_551910;
  wire [7:0] sel_551911;
  wire [7:0] add_551914;
  wire [7:0] sel_551915;
  wire [7:0] add_551918;
  wire [7:0] sel_551919;
  wire [7:0] add_551922;
  wire [7:0] sel_551923;
  wire [7:0] add_551926;
  wire [7:0] sel_551927;
  wire [7:0] add_551930;
  wire [7:0] sel_551931;
  wire [7:0] add_551934;
  wire [7:0] sel_551935;
  wire [7:0] add_551938;
  wire [7:0] sel_551939;
  wire [7:0] add_551942;
  wire [7:0] sel_551943;
  wire [7:0] add_551946;
  wire [7:0] sel_551947;
  wire [7:0] add_551950;
  wire [7:0] sel_551951;
  wire [7:0] add_551954;
  wire [7:0] sel_551955;
  wire [7:0] add_551958;
  wire [7:0] sel_551959;
  wire [7:0] add_551962;
  wire [7:0] sel_551963;
  wire [7:0] add_551967;
  wire [15:0] array_index_551968;
  wire [7:0] sel_551969;
  wire [7:0] add_551972;
  wire [7:0] sel_551973;
  wire [7:0] add_551976;
  wire [7:0] sel_551977;
  wire [7:0] add_551980;
  wire [7:0] sel_551981;
  wire [7:0] add_551984;
  wire [7:0] sel_551985;
  wire [7:0] add_551988;
  wire [7:0] sel_551989;
  wire [7:0] add_551992;
  wire [7:0] sel_551993;
  wire [7:0] add_551996;
  wire [7:0] sel_551997;
  wire [7:0] add_552000;
  wire [7:0] sel_552001;
  wire [7:0] add_552004;
  wire [7:0] sel_552005;
  wire [7:0] add_552008;
  wire [7:0] sel_552009;
  wire [7:0] add_552012;
  wire [7:0] sel_552013;
  wire [7:0] add_552016;
  wire [7:0] sel_552017;
  wire [7:0] add_552020;
  wire [7:0] sel_552021;
  wire [7:0] add_552024;
  wire [7:0] sel_552025;
  wire [7:0] add_552028;
  wire [7:0] sel_552029;
  wire [7:0] add_552032;
  wire [7:0] sel_552033;
  wire [7:0] add_552036;
  wire [7:0] sel_552037;
  wire [7:0] add_552040;
  wire [7:0] sel_552041;
  wire [7:0] add_552044;
  wire [7:0] sel_552045;
  wire [7:0] add_552048;
  wire [7:0] sel_552049;
  wire [7:0] add_552052;
  wire [7:0] sel_552053;
  wire [7:0] add_552056;
  wire [7:0] sel_552057;
  wire [7:0] add_552060;
  wire [7:0] sel_552061;
  wire [7:0] add_552064;
  wire [7:0] sel_552065;
  wire [7:0] add_552068;
  wire [7:0] sel_552069;
  wire [7:0] add_552072;
  wire [7:0] sel_552073;
  wire [7:0] add_552076;
  wire [7:0] sel_552077;
  wire [7:0] add_552080;
  wire [7:0] sel_552081;
  wire [7:0] add_552084;
  wire [7:0] sel_552085;
  wire [7:0] add_552088;
  wire [7:0] sel_552089;
  wire [7:0] add_552092;
  wire [7:0] sel_552093;
  wire [7:0] add_552096;
  wire [7:0] sel_552097;
  wire [7:0] add_552100;
  wire [7:0] sel_552101;
  wire [7:0] add_552104;
  wire [7:0] sel_552105;
  wire [7:0] add_552108;
  wire [7:0] sel_552109;
  wire [7:0] add_552112;
  wire [7:0] sel_552113;
  wire [7:0] add_552116;
  wire [7:0] sel_552117;
  wire [7:0] add_552120;
  wire [7:0] sel_552121;
  wire [7:0] add_552124;
  wire [7:0] sel_552125;
  wire [7:0] add_552128;
  wire [7:0] sel_552129;
  wire [7:0] add_552132;
  wire [7:0] sel_552133;
  wire [7:0] add_552136;
  wire [7:0] sel_552137;
  wire [7:0] add_552140;
  wire [7:0] sel_552141;
  wire [7:0] add_552144;
  wire [7:0] sel_552145;
  wire [7:0] add_552148;
  wire [7:0] sel_552149;
  wire [7:0] add_552152;
  wire [7:0] sel_552153;
  wire [7:0] add_552156;
  wire [7:0] sel_552157;
  wire [7:0] add_552160;
  wire [7:0] sel_552161;
  wire [7:0] add_552164;
  wire [7:0] sel_552165;
  wire [7:0] add_552168;
  wire [7:0] sel_552169;
  wire [7:0] add_552172;
  wire [7:0] sel_552173;
  wire [7:0] add_552176;
  wire [7:0] sel_552177;
  wire [7:0] add_552180;
  wire [7:0] sel_552181;
  wire [7:0] add_552184;
  wire [7:0] sel_552185;
  wire [7:0] add_552188;
  wire [7:0] sel_552189;
  wire [7:0] add_552192;
  wire [7:0] sel_552193;
  wire [7:0] add_552196;
  wire [7:0] sel_552197;
  wire [7:0] add_552200;
  wire [7:0] sel_552201;
  wire [7:0] add_552204;
  wire [7:0] sel_552205;
  wire [7:0] add_552208;
  wire [7:0] sel_552209;
  wire [7:0] add_552212;
  wire [7:0] sel_552213;
  wire [7:0] add_552216;
  wire [7:0] sel_552217;
  wire [7:0] add_552220;
  wire [7:0] sel_552221;
  wire [7:0] add_552224;
  wire [7:0] sel_552225;
  wire [7:0] add_552228;
  wire [7:0] sel_552229;
  wire [7:0] add_552232;
  wire [7:0] sel_552233;
  wire [7:0] add_552236;
  wire [7:0] sel_552237;
  wire [7:0] add_552240;
  wire [7:0] sel_552241;
  wire [7:0] add_552244;
  wire [7:0] sel_552245;
  wire [7:0] add_552248;
  wire [7:0] sel_552249;
  wire [7:0] add_552252;
  wire [7:0] sel_552253;
  wire [7:0] add_552256;
  wire [7:0] sel_552257;
  wire [7:0] add_552260;
  wire [7:0] sel_552261;
  wire [7:0] add_552264;
  wire [7:0] sel_552265;
  wire [7:0] add_552269;
  wire [15:0] array_index_552270;
  wire [7:0] sel_552271;
  wire [7:0] add_552274;
  wire [7:0] sel_552275;
  wire [7:0] add_552278;
  wire [7:0] sel_552279;
  wire [7:0] add_552282;
  wire [7:0] sel_552283;
  wire [7:0] add_552286;
  wire [7:0] sel_552287;
  wire [7:0] add_552290;
  wire [7:0] sel_552291;
  wire [7:0] add_552294;
  wire [7:0] sel_552295;
  wire [7:0] add_552298;
  wire [7:0] sel_552299;
  wire [7:0] add_552302;
  wire [7:0] sel_552303;
  wire [7:0] add_552306;
  wire [7:0] sel_552307;
  wire [7:0] add_552310;
  wire [7:0] sel_552311;
  wire [7:0] add_552314;
  wire [7:0] sel_552315;
  wire [7:0] add_552318;
  wire [7:0] sel_552319;
  wire [7:0] add_552322;
  wire [7:0] sel_552323;
  wire [7:0] add_552326;
  wire [7:0] sel_552327;
  wire [7:0] add_552330;
  wire [7:0] sel_552331;
  wire [7:0] add_552334;
  wire [7:0] sel_552335;
  wire [7:0] add_552338;
  wire [7:0] sel_552339;
  wire [7:0] add_552342;
  wire [7:0] sel_552343;
  wire [7:0] add_552346;
  wire [7:0] sel_552347;
  wire [7:0] add_552350;
  wire [7:0] sel_552351;
  wire [7:0] add_552354;
  wire [7:0] sel_552355;
  wire [7:0] add_552358;
  wire [7:0] sel_552359;
  wire [7:0] add_552362;
  wire [7:0] sel_552363;
  wire [7:0] add_552366;
  wire [7:0] sel_552367;
  wire [7:0] add_552370;
  wire [7:0] sel_552371;
  wire [7:0] add_552374;
  wire [7:0] sel_552375;
  wire [7:0] add_552378;
  wire [7:0] sel_552379;
  wire [7:0] add_552382;
  wire [7:0] sel_552383;
  wire [7:0] add_552386;
  wire [7:0] sel_552387;
  wire [7:0] add_552390;
  wire [7:0] sel_552391;
  wire [7:0] add_552394;
  wire [7:0] sel_552395;
  wire [7:0] add_552398;
  wire [7:0] sel_552399;
  wire [7:0] add_552402;
  wire [7:0] sel_552403;
  wire [7:0] add_552406;
  wire [7:0] sel_552407;
  wire [7:0] add_552410;
  wire [7:0] sel_552411;
  wire [7:0] add_552414;
  wire [7:0] sel_552415;
  wire [7:0] add_552418;
  wire [7:0] sel_552419;
  wire [7:0] add_552422;
  wire [7:0] sel_552423;
  wire [7:0] add_552426;
  wire [7:0] sel_552427;
  wire [7:0] add_552430;
  wire [7:0] sel_552431;
  wire [7:0] add_552434;
  wire [7:0] sel_552435;
  wire [7:0] add_552438;
  wire [7:0] sel_552439;
  wire [7:0] add_552442;
  wire [7:0] sel_552443;
  wire [7:0] add_552446;
  wire [7:0] sel_552447;
  wire [7:0] add_552450;
  wire [7:0] sel_552451;
  wire [7:0] add_552454;
  wire [7:0] sel_552455;
  wire [7:0] add_552458;
  wire [7:0] sel_552459;
  wire [7:0] add_552462;
  wire [7:0] sel_552463;
  wire [7:0] add_552466;
  wire [7:0] sel_552467;
  wire [7:0] add_552470;
  wire [7:0] sel_552471;
  wire [7:0] add_552474;
  wire [7:0] sel_552475;
  wire [7:0] add_552478;
  wire [7:0] sel_552479;
  wire [7:0] add_552482;
  wire [7:0] sel_552483;
  wire [7:0] add_552486;
  wire [7:0] sel_552487;
  wire [7:0] add_552490;
  wire [7:0] sel_552491;
  wire [7:0] add_552494;
  wire [7:0] sel_552495;
  wire [7:0] add_552498;
  wire [7:0] sel_552499;
  wire [7:0] add_552502;
  wire [7:0] sel_552503;
  wire [7:0] add_552506;
  wire [7:0] sel_552507;
  wire [7:0] add_552510;
  wire [7:0] sel_552511;
  wire [7:0] add_552514;
  wire [7:0] sel_552515;
  wire [7:0] add_552518;
  wire [7:0] sel_552519;
  wire [7:0] add_552522;
  wire [7:0] sel_552523;
  wire [7:0] add_552526;
  wire [7:0] sel_552527;
  wire [7:0] add_552530;
  wire [7:0] sel_552531;
  wire [7:0] add_552534;
  wire [7:0] sel_552535;
  wire [7:0] add_552538;
  wire [7:0] sel_552539;
  wire [7:0] add_552542;
  wire [7:0] sel_552543;
  wire [7:0] add_552546;
  wire [7:0] sel_552547;
  wire [7:0] add_552550;
  wire [7:0] sel_552551;
  wire [7:0] add_552554;
  wire [7:0] sel_552555;
  wire [7:0] add_552558;
  wire [7:0] sel_552559;
  wire [7:0] add_552562;
  wire [7:0] sel_552563;
  wire [7:0] add_552566;
  wire [7:0] sel_552567;
  wire [7:0] add_552571;
  wire [15:0] array_index_552572;
  wire [7:0] sel_552573;
  wire [7:0] add_552576;
  wire [7:0] sel_552577;
  wire [7:0] add_552580;
  wire [7:0] sel_552581;
  wire [7:0] add_552584;
  wire [7:0] sel_552585;
  wire [7:0] add_552588;
  wire [7:0] sel_552589;
  wire [7:0] add_552592;
  wire [7:0] sel_552593;
  wire [7:0] add_552596;
  wire [7:0] sel_552597;
  wire [7:0] add_552600;
  wire [7:0] sel_552601;
  wire [7:0] add_552604;
  wire [7:0] sel_552605;
  wire [7:0] add_552608;
  wire [7:0] sel_552609;
  wire [7:0] add_552612;
  wire [7:0] sel_552613;
  wire [7:0] add_552616;
  wire [7:0] sel_552617;
  wire [7:0] add_552620;
  wire [7:0] sel_552621;
  wire [7:0] add_552624;
  wire [7:0] sel_552625;
  wire [7:0] add_552628;
  wire [7:0] sel_552629;
  wire [7:0] add_552632;
  wire [7:0] sel_552633;
  wire [7:0] add_552636;
  wire [7:0] sel_552637;
  wire [7:0] add_552640;
  wire [7:0] sel_552641;
  wire [7:0] add_552644;
  wire [7:0] sel_552645;
  wire [7:0] add_552648;
  wire [7:0] sel_552649;
  wire [7:0] add_552652;
  wire [7:0] sel_552653;
  wire [7:0] add_552656;
  wire [7:0] sel_552657;
  wire [7:0] add_552660;
  wire [7:0] sel_552661;
  wire [7:0] add_552664;
  wire [7:0] sel_552665;
  wire [7:0] add_552668;
  wire [7:0] sel_552669;
  wire [7:0] add_552672;
  wire [7:0] sel_552673;
  wire [7:0] add_552676;
  wire [7:0] sel_552677;
  wire [7:0] add_552680;
  wire [7:0] sel_552681;
  wire [7:0] add_552684;
  wire [7:0] sel_552685;
  wire [7:0] add_552688;
  wire [7:0] sel_552689;
  wire [7:0] add_552692;
  wire [7:0] sel_552693;
  wire [7:0] add_552696;
  wire [7:0] sel_552697;
  wire [7:0] add_552700;
  wire [7:0] sel_552701;
  wire [7:0] add_552704;
  wire [7:0] sel_552705;
  wire [7:0] add_552708;
  wire [7:0] sel_552709;
  wire [7:0] add_552712;
  wire [7:0] sel_552713;
  wire [7:0] add_552716;
  wire [7:0] sel_552717;
  wire [7:0] add_552720;
  wire [7:0] sel_552721;
  wire [7:0] add_552724;
  wire [7:0] sel_552725;
  wire [7:0] add_552728;
  wire [7:0] sel_552729;
  wire [7:0] add_552732;
  wire [7:0] sel_552733;
  wire [7:0] add_552736;
  wire [7:0] sel_552737;
  wire [7:0] add_552740;
  wire [7:0] sel_552741;
  wire [7:0] add_552744;
  wire [7:0] sel_552745;
  wire [7:0] add_552748;
  wire [7:0] sel_552749;
  wire [7:0] add_552752;
  wire [7:0] sel_552753;
  wire [7:0] add_552756;
  wire [7:0] sel_552757;
  wire [7:0] add_552760;
  wire [7:0] sel_552761;
  wire [7:0] add_552764;
  wire [7:0] sel_552765;
  wire [7:0] add_552768;
  wire [7:0] sel_552769;
  wire [7:0] add_552772;
  wire [7:0] sel_552773;
  wire [7:0] add_552776;
  wire [7:0] sel_552777;
  wire [7:0] add_552780;
  wire [7:0] sel_552781;
  wire [7:0] add_552784;
  wire [7:0] sel_552785;
  wire [7:0] add_552788;
  wire [7:0] sel_552789;
  wire [7:0] add_552792;
  wire [7:0] sel_552793;
  wire [7:0] add_552796;
  wire [7:0] sel_552797;
  wire [7:0] add_552800;
  wire [7:0] sel_552801;
  wire [7:0] add_552804;
  wire [7:0] sel_552805;
  wire [7:0] add_552808;
  wire [7:0] sel_552809;
  wire [7:0] add_552812;
  wire [7:0] sel_552813;
  wire [7:0] add_552816;
  wire [7:0] sel_552817;
  wire [7:0] add_552820;
  wire [7:0] sel_552821;
  wire [7:0] add_552824;
  wire [7:0] sel_552825;
  wire [7:0] add_552828;
  wire [7:0] sel_552829;
  wire [7:0] add_552832;
  wire [7:0] sel_552833;
  wire [7:0] add_552836;
  wire [7:0] sel_552837;
  wire [7:0] add_552840;
  wire [7:0] sel_552841;
  wire [7:0] add_552844;
  wire [7:0] sel_552845;
  wire [7:0] add_552848;
  wire [7:0] sel_552849;
  wire [7:0] add_552852;
  wire [7:0] sel_552853;
  wire [7:0] add_552856;
  wire [7:0] sel_552857;
  wire [7:0] add_552860;
  wire [7:0] sel_552861;
  wire [7:0] add_552864;
  wire [7:0] sel_552865;
  wire [7:0] add_552868;
  wire [7:0] sel_552869;
  wire [7:0] add_552873;
  wire [15:0] array_index_552874;
  wire [7:0] sel_552875;
  wire [7:0] add_552878;
  wire [7:0] sel_552879;
  wire [7:0] add_552882;
  wire [7:0] sel_552883;
  wire [7:0] add_552886;
  wire [7:0] sel_552887;
  wire [7:0] add_552890;
  wire [7:0] sel_552891;
  wire [7:0] add_552894;
  wire [7:0] sel_552895;
  wire [7:0] add_552898;
  wire [7:0] sel_552899;
  wire [7:0] add_552902;
  wire [7:0] sel_552903;
  wire [7:0] add_552906;
  wire [7:0] sel_552907;
  wire [7:0] add_552910;
  wire [7:0] sel_552911;
  wire [7:0] add_552914;
  wire [7:0] sel_552915;
  wire [7:0] add_552918;
  wire [7:0] sel_552919;
  wire [7:0] add_552922;
  wire [7:0] sel_552923;
  wire [7:0] add_552926;
  wire [7:0] sel_552927;
  wire [7:0] add_552930;
  wire [7:0] sel_552931;
  wire [7:0] add_552934;
  wire [7:0] sel_552935;
  wire [7:0] add_552938;
  wire [7:0] sel_552939;
  wire [7:0] add_552942;
  wire [7:0] sel_552943;
  wire [7:0] add_552946;
  wire [7:0] sel_552947;
  wire [7:0] add_552950;
  wire [7:0] sel_552951;
  wire [7:0] add_552954;
  wire [7:0] sel_552955;
  wire [7:0] add_552958;
  wire [7:0] sel_552959;
  wire [7:0] add_552962;
  wire [7:0] sel_552963;
  wire [7:0] add_552966;
  wire [7:0] sel_552967;
  wire [7:0] add_552970;
  wire [7:0] sel_552971;
  wire [7:0] add_552974;
  wire [7:0] sel_552975;
  wire [7:0] add_552978;
  wire [7:0] sel_552979;
  wire [7:0] add_552982;
  wire [7:0] sel_552983;
  wire [7:0] add_552986;
  wire [7:0] sel_552987;
  wire [7:0] add_552990;
  wire [7:0] sel_552991;
  wire [7:0] add_552994;
  wire [7:0] sel_552995;
  wire [7:0] add_552998;
  wire [7:0] sel_552999;
  wire [7:0] add_553002;
  wire [7:0] sel_553003;
  wire [7:0] add_553006;
  wire [7:0] sel_553007;
  wire [7:0] add_553010;
  wire [7:0] sel_553011;
  wire [7:0] add_553014;
  wire [7:0] sel_553015;
  wire [7:0] add_553018;
  wire [7:0] sel_553019;
  wire [7:0] add_553022;
  wire [7:0] sel_553023;
  wire [7:0] add_553026;
  wire [7:0] sel_553027;
  wire [7:0] add_553030;
  wire [7:0] sel_553031;
  wire [7:0] add_553034;
  wire [7:0] sel_553035;
  wire [7:0] add_553038;
  wire [7:0] sel_553039;
  wire [7:0] add_553042;
  wire [7:0] sel_553043;
  wire [7:0] add_553046;
  wire [7:0] sel_553047;
  wire [7:0] add_553050;
  wire [7:0] sel_553051;
  wire [7:0] add_553054;
  wire [7:0] sel_553055;
  wire [7:0] add_553058;
  wire [7:0] sel_553059;
  wire [7:0] add_553062;
  wire [7:0] sel_553063;
  wire [7:0] add_553066;
  wire [7:0] sel_553067;
  wire [7:0] add_553070;
  wire [7:0] sel_553071;
  wire [7:0] add_553074;
  wire [7:0] sel_553075;
  wire [7:0] add_553078;
  wire [7:0] sel_553079;
  wire [7:0] add_553082;
  wire [7:0] sel_553083;
  wire [7:0] add_553086;
  wire [7:0] sel_553087;
  wire [7:0] add_553090;
  wire [7:0] sel_553091;
  wire [7:0] add_553094;
  wire [7:0] sel_553095;
  wire [7:0] add_553098;
  wire [7:0] sel_553099;
  wire [7:0] add_553102;
  wire [7:0] sel_553103;
  wire [7:0] add_553106;
  wire [7:0] sel_553107;
  wire [7:0] add_553110;
  wire [7:0] sel_553111;
  wire [7:0] add_553114;
  wire [7:0] sel_553115;
  wire [7:0] add_553118;
  wire [7:0] sel_553119;
  wire [7:0] add_553122;
  wire [7:0] sel_553123;
  wire [7:0] add_553126;
  wire [7:0] sel_553127;
  wire [7:0] add_553130;
  wire [7:0] sel_553131;
  wire [7:0] add_553134;
  wire [7:0] sel_553135;
  wire [7:0] add_553138;
  wire [7:0] sel_553139;
  wire [7:0] add_553142;
  wire [7:0] sel_553143;
  wire [7:0] add_553146;
  wire [7:0] sel_553147;
  wire [7:0] add_553150;
  wire [7:0] sel_553151;
  wire [7:0] add_553154;
  wire [7:0] sel_553155;
  wire [7:0] add_553158;
  wire [7:0] sel_553159;
  wire [7:0] add_553162;
  wire [7:0] sel_553163;
  wire [7:0] add_553166;
  wire [7:0] sel_553167;
  wire [7:0] add_553170;
  wire [7:0] sel_553171;
  wire [7:0] add_553175;
  wire [15:0] array_index_553176;
  wire [7:0] sel_553177;
  wire [7:0] add_553180;
  wire [7:0] sel_553181;
  wire [7:0] add_553184;
  wire [7:0] sel_553185;
  wire [7:0] add_553188;
  wire [7:0] sel_553189;
  wire [7:0] add_553192;
  wire [7:0] sel_553193;
  wire [7:0] add_553196;
  wire [7:0] sel_553197;
  wire [7:0] add_553200;
  wire [7:0] sel_553201;
  wire [7:0] add_553204;
  wire [7:0] sel_553205;
  wire [7:0] add_553208;
  wire [7:0] sel_553209;
  wire [7:0] add_553212;
  wire [7:0] sel_553213;
  wire [7:0] add_553216;
  wire [7:0] sel_553217;
  wire [7:0] add_553220;
  wire [7:0] sel_553221;
  wire [7:0] add_553224;
  wire [7:0] sel_553225;
  wire [7:0] add_553228;
  wire [7:0] sel_553229;
  wire [7:0] add_553232;
  wire [7:0] sel_553233;
  wire [7:0] add_553236;
  wire [7:0] sel_553237;
  wire [7:0] add_553240;
  wire [7:0] sel_553241;
  wire [7:0] add_553244;
  wire [7:0] sel_553245;
  wire [7:0] add_553248;
  wire [7:0] sel_553249;
  wire [7:0] add_553252;
  wire [7:0] sel_553253;
  wire [7:0] add_553256;
  wire [7:0] sel_553257;
  wire [7:0] add_553260;
  wire [7:0] sel_553261;
  wire [7:0] add_553264;
  wire [7:0] sel_553265;
  wire [7:0] add_553268;
  wire [7:0] sel_553269;
  wire [7:0] add_553272;
  wire [7:0] sel_553273;
  wire [7:0] add_553276;
  wire [7:0] sel_553277;
  wire [7:0] add_553280;
  wire [7:0] sel_553281;
  wire [7:0] add_553284;
  wire [7:0] sel_553285;
  wire [7:0] add_553288;
  wire [7:0] sel_553289;
  wire [7:0] add_553292;
  wire [7:0] sel_553293;
  wire [7:0] add_553296;
  wire [7:0] sel_553297;
  wire [7:0] add_553300;
  wire [7:0] sel_553301;
  wire [7:0] add_553304;
  wire [7:0] sel_553305;
  wire [7:0] add_553308;
  wire [7:0] sel_553309;
  wire [7:0] add_553312;
  wire [7:0] sel_553313;
  wire [7:0] add_553316;
  wire [7:0] sel_553317;
  wire [7:0] add_553320;
  wire [7:0] sel_553321;
  wire [7:0] add_553324;
  wire [7:0] sel_553325;
  wire [7:0] add_553328;
  wire [7:0] sel_553329;
  wire [7:0] add_553332;
  wire [7:0] sel_553333;
  wire [7:0] add_553336;
  wire [7:0] sel_553337;
  wire [7:0] add_553340;
  wire [7:0] sel_553341;
  wire [7:0] add_553344;
  wire [7:0] sel_553345;
  wire [7:0] add_553348;
  wire [7:0] sel_553349;
  wire [7:0] add_553352;
  wire [7:0] sel_553353;
  wire [7:0] add_553356;
  wire [7:0] sel_553357;
  wire [7:0] add_553360;
  wire [7:0] sel_553361;
  wire [7:0] add_553364;
  wire [7:0] sel_553365;
  wire [7:0] add_553368;
  wire [7:0] sel_553369;
  wire [7:0] add_553372;
  wire [7:0] sel_553373;
  wire [7:0] add_553376;
  wire [7:0] sel_553377;
  wire [7:0] add_553380;
  wire [7:0] sel_553381;
  wire [7:0] add_553384;
  wire [7:0] sel_553385;
  wire [7:0] add_553388;
  wire [7:0] sel_553389;
  wire [7:0] add_553392;
  wire [7:0] sel_553393;
  wire [7:0] add_553396;
  wire [7:0] sel_553397;
  wire [7:0] add_553400;
  wire [7:0] sel_553401;
  wire [7:0] add_553404;
  wire [7:0] sel_553405;
  wire [7:0] add_553408;
  wire [7:0] sel_553409;
  wire [7:0] add_553412;
  wire [7:0] sel_553413;
  wire [7:0] add_553416;
  wire [7:0] sel_553417;
  wire [7:0] add_553420;
  wire [7:0] sel_553421;
  wire [7:0] add_553424;
  wire [7:0] sel_553425;
  wire [7:0] add_553428;
  wire [7:0] sel_553429;
  wire [7:0] add_553432;
  wire [7:0] sel_553433;
  wire [7:0] add_553436;
  wire [7:0] sel_553437;
  wire [7:0] add_553440;
  wire [7:0] sel_553441;
  wire [7:0] add_553444;
  wire [7:0] sel_553445;
  wire [7:0] add_553448;
  wire [7:0] sel_553449;
  wire [7:0] add_553452;
  wire [7:0] sel_553453;
  wire [7:0] add_553456;
  wire [7:0] sel_553457;
  wire [7:0] add_553460;
  wire [7:0] sel_553461;
  wire [7:0] add_553464;
  wire [7:0] sel_553465;
  wire [7:0] add_553468;
  wire [7:0] sel_553469;
  wire [7:0] add_553472;
  wire [7:0] sel_553473;
  wire [7:0] add_553477;
  wire [15:0] array_index_553478;
  wire [7:0] sel_553479;
  wire [7:0] add_553482;
  wire [7:0] sel_553483;
  wire [7:0] add_553486;
  wire [7:0] sel_553487;
  wire [7:0] add_553490;
  wire [7:0] sel_553491;
  wire [7:0] add_553494;
  wire [7:0] sel_553495;
  wire [7:0] add_553498;
  wire [7:0] sel_553499;
  wire [7:0] add_553502;
  wire [7:0] sel_553503;
  wire [7:0] add_553506;
  wire [7:0] sel_553507;
  wire [7:0] add_553510;
  wire [7:0] sel_553511;
  wire [7:0] add_553514;
  wire [7:0] sel_553515;
  wire [7:0] add_553518;
  wire [7:0] sel_553519;
  wire [7:0] add_553522;
  wire [7:0] sel_553523;
  wire [7:0] add_553526;
  wire [7:0] sel_553527;
  wire [7:0] add_553530;
  wire [7:0] sel_553531;
  wire [7:0] add_553534;
  wire [7:0] sel_553535;
  wire [7:0] add_553538;
  wire [7:0] sel_553539;
  wire [7:0] add_553542;
  wire [7:0] sel_553543;
  wire [7:0] add_553546;
  wire [7:0] sel_553547;
  wire [7:0] add_553550;
  wire [7:0] sel_553551;
  wire [7:0] add_553554;
  wire [7:0] sel_553555;
  wire [7:0] add_553558;
  wire [7:0] sel_553559;
  wire [7:0] add_553562;
  wire [7:0] sel_553563;
  wire [7:0] add_553566;
  wire [7:0] sel_553567;
  wire [7:0] add_553570;
  wire [7:0] sel_553571;
  wire [7:0] add_553574;
  wire [7:0] sel_553575;
  wire [7:0] add_553578;
  wire [7:0] sel_553579;
  wire [7:0] add_553582;
  wire [7:0] sel_553583;
  wire [7:0] add_553586;
  wire [7:0] sel_553587;
  wire [7:0] add_553590;
  wire [7:0] sel_553591;
  wire [7:0] add_553594;
  wire [7:0] sel_553595;
  wire [7:0] add_553598;
  wire [7:0] sel_553599;
  wire [7:0] add_553602;
  wire [7:0] sel_553603;
  wire [7:0] add_553606;
  wire [7:0] sel_553607;
  wire [7:0] add_553610;
  wire [7:0] sel_553611;
  wire [7:0] add_553614;
  wire [7:0] sel_553615;
  wire [7:0] add_553618;
  wire [7:0] sel_553619;
  wire [7:0] add_553622;
  wire [7:0] sel_553623;
  wire [7:0] add_553626;
  wire [7:0] sel_553627;
  wire [7:0] add_553630;
  wire [7:0] sel_553631;
  wire [7:0] add_553634;
  wire [7:0] sel_553635;
  wire [7:0] add_553638;
  wire [7:0] sel_553639;
  wire [7:0] add_553642;
  wire [7:0] sel_553643;
  wire [7:0] add_553646;
  wire [7:0] sel_553647;
  wire [7:0] add_553650;
  wire [7:0] sel_553651;
  wire [7:0] add_553654;
  wire [7:0] sel_553655;
  wire [7:0] add_553658;
  wire [7:0] sel_553659;
  wire [7:0] add_553662;
  wire [7:0] sel_553663;
  wire [7:0] add_553666;
  wire [7:0] sel_553667;
  wire [7:0] add_553670;
  wire [7:0] sel_553671;
  wire [7:0] add_553674;
  wire [7:0] sel_553675;
  wire [7:0] add_553678;
  wire [7:0] sel_553679;
  wire [7:0] add_553682;
  wire [7:0] sel_553683;
  wire [7:0] add_553686;
  wire [7:0] sel_553687;
  wire [7:0] add_553690;
  wire [7:0] sel_553691;
  wire [7:0] add_553694;
  wire [7:0] sel_553695;
  wire [7:0] add_553698;
  wire [7:0] sel_553699;
  wire [7:0] add_553702;
  wire [7:0] sel_553703;
  wire [7:0] add_553706;
  wire [7:0] sel_553707;
  wire [7:0] add_553710;
  wire [7:0] sel_553711;
  wire [7:0] add_553714;
  wire [7:0] sel_553715;
  wire [7:0] add_553718;
  wire [7:0] sel_553719;
  wire [7:0] add_553722;
  wire [7:0] sel_553723;
  wire [7:0] add_553726;
  wire [7:0] sel_553727;
  wire [7:0] add_553730;
  wire [7:0] sel_553731;
  wire [7:0] add_553734;
  wire [7:0] sel_553735;
  wire [7:0] add_553738;
  wire [7:0] sel_553739;
  wire [7:0] add_553742;
  wire [7:0] sel_553743;
  wire [7:0] add_553746;
  wire [7:0] sel_553747;
  wire [7:0] add_553750;
  wire [7:0] sel_553751;
  wire [7:0] add_553754;
  wire [7:0] sel_553755;
  wire [7:0] add_553758;
  wire [7:0] sel_553759;
  wire [7:0] add_553762;
  wire [7:0] sel_553763;
  wire [7:0] add_553766;
  wire [7:0] sel_553767;
  wire [7:0] add_553770;
  wire [7:0] sel_553771;
  wire [7:0] add_553774;
  wire [7:0] sel_553775;
  wire [7:0] add_553779;
  wire [15:0] array_index_553780;
  wire [7:0] sel_553781;
  wire [7:0] add_553784;
  wire [7:0] sel_553785;
  wire [7:0] add_553788;
  wire [7:0] sel_553789;
  wire [7:0] add_553792;
  wire [7:0] sel_553793;
  wire [7:0] add_553796;
  wire [7:0] sel_553797;
  wire [7:0] add_553800;
  wire [7:0] sel_553801;
  wire [7:0] add_553804;
  wire [7:0] sel_553805;
  wire [7:0] add_553808;
  wire [7:0] sel_553809;
  wire [7:0] add_553812;
  wire [7:0] sel_553813;
  wire [7:0] add_553816;
  wire [7:0] sel_553817;
  wire [7:0] add_553820;
  wire [7:0] sel_553821;
  wire [7:0] add_553824;
  wire [7:0] sel_553825;
  wire [7:0] add_553828;
  wire [7:0] sel_553829;
  wire [7:0] add_553832;
  wire [7:0] sel_553833;
  wire [7:0] add_553836;
  wire [7:0] sel_553837;
  wire [7:0] add_553840;
  wire [7:0] sel_553841;
  wire [7:0] add_553844;
  wire [7:0] sel_553845;
  wire [7:0] add_553848;
  wire [7:0] sel_553849;
  wire [7:0] add_553852;
  wire [7:0] sel_553853;
  wire [7:0] add_553856;
  wire [7:0] sel_553857;
  wire [7:0] add_553860;
  wire [7:0] sel_553861;
  wire [7:0] add_553864;
  wire [7:0] sel_553865;
  wire [7:0] add_553868;
  wire [7:0] sel_553869;
  wire [7:0] add_553872;
  wire [7:0] sel_553873;
  wire [7:0] add_553876;
  wire [7:0] sel_553877;
  wire [7:0] add_553880;
  wire [7:0] sel_553881;
  wire [7:0] add_553884;
  wire [7:0] sel_553885;
  wire [7:0] add_553888;
  wire [7:0] sel_553889;
  wire [7:0] add_553892;
  wire [7:0] sel_553893;
  wire [7:0] add_553896;
  wire [7:0] sel_553897;
  wire [7:0] add_553900;
  wire [7:0] sel_553901;
  wire [7:0] add_553904;
  wire [7:0] sel_553905;
  wire [7:0] add_553908;
  wire [7:0] sel_553909;
  wire [7:0] add_553912;
  wire [7:0] sel_553913;
  wire [7:0] add_553916;
  wire [7:0] sel_553917;
  wire [7:0] add_553920;
  wire [7:0] sel_553921;
  wire [7:0] add_553924;
  wire [7:0] sel_553925;
  wire [7:0] add_553928;
  wire [7:0] sel_553929;
  wire [7:0] add_553932;
  wire [7:0] sel_553933;
  wire [7:0] add_553936;
  wire [7:0] sel_553937;
  wire [7:0] add_553940;
  wire [7:0] sel_553941;
  wire [7:0] add_553944;
  wire [7:0] sel_553945;
  wire [7:0] add_553948;
  wire [7:0] sel_553949;
  wire [7:0] add_553952;
  wire [7:0] sel_553953;
  wire [7:0] add_553956;
  wire [7:0] sel_553957;
  wire [7:0] add_553960;
  wire [7:0] sel_553961;
  wire [7:0] add_553964;
  wire [7:0] sel_553965;
  wire [7:0] add_553968;
  wire [7:0] sel_553969;
  wire [7:0] add_553972;
  wire [7:0] sel_553973;
  wire [7:0] add_553976;
  wire [7:0] sel_553977;
  wire [7:0] add_553980;
  wire [7:0] sel_553981;
  wire [7:0] add_553984;
  wire [7:0] sel_553985;
  wire [7:0] add_553988;
  wire [7:0] sel_553989;
  wire [7:0] add_553992;
  wire [7:0] sel_553993;
  wire [7:0] add_553996;
  wire [7:0] sel_553997;
  wire [7:0] add_554000;
  wire [7:0] sel_554001;
  wire [7:0] add_554004;
  wire [7:0] sel_554005;
  wire [7:0] add_554008;
  wire [7:0] sel_554009;
  wire [7:0] add_554012;
  wire [7:0] sel_554013;
  wire [7:0] add_554016;
  wire [7:0] sel_554017;
  wire [7:0] add_554020;
  wire [7:0] sel_554021;
  wire [7:0] add_554024;
  wire [7:0] sel_554025;
  wire [7:0] add_554028;
  wire [7:0] sel_554029;
  wire [7:0] add_554032;
  wire [7:0] sel_554033;
  wire [7:0] add_554036;
  wire [7:0] sel_554037;
  wire [7:0] add_554040;
  wire [7:0] sel_554041;
  wire [7:0] add_554044;
  wire [7:0] sel_554045;
  wire [7:0] add_554048;
  wire [7:0] sel_554049;
  wire [7:0] add_554052;
  wire [7:0] sel_554053;
  wire [7:0] add_554056;
  wire [7:0] sel_554057;
  wire [7:0] add_554060;
  wire [7:0] sel_554061;
  wire [7:0] add_554064;
  wire [7:0] sel_554065;
  wire [7:0] add_554068;
  wire [7:0] sel_554069;
  wire [7:0] add_554072;
  wire [7:0] sel_554073;
  wire [7:0] add_554076;
  wire [7:0] sel_554077;
  wire [7:0] add_554081;
  wire [15:0] array_index_554082;
  wire [7:0] sel_554083;
  wire [7:0] add_554086;
  wire [7:0] sel_554087;
  wire [7:0] add_554090;
  wire [7:0] sel_554091;
  wire [7:0] add_554094;
  wire [7:0] sel_554095;
  wire [7:0] add_554098;
  wire [7:0] sel_554099;
  wire [7:0] add_554102;
  wire [7:0] sel_554103;
  wire [7:0] add_554106;
  wire [7:0] sel_554107;
  wire [7:0] add_554110;
  wire [7:0] sel_554111;
  wire [7:0] add_554114;
  wire [7:0] sel_554115;
  wire [7:0] add_554118;
  wire [7:0] sel_554119;
  wire [7:0] add_554122;
  wire [7:0] sel_554123;
  wire [7:0] add_554126;
  wire [7:0] sel_554127;
  wire [7:0] add_554130;
  wire [7:0] sel_554131;
  wire [7:0] add_554134;
  wire [7:0] sel_554135;
  wire [7:0] add_554138;
  wire [7:0] sel_554139;
  wire [7:0] add_554142;
  wire [7:0] sel_554143;
  wire [7:0] add_554146;
  wire [7:0] sel_554147;
  wire [7:0] add_554150;
  wire [7:0] sel_554151;
  wire [7:0] add_554154;
  wire [7:0] sel_554155;
  wire [7:0] add_554158;
  wire [7:0] sel_554159;
  wire [7:0] add_554162;
  wire [7:0] sel_554163;
  wire [7:0] add_554166;
  wire [7:0] sel_554167;
  wire [7:0] add_554170;
  wire [7:0] sel_554171;
  wire [7:0] add_554174;
  wire [7:0] sel_554175;
  wire [7:0] add_554178;
  wire [7:0] sel_554179;
  wire [7:0] add_554182;
  wire [7:0] sel_554183;
  wire [7:0] add_554186;
  wire [7:0] sel_554187;
  wire [7:0] add_554190;
  wire [7:0] sel_554191;
  wire [7:0] add_554194;
  wire [7:0] sel_554195;
  wire [7:0] add_554198;
  wire [7:0] sel_554199;
  wire [7:0] add_554202;
  wire [7:0] sel_554203;
  wire [7:0] add_554206;
  wire [7:0] sel_554207;
  wire [7:0] add_554210;
  wire [7:0] sel_554211;
  wire [7:0] add_554214;
  wire [7:0] sel_554215;
  wire [7:0] add_554218;
  wire [7:0] sel_554219;
  wire [7:0] add_554222;
  wire [7:0] sel_554223;
  wire [7:0] add_554226;
  wire [7:0] sel_554227;
  wire [7:0] add_554230;
  wire [7:0] sel_554231;
  wire [7:0] add_554234;
  wire [7:0] sel_554235;
  wire [7:0] add_554238;
  wire [7:0] sel_554239;
  wire [7:0] add_554242;
  wire [7:0] sel_554243;
  wire [7:0] add_554246;
  wire [7:0] sel_554247;
  wire [7:0] add_554250;
  wire [7:0] sel_554251;
  wire [7:0] add_554254;
  wire [7:0] sel_554255;
  wire [7:0] add_554258;
  wire [7:0] sel_554259;
  wire [7:0] add_554262;
  wire [7:0] sel_554263;
  wire [7:0] add_554266;
  wire [7:0] sel_554267;
  wire [7:0] add_554270;
  wire [7:0] sel_554271;
  wire [7:0] add_554274;
  wire [7:0] sel_554275;
  wire [7:0] add_554278;
  wire [7:0] sel_554279;
  wire [7:0] add_554282;
  wire [7:0] sel_554283;
  wire [7:0] add_554286;
  wire [7:0] sel_554287;
  wire [7:0] add_554290;
  wire [7:0] sel_554291;
  wire [7:0] add_554294;
  wire [7:0] sel_554295;
  wire [7:0] add_554298;
  wire [7:0] sel_554299;
  wire [7:0] add_554302;
  wire [7:0] sel_554303;
  wire [7:0] add_554306;
  wire [7:0] sel_554307;
  wire [7:0] add_554310;
  wire [7:0] sel_554311;
  wire [7:0] add_554314;
  wire [7:0] sel_554315;
  wire [7:0] add_554318;
  wire [7:0] sel_554319;
  wire [7:0] add_554322;
  wire [7:0] sel_554323;
  wire [7:0] add_554326;
  wire [7:0] sel_554327;
  wire [7:0] add_554330;
  wire [7:0] sel_554331;
  wire [7:0] add_554334;
  wire [7:0] sel_554335;
  wire [7:0] add_554338;
  wire [7:0] sel_554339;
  wire [7:0] add_554342;
  wire [7:0] sel_554343;
  wire [7:0] add_554346;
  wire [7:0] sel_554347;
  wire [7:0] add_554350;
  wire [7:0] sel_554351;
  wire [7:0] add_554354;
  wire [7:0] sel_554355;
  wire [7:0] add_554358;
  wire [7:0] sel_554359;
  wire [7:0] add_554362;
  wire [7:0] sel_554363;
  wire [7:0] add_554366;
  wire [7:0] sel_554367;
  wire [7:0] add_554370;
  wire [7:0] sel_554371;
  wire [7:0] add_554374;
  wire [7:0] sel_554375;
  wire [7:0] add_554378;
  wire [7:0] sel_554379;
  wire [7:0] add_554383;
  wire [15:0] array_index_554384;
  wire [7:0] sel_554385;
  wire [7:0] add_554388;
  wire [7:0] sel_554389;
  wire [7:0] add_554392;
  wire [7:0] sel_554393;
  wire [7:0] add_554396;
  wire [7:0] sel_554397;
  wire [7:0] add_554400;
  wire [7:0] sel_554401;
  wire [7:0] add_554404;
  wire [7:0] sel_554405;
  wire [7:0] add_554408;
  wire [7:0] sel_554409;
  wire [7:0] add_554412;
  wire [7:0] sel_554413;
  wire [7:0] add_554416;
  wire [7:0] sel_554417;
  wire [7:0] add_554420;
  wire [7:0] sel_554421;
  wire [7:0] add_554424;
  wire [7:0] sel_554425;
  wire [7:0] add_554428;
  wire [7:0] sel_554429;
  wire [7:0] add_554432;
  wire [7:0] sel_554433;
  wire [7:0] add_554436;
  wire [7:0] sel_554437;
  wire [7:0] add_554440;
  wire [7:0] sel_554441;
  wire [7:0] add_554444;
  wire [7:0] sel_554445;
  wire [7:0] add_554448;
  wire [7:0] sel_554449;
  wire [7:0] add_554452;
  wire [7:0] sel_554453;
  wire [7:0] add_554456;
  wire [7:0] sel_554457;
  wire [7:0] add_554460;
  wire [7:0] sel_554461;
  wire [7:0] add_554464;
  wire [7:0] sel_554465;
  wire [7:0] add_554468;
  wire [7:0] sel_554469;
  wire [7:0] add_554472;
  wire [7:0] sel_554473;
  wire [7:0] add_554476;
  wire [7:0] sel_554477;
  wire [7:0] add_554480;
  wire [7:0] sel_554481;
  wire [7:0] add_554484;
  wire [7:0] sel_554485;
  wire [7:0] add_554488;
  wire [7:0] sel_554489;
  wire [7:0] add_554492;
  wire [7:0] sel_554493;
  wire [7:0] add_554496;
  wire [7:0] sel_554497;
  wire [7:0] add_554500;
  wire [7:0] sel_554501;
  wire [7:0] add_554504;
  wire [7:0] sel_554505;
  wire [7:0] add_554508;
  wire [7:0] sel_554509;
  wire [7:0] add_554512;
  wire [7:0] sel_554513;
  wire [7:0] add_554516;
  wire [7:0] sel_554517;
  wire [7:0] add_554520;
  wire [7:0] sel_554521;
  wire [7:0] add_554524;
  wire [7:0] sel_554525;
  wire [7:0] add_554528;
  wire [7:0] sel_554529;
  wire [7:0] add_554532;
  wire [7:0] sel_554533;
  wire [7:0] add_554536;
  wire [7:0] sel_554537;
  wire [7:0] add_554540;
  wire [7:0] sel_554541;
  wire [7:0] add_554544;
  wire [7:0] sel_554545;
  wire [7:0] add_554548;
  wire [7:0] sel_554549;
  wire [7:0] add_554552;
  wire [7:0] sel_554553;
  wire [7:0] add_554556;
  wire [7:0] sel_554557;
  wire [7:0] add_554560;
  wire [7:0] sel_554561;
  wire [7:0] add_554564;
  wire [7:0] sel_554565;
  wire [7:0] add_554568;
  wire [7:0] sel_554569;
  wire [7:0] add_554572;
  wire [7:0] sel_554573;
  wire [7:0] add_554576;
  wire [7:0] sel_554577;
  wire [7:0] add_554580;
  wire [7:0] sel_554581;
  wire [7:0] add_554584;
  wire [7:0] sel_554585;
  wire [7:0] add_554588;
  wire [7:0] sel_554589;
  wire [7:0] add_554592;
  wire [7:0] sel_554593;
  wire [7:0] add_554596;
  wire [7:0] sel_554597;
  wire [7:0] add_554600;
  wire [7:0] sel_554601;
  wire [7:0] add_554604;
  wire [7:0] sel_554605;
  wire [7:0] add_554608;
  wire [7:0] sel_554609;
  wire [7:0] add_554612;
  wire [7:0] sel_554613;
  wire [7:0] add_554616;
  wire [7:0] sel_554617;
  wire [7:0] add_554620;
  wire [7:0] sel_554621;
  wire [7:0] add_554624;
  wire [7:0] sel_554625;
  wire [7:0] add_554628;
  wire [7:0] sel_554629;
  wire [7:0] add_554632;
  wire [7:0] sel_554633;
  wire [7:0] add_554636;
  wire [7:0] sel_554637;
  wire [7:0] add_554640;
  wire [7:0] sel_554641;
  wire [7:0] add_554644;
  wire [7:0] sel_554645;
  wire [7:0] add_554648;
  wire [7:0] sel_554649;
  wire [7:0] add_554652;
  wire [7:0] sel_554653;
  wire [7:0] add_554656;
  wire [7:0] sel_554657;
  wire [7:0] add_554660;
  wire [7:0] sel_554661;
  wire [7:0] add_554664;
  wire [7:0] sel_554665;
  wire [7:0] add_554668;
  wire [7:0] sel_554669;
  wire [7:0] add_554672;
  wire [7:0] sel_554673;
  wire [7:0] add_554676;
  wire [7:0] sel_554677;
  wire [7:0] add_554680;
  wire [7:0] sel_554681;
  wire [7:0] add_554685;
  wire [15:0] array_index_554686;
  wire [7:0] sel_554687;
  wire [7:0] add_554690;
  wire [7:0] sel_554691;
  wire [7:0] add_554694;
  wire [7:0] sel_554695;
  wire [7:0] add_554698;
  wire [7:0] sel_554699;
  wire [7:0] add_554702;
  wire [7:0] sel_554703;
  wire [7:0] add_554706;
  wire [7:0] sel_554707;
  wire [7:0] add_554710;
  wire [7:0] sel_554711;
  wire [7:0] add_554714;
  wire [7:0] sel_554715;
  wire [7:0] add_554718;
  wire [7:0] sel_554719;
  wire [7:0] add_554722;
  wire [7:0] sel_554723;
  wire [7:0] add_554726;
  wire [7:0] sel_554727;
  wire [7:0] add_554730;
  wire [7:0] sel_554731;
  wire [7:0] add_554734;
  wire [7:0] sel_554735;
  wire [7:0] add_554738;
  wire [7:0] sel_554739;
  wire [7:0] add_554742;
  wire [7:0] sel_554743;
  wire [7:0] add_554746;
  wire [7:0] sel_554747;
  wire [7:0] add_554750;
  wire [7:0] sel_554751;
  wire [7:0] add_554754;
  wire [7:0] sel_554755;
  wire [7:0] add_554758;
  wire [7:0] sel_554759;
  wire [7:0] add_554762;
  wire [7:0] sel_554763;
  wire [7:0] add_554766;
  wire [7:0] sel_554767;
  wire [7:0] add_554770;
  wire [7:0] sel_554771;
  wire [7:0] add_554774;
  wire [7:0] sel_554775;
  wire [7:0] add_554778;
  wire [7:0] sel_554779;
  wire [7:0] add_554782;
  wire [7:0] sel_554783;
  wire [7:0] add_554786;
  wire [7:0] sel_554787;
  wire [7:0] add_554790;
  wire [7:0] sel_554791;
  wire [7:0] add_554794;
  wire [7:0] sel_554795;
  wire [7:0] add_554798;
  wire [7:0] sel_554799;
  wire [7:0] add_554802;
  wire [7:0] sel_554803;
  wire [7:0] add_554806;
  wire [7:0] sel_554807;
  wire [7:0] add_554810;
  wire [7:0] sel_554811;
  wire [7:0] add_554814;
  wire [7:0] sel_554815;
  wire [7:0] add_554818;
  wire [7:0] sel_554819;
  wire [7:0] add_554822;
  wire [7:0] sel_554823;
  wire [7:0] add_554826;
  wire [7:0] sel_554827;
  wire [7:0] add_554830;
  wire [7:0] sel_554831;
  wire [7:0] add_554834;
  wire [7:0] sel_554835;
  wire [7:0] add_554838;
  wire [7:0] sel_554839;
  wire [7:0] add_554842;
  wire [7:0] sel_554843;
  wire [7:0] add_554846;
  wire [7:0] sel_554847;
  wire [7:0] add_554850;
  wire [7:0] sel_554851;
  wire [7:0] add_554854;
  wire [7:0] sel_554855;
  wire [7:0] add_554858;
  wire [7:0] sel_554859;
  wire [7:0] add_554862;
  wire [7:0] sel_554863;
  wire [7:0] add_554866;
  wire [7:0] sel_554867;
  wire [7:0] add_554870;
  wire [7:0] sel_554871;
  wire [7:0] add_554874;
  wire [7:0] sel_554875;
  wire [7:0] add_554878;
  wire [7:0] sel_554879;
  wire [7:0] add_554882;
  wire [7:0] sel_554883;
  wire [7:0] add_554886;
  wire [7:0] sel_554887;
  wire [7:0] add_554890;
  wire [7:0] sel_554891;
  wire [7:0] add_554894;
  wire [7:0] sel_554895;
  wire [7:0] add_554898;
  wire [7:0] sel_554899;
  wire [7:0] add_554902;
  wire [7:0] sel_554903;
  wire [7:0] add_554906;
  wire [7:0] sel_554907;
  wire [7:0] add_554910;
  wire [7:0] sel_554911;
  wire [7:0] add_554914;
  wire [7:0] sel_554915;
  wire [7:0] add_554918;
  wire [7:0] sel_554919;
  wire [7:0] add_554922;
  wire [7:0] sel_554923;
  wire [7:0] add_554926;
  wire [7:0] sel_554927;
  wire [7:0] add_554930;
  wire [7:0] sel_554931;
  wire [7:0] add_554934;
  wire [7:0] sel_554935;
  wire [7:0] add_554938;
  wire [7:0] sel_554939;
  wire [7:0] add_554942;
  wire [7:0] sel_554943;
  wire [7:0] add_554946;
  wire [7:0] sel_554947;
  wire [7:0] add_554950;
  wire [7:0] sel_554951;
  wire [7:0] add_554954;
  wire [7:0] sel_554955;
  wire [7:0] add_554958;
  wire [7:0] sel_554959;
  wire [7:0] add_554962;
  wire [7:0] sel_554963;
  wire [7:0] add_554966;
  wire [7:0] sel_554967;
  wire [7:0] add_554970;
  wire [7:0] sel_554971;
  wire [7:0] add_554974;
  wire [7:0] sel_554975;
  wire [7:0] add_554978;
  wire [7:0] sel_554979;
  wire [7:0] add_554982;
  wire [7:0] sel_554983;
  wire [7:0] add_554987;
  wire [15:0] array_index_554988;
  wire [7:0] sel_554989;
  wire [7:0] add_554992;
  wire [7:0] sel_554993;
  wire [7:0] add_554996;
  wire [7:0] sel_554997;
  wire [7:0] add_555000;
  wire [7:0] sel_555001;
  wire [7:0] add_555004;
  wire [7:0] sel_555005;
  wire [7:0] add_555008;
  wire [7:0] sel_555009;
  wire [7:0] add_555012;
  wire [7:0] sel_555013;
  wire [7:0] add_555016;
  wire [7:0] sel_555017;
  wire [7:0] add_555020;
  wire [7:0] sel_555021;
  wire [7:0] add_555024;
  wire [7:0] sel_555025;
  wire [7:0] add_555028;
  wire [7:0] sel_555029;
  wire [7:0] add_555032;
  wire [7:0] sel_555033;
  wire [7:0] add_555036;
  wire [7:0] sel_555037;
  wire [7:0] add_555040;
  wire [7:0] sel_555041;
  wire [7:0] add_555044;
  wire [7:0] sel_555045;
  wire [7:0] add_555048;
  wire [7:0] sel_555049;
  wire [7:0] add_555052;
  wire [7:0] sel_555053;
  wire [7:0] add_555056;
  wire [7:0] sel_555057;
  wire [7:0] add_555060;
  wire [7:0] sel_555061;
  wire [7:0] add_555064;
  wire [7:0] sel_555065;
  wire [7:0] add_555068;
  wire [7:0] sel_555069;
  wire [7:0] add_555072;
  wire [7:0] sel_555073;
  wire [7:0] add_555076;
  wire [7:0] sel_555077;
  wire [7:0] add_555080;
  wire [7:0] sel_555081;
  wire [7:0] add_555084;
  wire [7:0] sel_555085;
  wire [7:0] add_555088;
  wire [7:0] sel_555089;
  wire [7:0] add_555092;
  wire [7:0] sel_555093;
  wire [7:0] add_555096;
  wire [7:0] sel_555097;
  wire [7:0] add_555100;
  wire [7:0] sel_555101;
  wire [7:0] add_555104;
  wire [7:0] sel_555105;
  wire [7:0] add_555108;
  wire [7:0] sel_555109;
  wire [7:0] add_555112;
  wire [7:0] sel_555113;
  wire [7:0] add_555116;
  wire [7:0] sel_555117;
  wire [7:0] add_555120;
  wire [7:0] sel_555121;
  wire [7:0] add_555124;
  wire [7:0] sel_555125;
  wire [7:0] add_555128;
  wire [7:0] sel_555129;
  wire [7:0] add_555132;
  wire [7:0] sel_555133;
  wire [7:0] add_555136;
  wire [7:0] sel_555137;
  wire [7:0] add_555140;
  wire [7:0] sel_555141;
  wire [7:0] add_555144;
  wire [7:0] sel_555145;
  wire [7:0] add_555148;
  wire [7:0] sel_555149;
  wire [7:0] add_555152;
  wire [7:0] sel_555153;
  wire [7:0] add_555156;
  wire [7:0] sel_555157;
  wire [7:0] add_555160;
  wire [7:0] sel_555161;
  wire [7:0] add_555164;
  wire [7:0] sel_555165;
  wire [7:0] add_555168;
  wire [7:0] sel_555169;
  wire [7:0] add_555172;
  wire [7:0] sel_555173;
  wire [7:0] add_555176;
  wire [7:0] sel_555177;
  wire [7:0] add_555180;
  wire [7:0] sel_555181;
  wire [7:0] add_555184;
  wire [7:0] sel_555185;
  wire [7:0] add_555188;
  wire [7:0] sel_555189;
  wire [7:0] add_555192;
  wire [7:0] sel_555193;
  wire [7:0] add_555196;
  wire [7:0] sel_555197;
  wire [7:0] add_555200;
  wire [7:0] sel_555201;
  wire [7:0] add_555204;
  wire [7:0] sel_555205;
  wire [7:0] add_555208;
  wire [7:0] sel_555209;
  wire [7:0] add_555212;
  wire [7:0] sel_555213;
  wire [7:0] add_555216;
  wire [7:0] sel_555217;
  wire [7:0] add_555220;
  wire [7:0] sel_555221;
  wire [7:0] add_555224;
  wire [7:0] sel_555225;
  wire [7:0] add_555228;
  wire [7:0] sel_555229;
  wire [7:0] add_555232;
  wire [7:0] sel_555233;
  wire [7:0] add_555236;
  wire [7:0] sel_555237;
  wire [7:0] add_555240;
  wire [7:0] sel_555241;
  wire [7:0] add_555244;
  wire [7:0] sel_555245;
  wire [7:0] add_555248;
  wire [7:0] sel_555249;
  wire [7:0] add_555252;
  wire [7:0] sel_555253;
  wire [7:0] add_555256;
  wire [7:0] sel_555257;
  wire [7:0] add_555260;
  wire [7:0] sel_555261;
  wire [7:0] add_555264;
  wire [7:0] sel_555265;
  wire [7:0] add_555268;
  wire [7:0] sel_555269;
  wire [7:0] add_555272;
  wire [7:0] sel_555273;
  wire [7:0] add_555276;
  wire [7:0] sel_555277;
  wire [7:0] add_555280;
  wire [7:0] sel_555281;
  wire [7:0] add_555284;
  wire [7:0] sel_555285;
  wire [7:0] add_555289;
  wire [15:0] array_index_555290;
  wire [7:0] sel_555291;
  wire [7:0] add_555294;
  wire [7:0] sel_555295;
  wire [7:0] add_555298;
  wire [7:0] sel_555299;
  wire [7:0] add_555302;
  wire [7:0] sel_555303;
  wire [7:0] add_555306;
  wire [7:0] sel_555307;
  wire [7:0] add_555310;
  wire [7:0] sel_555311;
  wire [7:0] add_555314;
  wire [7:0] sel_555315;
  wire [7:0] add_555318;
  wire [7:0] sel_555319;
  wire [7:0] add_555322;
  wire [7:0] sel_555323;
  wire [7:0] add_555326;
  wire [7:0] sel_555327;
  wire [7:0] add_555330;
  wire [7:0] sel_555331;
  wire [7:0] add_555334;
  wire [7:0] sel_555335;
  wire [7:0] add_555338;
  wire [7:0] sel_555339;
  wire [7:0] add_555342;
  wire [7:0] sel_555343;
  wire [7:0] add_555346;
  wire [7:0] sel_555347;
  wire [7:0] add_555350;
  wire [7:0] sel_555351;
  wire [7:0] add_555354;
  wire [7:0] sel_555355;
  wire [7:0] add_555358;
  wire [7:0] sel_555359;
  wire [7:0] add_555362;
  wire [7:0] sel_555363;
  wire [7:0] add_555366;
  wire [7:0] sel_555367;
  wire [7:0] add_555370;
  wire [7:0] sel_555371;
  wire [7:0] add_555374;
  wire [7:0] sel_555375;
  wire [7:0] add_555378;
  wire [7:0] sel_555379;
  wire [7:0] add_555382;
  wire [7:0] sel_555383;
  wire [7:0] add_555386;
  wire [7:0] sel_555387;
  wire [7:0] add_555390;
  wire [7:0] sel_555391;
  wire [7:0] add_555394;
  wire [7:0] sel_555395;
  wire [7:0] add_555398;
  wire [7:0] sel_555399;
  wire [7:0] add_555402;
  wire [7:0] sel_555403;
  wire [7:0] add_555406;
  wire [7:0] sel_555407;
  wire [7:0] add_555410;
  wire [7:0] sel_555411;
  wire [7:0] add_555414;
  wire [7:0] sel_555415;
  wire [7:0] add_555418;
  wire [7:0] sel_555419;
  wire [7:0] add_555422;
  wire [7:0] sel_555423;
  wire [7:0] add_555426;
  wire [7:0] sel_555427;
  wire [7:0] add_555430;
  wire [7:0] sel_555431;
  wire [7:0] add_555434;
  wire [7:0] sel_555435;
  wire [7:0] add_555438;
  wire [7:0] sel_555439;
  wire [7:0] add_555442;
  wire [7:0] sel_555443;
  wire [7:0] add_555446;
  wire [7:0] sel_555447;
  wire [7:0] add_555450;
  wire [7:0] sel_555451;
  wire [7:0] add_555454;
  wire [7:0] sel_555455;
  wire [7:0] add_555458;
  wire [7:0] sel_555459;
  wire [7:0] add_555462;
  wire [7:0] sel_555463;
  wire [7:0] add_555466;
  wire [7:0] sel_555467;
  wire [7:0] add_555470;
  wire [7:0] sel_555471;
  wire [7:0] add_555474;
  wire [7:0] sel_555475;
  wire [7:0] add_555478;
  wire [7:0] sel_555479;
  wire [7:0] add_555482;
  wire [7:0] sel_555483;
  wire [7:0] add_555486;
  wire [7:0] sel_555487;
  wire [7:0] add_555490;
  wire [7:0] sel_555491;
  wire [7:0] add_555494;
  wire [7:0] sel_555495;
  wire [7:0] add_555498;
  wire [7:0] sel_555499;
  wire [7:0] add_555502;
  wire [7:0] sel_555503;
  wire [7:0] add_555506;
  wire [7:0] sel_555507;
  wire [7:0] add_555510;
  wire [7:0] sel_555511;
  wire [7:0] add_555514;
  wire [7:0] sel_555515;
  wire [7:0] add_555518;
  wire [7:0] sel_555519;
  wire [7:0] add_555522;
  wire [7:0] sel_555523;
  wire [7:0] add_555526;
  wire [7:0] sel_555527;
  wire [7:0] add_555530;
  wire [7:0] sel_555531;
  wire [7:0] add_555534;
  wire [7:0] sel_555535;
  wire [7:0] add_555538;
  wire [7:0] sel_555539;
  wire [7:0] add_555542;
  wire [7:0] sel_555543;
  wire [7:0] add_555546;
  wire [7:0] sel_555547;
  wire [7:0] add_555550;
  wire [7:0] sel_555551;
  wire [7:0] add_555554;
  wire [7:0] sel_555555;
  wire [7:0] add_555558;
  wire [7:0] sel_555559;
  wire [7:0] add_555562;
  wire [7:0] sel_555563;
  wire [7:0] add_555566;
  wire [7:0] sel_555567;
  wire [7:0] add_555570;
  wire [7:0] sel_555571;
  wire [7:0] add_555574;
  wire [7:0] sel_555575;
  wire [7:0] add_555578;
  wire [7:0] sel_555579;
  wire [7:0] add_555582;
  wire [7:0] sel_555583;
  wire [7:0] add_555586;
  wire [7:0] sel_555587;
  wire [7:0] add_555591;
  wire [15:0] array_index_555592;
  wire [7:0] sel_555593;
  wire [7:0] add_555596;
  wire [7:0] sel_555597;
  wire [7:0] add_555600;
  wire [7:0] sel_555601;
  wire [7:0] add_555604;
  wire [7:0] sel_555605;
  wire [7:0] add_555608;
  wire [7:0] sel_555609;
  wire [7:0] add_555612;
  wire [7:0] sel_555613;
  wire [7:0] add_555616;
  wire [7:0] sel_555617;
  wire [7:0] add_555620;
  wire [7:0] sel_555621;
  wire [7:0] add_555624;
  wire [7:0] sel_555625;
  wire [7:0] add_555628;
  wire [7:0] sel_555629;
  wire [7:0] add_555632;
  wire [7:0] sel_555633;
  wire [7:0] add_555636;
  wire [7:0] sel_555637;
  wire [7:0] add_555640;
  wire [7:0] sel_555641;
  wire [7:0] add_555644;
  wire [7:0] sel_555645;
  wire [7:0] add_555648;
  wire [7:0] sel_555649;
  wire [7:0] add_555652;
  wire [7:0] sel_555653;
  wire [7:0] add_555656;
  wire [7:0] sel_555657;
  wire [7:0] add_555660;
  wire [7:0] sel_555661;
  wire [7:0] add_555664;
  wire [7:0] sel_555665;
  wire [7:0] add_555668;
  wire [7:0] sel_555669;
  wire [7:0] add_555672;
  wire [7:0] sel_555673;
  wire [7:0] add_555676;
  wire [7:0] sel_555677;
  wire [7:0] add_555680;
  wire [7:0] sel_555681;
  wire [7:0] add_555684;
  wire [7:0] sel_555685;
  wire [7:0] add_555688;
  wire [7:0] sel_555689;
  wire [7:0] add_555692;
  wire [7:0] sel_555693;
  wire [7:0] add_555696;
  wire [7:0] sel_555697;
  wire [7:0] add_555700;
  wire [7:0] sel_555701;
  wire [7:0] add_555704;
  wire [7:0] sel_555705;
  wire [7:0] add_555708;
  wire [7:0] sel_555709;
  wire [7:0] add_555712;
  wire [7:0] sel_555713;
  wire [7:0] add_555716;
  wire [7:0] sel_555717;
  wire [7:0] add_555720;
  wire [7:0] sel_555721;
  wire [7:0] add_555724;
  wire [7:0] sel_555725;
  wire [7:0] add_555728;
  wire [7:0] sel_555729;
  wire [7:0] add_555732;
  wire [7:0] sel_555733;
  wire [7:0] add_555736;
  wire [7:0] sel_555737;
  wire [7:0] add_555740;
  wire [7:0] sel_555741;
  wire [7:0] add_555744;
  wire [7:0] sel_555745;
  wire [7:0] add_555748;
  wire [7:0] sel_555749;
  wire [7:0] add_555752;
  wire [7:0] sel_555753;
  wire [7:0] add_555756;
  wire [7:0] sel_555757;
  wire [7:0] add_555760;
  wire [7:0] sel_555761;
  wire [7:0] add_555764;
  wire [7:0] sel_555765;
  wire [7:0] add_555768;
  wire [7:0] sel_555769;
  wire [7:0] add_555772;
  wire [7:0] sel_555773;
  wire [7:0] add_555776;
  wire [7:0] sel_555777;
  wire [7:0] add_555780;
  wire [7:0] sel_555781;
  wire [7:0] add_555784;
  wire [7:0] sel_555785;
  wire [7:0] add_555788;
  wire [7:0] sel_555789;
  wire [7:0] add_555792;
  wire [7:0] sel_555793;
  wire [7:0] add_555796;
  wire [7:0] sel_555797;
  wire [7:0] add_555800;
  wire [7:0] sel_555801;
  wire [7:0] add_555804;
  wire [7:0] sel_555805;
  wire [7:0] add_555808;
  wire [7:0] sel_555809;
  wire [7:0] add_555812;
  wire [7:0] sel_555813;
  wire [7:0] add_555816;
  wire [7:0] sel_555817;
  wire [7:0] add_555820;
  wire [7:0] sel_555821;
  wire [7:0] add_555824;
  wire [7:0] sel_555825;
  wire [7:0] add_555828;
  wire [7:0] sel_555829;
  wire [7:0] add_555832;
  wire [7:0] sel_555833;
  wire [7:0] add_555836;
  wire [7:0] sel_555837;
  wire [7:0] add_555840;
  wire [7:0] sel_555841;
  wire [7:0] add_555844;
  wire [7:0] sel_555845;
  wire [7:0] add_555848;
  wire [7:0] sel_555849;
  wire [7:0] add_555852;
  wire [7:0] sel_555853;
  wire [7:0] add_555856;
  wire [7:0] sel_555857;
  wire [7:0] add_555860;
  wire [7:0] sel_555861;
  wire [7:0] add_555864;
  wire [7:0] sel_555865;
  wire [7:0] add_555868;
  wire [7:0] sel_555869;
  wire [7:0] add_555872;
  wire [7:0] sel_555873;
  wire [7:0] add_555876;
  wire [7:0] sel_555877;
  wire [7:0] add_555880;
  wire [7:0] sel_555881;
  wire [7:0] add_555884;
  wire [7:0] sel_555885;
  wire [7:0] add_555888;
  wire [7:0] sel_555889;
  wire [7:0] add_555893;
  wire [15:0] array_index_555894;
  wire [7:0] sel_555895;
  wire [7:0] add_555898;
  wire [7:0] sel_555899;
  wire [7:0] add_555902;
  wire [7:0] sel_555903;
  wire [7:0] add_555906;
  wire [7:0] sel_555907;
  wire [7:0] add_555910;
  wire [7:0] sel_555911;
  wire [7:0] add_555914;
  wire [7:0] sel_555915;
  wire [7:0] add_555918;
  wire [7:0] sel_555919;
  wire [7:0] add_555922;
  wire [7:0] sel_555923;
  wire [7:0] add_555926;
  wire [7:0] sel_555927;
  wire [7:0] add_555930;
  wire [7:0] sel_555931;
  wire [7:0] add_555934;
  wire [7:0] sel_555935;
  wire [7:0] add_555938;
  wire [7:0] sel_555939;
  wire [7:0] add_555942;
  wire [7:0] sel_555943;
  wire [7:0] add_555946;
  wire [7:0] sel_555947;
  wire [7:0] add_555950;
  wire [7:0] sel_555951;
  wire [7:0] add_555954;
  wire [7:0] sel_555955;
  wire [7:0] add_555958;
  wire [7:0] sel_555959;
  wire [7:0] add_555962;
  wire [7:0] sel_555963;
  wire [7:0] add_555966;
  wire [7:0] sel_555967;
  wire [7:0] add_555970;
  wire [7:0] sel_555971;
  wire [7:0] add_555974;
  wire [7:0] sel_555975;
  wire [7:0] add_555978;
  wire [7:0] sel_555979;
  wire [7:0] add_555982;
  wire [7:0] sel_555983;
  wire [7:0] add_555986;
  wire [7:0] sel_555987;
  wire [7:0] add_555990;
  wire [7:0] sel_555991;
  wire [7:0] add_555994;
  wire [7:0] sel_555995;
  wire [7:0] add_555998;
  wire [7:0] sel_555999;
  wire [7:0] add_556002;
  wire [7:0] sel_556003;
  wire [7:0] add_556006;
  wire [7:0] sel_556007;
  wire [7:0] add_556010;
  wire [7:0] sel_556011;
  wire [7:0] add_556014;
  wire [7:0] sel_556015;
  wire [7:0] add_556018;
  wire [7:0] sel_556019;
  wire [7:0] add_556022;
  wire [7:0] sel_556023;
  wire [7:0] add_556026;
  wire [7:0] sel_556027;
  wire [7:0] add_556030;
  wire [7:0] sel_556031;
  wire [7:0] add_556034;
  wire [7:0] sel_556035;
  wire [7:0] add_556038;
  wire [7:0] sel_556039;
  wire [7:0] add_556042;
  wire [7:0] sel_556043;
  wire [7:0] add_556046;
  wire [7:0] sel_556047;
  wire [7:0] add_556050;
  wire [7:0] sel_556051;
  wire [7:0] add_556054;
  wire [7:0] sel_556055;
  wire [7:0] add_556058;
  wire [7:0] sel_556059;
  wire [7:0] add_556062;
  wire [7:0] sel_556063;
  wire [7:0] add_556066;
  wire [7:0] sel_556067;
  wire [7:0] add_556070;
  wire [7:0] sel_556071;
  wire [7:0] add_556074;
  wire [7:0] sel_556075;
  wire [7:0] add_556078;
  wire [7:0] sel_556079;
  wire [7:0] add_556082;
  wire [7:0] sel_556083;
  wire [7:0] add_556086;
  wire [7:0] sel_556087;
  wire [7:0] add_556090;
  wire [7:0] sel_556091;
  wire [7:0] add_556094;
  wire [7:0] sel_556095;
  wire [7:0] add_556098;
  wire [7:0] sel_556099;
  wire [7:0] add_556102;
  wire [7:0] sel_556103;
  wire [7:0] add_556106;
  wire [7:0] sel_556107;
  wire [7:0] add_556110;
  wire [7:0] sel_556111;
  wire [7:0] add_556114;
  wire [7:0] sel_556115;
  wire [7:0] add_556118;
  wire [7:0] sel_556119;
  wire [7:0] add_556122;
  wire [7:0] sel_556123;
  wire [7:0] add_556126;
  wire [7:0] sel_556127;
  wire [7:0] add_556130;
  wire [7:0] sel_556131;
  wire [7:0] add_556134;
  wire [7:0] sel_556135;
  wire [7:0] add_556138;
  wire [7:0] sel_556139;
  wire [7:0] add_556142;
  wire [7:0] sel_556143;
  wire [7:0] add_556146;
  wire [7:0] sel_556147;
  wire [7:0] add_556150;
  wire [7:0] sel_556151;
  wire [7:0] add_556154;
  wire [7:0] sel_556155;
  wire [7:0] add_556158;
  wire [7:0] sel_556159;
  wire [7:0] add_556162;
  wire [7:0] sel_556163;
  wire [7:0] add_556166;
  wire [7:0] sel_556167;
  wire [7:0] add_556170;
  wire [7:0] sel_556171;
  wire [7:0] add_556174;
  wire [7:0] sel_556175;
  wire [7:0] add_556178;
  wire [7:0] sel_556179;
  wire [7:0] add_556182;
  wire [7:0] sel_556183;
  wire [7:0] add_556186;
  wire [7:0] sel_556187;
  wire [7:0] add_556190;
  wire [7:0] sel_556191;
  wire [7:0] add_556195;
  wire [15:0] array_index_556196;
  wire [7:0] sel_556197;
  wire [7:0] add_556200;
  wire [7:0] sel_556201;
  wire [7:0] add_556204;
  wire [7:0] sel_556205;
  wire [7:0] add_556208;
  wire [7:0] sel_556209;
  wire [7:0] add_556212;
  wire [7:0] sel_556213;
  wire [7:0] add_556216;
  wire [7:0] sel_556217;
  wire [7:0] add_556220;
  wire [7:0] sel_556221;
  wire [7:0] add_556224;
  wire [7:0] sel_556225;
  wire [7:0] add_556228;
  wire [7:0] sel_556229;
  wire [7:0] add_556232;
  wire [7:0] sel_556233;
  wire [7:0] add_556236;
  wire [7:0] sel_556237;
  wire [7:0] add_556240;
  wire [7:0] sel_556241;
  wire [7:0] add_556244;
  wire [7:0] sel_556245;
  wire [7:0] add_556248;
  wire [7:0] sel_556249;
  wire [7:0] add_556252;
  wire [7:0] sel_556253;
  wire [7:0] add_556256;
  wire [7:0] sel_556257;
  wire [7:0] add_556260;
  wire [7:0] sel_556261;
  wire [7:0] add_556264;
  wire [7:0] sel_556265;
  wire [7:0] add_556268;
  wire [7:0] sel_556269;
  wire [7:0] add_556272;
  wire [7:0] sel_556273;
  wire [7:0] add_556276;
  wire [7:0] sel_556277;
  wire [7:0] add_556280;
  wire [7:0] sel_556281;
  wire [7:0] add_556284;
  wire [7:0] sel_556285;
  wire [7:0] add_556288;
  wire [7:0] sel_556289;
  wire [7:0] add_556292;
  wire [7:0] sel_556293;
  wire [7:0] add_556296;
  wire [7:0] sel_556297;
  wire [7:0] add_556300;
  wire [7:0] sel_556301;
  wire [7:0] add_556304;
  wire [7:0] sel_556305;
  wire [7:0] add_556308;
  wire [7:0] sel_556309;
  wire [7:0] add_556312;
  wire [7:0] sel_556313;
  wire [7:0] add_556316;
  wire [7:0] sel_556317;
  wire [7:0] add_556320;
  wire [7:0] sel_556321;
  wire [7:0] add_556324;
  wire [7:0] sel_556325;
  wire [7:0] add_556328;
  wire [7:0] sel_556329;
  wire [7:0] add_556332;
  wire [7:0] sel_556333;
  wire [7:0] add_556336;
  wire [7:0] sel_556337;
  wire [7:0] add_556340;
  wire [7:0] sel_556341;
  wire [7:0] add_556344;
  wire [7:0] sel_556345;
  wire [7:0] add_556348;
  wire [7:0] sel_556349;
  wire [7:0] add_556352;
  wire [7:0] sel_556353;
  wire [7:0] add_556356;
  wire [7:0] sel_556357;
  wire [7:0] add_556360;
  wire [7:0] sel_556361;
  wire [7:0] add_556364;
  wire [7:0] sel_556365;
  wire [7:0] add_556368;
  wire [7:0] sel_556369;
  wire [7:0] add_556372;
  wire [7:0] sel_556373;
  wire [7:0] add_556376;
  wire [7:0] sel_556377;
  wire [7:0] add_556380;
  wire [7:0] sel_556381;
  wire [7:0] add_556384;
  wire [7:0] sel_556385;
  wire [7:0] add_556388;
  wire [7:0] sel_556389;
  wire [7:0] add_556392;
  wire [7:0] sel_556393;
  wire [7:0] add_556396;
  wire [7:0] sel_556397;
  wire [7:0] add_556400;
  wire [7:0] sel_556401;
  wire [7:0] add_556404;
  wire [7:0] sel_556405;
  wire [7:0] add_556408;
  wire [7:0] sel_556409;
  wire [7:0] add_556412;
  wire [7:0] sel_556413;
  wire [7:0] add_556416;
  wire [7:0] sel_556417;
  wire [7:0] add_556420;
  wire [7:0] sel_556421;
  wire [7:0] add_556424;
  wire [7:0] sel_556425;
  wire [7:0] add_556428;
  wire [7:0] sel_556429;
  wire [7:0] add_556432;
  wire [7:0] sel_556433;
  wire [7:0] add_556436;
  wire [7:0] sel_556437;
  wire [7:0] add_556440;
  wire [7:0] sel_556441;
  wire [7:0] add_556444;
  wire [7:0] sel_556445;
  wire [7:0] add_556448;
  wire [7:0] sel_556449;
  wire [7:0] add_556452;
  wire [7:0] sel_556453;
  wire [7:0] add_556456;
  wire [7:0] sel_556457;
  wire [7:0] add_556460;
  wire [7:0] sel_556461;
  wire [7:0] add_556464;
  wire [7:0] sel_556465;
  wire [7:0] add_556468;
  wire [7:0] sel_556469;
  wire [7:0] add_556472;
  wire [7:0] sel_556473;
  wire [7:0] add_556476;
  wire [7:0] sel_556477;
  wire [7:0] add_556480;
  wire [7:0] sel_556481;
  wire [7:0] add_556484;
  wire [7:0] sel_556485;
  wire [7:0] add_556488;
  wire [7:0] sel_556489;
  wire [7:0] add_556492;
  wire [7:0] sel_556493;
  wire [7:0] add_556497;
  wire [15:0] array_index_556498;
  wire [7:0] sel_556499;
  wire [7:0] add_556502;
  wire [7:0] sel_556503;
  wire [7:0] add_556506;
  wire [7:0] sel_556507;
  wire [7:0] add_556510;
  wire [7:0] sel_556511;
  wire [7:0] add_556514;
  wire [7:0] sel_556515;
  wire [7:0] add_556518;
  wire [7:0] sel_556519;
  wire [7:0] add_556522;
  wire [7:0] sel_556523;
  wire [7:0] add_556526;
  wire [7:0] sel_556527;
  wire [7:0] add_556530;
  wire [7:0] sel_556531;
  wire [7:0] add_556534;
  wire [7:0] sel_556535;
  wire [7:0] add_556538;
  wire [7:0] sel_556539;
  wire [7:0] add_556542;
  wire [7:0] sel_556543;
  wire [7:0] add_556546;
  wire [7:0] sel_556547;
  wire [7:0] add_556550;
  wire [7:0] sel_556551;
  wire [7:0] add_556554;
  wire [7:0] sel_556555;
  wire [7:0] add_556558;
  wire [7:0] sel_556559;
  wire [7:0] add_556562;
  wire [7:0] sel_556563;
  wire [7:0] add_556566;
  wire [7:0] sel_556567;
  wire [7:0] add_556570;
  wire [7:0] sel_556571;
  wire [7:0] add_556574;
  wire [7:0] sel_556575;
  wire [7:0] add_556578;
  wire [7:0] sel_556579;
  wire [7:0] add_556582;
  wire [7:0] sel_556583;
  wire [7:0] add_556586;
  wire [7:0] sel_556587;
  wire [7:0] add_556590;
  wire [7:0] sel_556591;
  wire [7:0] add_556594;
  wire [7:0] sel_556595;
  wire [7:0] add_556598;
  wire [7:0] sel_556599;
  wire [7:0] add_556602;
  wire [7:0] sel_556603;
  wire [7:0] add_556606;
  wire [7:0] sel_556607;
  wire [7:0] add_556610;
  wire [7:0] sel_556611;
  wire [7:0] add_556614;
  wire [7:0] sel_556615;
  wire [7:0] add_556618;
  wire [7:0] sel_556619;
  wire [7:0] add_556622;
  wire [7:0] sel_556623;
  wire [7:0] add_556626;
  wire [7:0] sel_556627;
  wire [7:0] add_556630;
  wire [7:0] sel_556631;
  wire [7:0] add_556634;
  wire [7:0] sel_556635;
  wire [7:0] add_556638;
  wire [7:0] sel_556639;
  wire [7:0] add_556642;
  wire [7:0] sel_556643;
  wire [7:0] add_556646;
  wire [7:0] sel_556647;
  wire [7:0] add_556650;
  wire [7:0] sel_556651;
  wire [7:0] add_556654;
  wire [7:0] sel_556655;
  wire [7:0] add_556658;
  wire [7:0] sel_556659;
  wire [7:0] add_556662;
  wire [7:0] sel_556663;
  wire [7:0] add_556666;
  wire [7:0] sel_556667;
  wire [7:0] add_556670;
  wire [7:0] sel_556671;
  wire [7:0] add_556674;
  wire [7:0] sel_556675;
  wire [7:0] add_556678;
  wire [7:0] sel_556679;
  wire [7:0] add_556682;
  wire [7:0] sel_556683;
  wire [7:0] add_556686;
  wire [7:0] sel_556687;
  wire [7:0] add_556690;
  wire [7:0] sel_556691;
  wire [7:0] add_556694;
  wire [7:0] sel_556695;
  wire [7:0] add_556698;
  wire [7:0] sel_556699;
  wire [7:0] add_556702;
  wire [7:0] sel_556703;
  wire [7:0] add_556706;
  wire [7:0] sel_556707;
  wire [7:0] add_556710;
  wire [7:0] sel_556711;
  wire [7:0] add_556714;
  wire [7:0] sel_556715;
  wire [7:0] add_556718;
  wire [7:0] sel_556719;
  wire [7:0] add_556722;
  wire [7:0] sel_556723;
  wire [7:0] add_556726;
  wire [7:0] sel_556727;
  wire [7:0] add_556730;
  wire [7:0] sel_556731;
  wire [7:0] add_556734;
  wire [7:0] sel_556735;
  wire [7:0] add_556738;
  wire [7:0] sel_556739;
  wire [7:0] add_556742;
  wire [7:0] sel_556743;
  wire [7:0] add_556746;
  wire [7:0] sel_556747;
  wire [7:0] add_556750;
  wire [7:0] sel_556751;
  wire [7:0] add_556754;
  wire [7:0] sel_556755;
  wire [7:0] add_556758;
  wire [7:0] sel_556759;
  wire [7:0] add_556762;
  wire [7:0] sel_556763;
  wire [7:0] add_556766;
  wire [7:0] sel_556767;
  wire [7:0] add_556770;
  wire [7:0] sel_556771;
  wire [7:0] add_556774;
  wire [7:0] sel_556775;
  wire [7:0] add_556778;
  wire [7:0] sel_556779;
  wire [7:0] add_556782;
  wire [7:0] sel_556783;
  wire [7:0] add_556786;
  wire [7:0] sel_556787;
  wire [7:0] add_556790;
  wire [7:0] sel_556791;
  wire [7:0] add_556794;
  wire [7:0] sel_556795;
  wire [7:0] add_556799;
  wire [15:0] array_index_556800;
  wire [7:0] sel_556801;
  wire [7:0] add_556804;
  wire [7:0] sel_556805;
  wire [7:0] add_556808;
  wire [7:0] sel_556809;
  wire [7:0] add_556812;
  wire [7:0] sel_556813;
  wire [7:0] add_556816;
  wire [7:0] sel_556817;
  wire [7:0] add_556820;
  wire [7:0] sel_556821;
  wire [7:0] add_556824;
  wire [7:0] sel_556825;
  wire [7:0] add_556828;
  wire [7:0] sel_556829;
  wire [7:0] add_556832;
  wire [7:0] sel_556833;
  wire [7:0] add_556836;
  wire [7:0] sel_556837;
  wire [7:0] add_556840;
  wire [7:0] sel_556841;
  wire [7:0] add_556844;
  wire [7:0] sel_556845;
  wire [7:0] add_556848;
  wire [7:0] sel_556849;
  wire [7:0] add_556852;
  wire [7:0] sel_556853;
  wire [7:0] add_556856;
  wire [7:0] sel_556857;
  wire [7:0] add_556860;
  wire [7:0] sel_556861;
  wire [7:0] add_556864;
  wire [7:0] sel_556865;
  wire [7:0] add_556868;
  wire [7:0] sel_556869;
  wire [7:0] add_556872;
  wire [7:0] sel_556873;
  wire [7:0] add_556876;
  wire [7:0] sel_556877;
  wire [7:0] add_556880;
  wire [7:0] sel_556881;
  wire [7:0] add_556884;
  wire [7:0] sel_556885;
  wire [7:0] add_556888;
  wire [7:0] sel_556889;
  wire [7:0] add_556892;
  wire [7:0] sel_556893;
  wire [7:0] add_556896;
  wire [7:0] sel_556897;
  wire [7:0] add_556900;
  wire [7:0] sel_556901;
  wire [7:0] add_556904;
  wire [7:0] sel_556905;
  wire [7:0] add_556908;
  wire [7:0] sel_556909;
  wire [7:0] add_556912;
  wire [7:0] sel_556913;
  wire [7:0] add_556916;
  wire [7:0] sel_556917;
  wire [7:0] add_556920;
  wire [7:0] sel_556921;
  wire [7:0] add_556924;
  wire [7:0] sel_556925;
  wire [7:0] add_556928;
  wire [7:0] sel_556929;
  wire [7:0] add_556932;
  wire [7:0] sel_556933;
  wire [7:0] add_556936;
  wire [7:0] sel_556937;
  wire [7:0] add_556940;
  wire [7:0] sel_556941;
  wire [7:0] add_556944;
  wire [7:0] sel_556945;
  wire [7:0] add_556948;
  wire [7:0] sel_556949;
  wire [7:0] add_556952;
  wire [7:0] sel_556953;
  wire [7:0] add_556956;
  wire [7:0] sel_556957;
  wire [7:0] add_556960;
  wire [7:0] sel_556961;
  wire [7:0] add_556964;
  wire [7:0] sel_556965;
  wire [7:0] add_556968;
  wire [7:0] sel_556969;
  wire [7:0] add_556972;
  wire [7:0] sel_556973;
  wire [7:0] add_556976;
  wire [7:0] sel_556977;
  wire [7:0] add_556980;
  wire [7:0] sel_556981;
  wire [7:0] add_556984;
  wire [7:0] sel_556985;
  wire [7:0] add_556988;
  wire [7:0] sel_556989;
  wire [7:0] add_556992;
  wire [7:0] sel_556993;
  wire [7:0] add_556996;
  wire [7:0] sel_556997;
  wire [7:0] add_557000;
  wire [7:0] sel_557001;
  wire [7:0] add_557004;
  wire [7:0] sel_557005;
  wire [7:0] add_557008;
  wire [7:0] sel_557009;
  wire [7:0] add_557012;
  wire [7:0] sel_557013;
  wire [7:0] add_557016;
  wire [7:0] sel_557017;
  wire [7:0] add_557020;
  wire [7:0] sel_557021;
  wire [7:0] add_557024;
  wire [7:0] sel_557025;
  wire [7:0] add_557028;
  wire [7:0] sel_557029;
  wire [7:0] add_557032;
  wire [7:0] sel_557033;
  wire [7:0] add_557036;
  wire [7:0] sel_557037;
  wire [7:0] add_557040;
  wire [7:0] sel_557041;
  wire [7:0] add_557044;
  wire [7:0] sel_557045;
  wire [7:0] add_557048;
  wire [7:0] sel_557049;
  wire [7:0] add_557052;
  wire [7:0] sel_557053;
  wire [7:0] add_557056;
  wire [7:0] sel_557057;
  wire [7:0] add_557060;
  wire [7:0] sel_557061;
  wire [7:0] add_557064;
  wire [7:0] sel_557065;
  wire [7:0] add_557068;
  wire [7:0] sel_557069;
  wire [7:0] add_557072;
  wire [7:0] sel_557073;
  wire [7:0] add_557076;
  wire [7:0] sel_557077;
  wire [7:0] add_557080;
  wire [7:0] sel_557081;
  wire [7:0] add_557084;
  wire [7:0] sel_557085;
  wire [7:0] add_557088;
  wire [7:0] sel_557089;
  wire [7:0] add_557092;
  wire [7:0] sel_557093;
  wire [7:0] add_557096;
  wire [7:0] sel_557097;
  wire [7:0] add_557101;
  wire [15:0] array_index_557102;
  wire [7:0] sel_557103;
  wire [7:0] add_557106;
  wire [7:0] sel_557107;
  wire [7:0] add_557110;
  wire [7:0] sel_557111;
  wire [7:0] add_557114;
  wire [7:0] sel_557115;
  wire [7:0] add_557118;
  wire [7:0] sel_557119;
  wire [7:0] add_557122;
  wire [7:0] sel_557123;
  wire [7:0] add_557126;
  wire [7:0] sel_557127;
  wire [7:0] add_557130;
  wire [7:0] sel_557131;
  wire [7:0] add_557134;
  wire [7:0] sel_557135;
  wire [7:0] add_557138;
  wire [7:0] sel_557139;
  wire [7:0] add_557142;
  wire [7:0] sel_557143;
  wire [7:0] add_557146;
  wire [7:0] sel_557147;
  wire [7:0] add_557150;
  wire [7:0] sel_557151;
  wire [7:0] add_557154;
  wire [7:0] sel_557155;
  wire [7:0] add_557158;
  wire [7:0] sel_557159;
  wire [7:0] add_557162;
  wire [7:0] sel_557163;
  wire [7:0] add_557166;
  wire [7:0] sel_557167;
  wire [7:0] add_557170;
  wire [7:0] sel_557171;
  wire [7:0] add_557174;
  wire [7:0] sel_557175;
  wire [7:0] add_557178;
  wire [7:0] sel_557179;
  wire [7:0] add_557182;
  wire [7:0] sel_557183;
  wire [7:0] add_557186;
  wire [7:0] sel_557187;
  wire [7:0] add_557190;
  wire [7:0] sel_557191;
  wire [7:0] add_557194;
  wire [7:0] sel_557195;
  wire [7:0] add_557198;
  wire [7:0] sel_557199;
  wire [7:0] add_557202;
  wire [7:0] sel_557203;
  wire [7:0] add_557206;
  wire [7:0] sel_557207;
  wire [7:0] add_557210;
  wire [7:0] sel_557211;
  wire [7:0] add_557214;
  wire [7:0] sel_557215;
  wire [7:0] add_557218;
  wire [7:0] sel_557219;
  wire [7:0] add_557222;
  wire [7:0] sel_557223;
  wire [7:0] add_557226;
  wire [7:0] sel_557227;
  wire [7:0] add_557230;
  wire [7:0] sel_557231;
  wire [7:0] add_557234;
  wire [7:0] sel_557235;
  wire [7:0] add_557238;
  wire [7:0] sel_557239;
  wire [7:0] add_557242;
  wire [7:0] sel_557243;
  wire [7:0] add_557246;
  wire [7:0] sel_557247;
  wire [7:0] add_557250;
  wire [7:0] sel_557251;
  wire [7:0] add_557254;
  wire [7:0] sel_557255;
  wire [7:0] add_557258;
  wire [7:0] sel_557259;
  wire [7:0] add_557262;
  wire [7:0] sel_557263;
  wire [7:0] add_557266;
  wire [7:0] sel_557267;
  wire [7:0] add_557270;
  wire [7:0] sel_557271;
  wire [7:0] add_557274;
  wire [7:0] sel_557275;
  wire [7:0] add_557278;
  wire [7:0] sel_557279;
  wire [7:0] add_557282;
  wire [7:0] sel_557283;
  wire [7:0] add_557286;
  wire [7:0] sel_557287;
  wire [7:0] add_557290;
  wire [7:0] sel_557291;
  wire [7:0] add_557294;
  wire [7:0] sel_557295;
  wire [7:0] add_557298;
  wire [7:0] sel_557299;
  wire [7:0] add_557302;
  wire [7:0] sel_557303;
  wire [7:0] add_557306;
  wire [7:0] sel_557307;
  wire [7:0] add_557310;
  wire [7:0] sel_557311;
  wire [7:0] add_557314;
  wire [7:0] sel_557315;
  wire [7:0] add_557318;
  wire [7:0] sel_557319;
  wire [7:0] add_557322;
  wire [7:0] sel_557323;
  wire [7:0] add_557326;
  wire [7:0] sel_557327;
  wire [7:0] add_557330;
  wire [7:0] sel_557331;
  wire [7:0] add_557334;
  wire [7:0] sel_557335;
  wire [7:0] add_557338;
  wire [7:0] sel_557339;
  wire [7:0] add_557342;
  wire [7:0] sel_557343;
  wire [7:0] add_557346;
  wire [7:0] sel_557347;
  wire [7:0] add_557350;
  wire [7:0] sel_557351;
  wire [7:0] add_557354;
  wire [7:0] sel_557355;
  wire [7:0] add_557358;
  wire [7:0] sel_557359;
  wire [7:0] add_557362;
  wire [7:0] sel_557363;
  wire [7:0] add_557366;
  wire [7:0] sel_557367;
  wire [7:0] add_557370;
  wire [7:0] sel_557371;
  wire [7:0] add_557374;
  wire [7:0] sel_557375;
  wire [7:0] add_557378;
  wire [7:0] sel_557379;
  wire [7:0] add_557382;
  wire [7:0] sel_557383;
  wire [7:0] add_557386;
  wire [7:0] sel_557387;
  wire [7:0] add_557390;
  wire [7:0] sel_557391;
  wire [7:0] add_557394;
  wire [7:0] sel_557395;
  wire [7:0] add_557398;
  wire [7:0] sel_557399;
  wire [7:0] add_557403;
  wire [15:0] array_index_557404;
  wire [7:0] sel_557405;
  wire [7:0] add_557408;
  wire [7:0] sel_557409;
  wire [7:0] add_557412;
  wire [7:0] sel_557413;
  wire [7:0] add_557416;
  wire [7:0] sel_557417;
  wire [7:0] add_557420;
  wire [7:0] sel_557421;
  wire [7:0] add_557424;
  wire [7:0] sel_557425;
  wire [7:0] add_557428;
  wire [7:0] sel_557429;
  wire [7:0] add_557432;
  wire [7:0] sel_557433;
  wire [7:0] add_557436;
  wire [7:0] sel_557437;
  wire [7:0] add_557440;
  wire [7:0] sel_557441;
  wire [7:0] add_557444;
  wire [7:0] sel_557445;
  wire [7:0] add_557448;
  wire [7:0] sel_557449;
  wire [7:0] add_557452;
  wire [7:0] sel_557453;
  wire [7:0] add_557456;
  wire [7:0] sel_557457;
  wire [7:0] add_557460;
  wire [7:0] sel_557461;
  wire [7:0] add_557464;
  wire [7:0] sel_557465;
  wire [7:0] add_557468;
  wire [7:0] sel_557469;
  wire [7:0] add_557472;
  wire [7:0] sel_557473;
  wire [7:0] add_557476;
  wire [7:0] sel_557477;
  wire [7:0] add_557480;
  wire [7:0] sel_557481;
  wire [7:0] add_557484;
  wire [7:0] sel_557485;
  wire [7:0] add_557488;
  wire [7:0] sel_557489;
  wire [7:0] add_557492;
  wire [7:0] sel_557493;
  wire [7:0] add_557496;
  wire [7:0] sel_557497;
  wire [7:0] add_557500;
  wire [7:0] sel_557501;
  wire [7:0] add_557504;
  wire [7:0] sel_557505;
  wire [7:0] add_557508;
  wire [7:0] sel_557509;
  wire [7:0] add_557512;
  wire [7:0] sel_557513;
  wire [7:0] add_557516;
  wire [7:0] sel_557517;
  wire [7:0] add_557520;
  wire [7:0] sel_557521;
  wire [7:0] add_557524;
  wire [7:0] sel_557525;
  wire [7:0] add_557528;
  wire [7:0] sel_557529;
  wire [7:0] add_557532;
  wire [7:0] sel_557533;
  wire [7:0] add_557536;
  wire [7:0] sel_557537;
  wire [7:0] add_557540;
  wire [7:0] sel_557541;
  wire [7:0] add_557544;
  wire [7:0] sel_557545;
  wire [7:0] add_557548;
  wire [7:0] sel_557549;
  wire [7:0] add_557552;
  wire [7:0] sel_557553;
  wire [7:0] add_557556;
  wire [7:0] sel_557557;
  wire [7:0] add_557560;
  wire [7:0] sel_557561;
  wire [7:0] add_557564;
  wire [7:0] sel_557565;
  wire [7:0] add_557568;
  wire [7:0] sel_557569;
  wire [7:0] add_557572;
  wire [7:0] sel_557573;
  wire [7:0] add_557576;
  wire [7:0] sel_557577;
  wire [7:0] add_557580;
  wire [7:0] sel_557581;
  wire [7:0] add_557584;
  wire [7:0] sel_557585;
  wire [7:0] add_557588;
  wire [7:0] sel_557589;
  wire [7:0] add_557592;
  wire [7:0] sel_557593;
  wire [7:0] add_557596;
  wire [7:0] sel_557597;
  wire [7:0] add_557600;
  wire [7:0] sel_557601;
  wire [7:0] add_557604;
  wire [7:0] sel_557605;
  wire [7:0] add_557608;
  wire [7:0] sel_557609;
  wire [7:0] add_557612;
  wire [7:0] sel_557613;
  wire [7:0] add_557616;
  wire [7:0] sel_557617;
  wire [7:0] add_557620;
  wire [7:0] sel_557621;
  wire [7:0] add_557624;
  wire [7:0] sel_557625;
  wire [7:0] add_557628;
  wire [7:0] sel_557629;
  wire [7:0] add_557632;
  wire [7:0] sel_557633;
  wire [7:0] add_557636;
  wire [7:0] sel_557637;
  wire [7:0] add_557640;
  wire [7:0] sel_557641;
  wire [7:0] add_557644;
  wire [7:0] sel_557645;
  wire [7:0] add_557648;
  wire [7:0] sel_557649;
  wire [7:0] add_557652;
  wire [7:0] sel_557653;
  wire [7:0] add_557656;
  wire [7:0] sel_557657;
  wire [7:0] add_557660;
  wire [7:0] sel_557661;
  wire [7:0] add_557664;
  wire [7:0] sel_557665;
  wire [7:0] add_557668;
  wire [7:0] sel_557669;
  wire [7:0] add_557672;
  wire [7:0] sel_557673;
  wire [7:0] add_557676;
  wire [7:0] sel_557677;
  wire [7:0] add_557680;
  wire [7:0] sel_557681;
  wire [7:0] add_557684;
  wire [7:0] sel_557685;
  wire [7:0] add_557688;
  wire [7:0] sel_557689;
  wire [7:0] add_557692;
  wire [7:0] sel_557693;
  wire [7:0] add_557696;
  wire [7:0] sel_557697;
  wire [7:0] add_557700;
  wire [7:0] sel_557701;
  wire [7:0] add_557705;
  wire [15:0] array_index_557706;
  wire [7:0] sel_557707;
  wire [7:0] add_557710;
  wire [7:0] sel_557711;
  wire [7:0] add_557714;
  wire [7:0] sel_557715;
  wire [7:0] add_557718;
  wire [7:0] sel_557719;
  wire [7:0] add_557722;
  wire [7:0] sel_557723;
  wire [7:0] add_557726;
  wire [7:0] sel_557727;
  wire [7:0] add_557730;
  wire [7:0] sel_557731;
  wire [7:0] add_557734;
  wire [7:0] sel_557735;
  wire [7:0] add_557738;
  wire [7:0] sel_557739;
  wire [7:0] add_557742;
  wire [7:0] sel_557743;
  wire [7:0] add_557746;
  wire [7:0] sel_557747;
  wire [7:0] add_557750;
  wire [7:0] sel_557751;
  wire [7:0] add_557754;
  wire [7:0] sel_557755;
  wire [7:0] add_557758;
  wire [7:0] sel_557759;
  wire [7:0] add_557762;
  wire [7:0] sel_557763;
  wire [7:0] add_557766;
  wire [7:0] sel_557767;
  wire [7:0] add_557770;
  wire [7:0] sel_557771;
  wire [7:0] add_557774;
  wire [7:0] sel_557775;
  wire [7:0] add_557778;
  wire [7:0] sel_557779;
  wire [7:0] add_557782;
  wire [7:0] sel_557783;
  wire [7:0] add_557786;
  wire [7:0] sel_557787;
  wire [7:0] add_557790;
  wire [7:0] sel_557791;
  wire [7:0] add_557794;
  wire [7:0] sel_557795;
  wire [7:0] add_557798;
  wire [7:0] sel_557799;
  wire [7:0] add_557802;
  wire [7:0] sel_557803;
  wire [7:0] add_557806;
  wire [7:0] sel_557807;
  wire [7:0] add_557810;
  wire [7:0] sel_557811;
  wire [7:0] add_557814;
  wire [7:0] sel_557815;
  wire [7:0] add_557818;
  wire [7:0] sel_557819;
  wire [7:0] add_557822;
  wire [7:0] sel_557823;
  wire [7:0] add_557826;
  wire [7:0] sel_557827;
  wire [7:0] add_557830;
  wire [7:0] sel_557831;
  wire [7:0] add_557834;
  wire [7:0] sel_557835;
  wire [7:0] add_557838;
  wire [7:0] sel_557839;
  wire [7:0] add_557842;
  wire [7:0] sel_557843;
  wire [7:0] add_557846;
  wire [7:0] sel_557847;
  wire [7:0] add_557850;
  wire [7:0] sel_557851;
  wire [7:0] add_557854;
  wire [7:0] sel_557855;
  wire [7:0] add_557858;
  wire [7:0] sel_557859;
  wire [7:0] add_557862;
  wire [7:0] sel_557863;
  wire [7:0] add_557866;
  wire [7:0] sel_557867;
  wire [7:0] add_557870;
  wire [7:0] sel_557871;
  wire [7:0] add_557874;
  wire [7:0] sel_557875;
  wire [7:0] add_557878;
  wire [7:0] sel_557879;
  wire [7:0] add_557882;
  wire [7:0] sel_557883;
  wire [7:0] add_557886;
  wire [7:0] sel_557887;
  wire [7:0] add_557890;
  wire [7:0] sel_557891;
  wire [7:0] add_557894;
  wire [7:0] sel_557895;
  wire [7:0] add_557898;
  wire [7:0] sel_557899;
  wire [7:0] add_557902;
  wire [7:0] sel_557903;
  wire [7:0] add_557906;
  wire [7:0] sel_557907;
  wire [7:0] add_557910;
  wire [7:0] sel_557911;
  wire [7:0] add_557914;
  wire [7:0] sel_557915;
  wire [7:0] add_557918;
  wire [7:0] sel_557919;
  wire [7:0] add_557922;
  wire [7:0] sel_557923;
  wire [7:0] add_557926;
  wire [7:0] sel_557927;
  wire [7:0] add_557930;
  wire [7:0] sel_557931;
  wire [7:0] add_557934;
  wire [7:0] sel_557935;
  wire [7:0] add_557938;
  wire [7:0] sel_557939;
  wire [7:0] add_557942;
  wire [7:0] sel_557943;
  wire [7:0] add_557946;
  wire [7:0] sel_557947;
  wire [7:0] add_557950;
  wire [7:0] sel_557951;
  wire [7:0] add_557954;
  wire [7:0] sel_557955;
  wire [7:0] add_557958;
  wire [7:0] sel_557959;
  wire [7:0] add_557962;
  wire [7:0] sel_557963;
  wire [7:0] add_557966;
  wire [7:0] sel_557967;
  wire [7:0] add_557970;
  wire [7:0] sel_557971;
  wire [7:0] add_557974;
  wire [7:0] sel_557975;
  wire [7:0] add_557978;
  wire [7:0] sel_557979;
  wire [7:0] add_557982;
  wire [7:0] sel_557983;
  wire [7:0] add_557986;
  wire [7:0] sel_557987;
  wire [7:0] add_557990;
  wire [7:0] sel_557991;
  wire [7:0] add_557994;
  wire [7:0] sel_557995;
  wire [7:0] add_557998;
  wire [7:0] sel_557999;
  wire [7:0] add_558002;
  wire [7:0] sel_558003;
  wire [7:0] add_558007;
  wire [15:0] array_index_558008;
  wire [7:0] sel_558009;
  wire [7:0] add_558012;
  wire [7:0] sel_558013;
  wire [7:0] add_558016;
  wire [7:0] sel_558017;
  wire [7:0] add_558020;
  wire [7:0] sel_558021;
  wire [7:0] add_558024;
  wire [7:0] sel_558025;
  wire [7:0] add_558028;
  wire [7:0] sel_558029;
  wire [7:0] add_558032;
  wire [7:0] sel_558033;
  wire [7:0] add_558036;
  wire [7:0] sel_558037;
  wire [7:0] add_558040;
  wire [7:0] sel_558041;
  wire [7:0] add_558044;
  wire [7:0] sel_558045;
  wire [7:0] add_558048;
  wire [7:0] sel_558049;
  wire [7:0] add_558052;
  wire [7:0] sel_558053;
  wire [7:0] add_558056;
  wire [7:0] sel_558057;
  wire [7:0] add_558060;
  wire [7:0] sel_558061;
  wire [7:0] add_558064;
  wire [7:0] sel_558065;
  wire [7:0] add_558068;
  wire [7:0] sel_558069;
  wire [7:0] add_558072;
  wire [7:0] sel_558073;
  wire [7:0] add_558076;
  wire [7:0] sel_558077;
  wire [7:0] add_558080;
  wire [7:0] sel_558081;
  wire [7:0] add_558084;
  wire [7:0] sel_558085;
  wire [7:0] add_558088;
  wire [7:0] sel_558089;
  wire [7:0] add_558092;
  wire [7:0] sel_558093;
  wire [7:0] add_558096;
  wire [7:0] sel_558097;
  wire [7:0] add_558100;
  wire [7:0] sel_558101;
  wire [7:0] add_558104;
  wire [7:0] sel_558105;
  wire [7:0] add_558108;
  wire [7:0] sel_558109;
  wire [7:0] add_558112;
  wire [7:0] sel_558113;
  wire [7:0] add_558116;
  wire [7:0] sel_558117;
  wire [7:0] add_558120;
  wire [7:0] sel_558121;
  wire [7:0] add_558124;
  wire [7:0] sel_558125;
  wire [7:0] add_558128;
  wire [7:0] sel_558129;
  wire [7:0] add_558132;
  wire [7:0] sel_558133;
  wire [7:0] add_558136;
  wire [7:0] sel_558137;
  wire [7:0] add_558140;
  wire [7:0] sel_558141;
  wire [7:0] add_558144;
  wire [7:0] sel_558145;
  wire [7:0] add_558148;
  wire [7:0] sel_558149;
  wire [7:0] add_558152;
  wire [7:0] sel_558153;
  wire [7:0] add_558156;
  wire [7:0] sel_558157;
  wire [7:0] add_558160;
  wire [7:0] sel_558161;
  wire [7:0] add_558164;
  wire [7:0] sel_558165;
  wire [7:0] add_558168;
  wire [7:0] sel_558169;
  wire [7:0] add_558172;
  wire [7:0] sel_558173;
  wire [7:0] add_558176;
  wire [7:0] sel_558177;
  wire [7:0] add_558180;
  wire [7:0] sel_558181;
  wire [7:0] add_558184;
  wire [7:0] sel_558185;
  wire [7:0] add_558188;
  wire [7:0] sel_558189;
  wire [7:0] add_558192;
  wire [7:0] sel_558193;
  wire [7:0] add_558196;
  wire [7:0] sel_558197;
  wire [7:0] add_558200;
  wire [7:0] sel_558201;
  wire [7:0] add_558204;
  wire [7:0] sel_558205;
  wire [7:0] add_558208;
  wire [7:0] sel_558209;
  wire [7:0] add_558212;
  wire [7:0] sel_558213;
  wire [7:0] add_558216;
  wire [7:0] sel_558217;
  wire [7:0] add_558220;
  wire [7:0] sel_558221;
  wire [7:0] add_558224;
  wire [7:0] sel_558225;
  wire [7:0] add_558228;
  wire [7:0] sel_558229;
  wire [7:0] add_558232;
  wire [7:0] sel_558233;
  wire [7:0] add_558236;
  wire [7:0] sel_558237;
  wire [7:0] add_558240;
  wire [7:0] sel_558241;
  wire [7:0] add_558244;
  wire [7:0] sel_558245;
  wire [7:0] add_558248;
  wire [7:0] sel_558249;
  wire [7:0] add_558252;
  wire [7:0] sel_558253;
  wire [7:0] add_558256;
  wire [7:0] sel_558257;
  wire [7:0] add_558260;
  wire [7:0] sel_558261;
  wire [7:0] add_558264;
  wire [7:0] sel_558265;
  wire [7:0] add_558268;
  wire [7:0] sel_558269;
  wire [7:0] add_558272;
  wire [7:0] sel_558273;
  wire [7:0] add_558276;
  wire [7:0] sel_558277;
  wire [7:0] add_558280;
  wire [7:0] sel_558281;
  wire [7:0] add_558284;
  wire [7:0] sel_558285;
  wire [7:0] add_558288;
  wire [7:0] sel_558289;
  wire [7:0] add_558292;
  wire [7:0] sel_558293;
  wire [7:0] add_558296;
  wire [7:0] sel_558297;
  wire [7:0] add_558300;
  wire [7:0] sel_558301;
  wire [7:0] add_558304;
  wire [7:0] sel_558305;
  wire [7:0] add_558309;
  wire [15:0] array_index_558310;
  wire [7:0] sel_558311;
  wire [7:0] add_558314;
  wire [7:0] sel_558315;
  wire [7:0] add_558318;
  wire [7:0] sel_558319;
  wire [7:0] add_558322;
  wire [7:0] sel_558323;
  wire [7:0] add_558326;
  wire [7:0] sel_558327;
  wire [7:0] add_558330;
  wire [7:0] sel_558331;
  wire [7:0] add_558334;
  wire [7:0] sel_558335;
  wire [7:0] add_558338;
  wire [7:0] sel_558339;
  wire [7:0] add_558342;
  wire [7:0] sel_558343;
  wire [7:0] add_558346;
  wire [7:0] sel_558347;
  wire [7:0] add_558350;
  wire [7:0] sel_558351;
  wire [7:0] add_558354;
  wire [7:0] sel_558355;
  wire [7:0] add_558358;
  wire [7:0] sel_558359;
  wire [7:0] add_558362;
  wire [7:0] sel_558363;
  wire [7:0] add_558366;
  wire [7:0] sel_558367;
  wire [7:0] add_558370;
  wire [7:0] sel_558371;
  wire [7:0] add_558374;
  wire [7:0] sel_558375;
  wire [7:0] add_558378;
  wire [7:0] sel_558379;
  wire [7:0] add_558382;
  wire [7:0] sel_558383;
  wire [7:0] add_558386;
  wire [7:0] sel_558387;
  wire [7:0] add_558390;
  wire [7:0] sel_558391;
  wire [7:0] add_558394;
  wire [7:0] sel_558395;
  wire [7:0] add_558398;
  wire [7:0] sel_558399;
  wire [7:0] add_558402;
  wire [7:0] sel_558403;
  wire [7:0] add_558406;
  wire [7:0] sel_558407;
  wire [7:0] add_558410;
  wire [7:0] sel_558411;
  wire [7:0] add_558414;
  wire [7:0] sel_558415;
  wire [7:0] add_558418;
  wire [7:0] sel_558419;
  wire [7:0] add_558422;
  wire [7:0] sel_558423;
  wire [7:0] add_558426;
  wire [7:0] sel_558427;
  wire [7:0] add_558430;
  wire [7:0] sel_558431;
  wire [7:0] add_558434;
  wire [7:0] sel_558435;
  wire [7:0] add_558438;
  wire [7:0] sel_558439;
  wire [7:0] add_558442;
  wire [7:0] sel_558443;
  wire [7:0] add_558446;
  wire [7:0] sel_558447;
  wire [7:0] add_558450;
  wire [7:0] sel_558451;
  wire [7:0] add_558454;
  wire [7:0] sel_558455;
  wire [7:0] add_558458;
  wire [7:0] sel_558459;
  wire [7:0] add_558462;
  wire [7:0] sel_558463;
  wire [7:0] add_558466;
  wire [7:0] sel_558467;
  wire [7:0] add_558470;
  wire [7:0] sel_558471;
  wire [7:0] add_558474;
  wire [7:0] sel_558475;
  wire [7:0] add_558478;
  wire [7:0] sel_558479;
  wire [7:0] add_558482;
  wire [7:0] sel_558483;
  wire [7:0] add_558486;
  wire [7:0] sel_558487;
  wire [7:0] add_558490;
  wire [7:0] sel_558491;
  wire [7:0] add_558494;
  wire [7:0] sel_558495;
  wire [7:0] add_558498;
  wire [7:0] sel_558499;
  wire [7:0] add_558502;
  wire [7:0] sel_558503;
  wire [7:0] add_558506;
  wire [7:0] sel_558507;
  wire [7:0] add_558510;
  wire [7:0] sel_558511;
  wire [7:0] add_558514;
  wire [7:0] sel_558515;
  wire [7:0] add_558518;
  wire [7:0] sel_558519;
  wire [7:0] add_558522;
  wire [7:0] sel_558523;
  wire [7:0] add_558526;
  wire [7:0] sel_558527;
  wire [7:0] add_558530;
  wire [7:0] sel_558531;
  wire [7:0] add_558534;
  wire [7:0] sel_558535;
  wire [7:0] add_558538;
  wire [7:0] sel_558539;
  wire [7:0] add_558542;
  wire [7:0] sel_558543;
  wire [7:0] add_558546;
  wire [7:0] sel_558547;
  wire [7:0] add_558550;
  wire [7:0] sel_558551;
  wire [7:0] add_558554;
  wire [7:0] sel_558555;
  wire [7:0] add_558558;
  wire [7:0] sel_558559;
  wire [7:0] add_558562;
  wire [7:0] sel_558563;
  wire [7:0] add_558566;
  wire [7:0] sel_558567;
  wire [7:0] add_558570;
  wire [7:0] sel_558571;
  wire [7:0] add_558574;
  wire [7:0] sel_558575;
  wire [7:0] add_558578;
  wire [7:0] sel_558579;
  wire [7:0] add_558582;
  wire [7:0] sel_558583;
  wire [7:0] add_558586;
  wire [7:0] sel_558587;
  wire [7:0] add_558590;
  wire [7:0] sel_558591;
  wire [7:0] add_558594;
  wire [7:0] sel_558595;
  wire [7:0] add_558598;
  wire [7:0] sel_558599;
  wire [7:0] add_558602;
  wire [7:0] sel_558603;
  wire [7:0] add_558606;
  wire [7:0] sel_558607;
  wire [7:0] add_558611;
  wire [15:0] array_index_558612;
  wire [7:0] sel_558613;
  wire [7:0] add_558616;
  wire [7:0] sel_558617;
  wire [7:0] add_558620;
  wire [7:0] sel_558621;
  wire [7:0] add_558624;
  wire [7:0] sel_558625;
  wire [7:0] add_558628;
  wire [7:0] sel_558629;
  wire [7:0] add_558632;
  wire [7:0] sel_558633;
  wire [7:0] add_558636;
  wire [7:0] sel_558637;
  wire [7:0] add_558640;
  wire [7:0] sel_558641;
  wire [7:0] add_558644;
  wire [7:0] sel_558645;
  wire [7:0] add_558648;
  wire [7:0] sel_558649;
  wire [7:0] add_558652;
  wire [7:0] sel_558653;
  wire [7:0] add_558656;
  wire [7:0] sel_558657;
  wire [7:0] add_558660;
  wire [7:0] sel_558661;
  wire [7:0] add_558664;
  wire [7:0] sel_558665;
  wire [7:0] add_558668;
  wire [7:0] sel_558669;
  wire [7:0] add_558672;
  wire [7:0] sel_558673;
  wire [7:0] add_558676;
  wire [7:0] sel_558677;
  wire [7:0] add_558680;
  wire [7:0] sel_558681;
  wire [7:0] add_558684;
  wire [7:0] sel_558685;
  wire [7:0] add_558688;
  wire [7:0] sel_558689;
  wire [7:0] add_558692;
  wire [7:0] sel_558693;
  wire [7:0] add_558696;
  wire [7:0] sel_558697;
  wire [7:0] add_558700;
  wire [7:0] sel_558701;
  wire [7:0] add_558704;
  wire [7:0] sel_558705;
  wire [7:0] add_558708;
  wire [7:0] sel_558709;
  wire [7:0] add_558712;
  wire [7:0] sel_558713;
  wire [7:0] add_558716;
  wire [7:0] sel_558717;
  wire [7:0] add_558720;
  wire [7:0] sel_558721;
  wire [7:0] add_558724;
  wire [7:0] sel_558725;
  wire [7:0] add_558728;
  wire [7:0] sel_558729;
  wire [7:0] add_558732;
  wire [7:0] sel_558733;
  wire [7:0] add_558736;
  wire [7:0] sel_558737;
  wire [7:0] add_558740;
  wire [7:0] sel_558741;
  wire [7:0] add_558744;
  wire [7:0] sel_558745;
  wire [7:0] add_558748;
  wire [7:0] sel_558749;
  wire [7:0] add_558752;
  wire [7:0] sel_558753;
  wire [7:0] add_558756;
  wire [7:0] sel_558757;
  wire [7:0] add_558760;
  wire [7:0] sel_558761;
  wire [7:0] add_558764;
  wire [7:0] sel_558765;
  wire [7:0] add_558768;
  wire [7:0] sel_558769;
  wire [7:0] add_558772;
  wire [7:0] sel_558773;
  wire [7:0] add_558776;
  wire [7:0] sel_558777;
  wire [7:0] add_558780;
  wire [7:0] sel_558781;
  wire [7:0] add_558784;
  wire [7:0] sel_558785;
  wire [7:0] add_558788;
  wire [7:0] sel_558789;
  wire [7:0] add_558792;
  wire [7:0] sel_558793;
  wire [7:0] add_558796;
  wire [7:0] sel_558797;
  wire [7:0] add_558800;
  wire [7:0] sel_558801;
  wire [7:0] add_558804;
  wire [7:0] sel_558805;
  wire [7:0] add_558808;
  wire [7:0] sel_558809;
  wire [7:0] add_558812;
  wire [7:0] sel_558813;
  wire [7:0] add_558816;
  wire [7:0] sel_558817;
  wire [7:0] add_558820;
  wire [7:0] sel_558821;
  wire [7:0] add_558824;
  wire [7:0] sel_558825;
  wire [7:0] add_558828;
  wire [7:0] sel_558829;
  wire [7:0] add_558832;
  wire [7:0] sel_558833;
  wire [7:0] add_558836;
  wire [7:0] sel_558837;
  wire [7:0] add_558840;
  wire [7:0] sel_558841;
  wire [7:0] add_558844;
  wire [7:0] sel_558845;
  wire [7:0] add_558848;
  wire [7:0] sel_558849;
  wire [7:0] add_558852;
  wire [7:0] sel_558853;
  wire [7:0] add_558856;
  wire [7:0] sel_558857;
  wire [7:0] add_558860;
  wire [7:0] sel_558861;
  wire [7:0] add_558864;
  wire [7:0] sel_558865;
  wire [7:0] add_558868;
  wire [7:0] sel_558869;
  wire [7:0] add_558872;
  wire [7:0] sel_558873;
  wire [7:0] add_558876;
  wire [7:0] sel_558877;
  wire [7:0] add_558880;
  wire [7:0] sel_558881;
  wire [7:0] add_558884;
  wire [7:0] sel_558885;
  wire [7:0] add_558888;
  wire [7:0] sel_558889;
  wire [7:0] add_558892;
  wire [7:0] sel_558893;
  wire [7:0] add_558896;
  wire [7:0] sel_558897;
  wire [7:0] add_558900;
  wire [7:0] sel_558901;
  wire [7:0] add_558904;
  wire [7:0] sel_558905;
  wire [7:0] add_558908;
  wire [7:0] sel_558909;
  wire [7:0] add_558913;
  wire [15:0] array_index_558914;
  wire [7:0] sel_558915;
  wire [7:0] add_558918;
  wire [7:0] sel_558919;
  wire [7:0] add_558922;
  wire [7:0] sel_558923;
  wire [7:0] add_558926;
  wire [7:0] sel_558927;
  wire [7:0] add_558930;
  wire [7:0] sel_558931;
  wire [7:0] add_558934;
  wire [7:0] sel_558935;
  wire [7:0] add_558938;
  wire [7:0] sel_558939;
  wire [7:0] add_558942;
  wire [7:0] sel_558943;
  wire [7:0] add_558946;
  wire [7:0] sel_558947;
  wire [7:0] add_558950;
  wire [7:0] sel_558951;
  wire [7:0] add_558954;
  wire [7:0] sel_558955;
  wire [7:0] add_558958;
  wire [7:0] sel_558959;
  wire [7:0] add_558962;
  wire [7:0] sel_558963;
  wire [7:0] add_558966;
  wire [7:0] sel_558967;
  wire [7:0] add_558970;
  wire [7:0] sel_558971;
  wire [7:0] add_558974;
  wire [7:0] sel_558975;
  wire [7:0] add_558978;
  wire [7:0] sel_558979;
  wire [7:0] add_558982;
  wire [7:0] sel_558983;
  wire [7:0] add_558986;
  wire [7:0] sel_558987;
  wire [7:0] add_558990;
  wire [7:0] sel_558991;
  wire [7:0] add_558994;
  wire [7:0] sel_558995;
  wire [7:0] add_558998;
  wire [7:0] sel_558999;
  wire [7:0] add_559002;
  wire [7:0] sel_559003;
  wire [7:0] add_559006;
  wire [7:0] sel_559007;
  wire [7:0] add_559010;
  wire [7:0] sel_559011;
  wire [7:0] add_559014;
  wire [7:0] sel_559015;
  wire [7:0] add_559018;
  wire [7:0] sel_559019;
  wire [7:0] add_559022;
  wire [7:0] sel_559023;
  wire [7:0] add_559026;
  wire [7:0] sel_559027;
  wire [7:0] add_559030;
  wire [7:0] sel_559031;
  wire [7:0] add_559034;
  wire [7:0] sel_559035;
  wire [7:0] add_559038;
  wire [7:0] sel_559039;
  wire [7:0] add_559042;
  wire [7:0] sel_559043;
  wire [7:0] add_559046;
  wire [7:0] sel_559047;
  wire [7:0] add_559050;
  wire [7:0] sel_559051;
  wire [7:0] add_559054;
  wire [7:0] sel_559055;
  wire [7:0] add_559058;
  wire [7:0] sel_559059;
  wire [7:0] add_559062;
  wire [7:0] sel_559063;
  wire [7:0] add_559066;
  wire [7:0] sel_559067;
  wire [7:0] add_559070;
  wire [7:0] sel_559071;
  wire [7:0] add_559074;
  wire [7:0] sel_559075;
  wire [7:0] add_559078;
  wire [7:0] sel_559079;
  wire [7:0] add_559082;
  wire [7:0] sel_559083;
  wire [7:0] add_559086;
  wire [7:0] sel_559087;
  wire [7:0] add_559090;
  wire [7:0] sel_559091;
  wire [7:0] add_559094;
  wire [7:0] sel_559095;
  wire [7:0] add_559098;
  wire [7:0] sel_559099;
  wire [7:0] add_559102;
  wire [7:0] sel_559103;
  wire [7:0] add_559106;
  wire [7:0] sel_559107;
  wire [7:0] add_559110;
  wire [7:0] sel_559111;
  wire [7:0] add_559114;
  wire [7:0] sel_559115;
  wire [7:0] add_559118;
  wire [7:0] sel_559119;
  wire [7:0] add_559122;
  wire [7:0] sel_559123;
  wire [7:0] add_559126;
  wire [7:0] sel_559127;
  wire [7:0] add_559130;
  wire [7:0] sel_559131;
  wire [7:0] add_559134;
  wire [7:0] sel_559135;
  wire [7:0] add_559138;
  wire [7:0] sel_559139;
  wire [7:0] add_559142;
  wire [7:0] sel_559143;
  wire [7:0] add_559146;
  wire [7:0] sel_559147;
  wire [7:0] add_559150;
  wire [7:0] sel_559151;
  wire [7:0] add_559154;
  wire [7:0] sel_559155;
  wire [7:0] add_559158;
  wire [7:0] sel_559159;
  wire [7:0] add_559162;
  wire [7:0] sel_559163;
  wire [7:0] add_559166;
  wire [7:0] sel_559167;
  wire [7:0] add_559170;
  wire [7:0] sel_559171;
  wire [7:0] add_559174;
  wire [7:0] sel_559175;
  wire [7:0] add_559178;
  wire [7:0] sel_559179;
  wire [7:0] add_559182;
  wire [7:0] sel_559183;
  wire [7:0] add_559186;
  wire [7:0] sel_559187;
  wire [7:0] add_559190;
  wire [7:0] sel_559191;
  wire [7:0] add_559194;
  wire [7:0] sel_559195;
  wire [7:0] add_559198;
  wire [7:0] sel_559199;
  wire [7:0] add_559202;
  wire [7:0] sel_559203;
  wire [7:0] add_559206;
  wire [7:0] sel_559207;
  wire [7:0] add_559210;
  wire [7:0] sel_559211;
  wire [7:0] add_559215;
  wire [15:0] array_index_559216;
  wire [7:0] sel_559217;
  wire [7:0] add_559220;
  wire [7:0] sel_559221;
  wire [7:0] add_559224;
  wire [7:0] sel_559225;
  wire [7:0] add_559228;
  wire [7:0] sel_559229;
  wire [7:0] add_559232;
  wire [7:0] sel_559233;
  wire [7:0] add_559236;
  wire [7:0] sel_559237;
  wire [7:0] add_559240;
  wire [7:0] sel_559241;
  wire [7:0] add_559244;
  wire [7:0] sel_559245;
  wire [7:0] add_559248;
  wire [7:0] sel_559249;
  wire [7:0] add_559252;
  wire [7:0] sel_559253;
  wire [7:0] add_559256;
  wire [7:0] sel_559257;
  wire [7:0] add_559260;
  wire [7:0] sel_559261;
  wire [7:0] add_559264;
  wire [7:0] sel_559265;
  wire [7:0] add_559268;
  wire [7:0] sel_559269;
  wire [7:0] add_559272;
  wire [7:0] sel_559273;
  wire [7:0] add_559276;
  wire [7:0] sel_559277;
  wire [7:0] add_559280;
  wire [7:0] sel_559281;
  wire [7:0] add_559284;
  wire [7:0] sel_559285;
  wire [7:0] add_559288;
  wire [7:0] sel_559289;
  wire [7:0] add_559292;
  wire [7:0] sel_559293;
  wire [7:0] add_559296;
  wire [7:0] sel_559297;
  wire [7:0] add_559300;
  wire [7:0] sel_559301;
  wire [7:0] add_559304;
  wire [7:0] sel_559305;
  wire [7:0] add_559308;
  wire [7:0] sel_559309;
  wire [7:0] add_559312;
  wire [7:0] sel_559313;
  wire [7:0] add_559316;
  wire [7:0] sel_559317;
  wire [7:0] add_559320;
  wire [7:0] sel_559321;
  wire [7:0] add_559324;
  wire [7:0] sel_559325;
  wire [7:0] add_559328;
  wire [7:0] sel_559329;
  wire [7:0] add_559332;
  wire [7:0] sel_559333;
  wire [7:0] add_559336;
  wire [7:0] sel_559337;
  wire [7:0] add_559340;
  wire [7:0] sel_559341;
  wire [7:0] add_559344;
  wire [7:0] sel_559345;
  wire [7:0] add_559348;
  wire [7:0] sel_559349;
  wire [7:0] add_559352;
  wire [7:0] sel_559353;
  wire [7:0] add_559356;
  wire [7:0] sel_559357;
  wire [7:0] add_559360;
  wire [7:0] sel_559361;
  wire [7:0] add_559364;
  wire [7:0] sel_559365;
  wire [7:0] add_559368;
  wire [7:0] sel_559369;
  wire [7:0] add_559372;
  wire [7:0] sel_559373;
  wire [7:0] add_559376;
  wire [7:0] sel_559377;
  wire [7:0] add_559380;
  wire [7:0] sel_559381;
  wire [7:0] add_559384;
  wire [7:0] sel_559385;
  wire [7:0] add_559388;
  wire [7:0] sel_559389;
  wire [7:0] add_559392;
  wire [7:0] sel_559393;
  wire [7:0] add_559396;
  wire [7:0] sel_559397;
  wire [7:0] add_559400;
  wire [7:0] sel_559401;
  wire [7:0] add_559404;
  wire [7:0] sel_559405;
  wire [7:0] add_559408;
  wire [7:0] sel_559409;
  wire [7:0] add_559412;
  wire [7:0] sel_559413;
  wire [7:0] add_559416;
  wire [7:0] sel_559417;
  wire [7:0] add_559420;
  wire [7:0] sel_559421;
  wire [7:0] add_559424;
  wire [7:0] sel_559425;
  wire [7:0] add_559428;
  wire [7:0] sel_559429;
  wire [7:0] add_559432;
  wire [7:0] sel_559433;
  wire [7:0] add_559436;
  wire [7:0] sel_559437;
  wire [7:0] add_559440;
  wire [7:0] sel_559441;
  wire [7:0] add_559444;
  wire [7:0] sel_559445;
  wire [7:0] add_559448;
  wire [7:0] sel_559449;
  wire [7:0] add_559452;
  wire [7:0] sel_559453;
  wire [7:0] add_559456;
  wire [7:0] sel_559457;
  wire [7:0] add_559460;
  wire [7:0] sel_559461;
  wire [7:0] add_559464;
  wire [7:0] sel_559465;
  wire [7:0] add_559468;
  wire [7:0] sel_559469;
  wire [7:0] add_559472;
  wire [7:0] sel_559473;
  wire [7:0] add_559476;
  wire [7:0] sel_559477;
  wire [7:0] add_559480;
  wire [7:0] sel_559481;
  wire [7:0] add_559484;
  wire [7:0] sel_559485;
  wire [7:0] add_559488;
  wire [7:0] sel_559489;
  wire [7:0] add_559492;
  wire [7:0] sel_559493;
  wire [7:0] add_559496;
  wire [7:0] sel_559497;
  wire [7:0] add_559500;
  wire [7:0] sel_559501;
  wire [7:0] add_559504;
  wire [7:0] sel_559505;
  wire [7:0] add_559508;
  wire [7:0] sel_559509;
  wire [7:0] add_559512;
  wire [7:0] sel_559513;
  wire [7:0] add_559517;
  wire [15:0] array_index_559518;
  wire [7:0] sel_559519;
  wire [7:0] add_559522;
  wire [7:0] sel_559523;
  wire [7:0] add_559526;
  wire [7:0] sel_559527;
  wire [7:0] add_559530;
  wire [7:0] sel_559531;
  wire [7:0] add_559534;
  wire [7:0] sel_559535;
  wire [7:0] add_559538;
  wire [7:0] sel_559539;
  wire [7:0] add_559542;
  wire [7:0] sel_559543;
  wire [7:0] add_559546;
  wire [7:0] sel_559547;
  wire [7:0] add_559550;
  wire [7:0] sel_559551;
  wire [7:0] add_559554;
  wire [7:0] sel_559555;
  wire [7:0] add_559558;
  wire [7:0] sel_559559;
  wire [7:0] add_559562;
  wire [7:0] sel_559563;
  wire [7:0] add_559566;
  wire [7:0] sel_559567;
  wire [7:0] add_559570;
  wire [7:0] sel_559571;
  wire [7:0] add_559574;
  wire [7:0] sel_559575;
  wire [7:0] add_559578;
  wire [7:0] sel_559579;
  wire [7:0] add_559582;
  wire [7:0] sel_559583;
  wire [7:0] add_559586;
  wire [7:0] sel_559587;
  wire [7:0] add_559590;
  wire [7:0] sel_559591;
  wire [7:0] add_559594;
  wire [7:0] sel_559595;
  wire [7:0] add_559598;
  wire [7:0] sel_559599;
  wire [7:0] add_559602;
  wire [7:0] sel_559603;
  wire [7:0] add_559606;
  wire [7:0] sel_559607;
  wire [7:0] add_559610;
  wire [7:0] sel_559611;
  wire [7:0] add_559614;
  wire [7:0] sel_559615;
  wire [7:0] add_559618;
  wire [7:0] sel_559619;
  wire [7:0] add_559622;
  wire [7:0] sel_559623;
  wire [7:0] add_559626;
  wire [7:0] sel_559627;
  wire [7:0] add_559630;
  wire [7:0] sel_559631;
  wire [7:0] add_559634;
  wire [7:0] sel_559635;
  wire [7:0] add_559638;
  wire [7:0] sel_559639;
  wire [7:0] add_559642;
  wire [7:0] sel_559643;
  wire [7:0] add_559646;
  wire [7:0] sel_559647;
  wire [7:0] add_559650;
  wire [7:0] sel_559651;
  wire [7:0] add_559654;
  wire [7:0] sel_559655;
  wire [7:0] add_559658;
  wire [7:0] sel_559659;
  wire [7:0] add_559662;
  wire [7:0] sel_559663;
  wire [7:0] add_559666;
  wire [7:0] sel_559667;
  wire [7:0] add_559670;
  wire [7:0] sel_559671;
  wire [7:0] add_559674;
  wire [7:0] sel_559675;
  wire [7:0] add_559678;
  wire [7:0] sel_559679;
  wire [7:0] add_559682;
  wire [7:0] sel_559683;
  wire [7:0] add_559686;
  wire [7:0] sel_559687;
  wire [7:0] add_559690;
  wire [7:0] sel_559691;
  wire [7:0] add_559694;
  wire [7:0] sel_559695;
  wire [7:0] add_559698;
  wire [7:0] sel_559699;
  wire [7:0] add_559702;
  wire [7:0] sel_559703;
  wire [7:0] add_559706;
  wire [7:0] sel_559707;
  wire [7:0] add_559710;
  wire [7:0] sel_559711;
  wire [7:0] add_559714;
  wire [7:0] sel_559715;
  wire [7:0] add_559718;
  wire [7:0] sel_559719;
  wire [7:0] add_559722;
  wire [7:0] sel_559723;
  wire [7:0] add_559726;
  wire [7:0] sel_559727;
  wire [7:0] add_559730;
  wire [7:0] sel_559731;
  wire [7:0] add_559734;
  wire [7:0] sel_559735;
  wire [7:0] add_559738;
  wire [7:0] sel_559739;
  wire [7:0] add_559742;
  wire [7:0] sel_559743;
  wire [7:0] add_559746;
  wire [7:0] sel_559747;
  wire [7:0] add_559750;
  wire [7:0] sel_559751;
  wire [7:0] add_559754;
  wire [7:0] sel_559755;
  wire [7:0] add_559758;
  wire [7:0] sel_559759;
  wire [7:0] add_559762;
  wire [7:0] sel_559763;
  wire [7:0] add_559766;
  wire [7:0] sel_559767;
  wire [7:0] add_559770;
  wire [7:0] sel_559771;
  wire [7:0] add_559774;
  wire [7:0] sel_559775;
  wire [7:0] add_559778;
  wire [7:0] sel_559779;
  wire [7:0] add_559782;
  wire [7:0] sel_559783;
  wire [7:0] add_559786;
  wire [7:0] sel_559787;
  wire [7:0] add_559790;
  wire [7:0] sel_559791;
  wire [7:0] add_559794;
  wire [7:0] sel_559795;
  wire [7:0] add_559798;
  wire [7:0] sel_559799;
  wire [7:0] add_559802;
  wire [7:0] sel_559803;
  wire [7:0] add_559806;
  wire [7:0] sel_559807;
  wire [7:0] add_559810;
  wire [7:0] sel_559811;
  wire [7:0] add_559814;
  wire [7:0] sel_559815;
  wire [7:0] add_559818;
  assign array_index_537011 = set1_unflattened[7'h00];
  assign array_index_537012 = set2_unflattened[7'h00];
  assign array_index_537016 = set2_unflattened[7'h01];
  assign concat_537017 = {1'h0, array_index_537011 == array_index_537012};
  assign add_537020 = concat_537017 + 2'h1;
  assign array_index_537024 = set2_unflattened[7'h02];
  assign concat_537025 = {1'h0, array_index_537011 == array_index_537016 ? add_537020 : concat_537017};
  assign add_537028 = concat_537025 + 3'h1;
  assign array_index_537032 = set2_unflattened[7'h03];
  assign concat_537033 = {1'h0, array_index_537011 == array_index_537024 ? add_537028 : concat_537025};
  assign add_537036 = concat_537033 + 4'h1;
  assign array_index_537040 = set2_unflattened[7'h04];
  assign concat_537041 = {1'h0, array_index_537011 == array_index_537032 ? add_537036 : concat_537033};
  assign add_537044 = concat_537041 + 5'h01;
  assign array_index_537048 = set2_unflattened[7'h05];
  assign concat_537049 = {1'h0, array_index_537011 == array_index_537040 ? add_537044 : concat_537041};
  assign add_537052 = concat_537049 + 6'h01;
  assign array_index_537056 = set2_unflattened[7'h06];
  assign concat_537057 = {1'h0, array_index_537011 == array_index_537048 ? add_537052 : concat_537049};
  assign add_537060 = concat_537057 + 7'h01;
  assign array_index_537064 = set2_unflattened[7'h07];
  assign concat_537065 = {1'h0, array_index_537011 == array_index_537056 ? add_537060 : concat_537057};
  assign add_537069 = concat_537065 + 8'h01;
  assign array_index_537070 = set2_unflattened[7'h08];
  assign sel_537071 = array_index_537011 == array_index_537064 ? add_537069 : concat_537065;
  assign add_537075 = sel_537071 + 8'h01;
  assign array_index_537076 = set2_unflattened[7'h09];
  assign sel_537077 = array_index_537011 == array_index_537070 ? add_537075 : sel_537071;
  assign add_537081 = sel_537077 + 8'h01;
  assign array_index_537082 = set2_unflattened[7'h0a];
  assign sel_537083 = array_index_537011 == array_index_537076 ? add_537081 : sel_537077;
  assign add_537087 = sel_537083 + 8'h01;
  assign array_index_537088 = set2_unflattened[7'h0b];
  assign sel_537089 = array_index_537011 == array_index_537082 ? add_537087 : sel_537083;
  assign add_537093 = sel_537089 + 8'h01;
  assign array_index_537094 = set2_unflattened[7'h0c];
  assign sel_537095 = array_index_537011 == array_index_537088 ? add_537093 : sel_537089;
  assign add_537099 = sel_537095 + 8'h01;
  assign array_index_537100 = set2_unflattened[7'h0d];
  assign sel_537101 = array_index_537011 == array_index_537094 ? add_537099 : sel_537095;
  assign add_537105 = sel_537101 + 8'h01;
  assign array_index_537106 = set2_unflattened[7'h0e];
  assign sel_537107 = array_index_537011 == array_index_537100 ? add_537105 : sel_537101;
  assign add_537111 = sel_537107 + 8'h01;
  assign array_index_537112 = set2_unflattened[7'h0f];
  assign sel_537113 = array_index_537011 == array_index_537106 ? add_537111 : sel_537107;
  assign add_537117 = sel_537113 + 8'h01;
  assign array_index_537118 = set2_unflattened[7'h10];
  assign sel_537119 = array_index_537011 == array_index_537112 ? add_537117 : sel_537113;
  assign add_537123 = sel_537119 + 8'h01;
  assign array_index_537124 = set2_unflattened[7'h11];
  assign sel_537125 = array_index_537011 == array_index_537118 ? add_537123 : sel_537119;
  assign add_537129 = sel_537125 + 8'h01;
  assign array_index_537130 = set2_unflattened[7'h12];
  assign sel_537131 = array_index_537011 == array_index_537124 ? add_537129 : sel_537125;
  assign add_537135 = sel_537131 + 8'h01;
  assign array_index_537136 = set2_unflattened[7'h13];
  assign sel_537137 = array_index_537011 == array_index_537130 ? add_537135 : sel_537131;
  assign add_537141 = sel_537137 + 8'h01;
  assign array_index_537142 = set2_unflattened[7'h14];
  assign sel_537143 = array_index_537011 == array_index_537136 ? add_537141 : sel_537137;
  assign add_537147 = sel_537143 + 8'h01;
  assign array_index_537148 = set2_unflattened[7'h15];
  assign sel_537149 = array_index_537011 == array_index_537142 ? add_537147 : sel_537143;
  assign add_537153 = sel_537149 + 8'h01;
  assign array_index_537154 = set2_unflattened[7'h16];
  assign sel_537155 = array_index_537011 == array_index_537148 ? add_537153 : sel_537149;
  assign add_537159 = sel_537155 + 8'h01;
  assign array_index_537160 = set2_unflattened[7'h17];
  assign sel_537161 = array_index_537011 == array_index_537154 ? add_537159 : sel_537155;
  assign add_537165 = sel_537161 + 8'h01;
  assign array_index_537166 = set2_unflattened[7'h18];
  assign sel_537167 = array_index_537011 == array_index_537160 ? add_537165 : sel_537161;
  assign add_537171 = sel_537167 + 8'h01;
  assign array_index_537172 = set2_unflattened[7'h19];
  assign sel_537173 = array_index_537011 == array_index_537166 ? add_537171 : sel_537167;
  assign add_537177 = sel_537173 + 8'h01;
  assign array_index_537178 = set2_unflattened[7'h1a];
  assign sel_537179 = array_index_537011 == array_index_537172 ? add_537177 : sel_537173;
  assign add_537183 = sel_537179 + 8'h01;
  assign array_index_537184 = set2_unflattened[7'h1b];
  assign sel_537185 = array_index_537011 == array_index_537178 ? add_537183 : sel_537179;
  assign add_537189 = sel_537185 + 8'h01;
  assign array_index_537190 = set2_unflattened[7'h1c];
  assign sel_537191 = array_index_537011 == array_index_537184 ? add_537189 : sel_537185;
  assign add_537195 = sel_537191 + 8'h01;
  assign array_index_537196 = set2_unflattened[7'h1d];
  assign sel_537197 = array_index_537011 == array_index_537190 ? add_537195 : sel_537191;
  assign add_537201 = sel_537197 + 8'h01;
  assign array_index_537202 = set2_unflattened[7'h1e];
  assign sel_537203 = array_index_537011 == array_index_537196 ? add_537201 : sel_537197;
  assign add_537207 = sel_537203 + 8'h01;
  assign array_index_537208 = set2_unflattened[7'h1f];
  assign sel_537209 = array_index_537011 == array_index_537202 ? add_537207 : sel_537203;
  assign add_537213 = sel_537209 + 8'h01;
  assign array_index_537214 = set2_unflattened[7'h20];
  assign sel_537215 = array_index_537011 == array_index_537208 ? add_537213 : sel_537209;
  assign add_537219 = sel_537215 + 8'h01;
  assign array_index_537220 = set2_unflattened[7'h21];
  assign sel_537221 = array_index_537011 == array_index_537214 ? add_537219 : sel_537215;
  assign add_537225 = sel_537221 + 8'h01;
  assign array_index_537226 = set2_unflattened[7'h22];
  assign sel_537227 = array_index_537011 == array_index_537220 ? add_537225 : sel_537221;
  assign add_537231 = sel_537227 + 8'h01;
  assign array_index_537232 = set2_unflattened[7'h23];
  assign sel_537233 = array_index_537011 == array_index_537226 ? add_537231 : sel_537227;
  assign add_537237 = sel_537233 + 8'h01;
  assign array_index_537238 = set2_unflattened[7'h24];
  assign sel_537239 = array_index_537011 == array_index_537232 ? add_537237 : sel_537233;
  assign add_537243 = sel_537239 + 8'h01;
  assign array_index_537244 = set2_unflattened[7'h25];
  assign sel_537245 = array_index_537011 == array_index_537238 ? add_537243 : sel_537239;
  assign add_537249 = sel_537245 + 8'h01;
  assign array_index_537250 = set2_unflattened[7'h26];
  assign sel_537251 = array_index_537011 == array_index_537244 ? add_537249 : sel_537245;
  assign add_537255 = sel_537251 + 8'h01;
  assign array_index_537256 = set2_unflattened[7'h27];
  assign sel_537257 = array_index_537011 == array_index_537250 ? add_537255 : sel_537251;
  assign add_537261 = sel_537257 + 8'h01;
  assign array_index_537262 = set2_unflattened[7'h28];
  assign sel_537263 = array_index_537011 == array_index_537256 ? add_537261 : sel_537257;
  assign add_537267 = sel_537263 + 8'h01;
  assign array_index_537268 = set2_unflattened[7'h29];
  assign sel_537269 = array_index_537011 == array_index_537262 ? add_537267 : sel_537263;
  assign add_537273 = sel_537269 + 8'h01;
  assign array_index_537274 = set2_unflattened[7'h2a];
  assign sel_537275 = array_index_537011 == array_index_537268 ? add_537273 : sel_537269;
  assign add_537279 = sel_537275 + 8'h01;
  assign array_index_537280 = set2_unflattened[7'h2b];
  assign sel_537281 = array_index_537011 == array_index_537274 ? add_537279 : sel_537275;
  assign add_537285 = sel_537281 + 8'h01;
  assign array_index_537286 = set2_unflattened[7'h2c];
  assign sel_537287 = array_index_537011 == array_index_537280 ? add_537285 : sel_537281;
  assign add_537291 = sel_537287 + 8'h01;
  assign array_index_537292 = set2_unflattened[7'h2d];
  assign sel_537293 = array_index_537011 == array_index_537286 ? add_537291 : sel_537287;
  assign add_537297 = sel_537293 + 8'h01;
  assign array_index_537298 = set2_unflattened[7'h2e];
  assign sel_537299 = array_index_537011 == array_index_537292 ? add_537297 : sel_537293;
  assign add_537303 = sel_537299 + 8'h01;
  assign array_index_537304 = set2_unflattened[7'h2f];
  assign sel_537305 = array_index_537011 == array_index_537298 ? add_537303 : sel_537299;
  assign add_537309 = sel_537305 + 8'h01;
  assign array_index_537310 = set2_unflattened[7'h30];
  assign sel_537311 = array_index_537011 == array_index_537304 ? add_537309 : sel_537305;
  assign add_537315 = sel_537311 + 8'h01;
  assign array_index_537316 = set2_unflattened[7'h31];
  assign sel_537317 = array_index_537011 == array_index_537310 ? add_537315 : sel_537311;
  assign add_537321 = sel_537317 + 8'h01;
  assign array_index_537322 = set2_unflattened[7'h32];
  assign sel_537323 = array_index_537011 == array_index_537316 ? add_537321 : sel_537317;
  assign add_537327 = sel_537323 + 8'h01;
  assign array_index_537328 = set2_unflattened[7'h33];
  assign sel_537329 = array_index_537011 == array_index_537322 ? add_537327 : sel_537323;
  assign add_537333 = sel_537329 + 8'h01;
  assign array_index_537334 = set2_unflattened[7'h34];
  assign sel_537335 = array_index_537011 == array_index_537328 ? add_537333 : sel_537329;
  assign add_537339 = sel_537335 + 8'h01;
  assign array_index_537340 = set2_unflattened[7'h35];
  assign sel_537341 = array_index_537011 == array_index_537334 ? add_537339 : sel_537335;
  assign add_537345 = sel_537341 + 8'h01;
  assign array_index_537346 = set2_unflattened[7'h36];
  assign sel_537347 = array_index_537011 == array_index_537340 ? add_537345 : sel_537341;
  assign add_537351 = sel_537347 + 8'h01;
  assign array_index_537352 = set2_unflattened[7'h37];
  assign sel_537353 = array_index_537011 == array_index_537346 ? add_537351 : sel_537347;
  assign add_537357 = sel_537353 + 8'h01;
  assign array_index_537358 = set2_unflattened[7'h38];
  assign sel_537359 = array_index_537011 == array_index_537352 ? add_537357 : sel_537353;
  assign add_537363 = sel_537359 + 8'h01;
  assign array_index_537364 = set2_unflattened[7'h39];
  assign sel_537365 = array_index_537011 == array_index_537358 ? add_537363 : sel_537359;
  assign add_537369 = sel_537365 + 8'h01;
  assign array_index_537370 = set2_unflattened[7'h3a];
  assign sel_537371 = array_index_537011 == array_index_537364 ? add_537369 : sel_537365;
  assign add_537375 = sel_537371 + 8'h01;
  assign array_index_537376 = set2_unflattened[7'h3b];
  assign sel_537377 = array_index_537011 == array_index_537370 ? add_537375 : sel_537371;
  assign add_537381 = sel_537377 + 8'h01;
  assign array_index_537382 = set2_unflattened[7'h3c];
  assign sel_537383 = array_index_537011 == array_index_537376 ? add_537381 : sel_537377;
  assign add_537387 = sel_537383 + 8'h01;
  assign array_index_537388 = set2_unflattened[7'h3d];
  assign sel_537389 = array_index_537011 == array_index_537382 ? add_537387 : sel_537383;
  assign add_537393 = sel_537389 + 8'h01;
  assign array_index_537394 = set2_unflattened[7'h3e];
  assign sel_537395 = array_index_537011 == array_index_537388 ? add_537393 : sel_537389;
  assign add_537399 = sel_537395 + 8'h01;
  assign array_index_537400 = set2_unflattened[7'h3f];
  assign sel_537401 = array_index_537011 == array_index_537394 ? add_537399 : sel_537395;
  assign add_537405 = sel_537401 + 8'h01;
  assign array_index_537406 = set2_unflattened[7'h40];
  assign sel_537407 = array_index_537011 == array_index_537400 ? add_537405 : sel_537401;
  assign add_537411 = sel_537407 + 8'h01;
  assign array_index_537412 = set2_unflattened[7'h41];
  assign sel_537413 = array_index_537011 == array_index_537406 ? add_537411 : sel_537407;
  assign add_537417 = sel_537413 + 8'h01;
  assign array_index_537418 = set2_unflattened[7'h42];
  assign sel_537419 = array_index_537011 == array_index_537412 ? add_537417 : sel_537413;
  assign add_537423 = sel_537419 + 8'h01;
  assign array_index_537424 = set2_unflattened[7'h43];
  assign sel_537425 = array_index_537011 == array_index_537418 ? add_537423 : sel_537419;
  assign add_537429 = sel_537425 + 8'h01;
  assign array_index_537430 = set2_unflattened[7'h44];
  assign sel_537431 = array_index_537011 == array_index_537424 ? add_537429 : sel_537425;
  assign add_537435 = sel_537431 + 8'h01;
  assign array_index_537436 = set2_unflattened[7'h45];
  assign sel_537437 = array_index_537011 == array_index_537430 ? add_537435 : sel_537431;
  assign add_537441 = sel_537437 + 8'h01;
  assign array_index_537442 = set2_unflattened[7'h46];
  assign sel_537443 = array_index_537011 == array_index_537436 ? add_537441 : sel_537437;
  assign add_537447 = sel_537443 + 8'h01;
  assign array_index_537448 = set2_unflattened[7'h47];
  assign sel_537449 = array_index_537011 == array_index_537442 ? add_537447 : sel_537443;
  assign add_537453 = sel_537449 + 8'h01;
  assign array_index_537454 = set2_unflattened[7'h48];
  assign sel_537455 = array_index_537011 == array_index_537448 ? add_537453 : sel_537449;
  assign add_537459 = sel_537455 + 8'h01;
  assign array_index_537460 = set2_unflattened[7'h49];
  assign sel_537461 = array_index_537011 == array_index_537454 ? add_537459 : sel_537455;
  assign add_537465 = sel_537461 + 8'h01;
  assign array_index_537466 = set2_unflattened[7'h4a];
  assign sel_537467 = array_index_537011 == array_index_537460 ? add_537465 : sel_537461;
  assign add_537471 = sel_537467 + 8'h01;
  assign array_index_537472 = set1_unflattened[7'h01];
  assign sel_537473 = array_index_537011 == array_index_537466 ? add_537471 : sel_537467;
  assign add_537476 = sel_537473 + 8'h01;
  assign sel_537477 = array_index_537472 == array_index_537012 ? add_537476 : sel_537473;
  assign add_537480 = sel_537477 + 8'h01;
  assign sel_537481 = array_index_537472 == array_index_537016 ? add_537480 : sel_537477;
  assign add_537484 = sel_537481 + 8'h01;
  assign sel_537485 = array_index_537472 == array_index_537024 ? add_537484 : sel_537481;
  assign add_537488 = sel_537485 + 8'h01;
  assign sel_537489 = array_index_537472 == array_index_537032 ? add_537488 : sel_537485;
  assign add_537492 = sel_537489 + 8'h01;
  assign sel_537493 = array_index_537472 == array_index_537040 ? add_537492 : sel_537489;
  assign add_537496 = sel_537493 + 8'h01;
  assign sel_537497 = array_index_537472 == array_index_537048 ? add_537496 : sel_537493;
  assign add_537500 = sel_537497 + 8'h01;
  assign sel_537501 = array_index_537472 == array_index_537056 ? add_537500 : sel_537497;
  assign add_537504 = sel_537501 + 8'h01;
  assign sel_537505 = array_index_537472 == array_index_537064 ? add_537504 : sel_537501;
  assign add_537508 = sel_537505 + 8'h01;
  assign sel_537509 = array_index_537472 == array_index_537070 ? add_537508 : sel_537505;
  assign add_537512 = sel_537509 + 8'h01;
  assign sel_537513 = array_index_537472 == array_index_537076 ? add_537512 : sel_537509;
  assign add_537516 = sel_537513 + 8'h01;
  assign sel_537517 = array_index_537472 == array_index_537082 ? add_537516 : sel_537513;
  assign add_537520 = sel_537517 + 8'h01;
  assign sel_537521 = array_index_537472 == array_index_537088 ? add_537520 : sel_537517;
  assign add_537524 = sel_537521 + 8'h01;
  assign sel_537525 = array_index_537472 == array_index_537094 ? add_537524 : sel_537521;
  assign add_537528 = sel_537525 + 8'h01;
  assign sel_537529 = array_index_537472 == array_index_537100 ? add_537528 : sel_537525;
  assign add_537532 = sel_537529 + 8'h01;
  assign sel_537533 = array_index_537472 == array_index_537106 ? add_537532 : sel_537529;
  assign add_537536 = sel_537533 + 8'h01;
  assign sel_537537 = array_index_537472 == array_index_537112 ? add_537536 : sel_537533;
  assign add_537540 = sel_537537 + 8'h01;
  assign sel_537541 = array_index_537472 == array_index_537118 ? add_537540 : sel_537537;
  assign add_537544 = sel_537541 + 8'h01;
  assign sel_537545 = array_index_537472 == array_index_537124 ? add_537544 : sel_537541;
  assign add_537548 = sel_537545 + 8'h01;
  assign sel_537549 = array_index_537472 == array_index_537130 ? add_537548 : sel_537545;
  assign add_537552 = sel_537549 + 8'h01;
  assign sel_537553 = array_index_537472 == array_index_537136 ? add_537552 : sel_537549;
  assign add_537556 = sel_537553 + 8'h01;
  assign sel_537557 = array_index_537472 == array_index_537142 ? add_537556 : sel_537553;
  assign add_537560 = sel_537557 + 8'h01;
  assign sel_537561 = array_index_537472 == array_index_537148 ? add_537560 : sel_537557;
  assign add_537564 = sel_537561 + 8'h01;
  assign sel_537565 = array_index_537472 == array_index_537154 ? add_537564 : sel_537561;
  assign add_537568 = sel_537565 + 8'h01;
  assign sel_537569 = array_index_537472 == array_index_537160 ? add_537568 : sel_537565;
  assign add_537572 = sel_537569 + 8'h01;
  assign sel_537573 = array_index_537472 == array_index_537166 ? add_537572 : sel_537569;
  assign add_537576 = sel_537573 + 8'h01;
  assign sel_537577 = array_index_537472 == array_index_537172 ? add_537576 : sel_537573;
  assign add_537580 = sel_537577 + 8'h01;
  assign sel_537581 = array_index_537472 == array_index_537178 ? add_537580 : sel_537577;
  assign add_537584 = sel_537581 + 8'h01;
  assign sel_537585 = array_index_537472 == array_index_537184 ? add_537584 : sel_537581;
  assign add_537588 = sel_537585 + 8'h01;
  assign sel_537589 = array_index_537472 == array_index_537190 ? add_537588 : sel_537585;
  assign add_537592 = sel_537589 + 8'h01;
  assign sel_537593 = array_index_537472 == array_index_537196 ? add_537592 : sel_537589;
  assign add_537596 = sel_537593 + 8'h01;
  assign sel_537597 = array_index_537472 == array_index_537202 ? add_537596 : sel_537593;
  assign add_537600 = sel_537597 + 8'h01;
  assign sel_537601 = array_index_537472 == array_index_537208 ? add_537600 : sel_537597;
  assign add_537604 = sel_537601 + 8'h01;
  assign sel_537605 = array_index_537472 == array_index_537214 ? add_537604 : sel_537601;
  assign add_537608 = sel_537605 + 8'h01;
  assign sel_537609 = array_index_537472 == array_index_537220 ? add_537608 : sel_537605;
  assign add_537612 = sel_537609 + 8'h01;
  assign sel_537613 = array_index_537472 == array_index_537226 ? add_537612 : sel_537609;
  assign add_537616 = sel_537613 + 8'h01;
  assign sel_537617 = array_index_537472 == array_index_537232 ? add_537616 : sel_537613;
  assign add_537620 = sel_537617 + 8'h01;
  assign sel_537621 = array_index_537472 == array_index_537238 ? add_537620 : sel_537617;
  assign add_537624 = sel_537621 + 8'h01;
  assign sel_537625 = array_index_537472 == array_index_537244 ? add_537624 : sel_537621;
  assign add_537628 = sel_537625 + 8'h01;
  assign sel_537629 = array_index_537472 == array_index_537250 ? add_537628 : sel_537625;
  assign add_537632 = sel_537629 + 8'h01;
  assign sel_537633 = array_index_537472 == array_index_537256 ? add_537632 : sel_537629;
  assign add_537636 = sel_537633 + 8'h01;
  assign sel_537637 = array_index_537472 == array_index_537262 ? add_537636 : sel_537633;
  assign add_537640 = sel_537637 + 8'h01;
  assign sel_537641 = array_index_537472 == array_index_537268 ? add_537640 : sel_537637;
  assign add_537644 = sel_537641 + 8'h01;
  assign sel_537645 = array_index_537472 == array_index_537274 ? add_537644 : sel_537641;
  assign add_537648 = sel_537645 + 8'h01;
  assign sel_537649 = array_index_537472 == array_index_537280 ? add_537648 : sel_537645;
  assign add_537652 = sel_537649 + 8'h01;
  assign sel_537653 = array_index_537472 == array_index_537286 ? add_537652 : sel_537649;
  assign add_537656 = sel_537653 + 8'h01;
  assign sel_537657 = array_index_537472 == array_index_537292 ? add_537656 : sel_537653;
  assign add_537660 = sel_537657 + 8'h01;
  assign sel_537661 = array_index_537472 == array_index_537298 ? add_537660 : sel_537657;
  assign add_537664 = sel_537661 + 8'h01;
  assign sel_537665 = array_index_537472 == array_index_537304 ? add_537664 : sel_537661;
  assign add_537668 = sel_537665 + 8'h01;
  assign sel_537669 = array_index_537472 == array_index_537310 ? add_537668 : sel_537665;
  assign add_537672 = sel_537669 + 8'h01;
  assign sel_537673 = array_index_537472 == array_index_537316 ? add_537672 : sel_537669;
  assign add_537676 = sel_537673 + 8'h01;
  assign sel_537677 = array_index_537472 == array_index_537322 ? add_537676 : sel_537673;
  assign add_537680 = sel_537677 + 8'h01;
  assign sel_537681 = array_index_537472 == array_index_537328 ? add_537680 : sel_537677;
  assign add_537684 = sel_537681 + 8'h01;
  assign sel_537685 = array_index_537472 == array_index_537334 ? add_537684 : sel_537681;
  assign add_537688 = sel_537685 + 8'h01;
  assign sel_537689 = array_index_537472 == array_index_537340 ? add_537688 : sel_537685;
  assign add_537692 = sel_537689 + 8'h01;
  assign sel_537693 = array_index_537472 == array_index_537346 ? add_537692 : sel_537689;
  assign add_537696 = sel_537693 + 8'h01;
  assign sel_537697 = array_index_537472 == array_index_537352 ? add_537696 : sel_537693;
  assign add_537700 = sel_537697 + 8'h01;
  assign sel_537701 = array_index_537472 == array_index_537358 ? add_537700 : sel_537697;
  assign add_537704 = sel_537701 + 8'h01;
  assign sel_537705 = array_index_537472 == array_index_537364 ? add_537704 : sel_537701;
  assign add_537708 = sel_537705 + 8'h01;
  assign sel_537709 = array_index_537472 == array_index_537370 ? add_537708 : sel_537705;
  assign add_537712 = sel_537709 + 8'h01;
  assign sel_537713 = array_index_537472 == array_index_537376 ? add_537712 : sel_537709;
  assign add_537716 = sel_537713 + 8'h01;
  assign sel_537717 = array_index_537472 == array_index_537382 ? add_537716 : sel_537713;
  assign add_537720 = sel_537717 + 8'h01;
  assign sel_537721 = array_index_537472 == array_index_537388 ? add_537720 : sel_537717;
  assign add_537724 = sel_537721 + 8'h01;
  assign sel_537725 = array_index_537472 == array_index_537394 ? add_537724 : sel_537721;
  assign add_537728 = sel_537725 + 8'h01;
  assign sel_537729 = array_index_537472 == array_index_537400 ? add_537728 : sel_537725;
  assign add_537732 = sel_537729 + 8'h01;
  assign sel_537733 = array_index_537472 == array_index_537406 ? add_537732 : sel_537729;
  assign add_537736 = sel_537733 + 8'h01;
  assign sel_537737 = array_index_537472 == array_index_537412 ? add_537736 : sel_537733;
  assign add_537740 = sel_537737 + 8'h01;
  assign sel_537741 = array_index_537472 == array_index_537418 ? add_537740 : sel_537737;
  assign add_537744 = sel_537741 + 8'h01;
  assign sel_537745 = array_index_537472 == array_index_537424 ? add_537744 : sel_537741;
  assign add_537748 = sel_537745 + 8'h01;
  assign sel_537749 = array_index_537472 == array_index_537430 ? add_537748 : sel_537745;
  assign add_537752 = sel_537749 + 8'h01;
  assign sel_537753 = array_index_537472 == array_index_537436 ? add_537752 : sel_537749;
  assign add_537756 = sel_537753 + 8'h01;
  assign sel_537757 = array_index_537472 == array_index_537442 ? add_537756 : sel_537753;
  assign add_537760 = sel_537757 + 8'h01;
  assign sel_537761 = array_index_537472 == array_index_537448 ? add_537760 : sel_537757;
  assign add_537764 = sel_537761 + 8'h01;
  assign sel_537765 = array_index_537472 == array_index_537454 ? add_537764 : sel_537761;
  assign add_537768 = sel_537765 + 8'h01;
  assign sel_537769 = array_index_537472 == array_index_537460 ? add_537768 : sel_537765;
  assign add_537773 = sel_537769 + 8'h01;
  assign array_index_537774 = set1_unflattened[7'h02];
  assign sel_537775 = array_index_537472 == array_index_537466 ? add_537773 : sel_537769;
  assign add_537778 = sel_537775 + 8'h01;
  assign sel_537779 = array_index_537774 == array_index_537012 ? add_537778 : sel_537775;
  assign add_537782 = sel_537779 + 8'h01;
  assign sel_537783 = array_index_537774 == array_index_537016 ? add_537782 : sel_537779;
  assign add_537786 = sel_537783 + 8'h01;
  assign sel_537787 = array_index_537774 == array_index_537024 ? add_537786 : sel_537783;
  assign add_537790 = sel_537787 + 8'h01;
  assign sel_537791 = array_index_537774 == array_index_537032 ? add_537790 : sel_537787;
  assign add_537794 = sel_537791 + 8'h01;
  assign sel_537795 = array_index_537774 == array_index_537040 ? add_537794 : sel_537791;
  assign add_537798 = sel_537795 + 8'h01;
  assign sel_537799 = array_index_537774 == array_index_537048 ? add_537798 : sel_537795;
  assign add_537802 = sel_537799 + 8'h01;
  assign sel_537803 = array_index_537774 == array_index_537056 ? add_537802 : sel_537799;
  assign add_537806 = sel_537803 + 8'h01;
  assign sel_537807 = array_index_537774 == array_index_537064 ? add_537806 : sel_537803;
  assign add_537810 = sel_537807 + 8'h01;
  assign sel_537811 = array_index_537774 == array_index_537070 ? add_537810 : sel_537807;
  assign add_537814 = sel_537811 + 8'h01;
  assign sel_537815 = array_index_537774 == array_index_537076 ? add_537814 : sel_537811;
  assign add_537818 = sel_537815 + 8'h01;
  assign sel_537819 = array_index_537774 == array_index_537082 ? add_537818 : sel_537815;
  assign add_537822 = sel_537819 + 8'h01;
  assign sel_537823 = array_index_537774 == array_index_537088 ? add_537822 : sel_537819;
  assign add_537826 = sel_537823 + 8'h01;
  assign sel_537827 = array_index_537774 == array_index_537094 ? add_537826 : sel_537823;
  assign add_537830 = sel_537827 + 8'h01;
  assign sel_537831 = array_index_537774 == array_index_537100 ? add_537830 : sel_537827;
  assign add_537834 = sel_537831 + 8'h01;
  assign sel_537835 = array_index_537774 == array_index_537106 ? add_537834 : sel_537831;
  assign add_537838 = sel_537835 + 8'h01;
  assign sel_537839 = array_index_537774 == array_index_537112 ? add_537838 : sel_537835;
  assign add_537842 = sel_537839 + 8'h01;
  assign sel_537843 = array_index_537774 == array_index_537118 ? add_537842 : sel_537839;
  assign add_537846 = sel_537843 + 8'h01;
  assign sel_537847 = array_index_537774 == array_index_537124 ? add_537846 : sel_537843;
  assign add_537850 = sel_537847 + 8'h01;
  assign sel_537851 = array_index_537774 == array_index_537130 ? add_537850 : sel_537847;
  assign add_537854 = sel_537851 + 8'h01;
  assign sel_537855 = array_index_537774 == array_index_537136 ? add_537854 : sel_537851;
  assign add_537858 = sel_537855 + 8'h01;
  assign sel_537859 = array_index_537774 == array_index_537142 ? add_537858 : sel_537855;
  assign add_537862 = sel_537859 + 8'h01;
  assign sel_537863 = array_index_537774 == array_index_537148 ? add_537862 : sel_537859;
  assign add_537866 = sel_537863 + 8'h01;
  assign sel_537867 = array_index_537774 == array_index_537154 ? add_537866 : sel_537863;
  assign add_537870 = sel_537867 + 8'h01;
  assign sel_537871 = array_index_537774 == array_index_537160 ? add_537870 : sel_537867;
  assign add_537874 = sel_537871 + 8'h01;
  assign sel_537875 = array_index_537774 == array_index_537166 ? add_537874 : sel_537871;
  assign add_537878 = sel_537875 + 8'h01;
  assign sel_537879 = array_index_537774 == array_index_537172 ? add_537878 : sel_537875;
  assign add_537882 = sel_537879 + 8'h01;
  assign sel_537883 = array_index_537774 == array_index_537178 ? add_537882 : sel_537879;
  assign add_537886 = sel_537883 + 8'h01;
  assign sel_537887 = array_index_537774 == array_index_537184 ? add_537886 : sel_537883;
  assign add_537890 = sel_537887 + 8'h01;
  assign sel_537891 = array_index_537774 == array_index_537190 ? add_537890 : sel_537887;
  assign add_537894 = sel_537891 + 8'h01;
  assign sel_537895 = array_index_537774 == array_index_537196 ? add_537894 : sel_537891;
  assign add_537898 = sel_537895 + 8'h01;
  assign sel_537899 = array_index_537774 == array_index_537202 ? add_537898 : sel_537895;
  assign add_537902 = sel_537899 + 8'h01;
  assign sel_537903 = array_index_537774 == array_index_537208 ? add_537902 : sel_537899;
  assign add_537906 = sel_537903 + 8'h01;
  assign sel_537907 = array_index_537774 == array_index_537214 ? add_537906 : sel_537903;
  assign add_537910 = sel_537907 + 8'h01;
  assign sel_537911 = array_index_537774 == array_index_537220 ? add_537910 : sel_537907;
  assign add_537914 = sel_537911 + 8'h01;
  assign sel_537915 = array_index_537774 == array_index_537226 ? add_537914 : sel_537911;
  assign add_537918 = sel_537915 + 8'h01;
  assign sel_537919 = array_index_537774 == array_index_537232 ? add_537918 : sel_537915;
  assign add_537922 = sel_537919 + 8'h01;
  assign sel_537923 = array_index_537774 == array_index_537238 ? add_537922 : sel_537919;
  assign add_537926 = sel_537923 + 8'h01;
  assign sel_537927 = array_index_537774 == array_index_537244 ? add_537926 : sel_537923;
  assign add_537930 = sel_537927 + 8'h01;
  assign sel_537931 = array_index_537774 == array_index_537250 ? add_537930 : sel_537927;
  assign add_537934 = sel_537931 + 8'h01;
  assign sel_537935 = array_index_537774 == array_index_537256 ? add_537934 : sel_537931;
  assign add_537938 = sel_537935 + 8'h01;
  assign sel_537939 = array_index_537774 == array_index_537262 ? add_537938 : sel_537935;
  assign add_537942 = sel_537939 + 8'h01;
  assign sel_537943 = array_index_537774 == array_index_537268 ? add_537942 : sel_537939;
  assign add_537946 = sel_537943 + 8'h01;
  assign sel_537947 = array_index_537774 == array_index_537274 ? add_537946 : sel_537943;
  assign add_537950 = sel_537947 + 8'h01;
  assign sel_537951 = array_index_537774 == array_index_537280 ? add_537950 : sel_537947;
  assign add_537954 = sel_537951 + 8'h01;
  assign sel_537955 = array_index_537774 == array_index_537286 ? add_537954 : sel_537951;
  assign add_537958 = sel_537955 + 8'h01;
  assign sel_537959 = array_index_537774 == array_index_537292 ? add_537958 : sel_537955;
  assign add_537962 = sel_537959 + 8'h01;
  assign sel_537963 = array_index_537774 == array_index_537298 ? add_537962 : sel_537959;
  assign add_537966 = sel_537963 + 8'h01;
  assign sel_537967 = array_index_537774 == array_index_537304 ? add_537966 : sel_537963;
  assign add_537970 = sel_537967 + 8'h01;
  assign sel_537971 = array_index_537774 == array_index_537310 ? add_537970 : sel_537967;
  assign add_537974 = sel_537971 + 8'h01;
  assign sel_537975 = array_index_537774 == array_index_537316 ? add_537974 : sel_537971;
  assign add_537978 = sel_537975 + 8'h01;
  assign sel_537979 = array_index_537774 == array_index_537322 ? add_537978 : sel_537975;
  assign add_537982 = sel_537979 + 8'h01;
  assign sel_537983 = array_index_537774 == array_index_537328 ? add_537982 : sel_537979;
  assign add_537986 = sel_537983 + 8'h01;
  assign sel_537987 = array_index_537774 == array_index_537334 ? add_537986 : sel_537983;
  assign add_537990 = sel_537987 + 8'h01;
  assign sel_537991 = array_index_537774 == array_index_537340 ? add_537990 : sel_537987;
  assign add_537994 = sel_537991 + 8'h01;
  assign sel_537995 = array_index_537774 == array_index_537346 ? add_537994 : sel_537991;
  assign add_537998 = sel_537995 + 8'h01;
  assign sel_537999 = array_index_537774 == array_index_537352 ? add_537998 : sel_537995;
  assign add_538002 = sel_537999 + 8'h01;
  assign sel_538003 = array_index_537774 == array_index_537358 ? add_538002 : sel_537999;
  assign add_538006 = sel_538003 + 8'h01;
  assign sel_538007 = array_index_537774 == array_index_537364 ? add_538006 : sel_538003;
  assign add_538010 = sel_538007 + 8'h01;
  assign sel_538011 = array_index_537774 == array_index_537370 ? add_538010 : sel_538007;
  assign add_538014 = sel_538011 + 8'h01;
  assign sel_538015 = array_index_537774 == array_index_537376 ? add_538014 : sel_538011;
  assign add_538018 = sel_538015 + 8'h01;
  assign sel_538019 = array_index_537774 == array_index_537382 ? add_538018 : sel_538015;
  assign add_538022 = sel_538019 + 8'h01;
  assign sel_538023 = array_index_537774 == array_index_537388 ? add_538022 : sel_538019;
  assign add_538026 = sel_538023 + 8'h01;
  assign sel_538027 = array_index_537774 == array_index_537394 ? add_538026 : sel_538023;
  assign add_538030 = sel_538027 + 8'h01;
  assign sel_538031 = array_index_537774 == array_index_537400 ? add_538030 : sel_538027;
  assign add_538034 = sel_538031 + 8'h01;
  assign sel_538035 = array_index_537774 == array_index_537406 ? add_538034 : sel_538031;
  assign add_538038 = sel_538035 + 8'h01;
  assign sel_538039 = array_index_537774 == array_index_537412 ? add_538038 : sel_538035;
  assign add_538042 = sel_538039 + 8'h01;
  assign sel_538043 = array_index_537774 == array_index_537418 ? add_538042 : sel_538039;
  assign add_538046 = sel_538043 + 8'h01;
  assign sel_538047 = array_index_537774 == array_index_537424 ? add_538046 : sel_538043;
  assign add_538050 = sel_538047 + 8'h01;
  assign sel_538051 = array_index_537774 == array_index_537430 ? add_538050 : sel_538047;
  assign add_538054 = sel_538051 + 8'h01;
  assign sel_538055 = array_index_537774 == array_index_537436 ? add_538054 : sel_538051;
  assign add_538058 = sel_538055 + 8'h01;
  assign sel_538059 = array_index_537774 == array_index_537442 ? add_538058 : sel_538055;
  assign add_538062 = sel_538059 + 8'h01;
  assign sel_538063 = array_index_537774 == array_index_537448 ? add_538062 : sel_538059;
  assign add_538066 = sel_538063 + 8'h01;
  assign sel_538067 = array_index_537774 == array_index_537454 ? add_538066 : sel_538063;
  assign add_538070 = sel_538067 + 8'h01;
  assign sel_538071 = array_index_537774 == array_index_537460 ? add_538070 : sel_538067;
  assign add_538075 = sel_538071 + 8'h01;
  assign array_index_538076 = set1_unflattened[7'h03];
  assign sel_538077 = array_index_537774 == array_index_537466 ? add_538075 : sel_538071;
  assign add_538080 = sel_538077 + 8'h01;
  assign sel_538081 = array_index_538076 == array_index_537012 ? add_538080 : sel_538077;
  assign add_538084 = sel_538081 + 8'h01;
  assign sel_538085 = array_index_538076 == array_index_537016 ? add_538084 : sel_538081;
  assign add_538088 = sel_538085 + 8'h01;
  assign sel_538089 = array_index_538076 == array_index_537024 ? add_538088 : sel_538085;
  assign add_538092 = sel_538089 + 8'h01;
  assign sel_538093 = array_index_538076 == array_index_537032 ? add_538092 : sel_538089;
  assign add_538096 = sel_538093 + 8'h01;
  assign sel_538097 = array_index_538076 == array_index_537040 ? add_538096 : sel_538093;
  assign add_538100 = sel_538097 + 8'h01;
  assign sel_538101 = array_index_538076 == array_index_537048 ? add_538100 : sel_538097;
  assign add_538104 = sel_538101 + 8'h01;
  assign sel_538105 = array_index_538076 == array_index_537056 ? add_538104 : sel_538101;
  assign add_538108 = sel_538105 + 8'h01;
  assign sel_538109 = array_index_538076 == array_index_537064 ? add_538108 : sel_538105;
  assign add_538112 = sel_538109 + 8'h01;
  assign sel_538113 = array_index_538076 == array_index_537070 ? add_538112 : sel_538109;
  assign add_538116 = sel_538113 + 8'h01;
  assign sel_538117 = array_index_538076 == array_index_537076 ? add_538116 : sel_538113;
  assign add_538120 = sel_538117 + 8'h01;
  assign sel_538121 = array_index_538076 == array_index_537082 ? add_538120 : sel_538117;
  assign add_538124 = sel_538121 + 8'h01;
  assign sel_538125 = array_index_538076 == array_index_537088 ? add_538124 : sel_538121;
  assign add_538128 = sel_538125 + 8'h01;
  assign sel_538129 = array_index_538076 == array_index_537094 ? add_538128 : sel_538125;
  assign add_538132 = sel_538129 + 8'h01;
  assign sel_538133 = array_index_538076 == array_index_537100 ? add_538132 : sel_538129;
  assign add_538136 = sel_538133 + 8'h01;
  assign sel_538137 = array_index_538076 == array_index_537106 ? add_538136 : sel_538133;
  assign add_538140 = sel_538137 + 8'h01;
  assign sel_538141 = array_index_538076 == array_index_537112 ? add_538140 : sel_538137;
  assign add_538144 = sel_538141 + 8'h01;
  assign sel_538145 = array_index_538076 == array_index_537118 ? add_538144 : sel_538141;
  assign add_538148 = sel_538145 + 8'h01;
  assign sel_538149 = array_index_538076 == array_index_537124 ? add_538148 : sel_538145;
  assign add_538152 = sel_538149 + 8'h01;
  assign sel_538153 = array_index_538076 == array_index_537130 ? add_538152 : sel_538149;
  assign add_538156 = sel_538153 + 8'h01;
  assign sel_538157 = array_index_538076 == array_index_537136 ? add_538156 : sel_538153;
  assign add_538160 = sel_538157 + 8'h01;
  assign sel_538161 = array_index_538076 == array_index_537142 ? add_538160 : sel_538157;
  assign add_538164 = sel_538161 + 8'h01;
  assign sel_538165 = array_index_538076 == array_index_537148 ? add_538164 : sel_538161;
  assign add_538168 = sel_538165 + 8'h01;
  assign sel_538169 = array_index_538076 == array_index_537154 ? add_538168 : sel_538165;
  assign add_538172 = sel_538169 + 8'h01;
  assign sel_538173 = array_index_538076 == array_index_537160 ? add_538172 : sel_538169;
  assign add_538176 = sel_538173 + 8'h01;
  assign sel_538177 = array_index_538076 == array_index_537166 ? add_538176 : sel_538173;
  assign add_538180 = sel_538177 + 8'h01;
  assign sel_538181 = array_index_538076 == array_index_537172 ? add_538180 : sel_538177;
  assign add_538184 = sel_538181 + 8'h01;
  assign sel_538185 = array_index_538076 == array_index_537178 ? add_538184 : sel_538181;
  assign add_538188 = sel_538185 + 8'h01;
  assign sel_538189 = array_index_538076 == array_index_537184 ? add_538188 : sel_538185;
  assign add_538192 = sel_538189 + 8'h01;
  assign sel_538193 = array_index_538076 == array_index_537190 ? add_538192 : sel_538189;
  assign add_538196 = sel_538193 + 8'h01;
  assign sel_538197 = array_index_538076 == array_index_537196 ? add_538196 : sel_538193;
  assign add_538200 = sel_538197 + 8'h01;
  assign sel_538201 = array_index_538076 == array_index_537202 ? add_538200 : sel_538197;
  assign add_538204 = sel_538201 + 8'h01;
  assign sel_538205 = array_index_538076 == array_index_537208 ? add_538204 : sel_538201;
  assign add_538208 = sel_538205 + 8'h01;
  assign sel_538209 = array_index_538076 == array_index_537214 ? add_538208 : sel_538205;
  assign add_538212 = sel_538209 + 8'h01;
  assign sel_538213 = array_index_538076 == array_index_537220 ? add_538212 : sel_538209;
  assign add_538216 = sel_538213 + 8'h01;
  assign sel_538217 = array_index_538076 == array_index_537226 ? add_538216 : sel_538213;
  assign add_538220 = sel_538217 + 8'h01;
  assign sel_538221 = array_index_538076 == array_index_537232 ? add_538220 : sel_538217;
  assign add_538224 = sel_538221 + 8'h01;
  assign sel_538225 = array_index_538076 == array_index_537238 ? add_538224 : sel_538221;
  assign add_538228 = sel_538225 + 8'h01;
  assign sel_538229 = array_index_538076 == array_index_537244 ? add_538228 : sel_538225;
  assign add_538232 = sel_538229 + 8'h01;
  assign sel_538233 = array_index_538076 == array_index_537250 ? add_538232 : sel_538229;
  assign add_538236 = sel_538233 + 8'h01;
  assign sel_538237 = array_index_538076 == array_index_537256 ? add_538236 : sel_538233;
  assign add_538240 = sel_538237 + 8'h01;
  assign sel_538241 = array_index_538076 == array_index_537262 ? add_538240 : sel_538237;
  assign add_538244 = sel_538241 + 8'h01;
  assign sel_538245 = array_index_538076 == array_index_537268 ? add_538244 : sel_538241;
  assign add_538248 = sel_538245 + 8'h01;
  assign sel_538249 = array_index_538076 == array_index_537274 ? add_538248 : sel_538245;
  assign add_538252 = sel_538249 + 8'h01;
  assign sel_538253 = array_index_538076 == array_index_537280 ? add_538252 : sel_538249;
  assign add_538256 = sel_538253 + 8'h01;
  assign sel_538257 = array_index_538076 == array_index_537286 ? add_538256 : sel_538253;
  assign add_538260 = sel_538257 + 8'h01;
  assign sel_538261 = array_index_538076 == array_index_537292 ? add_538260 : sel_538257;
  assign add_538264 = sel_538261 + 8'h01;
  assign sel_538265 = array_index_538076 == array_index_537298 ? add_538264 : sel_538261;
  assign add_538268 = sel_538265 + 8'h01;
  assign sel_538269 = array_index_538076 == array_index_537304 ? add_538268 : sel_538265;
  assign add_538272 = sel_538269 + 8'h01;
  assign sel_538273 = array_index_538076 == array_index_537310 ? add_538272 : sel_538269;
  assign add_538276 = sel_538273 + 8'h01;
  assign sel_538277 = array_index_538076 == array_index_537316 ? add_538276 : sel_538273;
  assign add_538280 = sel_538277 + 8'h01;
  assign sel_538281 = array_index_538076 == array_index_537322 ? add_538280 : sel_538277;
  assign add_538284 = sel_538281 + 8'h01;
  assign sel_538285 = array_index_538076 == array_index_537328 ? add_538284 : sel_538281;
  assign add_538288 = sel_538285 + 8'h01;
  assign sel_538289 = array_index_538076 == array_index_537334 ? add_538288 : sel_538285;
  assign add_538292 = sel_538289 + 8'h01;
  assign sel_538293 = array_index_538076 == array_index_537340 ? add_538292 : sel_538289;
  assign add_538296 = sel_538293 + 8'h01;
  assign sel_538297 = array_index_538076 == array_index_537346 ? add_538296 : sel_538293;
  assign add_538300 = sel_538297 + 8'h01;
  assign sel_538301 = array_index_538076 == array_index_537352 ? add_538300 : sel_538297;
  assign add_538304 = sel_538301 + 8'h01;
  assign sel_538305 = array_index_538076 == array_index_537358 ? add_538304 : sel_538301;
  assign add_538308 = sel_538305 + 8'h01;
  assign sel_538309 = array_index_538076 == array_index_537364 ? add_538308 : sel_538305;
  assign add_538312 = sel_538309 + 8'h01;
  assign sel_538313 = array_index_538076 == array_index_537370 ? add_538312 : sel_538309;
  assign add_538316 = sel_538313 + 8'h01;
  assign sel_538317 = array_index_538076 == array_index_537376 ? add_538316 : sel_538313;
  assign add_538320 = sel_538317 + 8'h01;
  assign sel_538321 = array_index_538076 == array_index_537382 ? add_538320 : sel_538317;
  assign add_538324 = sel_538321 + 8'h01;
  assign sel_538325 = array_index_538076 == array_index_537388 ? add_538324 : sel_538321;
  assign add_538328 = sel_538325 + 8'h01;
  assign sel_538329 = array_index_538076 == array_index_537394 ? add_538328 : sel_538325;
  assign add_538332 = sel_538329 + 8'h01;
  assign sel_538333 = array_index_538076 == array_index_537400 ? add_538332 : sel_538329;
  assign add_538336 = sel_538333 + 8'h01;
  assign sel_538337 = array_index_538076 == array_index_537406 ? add_538336 : sel_538333;
  assign add_538340 = sel_538337 + 8'h01;
  assign sel_538341 = array_index_538076 == array_index_537412 ? add_538340 : sel_538337;
  assign add_538344 = sel_538341 + 8'h01;
  assign sel_538345 = array_index_538076 == array_index_537418 ? add_538344 : sel_538341;
  assign add_538348 = sel_538345 + 8'h01;
  assign sel_538349 = array_index_538076 == array_index_537424 ? add_538348 : sel_538345;
  assign add_538352 = sel_538349 + 8'h01;
  assign sel_538353 = array_index_538076 == array_index_537430 ? add_538352 : sel_538349;
  assign add_538356 = sel_538353 + 8'h01;
  assign sel_538357 = array_index_538076 == array_index_537436 ? add_538356 : sel_538353;
  assign add_538360 = sel_538357 + 8'h01;
  assign sel_538361 = array_index_538076 == array_index_537442 ? add_538360 : sel_538357;
  assign add_538364 = sel_538361 + 8'h01;
  assign sel_538365 = array_index_538076 == array_index_537448 ? add_538364 : sel_538361;
  assign add_538368 = sel_538365 + 8'h01;
  assign sel_538369 = array_index_538076 == array_index_537454 ? add_538368 : sel_538365;
  assign add_538372 = sel_538369 + 8'h01;
  assign sel_538373 = array_index_538076 == array_index_537460 ? add_538372 : sel_538369;
  assign add_538377 = sel_538373 + 8'h01;
  assign array_index_538378 = set1_unflattened[7'h04];
  assign sel_538379 = array_index_538076 == array_index_537466 ? add_538377 : sel_538373;
  assign add_538382 = sel_538379 + 8'h01;
  assign sel_538383 = array_index_538378 == array_index_537012 ? add_538382 : sel_538379;
  assign add_538386 = sel_538383 + 8'h01;
  assign sel_538387 = array_index_538378 == array_index_537016 ? add_538386 : sel_538383;
  assign add_538390 = sel_538387 + 8'h01;
  assign sel_538391 = array_index_538378 == array_index_537024 ? add_538390 : sel_538387;
  assign add_538394 = sel_538391 + 8'h01;
  assign sel_538395 = array_index_538378 == array_index_537032 ? add_538394 : sel_538391;
  assign add_538398 = sel_538395 + 8'h01;
  assign sel_538399 = array_index_538378 == array_index_537040 ? add_538398 : sel_538395;
  assign add_538402 = sel_538399 + 8'h01;
  assign sel_538403 = array_index_538378 == array_index_537048 ? add_538402 : sel_538399;
  assign add_538406 = sel_538403 + 8'h01;
  assign sel_538407 = array_index_538378 == array_index_537056 ? add_538406 : sel_538403;
  assign add_538410 = sel_538407 + 8'h01;
  assign sel_538411 = array_index_538378 == array_index_537064 ? add_538410 : sel_538407;
  assign add_538414 = sel_538411 + 8'h01;
  assign sel_538415 = array_index_538378 == array_index_537070 ? add_538414 : sel_538411;
  assign add_538418 = sel_538415 + 8'h01;
  assign sel_538419 = array_index_538378 == array_index_537076 ? add_538418 : sel_538415;
  assign add_538422 = sel_538419 + 8'h01;
  assign sel_538423 = array_index_538378 == array_index_537082 ? add_538422 : sel_538419;
  assign add_538426 = sel_538423 + 8'h01;
  assign sel_538427 = array_index_538378 == array_index_537088 ? add_538426 : sel_538423;
  assign add_538430 = sel_538427 + 8'h01;
  assign sel_538431 = array_index_538378 == array_index_537094 ? add_538430 : sel_538427;
  assign add_538434 = sel_538431 + 8'h01;
  assign sel_538435 = array_index_538378 == array_index_537100 ? add_538434 : sel_538431;
  assign add_538438 = sel_538435 + 8'h01;
  assign sel_538439 = array_index_538378 == array_index_537106 ? add_538438 : sel_538435;
  assign add_538442 = sel_538439 + 8'h01;
  assign sel_538443 = array_index_538378 == array_index_537112 ? add_538442 : sel_538439;
  assign add_538446 = sel_538443 + 8'h01;
  assign sel_538447 = array_index_538378 == array_index_537118 ? add_538446 : sel_538443;
  assign add_538450 = sel_538447 + 8'h01;
  assign sel_538451 = array_index_538378 == array_index_537124 ? add_538450 : sel_538447;
  assign add_538454 = sel_538451 + 8'h01;
  assign sel_538455 = array_index_538378 == array_index_537130 ? add_538454 : sel_538451;
  assign add_538458 = sel_538455 + 8'h01;
  assign sel_538459 = array_index_538378 == array_index_537136 ? add_538458 : sel_538455;
  assign add_538462 = sel_538459 + 8'h01;
  assign sel_538463 = array_index_538378 == array_index_537142 ? add_538462 : sel_538459;
  assign add_538466 = sel_538463 + 8'h01;
  assign sel_538467 = array_index_538378 == array_index_537148 ? add_538466 : sel_538463;
  assign add_538470 = sel_538467 + 8'h01;
  assign sel_538471 = array_index_538378 == array_index_537154 ? add_538470 : sel_538467;
  assign add_538474 = sel_538471 + 8'h01;
  assign sel_538475 = array_index_538378 == array_index_537160 ? add_538474 : sel_538471;
  assign add_538478 = sel_538475 + 8'h01;
  assign sel_538479 = array_index_538378 == array_index_537166 ? add_538478 : sel_538475;
  assign add_538482 = sel_538479 + 8'h01;
  assign sel_538483 = array_index_538378 == array_index_537172 ? add_538482 : sel_538479;
  assign add_538486 = sel_538483 + 8'h01;
  assign sel_538487 = array_index_538378 == array_index_537178 ? add_538486 : sel_538483;
  assign add_538490 = sel_538487 + 8'h01;
  assign sel_538491 = array_index_538378 == array_index_537184 ? add_538490 : sel_538487;
  assign add_538494 = sel_538491 + 8'h01;
  assign sel_538495 = array_index_538378 == array_index_537190 ? add_538494 : sel_538491;
  assign add_538498 = sel_538495 + 8'h01;
  assign sel_538499 = array_index_538378 == array_index_537196 ? add_538498 : sel_538495;
  assign add_538502 = sel_538499 + 8'h01;
  assign sel_538503 = array_index_538378 == array_index_537202 ? add_538502 : sel_538499;
  assign add_538506 = sel_538503 + 8'h01;
  assign sel_538507 = array_index_538378 == array_index_537208 ? add_538506 : sel_538503;
  assign add_538510 = sel_538507 + 8'h01;
  assign sel_538511 = array_index_538378 == array_index_537214 ? add_538510 : sel_538507;
  assign add_538514 = sel_538511 + 8'h01;
  assign sel_538515 = array_index_538378 == array_index_537220 ? add_538514 : sel_538511;
  assign add_538518 = sel_538515 + 8'h01;
  assign sel_538519 = array_index_538378 == array_index_537226 ? add_538518 : sel_538515;
  assign add_538522 = sel_538519 + 8'h01;
  assign sel_538523 = array_index_538378 == array_index_537232 ? add_538522 : sel_538519;
  assign add_538526 = sel_538523 + 8'h01;
  assign sel_538527 = array_index_538378 == array_index_537238 ? add_538526 : sel_538523;
  assign add_538530 = sel_538527 + 8'h01;
  assign sel_538531 = array_index_538378 == array_index_537244 ? add_538530 : sel_538527;
  assign add_538534 = sel_538531 + 8'h01;
  assign sel_538535 = array_index_538378 == array_index_537250 ? add_538534 : sel_538531;
  assign add_538538 = sel_538535 + 8'h01;
  assign sel_538539 = array_index_538378 == array_index_537256 ? add_538538 : sel_538535;
  assign add_538542 = sel_538539 + 8'h01;
  assign sel_538543 = array_index_538378 == array_index_537262 ? add_538542 : sel_538539;
  assign add_538546 = sel_538543 + 8'h01;
  assign sel_538547 = array_index_538378 == array_index_537268 ? add_538546 : sel_538543;
  assign add_538550 = sel_538547 + 8'h01;
  assign sel_538551 = array_index_538378 == array_index_537274 ? add_538550 : sel_538547;
  assign add_538554 = sel_538551 + 8'h01;
  assign sel_538555 = array_index_538378 == array_index_537280 ? add_538554 : sel_538551;
  assign add_538558 = sel_538555 + 8'h01;
  assign sel_538559 = array_index_538378 == array_index_537286 ? add_538558 : sel_538555;
  assign add_538562 = sel_538559 + 8'h01;
  assign sel_538563 = array_index_538378 == array_index_537292 ? add_538562 : sel_538559;
  assign add_538566 = sel_538563 + 8'h01;
  assign sel_538567 = array_index_538378 == array_index_537298 ? add_538566 : sel_538563;
  assign add_538570 = sel_538567 + 8'h01;
  assign sel_538571 = array_index_538378 == array_index_537304 ? add_538570 : sel_538567;
  assign add_538574 = sel_538571 + 8'h01;
  assign sel_538575 = array_index_538378 == array_index_537310 ? add_538574 : sel_538571;
  assign add_538578 = sel_538575 + 8'h01;
  assign sel_538579 = array_index_538378 == array_index_537316 ? add_538578 : sel_538575;
  assign add_538582 = sel_538579 + 8'h01;
  assign sel_538583 = array_index_538378 == array_index_537322 ? add_538582 : sel_538579;
  assign add_538586 = sel_538583 + 8'h01;
  assign sel_538587 = array_index_538378 == array_index_537328 ? add_538586 : sel_538583;
  assign add_538590 = sel_538587 + 8'h01;
  assign sel_538591 = array_index_538378 == array_index_537334 ? add_538590 : sel_538587;
  assign add_538594 = sel_538591 + 8'h01;
  assign sel_538595 = array_index_538378 == array_index_537340 ? add_538594 : sel_538591;
  assign add_538598 = sel_538595 + 8'h01;
  assign sel_538599 = array_index_538378 == array_index_537346 ? add_538598 : sel_538595;
  assign add_538602 = sel_538599 + 8'h01;
  assign sel_538603 = array_index_538378 == array_index_537352 ? add_538602 : sel_538599;
  assign add_538606 = sel_538603 + 8'h01;
  assign sel_538607 = array_index_538378 == array_index_537358 ? add_538606 : sel_538603;
  assign add_538610 = sel_538607 + 8'h01;
  assign sel_538611 = array_index_538378 == array_index_537364 ? add_538610 : sel_538607;
  assign add_538614 = sel_538611 + 8'h01;
  assign sel_538615 = array_index_538378 == array_index_537370 ? add_538614 : sel_538611;
  assign add_538618 = sel_538615 + 8'h01;
  assign sel_538619 = array_index_538378 == array_index_537376 ? add_538618 : sel_538615;
  assign add_538622 = sel_538619 + 8'h01;
  assign sel_538623 = array_index_538378 == array_index_537382 ? add_538622 : sel_538619;
  assign add_538626 = sel_538623 + 8'h01;
  assign sel_538627 = array_index_538378 == array_index_537388 ? add_538626 : sel_538623;
  assign add_538630 = sel_538627 + 8'h01;
  assign sel_538631 = array_index_538378 == array_index_537394 ? add_538630 : sel_538627;
  assign add_538634 = sel_538631 + 8'h01;
  assign sel_538635 = array_index_538378 == array_index_537400 ? add_538634 : sel_538631;
  assign add_538638 = sel_538635 + 8'h01;
  assign sel_538639 = array_index_538378 == array_index_537406 ? add_538638 : sel_538635;
  assign add_538642 = sel_538639 + 8'h01;
  assign sel_538643 = array_index_538378 == array_index_537412 ? add_538642 : sel_538639;
  assign add_538646 = sel_538643 + 8'h01;
  assign sel_538647 = array_index_538378 == array_index_537418 ? add_538646 : sel_538643;
  assign add_538650 = sel_538647 + 8'h01;
  assign sel_538651 = array_index_538378 == array_index_537424 ? add_538650 : sel_538647;
  assign add_538654 = sel_538651 + 8'h01;
  assign sel_538655 = array_index_538378 == array_index_537430 ? add_538654 : sel_538651;
  assign add_538658 = sel_538655 + 8'h01;
  assign sel_538659 = array_index_538378 == array_index_537436 ? add_538658 : sel_538655;
  assign add_538662 = sel_538659 + 8'h01;
  assign sel_538663 = array_index_538378 == array_index_537442 ? add_538662 : sel_538659;
  assign add_538666 = sel_538663 + 8'h01;
  assign sel_538667 = array_index_538378 == array_index_537448 ? add_538666 : sel_538663;
  assign add_538670 = sel_538667 + 8'h01;
  assign sel_538671 = array_index_538378 == array_index_537454 ? add_538670 : sel_538667;
  assign add_538674 = sel_538671 + 8'h01;
  assign sel_538675 = array_index_538378 == array_index_537460 ? add_538674 : sel_538671;
  assign add_538679 = sel_538675 + 8'h01;
  assign array_index_538680 = set1_unflattened[7'h05];
  assign sel_538681 = array_index_538378 == array_index_537466 ? add_538679 : sel_538675;
  assign add_538684 = sel_538681 + 8'h01;
  assign sel_538685 = array_index_538680 == array_index_537012 ? add_538684 : sel_538681;
  assign add_538688 = sel_538685 + 8'h01;
  assign sel_538689 = array_index_538680 == array_index_537016 ? add_538688 : sel_538685;
  assign add_538692 = sel_538689 + 8'h01;
  assign sel_538693 = array_index_538680 == array_index_537024 ? add_538692 : sel_538689;
  assign add_538696 = sel_538693 + 8'h01;
  assign sel_538697 = array_index_538680 == array_index_537032 ? add_538696 : sel_538693;
  assign add_538700 = sel_538697 + 8'h01;
  assign sel_538701 = array_index_538680 == array_index_537040 ? add_538700 : sel_538697;
  assign add_538704 = sel_538701 + 8'h01;
  assign sel_538705 = array_index_538680 == array_index_537048 ? add_538704 : sel_538701;
  assign add_538708 = sel_538705 + 8'h01;
  assign sel_538709 = array_index_538680 == array_index_537056 ? add_538708 : sel_538705;
  assign add_538712 = sel_538709 + 8'h01;
  assign sel_538713 = array_index_538680 == array_index_537064 ? add_538712 : sel_538709;
  assign add_538716 = sel_538713 + 8'h01;
  assign sel_538717 = array_index_538680 == array_index_537070 ? add_538716 : sel_538713;
  assign add_538720 = sel_538717 + 8'h01;
  assign sel_538721 = array_index_538680 == array_index_537076 ? add_538720 : sel_538717;
  assign add_538724 = sel_538721 + 8'h01;
  assign sel_538725 = array_index_538680 == array_index_537082 ? add_538724 : sel_538721;
  assign add_538728 = sel_538725 + 8'h01;
  assign sel_538729 = array_index_538680 == array_index_537088 ? add_538728 : sel_538725;
  assign add_538732 = sel_538729 + 8'h01;
  assign sel_538733 = array_index_538680 == array_index_537094 ? add_538732 : sel_538729;
  assign add_538736 = sel_538733 + 8'h01;
  assign sel_538737 = array_index_538680 == array_index_537100 ? add_538736 : sel_538733;
  assign add_538740 = sel_538737 + 8'h01;
  assign sel_538741 = array_index_538680 == array_index_537106 ? add_538740 : sel_538737;
  assign add_538744 = sel_538741 + 8'h01;
  assign sel_538745 = array_index_538680 == array_index_537112 ? add_538744 : sel_538741;
  assign add_538748 = sel_538745 + 8'h01;
  assign sel_538749 = array_index_538680 == array_index_537118 ? add_538748 : sel_538745;
  assign add_538752 = sel_538749 + 8'h01;
  assign sel_538753 = array_index_538680 == array_index_537124 ? add_538752 : sel_538749;
  assign add_538756 = sel_538753 + 8'h01;
  assign sel_538757 = array_index_538680 == array_index_537130 ? add_538756 : sel_538753;
  assign add_538760 = sel_538757 + 8'h01;
  assign sel_538761 = array_index_538680 == array_index_537136 ? add_538760 : sel_538757;
  assign add_538764 = sel_538761 + 8'h01;
  assign sel_538765 = array_index_538680 == array_index_537142 ? add_538764 : sel_538761;
  assign add_538768 = sel_538765 + 8'h01;
  assign sel_538769 = array_index_538680 == array_index_537148 ? add_538768 : sel_538765;
  assign add_538772 = sel_538769 + 8'h01;
  assign sel_538773 = array_index_538680 == array_index_537154 ? add_538772 : sel_538769;
  assign add_538776 = sel_538773 + 8'h01;
  assign sel_538777 = array_index_538680 == array_index_537160 ? add_538776 : sel_538773;
  assign add_538780 = sel_538777 + 8'h01;
  assign sel_538781 = array_index_538680 == array_index_537166 ? add_538780 : sel_538777;
  assign add_538784 = sel_538781 + 8'h01;
  assign sel_538785 = array_index_538680 == array_index_537172 ? add_538784 : sel_538781;
  assign add_538788 = sel_538785 + 8'h01;
  assign sel_538789 = array_index_538680 == array_index_537178 ? add_538788 : sel_538785;
  assign add_538792 = sel_538789 + 8'h01;
  assign sel_538793 = array_index_538680 == array_index_537184 ? add_538792 : sel_538789;
  assign add_538796 = sel_538793 + 8'h01;
  assign sel_538797 = array_index_538680 == array_index_537190 ? add_538796 : sel_538793;
  assign add_538800 = sel_538797 + 8'h01;
  assign sel_538801 = array_index_538680 == array_index_537196 ? add_538800 : sel_538797;
  assign add_538804 = sel_538801 + 8'h01;
  assign sel_538805 = array_index_538680 == array_index_537202 ? add_538804 : sel_538801;
  assign add_538808 = sel_538805 + 8'h01;
  assign sel_538809 = array_index_538680 == array_index_537208 ? add_538808 : sel_538805;
  assign add_538812 = sel_538809 + 8'h01;
  assign sel_538813 = array_index_538680 == array_index_537214 ? add_538812 : sel_538809;
  assign add_538816 = sel_538813 + 8'h01;
  assign sel_538817 = array_index_538680 == array_index_537220 ? add_538816 : sel_538813;
  assign add_538820 = sel_538817 + 8'h01;
  assign sel_538821 = array_index_538680 == array_index_537226 ? add_538820 : sel_538817;
  assign add_538824 = sel_538821 + 8'h01;
  assign sel_538825 = array_index_538680 == array_index_537232 ? add_538824 : sel_538821;
  assign add_538828 = sel_538825 + 8'h01;
  assign sel_538829 = array_index_538680 == array_index_537238 ? add_538828 : sel_538825;
  assign add_538832 = sel_538829 + 8'h01;
  assign sel_538833 = array_index_538680 == array_index_537244 ? add_538832 : sel_538829;
  assign add_538836 = sel_538833 + 8'h01;
  assign sel_538837 = array_index_538680 == array_index_537250 ? add_538836 : sel_538833;
  assign add_538840 = sel_538837 + 8'h01;
  assign sel_538841 = array_index_538680 == array_index_537256 ? add_538840 : sel_538837;
  assign add_538844 = sel_538841 + 8'h01;
  assign sel_538845 = array_index_538680 == array_index_537262 ? add_538844 : sel_538841;
  assign add_538848 = sel_538845 + 8'h01;
  assign sel_538849 = array_index_538680 == array_index_537268 ? add_538848 : sel_538845;
  assign add_538852 = sel_538849 + 8'h01;
  assign sel_538853 = array_index_538680 == array_index_537274 ? add_538852 : sel_538849;
  assign add_538856 = sel_538853 + 8'h01;
  assign sel_538857 = array_index_538680 == array_index_537280 ? add_538856 : sel_538853;
  assign add_538860 = sel_538857 + 8'h01;
  assign sel_538861 = array_index_538680 == array_index_537286 ? add_538860 : sel_538857;
  assign add_538864 = sel_538861 + 8'h01;
  assign sel_538865 = array_index_538680 == array_index_537292 ? add_538864 : sel_538861;
  assign add_538868 = sel_538865 + 8'h01;
  assign sel_538869 = array_index_538680 == array_index_537298 ? add_538868 : sel_538865;
  assign add_538872 = sel_538869 + 8'h01;
  assign sel_538873 = array_index_538680 == array_index_537304 ? add_538872 : sel_538869;
  assign add_538876 = sel_538873 + 8'h01;
  assign sel_538877 = array_index_538680 == array_index_537310 ? add_538876 : sel_538873;
  assign add_538880 = sel_538877 + 8'h01;
  assign sel_538881 = array_index_538680 == array_index_537316 ? add_538880 : sel_538877;
  assign add_538884 = sel_538881 + 8'h01;
  assign sel_538885 = array_index_538680 == array_index_537322 ? add_538884 : sel_538881;
  assign add_538888 = sel_538885 + 8'h01;
  assign sel_538889 = array_index_538680 == array_index_537328 ? add_538888 : sel_538885;
  assign add_538892 = sel_538889 + 8'h01;
  assign sel_538893 = array_index_538680 == array_index_537334 ? add_538892 : sel_538889;
  assign add_538896 = sel_538893 + 8'h01;
  assign sel_538897 = array_index_538680 == array_index_537340 ? add_538896 : sel_538893;
  assign add_538900 = sel_538897 + 8'h01;
  assign sel_538901 = array_index_538680 == array_index_537346 ? add_538900 : sel_538897;
  assign add_538904 = sel_538901 + 8'h01;
  assign sel_538905 = array_index_538680 == array_index_537352 ? add_538904 : sel_538901;
  assign add_538908 = sel_538905 + 8'h01;
  assign sel_538909 = array_index_538680 == array_index_537358 ? add_538908 : sel_538905;
  assign add_538912 = sel_538909 + 8'h01;
  assign sel_538913 = array_index_538680 == array_index_537364 ? add_538912 : sel_538909;
  assign add_538916 = sel_538913 + 8'h01;
  assign sel_538917 = array_index_538680 == array_index_537370 ? add_538916 : sel_538913;
  assign add_538920 = sel_538917 + 8'h01;
  assign sel_538921 = array_index_538680 == array_index_537376 ? add_538920 : sel_538917;
  assign add_538924 = sel_538921 + 8'h01;
  assign sel_538925 = array_index_538680 == array_index_537382 ? add_538924 : sel_538921;
  assign add_538928 = sel_538925 + 8'h01;
  assign sel_538929 = array_index_538680 == array_index_537388 ? add_538928 : sel_538925;
  assign add_538932 = sel_538929 + 8'h01;
  assign sel_538933 = array_index_538680 == array_index_537394 ? add_538932 : sel_538929;
  assign add_538936 = sel_538933 + 8'h01;
  assign sel_538937 = array_index_538680 == array_index_537400 ? add_538936 : sel_538933;
  assign add_538940 = sel_538937 + 8'h01;
  assign sel_538941 = array_index_538680 == array_index_537406 ? add_538940 : sel_538937;
  assign add_538944 = sel_538941 + 8'h01;
  assign sel_538945 = array_index_538680 == array_index_537412 ? add_538944 : sel_538941;
  assign add_538948 = sel_538945 + 8'h01;
  assign sel_538949 = array_index_538680 == array_index_537418 ? add_538948 : sel_538945;
  assign add_538952 = sel_538949 + 8'h01;
  assign sel_538953 = array_index_538680 == array_index_537424 ? add_538952 : sel_538949;
  assign add_538956 = sel_538953 + 8'h01;
  assign sel_538957 = array_index_538680 == array_index_537430 ? add_538956 : sel_538953;
  assign add_538960 = sel_538957 + 8'h01;
  assign sel_538961 = array_index_538680 == array_index_537436 ? add_538960 : sel_538957;
  assign add_538964 = sel_538961 + 8'h01;
  assign sel_538965 = array_index_538680 == array_index_537442 ? add_538964 : sel_538961;
  assign add_538968 = sel_538965 + 8'h01;
  assign sel_538969 = array_index_538680 == array_index_537448 ? add_538968 : sel_538965;
  assign add_538972 = sel_538969 + 8'h01;
  assign sel_538973 = array_index_538680 == array_index_537454 ? add_538972 : sel_538969;
  assign add_538976 = sel_538973 + 8'h01;
  assign sel_538977 = array_index_538680 == array_index_537460 ? add_538976 : sel_538973;
  assign add_538981 = sel_538977 + 8'h01;
  assign array_index_538982 = set1_unflattened[7'h06];
  assign sel_538983 = array_index_538680 == array_index_537466 ? add_538981 : sel_538977;
  assign add_538986 = sel_538983 + 8'h01;
  assign sel_538987 = array_index_538982 == array_index_537012 ? add_538986 : sel_538983;
  assign add_538990 = sel_538987 + 8'h01;
  assign sel_538991 = array_index_538982 == array_index_537016 ? add_538990 : sel_538987;
  assign add_538994 = sel_538991 + 8'h01;
  assign sel_538995 = array_index_538982 == array_index_537024 ? add_538994 : sel_538991;
  assign add_538998 = sel_538995 + 8'h01;
  assign sel_538999 = array_index_538982 == array_index_537032 ? add_538998 : sel_538995;
  assign add_539002 = sel_538999 + 8'h01;
  assign sel_539003 = array_index_538982 == array_index_537040 ? add_539002 : sel_538999;
  assign add_539006 = sel_539003 + 8'h01;
  assign sel_539007 = array_index_538982 == array_index_537048 ? add_539006 : sel_539003;
  assign add_539010 = sel_539007 + 8'h01;
  assign sel_539011 = array_index_538982 == array_index_537056 ? add_539010 : sel_539007;
  assign add_539014 = sel_539011 + 8'h01;
  assign sel_539015 = array_index_538982 == array_index_537064 ? add_539014 : sel_539011;
  assign add_539018 = sel_539015 + 8'h01;
  assign sel_539019 = array_index_538982 == array_index_537070 ? add_539018 : sel_539015;
  assign add_539022 = sel_539019 + 8'h01;
  assign sel_539023 = array_index_538982 == array_index_537076 ? add_539022 : sel_539019;
  assign add_539026 = sel_539023 + 8'h01;
  assign sel_539027 = array_index_538982 == array_index_537082 ? add_539026 : sel_539023;
  assign add_539030 = sel_539027 + 8'h01;
  assign sel_539031 = array_index_538982 == array_index_537088 ? add_539030 : sel_539027;
  assign add_539034 = sel_539031 + 8'h01;
  assign sel_539035 = array_index_538982 == array_index_537094 ? add_539034 : sel_539031;
  assign add_539038 = sel_539035 + 8'h01;
  assign sel_539039 = array_index_538982 == array_index_537100 ? add_539038 : sel_539035;
  assign add_539042 = sel_539039 + 8'h01;
  assign sel_539043 = array_index_538982 == array_index_537106 ? add_539042 : sel_539039;
  assign add_539046 = sel_539043 + 8'h01;
  assign sel_539047 = array_index_538982 == array_index_537112 ? add_539046 : sel_539043;
  assign add_539050 = sel_539047 + 8'h01;
  assign sel_539051 = array_index_538982 == array_index_537118 ? add_539050 : sel_539047;
  assign add_539054 = sel_539051 + 8'h01;
  assign sel_539055 = array_index_538982 == array_index_537124 ? add_539054 : sel_539051;
  assign add_539058 = sel_539055 + 8'h01;
  assign sel_539059 = array_index_538982 == array_index_537130 ? add_539058 : sel_539055;
  assign add_539062 = sel_539059 + 8'h01;
  assign sel_539063 = array_index_538982 == array_index_537136 ? add_539062 : sel_539059;
  assign add_539066 = sel_539063 + 8'h01;
  assign sel_539067 = array_index_538982 == array_index_537142 ? add_539066 : sel_539063;
  assign add_539070 = sel_539067 + 8'h01;
  assign sel_539071 = array_index_538982 == array_index_537148 ? add_539070 : sel_539067;
  assign add_539074 = sel_539071 + 8'h01;
  assign sel_539075 = array_index_538982 == array_index_537154 ? add_539074 : sel_539071;
  assign add_539078 = sel_539075 + 8'h01;
  assign sel_539079 = array_index_538982 == array_index_537160 ? add_539078 : sel_539075;
  assign add_539082 = sel_539079 + 8'h01;
  assign sel_539083 = array_index_538982 == array_index_537166 ? add_539082 : sel_539079;
  assign add_539086 = sel_539083 + 8'h01;
  assign sel_539087 = array_index_538982 == array_index_537172 ? add_539086 : sel_539083;
  assign add_539090 = sel_539087 + 8'h01;
  assign sel_539091 = array_index_538982 == array_index_537178 ? add_539090 : sel_539087;
  assign add_539094 = sel_539091 + 8'h01;
  assign sel_539095 = array_index_538982 == array_index_537184 ? add_539094 : sel_539091;
  assign add_539098 = sel_539095 + 8'h01;
  assign sel_539099 = array_index_538982 == array_index_537190 ? add_539098 : sel_539095;
  assign add_539102 = sel_539099 + 8'h01;
  assign sel_539103 = array_index_538982 == array_index_537196 ? add_539102 : sel_539099;
  assign add_539106 = sel_539103 + 8'h01;
  assign sel_539107 = array_index_538982 == array_index_537202 ? add_539106 : sel_539103;
  assign add_539110 = sel_539107 + 8'h01;
  assign sel_539111 = array_index_538982 == array_index_537208 ? add_539110 : sel_539107;
  assign add_539114 = sel_539111 + 8'h01;
  assign sel_539115 = array_index_538982 == array_index_537214 ? add_539114 : sel_539111;
  assign add_539118 = sel_539115 + 8'h01;
  assign sel_539119 = array_index_538982 == array_index_537220 ? add_539118 : sel_539115;
  assign add_539122 = sel_539119 + 8'h01;
  assign sel_539123 = array_index_538982 == array_index_537226 ? add_539122 : sel_539119;
  assign add_539126 = sel_539123 + 8'h01;
  assign sel_539127 = array_index_538982 == array_index_537232 ? add_539126 : sel_539123;
  assign add_539130 = sel_539127 + 8'h01;
  assign sel_539131 = array_index_538982 == array_index_537238 ? add_539130 : sel_539127;
  assign add_539134 = sel_539131 + 8'h01;
  assign sel_539135 = array_index_538982 == array_index_537244 ? add_539134 : sel_539131;
  assign add_539138 = sel_539135 + 8'h01;
  assign sel_539139 = array_index_538982 == array_index_537250 ? add_539138 : sel_539135;
  assign add_539142 = sel_539139 + 8'h01;
  assign sel_539143 = array_index_538982 == array_index_537256 ? add_539142 : sel_539139;
  assign add_539146 = sel_539143 + 8'h01;
  assign sel_539147 = array_index_538982 == array_index_537262 ? add_539146 : sel_539143;
  assign add_539150 = sel_539147 + 8'h01;
  assign sel_539151 = array_index_538982 == array_index_537268 ? add_539150 : sel_539147;
  assign add_539154 = sel_539151 + 8'h01;
  assign sel_539155 = array_index_538982 == array_index_537274 ? add_539154 : sel_539151;
  assign add_539158 = sel_539155 + 8'h01;
  assign sel_539159 = array_index_538982 == array_index_537280 ? add_539158 : sel_539155;
  assign add_539162 = sel_539159 + 8'h01;
  assign sel_539163 = array_index_538982 == array_index_537286 ? add_539162 : sel_539159;
  assign add_539166 = sel_539163 + 8'h01;
  assign sel_539167 = array_index_538982 == array_index_537292 ? add_539166 : sel_539163;
  assign add_539170 = sel_539167 + 8'h01;
  assign sel_539171 = array_index_538982 == array_index_537298 ? add_539170 : sel_539167;
  assign add_539174 = sel_539171 + 8'h01;
  assign sel_539175 = array_index_538982 == array_index_537304 ? add_539174 : sel_539171;
  assign add_539178 = sel_539175 + 8'h01;
  assign sel_539179 = array_index_538982 == array_index_537310 ? add_539178 : sel_539175;
  assign add_539182 = sel_539179 + 8'h01;
  assign sel_539183 = array_index_538982 == array_index_537316 ? add_539182 : sel_539179;
  assign add_539186 = sel_539183 + 8'h01;
  assign sel_539187 = array_index_538982 == array_index_537322 ? add_539186 : sel_539183;
  assign add_539190 = sel_539187 + 8'h01;
  assign sel_539191 = array_index_538982 == array_index_537328 ? add_539190 : sel_539187;
  assign add_539194 = sel_539191 + 8'h01;
  assign sel_539195 = array_index_538982 == array_index_537334 ? add_539194 : sel_539191;
  assign add_539198 = sel_539195 + 8'h01;
  assign sel_539199 = array_index_538982 == array_index_537340 ? add_539198 : sel_539195;
  assign add_539202 = sel_539199 + 8'h01;
  assign sel_539203 = array_index_538982 == array_index_537346 ? add_539202 : sel_539199;
  assign add_539206 = sel_539203 + 8'h01;
  assign sel_539207 = array_index_538982 == array_index_537352 ? add_539206 : sel_539203;
  assign add_539210 = sel_539207 + 8'h01;
  assign sel_539211 = array_index_538982 == array_index_537358 ? add_539210 : sel_539207;
  assign add_539214 = sel_539211 + 8'h01;
  assign sel_539215 = array_index_538982 == array_index_537364 ? add_539214 : sel_539211;
  assign add_539218 = sel_539215 + 8'h01;
  assign sel_539219 = array_index_538982 == array_index_537370 ? add_539218 : sel_539215;
  assign add_539222 = sel_539219 + 8'h01;
  assign sel_539223 = array_index_538982 == array_index_537376 ? add_539222 : sel_539219;
  assign add_539226 = sel_539223 + 8'h01;
  assign sel_539227 = array_index_538982 == array_index_537382 ? add_539226 : sel_539223;
  assign add_539230 = sel_539227 + 8'h01;
  assign sel_539231 = array_index_538982 == array_index_537388 ? add_539230 : sel_539227;
  assign add_539234 = sel_539231 + 8'h01;
  assign sel_539235 = array_index_538982 == array_index_537394 ? add_539234 : sel_539231;
  assign add_539238 = sel_539235 + 8'h01;
  assign sel_539239 = array_index_538982 == array_index_537400 ? add_539238 : sel_539235;
  assign add_539242 = sel_539239 + 8'h01;
  assign sel_539243 = array_index_538982 == array_index_537406 ? add_539242 : sel_539239;
  assign add_539246 = sel_539243 + 8'h01;
  assign sel_539247 = array_index_538982 == array_index_537412 ? add_539246 : sel_539243;
  assign add_539250 = sel_539247 + 8'h01;
  assign sel_539251 = array_index_538982 == array_index_537418 ? add_539250 : sel_539247;
  assign add_539254 = sel_539251 + 8'h01;
  assign sel_539255 = array_index_538982 == array_index_537424 ? add_539254 : sel_539251;
  assign add_539258 = sel_539255 + 8'h01;
  assign sel_539259 = array_index_538982 == array_index_537430 ? add_539258 : sel_539255;
  assign add_539262 = sel_539259 + 8'h01;
  assign sel_539263 = array_index_538982 == array_index_537436 ? add_539262 : sel_539259;
  assign add_539266 = sel_539263 + 8'h01;
  assign sel_539267 = array_index_538982 == array_index_537442 ? add_539266 : sel_539263;
  assign add_539270 = sel_539267 + 8'h01;
  assign sel_539271 = array_index_538982 == array_index_537448 ? add_539270 : sel_539267;
  assign add_539274 = sel_539271 + 8'h01;
  assign sel_539275 = array_index_538982 == array_index_537454 ? add_539274 : sel_539271;
  assign add_539278 = sel_539275 + 8'h01;
  assign sel_539279 = array_index_538982 == array_index_537460 ? add_539278 : sel_539275;
  assign add_539283 = sel_539279 + 8'h01;
  assign array_index_539284 = set1_unflattened[7'h07];
  assign sel_539285 = array_index_538982 == array_index_537466 ? add_539283 : sel_539279;
  assign add_539288 = sel_539285 + 8'h01;
  assign sel_539289 = array_index_539284 == array_index_537012 ? add_539288 : sel_539285;
  assign add_539292 = sel_539289 + 8'h01;
  assign sel_539293 = array_index_539284 == array_index_537016 ? add_539292 : sel_539289;
  assign add_539296 = sel_539293 + 8'h01;
  assign sel_539297 = array_index_539284 == array_index_537024 ? add_539296 : sel_539293;
  assign add_539300 = sel_539297 + 8'h01;
  assign sel_539301 = array_index_539284 == array_index_537032 ? add_539300 : sel_539297;
  assign add_539304 = sel_539301 + 8'h01;
  assign sel_539305 = array_index_539284 == array_index_537040 ? add_539304 : sel_539301;
  assign add_539308 = sel_539305 + 8'h01;
  assign sel_539309 = array_index_539284 == array_index_537048 ? add_539308 : sel_539305;
  assign add_539312 = sel_539309 + 8'h01;
  assign sel_539313 = array_index_539284 == array_index_537056 ? add_539312 : sel_539309;
  assign add_539316 = sel_539313 + 8'h01;
  assign sel_539317 = array_index_539284 == array_index_537064 ? add_539316 : sel_539313;
  assign add_539320 = sel_539317 + 8'h01;
  assign sel_539321 = array_index_539284 == array_index_537070 ? add_539320 : sel_539317;
  assign add_539324 = sel_539321 + 8'h01;
  assign sel_539325 = array_index_539284 == array_index_537076 ? add_539324 : sel_539321;
  assign add_539328 = sel_539325 + 8'h01;
  assign sel_539329 = array_index_539284 == array_index_537082 ? add_539328 : sel_539325;
  assign add_539332 = sel_539329 + 8'h01;
  assign sel_539333 = array_index_539284 == array_index_537088 ? add_539332 : sel_539329;
  assign add_539336 = sel_539333 + 8'h01;
  assign sel_539337 = array_index_539284 == array_index_537094 ? add_539336 : sel_539333;
  assign add_539340 = sel_539337 + 8'h01;
  assign sel_539341 = array_index_539284 == array_index_537100 ? add_539340 : sel_539337;
  assign add_539344 = sel_539341 + 8'h01;
  assign sel_539345 = array_index_539284 == array_index_537106 ? add_539344 : sel_539341;
  assign add_539348 = sel_539345 + 8'h01;
  assign sel_539349 = array_index_539284 == array_index_537112 ? add_539348 : sel_539345;
  assign add_539352 = sel_539349 + 8'h01;
  assign sel_539353 = array_index_539284 == array_index_537118 ? add_539352 : sel_539349;
  assign add_539356 = sel_539353 + 8'h01;
  assign sel_539357 = array_index_539284 == array_index_537124 ? add_539356 : sel_539353;
  assign add_539360 = sel_539357 + 8'h01;
  assign sel_539361 = array_index_539284 == array_index_537130 ? add_539360 : sel_539357;
  assign add_539364 = sel_539361 + 8'h01;
  assign sel_539365 = array_index_539284 == array_index_537136 ? add_539364 : sel_539361;
  assign add_539368 = sel_539365 + 8'h01;
  assign sel_539369 = array_index_539284 == array_index_537142 ? add_539368 : sel_539365;
  assign add_539372 = sel_539369 + 8'h01;
  assign sel_539373 = array_index_539284 == array_index_537148 ? add_539372 : sel_539369;
  assign add_539376 = sel_539373 + 8'h01;
  assign sel_539377 = array_index_539284 == array_index_537154 ? add_539376 : sel_539373;
  assign add_539380 = sel_539377 + 8'h01;
  assign sel_539381 = array_index_539284 == array_index_537160 ? add_539380 : sel_539377;
  assign add_539384 = sel_539381 + 8'h01;
  assign sel_539385 = array_index_539284 == array_index_537166 ? add_539384 : sel_539381;
  assign add_539388 = sel_539385 + 8'h01;
  assign sel_539389 = array_index_539284 == array_index_537172 ? add_539388 : sel_539385;
  assign add_539392 = sel_539389 + 8'h01;
  assign sel_539393 = array_index_539284 == array_index_537178 ? add_539392 : sel_539389;
  assign add_539396 = sel_539393 + 8'h01;
  assign sel_539397 = array_index_539284 == array_index_537184 ? add_539396 : sel_539393;
  assign add_539400 = sel_539397 + 8'h01;
  assign sel_539401 = array_index_539284 == array_index_537190 ? add_539400 : sel_539397;
  assign add_539404 = sel_539401 + 8'h01;
  assign sel_539405 = array_index_539284 == array_index_537196 ? add_539404 : sel_539401;
  assign add_539408 = sel_539405 + 8'h01;
  assign sel_539409 = array_index_539284 == array_index_537202 ? add_539408 : sel_539405;
  assign add_539412 = sel_539409 + 8'h01;
  assign sel_539413 = array_index_539284 == array_index_537208 ? add_539412 : sel_539409;
  assign add_539416 = sel_539413 + 8'h01;
  assign sel_539417 = array_index_539284 == array_index_537214 ? add_539416 : sel_539413;
  assign add_539420 = sel_539417 + 8'h01;
  assign sel_539421 = array_index_539284 == array_index_537220 ? add_539420 : sel_539417;
  assign add_539424 = sel_539421 + 8'h01;
  assign sel_539425 = array_index_539284 == array_index_537226 ? add_539424 : sel_539421;
  assign add_539428 = sel_539425 + 8'h01;
  assign sel_539429 = array_index_539284 == array_index_537232 ? add_539428 : sel_539425;
  assign add_539432 = sel_539429 + 8'h01;
  assign sel_539433 = array_index_539284 == array_index_537238 ? add_539432 : sel_539429;
  assign add_539436 = sel_539433 + 8'h01;
  assign sel_539437 = array_index_539284 == array_index_537244 ? add_539436 : sel_539433;
  assign add_539440 = sel_539437 + 8'h01;
  assign sel_539441 = array_index_539284 == array_index_537250 ? add_539440 : sel_539437;
  assign add_539444 = sel_539441 + 8'h01;
  assign sel_539445 = array_index_539284 == array_index_537256 ? add_539444 : sel_539441;
  assign add_539448 = sel_539445 + 8'h01;
  assign sel_539449 = array_index_539284 == array_index_537262 ? add_539448 : sel_539445;
  assign add_539452 = sel_539449 + 8'h01;
  assign sel_539453 = array_index_539284 == array_index_537268 ? add_539452 : sel_539449;
  assign add_539456 = sel_539453 + 8'h01;
  assign sel_539457 = array_index_539284 == array_index_537274 ? add_539456 : sel_539453;
  assign add_539460 = sel_539457 + 8'h01;
  assign sel_539461 = array_index_539284 == array_index_537280 ? add_539460 : sel_539457;
  assign add_539464 = sel_539461 + 8'h01;
  assign sel_539465 = array_index_539284 == array_index_537286 ? add_539464 : sel_539461;
  assign add_539468 = sel_539465 + 8'h01;
  assign sel_539469 = array_index_539284 == array_index_537292 ? add_539468 : sel_539465;
  assign add_539472 = sel_539469 + 8'h01;
  assign sel_539473 = array_index_539284 == array_index_537298 ? add_539472 : sel_539469;
  assign add_539476 = sel_539473 + 8'h01;
  assign sel_539477 = array_index_539284 == array_index_537304 ? add_539476 : sel_539473;
  assign add_539480 = sel_539477 + 8'h01;
  assign sel_539481 = array_index_539284 == array_index_537310 ? add_539480 : sel_539477;
  assign add_539484 = sel_539481 + 8'h01;
  assign sel_539485 = array_index_539284 == array_index_537316 ? add_539484 : sel_539481;
  assign add_539488 = sel_539485 + 8'h01;
  assign sel_539489 = array_index_539284 == array_index_537322 ? add_539488 : sel_539485;
  assign add_539492 = sel_539489 + 8'h01;
  assign sel_539493 = array_index_539284 == array_index_537328 ? add_539492 : sel_539489;
  assign add_539496 = sel_539493 + 8'h01;
  assign sel_539497 = array_index_539284 == array_index_537334 ? add_539496 : sel_539493;
  assign add_539500 = sel_539497 + 8'h01;
  assign sel_539501 = array_index_539284 == array_index_537340 ? add_539500 : sel_539497;
  assign add_539504 = sel_539501 + 8'h01;
  assign sel_539505 = array_index_539284 == array_index_537346 ? add_539504 : sel_539501;
  assign add_539508 = sel_539505 + 8'h01;
  assign sel_539509 = array_index_539284 == array_index_537352 ? add_539508 : sel_539505;
  assign add_539512 = sel_539509 + 8'h01;
  assign sel_539513 = array_index_539284 == array_index_537358 ? add_539512 : sel_539509;
  assign add_539516 = sel_539513 + 8'h01;
  assign sel_539517 = array_index_539284 == array_index_537364 ? add_539516 : sel_539513;
  assign add_539520 = sel_539517 + 8'h01;
  assign sel_539521 = array_index_539284 == array_index_537370 ? add_539520 : sel_539517;
  assign add_539524 = sel_539521 + 8'h01;
  assign sel_539525 = array_index_539284 == array_index_537376 ? add_539524 : sel_539521;
  assign add_539528 = sel_539525 + 8'h01;
  assign sel_539529 = array_index_539284 == array_index_537382 ? add_539528 : sel_539525;
  assign add_539532 = sel_539529 + 8'h01;
  assign sel_539533 = array_index_539284 == array_index_537388 ? add_539532 : sel_539529;
  assign add_539536 = sel_539533 + 8'h01;
  assign sel_539537 = array_index_539284 == array_index_537394 ? add_539536 : sel_539533;
  assign add_539540 = sel_539537 + 8'h01;
  assign sel_539541 = array_index_539284 == array_index_537400 ? add_539540 : sel_539537;
  assign add_539544 = sel_539541 + 8'h01;
  assign sel_539545 = array_index_539284 == array_index_537406 ? add_539544 : sel_539541;
  assign add_539548 = sel_539545 + 8'h01;
  assign sel_539549 = array_index_539284 == array_index_537412 ? add_539548 : sel_539545;
  assign add_539552 = sel_539549 + 8'h01;
  assign sel_539553 = array_index_539284 == array_index_537418 ? add_539552 : sel_539549;
  assign add_539556 = sel_539553 + 8'h01;
  assign sel_539557 = array_index_539284 == array_index_537424 ? add_539556 : sel_539553;
  assign add_539560 = sel_539557 + 8'h01;
  assign sel_539561 = array_index_539284 == array_index_537430 ? add_539560 : sel_539557;
  assign add_539564 = sel_539561 + 8'h01;
  assign sel_539565 = array_index_539284 == array_index_537436 ? add_539564 : sel_539561;
  assign add_539568 = sel_539565 + 8'h01;
  assign sel_539569 = array_index_539284 == array_index_537442 ? add_539568 : sel_539565;
  assign add_539572 = sel_539569 + 8'h01;
  assign sel_539573 = array_index_539284 == array_index_537448 ? add_539572 : sel_539569;
  assign add_539576 = sel_539573 + 8'h01;
  assign sel_539577 = array_index_539284 == array_index_537454 ? add_539576 : sel_539573;
  assign add_539580 = sel_539577 + 8'h01;
  assign sel_539581 = array_index_539284 == array_index_537460 ? add_539580 : sel_539577;
  assign add_539585 = sel_539581 + 8'h01;
  assign array_index_539586 = set1_unflattened[7'h08];
  assign sel_539587 = array_index_539284 == array_index_537466 ? add_539585 : sel_539581;
  assign add_539590 = sel_539587 + 8'h01;
  assign sel_539591 = array_index_539586 == array_index_537012 ? add_539590 : sel_539587;
  assign add_539594 = sel_539591 + 8'h01;
  assign sel_539595 = array_index_539586 == array_index_537016 ? add_539594 : sel_539591;
  assign add_539598 = sel_539595 + 8'h01;
  assign sel_539599 = array_index_539586 == array_index_537024 ? add_539598 : sel_539595;
  assign add_539602 = sel_539599 + 8'h01;
  assign sel_539603 = array_index_539586 == array_index_537032 ? add_539602 : sel_539599;
  assign add_539606 = sel_539603 + 8'h01;
  assign sel_539607 = array_index_539586 == array_index_537040 ? add_539606 : sel_539603;
  assign add_539610 = sel_539607 + 8'h01;
  assign sel_539611 = array_index_539586 == array_index_537048 ? add_539610 : sel_539607;
  assign add_539614 = sel_539611 + 8'h01;
  assign sel_539615 = array_index_539586 == array_index_537056 ? add_539614 : sel_539611;
  assign add_539618 = sel_539615 + 8'h01;
  assign sel_539619 = array_index_539586 == array_index_537064 ? add_539618 : sel_539615;
  assign add_539622 = sel_539619 + 8'h01;
  assign sel_539623 = array_index_539586 == array_index_537070 ? add_539622 : sel_539619;
  assign add_539626 = sel_539623 + 8'h01;
  assign sel_539627 = array_index_539586 == array_index_537076 ? add_539626 : sel_539623;
  assign add_539630 = sel_539627 + 8'h01;
  assign sel_539631 = array_index_539586 == array_index_537082 ? add_539630 : sel_539627;
  assign add_539634 = sel_539631 + 8'h01;
  assign sel_539635 = array_index_539586 == array_index_537088 ? add_539634 : sel_539631;
  assign add_539638 = sel_539635 + 8'h01;
  assign sel_539639 = array_index_539586 == array_index_537094 ? add_539638 : sel_539635;
  assign add_539642 = sel_539639 + 8'h01;
  assign sel_539643 = array_index_539586 == array_index_537100 ? add_539642 : sel_539639;
  assign add_539646 = sel_539643 + 8'h01;
  assign sel_539647 = array_index_539586 == array_index_537106 ? add_539646 : sel_539643;
  assign add_539650 = sel_539647 + 8'h01;
  assign sel_539651 = array_index_539586 == array_index_537112 ? add_539650 : sel_539647;
  assign add_539654 = sel_539651 + 8'h01;
  assign sel_539655 = array_index_539586 == array_index_537118 ? add_539654 : sel_539651;
  assign add_539658 = sel_539655 + 8'h01;
  assign sel_539659 = array_index_539586 == array_index_537124 ? add_539658 : sel_539655;
  assign add_539662 = sel_539659 + 8'h01;
  assign sel_539663 = array_index_539586 == array_index_537130 ? add_539662 : sel_539659;
  assign add_539666 = sel_539663 + 8'h01;
  assign sel_539667 = array_index_539586 == array_index_537136 ? add_539666 : sel_539663;
  assign add_539670 = sel_539667 + 8'h01;
  assign sel_539671 = array_index_539586 == array_index_537142 ? add_539670 : sel_539667;
  assign add_539674 = sel_539671 + 8'h01;
  assign sel_539675 = array_index_539586 == array_index_537148 ? add_539674 : sel_539671;
  assign add_539678 = sel_539675 + 8'h01;
  assign sel_539679 = array_index_539586 == array_index_537154 ? add_539678 : sel_539675;
  assign add_539682 = sel_539679 + 8'h01;
  assign sel_539683 = array_index_539586 == array_index_537160 ? add_539682 : sel_539679;
  assign add_539686 = sel_539683 + 8'h01;
  assign sel_539687 = array_index_539586 == array_index_537166 ? add_539686 : sel_539683;
  assign add_539690 = sel_539687 + 8'h01;
  assign sel_539691 = array_index_539586 == array_index_537172 ? add_539690 : sel_539687;
  assign add_539694 = sel_539691 + 8'h01;
  assign sel_539695 = array_index_539586 == array_index_537178 ? add_539694 : sel_539691;
  assign add_539698 = sel_539695 + 8'h01;
  assign sel_539699 = array_index_539586 == array_index_537184 ? add_539698 : sel_539695;
  assign add_539702 = sel_539699 + 8'h01;
  assign sel_539703 = array_index_539586 == array_index_537190 ? add_539702 : sel_539699;
  assign add_539706 = sel_539703 + 8'h01;
  assign sel_539707 = array_index_539586 == array_index_537196 ? add_539706 : sel_539703;
  assign add_539710 = sel_539707 + 8'h01;
  assign sel_539711 = array_index_539586 == array_index_537202 ? add_539710 : sel_539707;
  assign add_539714 = sel_539711 + 8'h01;
  assign sel_539715 = array_index_539586 == array_index_537208 ? add_539714 : sel_539711;
  assign add_539718 = sel_539715 + 8'h01;
  assign sel_539719 = array_index_539586 == array_index_537214 ? add_539718 : sel_539715;
  assign add_539722 = sel_539719 + 8'h01;
  assign sel_539723 = array_index_539586 == array_index_537220 ? add_539722 : sel_539719;
  assign add_539726 = sel_539723 + 8'h01;
  assign sel_539727 = array_index_539586 == array_index_537226 ? add_539726 : sel_539723;
  assign add_539730 = sel_539727 + 8'h01;
  assign sel_539731 = array_index_539586 == array_index_537232 ? add_539730 : sel_539727;
  assign add_539734 = sel_539731 + 8'h01;
  assign sel_539735 = array_index_539586 == array_index_537238 ? add_539734 : sel_539731;
  assign add_539738 = sel_539735 + 8'h01;
  assign sel_539739 = array_index_539586 == array_index_537244 ? add_539738 : sel_539735;
  assign add_539742 = sel_539739 + 8'h01;
  assign sel_539743 = array_index_539586 == array_index_537250 ? add_539742 : sel_539739;
  assign add_539746 = sel_539743 + 8'h01;
  assign sel_539747 = array_index_539586 == array_index_537256 ? add_539746 : sel_539743;
  assign add_539750 = sel_539747 + 8'h01;
  assign sel_539751 = array_index_539586 == array_index_537262 ? add_539750 : sel_539747;
  assign add_539754 = sel_539751 + 8'h01;
  assign sel_539755 = array_index_539586 == array_index_537268 ? add_539754 : sel_539751;
  assign add_539758 = sel_539755 + 8'h01;
  assign sel_539759 = array_index_539586 == array_index_537274 ? add_539758 : sel_539755;
  assign add_539762 = sel_539759 + 8'h01;
  assign sel_539763 = array_index_539586 == array_index_537280 ? add_539762 : sel_539759;
  assign add_539766 = sel_539763 + 8'h01;
  assign sel_539767 = array_index_539586 == array_index_537286 ? add_539766 : sel_539763;
  assign add_539770 = sel_539767 + 8'h01;
  assign sel_539771 = array_index_539586 == array_index_537292 ? add_539770 : sel_539767;
  assign add_539774 = sel_539771 + 8'h01;
  assign sel_539775 = array_index_539586 == array_index_537298 ? add_539774 : sel_539771;
  assign add_539778 = sel_539775 + 8'h01;
  assign sel_539779 = array_index_539586 == array_index_537304 ? add_539778 : sel_539775;
  assign add_539782 = sel_539779 + 8'h01;
  assign sel_539783 = array_index_539586 == array_index_537310 ? add_539782 : sel_539779;
  assign add_539786 = sel_539783 + 8'h01;
  assign sel_539787 = array_index_539586 == array_index_537316 ? add_539786 : sel_539783;
  assign add_539790 = sel_539787 + 8'h01;
  assign sel_539791 = array_index_539586 == array_index_537322 ? add_539790 : sel_539787;
  assign add_539794 = sel_539791 + 8'h01;
  assign sel_539795 = array_index_539586 == array_index_537328 ? add_539794 : sel_539791;
  assign add_539798 = sel_539795 + 8'h01;
  assign sel_539799 = array_index_539586 == array_index_537334 ? add_539798 : sel_539795;
  assign add_539802 = sel_539799 + 8'h01;
  assign sel_539803 = array_index_539586 == array_index_537340 ? add_539802 : sel_539799;
  assign add_539806 = sel_539803 + 8'h01;
  assign sel_539807 = array_index_539586 == array_index_537346 ? add_539806 : sel_539803;
  assign add_539810 = sel_539807 + 8'h01;
  assign sel_539811 = array_index_539586 == array_index_537352 ? add_539810 : sel_539807;
  assign add_539814 = sel_539811 + 8'h01;
  assign sel_539815 = array_index_539586 == array_index_537358 ? add_539814 : sel_539811;
  assign add_539818 = sel_539815 + 8'h01;
  assign sel_539819 = array_index_539586 == array_index_537364 ? add_539818 : sel_539815;
  assign add_539822 = sel_539819 + 8'h01;
  assign sel_539823 = array_index_539586 == array_index_537370 ? add_539822 : sel_539819;
  assign add_539826 = sel_539823 + 8'h01;
  assign sel_539827 = array_index_539586 == array_index_537376 ? add_539826 : sel_539823;
  assign add_539830 = sel_539827 + 8'h01;
  assign sel_539831 = array_index_539586 == array_index_537382 ? add_539830 : sel_539827;
  assign add_539834 = sel_539831 + 8'h01;
  assign sel_539835 = array_index_539586 == array_index_537388 ? add_539834 : sel_539831;
  assign add_539838 = sel_539835 + 8'h01;
  assign sel_539839 = array_index_539586 == array_index_537394 ? add_539838 : sel_539835;
  assign add_539842 = sel_539839 + 8'h01;
  assign sel_539843 = array_index_539586 == array_index_537400 ? add_539842 : sel_539839;
  assign add_539846 = sel_539843 + 8'h01;
  assign sel_539847 = array_index_539586 == array_index_537406 ? add_539846 : sel_539843;
  assign add_539850 = sel_539847 + 8'h01;
  assign sel_539851 = array_index_539586 == array_index_537412 ? add_539850 : sel_539847;
  assign add_539854 = sel_539851 + 8'h01;
  assign sel_539855 = array_index_539586 == array_index_537418 ? add_539854 : sel_539851;
  assign add_539858 = sel_539855 + 8'h01;
  assign sel_539859 = array_index_539586 == array_index_537424 ? add_539858 : sel_539855;
  assign add_539862 = sel_539859 + 8'h01;
  assign sel_539863 = array_index_539586 == array_index_537430 ? add_539862 : sel_539859;
  assign add_539866 = sel_539863 + 8'h01;
  assign sel_539867 = array_index_539586 == array_index_537436 ? add_539866 : sel_539863;
  assign add_539870 = sel_539867 + 8'h01;
  assign sel_539871 = array_index_539586 == array_index_537442 ? add_539870 : sel_539867;
  assign add_539874 = sel_539871 + 8'h01;
  assign sel_539875 = array_index_539586 == array_index_537448 ? add_539874 : sel_539871;
  assign add_539878 = sel_539875 + 8'h01;
  assign sel_539879 = array_index_539586 == array_index_537454 ? add_539878 : sel_539875;
  assign add_539882 = sel_539879 + 8'h01;
  assign sel_539883 = array_index_539586 == array_index_537460 ? add_539882 : sel_539879;
  assign add_539887 = sel_539883 + 8'h01;
  assign array_index_539888 = set1_unflattened[7'h09];
  assign sel_539889 = array_index_539586 == array_index_537466 ? add_539887 : sel_539883;
  assign add_539892 = sel_539889 + 8'h01;
  assign sel_539893 = array_index_539888 == array_index_537012 ? add_539892 : sel_539889;
  assign add_539896 = sel_539893 + 8'h01;
  assign sel_539897 = array_index_539888 == array_index_537016 ? add_539896 : sel_539893;
  assign add_539900 = sel_539897 + 8'h01;
  assign sel_539901 = array_index_539888 == array_index_537024 ? add_539900 : sel_539897;
  assign add_539904 = sel_539901 + 8'h01;
  assign sel_539905 = array_index_539888 == array_index_537032 ? add_539904 : sel_539901;
  assign add_539908 = sel_539905 + 8'h01;
  assign sel_539909 = array_index_539888 == array_index_537040 ? add_539908 : sel_539905;
  assign add_539912 = sel_539909 + 8'h01;
  assign sel_539913 = array_index_539888 == array_index_537048 ? add_539912 : sel_539909;
  assign add_539916 = sel_539913 + 8'h01;
  assign sel_539917 = array_index_539888 == array_index_537056 ? add_539916 : sel_539913;
  assign add_539920 = sel_539917 + 8'h01;
  assign sel_539921 = array_index_539888 == array_index_537064 ? add_539920 : sel_539917;
  assign add_539924 = sel_539921 + 8'h01;
  assign sel_539925 = array_index_539888 == array_index_537070 ? add_539924 : sel_539921;
  assign add_539928 = sel_539925 + 8'h01;
  assign sel_539929 = array_index_539888 == array_index_537076 ? add_539928 : sel_539925;
  assign add_539932 = sel_539929 + 8'h01;
  assign sel_539933 = array_index_539888 == array_index_537082 ? add_539932 : sel_539929;
  assign add_539936 = sel_539933 + 8'h01;
  assign sel_539937 = array_index_539888 == array_index_537088 ? add_539936 : sel_539933;
  assign add_539940 = sel_539937 + 8'h01;
  assign sel_539941 = array_index_539888 == array_index_537094 ? add_539940 : sel_539937;
  assign add_539944 = sel_539941 + 8'h01;
  assign sel_539945 = array_index_539888 == array_index_537100 ? add_539944 : sel_539941;
  assign add_539948 = sel_539945 + 8'h01;
  assign sel_539949 = array_index_539888 == array_index_537106 ? add_539948 : sel_539945;
  assign add_539952 = sel_539949 + 8'h01;
  assign sel_539953 = array_index_539888 == array_index_537112 ? add_539952 : sel_539949;
  assign add_539956 = sel_539953 + 8'h01;
  assign sel_539957 = array_index_539888 == array_index_537118 ? add_539956 : sel_539953;
  assign add_539960 = sel_539957 + 8'h01;
  assign sel_539961 = array_index_539888 == array_index_537124 ? add_539960 : sel_539957;
  assign add_539964 = sel_539961 + 8'h01;
  assign sel_539965 = array_index_539888 == array_index_537130 ? add_539964 : sel_539961;
  assign add_539968 = sel_539965 + 8'h01;
  assign sel_539969 = array_index_539888 == array_index_537136 ? add_539968 : sel_539965;
  assign add_539972 = sel_539969 + 8'h01;
  assign sel_539973 = array_index_539888 == array_index_537142 ? add_539972 : sel_539969;
  assign add_539976 = sel_539973 + 8'h01;
  assign sel_539977 = array_index_539888 == array_index_537148 ? add_539976 : sel_539973;
  assign add_539980 = sel_539977 + 8'h01;
  assign sel_539981 = array_index_539888 == array_index_537154 ? add_539980 : sel_539977;
  assign add_539984 = sel_539981 + 8'h01;
  assign sel_539985 = array_index_539888 == array_index_537160 ? add_539984 : sel_539981;
  assign add_539988 = sel_539985 + 8'h01;
  assign sel_539989 = array_index_539888 == array_index_537166 ? add_539988 : sel_539985;
  assign add_539992 = sel_539989 + 8'h01;
  assign sel_539993 = array_index_539888 == array_index_537172 ? add_539992 : sel_539989;
  assign add_539996 = sel_539993 + 8'h01;
  assign sel_539997 = array_index_539888 == array_index_537178 ? add_539996 : sel_539993;
  assign add_540000 = sel_539997 + 8'h01;
  assign sel_540001 = array_index_539888 == array_index_537184 ? add_540000 : sel_539997;
  assign add_540004 = sel_540001 + 8'h01;
  assign sel_540005 = array_index_539888 == array_index_537190 ? add_540004 : sel_540001;
  assign add_540008 = sel_540005 + 8'h01;
  assign sel_540009 = array_index_539888 == array_index_537196 ? add_540008 : sel_540005;
  assign add_540012 = sel_540009 + 8'h01;
  assign sel_540013 = array_index_539888 == array_index_537202 ? add_540012 : sel_540009;
  assign add_540016 = sel_540013 + 8'h01;
  assign sel_540017 = array_index_539888 == array_index_537208 ? add_540016 : sel_540013;
  assign add_540020 = sel_540017 + 8'h01;
  assign sel_540021 = array_index_539888 == array_index_537214 ? add_540020 : sel_540017;
  assign add_540024 = sel_540021 + 8'h01;
  assign sel_540025 = array_index_539888 == array_index_537220 ? add_540024 : sel_540021;
  assign add_540028 = sel_540025 + 8'h01;
  assign sel_540029 = array_index_539888 == array_index_537226 ? add_540028 : sel_540025;
  assign add_540032 = sel_540029 + 8'h01;
  assign sel_540033 = array_index_539888 == array_index_537232 ? add_540032 : sel_540029;
  assign add_540036 = sel_540033 + 8'h01;
  assign sel_540037 = array_index_539888 == array_index_537238 ? add_540036 : sel_540033;
  assign add_540040 = sel_540037 + 8'h01;
  assign sel_540041 = array_index_539888 == array_index_537244 ? add_540040 : sel_540037;
  assign add_540044 = sel_540041 + 8'h01;
  assign sel_540045 = array_index_539888 == array_index_537250 ? add_540044 : sel_540041;
  assign add_540048 = sel_540045 + 8'h01;
  assign sel_540049 = array_index_539888 == array_index_537256 ? add_540048 : sel_540045;
  assign add_540052 = sel_540049 + 8'h01;
  assign sel_540053 = array_index_539888 == array_index_537262 ? add_540052 : sel_540049;
  assign add_540056 = sel_540053 + 8'h01;
  assign sel_540057 = array_index_539888 == array_index_537268 ? add_540056 : sel_540053;
  assign add_540060 = sel_540057 + 8'h01;
  assign sel_540061 = array_index_539888 == array_index_537274 ? add_540060 : sel_540057;
  assign add_540064 = sel_540061 + 8'h01;
  assign sel_540065 = array_index_539888 == array_index_537280 ? add_540064 : sel_540061;
  assign add_540068 = sel_540065 + 8'h01;
  assign sel_540069 = array_index_539888 == array_index_537286 ? add_540068 : sel_540065;
  assign add_540072 = sel_540069 + 8'h01;
  assign sel_540073 = array_index_539888 == array_index_537292 ? add_540072 : sel_540069;
  assign add_540076 = sel_540073 + 8'h01;
  assign sel_540077 = array_index_539888 == array_index_537298 ? add_540076 : sel_540073;
  assign add_540080 = sel_540077 + 8'h01;
  assign sel_540081 = array_index_539888 == array_index_537304 ? add_540080 : sel_540077;
  assign add_540084 = sel_540081 + 8'h01;
  assign sel_540085 = array_index_539888 == array_index_537310 ? add_540084 : sel_540081;
  assign add_540088 = sel_540085 + 8'h01;
  assign sel_540089 = array_index_539888 == array_index_537316 ? add_540088 : sel_540085;
  assign add_540092 = sel_540089 + 8'h01;
  assign sel_540093 = array_index_539888 == array_index_537322 ? add_540092 : sel_540089;
  assign add_540096 = sel_540093 + 8'h01;
  assign sel_540097 = array_index_539888 == array_index_537328 ? add_540096 : sel_540093;
  assign add_540100 = sel_540097 + 8'h01;
  assign sel_540101 = array_index_539888 == array_index_537334 ? add_540100 : sel_540097;
  assign add_540104 = sel_540101 + 8'h01;
  assign sel_540105 = array_index_539888 == array_index_537340 ? add_540104 : sel_540101;
  assign add_540108 = sel_540105 + 8'h01;
  assign sel_540109 = array_index_539888 == array_index_537346 ? add_540108 : sel_540105;
  assign add_540112 = sel_540109 + 8'h01;
  assign sel_540113 = array_index_539888 == array_index_537352 ? add_540112 : sel_540109;
  assign add_540116 = sel_540113 + 8'h01;
  assign sel_540117 = array_index_539888 == array_index_537358 ? add_540116 : sel_540113;
  assign add_540120 = sel_540117 + 8'h01;
  assign sel_540121 = array_index_539888 == array_index_537364 ? add_540120 : sel_540117;
  assign add_540124 = sel_540121 + 8'h01;
  assign sel_540125 = array_index_539888 == array_index_537370 ? add_540124 : sel_540121;
  assign add_540128 = sel_540125 + 8'h01;
  assign sel_540129 = array_index_539888 == array_index_537376 ? add_540128 : sel_540125;
  assign add_540132 = sel_540129 + 8'h01;
  assign sel_540133 = array_index_539888 == array_index_537382 ? add_540132 : sel_540129;
  assign add_540136 = sel_540133 + 8'h01;
  assign sel_540137 = array_index_539888 == array_index_537388 ? add_540136 : sel_540133;
  assign add_540140 = sel_540137 + 8'h01;
  assign sel_540141 = array_index_539888 == array_index_537394 ? add_540140 : sel_540137;
  assign add_540144 = sel_540141 + 8'h01;
  assign sel_540145 = array_index_539888 == array_index_537400 ? add_540144 : sel_540141;
  assign add_540148 = sel_540145 + 8'h01;
  assign sel_540149 = array_index_539888 == array_index_537406 ? add_540148 : sel_540145;
  assign add_540152 = sel_540149 + 8'h01;
  assign sel_540153 = array_index_539888 == array_index_537412 ? add_540152 : sel_540149;
  assign add_540156 = sel_540153 + 8'h01;
  assign sel_540157 = array_index_539888 == array_index_537418 ? add_540156 : sel_540153;
  assign add_540160 = sel_540157 + 8'h01;
  assign sel_540161 = array_index_539888 == array_index_537424 ? add_540160 : sel_540157;
  assign add_540164 = sel_540161 + 8'h01;
  assign sel_540165 = array_index_539888 == array_index_537430 ? add_540164 : sel_540161;
  assign add_540168 = sel_540165 + 8'h01;
  assign sel_540169 = array_index_539888 == array_index_537436 ? add_540168 : sel_540165;
  assign add_540172 = sel_540169 + 8'h01;
  assign sel_540173 = array_index_539888 == array_index_537442 ? add_540172 : sel_540169;
  assign add_540176 = sel_540173 + 8'h01;
  assign sel_540177 = array_index_539888 == array_index_537448 ? add_540176 : sel_540173;
  assign add_540180 = sel_540177 + 8'h01;
  assign sel_540181 = array_index_539888 == array_index_537454 ? add_540180 : sel_540177;
  assign add_540184 = sel_540181 + 8'h01;
  assign sel_540185 = array_index_539888 == array_index_537460 ? add_540184 : sel_540181;
  assign add_540189 = sel_540185 + 8'h01;
  assign array_index_540190 = set1_unflattened[7'h0a];
  assign sel_540191 = array_index_539888 == array_index_537466 ? add_540189 : sel_540185;
  assign add_540194 = sel_540191 + 8'h01;
  assign sel_540195 = array_index_540190 == array_index_537012 ? add_540194 : sel_540191;
  assign add_540198 = sel_540195 + 8'h01;
  assign sel_540199 = array_index_540190 == array_index_537016 ? add_540198 : sel_540195;
  assign add_540202 = sel_540199 + 8'h01;
  assign sel_540203 = array_index_540190 == array_index_537024 ? add_540202 : sel_540199;
  assign add_540206 = sel_540203 + 8'h01;
  assign sel_540207 = array_index_540190 == array_index_537032 ? add_540206 : sel_540203;
  assign add_540210 = sel_540207 + 8'h01;
  assign sel_540211 = array_index_540190 == array_index_537040 ? add_540210 : sel_540207;
  assign add_540214 = sel_540211 + 8'h01;
  assign sel_540215 = array_index_540190 == array_index_537048 ? add_540214 : sel_540211;
  assign add_540218 = sel_540215 + 8'h01;
  assign sel_540219 = array_index_540190 == array_index_537056 ? add_540218 : sel_540215;
  assign add_540222 = sel_540219 + 8'h01;
  assign sel_540223 = array_index_540190 == array_index_537064 ? add_540222 : sel_540219;
  assign add_540226 = sel_540223 + 8'h01;
  assign sel_540227 = array_index_540190 == array_index_537070 ? add_540226 : sel_540223;
  assign add_540230 = sel_540227 + 8'h01;
  assign sel_540231 = array_index_540190 == array_index_537076 ? add_540230 : sel_540227;
  assign add_540234 = sel_540231 + 8'h01;
  assign sel_540235 = array_index_540190 == array_index_537082 ? add_540234 : sel_540231;
  assign add_540238 = sel_540235 + 8'h01;
  assign sel_540239 = array_index_540190 == array_index_537088 ? add_540238 : sel_540235;
  assign add_540242 = sel_540239 + 8'h01;
  assign sel_540243 = array_index_540190 == array_index_537094 ? add_540242 : sel_540239;
  assign add_540246 = sel_540243 + 8'h01;
  assign sel_540247 = array_index_540190 == array_index_537100 ? add_540246 : sel_540243;
  assign add_540250 = sel_540247 + 8'h01;
  assign sel_540251 = array_index_540190 == array_index_537106 ? add_540250 : sel_540247;
  assign add_540254 = sel_540251 + 8'h01;
  assign sel_540255 = array_index_540190 == array_index_537112 ? add_540254 : sel_540251;
  assign add_540258 = sel_540255 + 8'h01;
  assign sel_540259 = array_index_540190 == array_index_537118 ? add_540258 : sel_540255;
  assign add_540262 = sel_540259 + 8'h01;
  assign sel_540263 = array_index_540190 == array_index_537124 ? add_540262 : sel_540259;
  assign add_540266 = sel_540263 + 8'h01;
  assign sel_540267 = array_index_540190 == array_index_537130 ? add_540266 : sel_540263;
  assign add_540270 = sel_540267 + 8'h01;
  assign sel_540271 = array_index_540190 == array_index_537136 ? add_540270 : sel_540267;
  assign add_540274 = sel_540271 + 8'h01;
  assign sel_540275 = array_index_540190 == array_index_537142 ? add_540274 : sel_540271;
  assign add_540278 = sel_540275 + 8'h01;
  assign sel_540279 = array_index_540190 == array_index_537148 ? add_540278 : sel_540275;
  assign add_540282 = sel_540279 + 8'h01;
  assign sel_540283 = array_index_540190 == array_index_537154 ? add_540282 : sel_540279;
  assign add_540286 = sel_540283 + 8'h01;
  assign sel_540287 = array_index_540190 == array_index_537160 ? add_540286 : sel_540283;
  assign add_540290 = sel_540287 + 8'h01;
  assign sel_540291 = array_index_540190 == array_index_537166 ? add_540290 : sel_540287;
  assign add_540294 = sel_540291 + 8'h01;
  assign sel_540295 = array_index_540190 == array_index_537172 ? add_540294 : sel_540291;
  assign add_540298 = sel_540295 + 8'h01;
  assign sel_540299 = array_index_540190 == array_index_537178 ? add_540298 : sel_540295;
  assign add_540302 = sel_540299 + 8'h01;
  assign sel_540303 = array_index_540190 == array_index_537184 ? add_540302 : sel_540299;
  assign add_540306 = sel_540303 + 8'h01;
  assign sel_540307 = array_index_540190 == array_index_537190 ? add_540306 : sel_540303;
  assign add_540310 = sel_540307 + 8'h01;
  assign sel_540311 = array_index_540190 == array_index_537196 ? add_540310 : sel_540307;
  assign add_540314 = sel_540311 + 8'h01;
  assign sel_540315 = array_index_540190 == array_index_537202 ? add_540314 : sel_540311;
  assign add_540318 = sel_540315 + 8'h01;
  assign sel_540319 = array_index_540190 == array_index_537208 ? add_540318 : sel_540315;
  assign add_540322 = sel_540319 + 8'h01;
  assign sel_540323 = array_index_540190 == array_index_537214 ? add_540322 : sel_540319;
  assign add_540326 = sel_540323 + 8'h01;
  assign sel_540327 = array_index_540190 == array_index_537220 ? add_540326 : sel_540323;
  assign add_540330 = sel_540327 + 8'h01;
  assign sel_540331 = array_index_540190 == array_index_537226 ? add_540330 : sel_540327;
  assign add_540334 = sel_540331 + 8'h01;
  assign sel_540335 = array_index_540190 == array_index_537232 ? add_540334 : sel_540331;
  assign add_540338 = sel_540335 + 8'h01;
  assign sel_540339 = array_index_540190 == array_index_537238 ? add_540338 : sel_540335;
  assign add_540342 = sel_540339 + 8'h01;
  assign sel_540343 = array_index_540190 == array_index_537244 ? add_540342 : sel_540339;
  assign add_540346 = sel_540343 + 8'h01;
  assign sel_540347 = array_index_540190 == array_index_537250 ? add_540346 : sel_540343;
  assign add_540350 = sel_540347 + 8'h01;
  assign sel_540351 = array_index_540190 == array_index_537256 ? add_540350 : sel_540347;
  assign add_540354 = sel_540351 + 8'h01;
  assign sel_540355 = array_index_540190 == array_index_537262 ? add_540354 : sel_540351;
  assign add_540358 = sel_540355 + 8'h01;
  assign sel_540359 = array_index_540190 == array_index_537268 ? add_540358 : sel_540355;
  assign add_540362 = sel_540359 + 8'h01;
  assign sel_540363 = array_index_540190 == array_index_537274 ? add_540362 : sel_540359;
  assign add_540366 = sel_540363 + 8'h01;
  assign sel_540367 = array_index_540190 == array_index_537280 ? add_540366 : sel_540363;
  assign add_540370 = sel_540367 + 8'h01;
  assign sel_540371 = array_index_540190 == array_index_537286 ? add_540370 : sel_540367;
  assign add_540374 = sel_540371 + 8'h01;
  assign sel_540375 = array_index_540190 == array_index_537292 ? add_540374 : sel_540371;
  assign add_540378 = sel_540375 + 8'h01;
  assign sel_540379 = array_index_540190 == array_index_537298 ? add_540378 : sel_540375;
  assign add_540382 = sel_540379 + 8'h01;
  assign sel_540383 = array_index_540190 == array_index_537304 ? add_540382 : sel_540379;
  assign add_540386 = sel_540383 + 8'h01;
  assign sel_540387 = array_index_540190 == array_index_537310 ? add_540386 : sel_540383;
  assign add_540390 = sel_540387 + 8'h01;
  assign sel_540391 = array_index_540190 == array_index_537316 ? add_540390 : sel_540387;
  assign add_540394 = sel_540391 + 8'h01;
  assign sel_540395 = array_index_540190 == array_index_537322 ? add_540394 : sel_540391;
  assign add_540398 = sel_540395 + 8'h01;
  assign sel_540399 = array_index_540190 == array_index_537328 ? add_540398 : sel_540395;
  assign add_540402 = sel_540399 + 8'h01;
  assign sel_540403 = array_index_540190 == array_index_537334 ? add_540402 : sel_540399;
  assign add_540406 = sel_540403 + 8'h01;
  assign sel_540407 = array_index_540190 == array_index_537340 ? add_540406 : sel_540403;
  assign add_540410 = sel_540407 + 8'h01;
  assign sel_540411 = array_index_540190 == array_index_537346 ? add_540410 : sel_540407;
  assign add_540414 = sel_540411 + 8'h01;
  assign sel_540415 = array_index_540190 == array_index_537352 ? add_540414 : sel_540411;
  assign add_540418 = sel_540415 + 8'h01;
  assign sel_540419 = array_index_540190 == array_index_537358 ? add_540418 : sel_540415;
  assign add_540422 = sel_540419 + 8'h01;
  assign sel_540423 = array_index_540190 == array_index_537364 ? add_540422 : sel_540419;
  assign add_540426 = sel_540423 + 8'h01;
  assign sel_540427 = array_index_540190 == array_index_537370 ? add_540426 : sel_540423;
  assign add_540430 = sel_540427 + 8'h01;
  assign sel_540431 = array_index_540190 == array_index_537376 ? add_540430 : sel_540427;
  assign add_540434 = sel_540431 + 8'h01;
  assign sel_540435 = array_index_540190 == array_index_537382 ? add_540434 : sel_540431;
  assign add_540438 = sel_540435 + 8'h01;
  assign sel_540439 = array_index_540190 == array_index_537388 ? add_540438 : sel_540435;
  assign add_540442 = sel_540439 + 8'h01;
  assign sel_540443 = array_index_540190 == array_index_537394 ? add_540442 : sel_540439;
  assign add_540446 = sel_540443 + 8'h01;
  assign sel_540447 = array_index_540190 == array_index_537400 ? add_540446 : sel_540443;
  assign add_540450 = sel_540447 + 8'h01;
  assign sel_540451 = array_index_540190 == array_index_537406 ? add_540450 : sel_540447;
  assign add_540454 = sel_540451 + 8'h01;
  assign sel_540455 = array_index_540190 == array_index_537412 ? add_540454 : sel_540451;
  assign add_540458 = sel_540455 + 8'h01;
  assign sel_540459 = array_index_540190 == array_index_537418 ? add_540458 : sel_540455;
  assign add_540462 = sel_540459 + 8'h01;
  assign sel_540463 = array_index_540190 == array_index_537424 ? add_540462 : sel_540459;
  assign add_540466 = sel_540463 + 8'h01;
  assign sel_540467 = array_index_540190 == array_index_537430 ? add_540466 : sel_540463;
  assign add_540470 = sel_540467 + 8'h01;
  assign sel_540471 = array_index_540190 == array_index_537436 ? add_540470 : sel_540467;
  assign add_540474 = sel_540471 + 8'h01;
  assign sel_540475 = array_index_540190 == array_index_537442 ? add_540474 : sel_540471;
  assign add_540478 = sel_540475 + 8'h01;
  assign sel_540479 = array_index_540190 == array_index_537448 ? add_540478 : sel_540475;
  assign add_540482 = sel_540479 + 8'h01;
  assign sel_540483 = array_index_540190 == array_index_537454 ? add_540482 : sel_540479;
  assign add_540486 = sel_540483 + 8'h01;
  assign sel_540487 = array_index_540190 == array_index_537460 ? add_540486 : sel_540483;
  assign add_540491 = sel_540487 + 8'h01;
  assign array_index_540492 = set1_unflattened[7'h0b];
  assign sel_540493 = array_index_540190 == array_index_537466 ? add_540491 : sel_540487;
  assign add_540496 = sel_540493 + 8'h01;
  assign sel_540497 = array_index_540492 == array_index_537012 ? add_540496 : sel_540493;
  assign add_540500 = sel_540497 + 8'h01;
  assign sel_540501 = array_index_540492 == array_index_537016 ? add_540500 : sel_540497;
  assign add_540504 = sel_540501 + 8'h01;
  assign sel_540505 = array_index_540492 == array_index_537024 ? add_540504 : sel_540501;
  assign add_540508 = sel_540505 + 8'h01;
  assign sel_540509 = array_index_540492 == array_index_537032 ? add_540508 : sel_540505;
  assign add_540512 = sel_540509 + 8'h01;
  assign sel_540513 = array_index_540492 == array_index_537040 ? add_540512 : sel_540509;
  assign add_540516 = sel_540513 + 8'h01;
  assign sel_540517 = array_index_540492 == array_index_537048 ? add_540516 : sel_540513;
  assign add_540520 = sel_540517 + 8'h01;
  assign sel_540521 = array_index_540492 == array_index_537056 ? add_540520 : sel_540517;
  assign add_540524 = sel_540521 + 8'h01;
  assign sel_540525 = array_index_540492 == array_index_537064 ? add_540524 : sel_540521;
  assign add_540528 = sel_540525 + 8'h01;
  assign sel_540529 = array_index_540492 == array_index_537070 ? add_540528 : sel_540525;
  assign add_540532 = sel_540529 + 8'h01;
  assign sel_540533 = array_index_540492 == array_index_537076 ? add_540532 : sel_540529;
  assign add_540536 = sel_540533 + 8'h01;
  assign sel_540537 = array_index_540492 == array_index_537082 ? add_540536 : sel_540533;
  assign add_540540 = sel_540537 + 8'h01;
  assign sel_540541 = array_index_540492 == array_index_537088 ? add_540540 : sel_540537;
  assign add_540544 = sel_540541 + 8'h01;
  assign sel_540545 = array_index_540492 == array_index_537094 ? add_540544 : sel_540541;
  assign add_540548 = sel_540545 + 8'h01;
  assign sel_540549 = array_index_540492 == array_index_537100 ? add_540548 : sel_540545;
  assign add_540552 = sel_540549 + 8'h01;
  assign sel_540553 = array_index_540492 == array_index_537106 ? add_540552 : sel_540549;
  assign add_540556 = sel_540553 + 8'h01;
  assign sel_540557 = array_index_540492 == array_index_537112 ? add_540556 : sel_540553;
  assign add_540560 = sel_540557 + 8'h01;
  assign sel_540561 = array_index_540492 == array_index_537118 ? add_540560 : sel_540557;
  assign add_540564 = sel_540561 + 8'h01;
  assign sel_540565 = array_index_540492 == array_index_537124 ? add_540564 : sel_540561;
  assign add_540568 = sel_540565 + 8'h01;
  assign sel_540569 = array_index_540492 == array_index_537130 ? add_540568 : sel_540565;
  assign add_540572 = sel_540569 + 8'h01;
  assign sel_540573 = array_index_540492 == array_index_537136 ? add_540572 : sel_540569;
  assign add_540576 = sel_540573 + 8'h01;
  assign sel_540577 = array_index_540492 == array_index_537142 ? add_540576 : sel_540573;
  assign add_540580 = sel_540577 + 8'h01;
  assign sel_540581 = array_index_540492 == array_index_537148 ? add_540580 : sel_540577;
  assign add_540584 = sel_540581 + 8'h01;
  assign sel_540585 = array_index_540492 == array_index_537154 ? add_540584 : sel_540581;
  assign add_540588 = sel_540585 + 8'h01;
  assign sel_540589 = array_index_540492 == array_index_537160 ? add_540588 : sel_540585;
  assign add_540592 = sel_540589 + 8'h01;
  assign sel_540593 = array_index_540492 == array_index_537166 ? add_540592 : sel_540589;
  assign add_540596 = sel_540593 + 8'h01;
  assign sel_540597 = array_index_540492 == array_index_537172 ? add_540596 : sel_540593;
  assign add_540600 = sel_540597 + 8'h01;
  assign sel_540601 = array_index_540492 == array_index_537178 ? add_540600 : sel_540597;
  assign add_540604 = sel_540601 + 8'h01;
  assign sel_540605 = array_index_540492 == array_index_537184 ? add_540604 : sel_540601;
  assign add_540608 = sel_540605 + 8'h01;
  assign sel_540609 = array_index_540492 == array_index_537190 ? add_540608 : sel_540605;
  assign add_540612 = sel_540609 + 8'h01;
  assign sel_540613 = array_index_540492 == array_index_537196 ? add_540612 : sel_540609;
  assign add_540616 = sel_540613 + 8'h01;
  assign sel_540617 = array_index_540492 == array_index_537202 ? add_540616 : sel_540613;
  assign add_540620 = sel_540617 + 8'h01;
  assign sel_540621 = array_index_540492 == array_index_537208 ? add_540620 : sel_540617;
  assign add_540624 = sel_540621 + 8'h01;
  assign sel_540625 = array_index_540492 == array_index_537214 ? add_540624 : sel_540621;
  assign add_540628 = sel_540625 + 8'h01;
  assign sel_540629 = array_index_540492 == array_index_537220 ? add_540628 : sel_540625;
  assign add_540632 = sel_540629 + 8'h01;
  assign sel_540633 = array_index_540492 == array_index_537226 ? add_540632 : sel_540629;
  assign add_540636 = sel_540633 + 8'h01;
  assign sel_540637 = array_index_540492 == array_index_537232 ? add_540636 : sel_540633;
  assign add_540640 = sel_540637 + 8'h01;
  assign sel_540641 = array_index_540492 == array_index_537238 ? add_540640 : sel_540637;
  assign add_540644 = sel_540641 + 8'h01;
  assign sel_540645 = array_index_540492 == array_index_537244 ? add_540644 : sel_540641;
  assign add_540648 = sel_540645 + 8'h01;
  assign sel_540649 = array_index_540492 == array_index_537250 ? add_540648 : sel_540645;
  assign add_540652 = sel_540649 + 8'h01;
  assign sel_540653 = array_index_540492 == array_index_537256 ? add_540652 : sel_540649;
  assign add_540656 = sel_540653 + 8'h01;
  assign sel_540657 = array_index_540492 == array_index_537262 ? add_540656 : sel_540653;
  assign add_540660 = sel_540657 + 8'h01;
  assign sel_540661 = array_index_540492 == array_index_537268 ? add_540660 : sel_540657;
  assign add_540664 = sel_540661 + 8'h01;
  assign sel_540665 = array_index_540492 == array_index_537274 ? add_540664 : sel_540661;
  assign add_540668 = sel_540665 + 8'h01;
  assign sel_540669 = array_index_540492 == array_index_537280 ? add_540668 : sel_540665;
  assign add_540672 = sel_540669 + 8'h01;
  assign sel_540673 = array_index_540492 == array_index_537286 ? add_540672 : sel_540669;
  assign add_540676 = sel_540673 + 8'h01;
  assign sel_540677 = array_index_540492 == array_index_537292 ? add_540676 : sel_540673;
  assign add_540680 = sel_540677 + 8'h01;
  assign sel_540681 = array_index_540492 == array_index_537298 ? add_540680 : sel_540677;
  assign add_540684 = sel_540681 + 8'h01;
  assign sel_540685 = array_index_540492 == array_index_537304 ? add_540684 : sel_540681;
  assign add_540688 = sel_540685 + 8'h01;
  assign sel_540689 = array_index_540492 == array_index_537310 ? add_540688 : sel_540685;
  assign add_540692 = sel_540689 + 8'h01;
  assign sel_540693 = array_index_540492 == array_index_537316 ? add_540692 : sel_540689;
  assign add_540696 = sel_540693 + 8'h01;
  assign sel_540697 = array_index_540492 == array_index_537322 ? add_540696 : sel_540693;
  assign add_540700 = sel_540697 + 8'h01;
  assign sel_540701 = array_index_540492 == array_index_537328 ? add_540700 : sel_540697;
  assign add_540704 = sel_540701 + 8'h01;
  assign sel_540705 = array_index_540492 == array_index_537334 ? add_540704 : sel_540701;
  assign add_540708 = sel_540705 + 8'h01;
  assign sel_540709 = array_index_540492 == array_index_537340 ? add_540708 : sel_540705;
  assign add_540712 = sel_540709 + 8'h01;
  assign sel_540713 = array_index_540492 == array_index_537346 ? add_540712 : sel_540709;
  assign add_540716 = sel_540713 + 8'h01;
  assign sel_540717 = array_index_540492 == array_index_537352 ? add_540716 : sel_540713;
  assign add_540720 = sel_540717 + 8'h01;
  assign sel_540721 = array_index_540492 == array_index_537358 ? add_540720 : sel_540717;
  assign add_540724 = sel_540721 + 8'h01;
  assign sel_540725 = array_index_540492 == array_index_537364 ? add_540724 : sel_540721;
  assign add_540728 = sel_540725 + 8'h01;
  assign sel_540729 = array_index_540492 == array_index_537370 ? add_540728 : sel_540725;
  assign add_540732 = sel_540729 + 8'h01;
  assign sel_540733 = array_index_540492 == array_index_537376 ? add_540732 : sel_540729;
  assign add_540736 = sel_540733 + 8'h01;
  assign sel_540737 = array_index_540492 == array_index_537382 ? add_540736 : sel_540733;
  assign add_540740 = sel_540737 + 8'h01;
  assign sel_540741 = array_index_540492 == array_index_537388 ? add_540740 : sel_540737;
  assign add_540744 = sel_540741 + 8'h01;
  assign sel_540745 = array_index_540492 == array_index_537394 ? add_540744 : sel_540741;
  assign add_540748 = sel_540745 + 8'h01;
  assign sel_540749 = array_index_540492 == array_index_537400 ? add_540748 : sel_540745;
  assign add_540752 = sel_540749 + 8'h01;
  assign sel_540753 = array_index_540492 == array_index_537406 ? add_540752 : sel_540749;
  assign add_540756 = sel_540753 + 8'h01;
  assign sel_540757 = array_index_540492 == array_index_537412 ? add_540756 : sel_540753;
  assign add_540760 = sel_540757 + 8'h01;
  assign sel_540761 = array_index_540492 == array_index_537418 ? add_540760 : sel_540757;
  assign add_540764 = sel_540761 + 8'h01;
  assign sel_540765 = array_index_540492 == array_index_537424 ? add_540764 : sel_540761;
  assign add_540768 = sel_540765 + 8'h01;
  assign sel_540769 = array_index_540492 == array_index_537430 ? add_540768 : sel_540765;
  assign add_540772 = sel_540769 + 8'h01;
  assign sel_540773 = array_index_540492 == array_index_537436 ? add_540772 : sel_540769;
  assign add_540776 = sel_540773 + 8'h01;
  assign sel_540777 = array_index_540492 == array_index_537442 ? add_540776 : sel_540773;
  assign add_540780 = sel_540777 + 8'h01;
  assign sel_540781 = array_index_540492 == array_index_537448 ? add_540780 : sel_540777;
  assign add_540784 = sel_540781 + 8'h01;
  assign sel_540785 = array_index_540492 == array_index_537454 ? add_540784 : sel_540781;
  assign add_540788 = sel_540785 + 8'h01;
  assign sel_540789 = array_index_540492 == array_index_537460 ? add_540788 : sel_540785;
  assign add_540793 = sel_540789 + 8'h01;
  assign array_index_540794 = set1_unflattened[7'h0c];
  assign sel_540795 = array_index_540492 == array_index_537466 ? add_540793 : sel_540789;
  assign add_540798 = sel_540795 + 8'h01;
  assign sel_540799 = array_index_540794 == array_index_537012 ? add_540798 : sel_540795;
  assign add_540802 = sel_540799 + 8'h01;
  assign sel_540803 = array_index_540794 == array_index_537016 ? add_540802 : sel_540799;
  assign add_540806 = sel_540803 + 8'h01;
  assign sel_540807 = array_index_540794 == array_index_537024 ? add_540806 : sel_540803;
  assign add_540810 = sel_540807 + 8'h01;
  assign sel_540811 = array_index_540794 == array_index_537032 ? add_540810 : sel_540807;
  assign add_540814 = sel_540811 + 8'h01;
  assign sel_540815 = array_index_540794 == array_index_537040 ? add_540814 : sel_540811;
  assign add_540818 = sel_540815 + 8'h01;
  assign sel_540819 = array_index_540794 == array_index_537048 ? add_540818 : sel_540815;
  assign add_540822 = sel_540819 + 8'h01;
  assign sel_540823 = array_index_540794 == array_index_537056 ? add_540822 : sel_540819;
  assign add_540826 = sel_540823 + 8'h01;
  assign sel_540827 = array_index_540794 == array_index_537064 ? add_540826 : sel_540823;
  assign add_540830 = sel_540827 + 8'h01;
  assign sel_540831 = array_index_540794 == array_index_537070 ? add_540830 : sel_540827;
  assign add_540834 = sel_540831 + 8'h01;
  assign sel_540835 = array_index_540794 == array_index_537076 ? add_540834 : sel_540831;
  assign add_540838 = sel_540835 + 8'h01;
  assign sel_540839 = array_index_540794 == array_index_537082 ? add_540838 : sel_540835;
  assign add_540842 = sel_540839 + 8'h01;
  assign sel_540843 = array_index_540794 == array_index_537088 ? add_540842 : sel_540839;
  assign add_540846 = sel_540843 + 8'h01;
  assign sel_540847 = array_index_540794 == array_index_537094 ? add_540846 : sel_540843;
  assign add_540850 = sel_540847 + 8'h01;
  assign sel_540851 = array_index_540794 == array_index_537100 ? add_540850 : sel_540847;
  assign add_540854 = sel_540851 + 8'h01;
  assign sel_540855 = array_index_540794 == array_index_537106 ? add_540854 : sel_540851;
  assign add_540858 = sel_540855 + 8'h01;
  assign sel_540859 = array_index_540794 == array_index_537112 ? add_540858 : sel_540855;
  assign add_540862 = sel_540859 + 8'h01;
  assign sel_540863 = array_index_540794 == array_index_537118 ? add_540862 : sel_540859;
  assign add_540866 = sel_540863 + 8'h01;
  assign sel_540867 = array_index_540794 == array_index_537124 ? add_540866 : sel_540863;
  assign add_540870 = sel_540867 + 8'h01;
  assign sel_540871 = array_index_540794 == array_index_537130 ? add_540870 : sel_540867;
  assign add_540874 = sel_540871 + 8'h01;
  assign sel_540875 = array_index_540794 == array_index_537136 ? add_540874 : sel_540871;
  assign add_540878 = sel_540875 + 8'h01;
  assign sel_540879 = array_index_540794 == array_index_537142 ? add_540878 : sel_540875;
  assign add_540882 = sel_540879 + 8'h01;
  assign sel_540883 = array_index_540794 == array_index_537148 ? add_540882 : sel_540879;
  assign add_540886 = sel_540883 + 8'h01;
  assign sel_540887 = array_index_540794 == array_index_537154 ? add_540886 : sel_540883;
  assign add_540890 = sel_540887 + 8'h01;
  assign sel_540891 = array_index_540794 == array_index_537160 ? add_540890 : sel_540887;
  assign add_540894 = sel_540891 + 8'h01;
  assign sel_540895 = array_index_540794 == array_index_537166 ? add_540894 : sel_540891;
  assign add_540898 = sel_540895 + 8'h01;
  assign sel_540899 = array_index_540794 == array_index_537172 ? add_540898 : sel_540895;
  assign add_540902 = sel_540899 + 8'h01;
  assign sel_540903 = array_index_540794 == array_index_537178 ? add_540902 : sel_540899;
  assign add_540906 = sel_540903 + 8'h01;
  assign sel_540907 = array_index_540794 == array_index_537184 ? add_540906 : sel_540903;
  assign add_540910 = sel_540907 + 8'h01;
  assign sel_540911 = array_index_540794 == array_index_537190 ? add_540910 : sel_540907;
  assign add_540914 = sel_540911 + 8'h01;
  assign sel_540915 = array_index_540794 == array_index_537196 ? add_540914 : sel_540911;
  assign add_540918 = sel_540915 + 8'h01;
  assign sel_540919 = array_index_540794 == array_index_537202 ? add_540918 : sel_540915;
  assign add_540922 = sel_540919 + 8'h01;
  assign sel_540923 = array_index_540794 == array_index_537208 ? add_540922 : sel_540919;
  assign add_540926 = sel_540923 + 8'h01;
  assign sel_540927 = array_index_540794 == array_index_537214 ? add_540926 : sel_540923;
  assign add_540930 = sel_540927 + 8'h01;
  assign sel_540931 = array_index_540794 == array_index_537220 ? add_540930 : sel_540927;
  assign add_540934 = sel_540931 + 8'h01;
  assign sel_540935 = array_index_540794 == array_index_537226 ? add_540934 : sel_540931;
  assign add_540938 = sel_540935 + 8'h01;
  assign sel_540939 = array_index_540794 == array_index_537232 ? add_540938 : sel_540935;
  assign add_540942 = sel_540939 + 8'h01;
  assign sel_540943 = array_index_540794 == array_index_537238 ? add_540942 : sel_540939;
  assign add_540946 = sel_540943 + 8'h01;
  assign sel_540947 = array_index_540794 == array_index_537244 ? add_540946 : sel_540943;
  assign add_540950 = sel_540947 + 8'h01;
  assign sel_540951 = array_index_540794 == array_index_537250 ? add_540950 : sel_540947;
  assign add_540954 = sel_540951 + 8'h01;
  assign sel_540955 = array_index_540794 == array_index_537256 ? add_540954 : sel_540951;
  assign add_540958 = sel_540955 + 8'h01;
  assign sel_540959 = array_index_540794 == array_index_537262 ? add_540958 : sel_540955;
  assign add_540962 = sel_540959 + 8'h01;
  assign sel_540963 = array_index_540794 == array_index_537268 ? add_540962 : sel_540959;
  assign add_540966 = sel_540963 + 8'h01;
  assign sel_540967 = array_index_540794 == array_index_537274 ? add_540966 : sel_540963;
  assign add_540970 = sel_540967 + 8'h01;
  assign sel_540971 = array_index_540794 == array_index_537280 ? add_540970 : sel_540967;
  assign add_540974 = sel_540971 + 8'h01;
  assign sel_540975 = array_index_540794 == array_index_537286 ? add_540974 : sel_540971;
  assign add_540978 = sel_540975 + 8'h01;
  assign sel_540979 = array_index_540794 == array_index_537292 ? add_540978 : sel_540975;
  assign add_540982 = sel_540979 + 8'h01;
  assign sel_540983 = array_index_540794 == array_index_537298 ? add_540982 : sel_540979;
  assign add_540986 = sel_540983 + 8'h01;
  assign sel_540987 = array_index_540794 == array_index_537304 ? add_540986 : sel_540983;
  assign add_540990 = sel_540987 + 8'h01;
  assign sel_540991 = array_index_540794 == array_index_537310 ? add_540990 : sel_540987;
  assign add_540994 = sel_540991 + 8'h01;
  assign sel_540995 = array_index_540794 == array_index_537316 ? add_540994 : sel_540991;
  assign add_540998 = sel_540995 + 8'h01;
  assign sel_540999 = array_index_540794 == array_index_537322 ? add_540998 : sel_540995;
  assign add_541002 = sel_540999 + 8'h01;
  assign sel_541003 = array_index_540794 == array_index_537328 ? add_541002 : sel_540999;
  assign add_541006 = sel_541003 + 8'h01;
  assign sel_541007 = array_index_540794 == array_index_537334 ? add_541006 : sel_541003;
  assign add_541010 = sel_541007 + 8'h01;
  assign sel_541011 = array_index_540794 == array_index_537340 ? add_541010 : sel_541007;
  assign add_541014 = sel_541011 + 8'h01;
  assign sel_541015 = array_index_540794 == array_index_537346 ? add_541014 : sel_541011;
  assign add_541018 = sel_541015 + 8'h01;
  assign sel_541019 = array_index_540794 == array_index_537352 ? add_541018 : sel_541015;
  assign add_541022 = sel_541019 + 8'h01;
  assign sel_541023 = array_index_540794 == array_index_537358 ? add_541022 : sel_541019;
  assign add_541026 = sel_541023 + 8'h01;
  assign sel_541027 = array_index_540794 == array_index_537364 ? add_541026 : sel_541023;
  assign add_541030 = sel_541027 + 8'h01;
  assign sel_541031 = array_index_540794 == array_index_537370 ? add_541030 : sel_541027;
  assign add_541034 = sel_541031 + 8'h01;
  assign sel_541035 = array_index_540794 == array_index_537376 ? add_541034 : sel_541031;
  assign add_541038 = sel_541035 + 8'h01;
  assign sel_541039 = array_index_540794 == array_index_537382 ? add_541038 : sel_541035;
  assign add_541042 = sel_541039 + 8'h01;
  assign sel_541043 = array_index_540794 == array_index_537388 ? add_541042 : sel_541039;
  assign add_541046 = sel_541043 + 8'h01;
  assign sel_541047 = array_index_540794 == array_index_537394 ? add_541046 : sel_541043;
  assign add_541050 = sel_541047 + 8'h01;
  assign sel_541051 = array_index_540794 == array_index_537400 ? add_541050 : sel_541047;
  assign add_541054 = sel_541051 + 8'h01;
  assign sel_541055 = array_index_540794 == array_index_537406 ? add_541054 : sel_541051;
  assign add_541058 = sel_541055 + 8'h01;
  assign sel_541059 = array_index_540794 == array_index_537412 ? add_541058 : sel_541055;
  assign add_541062 = sel_541059 + 8'h01;
  assign sel_541063 = array_index_540794 == array_index_537418 ? add_541062 : sel_541059;
  assign add_541066 = sel_541063 + 8'h01;
  assign sel_541067 = array_index_540794 == array_index_537424 ? add_541066 : sel_541063;
  assign add_541070 = sel_541067 + 8'h01;
  assign sel_541071 = array_index_540794 == array_index_537430 ? add_541070 : sel_541067;
  assign add_541074 = sel_541071 + 8'h01;
  assign sel_541075 = array_index_540794 == array_index_537436 ? add_541074 : sel_541071;
  assign add_541078 = sel_541075 + 8'h01;
  assign sel_541079 = array_index_540794 == array_index_537442 ? add_541078 : sel_541075;
  assign add_541082 = sel_541079 + 8'h01;
  assign sel_541083 = array_index_540794 == array_index_537448 ? add_541082 : sel_541079;
  assign add_541086 = sel_541083 + 8'h01;
  assign sel_541087 = array_index_540794 == array_index_537454 ? add_541086 : sel_541083;
  assign add_541090 = sel_541087 + 8'h01;
  assign sel_541091 = array_index_540794 == array_index_537460 ? add_541090 : sel_541087;
  assign add_541095 = sel_541091 + 8'h01;
  assign array_index_541096 = set1_unflattened[7'h0d];
  assign sel_541097 = array_index_540794 == array_index_537466 ? add_541095 : sel_541091;
  assign add_541100 = sel_541097 + 8'h01;
  assign sel_541101 = array_index_541096 == array_index_537012 ? add_541100 : sel_541097;
  assign add_541104 = sel_541101 + 8'h01;
  assign sel_541105 = array_index_541096 == array_index_537016 ? add_541104 : sel_541101;
  assign add_541108 = sel_541105 + 8'h01;
  assign sel_541109 = array_index_541096 == array_index_537024 ? add_541108 : sel_541105;
  assign add_541112 = sel_541109 + 8'h01;
  assign sel_541113 = array_index_541096 == array_index_537032 ? add_541112 : sel_541109;
  assign add_541116 = sel_541113 + 8'h01;
  assign sel_541117 = array_index_541096 == array_index_537040 ? add_541116 : sel_541113;
  assign add_541120 = sel_541117 + 8'h01;
  assign sel_541121 = array_index_541096 == array_index_537048 ? add_541120 : sel_541117;
  assign add_541124 = sel_541121 + 8'h01;
  assign sel_541125 = array_index_541096 == array_index_537056 ? add_541124 : sel_541121;
  assign add_541128 = sel_541125 + 8'h01;
  assign sel_541129 = array_index_541096 == array_index_537064 ? add_541128 : sel_541125;
  assign add_541132 = sel_541129 + 8'h01;
  assign sel_541133 = array_index_541096 == array_index_537070 ? add_541132 : sel_541129;
  assign add_541136 = sel_541133 + 8'h01;
  assign sel_541137 = array_index_541096 == array_index_537076 ? add_541136 : sel_541133;
  assign add_541140 = sel_541137 + 8'h01;
  assign sel_541141 = array_index_541096 == array_index_537082 ? add_541140 : sel_541137;
  assign add_541144 = sel_541141 + 8'h01;
  assign sel_541145 = array_index_541096 == array_index_537088 ? add_541144 : sel_541141;
  assign add_541148 = sel_541145 + 8'h01;
  assign sel_541149 = array_index_541096 == array_index_537094 ? add_541148 : sel_541145;
  assign add_541152 = sel_541149 + 8'h01;
  assign sel_541153 = array_index_541096 == array_index_537100 ? add_541152 : sel_541149;
  assign add_541156 = sel_541153 + 8'h01;
  assign sel_541157 = array_index_541096 == array_index_537106 ? add_541156 : sel_541153;
  assign add_541160 = sel_541157 + 8'h01;
  assign sel_541161 = array_index_541096 == array_index_537112 ? add_541160 : sel_541157;
  assign add_541164 = sel_541161 + 8'h01;
  assign sel_541165 = array_index_541096 == array_index_537118 ? add_541164 : sel_541161;
  assign add_541168 = sel_541165 + 8'h01;
  assign sel_541169 = array_index_541096 == array_index_537124 ? add_541168 : sel_541165;
  assign add_541172 = sel_541169 + 8'h01;
  assign sel_541173 = array_index_541096 == array_index_537130 ? add_541172 : sel_541169;
  assign add_541176 = sel_541173 + 8'h01;
  assign sel_541177 = array_index_541096 == array_index_537136 ? add_541176 : sel_541173;
  assign add_541180 = sel_541177 + 8'h01;
  assign sel_541181 = array_index_541096 == array_index_537142 ? add_541180 : sel_541177;
  assign add_541184 = sel_541181 + 8'h01;
  assign sel_541185 = array_index_541096 == array_index_537148 ? add_541184 : sel_541181;
  assign add_541188 = sel_541185 + 8'h01;
  assign sel_541189 = array_index_541096 == array_index_537154 ? add_541188 : sel_541185;
  assign add_541192 = sel_541189 + 8'h01;
  assign sel_541193 = array_index_541096 == array_index_537160 ? add_541192 : sel_541189;
  assign add_541196 = sel_541193 + 8'h01;
  assign sel_541197 = array_index_541096 == array_index_537166 ? add_541196 : sel_541193;
  assign add_541200 = sel_541197 + 8'h01;
  assign sel_541201 = array_index_541096 == array_index_537172 ? add_541200 : sel_541197;
  assign add_541204 = sel_541201 + 8'h01;
  assign sel_541205 = array_index_541096 == array_index_537178 ? add_541204 : sel_541201;
  assign add_541208 = sel_541205 + 8'h01;
  assign sel_541209 = array_index_541096 == array_index_537184 ? add_541208 : sel_541205;
  assign add_541212 = sel_541209 + 8'h01;
  assign sel_541213 = array_index_541096 == array_index_537190 ? add_541212 : sel_541209;
  assign add_541216 = sel_541213 + 8'h01;
  assign sel_541217 = array_index_541096 == array_index_537196 ? add_541216 : sel_541213;
  assign add_541220 = sel_541217 + 8'h01;
  assign sel_541221 = array_index_541096 == array_index_537202 ? add_541220 : sel_541217;
  assign add_541224 = sel_541221 + 8'h01;
  assign sel_541225 = array_index_541096 == array_index_537208 ? add_541224 : sel_541221;
  assign add_541228 = sel_541225 + 8'h01;
  assign sel_541229 = array_index_541096 == array_index_537214 ? add_541228 : sel_541225;
  assign add_541232 = sel_541229 + 8'h01;
  assign sel_541233 = array_index_541096 == array_index_537220 ? add_541232 : sel_541229;
  assign add_541236 = sel_541233 + 8'h01;
  assign sel_541237 = array_index_541096 == array_index_537226 ? add_541236 : sel_541233;
  assign add_541240 = sel_541237 + 8'h01;
  assign sel_541241 = array_index_541096 == array_index_537232 ? add_541240 : sel_541237;
  assign add_541244 = sel_541241 + 8'h01;
  assign sel_541245 = array_index_541096 == array_index_537238 ? add_541244 : sel_541241;
  assign add_541248 = sel_541245 + 8'h01;
  assign sel_541249 = array_index_541096 == array_index_537244 ? add_541248 : sel_541245;
  assign add_541252 = sel_541249 + 8'h01;
  assign sel_541253 = array_index_541096 == array_index_537250 ? add_541252 : sel_541249;
  assign add_541256 = sel_541253 + 8'h01;
  assign sel_541257 = array_index_541096 == array_index_537256 ? add_541256 : sel_541253;
  assign add_541260 = sel_541257 + 8'h01;
  assign sel_541261 = array_index_541096 == array_index_537262 ? add_541260 : sel_541257;
  assign add_541264 = sel_541261 + 8'h01;
  assign sel_541265 = array_index_541096 == array_index_537268 ? add_541264 : sel_541261;
  assign add_541268 = sel_541265 + 8'h01;
  assign sel_541269 = array_index_541096 == array_index_537274 ? add_541268 : sel_541265;
  assign add_541272 = sel_541269 + 8'h01;
  assign sel_541273 = array_index_541096 == array_index_537280 ? add_541272 : sel_541269;
  assign add_541276 = sel_541273 + 8'h01;
  assign sel_541277 = array_index_541096 == array_index_537286 ? add_541276 : sel_541273;
  assign add_541280 = sel_541277 + 8'h01;
  assign sel_541281 = array_index_541096 == array_index_537292 ? add_541280 : sel_541277;
  assign add_541284 = sel_541281 + 8'h01;
  assign sel_541285 = array_index_541096 == array_index_537298 ? add_541284 : sel_541281;
  assign add_541288 = sel_541285 + 8'h01;
  assign sel_541289 = array_index_541096 == array_index_537304 ? add_541288 : sel_541285;
  assign add_541292 = sel_541289 + 8'h01;
  assign sel_541293 = array_index_541096 == array_index_537310 ? add_541292 : sel_541289;
  assign add_541296 = sel_541293 + 8'h01;
  assign sel_541297 = array_index_541096 == array_index_537316 ? add_541296 : sel_541293;
  assign add_541300 = sel_541297 + 8'h01;
  assign sel_541301 = array_index_541096 == array_index_537322 ? add_541300 : sel_541297;
  assign add_541304 = sel_541301 + 8'h01;
  assign sel_541305 = array_index_541096 == array_index_537328 ? add_541304 : sel_541301;
  assign add_541308 = sel_541305 + 8'h01;
  assign sel_541309 = array_index_541096 == array_index_537334 ? add_541308 : sel_541305;
  assign add_541312 = sel_541309 + 8'h01;
  assign sel_541313 = array_index_541096 == array_index_537340 ? add_541312 : sel_541309;
  assign add_541316 = sel_541313 + 8'h01;
  assign sel_541317 = array_index_541096 == array_index_537346 ? add_541316 : sel_541313;
  assign add_541320 = sel_541317 + 8'h01;
  assign sel_541321 = array_index_541096 == array_index_537352 ? add_541320 : sel_541317;
  assign add_541324 = sel_541321 + 8'h01;
  assign sel_541325 = array_index_541096 == array_index_537358 ? add_541324 : sel_541321;
  assign add_541328 = sel_541325 + 8'h01;
  assign sel_541329 = array_index_541096 == array_index_537364 ? add_541328 : sel_541325;
  assign add_541332 = sel_541329 + 8'h01;
  assign sel_541333 = array_index_541096 == array_index_537370 ? add_541332 : sel_541329;
  assign add_541336 = sel_541333 + 8'h01;
  assign sel_541337 = array_index_541096 == array_index_537376 ? add_541336 : sel_541333;
  assign add_541340 = sel_541337 + 8'h01;
  assign sel_541341 = array_index_541096 == array_index_537382 ? add_541340 : sel_541337;
  assign add_541344 = sel_541341 + 8'h01;
  assign sel_541345 = array_index_541096 == array_index_537388 ? add_541344 : sel_541341;
  assign add_541348 = sel_541345 + 8'h01;
  assign sel_541349 = array_index_541096 == array_index_537394 ? add_541348 : sel_541345;
  assign add_541352 = sel_541349 + 8'h01;
  assign sel_541353 = array_index_541096 == array_index_537400 ? add_541352 : sel_541349;
  assign add_541356 = sel_541353 + 8'h01;
  assign sel_541357 = array_index_541096 == array_index_537406 ? add_541356 : sel_541353;
  assign add_541360 = sel_541357 + 8'h01;
  assign sel_541361 = array_index_541096 == array_index_537412 ? add_541360 : sel_541357;
  assign add_541364 = sel_541361 + 8'h01;
  assign sel_541365 = array_index_541096 == array_index_537418 ? add_541364 : sel_541361;
  assign add_541368 = sel_541365 + 8'h01;
  assign sel_541369 = array_index_541096 == array_index_537424 ? add_541368 : sel_541365;
  assign add_541372 = sel_541369 + 8'h01;
  assign sel_541373 = array_index_541096 == array_index_537430 ? add_541372 : sel_541369;
  assign add_541376 = sel_541373 + 8'h01;
  assign sel_541377 = array_index_541096 == array_index_537436 ? add_541376 : sel_541373;
  assign add_541380 = sel_541377 + 8'h01;
  assign sel_541381 = array_index_541096 == array_index_537442 ? add_541380 : sel_541377;
  assign add_541384 = sel_541381 + 8'h01;
  assign sel_541385 = array_index_541096 == array_index_537448 ? add_541384 : sel_541381;
  assign add_541388 = sel_541385 + 8'h01;
  assign sel_541389 = array_index_541096 == array_index_537454 ? add_541388 : sel_541385;
  assign add_541392 = sel_541389 + 8'h01;
  assign sel_541393 = array_index_541096 == array_index_537460 ? add_541392 : sel_541389;
  assign add_541397 = sel_541393 + 8'h01;
  assign array_index_541398 = set1_unflattened[7'h0e];
  assign sel_541399 = array_index_541096 == array_index_537466 ? add_541397 : sel_541393;
  assign add_541402 = sel_541399 + 8'h01;
  assign sel_541403 = array_index_541398 == array_index_537012 ? add_541402 : sel_541399;
  assign add_541406 = sel_541403 + 8'h01;
  assign sel_541407 = array_index_541398 == array_index_537016 ? add_541406 : sel_541403;
  assign add_541410 = sel_541407 + 8'h01;
  assign sel_541411 = array_index_541398 == array_index_537024 ? add_541410 : sel_541407;
  assign add_541414 = sel_541411 + 8'h01;
  assign sel_541415 = array_index_541398 == array_index_537032 ? add_541414 : sel_541411;
  assign add_541418 = sel_541415 + 8'h01;
  assign sel_541419 = array_index_541398 == array_index_537040 ? add_541418 : sel_541415;
  assign add_541422 = sel_541419 + 8'h01;
  assign sel_541423 = array_index_541398 == array_index_537048 ? add_541422 : sel_541419;
  assign add_541426 = sel_541423 + 8'h01;
  assign sel_541427 = array_index_541398 == array_index_537056 ? add_541426 : sel_541423;
  assign add_541430 = sel_541427 + 8'h01;
  assign sel_541431 = array_index_541398 == array_index_537064 ? add_541430 : sel_541427;
  assign add_541434 = sel_541431 + 8'h01;
  assign sel_541435 = array_index_541398 == array_index_537070 ? add_541434 : sel_541431;
  assign add_541438 = sel_541435 + 8'h01;
  assign sel_541439 = array_index_541398 == array_index_537076 ? add_541438 : sel_541435;
  assign add_541442 = sel_541439 + 8'h01;
  assign sel_541443 = array_index_541398 == array_index_537082 ? add_541442 : sel_541439;
  assign add_541446 = sel_541443 + 8'h01;
  assign sel_541447 = array_index_541398 == array_index_537088 ? add_541446 : sel_541443;
  assign add_541450 = sel_541447 + 8'h01;
  assign sel_541451 = array_index_541398 == array_index_537094 ? add_541450 : sel_541447;
  assign add_541454 = sel_541451 + 8'h01;
  assign sel_541455 = array_index_541398 == array_index_537100 ? add_541454 : sel_541451;
  assign add_541458 = sel_541455 + 8'h01;
  assign sel_541459 = array_index_541398 == array_index_537106 ? add_541458 : sel_541455;
  assign add_541462 = sel_541459 + 8'h01;
  assign sel_541463 = array_index_541398 == array_index_537112 ? add_541462 : sel_541459;
  assign add_541466 = sel_541463 + 8'h01;
  assign sel_541467 = array_index_541398 == array_index_537118 ? add_541466 : sel_541463;
  assign add_541470 = sel_541467 + 8'h01;
  assign sel_541471 = array_index_541398 == array_index_537124 ? add_541470 : sel_541467;
  assign add_541474 = sel_541471 + 8'h01;
  assign sel_541475 = array_index_541398 == array_index_537130 ? add_541474 : sel_541471;
  assign add_541478 = sel_541475 + 8'h01;
  assign sel_541479 = array_index_541398 == array_index_537136 ? add_541478 : sel_541475;
  assign add_541482 = sel_541479 + 8'h01;
  assign sel_541483 = array_index_541398 == array_index_537142 ? add_541482 : sel_541479;
  assign add_541486 = sel_541483 + 8'h01;
  assign sel_541487 = array_index_541398 == array_index_537148 ? add_541486 : sel_541483;
  assign add_541490 = sel_541487 + 8'h01;
  assign sel_541491 = array_index_541398 == array_index_537154 ? add_541490 : sel_541487;
  assign add_541494 = sel_541491 + 8'h01;
  assign sel_541495 = array_index_541398 == array_index_537160 ? add_541494 : sel_541491;
  assign add_541498 = sel_541495 + 8'h01;
  assign sel_541499 = array_index_541398 == array_index_537166 ? add_541498 : sel_541495;
  assign add_541502 = sel_541499 + 8'h01;
  assign sel_541503 = array_index_541398 == array_index_537172 ? add_541502 : sel_541499;
  assign add_541506 = sel_541503 + 8'h01;
  assign sel_541507 = array_index_541398 == array_index_537178 ? add_541506 : sel_541503;
  assign add_541510 = sel_541507 + 8'h01;
  assign sel_541511 = array_index_541398 == array_index_537184 ? add_541510 : sel_541507;
  assign add_541514 = sel_541511 + 8'h01;
  assign sel_541515 = array_index_541398 == array_index_537190 ? add_541514 : sel_541511;
  assign add_541518 = sel_541515 + 8'h01;
  assign sel_541519 = array_index_541398 == array_index_537196 ? add_541518 : sel_541515;
  assign add_541522 = sel_541519 + 8'h01;
  assign sel_541523 = array_index_541398 == array_index_537202 ? add_541522 : sel_541519;
  assign add_541526 = sel_541523 + 8'h01;
  assign sel_541527 = array_index_541398 == array_index_537208 ? add_541526 : sel_541523;
  assign add_541530 = sel_541527 + 8'h01;
  assign sel_541531 = array_index_541398 == array_index_537214 ? add_541530 : sel_541527;
  assign add_541534 = sel_541531 + 8'h01;
  assign sel_541535 = array_index_541398 == array_index_537220 ? add_541534 : sel_541531;
  assign add_541538 = sel_541535 + 8'h01;
  assign sel_541539 = array_index_541398 == array_index_537226 ? add_541538 : sel_541535;
  assign add_541542 = sel_541539 + 8'h01;
  assign sel_541543 = array_index_541398 == array_index_537232 ? add_541542 : sel_541539;
  assign add_541546 = sel_541543 + 8'h01;
  assign sel_541547 = array_index_541398 == array_index_537238 ? add_541546 : sel_541543;
  assign add_541550 = sel_541547 + 8'h01;
  assign sel_541551 = array_index_541398 == array_index_537244 ? add_541550 : sel_541547;
  assign add_541554 = sel_541551 + 8'h01;
  assign sel_541555 = array_index_541398 == array_index_537250 ? add_541554 : sel_541551;
  assign add_541558 = sel_541555 + 8'h01;
  assign sel_541559 = array_index_541398 == array_index_537256 ? add_541558 : sel_541555;
  assign add_541562 = sel_541559 + 8'h01;
  assign sel_541563 = array_index_541398 == array_index_537262 ? add_541562 : sel_541559;
  assign add_541566 = sel_541563 + 8'h01;
  assign sel_541567 = array_index_541398 == array_index_537268 ? add_541566 : sel_541563;
  assign add_541570 = sel_541567 + 8'h01;
  assign sel_541571 = array_index_541398 == array_index_537274 ? add_541570 : sel_541567;
  assign add_541574 = sel_541571 + 8'h01;
  assign sel_541575 = array_index_541398 == array_index_537280 ? add_541574 : sel_541571;
  assign add_541578 = sel_541575 + 8'h01;
  assign sel_541579 = array_index_541398 == array_index_537286 ? add_541578 : sel_541575;
  assign add_541582 = sel_541579 + 8'h01;
  assign sel_541583 = array_index_541398 == array_index_537292 ? add_541582 : sel_541579;
  assign add_541586 = sel_541583 + 8'h01;
  assign sel_541587 = array_index_541398 == array_index_537298 ? add_541586 : sel_541583;
  assign add_541590 = sel_541587 + 8'h01;
  assign sel_541591 = array_index_541398 == array_index_537304 ? add_541590 : sel_541587;
  assign add_541594 = sel_541591 + 8'h01;
  assign sel_541595 = array_index_541398 == array_index_537310 ? add_541594 : sel_541591;
  assign add_541598 = sel_541595 + 8'h01;
  assign sel_541599 = array_index_541398 == array_index_537316 ? add_541598 : sel_541595;
  assign add_541602 = sel_541599 + 8'h01;
  assign sel_541603 = array_index_541398 == array_index_537322 ? add_541602 : sel_541599;
  assign add_541606 = sel_541603 + 8'h01;
  assign sel_541607 = array_index_541398 == array_index_537328 ? add_541606 : sel_541603;
  assign add_541610 = sel_541607 + 8'h01;
  assign sel_541611 = array_index_541398 == array_index_537334 ? add_541610 : sel_541607;
  assign add_541614 = sel_541611 + 8'h01;
  assign sel_541615 = array_index_541398 == array_index_537340 ? add_541614 : sel_541611;
  assign add_541618 = sel_541615 + 8'h01;
  assign sel_541619 = array_index_541398 == array_index_537346 ? add_541618 : sel_541615;
  assign add_541622 = sel_541619 + 8'h01;
  assign sel_541623 = array_index_541398 == array_index_537352 ? add_541622 : sel_541619;
  assign add_541626 = sel_541623 + 8'h01;
  assign sel_541627 = array_index_541398 == array_index_537358 ? add_541626 : sel_541623;
  assign add_541630 = sel_541627 + 8'h01;
  assign sel_541631 = array_index_541398 == array_index_537364 ? add_541630 : sel_541627;
  assign add_541634 = sel_541631 + 8'h01;
  assign sel_541635 = array_index_541398 == array_index_537370 ? add_541634 : sel_541631;
  assign add_541638 = sel_541635 + 8'h01;
  assign sel_541639 = array_index_541398 == array_index_537376 ? add_541638 : sel_541635;
  assign add_541642 = sel_541639 + 8'h01;
  assign sel_541643 = array_index_541398 == array_index_537382 ? add_541642 : sel_541639;
  assign add_541646 = sel_541643 + 8'h01;
  assign sel_541647 = array_index_541398 == array_index_537388 ? add_541646 : sel_541643;
  assign add_541650 = sel_541647 + 8'h01;
  assign sel_541651 = array_index_541398 == array_index_537394 ? add_541650 : sel_541647;
  assign add_541654 = sel_541651 + 8'h01;
  assign sel_541655 = array_index_541398 == array_index_537400 ? add_541654 : sel_541651;
  assign add_541658 = sel_541655 + 8'h01;
  assign sel_541659 = array_index_541398 == array_index_537406 ? add_541658 : sel_541655;
  assign add_541662 = sel_541659 + 8'h01;
  assign sel_541663 = array_index_541398 == array_index_537412 ? add_541662 : sel_541659;
  assign add_541666 = sel_541663 + 8'h01;
  assign sel_541667 = array_index_541398 == array_index_537418 ? add_541666 : sel_541663;
  assign add_541670 = sel_541667 + 8'h01;
  assign sel_541671 = array_index_541398 == array_index_537424 ? add_541670 : sel_541667;
  assign add_541674 = sel_541671 + 8'h01;
  assign sel_541675 = array_index_541398 == array_index_537430 ? add_541674 : sel_541671;
  assign add_541678 = sel_541675 + 8'h01;
  assign sel_541679 = array_index_541398 == array_index_537436 ? add_541678 : sel_541675;
  assign add_541682 = sel_541679 + 8'h01;
  assign sel_541683 = array_index_541398 == array_index_537442 ? add_541682 : sel_541679;
  assign add_541686 = sel_541683 + 8'h01;
  assign sel_541687 = array_index_541398 == array_index_537448 ? add_541686 : sel_541683;
  assign add_541690 = sel_541687 + 8'h01;
  assign sel_541691 = array_index_541398 == array_index_537454 ? add_541690 : sel_541687;
  assign add_541694 = sel_541691 + 8'h01;
  assign sel_541695 = array_index_541398 == array_index_537460 ? add_541694 : sel_541691;
  assign add_541699 = sel_541695 + 8'h01;
  assign array_index_541700 = set1_unflattened[7'h0f];
  assign sel_541701 = array_index_541398 == array_index_537466 ? add_541699 : sel_541695;
  assign add_541704 = sel_541701 + 8'h01;
  assign sel_541705 = array_index_541700 == array_index_537012 ? add_541704 : sel_541701;
  assign add_541708 = sel_541705 + 8'h01;
  assign sel_541709 = array_index_541700 == array_index_537016 ? add_541708 : sel_541705;
  assign add_541712 = sel_541709 + 8'h01;
  assign sel_541713 = array_index_541700 == array_index_537024 ? add_541712 : sel_541709;
  assign add_541716 = sel_541713 + 8'h01;
  assign sel_541717 = array_index_541700 == array_index_537032 ? add_541716 : sel_541713;
  assign add_541720 = sel_541717 + 8'h01;
  assign sel_541721 = array_index_541700 == array_index_537040 ? add_541720 : sel_541717;
  assign add_541724 = sel_541721 + 8'h01;
  assign sel_541725 = array_index_541700 == array_index_537048 ? add_541724 : sel_541721;
  assign add_541728 = sel_541725 + 8'h01;
  assign sel_541729 = array_index_541700 == array_index_537056 ? add_541728 : sel_541725;
  assign add_541732 = sel_541729 + 8'h01;
  assign sel_541733 = array_index_541700 == array_index_537064 ? add_541732 : sel_541729;
  assign add_541736 = sel_541733 + 8'h01;
  assign sel_541737 = array_index_541700 == array_index_537070 ? add_541736 : sel_541733;
  assign add_541740 = sel_541737 + 8'h01;
  assign sel_541741 = array_index_541700 == array_index_537076 ? add_541740 : sel_541737;
  assign add_541744 = sel_541741 + 8'h01;
  assign sel_541745 = array_index_541700 == array_index_537082 ? add_541744 : sel_541741;
  assign add_541748 = sel_541745 + 8'h01;
  assign sel_541749 = array_index_541700 == array_index_537088 ? add_541748 : sel_541745;
  assign add_541752 = sel_541749 + 8'h01;
  assign sel_541753 = array_index_541700 == array_index_537094 ? add_541752 : sel_541749;
  assign add_541756 = sel_541753 + 8'h01;
  assign sel_541757 = array_index_541700 == array_index_537100 ? add_541756 : sel_541753;
  assign add_541760 = sel_541757 + 8'h01;
  assign sel_541761 = array_index_541700 == array_index_537106 ? add_541760 : sel_541757;
  assign add_541764 = sel_541761 + 8'h01;
  assign sel_541765 = array_index_541700 == array_index_537112 ? add_541764 : sel_541761;
  assign add_541768 = sel_541765 + 8'h01;
  assign sel_541769 = array_index_541700 == array_index_537118 ? add_541768 : sel_541765;
  assign add_541772 = sel_541769 + 8'h01;
  assign sel_541773 = array_index_541700 == array_index_537124 ? add_541772 : sel_541769;
  assign add_541776 = sel_541773 + 8'h01;
  assign sel_541777 = array_index_541700 == array_index_537130 ? add_541776 : sel_541773;
  assign add_541780 = sel_541777 + 8'h01;
  assign sel_541781 = array_index_541700 == array_index_537136 ? add_541780 : sel_541777;
  assign add_541784 = sel_541781 + 8'h01;
  assign sel_541785 = array_index_541700 == array_index_537142 ? add_541784 : sel_541781;
  assign add_541788 = sel_541785 + 8'h01;
  assign sel_541789 = array_index_541700 == array_index_537148 ? add_541788 : sel_541785;
  assign add_541792 = sel_541789 + 8'h01;
  assign sel_541793 = array_index_541700 == array_index_537154 ? add_541792 : sel_541789;
  assign add_541796 = sel_541793 + 8'h01;
  assign sel_541797 = array_index_541700 == array_index_537160 ? add_541796 : sel_541793;
  assign add_541800 = sel_541797 + 8'h01;
  assign sel_541801 = array_index_541700 == array_index_537166 ? add_541800 : sel_541797;
  assign add_541804 = sel_541801 + 8'h01;
  assign sel_541805 = array_index_541700 == array_index_537172 ? add_541804 : sel_541801;
  assign add_541808 = sel_541805 + 8'h01;
  assign sel_541809 = array_index_541700 == array_index_537178 ? add_541808 : sel_541805;
  assign add_541812 = sel_541809 + 8'h01;
  assign sel_541813 = array_index_541700 == array_index_537184 ? add_541812 : sel_541809;
  assign add_541816 = sel_541813 + 8'h01;
  assign sel_541817 = array_index_541700 == array_index_537190 ? add_541816 : sel_541813;
  assign add_541820 = sel_541817 + 8'h01;
  assign sel_541821 = array_index_541700 == array_index_537196 ? add_541820 : sel_541817;
  assign add_541824 = sel_541821 + 8'h01;
  assign sel_541825 = array_index_541700 == array_index_537202 ? add_541824 : sel_541821;
  assign add_541828 = sel_541825 + 8'h01;
  assign sel_541829 = array_index_541700 == array_index_537208 ? add_541828 : sel_541825;
  assign add_541832 = sel_541829 + 8'h01;
  assign sel_541833 = array_index_541700 == array_index_537214 ? add_541832 : sel_541829;
  assign add_541836 = sel_541833 + 8'h01;
  assign sel_541837 = array_index_541700 == array_index_537220 ? add_541836 : sel_541833;
  assign add_541840 = sel_541837 + 8'h01;
  assign sel_541841 = array_index_541700 == array_index_537226 ? add_541840 : sel_541837;
  assign add_541844 = sel_541841 + 8'h01;
  assign sel_541845 = array_index_541700 == array_index_537232 ? add_541844 : sel_541841;
  assign add_541848 = sel_541845 + 8'h01;
  assign sel_541849 = array_index_541700 == array_index_537238 ? add_541848 : sel_541845;
  assign add_541852 = sel_541849 + 8'h01;
  assign sel_541853 = array_index_541700 == array_index_537244 ? add_541852 : sel_541849;
  assign add_541856 = sel_541853 + 8'h01;
  assign sel_541857 = array_index_541700 == array_index_537250 ? add_541856 : sel_541853;
  assign add_541860 = sel_541857 + 8'h01;
  assign sel_541861 = array_index_541700 == array_index_537256 ? add_541860 : sel_541857;
  assign add_541864 = sel_541861 + 8'h01;
  assign sel_541865 = array_index_541700 == array_index_537262 ? add_541864 : sel_541861;
  assign add_541868 = sel_541865 + 8'h01;
  assign sel_541869 = array_index_541700 == array_index_537268 ? add_541868 : sel_541865;
  assign add_541872 = sel_541869 + 8'h01;
  assign sel_541873 = array_index_541700 == array_index_537274 ? add_541872 : sel_541869;
  assign add_541876 = sel_541873 + 8'h01;
  assign sel_541877 = array_index_541700 == array_index_537280 ? add_541876 : sel_541873;
  assign add_541880 = sel_541877 + 8'h01;
  assign sel_541881 = array_index_541700 == array_index_537286 ? add_541880 : sel_541877;
  assign add_541884 = sel_541881 + 8'h01;
  assign sel_541885 = array_index_541700 == array_index_537292 ? add_541884 : sel_541881;
  assign add_541888 = sel_541885 + 8'h01;
  assign sel_541889 = array_index_541700 == array_index_537298 ? add_541888 : sel_541885;
  assign add_541892 = sel_541889 + 8'h01;
  assign sel_541893 = array_index_541700 == array_index_537304 ? add_541892 : sel_541889;
  assign add_541896 = sel_541893 + 8'h01;
  assign sel_541897 = array_index_541700 == array_index_537310 ? add_541896 : sel_541893;
  assign add_541900 = sel_541897 + 8'h01;
  assign sel_541901 = array_index_541700 == array_index_537316 ? add_541900 : sel_541897;
  assign add_541904 = sel_541901 + 8'h01;
  assign sel_541905 = array_index_541700 == array_index_537322 ? add_541904 : sel_541901;
  assign add_541908 = sel_541905 + 8'h01;
  assign sel_541909 = array_index_541700 == array_index_537328 ? add_541908 : sel_541905;
  assign add_541912 = sel_541909 + 8'h01;
  assign sel_541913 = array_index_541700 == array_index_537334 ? add_541912 : sel_541909;
  assign add_541916 = sel_541913 + 8'h01;
  assign sel_541917 = array_index_541700 == array_index_537340 ? add_541916 : sel_541913;
  assign add_541920 = sel_541917 + 8'h01;
  assign sel_541921 = array_index_541700 == array_index_537346 ? add_541920 : sel_541917;
  assign add_541924 = sel_541921 + 8'h01;
  assign sel_541925 = array_index_541700 == array_index_537352 ? add_541924 : sel_541921;
  assign add_541928 = sel_541925 + 8'h01;
  assign sel_541929 = array_index_541700 == array_index_537358 ? add_541928 : sel_541925;
  assign add_541932 = sel_541929 + 8'h01;
  assign sel_541933 = array_index_541700 == array_index_537364 ? add_541932 : sel_541929;
  assign add_541936 = sel_541933 + 8'h01;
  assign sel_541937 = array_index_541700 == array_index_537370 ? add_541936 : sel_541933;
  assign add_541940 = sel_541937 + 8'h01;
  assign sel_541941 = array_index_541700 == array_index_537376 ? add_541940 : sel_541937;
  assign add_541944 = sel_541941 + 8'h01;
  assign sel_541945 = array_index_541700 == array_index_537382 ? add_541944 : sel_541941;
  assign add_541948 = sel_541945 + 8'h01;
  assign sel_541949 = array_index_541700 == array_index_537388 ? add_541948 : sel_541945;
  assign add_541952 = sel_541949 + 8'h01;
  assign sel_541953 = array_index_541700 == array_index_537394 ? add_541952 : sel_541949;
  assign add_541956 = sel_541953 + 8'h01;
  assign sel_541957 = array_index_541700 == array_index_537400 ? add_541956 : sel_541953;
  assign add_541960 = sel_541957 + 8'h01;
  assign sel_541961 = array_index_541700 == array_index_537406 ? add_541960 : sel_541957;
  assign add_541964 = sel_541961 + 8'h01;
  assign sel_541965 = array_index_541700 == array_index_537412 ? add_541964 : sel_541961;
  assign add_541968 = sel_541965 + 8'h01;
  assign sel_541969 = array_index_541700 == array_index_537418 ? add_541968 : sel_541965;
  assign add_541972 = sel_541969 + 8'h01;
  assign sel_541973 = array_index_541700 == array_index_537424 ? add_541972 : sel_541969;
  assign add_541976 = sel_541973 + 8'h01;
  assign sel_541977 = array_index_541700 == array_index_537430 ? add_541976 : sel_541973;
  assign add_541980 = sel_541977 + 8'h01;
  assign sel_541981 = array_index_541700 == array_index_537436 ? add_541980 : sel_541977;
  assign add_541984 = sel_541981 + 8'h01;
  assign sel_541985 = array_index_541700 == array_index_537442 ? add_541984 : sel_541981;
  assign add_541988 = sel_541985 + 8'h01;
  assign sel_541989 = array_index_541700 == array_index_537448 ? add_541988 : sel_541985;
  assign add_541992 = sel_541989 + 8'h01;
  assign sel_541993 = array_index_541700 == array_index_537454 ? add_541992 : sel_541989;
  assign add_541996 = sel_541993 + 8'h01;
  assign sel_541997 = array_index_541700 == array_index_537460 ? add_541996 : sel_541993;
  assign add_542001 = sel_541997 + 8'h01;
  assign array_index_542002 = set1_unflattened[7'h10];
  assign sel_542003 = array_index_541700 == array_index_537466 ? add_542001 : sel_541997;
  assign add_542006 = sel_542003 + 8'h01;
  assign sel_542007 = array_index_542002 == array_index_537012 ? add_542006 : sel_542003;
  assign add_542010 = sel_542007 + 8'h01;
  assign sel_542011 = array_index_542002 == array_index_537016 ? add_542010 : sel_542007;
  assign add_542014 = sel_542011 + 8'h01;
  assign sel_542015 = array_index_542002 == array_index_537024 ? add_542014 : sel_542011;
  assign add_542018 = sel_542015 + 8'h01;
  assign sel_542019 = array_index_542002 == array_index_537032 ? add_542018 : sel_542015;
  assign add_542022 = sel_542019 + 8'h01;
  assign sel_542023 = array_index_542002 == array_index_537040 ? add_542022 : sel_542019;
  assign add_542026 = sel_542023 + 8'h01;
  assign sel_542027 = array_index_542002 == array_index_537048 ? add_542026 : sel_542023;
  assign add_542030 = sel_542027 + 8'h01;
  assign sel_542031 = array_index_542002 == array_index_537056 ? add_542030 : sel_542027;
  assign add_542034 = sel_542031 + 8'h01;
  assign sel_542035 = array_index_542002 == array_index_537064 ? add_542034 : sel_542031;
  assign add_542038 = sel_542035 + 8'h01;
  assign sel_542039 = array_index_542002 == array_index_537070 ? add_542038 : sel_542035;
  assign add_542042 = sel_542039 + 8'h01;
  assign sel_542043 = array_index_542002 == array_index_537076 ? add_542042 : sel_542039;
  assign add_542046 = sel_542043 + 8'h01;
  assign sel_542047 = array_index_542002 == array_index_537082 ? add_542046 : sel_542043;
  assign add_542050 = sel_542047 + 8'h01;
  assign sel_542051 = array_index_542002 == array_index_537088 ? add_542050 : sel_542047;
  assign add_542054 = sel_542051 + 8'h01;
  assign sel_542055 = array_index_542002 == array_index_537094 ? add_542054 : sel_542051;
  assign add_542058 = sel_542055 + 8'h01;
  assign sel_542059 = array_index_542002 == array_index_537100 ? add_542058 : sel_542055;
  assign add_542062 = sel_542059 + 8'h01;
  assign sel_542063 = array_index_542002 == array_index_537106 ? add_542062 : sel_542059;
  assign add_542066 = sel_542063 + 8'h01;
  assign sel_542067 = array_index_542002 == array_index_537112 ? add_542066 : sel_542063;
  assign add_542070 = sel_542067 + 8'h01;
  assign sel_542071 = array_index_542002 == array_index_537118 ? add_542070 : sel_542067;
  assign add_542074 = sel_542071 + 8'h01;
  assign sel_542075 = array_index_542002 == array_index_537124 ? add_542074 : sel_542071;
  assign add_542078 = sel_542075 + 8'h01;
  assign sel_542079 = array_index_542002 == array_index_537130 ? add_542078 : sel_542075;
  assign add_542082 = sel_542079 + 8'h01;
  assign sel_542083 = array_index_542002 == array_index_537136 ? add_542082 : sel_542079;
  assign add_542086 = sel_542083 + 8'h01;
  assign sel_542087 = array_index_542002 == array_index_537142 ? add_542086 : sel_542083;
  assign add_542090 = sel_542087 + 8'h01;
  assign sel_542091 = array_index_542002 == array_index_537148 ? add_542090 : sel_542087;
  assign add_542094 = sel_542091 + 8'h01;
  assign sel_542095 = array_index_542002 == array_index_537154 ? add_542094 : sel_542091;
  assign add_542098 = sel_542095 + 8'h01;
  assign sel_542099 = array_index_542002 == array_index_537160 ? add_542098 : sel_542095;
  assign add_542102 = sel_542099 + 8'h01;
  assign sel_542103 = array_index_542002 == array_index_537166 ? add_542102 : sel_542099;
  assign add_542106 = sel_542103 + 8'h01;
  assign sel_542107 = array_index_542002 == array_index_537172 ? add_542106 : sel_542103;
  assign add_542110 = sel_542107 + 8'h01;
  assign sel_542111 = array_index_542002 == array_index_537178 ? add_542110 : sel_542107;
  assign add_542114 = sel_542111 + 8'h01;
  assign sel_542115 = array_index_542002 == array_index_537184 ? add_542114 : sel_542111;
  assign add_542118 = sel_542115 + 8'h01;
  assign sel_542119 = array_index_542002 == array_index_537190 ? add_542118 : sel_542115;
  assign add_542122 = sel_542119 + 8'h01;
  assign sel_542123 = array_index_542002 == array_index_537196 ? add_542122 : sel_542119;
  assign add_542126 = sel_542123 + 8'h01;
  assign sel_542127 = array_index_542002 == array_index_537202 ? add_542126 : sel_542123;
  assign add_542130 = sel_542127 + 8'h01;
  assign sel_542131 = array_index_542002 == array_index_537208 ? add_542130 : sel_542127;
  assign add_542134 = sel_542131 + 8'h01;
  assign sel_542135 = array_index_542002 == array_index_537214 ? add_542134 : sel_542131;
  assign add_542138 = sel_542135 + 8'h01;
  assign sel_542139 = array_index_542002 == array_index_537220 ? add_542138 : sel_542135;
  assign add_542142 = sel_542139 + 8'h01;
  assign sel_542143 = array_index_542002 == array_index_537226 ? add_542142 : sel_542139;
  assign add_542146 = sel_542143 + 8'h01;
  assign sel_542147 = array_index_542002 == array_index_537232 ? add_542146 : sel_542143;
  assign add_542150 = sel_542147 + 8'h01;
  assign sel_542151 = array_index_542002 == array_index_537238 ? add_542150 : sel_542147;
  assign add_542154 = sel_542151 + 8'h01;
  assign sel_542155 = array_index_542002 == array_index_537244 ? add_542154 : sel_542151;
  assign add_542158 = sel_542155 + 8'h01;
  assign sel_542159 = array_index_542002 == array_index_537250 ? add_542158 : sel_542155;
  assign add_542162 = sel_542159 + 8'h01;
  assign sel_542163 = array_index_542002 == array_index_537256 ? add_542162 : sel_542159;
  assign add_542166 = sel_542163 + 8'h01;
  assign sel_542167 = array_index_542002 == array_index_537262 ? add_542166 : sel_542163;
  assign add_542170 = sel_542167 + 8'h01;
  assign sel_542171 = array_index_542002 == array_index_537268 ? add_542170 : sel_542167;
  assign add_542174 = sel_542171 + 8'h01;
  assign sel_542175 = array_index_542002 == array_index_537274 ? add_542174 : sel_542171;
  assign add_542178 = sel_542175 + 8'h01;
  assign sel_542179 = array_index_542002 == array_index_537280 ? add_542178 : sel_542175;
  assign add_542182 = sel_542179 + 8'h01;
  assign sel_542183 = array_index_542002 == array_index_537286 ? add_542182 : sel_542179;
  assign add_542186 = sel_542183 + 8'h01;
  assign sel_542187 = array_index_542002 == array_index_537292 ? add_542186 : sel_542183;
  assign add_542190 = sel_542187 + 8'h01;
  assign sel_542191 = array_index_542002 == array_index_537298 ? add_542190 : sel_542187;
  assign add_542194 = sel_542191 + 8'h01;
  assign sel_542195 = array_index_542002 == array_index_537304 ? add_542194 : sel_542191;
  assign add_542198 = sel_542195 + 8'h01;
  assign sel_542199 = array_index_542002 == array_index_537310 ? add_542198 : sel_542195;
  assign add_542202 = sel_542199 + 8'h01;
  assign sel_542203 = array_index_542002 == array_index_537316 ? add_542202 : sel_542199;
  assign add_542206 = sel_542203 + 8'h01;
  assign sel_542207 = array_index_542002 == array_index_537322 ? add_542206 : sel_542203;
  assign add_542210 = sel_542207 + 8'h01;
  assign sel_542211 = array_index_542002 == array_index_537328 ? add_542210 : sel_542207;
  assign add_542214 = sel_542211 + 8'h01;
  assign sel_542215 = array_index_542002 == array_index_537334 ? add_542214 : sel_542211;
  assign add_542218 = sel_542215 + 8'h01;
  assign sel_542219 = array_index_542002 == array_index_537340 ? add_542218 : sel_542215;
  assign add_542222 = sel_542219 + 8'h01;
  assign sel_542223 = array_index_542002 == array_index_537346 ? add_542222 : sel_542219;
  assign add_542226 = sel_542223 + 8'h01;
  assign sel_542227 = array_index_542002 == array_index_537352 ? add_542226 : sel_542223;
  assign add_542230 = sel_542227 + 8'h01;
  assign sel_542231 = array_index_542002 == array_index_537358 ? add_542230 : sel_542227;
  assign add_542234 = sel_542231 + 8'h01;
  assign sel_542235 = array_index_542002 == array_index_537364 ? add_542234 : sel_542231;
  assign add_542238 = sel_542235 + 8'h01;
  assign sel_542239 = array_index_542002 == array_index_537370 ? add_542238 : sel_542235;
  assign add_542242 = sel_542239 + 8'h01;
  assign sel_542243 = array_index_542002 == array_index_537376 ? add_542242 : sel_542239;
  assign add_542246 = sel_542243 + 8'h01;
  assign sel_542247 = array_index_542002 == array_index_537382 ? add_542246 : sel_542243;
  assign add_542250 = sel_542247 + 8'h01;
  assign sel_542251 = array_index_542002 == array_index_537388 ? add_542250 : sel_542247;
  assign add_542254 = sel_542251 + 8'h01;
  assign sel_542255 = array_index_542002 == array_index_537394 ? add_542254 : sel_542251;
  assign add_542258 = sel_542255 + 8'h01;
  assign sel_542259 = array_index_542002 == array_index_537400 ? add_542258 : sel_542255;
  assign add_542262 = sel_542259 + 8'h01;
  assign sel_542263 = array_index_542002 == array_index_537406 ? add_542262 : sel_542259;
  assign add_542266 = sel_542263 + 8'h01;
  assign sel_542267 = array_index_542002 == array_index_537412 ? add_542266 : sel_542263;
  assign add_542270 = sel_542267 + 8'h01;
  assign sel_542271 = array_index_542002 == array_index_537418 ? add_542270 : sel_542267;
  assign add_542274 = sel_542271 + 8'h01;
  assign sel_542275 = array_index_542002 == array_index_537424 ? add_542274 : sel_542271;
  assign add_542278 = sel_542275 + 8'h01;
  assign sel_542279 = array_index_542002 == array_index_537430 ? add_542278 : sel_542275;
  assign add_542282 = sel_542279 + 8'h01;
  assign sel_542283 = array_index_542002 == array_index_537436 ? add_542282 : sel_542279;
  assign add_542286 = sel_542283 + 8'h01;
  assign sel_542287 = array_index_542002 == array_index_537442 ? add_542286 : sel_542283;
  assign add_542290 = sel_542287 + 8'h01;
  assign sel_542291 = array_index_542002 == array_index_537448 ? add_542290 : sel_542287;
  assign add_542294 = sel_542291 + 8'h01;
  assign sel_542295 = array_index_542002 == array_index_537454 ? add_542294 : sel_542291;
  assign add_542298 = sel_542295 + 8'h01;
  assign sel_542299 = array_index_542002 == array_index_537460 ? add_542298 : sel_542295;
  assign add_542303 = sel_542299 + 8'h01;
  assign array_index_542304 = set1_unflattened[7'h11];
  assign sel_542305 = array_index_542002 == array_index_537466 ? add_542303 : sel_542299;
  assign add_542308 = sel_542305 + 8'h01;
  assign sel_542309 = array_index_542304 == array_index_537012 ? add_542308 : sel_542305;
  assign add_542312 = sel_542309 + 8'h01;
  assign sel_542313 = array_index_542304 == array_index_537016 ? add_542312 : sel_542309;
  assign add_542316 = sel_542313 + 8'h01;
  assign sel_542317 = array_index_542304 == array_index_537024 ? add_542316 : sel_542313;
  assign add_542320 = sel_542317 + 8'h01;
  assign sel_542321 = array_index_542304 == array_index_537032 ? add_542320 : sel_542317;
  assign add_542324 = sel_542321 + 8'h01;
  assign sel_542325 = array_index_542304 == array_index_537040 ? add_542324 : sel_542321;
  assign add_542328 = sel_542325 + 8'h01;
  assign sel_542329 = array_index_542304 == array_index_537048 ? add_542328 : sel_542325;
  assign add_542332 = sel_542329 + 8'h01;
  assign sel_542333 = array_index_542304 == array_index_537056 ? add_542332 : sel_542329;
  assign add_542336 = sel_542333 + 8'h01;
  assign sel_542337 = array_index_542304 == array_index_537064 ? add_542336 : sel_542333;
  assign add_542340 = sel_542337 + 8'h01;
  assign sel_542341 = array_index_542304 == array_index_537070 ? add_542340 : sel_542337;
  assign add_542344 = sel_542341 + 8'h01;
  assign sel_542345 = array_index_542304 == array_index_537076 ? add_542344 : sel_542341;
  assign add_542348 = sel_542345 + 8'h01;
  assign sel_542349 = array_index_542304 == array_index_537082 ? add_542348 : sel_542345;
  assign add_542352 = sel_542349 + 8'h01;
  assign sel_542353 = array_index_542304 == array_index_537088 ? add_542352 : sel_542349;
  assign add_542356 = sel_542353 + 8'h01;
  assign sel_542357 = array_index_542304 == array_index_537094 ? add_542356 : sel_542353;
  assign add_542360 = sel_542357 + 8'h01;
  assign sel_542361 = array_index_542304 == array_index_537100 ? add_542360 : sel_542357;
  assign add_542364 = sel_542361 + 8'h01;
  assign sel_542365 = array_index_542304 == array_index_537106 ? add_542364 : sel_542361;
  assign add_542368 = sel_542365 + 8'h01;
  assign sel_542369 = array_index_542304 == array_index_537112 ? add_542368 : sel_542365;
  assign add_542372 = sel_542369 + 8'h01;
  assign sel_542373 = array_index_542304 == array_index_537118 ? add_542372 : sel_542369;
  assign add_542376 = sel_542373 + 8'h01;
  assign sel_542377 = array_index_542304 == array_index_537124 ? add_542376 : sel_542373;
  assign add_542380 = sel_542377 + 8'h01;
  assign sel_542381 = array_index_542304 == array_index_537130 ? add_542380 : sel_542377;
  assign add_542384 = sel_542381 + 8'h01;
  assign sel_542385 = array_index_542304 == array_index_537136 ? add_542384 : sel_542381;
  assign add_542388 = sel_542385 + 8'h01;
  assign sel_542389 = array_index_542304 == array_index_537142 ? add_542388 : sel_542385;
  assign add_542392 = sel_542389 + 8'h01;
  assign sel_542393 = array_index_542304 == array_index_537148 ? add_542392 : sel_542389;
  assign add_542396 = sel_542393 + 8'h01;
  assign sel_542397 = array_index_542304 == array_index_537154 ? add_542396 : sel_542393;
  assign add_542400 = sel_542397 + 8'h01;
  assign sel_542401 = array_index_542304 == array_index_537160 ? add_542400 : sel_542397;
  assign add_542404 = sel_542401 + 8'h01;
  assign sel_542405 = array_index_542304 == array_index_537166 ? add_542404 : sel_542401;
  assign add_542408 = sel_542405 + 8'h01;
  assign sel_542409 = array_index_542304 == array_index_537172 ? add_542408 : sel_542405;
  assign add_542412 = sel_542409 + 8'h01;
  assign sel_542413 = array_index_542304 == array_index_537178 ? add_542412 : sel_542409;
  assign add_542416 = sel_542413 + 8'h01;
  assign sel_542417 = array_index_542304 == array_index_537184 ? add_542416 : sel_542413;
  assign add_542420 = sel_542417 + 8'h01;
  assign sel_542421 = array_index_542304 == array_index_537190 ? add_542420 : sel_542417;
  assign add_542424 = sel_542421 + 8'h01;
  assign sel_542425 = array_index_542304 == array_index_537196 ? add_542424 : sel_542421;
  assign add_542428 = sel_542425 + 8'h01;
  assign sel_542429 = array_index_542304 == array_index_537202 ? add_542428 : sel_542425;
  assign add_542432 = sel_542429 + 8'h01;
  assign sel_542433 = array_index_542304 == array_index_537208 ? add_542432 : sel_542429;
  assign add_542436 = sel_542433 + 8'h01;
  assign sel_542437 = array_index_542304 == array_index_537214 ? add_542436 : sel_542433;
  assign add_542440 = sel_542437 + 8'h01;
  assign sel_542441 = array_index_542304 == array_index_537220 ? add_542440 : sel_542437;
  assign add_542444 = sel_542441 + 8'h01;
  assign sel_542445 = array_index_542304 == array_index_537226 ? add_542444 : sel_542441;
  assign add_542448 = sel_542445 + 8'h01;
  assign sel_542449 = array_index_542304 == array_index_537232 ? add_542448 : sel_542445;
  assign add_542452 = sel_542449 + 8'h01;
  assign sel_542453 = array_index_542304 == array_index_537238 ? add_542452 : sel_542449;
  assign add_542456 = sel_542453 + 8'h01;
  assign sel_542457 = array_index_542304 == array_index_537244 ? add_542456 : sel_542453;
  assign add_542460 = sel_542457 + 8'h01;
  assign sel_542461 = array_index_542304 == array_index_537250 ? add_542460 : sel_542457;
  assign add_542464 = sel_542461 + 8'h01;
  assign sel_542465 = array_index_542304 == array_index_537256 ? add_542464 : sel_542461;
  assign add_542468 = sel_542465 + 8'h01;
  assign sel_542469 = array_index_542304 == array_index_537262 ? add_542468 : sel_542465;
  assign add_542472 = sel_542469 + 8'h01;
  assign sel_542473 = array_index_542304 == array_index_537268 ? add_542472 : sel_542469;
  assign add_542476 = sel_542473 + 8'h01;
  assign sel_542477 = array_index_542304 == array_index_537274 ? add_542476 : sel_542473;
  assign add_542480 = sel_542477 + 8'h01;
  assign sel_542481 = array_index_542304 == array_index_537280 ? add_542480 : sel_542477;
  assign add_542484 = sel_542481 + 8'h01;
  assign sel_542485 = array_index_542304 == array_index_537286 ? add_542484 : sel_542481;
  assign add_542488 = sel_542485 + 8'h01;
  assign sel_542489 = array_index_542304 == array_index_537292 ? add_542488 : sel_542485;
  assign add_542492 = sel_542489 + 8'h01;
  assign sel_542493 = array_index_542304 == array_index_537298 ? add_542492 : sel_542489;
  assign add_542496 = sel_542493 + 8'h01;
  assign sel_542497 = array_index_542304 == array_index_537304 ? add_542496 : sel_542493;
  assign add_542500 = sel_542497 + 8'h01;
  assign sel_542501 = array_index_542304 == array_index_537310 ? add_542500 : sel_542497;
  assign add_542504 = sel_542501 + 8'h01;
  assign sel_542505 = array_index_542304 == array_index_537316 ? add_542504 : sel_542501;
  assign add_542508 = sel_542505 + 8'h01;
  assign sel_542509 = array_index_542304 == array_index_537322 ? add_542508 : sel_542505;
  assign add_542512 = sel_542509 + 8'h01;
  assign sel_542513 = array_index_542304 == array_index_537328 ? add_542512 : sel_542509;
  assign add_542516 = sel_542513 + 8'h01;
  assign sel_542517 = array_index_542304 == array_index_537334 ? add_542516 : sel_542513;
  assign add_542520 = sel_542517 + 8'h01;
  assign sel_542521 = array_index_542304 == array_index_537340 ? add_542520 : sel_542517;
  assign add_542524 = sel_542521 + 8'h01;
  assign sel_542525 = array_index_542304 == array_index_537346 ? add_542524 : sel_542521;
  assign add_542528 = sel_542525 + 8'h01;
  assign sel_542529 = array_index_542304 == array_index_537352 ? add_542528 : sel_542525;
  assign add_542532 = sel_542529 + 8'h01;
  assign sel_542533 = array_index_542304 == array_index_537358 ? add_542532 : sel_542529;
  assign add_542536 = sel_542533 + 8'h01;
  assign sel_542537 = array_index_542304 == array_index_537364 ? add_542536 : sel_542533;
  assign add_542540 = sel_542537 + 8'h01;
  assign sel_542541 = array_index_542304 == array_index_537370 ? add_542540 : sel_542537;
  assign add_542544 = sel_542541 + 8'h01;
  assign sel_542545 = array_index_542304 == array_index_537376 ? add_542544 : sel_542541;
  assign add_542548 = sel_542545 + 8'h01;
  assign sel_542549 = array_index_542304 == array_index_537382 ? add_542548 : sel_542545;
  assign add_542552 = sel_542549 + 8'h01;
  assign sel_542553 = array_index_542304 == array_index_537388 ? add_542552 : sel_542549;
  assign add_542556 = sel_542553 + 8'h01;
  assign sel_542557 = array_index_542304 == array_index_537394 ? add_542556 : sel_542553;
  assign add_542560 = sel_542557 + 8'h01;
  assign sel_542561 = array_index_542304 == array_index_537400 ? add_542560 : sel_542557;
  assign add_542564 = sel_542561 + 8'h01;
  assign sel_542565 = array_index_542304 == array_index_537406 ? add_542564 : sel_542561;
  assign add_542568 = sel_542565 + 8'h01;
  assign sel_542569 = array_index_542304 == array_index_537412 ? add_542568 : sel_542565;
  assign add_542572 = sel_542569 + 8'h01;
  assign sel_542573 = array_index_542304 == array_index_537418 ? add_542572 : sel_542569;
  assign add_542576 = sel_542573 + 8'h01;
  assign sel_542577 = array_index_542304 == array_index_537424 ? add_542576 : sel_542573;
  assign add_542580 = sel_542577 + 8'h01;
  assign sel_542581 = array_index_542304 == array_index_537430 ? add_542580 : sel_542577;
  assign add_542584 = sel_542581 + 8'h01;
  assign sel_542585 = array_index_542304 == array_index_537436 ? add_542584 : sel_542581;
  assign add_542588 = sel_542585 + 8'h01;
  assign sel_542589 = array_index_542304 == array_index_537442 ? add_542588 : sel_542585;
  assign add_542592 = sel_542589 + 8'h01;
  assign sel_542593 = array_index_542304 == array_index_537448 ? add_542592 : sel_542589;
  assign add_542596 = sel_542593 + 8'h01;
  assign sel_542597 = array_index_542304 == array_index_537454 ? add_542596 : sel_542593;
  assign add_542600 = sel_542597 + 8'h01;
  assign sel_542601 = array_index_542304 == array_index_537460 ? add_542600 : sel_542597;
  assign add_542605 = sel_542601 + 8'h01;
  assign array_index_542606 = set1_unflattened[7'h12];
  assign sel_542607 = array_index_542304 == array_index_537466 ? add_542605 : sel_542601;
  assign add_542610 = sel_542607 + 8'h01;
  assign sel_542611 = array_index_542606 == array_index_537012 ? add_542610 : sel_542607;
  assign add_542614 = sel_542611 + 8'h01;
  assign sel_542615 = array_index_542606 == array_index_537016 ? add_542614 : sel_542611;
  assign add_542618 = sel_542615 + 8'h01;
  assign sel_542619 = array_index_542606 == array_index_537024 ? add_542618 : sel_542615;
  assign add_542622 = sel_542619 + 8'h01;
  assign sel_542623 = array_index_542606 == array_index_537032 ? add_542622 : sel_542619;
  assign add_542626 = sel_542623 + 8'h01;
  assign sel_542627 = array_index_542606 == array_index_537040 ? add_542626 : sel_542623;
  assign add_542630 = sel_542627 + 8'h01;
  assign sel_542631 = array_index_542606 == array_index_537048 ? add_542630 : sel_542627;
  assign add_542634 = sel_542631 + 8'h01;
  assign sel_542635 = array_index_542606 == array_index_537056 ? add_542634 : sel_542631;
  assign add_542638 = sel_542635 + 8'h01;
  assign sel_542639 = array_index_542606 == array_index_537064 ? add_542638 : sel_542635;
  assign add_542642 = sel_542639 + 8'h01;
  assign sel_542643 = array_index_542606 == array_index_537070 ? add_542642 : sel_542639;
  assign add_542646 = sel_542643 + 8'h01;
  assign sel_542647 = array_index_542606 == array_index_537076 ? add_542646 : sel_542643;
  assign add_542650 = sel_542647 + 8'h01;
  assign sel_542651 = array_index_542606 == array_index_537082 ? add_542650 : sel_542647;
  assign add_542654 = sel_542651 + 8'h01;
  assign sel_542655 = array_index_542606 == array_index_537088 ? add_542654 : sel_542651;
  assign add_542658 = sel_542655 + 8'h01;
  assign sel_542659 = array_index_542606 == array_index_537094 ? add_542658 : sel_542655;
  assign add_542662 = sel_542659 + 8'h01;
  assign sel_542663 = array_index_542606 == array_index_537100 ? add_542662 : sel_542659;
  assign add_542666 = sel_542663 + 8'h01;
  assign sel_542667 = array_index_542606 == array_index_537106 ? add_542666 : sel_542663;
  assign add_542670 = sel_542667 + 8'h01;
  assign sel_542671 = array_index_542606 == array_index_537112 ? add_542670 : sel_542667;
  assign add_542674 = sel_542671 + 8'h01;
  assign sel_542675 = array_index_542606 == array_index_537118 ? add_542674 : sel_542671;
  assign add_542678 = sel_542675 + 8'h01;
  assign sel_542679 = array_index_542606 == array_index_537124 ? add_542678 : sel_542675;
  assign add_542682 = sel_542679 + 8'h01;
  assign sel_542683 = array_index_542606 == array_index_537130 ? add_542682 : sel_542679;
  assign add_542686 = sel_542683 + 8'h01;
  assign sel_542687 = array_index_542606 == array_index_537136 ? add_542686 : sel_542683;
  assign add_542690 = sel_542687 + 8'h01;
  assign sel_542691 = array_index_542606 == array_index_537142 ? add_542690 : sel_542687;
  assign add_542694 = sel_542691 + 8'h01;
  assign sel_542695 = array_index_542606 == array_index_537148 ? add_542694 : sel_542691;
  assign add_542698 = sel_542695 + 8'h01;
  assign sel_542699 = array_index_542606 == array_index_537154 ? add_542698 : sel_542695;
  assign add_542702 = sel_542699 + 8'h01;
  assign sel_542703 = array_index_542606 == array_index_537160 ? add_542702 : sel_542699;
  assign add_542706 = sel_542703 + 8'h01;
  assign sel_542707 = array_index_542606 == array_index_537166 ? add_542706 : sel_542703;
  assign add_542710 = sel_542707 + 8'h01;
  assign sel_542711 = array_index_542606 == array_index_537172 ? add_542710 : sel_542707;
  assign add_542714 = sel_542711 + 8'h01;
  assign sel_542715 = array_index_542606 == array_index_537178 ? add_542714 : sel_542711;
  assign add_542718 = sel_542715 + 8'h01;
  assign sel_542719 = array_index_542606 == array_index_537184 ? add_542718 : sel_542715;
  assign add_542722 = sel_542719 + 8'h01;
  assign sel_542723 = array_index_542606 == array_index_537190 ? add_542722 : sel_542719;
  assign add_542726 = sel_542723 + 8'h01;
  assign sel_542727 = array_index_542606 == array_index_537196 ? add_542726 : sel_542723;
  assign add_542730 = sel_542727 + 8'h01;
  assign sel_542731 = array_index_542606 == array_index_537202 ? add_542730 : sel_542727;
  assign add_542734 = sel_542731 + 8'h01;
  assign sel_542735 = array_index_542606 == array_index_537208 ? add_542734 : sel_542731;
  assign add_542738 = sel_542735 + 8'h01;
  assign sel_542739 = array_index_542606 == array_index_537214 ? add_542738 : sel_542735;
  assign add_542742 = sel_542739 + 8'h01;
  assign sel_542743 = array_index_542606 == array_index_537220 ? add_542742 : sel_542739;
  assign add_542746 = sel_542743 + 8'h01;
  assign sel_542747 = array_index_542606 == array_index_537226 ? add_542746 : sel_542743;
  assign add_542750 = sel_542747 + 8'h01;
  assign sel_542751 = array_index_542606 == array_index_537232 ? add_542750 : sel_542747;
  assign add_542754 = sel_542751 + 8'h01;
  assign sel_542755 = array_index_542606 == array_index_537238 ? add_542754 : sel_542751;
  assign add_542758 = sel_542755 + 8'h01;
  assign sel_542759 = array_index_542606 == array_index_537244 ? add_542758 : sel_542755;
  assign add_542762 = sel_542759 + 8'h01;
  assign sel_542763 = array_index_542606 == array_index_537250 ? add_542762 : sel_542759;
  assign add_542766 = sel_542763 + 8'h01;
  assign sel_542767 = array_index_542606 == array_index_537256 ? add_542766 : sel_542763;
  assign add_542770 = sel_542767 + 8'h01;
  assign sel_542771 = array_index_542606 == array_index_537262 ? add_542770 : sel_542767;
  assign add_542774 = sel_542771 + 8'h01;
  assign sel_542775 = array_index_542606 == array_index_537268 ? add_542774 : sel_542771;
  assign add_542778 = sel_542775 + 8'h01;
  assign sel_542779 = array_index_542606 == array_index_537274 ? add_542778 : sel_542775;
  assign add_542782 = sel_542779 + 8'h01;
  assign sel_542783 = array_index_542606 == array_index_537280 ? add_542782 : sel_542779;
  assign add_542786 = sel_542783 + 8'h01;
  assign sel_542787 = array_index_542606 == array_index_537286 ? add_542786 : sel_542783;
  assign add_542790 = sel_542787 + 8'h01;
  assign sel_542791 = array_index_542606 == array_index_537292 ? add_542790 : sel_542787;
  assign add_542794 = sel_542791 + 8'h01;
  assign sel_542795 = array_index_542606 == array_index_537298 ? add_542794 : sel_542791;
  assign add_542798 = sel_542795 + 8'h01;
  assign sel_542799 = array_index_542606 == array_index_537304 ? add_542798 : sel_542795;
  assign add_542802 = sel_542799 + 8'h01;
  assign sel_542803 = array_index_542606 == array_index_537310 ? add_542802 : sel_542799;
  assign add_542806 = sel_542803 + 8'h01;
  assign sel_542807 = array_index_542606 == array_index_537316 ? add_542806 : sel_542803;
  assign add_542810 = sel_542807 + 8'h01;
  assign sel_542811 = array_index_542606 == array_index_537322 ? add_542810 : sel_542807;
  assign add_542814 = sel_542811 + 8'h01;
  assign sel_542815 = array_index_542606 == array_index_537328 ? add_542814 : sel_542811;
  assign add_542818 = sel_542815 + 8'h01;
  assign sel_542819 = array_index_542606 == array_index_537334 ? add_542818 : sel_542815;
  assign add_542822 = sel_542819 + 8'h01;
  assign sel_542823 = array_index_542606 == array_index_537340 ? add_542822 : sel_542819;
  assign add_542826 = sel_542823 + 8'h01;
  assign sel_542827 = array_index_542606 == array_index_537346 ? add_542826 : sel_542823;
  assign add_542830 = sel_542827 + 8'h01;
  assign sel_542831 = array_index_542606 == array_index_537352 ? add_542830 : sel_542827;
  assign add_542834 = sel_542831 + 8'h01;
  assign sel_542835 = array_index_542606 == array_index_537358 ? add_542834 : sel_542831;
  assign add_542838 = sel_542835 + 8'h01;
  assign sel_542839 = array_index_542606 == array_index_537364 ? add_542838 : sel_542835;
  assign add_542842 = sel_542839 + 8'h01;
  assign sel_542843 = array_index_542606 == array_index_537370 ? add_542842 : sel_542839;
  assign add_542846 = sel_542843 + 8'h01;
  assign sel_542847 = array_index_542606 == array_index_537376 ? add_542846 : sel_542843;
  assign add_542850 = sel_542847 + 8'h01;
  assign sel_542851 = array_index_542606 == array_index_537382 ? add_542850 : sel_542847;
  assign add_542854 = sel_542851 + 8'h01;
  assign sel_542855 = array_index_542606 == array_index_537388 ? add_542854 : sel_542851;
  assign add_542858 = sel_542855 + 8'h01;
  assign sel_542859 = array_index_542606 == array_index_537394 ? add_542858 : sel_542855;
  assign add_542862 = sel_542859 + 8'h01;
  assign sel_542863 = array_index_542606 == array_index_537400 ? add_542862 : sel_542859;
  assign add_542866 = sel_542863 + 8'h01;
  assign sel_542867 = array_index_542606 == array_index_537406 ? add_542866 : sel_542863;
  assign add_542870 = sel_542867 + 8'h01;
  assign sel_542871 = array_index_542606 == array_index_537412 ? add_542870 : sel_542867;
  assign add_542874 = sel_542871 + 8'h01;
  assign sel_542875 = array_index_542606 == array_index_537418 ? add_542874 : sel_542871;
  assign add_542878 = sel_542875 + 8'h01;
  assign sel_542879 = array_index_542606 == array_index_537424 ? add_542878 : sel_542875;
  assign add_542882 = sel_542879 + 8'h01;
  assign sel_542883 = array_index_542606 == array_index_537430 ? add_542882 : sel_542879;
  assign add_542886 = sel_542883 + 8'h01;
  assign sel_542887 = array_index_542606 == array_index_537436 ? add_542886 : sel_542883;
  assign add_542890 = sel_542887 + 8'h01;
  assign sel_542891 = array_index_542606 == array_index_537442 ? add_542890 : sel_542887;
  assign add_542894 = sel_542891 + 8'h01;
  assign sel_542895 = array_index_542606 == array_index_537448 ? add_542894 : sel_542891;
  assign add_542898 = sel_542895 + 8'h01;
  assign sel_542899 = array_index_542606 == array_index_537454 ? add_542898 : sel_542895;
  assign add_542902 = sel_542899 + 8'h01;
  assign sel_542903 = array_index_542606 == array_index_537460 ? add_542902 : sel_542899;
  assign add_542907 = sel_542903 + 8'h01;
  assign array_index_542908 = set1_unflattened[7'h13];
  assign sel_542909 = array_index_542606 == array_index_537466 ? add_542907 : sel_542903;
  assign add_542912 = sel_542909 + 8'h01;
  assign sel_542913 = array_index_542908 == array_index_537012 ? add_542912 : sel_542909;
  assign add_542916 = sel_542913 + 8'h01;
  assign sel_542917 = array_index_542908 == array_index_537016 ? add_542916 : sel_542913;
  assign add_542920 = sel_542917 + 8'h01;
  assign sel_542921 = array_index_542908 == array_index_537024 ? add_542920 : sel_542917;
  assign add_542924 = sel_542921 + 8'h01;
  assign sel_542925 = array_index_542908 == array_index_537032 ? add_542924 : sel_542921;
  assign add_542928 = sel_542925 + 8'h01;
  assign sel_542929 = array_index_542908 == array_index_537040 ? add_542928 : sel_542925;
  assign add_542932 = sel_542929 + 8'h01;
  assign sel_542933 = array_index_542908 == array_index_537048 ? add_542932 : sel_542929;
  assign add_542936 = sel_542933 + 8'h01;
  assign sel_542937 = array_index_542908 == array_index_537056 ? add_542936 : sel_542933;
  assign add_542940 = sel_542937 + 8'h01;
  assign sel_542941 = array_index_542908 == array_index_537064 ? add_542940 : sel_542937;
  assign add_542944 = sel_542941 + 8'h01;
  assign sel_542945 = array_index_542908 == array_index_537070 ? add_542944 : sel_542941;
  assign add_542948 = sel_542945 + 8'h01;
  assign sel_542949 = array_index_542908 == array_index_537076 ? add_542948 : sel_542945;
  assign add_542952 = sel_542949 + 8'h01;
  assign sel_542953 = array_index_542908 == array_index_537082 ? add_542952 : sel_542949;
  assign add_542956 = sel_542953 + 8'h01;
  assign sel_542957 = array_index_542908 == array_index_537088 ? add_542956 : sel_542953;
  assign add_542960 = sel_542957 + 8'h01;
  assign sel_542961 = array_index_542908 == array_index_537094 ? add_542960 : sel_542957;
  assign add_542964 = sel_542961 + 8'h01;
  assign sel_542965 = array_index_542908 == array_index_537100 ? add_542964 : sel_542961;
  assign add_542968 = sel_542965 + 8'h01;
  assign sel_542969 = array_index_542908 == array_index_537106 ? add_542968 : sel_542965;
  assign add_542972 = sel_542969 + 8'h01;
  assign sel_542973 = array_index_542908 == array_index_537112 ? add_542972 : sel_542969;
  assign add_542976 = sel_542973 + 8'h01;
  assign sel_542977 = array_index_542908 == array_index_537118 ? add_542976 : sel_542973;
  assign add_542980 = sel_542977 + 8'h01;
  assign sel_542981 = array_index_542908 == array_index_537124 ? add_542980 : sel_542977;
  assign add_542984 = sel_542981 + 8'h01;
  assign sel_542985 = array_index_542908 == array_index_537130 ? add_542984 : sel_542981;
  assign add_542988 = sel_542985 + 8'h01;
  assign sel_542989 = array_index_542908 == array_index_537136 ? add_542988 : sel_542985;
  assign add_542992 = sel_542989 + 8'h01;
  assign sel_542993 = array_index_542908 == array_index_537142 ? add_542992 : sel_542989;
  assign add_542996 = sel_542993 + 8'h01;
  assign sel_542997 = array_index_542908 == array_index_537148 ? add_542996 : sel_542993;
  assign add_543000 = sel_542997 + 8'h01;
  assign sel_543001 = array_index_542908 == array_index_537154 ? add_543000 : sel_542997;
  assign add_543004 = sel_543001 + 8'h01;
  assign sel_543005 = array_index_542908 == array_index_537160 ? add_543004 : sel_543001;
  assign add_543008 = sel_543005 + 8'h01;
  assign sel_543009 = array_index_542908 == array_index_537166 ? add_543008 : sel_543005;
  assign add_543012 = sel_543009 + 8'h01;
  assign sel_543013 = array_index_542908 == array_index_537172 ? add_543012 : sel_543009;
  assign add_543016 = sel_543013 + 8'h01;
  assign sel_543017 = array_index_542908 == array_index_537178 ? add_543016 : sel_543013;
  assign add_543020 = sel_543017 + 8'h01;
  assign sel_543021 = array_index_542908 == array_index_537184 ? add_543020 : sel_543017;
  assign add_543024 = sel_543021 + 8'h01;
  assign sel_543025 = array_index_542908 == array_index_537190 ? add_543024 : sel_543021;
  assign add_543028 = sel_543025 + 8'h01;
  assign sel_543029 = array_index_542908 == array_index_537196 ? add_543028 : sel_543025;
  assign add_543032 = sel_543029 + 8'h01;
  assign sel_543033 = array_index_542908 == array_index_537202 ? add_543032 : sel_543029;
  assign add_543036 = sel_543033 + 8'h01;
  assign sel_543037 = array_index_542908 == array_index_537208 ? add_543036 : sel_543033;
  assign add_543040 = sel_543037 + 8'h01;
  assign sel_543041 = array_index_542908 == array_index_537214 ? add_543040 : sel_543037;
  assign add_543044 = sel_543041 + 8'h01;
  assign sel_543045 = array_index_542908 == array_index_537220 ? add_543044 : sel_543041;
  assign add_543048 = sel_543045 + 8'h01;
  assign sel_543049 = array_index_542908 == array_index_537226 ? add_543048 : sel_543045;
  assign add_543052 = sel_543049 + 8'h01;
  assign sel_543053 = array_index_542908 == array_index_537232 ? add_543052 : sel_543049;
  assign add_543056 = sel_543053 + 8'h01;
  assign sel_543057 = array_index_542908 == array_index_537238 ? add_543056 : sel_543053;
  assign add_543060 = sel_543057 + 8'h01;
  assign sel_543061 = array_index_542908 == array_index_537244 ? add_543060 : sel_543057;
  assign add_543064 = sel_543061 + 8'h01;
  assign sel_543065 = array_index_542908 == array_index_537250 ? add_543064 : sel_543061;
  assign add_543068 = sel_543065 + 8'h01;
  assign sel_543069 = array_index_542908 == array_index_537256 ? add_543068 : sel_543065;
  assign add_543072 = sel_543069 + 8'h01;
  assign sel_543073 = array_index_542908 == array_index_537262 ? add_543072 : sel_543069;
  assign add_543076 = sel_543073 + 8'h01;
  assign sel_543077 = array_index_542908 == array_index_537268 ? add_543076 : sel_543073;
  assign add_543080 = sel_543077 + 8'h01;
  assign sel_543081 = array_index_542908 == array_index_537274 ? add_543080 : sel_543077;
  assign add_543084 = sel_543081 + 8'h01;
  assign sel_543085 = array_index_542908 == array_index_537280 ? add_543084 : sel_543081;
  assign add_543088 = sel_543085 + 8'h01;
  assign sel_543089 = array_index_542908 == array_index_537286 ? add_543088 : sel_543085;
  assign add_543092 = sel_543089 + 8'h01;
  assign sel_543093 = array_index_542908 == array_index_537292 ? add_543092 : sel_543089;
  assign add_543096 = sel_543093 + 8'h01;
  assign sel_543097 = array_index_542908 == array_index_537298 ? add_543096 : sel_543093;
  assign add_543100 = sel_543097 + 8'h01;
  assign sel_543101 = array_index_542908 == array_index_537304 ? add_543100 : sel_543097;
  assign add_543104 = sel_543101 + 8'h01;
  assign sel_543105 = array_index_542908 == array_index_537310 ? add_543104 : sel_543101;
  assign add_543108 = sel_543105 + 8'h01;
  assign sel_543109 = array_index_542908 == array_index_537316 ? add_543108 : sel_543105;
  assign add_543112 = sel_543109 + 8'h01;
  assign sel_543113 = array_index_542908 == array_index_537322 ? add_543112 : sel_543109;
  assign add_543116 = sel_543113 + 8'h01;
  assign sel_543117 = array_index_542908 == array_index_537328 ? add_543116 : sel_543113;
  assign add_543120 = sel_543117 + 8'h01;
  assign sel_543121 = array_index_542908 == array_index_537334 ? add_543120 : sel_543117;
  assign add_543124 = sel_543121 + 8'h01;
  assign sel_543125 = array_index_542908 == array_index_537340 ? add_543124 : sel_543121;
  assign add_543128 = sel_543125 + 8'h01;
  assign sel_543129 = array_index_542908 == array_index_537346 ? add_543128 : sel_543125;
  assign add_543132 = sel_543129 + 8'h01;
  assign sel_543133 = array_index_542908 == array_index_537352 ? add_543132 : sel_543129;
  assign add_543136 = sel_543133 + 8'h01;
  assign sel_543137 = array_index_542908 == array_index_537358 ? add_543136 : sel_543133;
  assign add_543140 = sel_543137 + 8'h01;
  assign sel_543141 = array_index_542908 == array_index_537364 ? add_543140 : sel_543137;
  assign add_543144 = sel_543141 + 8'h01;
  assign sel_543145 = array_index_542908 == array_index_537370 ? add_543144 : sel_543141;
  assign add_543148 = sel_543145 + 8'h01;
  assign sel_543149 = array_index_542908 == array_index_537376 ? add_543148 : sel_543145;
  assign add_543152 = sel_543149 + 8'h01;
  assign sel_543153 = array_index_542908 == array_index_537382 ? add_543152 : sel_543149;
  assign add_543156 = sel_543153 + 8'h01;
  assign sel_543157 = array_index_542908 == array_index_537388 ? add_543156 : sel_543153;
  assign add_543160 = sel_543157 + 8'h01;
  assign sel_543161 = array_index_542908 == array_index_537394 ? add_543160 : sel_543157;
  assign add_543164 = sel_543161 + 8'h01;
  assign sel_543165 = array_index_542908 == array_index_537400 ? add_543164 : sel_543161;
  assign add_543168 = sel_543165 + 8'h01;
  assign sel_543169 = array_index_542908 == array_index_537406 ? add_543168 : sel_543165;
  assign add_543172 = sel_543169 + 8'h01;
  assign sel_543173 = array_index_542908 == array_index_537412 ? add_543172 : sel_543169;
  assign add_543176 = sel_543173 + 8'h01;
  assign sel_543177 = array_index_542908 == array_index_537418 ? add_543176 : sel_543173;
  assign add_543180 = sel_543177 + 8'h01;
  assign sel_543181 = array_index_542908 == array_index_537424 ? add_543180 : sel_543177;
  assign add_543184 = sel_543181 + 8'h01;
  assign sel_543185 = array_index_542908 == array_index_537430 ? add_543184 : sel_543181;
  assign add_543188 = sel_543185 + 8'h01;
  assign sel_543189 = array_index_542908 == array_index_537436 ? add_543188 : sel_543185;
  assign add_543192 = sel_543189 + 8'h01;
  assign sel_543193 = array_index_542908 == array_index_537442 ? add_543192 : sel_543189;
  assign add_543196 = sel_543193 + 8'h01;
  assign sel_543197 = array_index_542908 == array_index_537448 ? add_543196 : sel_543193;
  assign add_543200 = sel_543197 + 8'h01;
  assign sel_543201 = array_index_542908 == array_index_537454 ? add_543200 : sel_543197;
  assign add_543204 = sel_543201 + 8'h01;
  assign sel_543205 = array_index_542908 == array_index_537460 ? add_543204 : sel_543201;
  assign add_543209 = sel_543205 + 8'h01;
  assign array_index_543210 = set1_unflattened[7'h14];
  assign sel_543211 = array_index_542908 == array_index_537466 ? add_543209 : sel_543205;
  assign add_543214 = sel_543211 + 8'h01;
  assign sel_543215 = array_index_543210 == array_index_537012 ? add_543214 : sel_543211;
  assign add_543218 = sel_543215 + 8'h01;
  assign sel_543219 = array_index_543210 == array_index_537016 ? add_543218 : sel_543215;
  assign add_543222 = sel_543219 + 8'h01;
  assign sel_543223 = array_index_543210 == array_index_537024 ? add_543222 : sel_543219;
  assign add_543226 = sel_543223 + 8'h01;
  assign sel_543227 = array_index_543210 == array_index_537032 ? add_543226 : sel_543223;
  assign add_543230 = sel_543227 + 8'h01;
  assign sel_543231 = array_index_543210 == array_index_537040 ? add_543230 : sel_543227;
  assign add_543234 = sel_543231 + 8'h01;
  assign sel_543235 = array_index_543210 == array_index_537048 ? add_543234 : sel_543231;
  assign add_543238 = sel_543235 + 8'h01;
  assign sel_543239 = array_index_543210 == array_index_537056 ? add_543238 : sel_543235;
  assign add_543242 = sel_543239 + 8'h01;
  assign sel_543243 = array_index_543210 == array_index_537064 ? add_543242 : sel_543239;
  assign add_543246 = sel_543243 + 8'h01;
  assign sel_543247 = array_index_543210 == array_index_537070 ? add_543246 : sel_543243;
  assign add_543250 = sel_543247 + 8'h01;
  assign sel_543251 = array_index_543210 == array_index_537076 ? add_543250 : sel_543247;
  assign add_543254 = sel_543251 + 8'h01;
  assign sel_543255 = array_index_543210 == array_index_537082 ? add_543254 : sel_543251;
  assign add_543258 = sel_543255 + 8'h01;
  assign sel_543259 = array_index_543210 == array_index_537088 ? add_543258 : sel_543255;
  assign add_543262 = sel_543259 + 8'h01;
  assign sel_543263 = array_index_543210 == array_index_537094 ? add_543262 : sel_543259;
  assign add_543266 = sel_543263 + 8'h01;
  assign sel_543267 = array_index_543210 == array_index_537100 ? add_543266 : sel_543263;
  assign add_543270 = sel_543267 + 8'h01;
  assign sel_543271 = array_index_543210 == array_index_537106 ? add_543270 : sel_543267;
  assign add_543274 = sel_543271 + 8'h01;
  assign sel_543275 = array_index_543210 == array_index_537112 ? add_543274 : sel_543271;
  assign add_543278 = sel_543275 + 8'h01;
  assign sel_543279 = array_index_543210 == array_index_537118 ? add_543278 : sel_543275;
  assign add_543282 = sel_543279 + 8'h01;
  assign sel_543283 = array_index_543210 == array_index_537124 ? add_543282 : sel_543279;
  assign add_543286 = sel_543283 + 8'h01;
  assign sel_543287 = array_index_543210 == array_index_537130 ? add_543286 : sel_543283;
  assign add_543290 = sel_543287 + 8'h01;
  assign sel_543291 = array_index_543210 == array_index_537136 ? add_543290 : sel_543287;
  assign add_543294 = sel_543291 + 8'h01;
  assign sel_543295 = array_index_543210 == array_index_537142 ? add_543294 : sel_543291;
  assign add_543298 = sel_543295 + 8'h01;
  assign sel_543299 = array_index_543210 == array_index_537148 ? add_543298 : sel_543295;
  assign add_543302 = sel_543299 + 8'h01;
  assign sel_543303 = array_index_543210 == array_index_537154 ? add_543302 : sel_543299;
  assign add_543306 = sel_543303 + 8'h01;
  assign sel_543307 = array_index_543210 == array_index_537160 ? add_543306 : sel_543303;
  assign add_543310 = sel_543307 + 8'h01;
  assign sel_543311 = array_index_543210 == array_index_537166 ? add_543310 : sel_543307;
  assign add_543314 = sel_543311 + 8'h01;
  assign sel_543315 = array_index_543210 == array_index_537172 ? add_543314 : sel_543311;
  assign add_543318 = sel_543315 + 8'h01;
  assign sel_543319 = array_index_543210 == array_index_537178 ? add_543318 : sel_543315;
  assign add_543322 = sel_543319 + 8'h01;
  assign sel_543323 = array_index_543210 == array_index_537184 ? add_543322 : sel_543319;
  assign add_543326 = sel_543323 + 8'h01;
  assign sel_543327 = array_index_543210 == array_index_537190 ? add_543326 : sel_543323;
  assign add_543330 = sel_543327 + 8'h01;
  assign sel_543331 = array_index_543210 == array_index_537196 ? add_543330 : sel_543327;
  assign add_543334 = sel_543331 + 8'h01;
  assign sel_543335 = array_index_543210 == array_index_537202 ? add_543334 : sel_543331;
  assign add_543338 = sel_543335 + 8'h01;
  assign sel_543339 = array_index_543210 == array_index_537208 ? add_543338 : sel_543335;
  assign add_543342 = sel_543339 + 8'h01;
  assign sel_543343 = array_index_543210 == array_index_537214 ? add_543342 : sel_543339;
  assign add_543346 = sel_543343 + 8'h01;
  assign sel_543347 = array_index_543210 == array_index_537220 ? add_543346 : sel_543343;
  assign add_543350 = sel_543347 + 8'h01;
  assign sel_543351 = array_index_543210 == array_index_537226 ? add_543350 : sel_543347;
  assign add_543354 = sel_543351 + 8'h01;
  assign sel_543355 = array_index_543210 == array_index_537232 ? add_543354 : sel_543351;
  assign add_543358 = sel_543355 + 8'h01;
  assign sel_543359 = array_index_543210 == array_index_537238 ? add_543358 : sel_543355;
  assign add_543362 = sel_543359 + 8'h01;
  assign sel_543363 = array_index_543210 == array_index_537244 ? add_543362 : sel_543359;
  assign add_543366 = sel_543363 + 8'h01;
  assign sel_543367 = array_index_543210 == array_index_537250 ? add_543366 : sel_543363;
  assign add_543370 = sel_543367 + 8'h01;
  assign sel_543371 = array_index_543210 == array_index_537256 ? add_543370 : sel_543367;
  assign add_543374 = sel_543371 + 8'h01;
  assign sel_543375 = array_index_543210 == array_index_537262 ? add_543374 : sel_543371;
  assign add_543378 = sel_543375 + 8'h01;
  assign sel_543379 = array_index_543210 == array_index_537268 ? add_543378 : sel_543375;
  assign add_543382 = sel_543379 + 8'h01;
  assign sel_543383 = array_index_543210 == array_index_537274 ? add_543382 : sel_543379;
  assign add_543386 = sel_543383 + 8'h01;
  assign sel_543387 = array_index_543210 == array_index_537280 ? add_543386 : sel_543383;
  assign add_543390 = sel_543387 + 8'h01;
  assign sel_543391 = array_index_543210 == array_index_537286 ? add_543390 : sel_543387;
  assign add_543394 = sel_543391 + 8'h01;
  assign sel_543395 = array_index_543210 == array_index_537292 ? add_543394 : sel_543391;
  assign add_543398 = sel_543395 + 8'h01;
  assign sel_543399 = array_index_543210 == array_index_537298 ? add_543398 : sel_543395;
  assign add_543402 = sel_543399 + 8'h01;
  assign sel_543403 = array_index_543210 == array_index_537304 ? add_543402 : sel_543399;
  assign add_543406 = sel_543403 + 8'h01;
  assign sel_543407 = array_index_543210 == array_index_537310 ? add_543406 : sel_543403;
  assign add_543410 = sel_543407 + 8'h01;
  assign sel_543411 = array_index_543210 == array_index_537316 ? add_543410 : sel_543407;
  assign add_543414 = sel_543411 + 8'h01;
  assign sel_543415 = array_index_543210 == array_index_537322 ? add_543414 : sel_543411;
  assign add_543418 = sel_543415 + 8'h01;
  assign sel_543419 = array_index_543210 == array_index_537328 ? add_543418 : sel_543415;
  assign add_543422 = sel_543419 + 8'h01;
  assign sel_543423 = array_index_543210 == array_index_537334 ? add_543422 : sel_543419;
  assign add_543426 = sel_543423 + 8'h01;
  assign sel_543427 = array_index_543210 == array_index_537340 ? add_543426 : sel_543423;
  assign add_543430 = sel_543427 + 8'h01;
  assign sel_543431 = array_index_543210 == array_index_537346 ? add_543430 : sel_543427;
  assign add_543434 = sel_543431 + 8'h01;
  assign sel_543435 = array_index_543210 == array_index_537352 ? add_543434 : sel_543431;
  assign add_543438 = sel_543435 + 8'h01;
  assign sel_543439 = array_index_543210 == array_index_537358 ? add_543438 : sel_543435;
  assign add_543442 = sel_543439 + 8'h01;
  assign sel_543443 = array_index_543210 == array_index_537364 ? add_543442 : sel_543439;
  assign add_543446 = sel_543443 + 8'h01;
  assign sel_543447 = array_index_543210 == array_index_537370 ? add_543446 : sel_543443;
  assign add_543450 = sel_543447 + 8'h01;
  assign sel_543451 = array_index_543210 == array_index_537376 ? add_543450 : sel_543447;
  assign add_543454 = sel_543451 + 8'h01;
  assign sel_543455 = array_index_543210 == array_index_537382 ? add_543454 : sel_543451;
  assign add_543458 = sel_543455 + 8'h01;
  assign sel_543459 = array_index_543210 == array_index_537388 ? add_543458 : sel_543455;
  assign add_543462 = sel_543459 + 8'h01;
  assign sel_543463 = array_index_543210 == array_index_537394 ? add_543462 : sel_543459;
  assign add_543466 = sel_543463 + 8'h01;
  assign sel_543467 = array_index_543210 == array_index_537400 ? add_543466 : sel_543463;
  assign add_543470 = sel_543467 + 8'h01;
  assign sel_543471 = array_index_543210 == array_index_537406 ? add_543470 : sel_543467;
  assign add_543474 = sel_543471 + 8'h01;
  assign sel_543475 = array_index_543210 == array_index_537412 ? add_543474 : sel_543471;
  assign add_543478 = sel_543475 + 8'h01;
  assign sel_543479 = array_index_543210 == array_index_537418 ? add_543478 : sel_543475;
  assign add_543482 = sel_543479 + 8'h01;
  assign sel_543483 = array_index_543210 == array_index_537424 ? add_543482 : sel_543479;
  assign add_543486 = sel_543483 + 8'h01;
  assign sel_543487 = array_index_543210 == array_index_537430 ? add_543486 : sel_543483;
  assign add_543490 = sel_543487 + 8'h01;
  assign sel_543491 = array_index_543210 == array_index_537436 ? add_543490 : sel_543487;
  assign add_543494 = sel_543491 + 8'h01;
  assign sel_543495 = array_index_543210 == array_index_537442 ? add_543494 : sel_543491;
  assign add_543498 = sel_543495 + 8'h01;
  assign sel_543499 = array_index_543210 == array_index_537448 ? add_543498 : sel_543495;
  assign add_543502 = sel_543499 + 8'h01;
  assign sel_543503 = array_index_543210 == array_index_537454 ? add_543502 : sel_543499;
  assign add_543506 = sel_543503 + 8'h01;
  assign sel_543507 = array_index_543210 == array_index_537460 ? add_543506 : sel_543503;
  assign add_543511 = sel_543507 + 8'h01;
  assign array_index_543512 = set1_unflattened[7'h15];
  assign sel_543513 = array_index_543210 == array_index_537466 ? add_543511 : sel_543507;
  assign add_543516 = sel_543513 + 8'h01;
  assign sel_543517 = array_index_543512 == array_index_537012 ? add_543516 : sel_543513;
  assign add_543520 = sel_543517 + 8'h01;
  assign sel_543521 = array_index_543512 == array_index_537016 ? add_543520 : sel_543517;
  assign add_543524 = sel_543521 + 8'h01;
  assign sel_543525 = array_index_543512 == array_index_537024 ? add_543524 : sel_543521;
  assign add_543528 = sel_543525 + 8'h01;
  assign sel_543529 = array_index_543512 == array_index_537032 ? add_543528 : sel_543525;
  assign add_543532 = sel_543529 + 8'h01;
  assign sel_543533 = array_index_543512 == array_index_537040 ? add_543532 : sel_543529;
  assign add_543536 = sel_543533 + 8'h01;
  assign sel_543537 = array_index_543512 == array_index_537048 ? add_543536 : sel_543533;
  assign add_543540 = sel_543537 + 8'h01;
  assign sel_543541 = array_index_543512 == array_index_537056 ? add_543540 : sel_543537;
  assign add_543544 = sel_543541 + 8'h01;
  assign sel_543545 = array_index_543512 == array_index_537064 ? add_543544 : sel_543541;
  assign add_543548 = sel_543545 + 8'h01;
  assign sel_543549 = array_index_543512 == array_index_537070 ? add_543548 : sel_543545;
  assign add_543552 = sel_543549 + 8'h01;
  assign sel_543553 = array_index_543512 == array_index_537076 ? add_543552 : sel_543549;
  assign add_543556 = sel_543553 + 8'h01;
  assign sel_543557 = array_index_543512 == array_index_537082 ? add_543556 : sel_543553;
  assign add_543560 = sel_543557 + 8'h01;
  assign sel_543561 = array_index_543512 == array_index_537088 ? add_543560 : sel_543557;
  assign add_543564 = sel_543561 + 8'h01;
  assign sel_543565 = array_index_543512 == array_index_537094 ? add_543564 : sel_543561;
  assign add_543568 = sel_543565 + 8'h01;
  assign sel_543569 = array_index_543512 == array_index_537100 ? add_543568 : sel_543565;
  assign add_543572 = sel_543569 + 8'h01;
  assign sel_543573 = array_index_543512 == array_index_537106 ? add_543572 : sel_543569;
  assign add_543576 = sel_543573 + 8'h01;
  assign sel_543577 = array_index_543512 == array_index_537112 ? add_543576 : sel_543573;
  assign add_543580 = sel_543577 + 8'h01;
  assign sel_543581 = array_index_543512 == array_index_537118 ? add_543580 : sel_543577;
  assign add_543584 = sel_543581 + 8'h01;
  assign sel_543585 = array_index_543512 == array_index_537124 ? add_543584 : sel_543581;
  assign add_543588 = sel_543585 + 8'h01;
  assign sel_543589 = array_index_543512 == array_index_537130 ? add_543588 : sel_543585;
  assign add_543592 = sel_543589 + 8'h01;
  assign sel_543593 = array_index_543512 == array_index_537136 ? add_543592 : sel_543589;
  assign add_543596 = sel_543593 + 8'h01;
  assign sel_543597 = array_index_543512 == array_index_537142 ? add_543596 : sel_543593;
  assign add_543600 = sel_543597 + 8'h01;
  assign sel_543601 = array_index_543512 == array_index_537148 ? add_543600 : sel_543597;
  assign add_543604 = sel_543601 + 8'h01;
  assign sel_543605 = array_index_543512 == array_index_537154 ? add_543604 : sel_543601;
  assign add_543608 = sel_543605 + 8'h01;
  assign sel_543609 = array_index_543512 == array_index_537160 ? add_543608 : sel_543605;
  assign add_543612 = sel_543609 + 8'h01;
  assign sel_543613 = array_index_543512 == array_index_537166 ? add_543612 : sel_543609;
  assign add_543616 = sel_543613 + 8'h01;
  assign sel_543617 = array_index_543512 == array_index_537172 ? add_543616 : sel_543613;
  assign add_543620 = sel_543617 + 8'h01;
  assign sel_543621 = array_index_543512 == array_index_537178 ? add_543620 : sel_543617;
  assign add_543624 = sel_543621 + 8'h01;
  assign sel_543625 = array_index_543512 == array_index_537184 ? add_543624 : sel_543621;
  assign add_543628 = sel_543625 + 8'h01;
  assign sel_543629 = array_index_543512 == array_index_537190 ? add_543628 : sel_543625;
  assign add_543632 = sel_543629 + 8'h01;
  assign sel_543633 = array_index_543512 == array_index_537196 ? add_543632 : sel_543629;
  assign add_543636 = sel_543633 + 8'h01;
  assign sel_543637 = array_index_543512 == array_index_537202 ? add_543636 : sel_543633;
  assign add_543640 = sel_543637 + 8'h01;
  assign sel_543641 = array_index_543512 == array_index_537208 ? add_543640 : sel_543637;
  assign add_543644 = sel_543641 + 8'h01;
  assign sel_543645 = array_index_543512 == array_index_537214 ? add_543644 : sel_543641;
  assign add_543648 = sel_543645 + 8'h01;
  assign sel_543649 = array_index_543512 == array_index_537220 ? add_543648 : sel_543645;
  assign add_543652 = sel_543649 + 8'h01;
  assign sel_543653 = array_index_543512 == array_index_537226 ? add_543652 : sel_543649;
  assign add_543656 = sel_543653 + 8'h01;
  assign sel_543657 = array_index_543512 == array_index_537232 ? add_543656 : sel_543653;
  assign add_543660 = sel_543657 + 8'h01;
  assign sel_543661 = array_index_543512 == array_index_537238 ? add_543660 : sel_543657;
  assign add_543664 = sel_543661 + 8'h01;
  assign sel_543665 = array_index_543512 == array_index_537244 ? add_543664 : sel_543661;
  assign add_543668 = sel_543665 + 8'h01;
  assign sel_543669 = array_index_543512 == array_index_537250 ? add_543668 : sel_543665;
  assign add_543672 = sel_543669 + 8'h01;
  assign sel_543673 = array_index_543512 == array_index_537256 ? add_543672 : sel_543669;
  assign add_543676 = sel_543673 + 8'h01;
  assign sel_543677 = array_index_543512 == array_index_537262 ? add_543676 : sel_543673;
  assign add_543680 = sel_543677 + 8'h01;
  assign sel_543681 = array_index_543512 == array_index_537268 ? add_543680 : sel_543677;
  assign add_543684 = sel_543681 + 8'h01;
  assign sel_543685 = array_index_543512 == array_index_537274 ? add_543684 : sel_543681;
  assign add_543688 = sel_543685 + 8'h01;
  assign sel_543689 = array_index_543512 == array_index_537280 ? add_543688 : sel_543685;
  assign add_543692 = sel_543689 + 8'h01;
  assign sel_543693 = array_index_543512 == array_index_537286 ? add_543692 : sel_543689;
  assign add_543696 = sel_543693 + 8'h01;
  assign sel_543697 = array_index_543512 == array_index_537292 ? add_543696 : sel_543693;
  assign add_543700 = sel_543697 + 8'h01;
  assign sel_543701 = array_index_543512 == array_index_537298 ? add_543700 : sel_543697;
  assign add_543704 = sel_543701 + 8'h01;
  assign sel_543705 = array_index_543512 == array_index_537304 ? add_543704 : sel_543701;
  assign add_543708 = sel_543705 + 8'h01;
  assign sel_543709 = array_index_543512 == array_index_537310 ? add_543708 : sel_543705;
  assign add_543712 = sel_543709 + 8'h01;
  assign sel_543713 = array_index_543512 == array_index_537316 ? add_543712 : sel_543709;
  assign add_543716 = sel_543713 + 8'h01;
  assign sel_543717 = array_index_543512 == array_index_537322 ? add_543716 : sel_543713;
  assign add_543720 = sel_543717 + 8'h01;
  assign sel_543721 = array_index_543512 == array_index_537328 ? add_543720 : sel_543717;
  assign add_543724 = sel_543721 + 8'h01;
  assign sel_543725 = array_index_543512 == array_index_537334 ? add_543724 : sel_543721;
  assign add_543728 = sel_543725 + 8'h01;
  assign sel_543729 = array_index_543512 == array_index_537340 ? add_543728 : sel_543725;
  assign add_543732 = sel_543729 + 8'h01;
  assign sel_543733 = array_index_543512 == array_index_537346 ? add_543732 : sel_543729;
  assign add_543736 = sel_543733 + 8'h01;
  assign sel_543737 = array_index_543512 == array_index_537352 ? add_543736 : sel_543733;
  assign add_543740 = sel_543737 + 8'h01;
  assign sel_543741 = array_index_543512 == array_index_537358 ? add_543740 : sel_543737;
  assign add_543744 = sel_543741 + 8'h01;
  assign sel_543745 = array_index_543512 == array_index_537364 ? add_543744 : sel_543741;
  assign add_543748 = sel_543745 + 8'h01;
  assign sel_543749 = array_index_543512 == array_index_537370 ? add_543748 : sel_543745;
  assign add_543752 = sel_543749 + 8'h01;
  assign sel_543753 = array_index_543512 == array_index_537376 ? add_543752 : sel_543749;
  assign add_543756 = sel_543753 + 8'h01;
  assign sel_543757 = array_index_543512 == array_index_537382 ? add_543756 : sel_543753;
  assign add_543760 = sel_543757 + 8'h01;
  assign sel_543761 = array_index_543512 == array_index_537388 ? add_543760 : sel_543757;
  assign add_543764 = sel_543761 + 8'h01;
  assign sel_543765 = array_index_543512 == array_index_537394 ? add_543764 : sel_543761;
  assign add_543768 = sel_543765 + 8'h01;
  assign sel_543769 = array_index_543512 == array_index_537400 ? add_543768 : sel_543765;
  assign add_543772 = sel_543769 + 8'h01;
  assign sel_543773 = array_index_543512 == array_index_537406 ? add_543772 : sel_543769;
  assign add_543776 = sel_543773 + 8'h01;
  assign sel_543777 = array_index_543512 == array_index_537412 ? add_543776 : sel_543773;
  assign add_543780 = sel_543777 + 8'h01;
  assign sel_543781 = array_index_543512 == array_index_537418 ? add_543780 : sel_543777;
  assign add_543784 = sel_543781 + 8'h01;
  assign sel_543785 = array_index_543512 == array_index_537424 ? add_543784 : sel_543781;
  assign add_543788 = sel_543785 + 8'h01;
  assign sel_543789 = array_index_543512 == array_index_537430 ? add_543788 : sel_543785;
  assign add_543792 = sel_543789 + 8'h01;
  assign sel_543793 = array_index_543512 == array_index_537436 ? add_543792 : sel_543789;
  assign add_543796 = sel_543793 + 8'h01;
  assign sel_543797 = array_index_543512 == array_index_537442 ? add_543796 : sel_543793;
  assign add_543800 = sel_543797 + 8'h01;
  assign sel_543801 = array_index_543512 == array_index_537448 ? add_543800 : sel_543797;
  assign add_543804 = sel_543801 + 8'h01;
  assign sel_543805 = array_index_543512 == array_index_537454 ? add_543804 : sel_543801;
  assign add_543808 = sel_543805 + 8'h01;
  assign sel_543809 = array_index_543512 == array_index_537460 ? add_543808 : sel_543805;
  assign add_543813 = sel_543809 + 8'h01;
  assign array_index_543814 = set1_unflattened[7'h16];
  assign sel_543815 = array_index_543512 == array_index_537466 ? add_543813 : sel_543809;
  assign add_543818 = sel_543815 + 8'h01;
  assign sel_543819 = array_index_543814 == array_index_537012 ? add_543818 : sel_543815;
  assign add_543822 = sel_543819 + 8'h01;
  assign sel_543823 = array_index_543814 == array_index_537016 ? add_543822 : sel_543819;
  assign add_543826 = sel_543823 + 8'h01;
  assign sel_543827 = array_index_543814 == array_index_537024 ? add_543826 : sel_543823;
  assign add_543830 = sel_543827 + 8'h01;
  assign sel_543831 = array_index_543814 == array_index_537032 ? add_543830 : sel_543827;
  assign add_543834 = sel_543831 + 8'h01;
  assign sel_543835 = array_index_543814 == array_index_537040 ? add_543834 : sel_543831;
  assign add_543838 = sel_543835 + 8'h01;
  assign sel_543839 = array_index_543814 == array_index_537048 ? add_543838 : sel_543835;
  assign add_543842 = sel_543839 + 8'h01;
  assign sel_543843 = array_index_543814 == array_index_537056 ? add_543842 : sel_543839;
  assign add_543846 = sel_543843 + 8'h01;
  assign sel_543847 = array_index_543814 == array_index_537064 ? add_543846 : sel_543843;
  assign add_543850 = sel_543847 + 8'h01;
  assign sel_543851 = array_index_543814 == array_index_537070 ? add_543850 : sel_543847;
  assign add_543854 = sel_543851 + 8'h01;
  assign sel_543855 = array_index_543814 == array_index_537076 ? add_543854 : sel_543851;
  assign add_543858 = sel_543855 + 8'h01;
  assign sel_543859 = array_index_543814 == array_index_537082 ? add_543858 : sel_543855;
  assign add_543862 = sel_543859 + 8'h01;
  assign sel_543863 = array_index_543814 == array_index_537088 ? add_543862 : sel_543859;
  assign add_543866 = sel_543863 + 8'h01;
  assign sel_543867 = array_index_543814 == array_index_537094 ? add_543866 : sel_543863;
  assign add_543870 = sel_543867 + 8'h01;
  assign sel_543871 = array_index_543814 == array_index_537100 ? add_543870 : sel_543867;
  assign add_543874 = sel_543871 + 8'h01;
  assign sel_543875 = array_index_543814 == array_index_537106 ? add_543874 : sel_543871;
  assign add_543878 = sel_543875 + 8'h01;
  assign sel_543879 = array_index_543814 == array_index_537112 ? add_543878 : sel_543875;
  assign add_543882 = sel_543879 + 8'h01;
  assign sel_543883 = array_index_543814 == array_index_537118 ? add_543882 : sel_543879;
  assign add_543886 = sel_543883 + 8'h01;
  assign sel_543887 = array_index_543814 == array_index_537124 ? add_543886 : sel_543883;
  assign add_543890 = sel_543887 + 8'h01;
  assign sel_543891 = array_index_543814 == array_index_537130 ? add_543890 : sel_543887;
  assign add_543894 = sel_543891 + 8'h01;
  assign sel_543895 = array_index_543814 == array_index_537136 ? add_543894 : sel_543891;
  assign add_543898 = sel_543895 + 8'h01;
  assign sel_543899 = array_index_543814 == array_index_537142 ? add_543898 : sel_543895;
  assign add_543902 = sel_543899 + 8'h01;
  assign sel_543903 = array_index_543814 == array_index_537148 ? add_543902 : sel_543899;
  assign add_543906 = sel_543903 + 8'h01;
  assign sel_543907 = array_index_543814 == array_index_537154 ? add_543906 : sel_543903;
  assign add_543910 = sel_543907 + 8'h01;
  assign sel_543911 = array_index_543814 == array_index_537160 ? add_543910 : sel_543907;
  assign add_543914 = sel_543911 + 8'h01;
  assign sel_543915 = array_index_543814 == array_index_537166 ? add_543914 : sel_543911;
  assign add_543918 = sel_543915 + 8'h01;
  assign sel_543919 = array_index_543814 == array_index_537172 ? add_543918 : sel_543915;
  assign add_543922 = sel_543919 + 8'h01;
  assign sel_543923 = array_index_543814 == array_index_537178 ? add_543922 : sel_543919;
  assign add_543926 = sel_543923 + 8'h01;
  assign sel_543927 = array_index_543814 == array_index_537184 ? add_543926 : sel_543923;
  assign add_543930 = sel_543927 + 8'h01;
  assign sel_543931 = array_index_543814 == array_index_537190 ? add_543930 : sel_543927;
  assign add_543934 = sel_543931 + 8'h01;
  assign sel_543935 = array_index_543814 == array_index_537196 ? add_543934 : sel_543931;
  assign add_543938 = sel_543935 + 8'h01;
  assign sel_543939 = array_index_543814 == array_index_537202 ? add_543938 : sel_543935;
  assign add_543942 = sel_543939 + 8'h01;
  assign sel_543943 = array_index_543814 == array_index_537208 ? add_543942 : sel_543939;
  assign add_543946 = sel_543943 + 8'h01;
  assign sel_543947 = array_index_543814 == array_index_537214 ? add_543946 : sel_543943;
  assign add_543950 = sel_543947 + 8'h01;
  assign sel_543951 = array_index_543814 == array_index_537220 ? add_543950 : sel_543947;
  assign add_543954 = sel_543951 + 8'h01;
  assign sel_543955 = array_index_543814 == array_index_537226 ? add_543954 : sel_543951;
  assign add_543958 = sel_543955 + 8'h01;
  assign sel_543959 = array_index_543814 == array_index_537232 ? add_543958 : sel_543955;
  assign add_543962 = sel_543959 + 8'h01;
  assign sel_543963 = array_index_543814 == array_index_537238 ? add_543962 : sel_543959;
  assign add_543966 = sel_543963 + 8'h01;
  assign sel_543967 = array_index_543814 == array_index_537244 ? add_543966 : sel_543963;
  assign add_543970 = sel_543967 + 8'h01;
  assign sel_543971 = array_index_543814 == array_index_537250 ? add_543970 : sel_543967;
  assign add_543974 = sel_543971 + 8'h01;
  assign sel_543975 = array_index_543814 == array_index_537256 ? add_543974 : sel_543971;
  assign add_543978 = sel_543975 + 8'h01;
  assign sel_543979 = array_index_543814 == array_index_537262 ? add_543978 : sel_543975;
  assign add_543982 = sel_543979 + 8'h01;
  assign sel_543983 = array_index_543814 == array_index_537268 ? add_543982 : sel_543979;
  assign add_543986 = sel_543983 + 8'h01;
  assign sel_543987 = array_index_543814 == array_index_537274 ? add_543986 : sel_543983;
  assign add_543990 = sel_543987 + 8'h01;
  assign sel_543991 = array_index_543814 == array_index_537280 ? add_543990 : sel_543987;
  assign add_543994 = sel_543991 + 8'h01;
  assign sel_543995 = array_index_543814 == array_index_537286 ? add_543994 : sel_543991;
  assign add_543998 = sel_543995 + 8'h01;
  assign sel_543999 = array_index_543814 == array_index_537292 ? add_543998 : sel_543995;
  assign add_544002 = sel_543999 + 8'h01;
  assign sel_544003 = array_index_543814 == array_index_537298 ? add_544002 : sel_543999;
  assign add_544006 = sel_544003 + 8'h01;
  assign sel_544007 = array_index_543814 == array_index_537304 ? add_544006 : sel_544003;
  assign add_544010 = sel_544007 + 8'h01;
  assign sel_544011 = array_index_543814 == array_index_537310 ? add_544010 : sel_544007;
  assign add_544014 = sel_544011 + 8'h01;
  assign sel_544015 = array_index_543814 == array_index_537316 ? add_544014 : sel_544011;
  assign add_544018 = sel_544015 + 8'h01;
  assign sel_544019 = array_index_543814 == array_index_537322 ? add_544018 : sel_544015;
  assign add_544022 = sel_544019 + 8'h01;
  assign sel_544023 = array_index_543814 == array_index_537328 ? add_544022 : sel_544019;
  assign add_544026 = sel_544023 + 8'h01;
  assign sel_544027 = array_index_543814 == array_index_537334 ? add_544026 : sel_544023;
  assign add_544030 = sel_544027 + 8'h01;
  assign sel_544031 = array_index_543814 == array_index_537340 ? add_544030 : sel_544027;
  assign add_544034 = sel_544031 + 8'h01;
  assign sel_544035 = array_index_543814 == array_index_537346 ? add_544034 : sel_544031;
  assign add_544038 = sel_544035 + 8'h01;
  assign sel_544039 = array_index_543814 == array_index_537352 ? add_544038 : sel_544035;
  assign add_544042 = sel_544039 + 8'h01;
  assign sel_544043 = array_index_543814 == array_index_537358 ? add_544042 : sel_544039;
  assign add_544046 = sel_544043 + 8'h01;
  assign sel_544047 = array_index_543814 == array_index_537364 ? add_544046 : sel_544043;
  assign add_544050 = sel_544047 + 8'h01;
  assign sel_544051 = array_index_543814 == array_index_537370 ? add_544050 : sel_544047;
  assign add_544054 = sel_544051 + 8'h01;
  assign sel_544055 = array_index_543814 == array_index_537376 ? add_544054 : sel_544051;
  assign add_544058 = sel_544055 + 8'h01;
  assign sel_544059 = array_index_543814 == array_index_537382 ? add_544058 : sel_544055;
  assign add_544062 = sel_544059 + 8'h01;
  assign sel_544063 = array_index_543814 == array_index_537388 ? add_544062 : sel_544059;
  assign add_544066 = sel_544063 + 8'h01;
  assign sel_544067 = array_index_543814 == array_index_537394 ? add_544066 : sel_544063;
  assign add_544070 = sel_544067 + 8'h01;
  assign sel_544071 = array_index_543814 == array_index_537400 ? add_544070 : sel_544067;
  assign add_544074 = sel_544071 + 8'h01;
  assign sel_544075 = array_index_543814 == array_index_537406 ? add_544074 : sel_544071;
  assign add_544078 = sel_544075 + 8'h01;
  assign sel_544079 = array_index_543814 == array_index_537412 ? add_544078 : sel_544075;
  assign add_544082 = sel_544079 + 8'h01;
  assign sel_544083 = array_index_543814 == array_index_537418 ? add_544082 : sel_544079;
  assign add_544086 = sel_544083 + 8'h01;
  assign sel_544087 = array_index_543814 == array_index_537424 ? add_544086 : sel_544083;
  assign add_544090 = sel_544087 + 8'h01;
  assign sel_544091 = array_index_543814 == array_index_537430 ? add_544090 : sel_544087;
  assign add_544094 = sel_544091 + 8'h01;
  assign sel_544095 = array_index_543814 == array_index_537436 ? add_544094 : sel_544091;
  assign add_544098 = sel_544095 + 8'h01;
  assign sel_544099 = array_index_543814 == array_index_537442 ? add_544098 : sel_544095;
  assign add_544102 = sel_544099 + 8'h01;
  assign sel_544103 = array_index_543814 == array_index_537448 ? add_544102 : sel_544099;
  assign add_544106 = sel_544103 + 8'h01;
  assign sel_544107 = array_index_543814 == array_index_537454 ? add_544106 : sel_544103;
  assign add_544110 = sel_544107 + 8'h01;
  assign sel_544111 = array_index_543814 == array_index_537460 ? add_544110 : sel_544107;
  assign add_544115 = sel_544111 + 8'h01;
  assign array_index_544116 = set1_unflattened[7'h17];
  assign sel_544117 = array_index_543814 == array_index_537466 ? add_544115 : sel_544111;
  assign add_544120 = sel_544117 + 8'h01;
  assign sel_544121 = array_index_544116 == array_index_537012 ? add_544120 : sel_544117;
  assign add_544124 = sel_544121 + 8'h01;
  assign sel_544125 = array_index_544116 == array_index_537016 ? add_544124 : sel_544121;
  assign add_544128 = sel_544125 + 8'h01;
  assign sel_544129 = array_index_544116 == array_index_537024 ? add_544128 : sel_544125;
  assign add_544132 = sel_544129 + 8'h01;
  assign sel_544133 = array_index_544116 == array_index_537032 ? add_544132 : sel_544129;
  assign add_544136 = sel_544133 + 8'h01;
  assign sel_544137 = array_index_544116 == array_index_537040 ? add_544136 : sel_544133;
  assign add_544140 = sel_544137 + 8'h01;
  assign sel_544141 = array_index_544116 == array_index_537048 ? add_544140 : sel_544137;
  assign add_544144 = sel_544141 + 8'h01;
  assign sel_544145 = array_index_544116 == array_index_537056 ? add_544144 : sel_544141;
  assign add_544148 = sel_544145 + 8'h01;
  assign sel_544149 = array_index_544116 == array_index_537064 ? add_544148 : sel_544145;
  assign add_544152 = sel_544149 + 8'h01;
  assign sel_544153 = array_index_544116 == array_index_537070 ? add_544152 : sel_544149;
  assign add_544156 = sel_544153 + 8'h01;
  assign sel_544157 = array_index_544116 == array_index_537076 ? add_544156 : sel_544153;
  assign add_544160 = sel_544157 + 8'h01;
  assign sel_544161 = array_index_544116 == array_index_537082 ? add_544160 : sel_544157;
  assign add_544164 = sel_544161 + 8'h01;
  assign sel_544165 = array_index_544116 == array_index_537088 ? add_544164 : sel_544161;
  assign add_544168 = sel_544165 + 8'h01;
  assign sel_544169 = array_index_544116 == array_index_537094 ? add_544168 : sel_544165;
  assign add_544172 = sel_544169 + 8'h01;
  assign sel_544173 = array_index_544116 == array_index_537100 ? add_544172 : sel_544169;
  assign add_544176 = sel_544173 + 8'h01;
  assign sel_544177 = array_index_544116 == array_index_537106 ? add_544176 : sel_544173;
  assign add_544180 = sel_544177 + 8'h01;
  assign sel_544181 = array_index_544116 == array_index_537112 ? add_544180 : sel_544177;
  assign add_544184 = sel_544181 + 8'h01;
  assign sel_544185 = array_index_544116 == array_index_537118 ? add_544184 : sel_544181;
  assign add_544188 = sel_544185 + 8'h01;
  assign sel_544189 = array_index_544116 == array_index_537124 ? add_544188 : sel_544185;
  assign add_544192 = sel_544189 + 8'h01;
  assign sel_544193 = array_index_544116 == array_index_537130 ? add_544192 : sel_544189;
  assign add_544196 = sel_544193 + 8'h01;
  assign sel_544197 = array_index_544116 == array_index_537136 ? add_544196 : sel_544193;
  assign add_544200 = sel_544197 + 8'h01;
  assign sel_544201 = array_index_544116 == array_index_537142 ? add_544200 : sel_544197;
  assign add_544204 = sel_544201 + 8'h01;
  assign sel_544205 = array_index_544116 == array_index_537148 ? add_544204 : sel_544201;
  assign add_544208 = sel_544205 + 8'h01;
  assign sel_544209 = array_index_544116 == array_index_537154 ? add_544208 : sel_544205;
  assign add_544212 = sel_544209 + 8'h01;
  assign sel_544213 = array_index_544116 == array_index_537160 ? add_544212 : sel_544209;
  assign add_544216 = sel_544213 + 8'h01;
  assign sel_544217 = array_index_544116 == array_index_537166 ? add_544216 : sel_544213;
  assign add_544220 = sel_544217 + 8'h01;
  assign sel_544221 = array_index_544116 == array_index_537172 ? add_544220 : sel_544217;
  assign add_544224 = sel_544221 + 8'h01;
  assign sel_544225 = array_index_544116 == array_index_537178 ? add_544224 : sel_544221;
  assign add_544228 = sel_544225 + 8'h01;
  assign sel_544229 = array_index_544116 == array_index_537184 ? add_544228 : sel_544225;
  assign add_544232 = sel_544229 + 8'h01;
  assign sel_544233 = array_index_544116 == array_index_537190 ? add_544232 : sel_544229;
  assign add_544236 = sel_544233 + 8'h01;
  assign sel_544237 = array_index_544116 == array_index_537196 ? add_544236 : sel_544233;
  assign add_544240 = sel_544237 + 8'h01;
  assign sel_544241 = array_index_544116 == array_index_537202 ? add_544240 : sel_544237;
  assign add_544244 = sel_544241 + 8'h01;
  assign sel_544245 = array_index_544116 == array_index_537208 ? add_544244 : sel_544241;
  assign add_544248 = sel_544245 + 8'h01;
  assign sel_544249 = array_index_544116 == array_index_537214 ? add_544248 : sel_544245;
  assign add_544252 = sel_544249 + 8'h01;
  assign sel_544253 = array_index_544116 == array_index_537220 ? add_544252 : sel_544249;
  assign add_544256 = sel_544253 + 8'h01;
  assign sel_544257 = array_index_544116 == array_index_537226 ? add_544256 : sel_544253;
  assign add_544260 = sel_544257 + 8'h01;
  assign sel_544261 = array_index_544116 == array_index_537232 ? add_544260 : sel_544257;
  assign add_544264 = sel_544261 + 8'h01;
  assign sel_544265 = array_index_544116 == array_index_537238 ? add_544264 : sel_544261;
  assign add_544268 = sel_544265 + 8'h01;
  assign sel_544269 = array_index_544116 == array_index_537244 ? add_544268 : sel_544265;
  assign add_544272 = sel_544269 + 8'h01;
  assign sel_544273 = array_index_544116 == array_index_537250 ? add_544272 : sel_544269;
  assign add_544276 = sel_544273 + 8'h01;
  assign sel_544277 = array_index_544116 == array_index_537256 ? add_544276 : sel_544273;
  assign add_544280 = sel_544277 + 8'h01;
  assign sel_544281 = array_index_544116 == array_index_537262 ? add_544280 : sel_544277;
  assign add_544284 = sel_544281 + 8'h01;
  assign sel_544285 = array_index_544116 == array_index_537268 ? add_544284 : sel_544281;
  assign add_544288 = sel_544285 + 8'h01;
  assign sel_544289 = array_index_544116 == array_index_537274 ? add_544288 : sel_544285;
  assign add_544292 = sel_544289 + 8'h01;
  assign sel_544293 = array_index_544116 == array_index_537280 ? add_544292 : sel_544289;
  assign add_544296 = sel_544293 + 8'h01;
  assign sel_544297 = array_index_544116 == array_index_537286 ? add_544296 : sel_544293;
  assign add_544300 = sel_544297 + 8'h01;
  assign sel_544301 = array_index_544116 == array_index_537292 ? add_544300 : sel_544297;
  assign add_544304 = sel_544301 + 8'h01;
  assign sel_544305 = array_index_544116 == array_index_537298 ? add_544304 : sel_544301;
  assign add_544308 = sel_544305 + 8'h01;
  assign sel_544309 = array_index_544116 == array_index_537304 ? add_544308 : sel_544305;
  assign add_544312 = sel_544309 + 8'h01;
  assign sel_544313 = array_index_544116 == array_index_537310 ? add_544312 : sel_544309;
  assign add_544316 = sel_544313 + 8'h01;
  assign sel_544317 = array_index_544116 == array_index_537316 ? add_544316 : sel_544313;
  assign add_544320 = sel_544317 + 8'h01;
  assign sel_544321 = array_index_544116 == array_index_537322 ? add_544320 : sel_544317;
  assign add_544324 = sel_544321 + 8'h01;
  assign sel_544325 = array_index_544116 == array_index_537328 ? add_544324 : sel_544321;
  assign add_544328 = sel_544325 + 8'h01;
  assign sel_544329 = array_index_544116 == array_index_537334 ? add_544328 : sel_544325;
  assign add_544332 = sel_544329 + 8'h01;
  assign sel_544333 = array_index_544116 == array_index_537340 ? add_544332 : sel_544329;
  assign add_544336 = sel_544333 + 8'h01;
  assign sel_544337 = array_index_544116 == array_index_537346 ? add_544336 : sel_544333;
  assign add_544340 = sel_544337 + 8'h01;
  assign sel_544341 = array_index_544116 == array_index_537352 ? add_544340 : sel_544337;
  assign add_544344 = sel_544341 + 8'h01;
  assign sel_544345 = array_index_544116 == array_index_537358 ? add_544344 : sel_544341;
  assign add_544348 = sel_544345 + 8'h01;
  assign sel_544349 = array_index_544116 == array_index_537364 ? add_544348 : sel_544345;
  assign add_544352 = sel_544349 + 8'h01;
  assign sel_544353 = array_index_544116 == array_index_537370 ? add_544352 : sel_544349;
  assign add_544356 = sel_544353 + 8'h01;
  assign sel_544357 = array_index_544116 == array_index_537376 ? add_544356 : sel_544353;
  assign add_544360 = sel_544357 + 8'h01;
  assign sel_544361 = array_index_544116 == array_index_537382 ? add_544360 : sel_544357;
  assign add_544364 = sel_544361 + 8'h01;
  assign sel_544365 = array_index_544116 == array_index_537388 ? add_544364 : sel_544361;
  assign add_544368 = sel_544365 + 8'h01;
  assign sel_544369 = array_index_544116 == array_index_537394 ? add_544368 : sel_544365;
  assign add_544372 = sel_544369 + 8'h01;
  assign sel_544373 = array_index_544116 == array_index_537400 ? add_544372 : sel_544369;
  assign add_544376 = sel_544373 + 8'h01;
  assign sel_544377 = array_index_544116 == array_index_537406 ? add_544376 : sel_544373;
  assign add_544380 = sel_544377 + 8'h01;
  assign sel_544381 = array_index_544116 == array_index_537412 ? add_544380 : sel_544377;
  assign add_544384 = sel_544381 + 8'h01;
  assign sel_544385 = array_index_544116 == array_index_537418 ? add_544384 : sel_544381;
  assign add_544388 = sel_544385 + 8'h01;
  assign sel_544389 = array_index_544116 == array_index_537424 ? add_544388 : sel_544385;
  assign add_544392 = sel_544389 + 8'h01;
  assign sel_544393 = array_index_544116 == array_index_537430 ? add_544392 : sel_544389;
  assign add_544396 = sel_544393 + 8'h01;
  assign sel_544397 = array_index_544116 == array_index_537436 ? add_544396 : sel_544393;
  assign add_544400 = sel_544397 + 8'h01;
  assign sel_544401 = array_index_544116 == array_index_537442 ? add_544400 : sel_544397;
  assign add_544404 = sel_544401 + 8'h01;
  assign sel_544405 = array_index_544116 == array_index_537448 ? add_544404 : sel_544401;
  assign add_544408 = sel_544405 + 8'h01;
  assign sel_544409 = array_index_544116 == array_index_537454 ? add_544408 : sel_544405;
  assign add_544412 = sel_544409 + 8'h01;
  assign sel_544413 = array_index_544116 == array_index_537460 ? add_544412 : sel_544409;
  assign add_544417 = sel_544413 + 8'h01;
  assign array_index_544418 = set1_unflattened[7'h18];
  assign sel_544419 = array_index_544116 == array_index_537466 ? add_544417 : sel_544413;
  assign add_544422 = sel_544419 + 8'h01;
  assign sel_544423 = array_index_544418 == array_index_537012 ? add_544422 : sel_544419;
  assign add_544426 = sel_544423 + 8'h01;
  assign sel_544427 = array_index_544418 == array_index_537016 ? add_544426 : sel_544423;
  assign add_544430 = sel_544427 + 8'h01;
  assign sel_544431 = array_index_544418 == array_index_537024 ? add_544430 : sel_544427;
  assign add_544434 = sel_544431 + 8'h01;
  assign sel_544435 = array_index_544418 == array_index_537032 ? add_544434 : sel_544431;
  assign add_544438 = sel_544435 + 8'h01;
  assign sel_544439 = array_index_544418 == array_index_537040 ? add_544438 : sel_544435;
  assign add_544442 = sel_544439 + 8'h01;
  assign sel_544443 = array_index_544418 == array_index_537048 ? add_544442 : sel_544439;
  assign add_544446 = sel_544443 + 8'h01;
  assign sel_544447 = array_index_544418 == array_index_537056 ? add_544446 : sel_544443;
  assign add_544450 = sel_544447 + 8'h01;
  assign sel_544451 = array_index_544418 == array_index_537064 ? add_544450 : sel_544447;
  assign add_544454 = sel_544451 + 8'h01;
  assign sel_544455 = array_index_544418 == array_index_537070 ? add_544454 : sel_544451;
  assign add_544458 = sel_544455 + 8'h01;
  assign sel_544459 = array_index_544418 == array_index_537076 ? add_544458 : sel_544455;
  assign add_544462 = sel_544459 + 8'h01;
  assign sel_544463 = array_index_544418 == array_index_537082 ? add_544462 : sel_544459;
  assign add_544466 = sel_544463 + 8'h01;
  assign sel_544467 = array_index_544418 == array_index_537088 ? add_544466 : sel_544463;
  assign add_544470 = sel_544467 + 8'h01;
  assign sel_544471 = array_index_544418 == array_index_537094 ? add_544470 : sel_544467;
  assign add_544474 = sel_544471 + 8'h01;
  assign sel_544475 = array_index_544418 == array_index_537100 ? add_544474 : sel_544471;
  assign add_544478 = sel_544475 + 8'h01;
  assign sel_544479 = array_index_544418 == array_index_537106 ? add_544478 : sel_544475;
  assign add_544482 = sel_544479 + 8'h01;
  assign sel_544483 = array_index_544418 == array_index_537112 ? add_544482 : sel_544479;
  assign add_544486 = sel_544483 + 8'h01;
  assign sel_544487 = array_index_544418 == array_index_537118 ? add_544486 : sel_544483;
  assign add_544490 = sel_544487 + 8'h01;
  assign sel_544491 = array_index_544418 == array_index_537124 ? add_544490 : sel_544487;
  assign add_544494 = sel_544491 + 8'h01;
  assign sel_544495 = array_index_544418 == array_index_537130 ? add_544494 : sel_544491;
  assign add_544498 = sel_544495 + 8'h01;
  assign sel_544499 = array_index_544418 == array_index_537136 ? add_544498 : sel_544495;
  assign add_544502 = sel_544499 + 8'h01;
  assign sel_544503 = array_index_544418 == array_index_537142 ? add_544502 : sel_544499;
  assign add_544506 = sel_544503 + 8'h01;
  assign sel_544507 = array_index_544418 == array_index_537148 ? add_544506 : sel_544503;
  assign add_544510 = sel_544507 + 8'h01;
  assign sel_544511 = array_index_544418 == array_index_537154 ? add_544510 : sel_544507;
  assign add_544514 = sel_544511 + 8'h01;
  assign sel_544515 = array_index_544418 == array_index_537160 ? add_544514 : sel_544511;
  assign add_544518 = sel_544515 + 8'h01;
  assign sel_544519 = array_index_544418 == array_index_537166 ? add_544518 : sel_544515;
  assign add_544522 = sel_544519 + 8'h01;
  assign sel_544523 = array_index_544418 == array_index_537172 ? add_544522 : sel_544519;
  assign add_544526 = sel_544523 + 8'h01;
  assign sel_544527 = array_index_544418 == array_index_537178 ? add_544526 : sel_544523;
  assign add_544530 = sel_544527 + 8'h01;
  assign sel_544531 = array_index_544418 == array_index_537184 ? add_544530 : sel_544527;
  assign add_544534 = sel_544531 + 8'h01;
  assign sel_544535 = array_index_544418 == array_index_537190 ? add_544534 : sel_544531;
  assign add_544538 = sel_544535 + 8'h01;
  assign sel_544539 = array_index_544418 == array_index_537196 ? add_544538 : sel_544535;
  assign add_544542 = sel_544539 + 8'h01;
  assign sel_544543 = array_index_544418 == array_index_537202 ? add_544542 : sel_544539;
  assign add_544546 = sel_544543 + 8'h01;
  assign sel_544547 = array_index_544418 == array_index_537208 ? add_544546 : sel_544543;
  assign add_544550 = sel_544547 + 8'h01;
  assign sel_544551 = array_index_544418 == array_index_537214 ? add_544550 : sel_544547;
  assign add_544554 = sel_544551 + 8'h01;
  assign sel_544555 = array_index_544418 == array_index_537220 ? add_544554 : sel_544551;
  assign add_544558 = sel_544555 + 8'h01;
  assign sel_544559 = array_index_544418 == array_index_537226 ? add_544558 : sel_544555;
  assign add_544562 = sel_544559 + 8'h01;
  assign sel_544563 = array_index_544418 == array_index_537232 ? add_544562 : sel_544559;
  assign add_544566 = sel_544563 + 8'h01;
  assign sel_544567 = array_index_544418 == array_index_537238 ? add_544566 : sel_544563;
  assign add_544570 = sel_544567 + 8'h01;
  assign sel_544571 = array_index_544418 == array_index_537244 ? add_544570 : sel_544567;
  assign add_544574 = sel_544571 + 8'h01;
  assign sel_544575 = array_index_544418 == array_index_537250 ? add_544574 : sel_544571;
  assign add_544578 = sel_544575 + 8'h01;
  assign sel_544579 = array_index_544418 == array_index_537256 ? add_544578 : sel_544575;
  assign add_544582 = sel_544579 + 8'h01;
  assign sel_544583 = array_index_544418 == array_index_537262 ? add_544582 : sel_544579;
  assign add_544586 = sel_544583 + 8'h01;
  assign sel_544587 = array_index_544418 == array_index_537268 ? add_544586 : sel_544583;
  assign add_544590 = sel_544587 + 8'h01;
  assign sel_544591 = array_index_544418 == array_index_537274 ? add_544590 : sel_544587;
  assign add_544594 = sel_544591 + 8'h01;
  assign sel_544595 = array_index_544418 == array_index_537280 ? add_544594 : sel_544591;
  assign add_544598 = sel_544595 + 8'h01;
  assign sel_544599 = array_index_544418 == array_index_537286 ? add_544598 : sel_544595;
  assign add_544602 = sel_544599 + 8'h01;
  assign sel_544603 = array_index_544418 == array_index_537292 ? add_544602 : sel_544599;
  assign add_544606 = sel_544603 + 8'h01;
  assign sel_544607 = array_index_544418 == array_index_537298 ? add_544606 : sel_544603;
  assign add_544610 = sel_544607 + 8'h01;
  assign sel_544611 = array_index_544418 == array_index_537304 ? add_544610 : sel_544607;
  assign add_544614 = sel_544611 + 8'h01;
  assign sel_544615 = array_index_544418 == array_index_537310 ? add_544614 : sel_544611;
  assign add_544618 = sel_544615 + 8'h01;
  assign sel_544619 = array_index_544418 == array_index_537316 ? add_544618 : sel_544615;
  assign add_544622 = sel_544619 + 8'h01;
  assign sel_544623 = array_index_544418 == array_index_537322 ? add_544622 : sel_544619;
  assign add_544626 = sel_544623 + 8'h01;
  assign sel_544627 = array_index_544418 == array_index_537328 ? add_544626 : sel_544623;
  assign add_544630 = sel_544627 + 8'h01;
  assign sel_544631 = array_index_544418 == array_index_537334 ? add_544630 : sel_544627;
  assign add_544634 = sel_544631 + 8'h01;
  assign sel_544635 = array_index_544418 == array_index_537340 ? add_544634 : sel_544631;
  assign add_544638 = sel_544635 + 8'h01;
  assign sel_544639 = array_index_544418 == array_index_537346 ? add_544638 : sel_544635;
  assign add_544642 = sel_544639 + 8'h01;
  assign sel_544643 = array_index_544418 == array_index_537352 ? add_544642 : sel_544639;
  assign add_544646 = sel_544643 + 8'h01;
  assign sel_544647 = array_index_544418 == array_index_537358 ? add_544646 : sel_544643;
  assign add_544650 = sel_544647 + 8'h01;
  assign sel_544651 = array_index_544418 == array_index_537364 ? add_544650 : sel_544647;
  assign add_544654 = sel_544651 + 8'h01;
  assign sel_544655 = array_index_544418 == array_index_537370 ? add_544654 : sel_544651;
  assign add_544658 = sel_544655 + 8'h01;
  assign sel_544659 = array_index_544418 == array_index_537376 ? add_544658 : sel_544655;
  assign add_544662 = sel_544659 + 8'h01;
  assign sel_544663 = array_index_544418 == array_index_537382 ? add_544662 : sel_544659;
  assign add_544666 = sel_544663 + 8'h01;
  assign sel_544667 = array_index_544418 == array_index_537388 ? add_544666 : sel_544663;
  assign add_544670 = sel_544667 + 8'h01;
  assign sel_544671 = array_index_544418 == array_index_537394 ? add_544670 : sel_544667;
  assign add_544674 = sel_544671 + 8'h01;
  assign sel_544675 = array_index_544418 == array_index_537400 ? add_544674 : sel_544671;
  assign add_544678 = sel_544675 + 8'h01;
  assign sel_544679 = array_index_544418 == array_index_537406 ? add_544678 : sel_544675;
  assign add_544682 = sel_544679 + 8'h01;
  assign sel_544683 = array_index_544418 == array_index_537412 ? add_544682 : sel_544679;
  assign add_544686 = sel_544683 + 8'h01;
  assign sel_544687 = array_index_544418 == array_index_537418 ? add_544686 : sel_544683;
  assign add_544690 = sel_544687 + 8'h01;
  assign sel_544691 = array_index_544418 == array_index_537424 ? add_544690 : sel_544687;
  assign add_544694 = sel_544691 + 8'h01;
  assign sel_544695 = array_index_544418 == array_index_537430 ? add_544694 : sel_544691;
  assign add_544698 = sel_544695 + 8'h01;
  assign sel_544699 = array_index_544418 == array_index_537436 ? add_544698 : sel_544695;
  assign add_544702 = sel_544699 + 8'h01;
  assign sel_544703 = array_index_544418 == array_index_537442 ? add_544702 : sel_544699;
  assign add_544706 = sel_544703 + 8'h01;
  assign sel_544707 = array_index_544418 == array_index_537448 ? add_544706 : sel_544703;
  assign add_544710 = sel_544707 + 8'h01;
  assign sel_544711 = array_index_544418 == array_index_537454 ? add_544710 : sel_544707;
  assign add_544714 = sel_544711 + 8'h01;
  assign sel_544715 = array_index_544418 == array_index_537460 ? add_544714 : sel_544711;
  assign add_544719 = sel_544715 + 8'h01;
  assign array_index_544720 = set1_unflattened[7'h19];
  assign sel_544721 = array_index_544418 == array_index_537466 ? add_544719 : sel_544715;
  assign add_544724 = sel_544721 + 8'h01;
  assign sel_544725 = array_index_544720 == array_index_537012 ? add_544724 : sel_544721;
  assign add_544728 = sel_544725 + 8'h01;
  assign sel_544729 = array_index_544720 == array_index_537016 ? add_544728 : sel_544725;
  assign add_544732 = sel_544729 + 8'h01;
  assign sel_544733 = array_index_544720 == array_index_537024 ? add_544732 : sel_544729;
  assign add_544736 = sel_544733 + 8'h01;
  assign sel_544737 = array_index_544720 == array_index_537032 ? add_544736 : sel_544733;
  assign add_544740 = sel_544737 + 8'h01;
  assign sel_544741 = array_index_544720 == array_index_537040 ? add_544740 : sel_544737;
  assign add_544744 = sel_544741 + 8'h01;
  assign sel_544745 = array_index_544720 == array_index_537048 ? add_544744 : sel_544741;
  assign add_544748 = sel_544745 + 8'h01;
  assign sel_544749 = array_index_544720 == array_index_537056 ? add_544748 : sel_544745;
  assign add_544752 = sel_544749 + 8'h01;
  assign sel_544753 = array_index_544720 == array_index_537064 ? add_544752 : sel_544749;
  assign add_544756 = sel_544753 + 8'h01;
  assign sel_544757 = array_index_544720 == array_index_537070 ? add_544756 : sel_544753;
  assign add_544760 = sel_544757 + 8'h01;
  assign sel_544761 = array_index_544720 == array_index_537076 ? add_544760 : sel_544757;
  assign add_544764 = sel_544761 + 8'h01;
  assign sel_544765 = array_index_544720 == array_index_537082 ? add_544764 : sel_544761;
  assign add_544768 = sel_544765 + 8'h01;
  assign sel_544769 = array_index_544720 == array_index_537088 ? add_544768 : sel_544765;
  assign add_544772 = sel_544769 + 8'h01;
  assign sel_544773 = array_index_544720 == array_index_537094 ? add_544772 : sel_544769;
  assign add_544776 = sel_544773 + 8'h01;
  assign sel_544777 = array_index_544720 == array_index_537100 ? add_544776 : sel_544773;
  assign add_544780 = sel_544777 + 8'h01;
  assign sel_544781 = array_index_544720 == array_index_537106 ? add_544780 : sel_544777;
  assign add_544784 = sel_544781 + 8'h01;
  assign sel_544785 = array_index_544720 == array_index_537112 ? add_544784 : sel_544781;
  assign add_544788 = sel_544785 + 8'h01;
  assign sel_544789 = array_index_544720 == array_index_537118 ? add_544788 : sel_544785;
  assign add_544792 = sel_544789 + 8'h01;
  assign sel_544793 = array_index_544720 == array_index_537124 ? add_544792 : sel_544789;
  assign add_544796 = sel_544793 + 8'h01;
  assign sel_544797 = array_index_544720 == array_index_537130 ? add_544796 : sel_544793;
  assign add_544800 = sel_544797 + 8'h01;
  assign sel_544801 = array_index_544720 == array_index_537136 ? add_544800 : sel_544797;
  assign add_544804 = sel_544801 + 8'h01;
  assign sel_544805 = array_index_544720 == array_index_537142 ? add_544804 : sel_544801;
  assign add_544808 = sel_544805 + 8'h01;
  assign sel_544809 = array_index_544720 == array_index_537148 ? add_544808 : sel_544805;
  assign add_544812 = sel_544809 + 8'h01;
  assign sel_544813 = array_index_544720 == array_index_537154 ? add_544812 : sel_544809;
  assign add_544816 = sel_544813 + 8'h01;
  assign sel_544817 = array_index_544720 == array_index_537160 ? add_544816 : sel_544813;
  assign add_544820 = sel_544817 + 8'h01;
  assign sel_544821 = array_index_544720 == array_index_537166 ? add_544820 : sel_544817;
  assign add_544824 = sel_544821 + 8'h01;
  assign sel_544825 = array_index_544720 == array_index_537172 ? add_544824 : sel_544821;
  assign add_544828 = sel_544825 + 8'h01;
  assign sel_544829 = array_index_544720 == array_index_537178 ? add_544828 : sel_544825;
  assign add_544832 = sel_544829 + 8'h01;
  assign sel_544833 = array_index_544720 == array_index_537184 ? add_544832 : sel_544829;
  assign add_544836 = sel_544833 + 8'h01;
  assign sel_544837 = array_index_544720 == array_index_537190 ? add_544836 : sel_544833;
  assign add_544840 = sel_544837 + 8'h01;
  assign sel_544841 = array_index_544720 == array_index_537196 ? add_544840 : sel_544837;
  assign add_544844 = sel_544841 + 8'h01;
  assign sel_544845 = array_index_544720 == array_index_537202 ? add_544844 : sel_544841;
  assign add_544848 = sel_544845 + 8'h01;
  assign sel_544849 = array_index_544720 == array_index_537208 ? add_544848 : sel_544845;
  assign add_544852 = sel_544849 + 8'h01;
  assign sel_544853 = array_index_544720 == array_index_537214 ? add_544852 : sel_544849;
  assign add_544856 = sel_544853 + 8'h01;
  assign sel_544857 = array_index_544720 == array_index_537220 ? add_544856 : sel_544853;
  assign add_544860 = sel_544857 + 8'h01;
  assign sel_544861 = array_index_544720 == array_index_537226 ? add_544860 : sel_544857;
  assign add_544864 = sel_544861 + 8'h01;
  assign sel_544865 = array_index_544720 == array_index_537232 ? add_544864 : sel_544861;
  assign add_544868 = sel_544865 + 8'h01;
  assign sel_544869 = array_index_544720 == array_index_537238 ? add_544868 : sel_544865;
  assign add_544872 = sel_544869 + 8'h01;
  assign sel_544873 = array_index_544720 == array_index_537244 ? add_544872 : sel_544869;
  assign add_544876 = sel_544873 + 8'h01;
  assign sel_544877 = array_index_544720 == array_index_537250 ? add_544876 : sel_544873;
  assign add_544880 = sel_544877 + 8'h01;
  assign sel_544881 = array_index_544720 == array_index_537256 ? add_544880 : sel_544877;
  assign add_544884 = sel_544881 + 8'h01;
  assign sel_544885 = array_index_544720 == array_index_537262 ? add_544884 : sel_544881;
  assign add_544888 = sel_544885 + 8'h01;
  assign sel_544889 = array_index_544720 == array_index_537268 ? add_544888 : sel_544885;
  assign add_544892 = sel_544889 + 8'h01;
  assign sel_544893 = array_index_544720 == array_index_537274 ? add_544892 : sel_544889;
  assign add_544896 = sel_544893 + 8'h01;
  assign sel_544897 = array_index_544720 == array_index_537280 ? add_544896 : sel_544893;
  assign add_544900 = sel_544897 + 8'h01;
  assign sel_544901 = array_index_544720 == array_index_537286 ? add_544900 : sel_544897;
  assign add_544904 = sel_544901 + 8'h01;
  assign sel_544905 = array_index_544720 == array_index_537292 ? add_544904 : sel_544901;
  assign add_544908 = sel_544905 + 8'h01;
  assign sel_544909 = array_index_544720 == array_index_537298 ? add_544908 : sel_544905;
  assign add_544912 = sel_544909 + 8'h01;
  assign sel_544913 = array_index_544720 == array_index_537304 ? add_544912 : sel_544909;
  assign add_544916 = sel_544913 + 8'h01;
  assign sel_544917 = array_index_544720 == array_index_537310 ? add_544916 : sel_544913;
  assign add_544920 = sel_544917 + 8'h01;
  assign sel_544921 = array_index_544720 == array_index_537316 ? add_544920 : sel_544917;
  assign add_544924 = sel_544921 + 8'h01;
  assign sel_544925 = array_index_544720 == array_index_537322 ? add_544924 : sel_544921;
  assign add_544928 = sel_544925 + 8'h01;
  assign sel_544929 = array_index_544720 == array_index_537328 ? add_544928 : sel_544925;
  assign add_544932 = sel_544929 + 8'h01;
  assign sel_544933 = array_index_544720 == array_index_537334 ? add_544932 : sel_544929;
  assign add_544936 = sel_544933 + 8'h01;
  assign sel_544937 = array_index_544720 == array_index_537340 ? add_544936 : sel_544933;
  assign add_544940 = sel_544937 + 8'h01;
  assign sel_544941 = array_index_544720 == array_index_537346 ? add_544940 : sel_544937;
  assign add_544944 = sel_544941 + 8'h01;
  assign sel_544945 = array_index_544720 == array_index_537352 ? add_544944 : sel_544941;
  assign add_544948 = sel_544945 + 8'h01;
  assign sel_544949 = array_index_544720 == array_index_537358 ? add_544948 : sel_544945;
  assign add_544952 = sel_544949 + 8'h01;
  assign sel_544953 = array_index_544720 == array_index_537364 ? add_544952 : sel_544949;
  assign add_544956 = sel_544953 + 8'h01;
  assign sel_544957 = array_index_544720 == array_index_537370 ? add_544956 : sel_544953;
  assign add_544960 = sel_544957 + 8'h01;
  assign sel_544961 = array_index_544720 == array_index_537376 ? add_544960 : sel_544957;
  assign add_544964 = sel_544961 + 8'h01;
  assign sel_544965 = array_index_544720 == array_index_537382 ? add_544964 : sel_544961;
  assign add_544968 = sel_544965 + 8'h01;
  assign sel_544969 = array_index_544720 == array_index_537388 ? add_544968 : sel_544965;
  assign add_544972 = sel_544969 + 8'h01;
  assign sel_544973 = array_index_544720 == array_index_537394 ? add_544972 : sel_544969;
  assign add_544976 = sel_544973 + 8'h01;
  assign sel_544977 = array_index_544720 == array_index_537400 ? add_544976 : sel_544973;
  assign add_544980 = sel_544977 + 8'h01;
  assign sel_544981 = array_index_544720 == array_index_537406 ? add_544980 : sel_544977;
  assign add_544984 = sel_544981 + 8'h01;
  assign sel_544985 = array_index_544720 == array_index_537412 ? add_544984 : sel_544981;
  assign add_544988 = sel_544985 + 8'h01;
  assign sel_544989 = array_index_544720 == array_index_537418 ? add_544988 : sel_544985;
  assign add_544992 = sel_544989 + 8'h01;
  assign sel_544993 = array_index_544720 == array_index_537424 ? add_544992 : sel_544989;
  assign add_544996 = sel_544993 + 8'h01;
  assign sel_544997 = array_index_544720 == array_index_537430 ? add_544996 : sel_544993;
  assign add_545000 = sel_544997 + 8'h01;
  assign sel_545001 = array_index_544720 == array_index_537436 ? add_545000 : sel_544997;
  assign add_545004 = sel_545001 + 8'h01;
  assign sel_545005 = array_index_544720 == array_index_537442 ? add_545004 : sel_545001;
  assign add_545008 = sel_545005 + 8'h01;
  assign sel_545009 = array_index_544720 == array_index_537448 ? add_545008 : sel_545005;
  assign add_545012 = sel_545009 + 8'h01;
  assign sel_545013 = array_index_544720 == array_index_537454 ? add_545012 : sel_545009;
  assign add_545016 = sel_545013 + 8'h01;
  assign sel_545017 = array_index_544720 == array_index_537460 ? add_545016 : sel_545013;
  assign add_545021 = sel_545017 + 8'h01;
  assign array_index_545022 = set1_unflattened[7'h1a];
  assign sel_545023 = array_index_544720 == array_index_537466 ? add_545021 : sel_545017;
  assign add_545026 = sel_545023 + 8'h01;
  assign sel_545027 = array_index_545022 == array_index_537012 ? add_545026 : sel_545023;
  assign add_545030 = sel_545027 + 8'h01;
  assign sel_545031 = array_index_545022 == array_index_537016 ? add_545030 : sel_545027;
  assign add_545034 = sel_545031 + 8'h01;
  assign sel_545035 = array_index_545022 == array_index_537024 ? add_545034 : sel_545031;
  assign add_545038 = sel_545035 + 8'h01;
  assign sel_545039 = array_index_545022 == array_index_537032 ? add_545038 : sel_545035;
  assign add_545042 = sel_545039 + 8'h01;
  assign sel_545043 = array_index_545022 == array_index_537040 ? add_545042 : sel_545039;
  assign add_545046 = sel_545043 + 8'h01;
  assign sel_545047 = array_index_545022 == array_index_537048 ? add_545046 : sel_545043;
  assign add_545050 = sel_545047 + 8'h01;
  assign sel_545051 = array_index_545022 == array_index_537056 ? add_545050 : sel_545047;
  assign add_545054 = sel_545051 + 8'h01;
  assign sel_545055 = array_index_545022 == array_index_537064 ? add_545054 : sel_545051;
  assign add_545058 = sel_545055 + 8'h01;
  assign sel_545059 = array_index_545022 == array_index_537070 ? add_545058 : sel_545055;
  assign add_545062 = sel_545059 + 8'h01;
  assign sel_545063 = array_index_545022 == array_index_537076 ? add_545062 : sel_545059;
  assign add_545066 = sel_545063 + 8'h01;
  assign sel_545067 = array_index_545022 == array_index_537082 ? add_545066 : sel_545063;
  assign add_545070 = sel_545067 + 8'h01;
  assign sel_545071 = array_index_545022 == array_index_537088 ? add_545070 : sel_545067;
  assign add_545074 = sel_545071 + 8'h01;
  assign sel_545075 = array_index_545022 == array_index_537094 ? add_545074 : sel_545071;
  assign add_545078 = sel_545075 + 8'h01;
  assign sel_545079 = array_index_545022 == array_index_537100 ? add_545078 : sel_545075;
  assign add_545082 = sel_545079 + 8'h01;
  assign sel_545083 = array_index_545022 == array_index_537106 ? add_545082 : sel_545079;
  assign add_545086 = sel_545083 + 8'h01;
  assign sel_545087 = array_index_545022 == array_index_537112 ? add_545086 : sel_545083;
  assign add_545090 = sel_545087 + 8'h01;
  assign sel_545091 = array_index_545022 == array_index_537118 ? add_545090 : sel_545087;
  assign add_545094 = sel_545091 + 8'h01;
  assign sel_545095 = array_index_545022 == array_index_537124 ? add_545094 : sel_545091;
  assign add_545098 = sel_545095 + 8'h01;
  assign sel_545099 = array_index_545022 == array_index_537130 ? add_545098 : sel_545095;
  assign add_545102 = sel_545099 + 8'h01;
  assign sel_545103 = array_index_545022 == array_index_537136 ? add_545102 : sel_545099;
  assign add_545106 = sel_545103 + 8'h01;
  assign sel_545107 = array_index_545022 == array_index_537142 ? add_545106 : sel_545103;
  assign add_545110 = sel_545107 + 8'h01;
  assign sel_545111 = array_index_545022 == array_index_537148 ? add_545110 : sel_545107;
  assign add_545114 = sel_545111 + 8'h01;
  assign sel_545115 = array_index_545022 == array_index_537154 ? add_545114 : sel_545111;
  assign add_545118 = sel_545115 + 8'h01;
  assign sel_545119 = array_index_545022 == array_index_537160 ? add_545118 : sel_545115;
  assign add_545122 = sel_545119 + 8'h01;
  assign sel_545123 = array_index_545022 == array_index_537166 ? add_545122 : sel_545119;
  assign add_545126 = sel_545123 + 8'h01;
  assign sel_545127 = array_index_545022 == array_index_537172 ? add_545126 : sel_545123;
  assign add_545130 = sel_545127 + 8'h01;
  assign sel_545131 = array_index_545022 == array_index_537178 ? add_545130 : sel_545127;
  assign add_545134 = sel_545131 + 8'h01;
  assign sel_545135 = array_index_545022 == array_index_537184 ? add_545134 : sel_545131;
  assign add_545138 = sel_545135 + 8'h01;
  assign sel_545139 = array_index_545022 == array_index_537190 ? add_545138 : sel_545135;
  assign add_545142 = sel_545139 + 8'h01;
  assign sel_545143 = array_index_545022 == array_index_537196 ? add_545142 : sel_545139;
  assign add_545146 = sel_545143 + 8'h01;
  assign sel_545147 = array_index_545022 == array_index_537202 ? add_545146 : sel_545143;
  assign add_545150 = sel_545147 + 8'h01;
  assign sel_545151 = array_index_545022 == array_index_537208 ? add_545150 : sel_545147;
  assign add_545154 = sel_545151 + 8'h01;
  assign sel_545155 = array_index_545022 == array_index_537214 ? add_545154 : sel_545151;
  assign add_545158 = sel_545155 + 8'h01;
  assign sel_545159 = array_index_545022 == array_index_537220 ? add_545158 : sel_545155;
  assign add_545162 = sel_545159 + 8'h01;
  assign sel_545163 = array_index_545022 == array_index_537226 ? add_545162 : sel_545159;
  assign add_545166 = sel_545163 + 8'h01;
  assign sel_545167 = array_index_545022 == array_index_537232 ? add_545166 : sel_545163;
  assign add_545170 = sel_545167 + 8'h01;
  assign sel_545171 = array_index_545022 == array_index_537238 ? add_545170 : sel_545167;
  assign add_545174 = sel_545171 + 8'h01;
  assign sel_545175 = array_index_545022 == array_index_537244 ? add_545174 : sel_545171;
  assign add_545178 = sel_545175 + 8'h01;
  assign sel_545179 = array_index_545022 == array_index_537250 ? add_545178 : sel_545175;
  assign add_545182 = sel_545179 + 8'h01;
  assign sel_545183 = array_index_545022 == array_index_537256 ? add_545182 : sel_545179;
  assign add_545186 = sel_545183 + 8'h01;
  assign sel_545187 = array_index_545022 == array_index_537262 ? add_545186 : sel_545183;
  assign add_545190 = sel_545187 + 8'h01;
  assign sel_545191 = array_index_545022 == array_index_537268 ? add_545190 : sel_545187;
  assign add_545194 = sel_545191 + 8'h01;
  assign sel_545195 = array_index_545022 == array_index_537274 ? add_545194 : sel_545191;
  assign add_545198 = sel_545195 + 8'h01;
  assign sel_545199 = array_index_545022 == array_index_537280 ? add_545198 : sel_545195;
  assign add_545202 = sel_545199 + 8'h01;
  assign sel_545203 = array_index_545022 == array_index_537286 ? add_545202 : sel_545199;
  assign add_545206 = sel_545203 + 8'h01;
  assign sel_545207 = array_index_545022 == array_index_537292 ? add_545206 : sel_545203;
  assign add_545210 = sel_545207 + 8'h01;
  assign sel_545211 = array_index_545022 == array_index_537298 ? add_545210 : sel_545207;
  assign add_545214 = sel_545211 + 8'h01;
  assign sel_545215 = array_index_545022 == array_index_537304 ? add_545214 : sel_545211;
  assign add_545218 = sel_545215 + 8'h01;
  assign sel_545219 = array_index_545022 == array_index_537310 ? add_545218 : sel_545215;
  assign add_545222 = sel_545219 + 8'h01;
  assign sel_545223 = array_index_545022 == array_index_537316 ? add_545222 : sel_545219;
  assign add_545226 = sel_545223 + 8'h01;
  assign sel_545227 = array_index_545022 == array_index_537322 ? add_545226 : sel_545223;
  assign add_545230 = sel_545227 + 8'h01;
  assign sel_545231 = array_index_545022 == array_index_537328 ? add_545230 : sel_545227;
  assign add_545234 = sel_545231 + 8'h01;
  assign sel_545235 = array_index_545022 == array_index_537334 ? add_545234 : sel_545231;
  assign add_545238 = sel_545235 + 8'h01;
  assign sel_545239 = array_index_545022 == array_index_537340 ? add_545238 : sel_545235;
  assign add_545242 = sel_545239 + 8'h01;
  assign sel_545243 = array_index_545022 == array_index_537346 ? add_545242 : sel_545239;
  assign add_545246 = sel_545243 + 8'h01;
  assign sel_545247 = array_index_545022 == array_index_537352 ? add_545246 : sel_545243;
  assign add_545250 = sel_545247 + 8'h01;
  assign sel_545251 = array_index_545022 == array_index_537358 ? add_545250 : sel_545247;
  assign add_545254 = sel_545251 + 8'h01;
  assign sel_545255 = array_index_545022 == array_index_537364 ? add_545254 : sel_545251;
  assign add_545258 = sel_545255 + 8'h01;
  assign sel_545259 = array_index_545022 == array_index_537370 ? add_545258 : sel_545255;
  assign add_545262 = sel_545259 + 8'h01;
  assign sel_545263 = array_index_545022 == array_index_537376 ? add_545262 : sel_545259;
  assign add_545266 = sel_545263 + 8'h01;
  assign sel_545267 = array_index_545022 == array_index_537382 ? add_545266 : sel_545263;
  assign add_545270 = sel_545267 + 8'h01;
  assign sel_545271 = array_index_545022 == array_index_537388 ? add_545270 : sel_545267;
  assign add_545274 = sel_545271 + 8'h01;
  assign sel_545275 = array_index_545022 == array_index_537394 ? add_545274 : sel_545271;
  assign add_545278 = sel_545275 + 8'h01;
  assign sel_545279 = array_index_545022 == array_index_537400 ? add_545278 : sel_545275;
  assign add_545282 = sel_545279 + 8'h01;
  assign sel_545283 = array_index_545022 == array_index_537406 ? add_545282 : sel_545279;
  assign add_545286 = sel_545283 + 8'h01;
  assign sel_545287 = array_index_545022 == array_index_537412 ? add_545286 : sel_545283;
  assign add_545290 = sel_545287 + 8'h01;
  assign sel_545291 = array_index_545022 == array_index_537418 ? add_545290 : sel_545287;
  assign add_545294 = sel_545291 + 8'h01;
  assign sel_545295 = array_index_545022 == array_index_537424 ? add_545294 : sel_545291;
  assign add_545298 = sel_545295 + 8'h01;
  assign sel_545299 = array_index_545022 == array_index_537430 ? add_545298 : sel_545295;
  assign add_545302 = sel_545299 + 8'h01;
  assign sel_545303 = array_index_545022 == array_index_537436 ? add_545302 : sel_545299;
  assign add_545306 = sel_545303 + 8'h01;
  assign sel_545307 = array_index_545022 == array_index_537442 ? add_545306 : sel_545303;
  assign add_545310 = sel_545307 + 8'h01;
  assign sel_545311 = array_index_545022 == array_index_537448 ? add_545310 : sel_545307;
  assign add_545314 = sel_545311 + 8'h01;
  assign sel_545315 = array_index_545022 == array_index_537454 ? add_545314 : sel_545311;
  assign add_545318 = sel_545315 + 8'h01;
  assign sel_545319 = array_index_545022 == array_index_537460 ? add_545318 : sel_545315;
  assign add_545323 = sel_545319 + 8'h01;
  assign array_index_545324 = set1_unflattened[7'h1b];
  assign sel_545325 = array_index_545022 == array_index_537466 ? add_545323 : sel_545319;
  assign add_545328 = sel_545325 + 8'h01;
  assign sel_545329 = array_index_545324 == array_index_537012 ? add_545328 : sel_545325;
  assign add_545332 = sel_545329 + 8'h01;
  assign sel_545333 = array_index_545324 == array_index_537016 ? add_545332 : sel_545329;
  assign add_545336 = sel_545333 + 8'h01;
  assign sel_545337 = array_index_545324 == array_index_537024 ? add_545336 : sel_545333;
  assign add_545340 = sel_545337 + 8'h01;
  assign sel_545341 = array_index_545324 == array_index_537032 ? add_545340 : sel_545337;
  assign add_545344 = sel_545341 + 8'h01;
  assign sel_545345 = array_index_545324 == array_index_537040 ? add_545344 : sel_545341;
  assign add_545348 = sel_545345 + 8'h01;
  assign sel_545349 = array_index_545324 == array_index_537048 ? add_545348 : sel_545345;
  assign add_545352 = sel_545349 + 8'h01;
  assign sel_545353 = array_index_545324 == array_index_537056 ? add_545352 : sel_545349;
  assign add_545356 = sel_545353 + 8'h01;
  assign sel_545357 = array_index_545324 == array_index_537064 ? add_545356 : sel_545353;
  assign add_545360 = sel_545357 + 8'h01;
  assign sel_545361 = array_index_545324 == array_index_537070 ? add_545360 : sel_545357;
  assign add_545364 = sel_545361 + 8'h01;
  assign sel_545365 = array_index_545324 == array_index_537076 ? add_545364 : sel_545361;
  assign add_545368 = sel_545365 + 8'h01;
  assign sel_545369 = array_index_545324 == array_index_537082 ? add_545368 : sel_545365;
  assign add_545372 = sel_545369 + 8'h01;
  assign sel_545373 = array_index_545324 == array_index_537088 ? add_545372 : sel_545369;
  assign add_545376 = sel_545373 + 8'h01;
  assign sel_545377 = array_index_545324 == array_index_537094 ? add_545376 : sel_545373;
  assign add_545380 = sel_545377 + 8'h01;
  assign sel_545381 = array_index_545324 == array_index_537100 ? add_545380 : sel_545377;
  assign add_545384 = sel_545381 + 8'h01;
  assign sel_545385 = array_index_545324 == array_index_537106 ? add_545384 : sel_545381;
  assign add_545388 = sel_545385 + 8'h01;
  assign sel_545389 = array_index_545324 == array_index_537112 ? add_545388 : sel_545385;
  assign add_545392 = sel_545389 + 8'h01;
  assign sel_545393 = array_index_545324 == array_index_537118 ? add_545392 : sel_545389;
  assign add_545396 = sel_545393 + 8'h01;
  assign sel_545397 = array_index_545324 == array_index_537124 ? add_545396 : sel_545393;
  assign add_545400 = sel_545397 + 8'h01;
  assign sel_545401 = array_index_545324 == array_index_537130 ? add_545400 : sel_545397;
  assign add_545404 = sel_545401 + 8'h01;
  assign sel_545405 = array_index_545324 == array_index_537136 ? add_545404 : sel_545401;
  assign add_545408 = sel_545405 + 8'h01;
  assign sel_545409 = array_index_545324 == array_index_537142 ? add_545408 : sel_545405;
  assign add_545412 = sel_545409 + 8'h01;
  assign sel_545413 = array_index_545324 == array_index_537148 ? add_545412 : sel_545409;
  assign add_545416 = sel_545413 + 8'h01;
  assign sel_545417 = array_index_545324 == array_index_537154 ? add_545416 : sel_545413;
  assign add_545420 = sel_545417 + 8'h01;
  assign sel_545421 = array_index_545324 == array_index_537160 ? add_545420 : sel_545417;
  assign add_545424 = sel_545421 + 8'h01;
  assign sel_545425 = array_index_545324 == array_index_537166 ? add_545424 : sel_545421;
  assign add_545428 = sel_545425 + 8'h01;
  assign sel_545429 = array_index_545324 == array_index_537172 ? add_545428 : sel_545425;
  assign add_545432 = sel_545429 + 8'h01;
  assign sel_545433 = array_index_545324 == array_index_537178 ? add_545432 : sel_545429;
  assign add_545436 = sel_545433 + 8'h01;
  assign sel_545437 = array_index_545324 == array_index_537184 ? add_545436 : sel_545433;
  assign add_545440 = sel_545437 + 8'h01;
  assign sel_545441 = array_index_545324 == array_index_537190 ? add_545440 : sel_545437;
  assign add_545444 = sel_545441 + 8'h01;
  assign sel_545445 = array_index_545324 == array_index_537196 ? add_545444 : sel_545441;
  assign add_545448 = sel_545445 + 8'h01;
  assign sel_545449 = array_index_545324 == array_index_537202 ? add_545448 : sel_545445;
  assign add_545452 = sel_545449 + 8'h01;
  assign sel_545453 = array_index_545324 == array_index_537208 ? add_545452 : sel_545449;
  assign add_545456 = sel_545453 + 8'h01;
  assign sel_545457 = array_index_545324 == array_index_537214 ? add_545456 : sel_545453;
  assign add_545460 = sel_545457 + 8'h01;
  assign sel_545461 = array_index_545324 == array_index_537220 ? add_545460 : sel_545457;
  assign add_545464 = sel_545461 + 8'h01;
  assign sel_545465 = array_index_545324 == array_index_537226 ? add_545464 : sel_545461;
  assign add_545468 = sel_545465 + 8'h01;
  assign sel_545469 = array_index_545324 == array_index_537232 ? add_545468 : sel_545465;
  assign add_545472 = sel_545469 + 8'h01;
  assign sel_545473 = array_index_545324 == array_index_537238 ? add_545472 : sel_545469;
  assign add_545476 = sel_545473 + 8'h01;
  assign sel_545477 = array_index_545324 == array_index_537244 ? add_545476 : sel_545473;
  assign add_545480 = sel_545477 + 8'h01;
  assign sel_545481 = array_index_545324 == array_index_537250 ? add_545480 : sel_545477;
  assign add_545484 = sel_545481 + 8'h01;
  assign sel_545485 = array_index_545324 == array_index_537256 ? add_545484 : sel_545481;
  assign add_545488 = sel_545485 + 8'h01;
  assign sel_545489 = array_index_545324 == array_index_537262 ? add_545488 : sel_545485;
  assign add_545492 = sel_545489 + 8'h01;
  assign sel_545493 = array_index_545324 == array_index_537268 ? add_545492 : sel_545489;
  assign add_545496 = sel_545493 + 8'h01;
  assign sel_545497 = array_index_545324 == array_index_537274 ? add_545496 : sel_545493;
  assign add_545500 = sel_545497 + 8'h01;
  assign sel_545501 = array_index_545324 == array_index_537280 ? add_545500 : sel_545497;
  assign add_545504 = sel_545501 + 8'h01;
  assign sel_545505 = array_index_545324 == array_index_537286 ? add_545504 : sel_545501;
  assign add_545508 = sel_545505 + 8'h01;
  assign sel_545509 = array_index_545324 == array_index_537292 ? add_545508 : sel_545505;
  assign add_545512 = sel_545509 + 8'h01;
  assign sel_545513 = array_index_545324 == array_index_537298 ? add_545512 : sel_545509;
  assign add_545516 = sel_545513 + 8'h01;
  assign sel_545517 = array_index_545324 == array_index_537304 ? add_545516 : sel_545513;
  assign add_545520 = sel_545517 + 8'h01;
  assign sel_545521 = array_index_545324 == array_index_537310 ? add_545520 : sel_545517;
  assign add_545524 = sel_545521 + 8'h01;
  assign sel_545525 = array_index_545324 == array_index_537316 ? add_545524 : sel_545521;
  assign add_545528 = sel_545525 + 8'h01;
  assign sel_545529 = array_index_545324 == array_index_537322 ? add_545528 : sel_545525;
  assign add_545532 = sel_545529 + 8'h01;
  assign sel_545533 = array_index_545324 == array_index_537328 ? add_545532 : sel_545529;
  assign add_545536 = sel_545533 + 8'h01;
  assign sel_545537 = array_index_545324 == array_index_537334 ? add_545536 : sel_545533;
  assign add_545540 = sel_545537 + 8'h01;
  assign sel_545541 = array_index_545324 == array_index_537340 ? add_545540 : sel_545537;
  assign add_545544 = sel_545541 + 8'h01;
  assign sel_545545 = array_index_545324 == array_index_537346 ? add_545544 : sel_545541;
  assign add_545548 = sel_545545 + 8'h01;
  assign sel_545549 = array_index_545324 == array_index_537352 ? add_545548 : sel_545545;
  assign add_545552 = sel_545549 + 8'h01;
  assign sel_545553 = array_index_545324 == array_index_537358 ? add_545552 : sel_545549;
  assign add_545556 = sel_545553 + 8'h01;
  assign sel_545557 = array_index_545324 == array_index_537364 ? add_545556 : sel_545553;
  assign add_545560 = sel_545557 + 8'h01;
  assign sel_545561 = array_index_545324 == array_index_537370 ? add_545560 : sel_545557;
  assign add_545564 = sel_545561 + 8'h01;
  assign sel_545565 = array_index_545324 == array_index_537376 ? add_545564 : sel_545561;
  assign add_545568 = sel_545565 + 8'h01;
  assign sel_545569 = array_index_545324 == array_index_537382 ? add_545568 : sel_545565;
  assign add_545572 = sel_545569 + 8'h01;
  assign sel_545573 = array_index_545324 == array_index_537388 ? add_545572 : sel_545569;
  assign add_545576 = sel_545573 + 8'h01;
  assign sel_545577 = array_index_545324 == array_index_537394 ? add_545576 : sel_545573;
  assign add_545580 = sel_545577 + 8'h01;
  assign sel_545581 = array_index_545324 == array_index_537400 ? add_545580 : sel_545577;
  assign add_545584 = sel_545581 + 8'h01;
  assign sel_545585 = array_index_545324 == array_index_537406 ? add_545584 : sel_545581;
  assign add_545588 = sel_545585 + 8'h01;
  assign sel_545589 = array_index_545324 == array_index_537412 ? add_545588 : sel_545585;
  assign add_545592 = sel_545589 + 8'h01;
  assign sel_545593 = array_index_545324 == array_index_537418 ? add_545592 : sel_545589;
  assign add_545596 = sel_545593 + 8'h01;
  assign sel_545597 = array_index_545324 == array_index_537424 ? add_545596 : sel_545593;
  assign add_545600 = sel_545597 + 8'h01;
  assign sel_545601 = array_index_545324 == array_index_537430 ? add_545600 : sel_545597;
  assign add_545604 = sel_545601 + 8'h01;
  assign sel_545605 = array_index_545324 == array_index_537436 ? add_545604 : sel_545601;
  assign add_545608 = sel_545605 + 8'h01;
  assign sel_545609 = array_index_545324 == array_index_537442 ? add_545608 : sel_545605;
  assign add_545612 = sel_545609 + 8'h01;
  assign sel_545613 = array_index_545324 == array_index_537448 ? add_545612 : sel_545609;
  assign add_545616 = sel_545613 + 8'h01;
  assign sel_545617 = array_index_545324 == array_index_537454 ? add_545616 : sel_545613;
  assign add_545620 = sel_545617 + 8'h01;
  assign sel_545621 = array_index_545324 == array_index_537460 ? add_545620 : sel_545617;
  assign add_545625 = sel_545621 + 8'h01;
  assign array_index_545626 = set1_unflattened[7'h1c];
  assign sel_545627 = array_index_545324 == array_index_537466 ? add_545625 : sel_545621;
  assign add_545630 = sel_545627 + 8'h01;
  assign sel_545631 = array_index_545626 == array_index_537012 ? add_545630 : sel_545627;
  assign add_545634 = sel_545631 + 8'h01;
  assign sel_545635 = array_index_545626 == array_index_537016 ? add_545634 : sel_545631;
  assign add_545638 = sel_545635 + 8'h01;
  assign sel_545639 = array_index_545626 == array_index_537024 ? add_545638 : sel_545635;
  assign add_545642 = sel_545639 + 8'h01;
  assign sel_545643 = array_index_545626 == array_index_537032 ? add_545642 : sel_545639;
  assign add_545646 = sel_545643 + 8'h01;
  assign sel_545647 = array_index_545626 == array_index_537040 ? add_545646 : sel_545643;
  assign add_545650 = sel_545647 + 8'h01;
  assign sel_545651 = array_index_545626 == array_index_537048 ? add_545650 : sel_545647;
  assign add_545654 = sel_545651 + 8'h01;
  assign sel_545655 = array_index_545626 == array_index_537056 ? add_545654 : sel_545651;
  assign add_545658 = sel_545655 + 8'h01;
  assign sel_545659 = array_index_545626 == array_index_537064 ? add_545658 : sel_545655;
  assign add_545662 = sel_545659 + 8'h01;
  assign sel_545663 = array_index_545626 == array_index_537070 ? add_545662 : sel_545659;
  assign add_545666 = sel_545663 + 8'h01;
  assign sel_545667 = array_index_545626 == array_index_537076 ? add_545666 : sel_545663;
  assign add_545670 = sel_545667 + 8'h01;
  assign sel_545671 = array_index_545626 == array_index_537082 ? add_545670 : sel_545667;
  assign add_545674 = sel_545671 + 8'h01;
  assign sel_545675 = array_index_545626 == array_index_537088 ? add_545674 : sel_545671;
  assign add_545678 = sel_545675 + 8'h01;
  assign sel_545679 = array_index_545626 == array_index_537094 ? add_545678 : sel_545675;
  assign add_545682 = sel_545679 + 8'h01;
  assign sel_545683 = array_index_545626 == array_index_537100 ? add_545682 : sel_545679;
  assign add_545686 = sel_545683 + 8'h01;
  assign sel_545687 = array_index_545626 == array_index_537106 ? add_545686 : sel_545683;
  assign add_545690 = sel_545687 + 8'h01;
  assign sel_545691 = array_index_545626 == array_index_537112 ? add_545690 : sel_545687;
  assign add_545694 = sel_545691 + 8'h01;
  assign sel_545695 = array_index_545626 == array_index_537118 ? add_545694 : sel_545691;
  assign add_545698 = sel_545695 + 8'h01;
  assign sel_545699 = array_index_545626 == array_index_537124 ? add_545698 : sel_545695;
  assign add_545702 = sel_545699 + 8'h01;
  assign sel_545703 = array_index_545626 == array_index_537130 ? add_545702 : sel_545699;
  assign add_545706 = sel_545703 + 8'h01;
  assign sel_545707 = array_index_545626 == array_index_537136 ? add_545706 : sel_545703;
  assign add_545710 = sel_545707 + 8'h01;
  assign sel_545711 = array_index_545626 == array_index_537142 ? add_545710 : sel_545707;
  assign add_545714 = sel_545711 + 8'h01;
  assign sel_545715 = array_index_545626 == array_index_537148 ? add_545714 : sel_545711;
  assign add_545718 = sel_545715 + 8'h01;
  assign sel_545719 = array_index_545626 == array_index_537154 ? add_545718 : sel_545715;
  assign add_545722 = sel_545719 + 8'h01;
  assign sel_545723 = array_index_545626 == array_index_537160 ? add_545722 : sel_545719;
  assign add_545726 = sel_545723 + 8'h01;
  assign sel_545727 = array_index_545626 == array_index_537166 ? add_545726 : sel_545723;
  assign add_545730 = sel_545727 + 8'h01;
  assign sel_545731 = array_index_545626 == array_index_537172 ? add_545730 : sel_545727;
  assign add_545734 = sel_545731 + 8'h01;
  assign sel_545735 = array_index_545626 == array_index_537178 ? add_545734 : sel_545731;
  assign add_545738 = sel_545735 + 8'h01;
  assign sel_545739 = array_index_545626 == array_index_537184 ? add_545738 : sel_545735;
  assign add_545742 = sel_545739 + 8'h01;
  assign sel_545743 = array_index_545626 == array_index_537190 ? add_545742 : sel_545739;
  assign add_545746 = sel_545743 + 8'h01;
  assign sel_545747 = array_index_545626 == array_index_537196 ? add_545746 : sel_545743;
  assign add_545750 = sel_545747 + 8'h01;
  assign sel_545751 = array_index_545626 == array_index_537202 ? add_545750 : sel_545747;
  assign add_545754 = sel_545751 + 8'h01;
  assign sel_545755 = array_index_545626 == array_index_537208 ? add_545754 : sel_545751;
  assign add_545758 = sel_545755 + 8'h01;
  assign sel_545759 = array_index_545626 == array_index_537214 ? add_545758 : sel_545755;
  assign add_545762 = sel_545759 + 8'h01;
  assign sel_545763 = array_index_545626 == array_index_537220 ? add_545762 : sel_545759;
  assign add_545766 = sel_545763 + 8'h01;
  assign sel_545767 = array_index_545626 == array_index_537226 ? add_545766 : sel_545763;
  assign add_545770 = sel_545767 + 8'h01;
  assign sel_545771 = array_index_545626 == array_index_537232 ? add_545770 : sel_545767;
  assign add_545774 = sel_545771 + 8'h01;
  assign sel_545775 = array_index_545626 == array_index_537238 ? add_545774 : sel_545771;
  assign add_545778 = sel_545775 + 8'h01;
  assign sel_545779 = array_index_545626 == array_index_537244 ? add_545778 : sel_545775;
  assign add_545782 = sel_545779 + 8'h01;
  assign sel_545783 = array_index_545626 == array_index_537250 ? add_545782 : sel_545779;
  assign add_545786 = sel_545783 + 8'h01;
  assign sel_545787 = array_index_545626 == array_index_537256 ? add_545786 : sel_545783;
  assign add_545790 = sel_545787 + 8'h01;
  assign sel_545791 = array_index_545626 == array_index_537262 ? add_545790 : sel_545787;
  assign add_545794 = sel_545791 + 8'h01;
  assign sel_545795 = array_index_545626 == array_index_537268 ? add_545794 : sel_545791;
  assign add_545798 = sel_545795 + 8'h01;
  assign sel_545799 = array_index_545626 == array_index_537274 ? add_545798 : sel_545795;
  assign add_545802 = sel_545799 + 8'h01;
  assign sel_545803 = array_index_545626 == array_index_537280 ? add_545802 : sel_545799;
  assign add_545806 = sel_545803 + 8'h01;
  assign sel_545807 = array_index_545626 == array_index_537286 ? add_545806 : sel_545803;
  assign add_545810 = sel_545807 + 8'h01;
  assign sel_545811 = array_index_545626 == array_index_537292 ? add_545810 : sel_545807;
  assign add_545814 = sel_545811 + 8'h01;
  assign sel_545815 = array_index_545626 == array_index_537298 ? add_545814 : sel_545811;
  assign add_545818 = sel_545815 + 8'h01;
  assign sel_545819 = array_index_545626 == array_index_537304 ? add_545818 : sel_545815;
  assign add_545822 = sel_545819 + 8'h01;
  assign sel_545823 = array_index_545626 == array_index_537310 ? add_545822 : sel_545819;
  assign add_545826 = sel_545823 + 8'h01;
  assign sel_545827 = array_index_545626 == array_index_537316 ? add_545826 : sel_545823;
  assign add_545830 = sel_545827 + 8'h01;
  assign sel_545831 = array_index_545626 == array_index_537322 ? add_545830 : sel_545827;
  assign add_545834 = sel_545831 + 8'h01;
  assign sel_545835 = array_index_545626 == array_index_537328 ? add_545834 : sel_545831;
  assign add_545838 = sel_545835 + 8'h01;
  assign sel_545839 = array_index_545626 == array_index_537334 ? add_545838 : sel_545835;
  assign add_545842 = sel_545839 + 8'h01;
  assign sel_545843 = array_index_545626 == array_index_537340 ? add_545842 : sel_545839;
  assign add_545846 = sel_545843 + 8'h01;
  assign sel_545847 = array_index_545626 == array_index_537346 ? add_545846 : sel_545843;
  assign add_545850 = sel_545847 + 8'h01;
  assign sel_545851 = array_index_545626 == array_index_537352 ? add_545850 : sel_545847;
  assign add_545854 = sel_545851 + 8'h01;
  assign sel_545855 = array_index_545626 == array_index_537358 ? add_545854 : sel_545851;
  assign add_545858 = sel_545855 + 8'h01;
  assign sel_545859 = array_index_545626 == array_index_537364 ? add_545858 : sel_545855;
  assign add_545862 = sel_545859 + 8'h01;
  assign sel_545863 = array_index_545626 == array_index_537370 ? add_545862 : sel_545859;
  assign add_545866 = sel_545863 + 8'h01;
  assign sel_545867 = array_index_545626 == array_index_537376 ? add_545866 : sel_545863;
  assign add_545870 = sel_545867 + 8'h01;
  assign sel_545871 = array_index_545626 == array_index_537382 ? add_545870 : sel_545867;
  assign add_545874 = sel_545871 + 8'h01;
  assign sel_545875 = array_index_545626 == array_index_537388 ? add_545874 : sel_545871;
  assign add_545878 = sel_545875 + 8'h01;
  assign sel_545879 = array_index_545626 == array_index_537394 ? add_545878 : sel_545875;
  assign add_545882 = sel_545879 + 8'h01;
  assign sel_545883 = array_index_545626 == array_index_537400 ? add_545882 : sel_545879;
  assign add_545886 = sel_545883 + 8'h01;
  assign sel_545887 = array_index_545626 == array_index_537406 ? add_545886 : sel_545883;
  assign add_545890 = sel_545887 + 8'h01;
  assign sel_545891 = array_index_545626 == array_index_537412 ? add_545890 : sel_545887;
  assign add_545894 = sel_545891 + 8'h01;
  assign sel_545895 = array_index_545626 == array_index_537418 ? add_545894 : sel_545891;
  assign add_545898 = sel_545895 + 8'h01;
  assign sel_545899 = array_index_545626 == array_index_537424 ? add_545898 : sel_545895;
  assign add_545902 = sel_545899 + 8'h01;
  assign sel_545903 = array_index_545626 == array_index_537430 ? add_545902 : sel_545899;
  assign add_545906 = sel_545903 + 8'h01;
  assign sel_545907 = array_index_545626 == array_index_537436 ? add_545906 : sel_545903;
  assign add_545910 = sel_545907 + 8'h01;
  assign sel_545911 = array_index_545626 == array_index_537442 ? add_545910 : sel_545907;
  assign add_545914 = sel_545911 + 8'h01;
  assign sel_545915 = array_index_545626 == array_index_537448 ? add_545914 : sel_545911;
  assign add_545918 = sel_545915 + 8'h01;
  assign sel_545919 = array_index_545626 == array_index_537454 ? add_545918 : sel_545915;
  assign add_545922 = sel_545919 + 8'h01;
  assign sel_545923 = array_index_545626 == array_index_537460 ? add_545922 : sel_545919;
  assign add_545927 = sel_545923 + 8'h01;
  assign array_index_545928 = set1_unflattened[7'h1d];
  assign sel_545929 = array_index_545626 == array_index_537466 ? add_545927 : sel_545923;
  assign add_545932 = sel_545929 + 8'h01;
  assign sel_545933 = array_index_545928 == array_index_537012 ? add_545932 : sel_545929;
  assign add_545936 = sel_545933 + 8'h01;
  assign sel_545937 = array_index_545928 == array_index_537016 ? add_545936 : sel_545933;
  assign add_545940 = sel_545937 + 8'h01;
  assign sel_545941 = array_index_545928 == array_index_537024 ? add_545940 : sel_545937;
  assign add_545944 = sel_545941 + 8'h01;
  assign sel_545945 = array_index_545928 == array_index_537032 ? add_545944 : sel_545941;
  assign add_545948 = sel_545945 + 8'h01;
  assign sel_545949 = array_index_545928 == array_index_537040 ? add_545948 : sel_545945;
  assign add_545952 = sel_545949 + 8'h01;
  assign sel_545953 = array_index_545928 == array_index_537048 ? add_545952 : sel_545949;
  assign add_545956 = sel_545953 + 8'h01;
  assign sel_545957 = array_index_545928 == array_index_537056 ? add_545956 : sel_545953;
  assign add_545960 = sel_545957 + 8'h01;
  assign sel_545961 = array_index_545928 == array_index_537064 ? add_545960 : sel_545957;
  assign add_545964 = sel_545961 + 8'h01;
  assign sel_545965 = array_index_545928 == array_index_537070 ? add_545964 : sel_545961;
  assign add_545968 = sel_545965 + 8'h01;
  assign sel_545969 = array_index_545928 == array_index_537076 ? add_545968 : sel_545965;
  assign add_545972 = sel_545969 + 8'h01;
  assign sel_545973 = array_index_545928 == array_index_537082 ? add_545972 : sel_545969;
  assign add_545976 = sel_545973 + 8'h01;
  assign sel_545977 = array_index_545928 == array_index_537088 ? add_545976 : sel_545973;
  assign add_545980 = sel_545977 + 8'h01;
  assign sel_545981 = array_index_545928 == array_index_537094 ? add_545980 : sel_545977;
  assign add_545984 = sel_545981 + 8'h01;
  assign sel_545985 = array_index_545928 == array_index_537100 ? add_545984 : sel_545981;
  assign add_545988 = sel_545985 + 8'h01;
  assign sel_545989 = array_index_545928 == array_index_537106 ? add_545988 : sel_545985;
  assign add_545992 = sel_545989 + 8'h01;
  assign sel_545993 = array_index_545928 == array_index_537112 ? add_545992 : sel_545989;
  assign add_545996 = sel_545993 + 8'h01;
  assign sel_545997 = array_index_545928 == array_index_537118 ? add_545996 : sel_545993;
  assign add_546000 = sel_545997 + 8'h01;
  assign sel_546001 = array_index_545928 == array_index_537124 ? add_546000 : sel_545997;
  assign add_546004 = sel_546001 + 8'h01;
  assign sel_546005 = array_index_545928 == array_index_537130 ? add_546004 : sel_546001;
  assign add_546008 = sel_546005 + 8'h01;
  assign sel_546009 = array_index_545928 == array_index_537136 ? add_546008 : sel_546005;
  assign add_546012 = sel_546009 + 8'h01;
  assign sel_546013 = array_index_545928 == array_index_537142 ? add_546012 : sel_546009;
  assign add_546016 = sel_546013 + 8'h01;
  assign sel_546017 = array_index_545928 == array_index_537148 ? add_546016 : sel_546013;
  assign add_546020 = sel_546017 + 8'h01;
  assign sel_546021 = array_index_545928 == array_index_537154 ? add_546020 : sel_546017;
  assign add_546024 = sel_546021 + 8'h01;
  assign sel_546025 = array_index_545928 == array_index_537160 ? add_546024 : sel_546021;
  assign add_546028 = sel_546025 + 8'h01;
  assign sel_546029 = array_index_545928 == array_index_537166 ? add_546028 : sel_546025;
  assign add_546032 = sel_546029 + 8'h01;
  assign sel_546033 = array_index_545928 == array_index_537172 ? add_546032 : sel_546029;
  assign add_546036 = sel_546033 + 8'h01;
  assign sel_546037 = array_index_545928 == array_index_537178 ? add_546036 : sel_546033;
  assign add_546040 = sel_546037 + 8'h01;
  assign sel_546041 = array_index_545928 == array_index_537184 ? add_546040 : sel_546037;
  assign add_546044 = sel_546041 + 8'h01;
  assign sel_546045 = array_index_545928 == array_index_537190 ? add_546044 : sel_546041;
  assign add_546048 = sel_546045 + 8'h01;
  assign sel_546049 = array_index_545928 == array_index_537196 ? add_546048 : sel_546045;
  assign add_546052 = sel_546049 + 8'h01;
  assign sel_546053 = array_index_545928 == array_index_537202 ? add_546052 : sel_546049;
  assign add_546056 = sel_546053 + 8'h01;
  assign sel_546057 = array_index_545928 == array_index_537208 ? add_546056 : sel_546053;
  assign add_546060 = sel_546057 + 8'h01;
  assign sel_546061 = array_index_545928 == array_index_537214 ? add_546060 : sel_546057;
  assign add_546064 = sel_546061 + 8'h01;
  assign sel_546065 = array_index_545928 == array_index_537220 ? add_546064 : sel_546061;
  assign add_546068 = sel_546065 + 8'h01;
  assign sel_546069 = array_index_545928 == array_index_537226 ? add_546068 : sel_546065;
  assign add_546072 = sel_546069 + 8'h01;
  assign sel_546073 = array_index_545928 == array_index_537232 ? add_546072 : sel_546069;
  assign add_546076 = sel_546073 + 8'h01;
  assign sel_546077 = array_index_545928 == array_index_537238 ? add_546076 : sel_546073;
  assign add_546080 = sel_546077 + 8'h01;
  assign sel_546081 = array_index_545928 == array_index_537244 ? add_546080 : sel_546077;
  assign add_546084 = sel_546081 + 8'h01;
  assign sel_546085 = array_index_545928 == array_index_537250 ? add_546084 : sel_546081;
  assign add_546088 = sel_546085 + 8'h01;
  assign sel_546089 = array_index_545928 == array_index_537256 ? add_546088 : sel_546085;
  assign add_546092 = sel_546089 + 8'h01;
  assign sel_546093 = array_index_545928 == array_index_537262 ? add_546092 : sel_546089;
  assign add_546096 = sel_546093 + 8'h01;
  assign sel_546097 = array_index_545928 == array_index_537268 ? add_546096 : sel_546093;
  assign add_546100 = sel_546097 + 8'h01;
  assign sel_546101 = array_index_545928 == array_index_537274 ? add_546100 : sel_546097;
  assign add_546104 = sel_546101 + 8'h01;
  assign sel_546105 = array_index_545928 == array_index_537280 ? add_546104 : sel_546101;
  assign add_546108 = sel_546105 + 8'h01;
  assign sel_546109 = array_index_545928 == array_index_537286 ? add_546108 : sel_546105;
  assign add_546112 = sel_546109 + 8'h01;
  assign sel_546113 = array_index_545928 == array_index_537292 ? add_546112 : sel_546109;
  assign add_546116 = sel_546113 + 8'h01;
  assign sel_546117 = array_index_545928 == array_index_537298 ? add_546116 : sel_546113;
  assign add_546120 = sel_546117 + 8'h01;
  assign sel_546121 = array_index_545928 == array_index_537304 ? add_546120 : sel_546117;
  assign add_546124 = sel_546121 + 8'h01;
  assign sel_546125 = array_index_545928 == array_index_537310 ? add_546124 : sel_546121;
  assign add_546128 = sel_546125 + 8'h01;
  assign sel_546129 = array_index_545928 == array_index_537316 ? add_546128 : sel_546125;
  assign add_546132 = sel_546129 + 8'h01;
  assign sel_546133 = array_index_545928 == array_index_537322 ? add_546132 : sel_546129;
  assign add_546136 = sel_546133 + 8'h01;
  assign sel_546137 = array_index_545928 == array_index_537328 ? add_546136 : sel_546133;
  assign add_546140 = sel_546137 + 8'h01;
  assign sel_546141 = array_index_545928 == array_index_537334 ? add_546140 : sel_546137;
  assign add_546144 = sel_546141 + 8'h01;
  assign sel_546145 = array_index_545928 == array_index_537340 ? add_546144 : sel_546141;
  assign add_546148 = sel_546145 + 8'h01;
  assign sel_546149 = array_index_545928 == array_index_537346 ? add_546148 : sel_546145;
  assign add_546152 = sel_546149 + 8'h01;
  assign sel_546153 = array_index_545928 == array_index_537352 ? add_546152 : sel_546149;
  assign add_546156 = sel_546153 + 8'h01;
  assign sel_546157 = array_index_545928 == array_index_537358 ? add_546156 : sel_546153;
  assign add_546160 = sel_546157 + 8'h01;
  assign sel_546161 = array_index_545928 == array_index_537364 ? add_546160 : sel_546157;
  assign add_546164 = sel_546161 + 8'h01;
  assign sel_546165 = array_index_545928 == array_index_537370 ? add_546164 : sel_546161;
  assign add_546168 = sel_546165 + 8'h01;
  assign sel_546169 = array_index_545928 == array_index_537376 ? add_546168 : sel_546165;
  assign add_546172 = sel_546169 + 8'h01;
  assign sel_546173 = array_index_545928 == array_index_537382 ? add_546172 : sel_546169;
  assign add_546176 = sel_546173 + 8'h01;
  assign sel_546177 = array_index_545928 == array_index_537388 ? add_546176 : sel_546173;
  assign add_546180 = sel_546177 + 8'h01;
  assign sel_546181 = array_index_545928 == array_index_537394 ? add_546180 : sel_546177;
  assign add_546184 = sel_546181 + 8'h01;
  assign sel_546185 = array_index_545928 == array_index_537400 ? add_546184 : sel_546181;
  assign add_546188 = sel_546185 + 8'h01;
  assign sel_546189 = array_index_545928 == array_index_537406 ? add_546188 : sel_546185;
  assign add_546192 = sel_546189 + 8'h01;
  assign sel_546193 = array_index_545928 == array_index_537412 ? add_546192 : sel_546189;
  assign add_546196 = sel_546193 + 8'h01;
  assign sel_546197 = array_index_545928 == array_index_537418 ? add_546196 : sel_546193;
  assign add_546200 = sel_546197 + 8'h01;
  assign sel_546201 = array_index_545928 == array_index_537424 ? add_546200 : sel_546197;
  assign add_546204 = sel_546201 + 8'h01;
  assign sel_546205 = array_index_545928 == array_index_537430 ? add_546204 : sel_546201;
  assign add_546208 = sel_546205 + 8'h01;
  assign sel_546209 = array_index_545928 == array_index_537436 ? add_546208 : sel_546205;
  assign add_546212 = sel_546209 + 8'h01;
  assign sel_546213 = array_index_545928 == array_index_537442 ? add_546212 : sel_546209;
  assign add_546216 = sel_546213 + 8'h01;
  assign sel_546217 = array_index_545928 == array_index_537448 ? add_546216 : sel_546213;
  assign add_546220 = sel_546217 + 8'h01;
  assign sel_546221 = array_index_545928 == array_index_537454 ? add_546220 : sel_546217;
  assign add_546224 = sel_546221 + 8'h01;
  assign sel_546225 = array_index_545928 == array_index_537460 ? add_546224 : sel_546221;
  assign add_546229 = sel_546225 + 8'h01;
  assign array_index_546230 = set1_unflattened[7'h1e];
  assign sel_546231 = array_index_545928 == array_index_537466 ? add_546229 : sel_546225;
  assign add_546234 = sel_546231 + 8'h01;
  assign sel_546235 = array_index_546230 == array_index_537012 ? add_546234 : sel_546231;
  assign add_546238 = sel_546235 + 8'h01;
  assign sel_546239 = array_index_546230 == array_index_537016 ? add_546238 : sel_546235;
  assign add_546242 = sel_546239 + 8'h01;
  assign sel_546243 = array_index_546230 == array_index_537024 ? add_546242 : sel_546239;
  assign add_546246 = sel_546243 + 8'h01;
  assign sel_546247 = array_index_546230 == array_index_537032 ? add_546246 : sel_546243;
  assign add_546250 = sel_546247 + 8'h01;
  assign sel_546251 = array_index_546230 == array_index_537040 ? add_546250 : sel_546247;
  assign add_546254 = sel_546251 + 8'h01;
  assign sel_546255 = array_index_546230 == array_index_537048 ? add_546254 : sel_546251;
  assign add_546258 = sel_546255 + 8'h01;
  assign sel_546259 = array_index_546230 == array_index_537056 ? add_546258 : sel_546255;
  assign add_546262 = sel_546259 + 8'h01;
  assign sel_546263 = array_index_546230 == array_index_537064 ? add_546262 : sel_546259;
  assign add_546266 = sel_546263 + 8'h01;
  assign sel_546267 = array_index_546230 == array_index_537070 ? add_546266 : sel_546263;
  assign add_546270 = sel_546267 + 8'h01;
  assign sel_546271 = array_index_546230 == array_index_537076 ? add_546270 : sel_546267;
  assign add_546274 = sel_546271 + 8'h01;
  assign sel_546275 = array_index_546230 == array_index_537082 ? add_546274 : sel_546271;
  assign add_546278 = sel_546275 + 8'h01;
  assign sel_546279 = array_index_546230 == array_index_537088 ? add_546278 : sel_546275;
  assign add_546282 = sel_546279 + 8'h01;
  assign sel_546283 = array_index_546230 == array_index_537094 ? add_546282 : sel_546279;
  assign add_546286 = sel_546283 + 8'h01;
  assign sel_546287 = array_index_546230 == array_index_537100 ? add_546286 : sel_546283;
  assign add_546290 = sel_546287 + 8'h01;
  assign sel_546291 = array_index_546230 == array_index_537106 ? add_546290 : sel_546287;
  assign add_546294 = sel_546291 + 8'h01;
  assign sel_546295 = array_index_546230 == array_index_537112 ? add_546294 : sel_546291;
  assign add_546298 = sel_546295 + 8'h01;
  assign sel_546299 = array_index_546230 == array_index_537118 ? add_546298 : sel_546295;
  assign add_546302 = sel_546299 + 8'h01;
  assign sel_546303 = array_index_546230 == array_index_537124 ? add_546302 : sel_546299;
  assign add_546306 = sel_546303 + 8'h01;
  assign sel_546307 = array_index_546230 == array_index_537130 ? add_546306 : sel_546303;
  assign add_546310 = sel_546307 + 8'h01;
  assign sel_546311 = array_index_546230 == array_index_537136 ? add_546310 : sel_546307;
  assign add_546314 = sel_546311 + 8'h01;
  assign sel_546315 = array_index_546230 == array_index_537142 ? add_546314 : sel_546311;
  assign add_546318 = sel_546315 + 8'h01;
  assign sel_546319 = array_index_546230 == array_index_537148 ? add_546318 : sel_546315;
  assign add_546322 = sel_546319 + 8'h01;
  assign sel_546323 = array_index_546230 == array_index_537154 ? add_546322 : sel_546319;
  assign add_546326 = sel_546323 + 8'h01;
  assign sel_546327 = array_index_546230 == array_index_537160 ? add_546326 : sel_546323;
  assign add_546330 = sel_546327 + 8'h01;
  assign sel_546331 = array_index_546230 == array_index_537166 ? add_546330 : sel_546327;
  assign add_546334 = sel_546331 + 8'h01;
  assign sel_546335 = array_index_546230 == array_index_537172 ? add_546334 : sel_546331;
  assign add_546338 = sel_546335 + 8'h01;
  assign sel_546339 = array_index_546230 == array_index_537178 ? add_546338 : sel_546335;
  assign add_546342 = sel_546339 + 8'h01;
  assign sel_546343 = array_index_546230 == array_index_537184 ? add_546342 : sel_546339;
  assign add_546346 = sel_546343 + 8'h01;
  assign sel_546347 = array_index_546230 == array_index_537190 ? add_546346 : sel_546343;
  assign add_546350 = sel_546347 + 8'h01;
  assign sel_546351 = array_index_546230 == array_index_537196 ? add_546350 : sel_546347;
  assign add_546354 = sel_546351 + 8'h01;
  assign sel_546355 = array_index_546230 == array_index_537202 ? add_546354 : sel_546351;
  assign add_546358 = sel_546355 + 8'h01;
  assign sel_546359 = array_index_546230 == array_index_537208 ? add_546358 : sel_546355;
  assign add_546362 = sel_546359 + 8'h01;
  assign sel_546363 = array_index_546230 == array_index_537214 ? add_546362 : sel_546359;
  assign add_546366 = sel_546363 + 8'h01;
  assign sel_546367 = array_index_546230 == array_index_537220 ? add_546366 : sel_546363;
  assign add_546370 = sel_546367 + 8'h01;
  assign sel_546371 = array_index_546230 == array_index_537226 ? add_546370 : sel_546367;
  assign add_546374 = sel_546371 + 8'h01;
  assign sel_546375 = array_index_546230 == array_index_537232 ? add_546374 : sel_546371;
  assign add_546378 = sel_546375 + 8'h01;
  assign sel_546379 = array_index_546230 == array_index_537238 ? add_546378 : sel_546375;
  assign add_546382 = sel_546379 + 8'h01;
  assign sel_546383 = array_index_546230 == array_index_537244 ? add_546382 : sel_546379;
  assign add_546386 = sel_546383 + 8'h01;
  assign sel_546387 = array_index_546230 == array_index_537250 ? add_546386 : sel_546383;
  assign add_546390 = sel_546387 + 8'h01;
  assign sel_546391 = array_index_546230 == array_index_537256 ? add_546390 : sel_546387;
  assign add_546394 = sel_546391 + 8'h01;
  assign sel_546395 = array_index_546230 == array_index_537262 ? add_546394 : sel_546391;
  assign add_546398 = sel_546395 + 8'h01;
  assign sel_546399 = array_index_546230 == array_index_537268 ? add_546398 : sel_546395;
  assign add_546402 = sel_546399 + 8'h01;
  assign sel_546403 = array_index_546230 == array_index_537274 ? add_546402 : sel_546399;
  assign add_546406 = sel_546403 + 8'h01;
  assign sel_546407 = array_index_546230 == array_index_537280 ? add_546406 : sel_546403;
  assign add_546410 = sel_546407 + 8'h01;
  assign sel_546411 = array_index_546230 == array_index_537286 ? add_546410 : sel_546407;
  assign add_546414 = sel_546411 + 8'h01;
  assign sel_546415 = array_index_546230 == array_index_537292 ? add_546414 : sel_546411;
  assign add_546418 = sel_546415 + 8'h01;
  assign sel_546419 = array_index_546230 == array_index_537298 ? add_546418 : sel_546415;
  assign add_546422 = sel_546419 + 8'h01;
  assign sel_546423 = array_index_546230 == array_index_537304 ? add_546422 : sel_546419;
  assign add_546426 = sel_546423 + 8'h01;
  assign sel_546427 = array_index_546230 == array_index_537310 ? add_546426 : sel_546423;
  assign add_546430 = sel_546427 + 8'h01;
  assign sel_546431 = array_index_546230 == array_index_537316 ? add_546430 : sel_546427;
  assign add_546434 = sel_546431 + 8'h01;
  assign sel_546435 = array_index_546230 == array_index_537322 ? add_546434 : sel_546431;
  assign add_546438 = sel_546435 + 8'h01;
  assign sel_546439 = array_index_546230 == array_index_537328 ? add_546438 : sel_546435;
  assign add_546442 = sel_546439 + 8'h01;
  assign sel_546443 = array_index_546230 == array_index_537334 ? add_546442 : sel_546439;
  assign add_546446 = sel_546443 + 8'h01;
  assign sel_546447 = array_index_546230 == array_index_537340 ? add_546446 : sel_546443;
  assign add_546450 = sel_546447 + 8'h01;
  assign sel_546451 = array_index_546230 == array_index_537346 ? add_546450 : sel_546447;
  assign add_546454 = sel_546451 + 8'h01;
  assign sel_546455 = array_index_546230 == array_index_537352 ? add_546454 : sel_546451;
  assign add_546458 = sel_546455 + 8'h01;
  assign sel_546459 = array_index_546230 == array_index_537358 ? add_546458 : sel_546455;
  assign add_546462 = sel_546459 + 8'h01;
  assign sel_546463 = array_index_546230 == array_index_537364 ? add_546462 : sel_546459;
  assign add_546466 = sel_546463 + 8'h01;
  assign sel_546467 = array_index_546230 == array_index_537370 ? add_546466 : sel_546463;
  assign add_546470 = sel_546467 + 8'h01;
  assign sel_546471 = array_index_546230 == array_index_537376 ? add_546470 : sel_546467;
  assign add_546474 = sel_546471 + 8'h01;
  assign sel_546475 = array_index_546230 == array_index_537382 ? add_546474 : sel_546471;
  assign add_546478 = sel_546475 + 8'h01;
  assign sel_546479 = array_index_546230 == array_index_537388 ? add_546478 : sel_546475;
  assign add_546482 = sel_546479 + 8'h01;
  assign sel_546483 = array_index_546230 == array_index_537394 ? add_546482 : sel_546479;
  assign add_546486 = sel_546483 + 8'h01;
  assign sel_546487 = array_index_546230 == array_index_537400 ? add_546486 : sel_546483;
  assign add_546490 = sel_546487 + 8'h01;
  assign sel_546491 = array_index_546230 == array_index_537406 ? add_546490 : sel_546487;
  assign add_546494 = sel_546491 + 8'h01;
  assign sel_546495 = array_index_546230 == array_index_537412 ? add_546494 : sel_546491;
  assign add_546498 = sel_546495 + 8'h01;
  assign sel_546499 = array_index_546230 == array_index_537418 ? add_546498 : sel_546495;
  assign add_546502 = sel_546499 + 8'h01;
  assign sel_546503 = array_index_546230 == array_index_537424 ? add_546502 : sel_546499;
  assign add_546506 = sel_546503 + 8'h01;
  assign sel_546507 = array_index_546230 == array_index_537430 ? add_546506 : sel_546503;
  assign add_546510 = sel_546507 + 8'h01;
  assign sel_546511 = array_index_546230 == array_index_537436 ? add_546510 : sel_546507;
  assign add_546514 = sel_546511 + 8'h01;
  assign sel_546515 = array_index_546230 == array_index_537442 ? add_546514 : sel_546511;
  assign add_546518 = sel_546515 + 8'h01;
  assign sel_546519 = array_index_546230 == array_index_537448 ? add_546518 : sel_546515;
  assign add_546522 = sel_546519 + 8'h01;
  assign sel_546523 = array_index_546230 == array_index_537454 ? add_546522 : sel_546519;
  assign add_546526 = sel_546523 + 8'h01;
  assign sel_546527 = array_index_546230 == array_index_537460 ? add_546526 : sel_546523;
  assign add_546531 = sel_546527 + 8'h01;
  assign array_index_546532 = set1_unflattened[7'h1f];
  assign sel_546533 = array_index_546230 == array_index_537466 ? add_546531 : sel_546527;
  assign add_546536 = sel_546533 + 8'h01;
  assign sel_546537 = array_index_546532 == array_index_537012 ? add_546536 : sel_546533;
  assign add_546540 = sel_546537 + 8'h01;
  assign sel_546541 = array_index_546532 == array_index_537016 ? add_546540 : sel_546537;
  assign add_546544 = sel_546541 + 8'h01;
  assign sel_546545 = array_index_546532 == array_index_537024 ? add_546544 : sel_546541;
  assign add_546548 = sel_546545 + 8'h01;
  assign sel_546549 = array_index_546532 == array_index_537032 ? add_546548 : sel_546545;
  assign add_546552 = sel_546549 + 8'h01;
  assign sel_546553 = array_index_546532 == array_index_537040 ? add_546552 : sel_546549;
  assign add_546556 = sel_546553 + 8'h01;
  assign sel_546557 = array_index_546532 == array_index_537048 ? add_546556 : sel_546553;
  assign add_546560 = sel_546557 + 8'h01;
  assign sel_546561 = array_index_546532 == array_index_537056 ? add_546560 : sel_546557;
  assign add_546564 = sel_546561 + 8'h01;
  assign sel_546565 = array_index_546532 == array_index_537064 ? add_546564 : sel_546561;
  assign add_546568 = sel_546565 + 8'h01;
  assign sel_546569 = array_index_546532 == array_index_537070 ? add_546568 : sel_546565;
  assign add_546572 = sel_546569 + 8'h01;
  assign sel_546573 = array_index_546532 == array_index_537076 ? add_546572 : sel_546569;
  assign add_546576 = sel_546573 + 8'h01;
  assign sel_546577 = array_index_546532 == array_index_537082 ? add_546576 : sel_546573;
  assign add_546580 = sel_546577 + 8'h01;
  assign sel_546581 = array_index_546532 == array_index_537088 ? add_546580 : sel_546577;
  assign add_546584 = sel_546581 + 8'h01;
  assign sel_546585 = array_index_546532 == array_index_537094 ? add_546584 : sel_546581;
  assign add_546588 = sel_546585 + 8'h01;
  assign sel_546589 = array_index_546532 == array_index_537100 ? add_546588 : sel_546585;
  assign add_546592 = sel_546589 + 8'h01;
  assign sel_546593 = array_index_546532 == array_index_537106 ? add_546592 : sel_546589;
  assign add_546596 = sel_546593 + 8'h01;
  assign sel_546597 = array_index_546532 == array_index_537112 ? add_546596 : sel_546593;
  assign add_546600 = sel_546597 + 8'h01;
  assign sel_546601 = array_index_546532 == array_index_537118 ? add_546600 : sel_546597;
  assign add_546604 = sel_546601 + 8'h01;
  assign sel_546605 = array_index_546532 == array_index_537124 ? add_546604 : sel_546601;
  assign add_546608 = sel_546605 + 8'h01;
  assign sel_546609 = array_index_546532 == array_index_537130 ? add_546608 : sel_546605;
  assign add_546612 = sel_546609 + 8'h01;
  assign sel_546613 = array_index_546532 == array_index_537136 ? add_546612 : sel_546609;
  assign add_546616 = sel_546613 + 8'h01;
  assign sel_546617 = array_index_546532 == array_index_537142 ? add_546616 : sel_546613;
  assign add_546620 = sel_546617 + 8'h01;
  assign sel_546621 = array_index_546532 == array_index_537148 ? add_546620 : sel_546617;
  assign add_546624 = sel_546621 + 8'h01;
  assign sel_546625 = array_index_546532 == array_index_537154 ? add_546624 : sel_546621;
  assign add_546628 = sel_546625 + 8'h01;
  assign sel_546629 = array_index_546532 == array_index_537160 ? add_546628 : sel_546625;
  assign add_546632 = sel_546629 + 8'h01;
  assign sel_546633 = array_index_546532 == array_index_537166 ? add_546632 : sel_546629;
  assign add_546636 = sel_546633 + 8'h01;
  assign sel_546637 = array_index_546532 == array_index_537172 ? add_546636 : sel_546633;
  assign add_546640 = sel_546637 + 8'h01;
  assign sel_546641 = array_index_546532 == array_index_537178 ? add_546640 : sel_546637;
  assign add_546644 = sel_546641 + 8'h01;
  assign sel_546645 = array_index_546532 == array_index_537184 ? add_546644 : sel_546641;
  assign add_546648 = sel_546645 + 8'h01;
  assign sel_546649 = array_index_546532 == array_index_537190 ? add_546648 : sel_546645;
  assign add_546652 = sel_546649 + 8'h01;
  assign sel_546653 = array_index_546532 == array_index_537196 ? add_546652 : sel_546649;
  assign add_546656 = sel_546653 + 8'h01;
  assign sel_546657 = array_index_546532 == array_index_537202 ? add_546656 : sel_546653;
  assign add_546660 = sel_546657 + 8'h01;
  assign sel_546661 = array_index_546532 == array_index_537208 ? add_546660 : sel_546657;
  assign add_546664 = sel_546661 + 8'h01;
  assign sel_546665 = array_index_546532 == array_index_537214 ? add_546664 : sel_546661;
  assign add_546668 = sel_546665 + 8'h01;
  assign sel_546669 = array_index_546532 == array_index_537220 ? add_546668 : sel_546665;
  assign add_546672 = sel_546669 + 8'h01;
  assign sel_546673 = array_index_546532 == array_index_537226 ? add_546672 : sel_546669;
  assign add_546676 = sel_546673 + 8'h01;
  assign sel_546677 = array_index_546532 == array_index_537232 ? add_546676 : sel_546673;
  assign add_546680 = sel_546677 + 8'h01;
  assign sel_546681 = array_index_546532 == array_index_537238 ? add_546680 : sel_546677;
  assign add_546684 = sel_546681 + 8'h01;
  assign sel_546685 = array_index_546532 == array_index_537244 ? add_546684 : sel_546681;
  assign add_546688 = sel_546685 + 8'h01;
  assign sel_546689 = array_index_546532 == array_index_537250 ? add_546688 : sel_546685;
  assign add_546692 = sel_546689 + 8'h01;
  assign sel_546693 = array_index_546532 == array_index_537256 ? add_546692 : sel_546689;
  assign add_546696 = sel_546693 + 8'h01;
  assign sel_546697 = array_index_546532 == array_index_537262 ? add_546696 : sel_546693;
  assign add_546700 = sel_546697 + 8'h01;
  assign sel_546701 = array_index_546532 == array_index_537268 ? add_546700 : sel_546697;
  assign add_546704 = sel_546701 + 8'h01;
  assign sel_546705 = array_index_546532 == array_index_537274 ? add_546704 : sel_546701;
  assign add_546708 = sel_546705 + 8'h01;
  assign sel_546709 = array_index_546532 == array_index_537280 ? add_546708 : sel_546705;
  assign add_546712 = sel_546709 + 8'h01;
  assign sel_546713 = array_index_546532 == array_index_537286 ? add_546712 : sel_546709;
  assign add_546716 = sel_546713 + 8'h01;
  assign sel_546717 = array_index_546532 == array_index_537292 ? add_546716 : sel_546713;
  assign add_546720 = sel_546717 + 8'h01;
  assign sel_546721 = array_index_546532 == array_index_537298 ? add_546720 : sel_546717;
  assign add_546724 = sel_546721 + 8'h01;
  assign sel_546725 = array_index_546532 == array_index_537304 ? add_546724 : sel_546721;
  assign add_546728 = sel_546725 + 8'h01;
  assign sel_546729 = array_index_546532 == array_index_537310 ? add_546728 : sel_546725;
  assign add_546732 = sel_546729 + 8'h01;
  assign sel_546733 = array_index_546532 == array_index_537316 ? add_546732 : sel_546729;
  assign add_546736 = sel_546733 + 8'h01;
  assign sel_546737 = array_index_546532 == array_index_537322 ? add_546736 : sel_546733;
  assign add_546740 = sel_546737 + 8'h01;
  assign sel_546741 = array_index_546532 == array_index_537328 ? add_546740 : sel_546737;
  assign add_546744 = sel_546741 + 8'h01;
  assign sel_546745 = array_index_546532 == array_index_537334 ? add_546744 : sel_546741;
  assign add_546748 = sel_546745 + 8'h01;
  assign sel_546749 = array_index_546532 == array_index_537340 ? add_546748 : sel_546745;
  assign add_546752 = sel_546749 + 8'h01;
  assign sel_546753 = array_index_546532 == array_index_537346 ? add_546752 : sel_546749;
  assign add_546756 = sel_546753 + 8'h01;
  assign sel_546757 = array_index_546532 == array_index_537352 ? add_546756 : sel_546753;
  assign add_546760 = sel_546757 + 8'h01;
  assign sel_546761 = array_index_546532 == array_index_537358 ? add_546760 : sel_546757;
  assign add_546764 = sel_546761 + 8'h01;
  assign sel_546765 = array_index_546532 == array_index_537364 ? add_546764 : sel_546761;
  assign add_546768 = sel_546765 + 8'h01;
  assign sel_546769 = array_index_546532 == array_index_537370 ? add_546768 : sel_546765;
  assign add_546772 = sel_546769 + 8'h01;
  assign sel_546773 = array_index_546532 == array_index_537376 ? add_546772 : sel_546769;
  assign add_546776 = sel_546773 + 8'h01;
  assign sel_546777 = array_index_546532 == array_index_537382 ? add_546776 : sel_546773;
  assign add_546780 = sel_546777 + 8'h01;
  assign sel_546781 = array_index_546532 == array_index_537388 ? add_546780 : sel_546777;
  assign add_546784 = sel_546781 + 8'h01;
  assign sel_546785 = array_index_546532 == array_index_537394 ? add_546784 : sel_546781;
  assign add_546788 = sel_546785 + 8'h01;
  assign sel_546789 = array_index_546532 == array_index_537400 ? add_546788 : sel_546785;
  assign add_546792 = sel_546789 + 8'h01;
  assign sel_546793 = array_index_546532 == array_index_537406 ? add_546792 : sel_546789;
  assign add_546796 = sel_546793 + 8'h01;
  assign sel_546797 = array_index_546532 == array_index_537412 ? add_546796 : sel_546793;
  assign add_546800 = sel_546797 + 8'h01;
  assign sel_546801 = array_index_546532 == array_index_537418 ? add_546800 : sel_546797;
  assign add_546804 = sel_546801 + 8'h01;
  assign sel_546805 = array_index_546532 == array_index_537424 ? add_546804 : sel_546801;
  assign add_546808 = sel_546805 + 8'h01;
  assign sel_546809 = array_index_546532 == array_index_537430 ? add_546808 : sel_546805;
  assign add_546812 = sel_546809 + 8'h01;
  assign sel_546813 = array_index_546532 == array_index_537436 ? add_546812 : sel_546809;
  assign add_546816 = sel_546813 + 8'h01;
  assign sel_546817 = array_index_546532 == array_index_537442 ? add_546816 : sel_546813;
  assign add_546820 = sel_546817 + 8'h01;
  assign sel_546821 = array_index_546532 == array_index_537448 ? add_546820 : sel_546817;
  assign add_546824 = sel_546821 + 8'h01;
  assign sel_546825 = array_index_546532 == array_index_537454 ? add_546824 : sel_546821;
  assign add_546828 = sel_546825 + 8'h01;
  assign sel_546829 = array_index_546532 == array_index_537460 ? add_546828 : sel_546825;
  assign add_546833 = sel_546829 + 8'h01;
  assign array_index_546834 = set1_unflattened[7'h20];
  assign sel_546835 = array_index_546532 == array_index_537466 ? add_546833 : sel_546829;
  assign add_546838 = sel_546835 + 8'h01;
  assign sel_546839 = array_index_546834 == array_index_537012 ? add_546838 : sel_546835;
  assign add_546842 = sel_546839 + 8'h01;
  assign sel_546843 = array_index_546834 == array_index_537016 ? add_546842 : sel_546839;
  assign add_546846 = sel_546843 + 8'h01;
  assign sel_546847 = array_index_546834 == array_index_537024 ? add_546846 : sel_546843;
  assign add_546850 = sel_546847 + 8'h01;
  assign sel_546851 = array_index_546834 == array_index_537032 ? add_546850 : sel_546847;
  assign add_546854 = sel_546851 + 8'h01;
  assign sel_546855 = array_index_546834 == array_index_537040 ? add_546854 : sel_546851;
  assign add_546858 = sel_546855 + 8'h01;
  assign sel_546859 = array_index_546834 == array_index_537048 ? add_546858 : sel_546855;
  assign add_546862 = sel_546859 + 8'h01;
  assign sel_546863 = array_index_546834 == array_index_537056 ? add_546862 : sel_546859;
  assign add_546866 = sel_546863 + 8'h01;
  assign sel_546867 = array_index_546834 == array_index_537064 ? add_546866 : sel_546863;
  assign add_546870 = sel_546867 + 8'h01;
  assign sel_546871 = array_index_546834 == array_index_537070 ? add_546870 : sel_546867;
  assign add_546874 = sel_546871 + 8'h01;
  assign sel_546875 = array_index_546834 == array_index_537076 ? add_546874 : sel_546871;
  assign add_546878 = sel_546875 + 8'h01;
  assign sel_546879 = array_index_546834 == array_index_537082 ? add_546878 : sel_546875;
  assign add_546882 = sel_546879 + 8'h01;
  assign sel_546883 = array_index_546834 == array_index_537088 ? add_546882 : sel_546879;
  assign add_546886 = sel_546883 + 8'h01;
  assign sel_546887 = array_index_546834 == array_index_537094 ? add_546886 : sel_546883;
  assign add_546890 = sel_546887 + 8'h01;
  assign sel_546891 = array_index_546834 == array_index_537100 ? add_546890 : sel_546887;
  assign add_546894 = sel_546891 + 8'h01;
  assign sel_546895 = array_index_546834 == array_index_537106 ? add_546894 : sel_546891;
  assign add_546898 = sel_546895 + 8'h01;
  assign sel_546899 = array_index_546834 == array_index_537112 ? add_546898 : sel_546895;
  assign add_546902 = sel_546899 + 8'h01;
  assign sel_546903 = array_index_546834 == array_index_537118 ? add_546902 : sel_546899;
  assign add_546906 = sel_546903 + 8'h01;
  assign sel_546907 = array_index_546834 == array_index_537124 ? add_546906 : sel_546903;
  assign add_546910 = sel_546907 + 8'h01;
  assign sel_546911 = array_index_546834 == array_index_537130 ? add_546910 : sel_546907;
  assign add_546914 = sel_546911 + 8'h01;
  assign sel_546915 = array_index_546834 == array_index_537136 ? add_546914 : sel_546911;
  assign add_546918 = sel_546915 + 8'h01;
  assign sel_546919 = array_index_546834 == array_index_537142 ? add_546918 : sel_546915;
  assign add_546922 = sel_546919 + 8'h01;
  assign sel_546923 = array_index_546834 == array_index_537148 ? add_546922 : sel_546919;
  assign add_546926 = sel_546923 + 8'h01;
  assign sel_546927 = array_index_546834 == array_index_537154 ? add_546926 : sel_546923;
  assign add_546930 = sel_546927 + 8'h01;
  assign sel_546931 = array_index_546834 == array_index_537160 ? add_546930 : sel_546927;
  assign add_546934 = sel_546931 + 8'h01;
  assign sel_546935 = array_index_546834 == array_index_537166 ? add_546934 : sel_546931;
  assign add_546938 = sel_546935 + 8'h01;
  assign sel_546939 = array_index_546834 == array_index_537172 ? add_546938 : sel_546935;
  assign add_546942 = sel_546939 + 8'h01;
  assign sel_546943 = array_index_546834 == array_index_537178 ? add_546942 : sel_546939;
  assign add_546946 = sel_546943 + 8'h01;
  assign sel_546947 = array_index_546834 == array_index_537184 ? add_546946 : sel_546943;
  assign add_546950 = sel_546947 + 8'h01;
  assign sel_546951 = array_index_546834 == array_index_537190 ? add_546950 : sel_546947;
  assign add_546954 = sel_546951 + 8'h01;
  assign sel_546955 = array_index_546834 == array_index_537196 ? add_546954 : sel_546951;
  assign add_546958 = sel_546955 + 8'h01;
  assign sel_546959 = array_index_546834 == array_index_537202 ? add_546958 : sel_546955;
  assign add_546962 = sel_546959 + 8'h01;
  assign sel_546963 = array_index_546834 == array_index_537208 ? add_546962 : sel_546959;
  assign add_546966 = sel_546963 + 8'h01;
  assign sel_546967 = array_index_546834 == array_index_537214 ? add_546966 : sel_546963;
  assign add_546970 = sel_546967 + 8'h01;
  assign sel_546971 = array_index_546834 == array_index_537220 ? add_546970 : sel_546967;
  assign add_546974 = sel_546971 + 8'h01;
  assign sel_546975 = array_index_546834 == array_index_537226 ? add_546974 : sel_546971;
  assign add_546978 = sel_546975 + 8'h01;
  assign sel_546979 = array_index_546834 == array_index_537232 ? add_546978 : sel_546975;
  assign add_546982 = sel_546979 + 8'h01;
  assign sel_546983 = array_index_546834 == array_index_537238 ? add_546982 : sel_546979;
  assign add_546986 = sel_546983 + 8'h01;
  assign sel_546987 = array_index_546834 == array_index_537244 ? add_546986 : sel_546983;
  assign add_546990 = sel_546987 + 8'h01;
  assign sel_546991 = array_index_546834 == array_index_537250 ? add_546990 : sel_546987;
  assign add_546994 = sel_546991 + 8'h01;
  assign sel_546995 = array_index_546834 == array_index_537256 ? add_546994 : sel_546991;
  assign add_546998 = sel_546995 + 8'h01;
  assign sel_546999 = array_index_546834 == array_index_537262 ? add_546998 : sel_546995;
  assign add_547002 = sel_546999 + 8'h01;
  assign sel_547003 = array_index_546834 == array_index_537268 ? add_547002 : sel_546999;
  assign add_547006 = sel_547003 + 8'h01;
  assign sel_547007 = array_index_546834 == array_index_537274 ? add_547006 : sel_547003;
  assign add_547010 = sel_547007 + 8'h01;
  assign sel_547011 = array_index_546834 == array_index_537280 ? add_547010 : sel_547007;
  assign add_547014 = sel_547011 + 8'h01;
  assign sel_547015 = array_index_546834 == array_index_537286 ? add_547014 : sel_547011;
  assign add_547018 = sel_547015 + 8'h01;
  assign sel_547019 = array_index_546834 == array_index_537292 ? add_547018 : sel_547015;
  assign add_547022 = sel_547019 + 8'h01;
  assign sel_547023 = array_index_546834 == array_index_537298 ? add_547022 : sel_547019;
  assign add_547026 = sel_547023 + 8'h01;
  assign sel_547027 = array_index_546834 == array_index_537304 ? add_547026 : sel_547023;
  assign add_547030 = sel_547027 + 8'h01;
  assign sel_547031 = array_index_546834 == array_index_537310 ? add_547030 : sel_547027;
  assign add_547034 = sel_547031 + 8'h01;
  assign sel_547035 = array_index_546834 == array_index_537316 ? add_547034 : sel_547031;
  assign add_547038 = sel_547035 + 8'h01;
  assign sel_547039 = array_index_546834 == array_index_537322 ? add_547038 : sel_547035;
  assign add_547042 = sel_547039 + 8'h01;
  assign sel_547043 = array_index_546834 == array_index_537328 ? add_547042 : sel_547039;
  assign add_547046 = sel_547043 + 8'h01;
  assign sel_547047 = array_index_546834 == array_index_537334 ? add_547046 : sel_547043;
  assign add_547050 = sel_547047 + 8'h01;
  assign sel_547051 = array_index_546834 == array_index_537340 ? add_547050 : sel_547047;
  assign add_547054 = sel_547051 + 8'h01;
  assign sel_547055 = array_index_546834 == array_index_537346 ? add_547054 : sel_547051;
  assign add_547058 = sel_547055 + 8'h01;
  assign sel_547059 = array_index_546834 == array_index_537352 ? add_547058 : sel_547055;
  assign add_547062 = sel_547059 + 8'h01;
  assign sel_547063 = array_index_546834 == array_index_537358 ? add_547062 : sel_547059;
  assign add_547066 = sel_547063 + 8'h01;
  assign sel_547067 = array_index_546834 == array_index_537364 ? add_547066 : sel_547063;
  assign add_547070 = sel_547067 + 8'h01;
  assign sel_547071 = array_index_546834 == array_index_537370 ? add_547070 : sel_547067;
  assign add_547074 = sel_547071 + 8'h01;
  assign sel_547075 = array_index_546834 == array_index_537376 ? add_547074 : sel_547071;
  assign add_547078 = sel_547075 + 8'h01;
  assign sel_547079 = array_index_546834 == array_index_537382 ? add_547078 : sel_547075;
  assign add_547082 = sel_547079 + 8'h01;
  assign sel_547083 = array_index_546834 == array_index_537388 ? add_547082 : sel_547079;
  assign add_547086 = sel_547083 + 8'h01;
  assign sel_547087 = array_index_546834 == array_index_537394 ? add_547086 : sel_547083;
  assign add_547090 = sel_547087 + 8'h01;
  assign sel_547091 = array_index_546834 == array_index_537400 ? add_547090 : sel_547087;
  assign add_547094 = sel_547091 + 8'h01;
  assign sel_547095 = array_index_546834 == array_index_537406 ? add_547094 : sel_547091;
  assign add_547098 = sel_547095 + 8'h01;
  assign sel_547099 = array_index_546834 == array_index_537412 ? add_547098 : sel_547095;
  assign add_547102 = sel_547099 + 8'h01;
  assign sel_547103 = array_index_546834 == array_index_537418 ? add_547102 : sel_547099;
  assign add_547106 = sel_547103 + 8'h01;
  assign sel_547107 = array_index_546834 == array_index_537424 ? add_547106 : sel_547103;
  assign add_547110 = sel_547107 + 8'h01;
  assign sel_547111 = array_index_546834 == array_index_537430 ? add_547110 : sel_547107;
  assign add_547114 = sel_547111 + 8'h01;
  assign sel_547115 = array_index_546834 == array_index_537436 ? add_547114 : sel_547111;
  assign add_547118 = sel_547115 + 8'h01;
  assign sel_547119 = array_index_546834 == array_index_537442 ? add_547118 : sel_547115;
  assign add_547122 = sel_547119 + 8'h01;
  assign sel_547123 = array_index_546834 == array_index_537448 ? add_547122 : sel_547119;
  assign add_547126 = sel_547123 + 8'h01;
  assign sel_547127 = array_index_546834 == array_index_537454 ? add_547126 : sel_547123;
  assign add_547130 = sel_547127 + 8'h01;
  assign sel_547131 = array_index_546834 == array_index_537460 ? add_547130 : sel_547127;
  assign add_547135 = sel_547131 + 8'h01;
  assign array_index_547136 = set1_unflattened[7'h21];
  assign sel_547137 = array_index_546834 == array_index_537466 ? add_547135 : sel_547131;
  assign add_547140 = sel_547137 + 8'h01;
  assign sel_547141 = array_index_547136 == array_index_537012 ? add_547140 : sel_547137;
  assign add_547144 = sel_547141 + 8'h01;
  assign sel_547145 = array_index_547136 == array_index_537016 ? add_547144 : sel_547141;
  assign add_547148 = sel_547145 + 8'h01;
  assign sel_547149 = array_index_547136 == array_index_537024 ? add_547148 : sel_547145;
  assign add_547152 = sel_547149 + 8'h01;
  assign sel_547153 = array_index_547136 == array_index_537032 ? add_547152 : sel_547149;
  assign add_547156 = sel_547153 + 8'h01;
  assign sel_547157 = array_index_547136 == array_index_537040 ? add_547156 : sel_547153;
  assign add_547160 = sel_547157 + 8'h01;
  assign sel_547161 = array_index_547136 == array_index_537048 ? add_547160 : sel_547157;
  assign add_547164 = sel_547161 + 8'h01;
  assign sel_547165 = array_index_547136 == array_index_537056 ? add_547164 : sel_547161;
  assign add_547168 = sel_547165 + 8'h01;
  assign sel_547169 = array_index_547136 == array_index_537064 ? add_547168 : sel_547165;
  assign add_547172 = sel_547169 + 8'h01;
  assign sel_547173 = array_index_547136 == array_index_537070 ? add_547172 : sel_547169;
  assign add_547176 = sel_547173 + 8'h01;
  assign sel_547177 = array_index_547136 == array_index_537076 ? add_547176 : sel_547173;
  assign add_547180 = sel_547177 + 8'h01;
  assign sel_547181 = array_index_547136 == array_index_537082 ? add_547180 : sel_547177;
  assign add_547184 = sel_547181 + 8'h01;
  assign sel_547185 = array_index_547136 == array_index_537088 ? add_547184 : sel_547181;
  assign add_547188 = sel_547185 + 8'h01;
  assign sel_547189 = array_index_547136 == array_index_537094 ? add_547188 : sel_547185;
  assign add_547192 = sel_547189 + 8'h01;
  assign sel_547193 = array_index_547136 == array_index_537100 ? add_547192 : sel_547189;
  assign add_547196 = sel_547193 + 8'h01;
  assign sel_547197 = array_index_547136 == array_index_537106 ? add_547196 : sel_547193;
  assign add_547200 = sel_547197 + 8'h01;
  assign sel_547201 = array_index_547136 == array_index_537112 ? add_547200 : sel_547197;
  assign add_547204 = sel_547201 + 8'h01;
  assign sel_547205 = array_index_547136 == array_index_537118 ? add_547204 : sel_547201;
  assign add_547208 = sel_547205 + 8'h01;
  assign sel_547209 = array_index_547136 == array_index_537124 ? add_547208 : sel_547205;
  assign add_547212 = sel_547209 + 8'h01;
  assign sel_547213 = array_index_547136 == array_index_537130 ? add_547212 : sel_547209;
  assign add_547216 = sel_547213 + 8'h01;
  assign sel_547217 = array_index_547136 == array_index_537136 ? add_547216 : sel_547213;
  assign add_547220 = sel_547217 + 8'h01;
  assign sel_547221 = array_index_547136 == array_index_537142 ? add_547220 : sel_547217;
  assign add_547224 = sel_547221 + 8'h01;
  assign sel_547225 = array_index_547136 == array_index_537148 ? add_547224 : sel_547221;
  assign add_547228 = sel_547225 + 8'h01;
  assign sel_547229 = array_index_547136 == array_index_537154 ? add_547228 : sel_547225;
  assign add_547232 = sel_547229 + 8'h01;
  assign sel_547233 = array_index_547136 == array_index_537160 ? add_547232 : sel_547229;
  assign add_547236 = sel_547233 + 8'h01;
  assign sel_547237 = array_index_547136 == array_index_537166 ? add_547236 : sel_547233;
  assign add_547240 = sel_547237 + 8'h01;
  assign sel_547241 = array_index_547136 == array_index_537172 ? add_547240 : sel_547237;
  assign add_547244 = sel_547241 + 8'h01;
  assign sel_547245 = array_index_547136 == array_index_537178 ? add_547244 : sel_547241;
  assign add_547248 = sel_547245 + 8'h01;
  assign sel_547249 = array_index_547136 == array_index_537184 ? add_547248 : sel_547245;
  assign add_547252 = sel_547249 + 8'h01;
  assign sel_547253 = array_index_547136 == array_index_537190 ? add_547252 : sel_547249;
  assign add_547256 = sel_547253 + 8'h01;
  assign sel_547257 = array_index_547136 == array_index_537196 ? add_547256 : sel_547253;
  assign add_547260 = sel_547257 + 8'h01;
  assign sel_547261 = array_index_547136 == array_index_537202 ? add_547260 : sel_547257;
  assign add_547264 = sel_547261 + 8'h01;
  assign sel_547265 = array_index_547136 == array_index_537208 ? add_547264 : sel_547261;
  assign add_547268 = sel_547265 + 8'h01;
  assign sel_547269 = array_index_547136 == array_index_537214 ? add_547268 : sel_547265;
  assign add_547272 = sel_547269 + 8'h01;
  assign sel_547273 = array_index_547136 == array_index_537220 ? add_547272 : sel_547269;
  assign add_547276 = sel_547273 + 8'h01;
  assign sel_547277 = array_index_547136 == array_index_537226 ? add_547276 : sel_547273;
  assign add_547280 = sel_547277 + 8'h01;
  assign sel_547281 = array_index_547136 == array_index_537232 ? add_547280 : sel_547277;
  assign add_547284 = sel_547281 + 8'h01;
  assign sel_547285 = array_index_547136 == array_index_537238 ? add_547284 : sel_547281;
  assign add_547288 = sel_547285 + 8'h01;
  assign sel_547289 = array_index_547136 == array_index_537244 ? add_547288 : sel_547285;
  assign add_547292 = sel_547289 + 8'h01;
  assign sel_547293 = array_index_547136 == array_index_537250 ? add_547292 : sel_547289;
  assign add_547296 = sel_547293 + 8'h01;
  assign sel_547297 = array_index_547136 == array_index_537256 ? add_547296 : sel_547293;
  assign add_547300 = sel_547297 + 8'h01;
  assign sel_547301 = array_index_547136 == array_index_537262 ? add_547300 : sel_547297;
  assign add_547304 = sel_547301 + 8'h01;
  assign sel_547305 = array_index_547136 == array_index_537268 ? add_547304 : sel_547301;
  assign add_547308 = sel_547305 + 8'h01;
  assign sel_547309 = array_index_547136 == array_index_537274 ? add_547308 : sel_547305;
  assign add_547312 = sel_547309 + 8'h01;
  assign sel_547313 = array_index_547136 == array_index_537280 ? add_547312 : sel_547309;
  assign add_547316 = sel_547313 + 8'h01;
  assign sel_547317 = array_index_547136 == array_index_537286 ? add_547316 : sel_547313;
  assign add_547320 = sel_547317 + 8'h01;
  assign sel_547321 = array_index_547136 == array_index_537292 ? add_547320 : sel_547317;
  assign add_547324 = sel_547321 + 8'h01;
  assign sel_547325 = array_index_547136 == array_index_537298 ? add_547324 : sel_547321;
  assign add_547328 = sel_547325 + 8'h01;
  assign sel_547329 = array_index_547136 == array_index_537304 ? add_547328 : sel_547325;
  assign add_547332 = sel_547329 + 8'h01;
  assign sel_547333 = array_index_547136 == array_index_537310 ? add_547332 : sel_547329;
  assign add_547336 = sel_547333 + 8'h01;
  assign sel_547337 = array_index_547136 == array_index_537316 ? add_547336 : sel_547333;
  assign add_547340 = sel_547337 + 8'h01;
  assign sel_547341 = array_index_547136 == array_index_537322 ? add_547340 : sel_547337;
  assign add_547344 = sel_547341 + 8'h01;
  assign sel_547345 = array_index_547136 == array_index_537328 ? add_547344 : sel_547341;
  assign add_547348 = sel_547345 + 8'h01;
  assign sel_547349 = array_index_547136 == array_index_537334 ? add_547348 : sel_547345;
  assign add_547352 = sel_547349 + 8'h01;
  assign sel_547353 = array_index_547136 == array_index_537340 ? add_547352 : sel_547349;
  assign add_547356 = sel_547353 + 8'h01;
  assign sel_547357 = array_index_547136 == array_index_537346 ? add_547356 : sel_547353;
  assign add_547360 = sel_547357 + 8'h01;
  assign sel_547361 = array_index_547136 == array_index_537352 ? add_547360 : sel_547357;
  assign add_547364 = sel_547361 + 8'h01;
  assign sel_547365 = array_index_547136 == array_index_537358 ? add_547364 : sel_547361;
  assign add_547368 = sel_547365 + 8'h01;
  assign sel_547369 = array_index_547136 == array_index_537364 ? add_547368 : sel_547365;
  assign add_547372 = sel_547369 + 8'h01;
  assign sel_547373 = array_index_547136 == array_index_537370 ? add_547372 : sel_547369;
  assign add_547376 = sel_547373 + 8'h01;
  assign sel_547377 = array_index_547136 == array_index_537376 ? add_547376 : sel_547373;
  assign add_547380 = sel_547377 + 8'h01;
  assign sel_547381 = array_index_547136 == array_index_537382 ? add_547380 : sel_547377;
  assign add_547384 = sel_547381 + 8'h01;
  assign sel_547385 = array_index_547136 == array_index_537388 ? add_547384 : sel_547381;
  assign add_547388 = sel_547385 + 8'h01;
  assign sel_547389 = array_index_547136 == array_index_537394 ? add_547388 : sel_547385;
  assign add_547392 = sel_547389 + 8'h01;
  assign sel_547393 = array_index_547136 == array_index_537400 ? add_547392 : sel_547389;
  assign add_547396 = sel_547393 + 8'h01;
  assign sel_547397 = array_index_547136 == array_index_537406 ? add_547396 : sel_547393;
  assign add_547400 = sel_547397 + 8'h01;
  assign sel_547401 = array_index_547136 == array_index_537412 ? add_547400 : sel_547397;
  assign add_547404 = sel_547401 + 8'h01;
  assign sel_547405 = array_index_547136 == array_index_537418 ? add_547404 : sel_547401;
  assign add_547408 = sel_547405 + 8'h01;
  assign sel_547409 = array_index_547136 == array_index_537424 ? add_547408 : sel_547405;
  assign add_547412 = sel_547409 + 8'h01;
  assign sel_547413 = array_index_547136 == array_index_537430 ? add_547412 : sel_547409;
  assign add_547416 = sel_547413 + 8'h01;
  assign sel_547417 = array_index_547136 == array_index_537436 ? add_547416 : sel_547413;
  assign add_547420 = sel_547417 + 8'h01;
  assign sel_547421 = array_index_547136 == array_index_537442 ? add_547420 : sel_547417;
  assign add_547424 = sel_547421 + 8'h01;
  assign sel_547425 = array_index_547136 == array_index_537448 ? add_547424 : sel_547421;
  assign add_547428 = sel_547425 + 8'h01;
  assign sel_547429 = array_index_547136 == array_index_537454 ? add_547428 : sel_547425;
  assign add_547432 = sel_547429 + 8'h01;
  assign sel_547433 = array_index_547136 == array_index_537460 ? add_547432 : sel_547429;
  assign add_547437 = sel_547433 + 8'h01;
  assign array_index_547438 = set1_unflattened[7'h22];
  assign sel_547439 = array_index_547136 == array_index_537466 ? add_547437 : sel_547433;
  assign add_547442 = sel_547439 + 8'h01;
  assign sel_547443 = array_index_547438 == array_index_537012 ? add_547442 : sel_547439;
  assign add_547446 = sel_547443 + 8'h01;
  assign sel_547447 = array_index_547438 == array_index_537016 ? add_547446 : sel_547443;
  assign add_547450 = sel_547447 + 8'h01;
  assign sel_547451 = array_index_547438 == array_index_537024 ? add_547450 : sel_547447;
  assign add_547454 = sel_547451 + 8'h01;
  assign sel_547455 = array_index_547438 == array_index_537032 ? add_547454 : sel_547451;
  assign add_547458 = sel_547455 + 8'h01;
  assign sel_547459 = array_index_547438 == array_index_537040 ? add_547458 : sel_547455;
  assign add_547462 = sel_547459 + 8'h01;
  assign sel_547463 = array_index_547438 == array_index_537048 ? add_547462 : sel_547459;
  assign add_547466 = sel_547463 + 8'h01;
  assign sel_547467 = array_index_547438 == array_index_537056 ? add_547466 : sel_547463;
  assign add_547470 = sel_547467 + 8'h01;
  assign sel_547471 = array_index_547438 == array_index_537064 ? add_547470 : sel_547467;
  assign add_547474 = sel_547471 + 8'h01;
  assign sel_547475 = array_index_547438 == array_index_537070 ? add_547474 : sel_547471;
  assign add_547478 = sel_547475 + 8'h01;
  assign sel_547479 = array_index_547438 == array_index_537076 ? add_547478 : sel_547475;
  assign add_547482 = sel_547479 + 8'h01;
  assign sel_547483 = array_index_547438 == array_index_537082 ? add_547482 : sel_547479;
  assign add_547486 = sel_547483 + 8'h01;
  assign sel_547487 = array_index_547438 == array_index_537088 ? add_547486 : sel_547483;
  assign add_547490 = sel_547487 + 8'h01;
  assign sel_547491 = array_index_547438 == array_index_537094 ? add_547490 : sel_547487;
  assign add_547494 = sel_547491 + 8'h01;
  assign sel_547495 = array_index_547438 == array_index_537100 ? add_547494 : sel_547491;
  assign add_547498 = sel_547495 + 8'h01;
  assign sel_547499 = array_index_547438 == array_index_537106 ? add_547498 : sel_547495;
  assign add_547502 = sel_547499 + 8'h01;
  assign sel_547503 = array_index_547438 == array_index_537112 ? add_547502 : sel_547499;
  assign add_547506 = sel_547503 + 8'h01;
  assign sel_547507 = array_index_547438 == array_index_537118 ? add_547506 : sel_547503;
  assign add_547510 = sel_547507 + 8'h01;
  assign sel_547511 = array_index_547438 == array_index_537124 ? add_547510 : sel_547507;
  assign add_547514 = sel_547511 + 8'h01;
  assign sel_547515 = array_index_547438 == array_index_537130 ? add_547514 : sel_547511;
  assign add_547518 = sel_547515 + 8'h01;
  assign sel_547519 = array_index_547438 == array_index_537136 ? add_547518 : sel_547515;
  assign add_547522 = sel_547519 + 8'h01;
  assign sel_547523 = array_index_547438 == array_index_537142 ? add_547522 : sel_547519;
  assign add_547526 = sel_547523 + 8'h01;
  assign sel_547527 = array_index_547438 == array_index_537148 ? add_547526 : sel_547523;
  assign add_547530 = sel_547527 + 8'h01;
  assign sel_547531 = array_index_547438 == array_index_537154 ? add_547530 : sel_547527;
  assign add_547534 = sel_547531 + 8'h01;
  assign sel_547535 = array_index_547438 == array_index_537160 ? add_547534 : sel_547531;
  assign add_547538 = sel_547535 + 8'h01;
  assign sel_547539 = array_index_547438 == array_index_537166 ? add_547538 : sel_547535;
  assign add_547542 = sel_547539 + 8'h01;
  assign sel_547543 = array_index_547438 == array_index_537172 ? add_547542 : sel_547539;
  assign add_547546 = sel_547543 + 8'h01;
  assign sel_547547 = array_index_547438 == array_index_537178 ? add_547546 : sel_547543;
  assign add_547550 = sel_547547 + 8'h01;
  assign sel_547551 = array_index_547438 == array_index_537184 ? add_547550 : sel_547547;
  assign add_547554 = sel_547551 + 8'h01;
  assign sel_547555 = array_index_547438 == array_index_537190 ? add_547554 : sel_547551;
  assign add_547558 = sel_547555 + 8'h01;
  assign sel_547559 = array_index_547438 == array_index_537196 ? add_547558 : sel_547555;
  assign add_547562 = sel_547559 + 8'h01;
  assign sel_547563 = array_index_547438 == array_index_537202 ? add_547562 : sel_547559;
  assign add_547566 = sel_547563 + 8'h01;
  assign sel_547567 = array_index_547438 == array_index_537208 ? add_547566 : sel_547563;
  assign add_547570 = sel_547567 + 8'h01;
  assign sel_547571 = array_index_547438 == array_index_537214 ? add_547570 : sel_547567;
  assign add_547574 = sel_547571 + 8'h01;
  assign sel_547575 = array_index_547438 == array_index_537220 ? add_547574 : sel_547571;
  assign add_547578 = sel_547575 + 8'h01;
  assign sel_547579 = array_index_547438 == array_index_537226 ? add_547578 : sel_547575;
  assign add_547582 = sel_547579 + 8'h01;
  assign sel_547583 = array_index_547438 == array_index_537232 ? add_547582 : sel_547579;
  assign add_547586 = sel_547583 + 8'h01;
  assign sel_547587 = array_index_547438 == array_index_537238 ? add_547586 : sel_547583;
  assign add_547590 = sel_547587 + 8'h01;
  assign sel_547591 = array_index_547438 == array_index_537244 ? add_547590 : sel_547587;
  assign add_547594 = sel_547591 + 8'h01;
  assign sel_547595 = array_index_547438 == array_index_537250 ? add_547594 : sel_547591;
  assign add_547598 = sel_547595 + 8'h01;
  assign sel_547599 = array_index_547438 == array_index_537256 ? add_547598 : sel_547595;
  assign add_547602 = sel_547599 + 8'h01;
  assign sel_547603 = array_index_547438 == array_index_537262 ? add_547602 : sel_547599;
  assign add_547606 = sel_547603 + 8'h01;
  assign sel_547607 = array_index_547438 == array_index_537268 ? add_547606 : sel_547603;
  assign add_547610 = sel_547607 + 8'h01;
  assign sel_547611 = array_index_547438 == array_index_537274 ? add_547610 : sel_547607;
  assign add_547614 = sel_547611 + 8'h01;
  assign sel_547615 = array_index_547438 == array_index_537280 ? add_547614 : sel_547611;
  assign add_547618 = sel_547615 + 8'h01;
  assign sel_547619 = array_index_547438 == array_index_537286 ? add_547618 : sel_547615;
  assign add_547622 = sel_547619 + 8'h01;
  assign sel_547623 = array_index_547438 == array_index_537292 ? add_547622 : sel_547619;
  assign add_547626 = sel_547623 + 8'h01;
  assign sel_547627 = array_index_547438 == array_index_537298 ? add_547626 : sel_547623;
  assign add_547630 = sel_547627 + 8'h01;
  assign sel_547631 = array_index_547438 == array_index_537304 ? add_547630 : sel_547627;
  assign add_547634 = sel_547631 + 8'h01;
  assign sel_547635 = array_index_547438 == array_index_537310 ? add_547634 : sel_547631;
  assign add_547638 = sel_547635 + 8'h01;
  assign sel_547639 = array_index_547438 == array_index_537316 ? add_547638 : sel_547635;
  assign add_547642 = sel_547639 + 8'h01;
  assign sel_547643 = array_index_547438 == array_index_537322 ? add_547642 : sel_547639;
  assign add_547646 = sel_547643 + 8'h01;
  assign sel_547647 = array_index_547438 == array_index_537328 ? add_547646 : sel_547643;
  assign add_547650 = sel_547647 + 8'h01;
  assign sel_547651 = array_index_547438 == array_index_537334 ? add_547650 : sel_547647;
  assign add_547654 = sel_547651 + 8'h01;
  assign sel_547655 = array_index_547438 == array_index_537340 ? add_547654 : sel_547651;
  assign add_547658 = sel_547655 + 8'h01;
  assign sel_547659 = array_index_547438 == array_index_537346 ? add_547658 : sel_547655;
  assign add_547662 = sel_547659 + 8'h01;
  assign sel_547663 = array_index_547438 == array_index_537352 ? add_547662 : sel_547659;
  assign add_547666 = sel_547663 + 8'h01;
  assign sel_547667 = array_index_547438 == array_index_537358 ? add_547666 : sel_547663;
  assign add_547670 = sel_547667 + 8'h01;
  assign sel_547671 = array_index_547438 == array_index_537364 ? add_547670 : sel_547667;
  assign add_547674 = sel_547671 + 8'h01;
  assign sel_547675 = array_index_547438 == array_index_537370 ? add_547674 : sel_547671;
  assign add_547678 = sel_547675 + 8'h01;
  assign sel_547679 = array_index_547438 == array_index_537376 ? add_547678 : sel_547675;
  assign add_547682 = sel_547679 + 8'h01;
  assign sel_547683 = array_index_547438 == array_index_537382 ? add_547682 : sel_547679;
  assign add_547686 = sel_547683 + 8'h01;
  assign sel_547687 = array_index_547438 == array_index_537388 ? add_547686 : sel_547683;
  assign add_547690 = sel_547687 + 8'h01;
  assign sel_547691 = array_index_547438 == array_index_537394 ? add_547690 : sel_547687;
  assign add_547694 = sel_547691 + 8'h01;
  assign sel_547695 = array_index_547438 == array_index_537400 ? add_547694 : sel_547691;
  assign add_547698 = sel_547695 + 8'h01;
  assign sel_547699 = array_index_547438 == array_index_537406 ? add_547698 : sel_547695;
  assign add_547702 = sel_547699 + 8'h01;
  assign sel_547703 = array_index_547438 == array_index_537412 ? add_547702 : sel_547699;
  assign add_547706 = sel_547703 + 8'h01;
  assign sel_547707 = array_index_547438 == array_index_537418 ? add_547706 : sel_547703;
  assign add_547710 = sel_547707 + 8'h01;
  assign sel_547711 = array_index_547438 == array_index_537424 ? add_547710 : sel_547707;
  assign add_547714 = sel_547711 + 8'h01;
  assign sel_547715 = array_index_547438 == array_index_537430 ? add_547714 : sel_547711;
  assign add_547718 = sel_547715 + 8'h01;
  assign sel_547719 = array_index_547438 == array_index_537436 ? add_547718 : sel_547715;
  assign add_547722 = sel_547719 + 8'h01;
  assign sel_547723 = array_index_547438 == array_index_537442 ? add_547722 : sel_547719;
  assign add_547726 = sel_547723 + 8'h01;
  assign sel_547727 = array_index_547438 == array_index_537448 ? add_547726 : sel_547723;
  assign add_547730 = sel_547727 + 8'h01;
  assign sel_547731 = array_index_547438 == array_index_537454 ? add_547730 : sel_547727;
  assign add_547734 = sel_547731 + 8'h01;
  assign sel_547735 = array_index_547438 == array_index_537460 ? add_547734 : sel_547731;
  assign add_547739 = sel_547735 + 8'h01;
  assign array_index_547740 = set1_unflattened[7'h23];
  assign sel_547741 = array_index_547438 == array_index_537466 ? add_547739 : sel_547735;
  assign add_547744 = sel_547741 + 8'h01;
  assign sel_547745 = array_index_547740 == array_index_537012 ? add_547744 : sel_547741;
  assign add_547748 = sel_547745 + 8'h01;
  assign sel_547749 = array_index_547740 == array_index_537016 ? add_547748 : sel_547745;
  assign add_547752 = sel_547749 + 8'h01;
  assign sel_547753 = array_index_547740 == array_index_537024 ? add_547752 : sel_547749;
  assign add_547756 = sel_547753 + 8'h01;
  assign sel_547757 = array_index_547740 == array_index_537032 ? add_547756 : sel_547753;
  assign add_547760 = sel_547757 + 8'h01;
  assign sel_547761 = array_index_547740 == array_index_537040 ? add_547760 : sel_547757;
  assign add_547764 = sel_547761 + 8'h01;
  assign sel_547765 = array_index_547740 == array_index_537048 ? add_547764 : sel_547761;
  assign add_547768 = sel_547765 + 8'h01;
  assign sel_547769 = array_index_547740 == array_index_537056 ? add_547768 : sel_547765;
  assign add_547772 = sel_547769 + 8'h01;
  assign sel_547773 = array_index_547740 == array_index_537064 ? add_547772 : sel_547769;
  assign add_547776 = sel_547773 + 8'h01;
  assign sel_547777 = array_index_547740 == array_index_537070 ? add_547776 : sel_547773;
  assign add_547780 = sel_547777 + 8'h01;
  assign sel_547781 = array_index_547740 == array_index_537076 ? add_547780 : sel_547777;
  assign add_547784 = sel_547781 + 8'h01;
  assign sel_547785 = array_index_547740 == array_index_537082 ? add_547784 : sel_547781;
  assign add_547788 = sel_547785 + 8'h01;
  assign sel_547789 = array_index_547740 == array_index_537088 ? add_547788 : sel_547785;
  assign add_547792 = sel_547789 + 8'h01;
  assign sel_547793 = array_index_547740 == array_index_537094 ? add_547792 : sel_547789;
  assign add_547796 = sel_547793 + 8'h01;
  assign sel_547797 = array_index_547740 == array_index_537100 ? add_547796 : sel_547793;
  assign add_547800 = sel_547797 + 8'h01;
  assign sel_547801 = array_index_547740 == array_index_537106 ? add_547800 : sel_547797;
  assign add_547804 = sel_547801 + 8'h01;
  assign sel_547805 = array_index_547740 == array_index_537112 ? add_547804 : sel_547801;
  assign add_547808 = sel_547805 + 8'h01;
  assign sel_547809 = array_index_547740 == array_index_537118 ? add_547808 : sel_547805;
  assign add_547812 = sel_547809 + 8'h01;
  assign sel_547813 = array_index_547740 == array_index_537124 ? add_547812 : sel_547809;
  assign add_547816 = sel_547813 + 8'h01;
  assign sel_547817 = array_index_547740 == array_index_537130 ? add_547816 : sel_547813;
  assign add_547820 = sel_547817 + 8'h01;
  assign sel_547821 = array_index_547740 == array_index_537136 ? add_547820 : sel_547817;
  assign add_547824 = sel_547821 + 8'h01;
  assign sel_547825 = array_index_547740 == array_index_537142 ? add_547824 : sel_547821;
  assign add_547828 = sel_547825 + 8'h01;
  assign sel_547829 = array_index_547740 == array_index_537148 ? add_547828 : sel_547825;
  assign add_547832 = sel_547829 + 8'h01;
  assign sel_547833 = array_index_547740 == array_index_537154 ? add_547832 : sel_547829;
  assign add_547836 = sel_547833 + 8'h01;
  assign sel_547837 = array_index_547740 == array_index_537160 ? add_547836 : sel_547833;
  assign add_547840 = sel_547837 + 8'h01;
  assign sel_547841 = array_index_547740 == array_index_537166 ? add_547840 : sel_547837;
  assign add_547844 = sel_547841 + 8'h01;
  assign sel_547845 = array_index_547740 == array_index_537172 ? add_547844 : sel_547841;
  assign add_547848 = sel_547845 + 8'h01;
  assign sel_547849 = array_index_547740 == array_index_537178 ? add_547848 : sel_547845;
  assign add_547852 = sel_547849 + 8'h01;
  assign sel_547853 = array_index_547740 == array_index_537184 ? add_547852 : sel_547849;
  assign add_547856 = sel_547853 + 8'h01;
  assign sel_547857 = array_index_547740 == array_index_537190 ? add_547856 : sel_547853;
  assign add_547860 = sel_547857 + 8'h01;
  assign sel_547861 = array_index_547740 == array_index_537196 ? add_547860 : sel_547857;
  assign add_547864 = sel_547861 + 8'h01;
  assign sel_547865 = array_index_547740 == array_index_537202 ? add_547864 : sel_547861;
  assign add_547868 = sel_547865 + 8'h01;
  assign sel_547869 = array_index_547740 == array_index_537208 ? add_547868 : sel_547865;
  assign add_547872 = sel_547869 + 8'h01;
  assign sel_547873 = array_index_547740 == array_index_537214 ? add_547872 : sel_547869;
  assign add_547876 = sel_547873 + 8'h01;
  assign sel_547877 = array_index_547740 == array_index_537220 ? add_547876 : sel_547873;
  assign add_547880 = sel_547877 + 8'h01;
  assign sel_547881 = array_index_547740 == array_index_537226 ? add_547880 : sel_547877;
  assign add_547884 = sel_547881 + 8'h01;
  assign sel_547885 = array_index_547740 == array_index_537232 ? add_547884 : sel_547881;
  assign add_547888 = sel_547885 + 8'h01;
  assign sel_547889 = array_index_547740 == array_index_537238 ? add_547888 : sel_547885;
  assign add_547892 = sel_547889 + 8'h01;
  assign sel_547893 = array_index_547740 == array_index_537244 ? add_547892 : sel_547889;
  assign add_547896 = sel_547893 + 8'h01;
  assign sel_547897 = array_index_547740 == array_index_537250 ? add_547896 : sel_547893;
  assign add_547900 = sel_547897 + 8'h01;
  assign sel_547901 = array_index_547740 == array_index_537256 ? add_547900 : sel_547897;
  assign add_547904 = sel_547901 + 8'h01;
  assign sel_547905 = array_index_547740 == array_index_537262 ? add_547904 : sel_547901;
  assign add_547908 = sel_547905 + 8'h01;
  assign sel_547909 = array_index_547740 == array_index_537268 ? add_547908 : sel_547905;
  assign add_547912 = sel_547909 + 8'h01;
  assign sel_547913 = array_index_547740 == array_index_537274 ? add_547912 : sel_547909;
  assign add_547916 = sel_547913 + 8'h01;
  assign sel_547917 = array_index_547740 == array_index_537280 ? add_547916 : sel_547913;
  assign add_547920 = sel_547917 + 8'h01;
  assign sel_547921 = array_index_547740 == array_index_537286 ? add_547920 : sel_547917;
  assign add_547924 = sel_547921 + 8'h01;
  assign sel_547925 = array_index_547740 == array_index_537292 ? add_547924 : sel_547921;
  assign add_547928 = sel_547925 + 8'h01;
  assign sel_547929 = array_index_547740 == array_index_537298 ? add_547928 : sel_547925;
  assign add_547932 = sel_547929 + 8'h01;
  assign sel_547933 = array_index_547740 == array_index_537304 ? add_547932 : sel_547929;
  assign add_547936 = sel_547933 + 8'h01;
  assign sel_547937 = array_index_547740 == array_index_537310 ? add_547936 : sel_547933;
  assign add_547940 = sel_547937 + 8'h01;
  assign sel_547941 = array_index_547740 == array_index_537316 ? add_547940 : sel_547937;
  assign add_547944 = sel_547941 + 8'h01;
  assign sel_547945 = array_index_547740 == array_index_537322 ? add_547944 : sel_547941;
  assign add_547948 = sel_547945 + 8'h01;
  assign sel_547949 = array_index_547740 == array_index_537328 ? add_547948 : sel_547945;
  assign add_547952 = sel_547949 + 8'h01;
  assign sel_547953 = array_index_547740 == array_index_537334 ? add_547952 : sel_547949;
  assign add_547956 = sel_547953 + 8'h01;
  assign sel_547957 = array_index_547740 == array_index_537340 ? add_547956 : sel_547953;
  assign add_547960 = sel_547957 + 8'h01;
  assign sel_547961 = array_index_547740 == array_index_537346 ? add_547960 : sel_547957;
  assign add_547964 = sel_547961 + 8'h01;
  assign sel_547965 = array_index_547740 == array_index_537352 ? add_547964 : sel_547961;
  assign add_547968 = sel_547965 + 8'h01;
  assign sel_547969 = array_index_547740 == array_index_537358 ? add_547968 : sel_547965;
  assign add_547972 = sel_547969 + 8'h01;
  assign sel_547973 = array_index_547740 == array_index_537364 ? add_547972 : sel_547969;
  assign add_547976 = sel_547973 + 8'h01;
  assign sel_547977 = array_index_547740 == array_index_537370 ? add_547976 : sel_547973;
  assign add_547980 = sel_547977 + 8'h01;
  assign sel_547981 = array_index_547740 == array_index_537376 ? add_547980 : sel_547977;
  assign add_547984 = sel_547981 + 8'h01;
  assign sel_547985 = array_index_547740 == array_index_537382 ? add_547984 : sel_547981;
  assign add_547988 = sel_547985 + 8'h01;
  assign sel_547989 = array_index_547740 == array_index_537388 ? add_547988 : sel_547985;
  assign add_547992 = sel_547989 + 8'h01;
  assign sel_547993 = array_index_547740 == array_index_537394 ? add_547992 : sel_547989;
  assign add_547996 = sel_547993 + 8'h01;
  assign sel_547997 = array_index_547740 == array_index_537400 ? add_547996 : sel_547993;
  assign add_548000 = sel_547997 + 8'h01;
  assign sel_548001 = array_index_547740 == array_index_537406 ? add_548000 : sel_547997;
  assign add_548004 = sel_548001 + 8'h01;
  assign sel_548005 = array_index_547740 == array_index_537412 ? add_548004 : sel_548001;
  assign add_548008 = sel_548005 + 8'h01;
  assign sel_548009 = array_index_547740 == array_index_537418 ? add_548008 : sel_548005;
  assign add_548012 = sel_548009 + 8'h01;
  assign sel_548013 = array_index_547740 == array_index_537424 ? add_548012 : sel_548009;
  assign add_548016 = sel_548013 + 8'h01;
  assign sel_548017 = array_index_547740 == array_index_537430 ? add_548016 : sel_548013;
  assign add_548020 = sel_548017 + 8'h01;
  assign sel_548021 = array_index_547740 == array_index_537436 ? add_548020 : sel_548017;
  assign add_548024 = sel_548021 + 8'h01;
  assign sel_548025 = array_index_547740 == array_index_537442 ? add_548024 : sel_548021;
  assign add_548028 = sel_548025 + 8'h01;
  assign sel_548029 = array_index_547740 == array_index_537448 ? add_548028 : sel_548025;
  assign add_548032 = sel_548029 + 8'h01;
  assign sel_548033 = array_index_547740 == array_index_537454 ? add_548032 : sel_548029;
  assign add_548036 = sel_548033 + 8'h01;
  assign sel_548037 = array_index_547740 == array_index_537460 ? add_548036 : sel_548033;
  assign add_548041 = sel_548037 + 8'h01;
  assign array_index_548042 = set1_unflattened[7'h24];
  assign sel_548043 = array_index_547740 == array_index_537466 ? add_548041 : sel_548037;
  assign add_548046 = sel_548043 + 8'h01;
  assign sel_548047 = array_index_548042 == array_index_537012 ? add_548046 : sel_548043;
  assign add_548050 = sel_548047 + 8'h01;
  assign sel_548051 = array_index_548042 == array_index_537016 ? add_548050 : sel_548047;
  assign add_548054 = sel_548051 + 8'h01;
  assign sel_548055 = array_index_548042 == array_index_537024 ? add_548054 : sel_548051;
  assign add_548058 = sel_548055 + 8'h01;
  assign sel_548059 = array_index_548042 == array_index_537032 ? add_548058 : sel_548055;
  assign add_548062 = sel_548059 + 8'h01;
  assign sel_548063 = array_index_548042 == array_index_537040 ? add_548062 : sel_548059;
  assign add_548066 = sel_548063 + 8'h01;
  assign sel_548067 = array_index_548042 == array_index_537048 ? add_548066 : sel_548063;
  assign add_548070 = sel_548067 + 8'h01;
  assign sel_548071 = array_index_548042 == array_index_537056 ? add_548070 : sel_548067;
  assign add_548074 = sel_548071 + 8'h01;
  assign sel_548075 = array_index_548042 == array_index_537064 ? add_548074 : sel_548071;
  assign add_548078 = sel_548075 + 8'h01;
  assign sel_548079 = array_index_548042 == array_index_537070 ? add_548078 : sel_548075;
  assign add_548082 = sel_548079 + 8'h01;
  assign sel_548083 = array_index_548042 == array_index_537076 ? add_548082 : sel_548079;
  assign add_548086 = sel_548083 + 8'h01;
  assign sel_548087 = array_index_548042 == array_index_537082 ? add_548086 : sel_548083;
  assign add_548090 = sel_548087 + 8'h01;
  assign sel_548091 = array_index_548042 == array_index_537088 ? add_548090 : sel_548087;
  assign add_548094 = sel_548091 + 8'h01;
  assign sel_548095 = array_index_548042 == array_index_537094 ? add_548094 : sel_548091;
  assign add_548098 = sel_548095 + 8'h01;
  assign sel_548099 = array_index_548042 == array_index_537100 ? add_548098 : sel_548095;
  assign add_548102 = sel_548099 + 8'h01;
  assign sel_548103 = array_index_548042 == array_index_537106 ? add_548102 : sel_548099;
  assign add_548106 = sel_548103 + 8'h01;
  assign sel_548107 = array_index_548042 == array_index_537112 ? add_548106 : sel_548103;
  assign add_548110 = sel_548107 + 8'h01;
  assign sel_548111 = array_index_548042 == array_index_537118 ? add_548110 : sel_548107;
  assign add_548114 = sel_548111 + 8'h01;
  assign sel_548115 = array_index_548042 == array_index_537124 ? add_548114 : sel_548111;
  assign add_548118 = sel_548115 + 8'h01;
  assign sel_548119 = array_index_548042 == array_index_537130 ? add_548118 : sel_548115;
  assign add_548122 = sel_548119 + 8'h01;
  assign sel_548123 = array_index_548042 == array_index_537136 ? add_548122 : sel_548119;
  assign add_548126 = sel_548123 + 8'h01;
  assign sel_548127 = array_index_548042 == array_index_537142 ? add_548126 : sel_548123;
  assign add_548130 = sel_548127 + 8'h01;
  assign sel_548131 = array_index_548042 == array_index_537148 ? add_548130 : sel_548127;
  assign add_548134 = sel_548131 + 8'h01;
  assign sel_548135 = array_index_548042 == array_index_537154 ? add_548134 : sel_548131;
  assign add_548138 = sel_548135 + 8'h01;
  assign sel_548139 = array_index_548042 == array_index_537160 ? add_548138 : sel_548135;
  assign add_548142 = sel_548139 + 8'h01;
  assign sel_548143 = array_index_548042 == array_index_537166 ? add_548142 : sel_548139;
  assign add_548146 = sel_548143 + 8'h01;
  assign sel_548147 = array_index_548042 == array_index_537172 ? add_548146 : sel_548143;
  assign add_548150 = sel_548147 + 8'h01;
  assign sel_548151 = array_index_548042 == array_index_537178 ? add_548150 : sel_548147;
  assign add_548154 = sel_548151 + 8'h01;
  assign sel_548155 = array_index_548042 == array_index_537184 ? add_548154 : sel_548151;
  assign add_548158 = sel_548155 + 8'h01;
  assign sel_548159 = array_index_548042 == array_index_537190 ? add_548158 : sel_548155;
  assign add_548162 = sel_548159 + 8'h01;
  assign sel_548163 = array_index_548042 == array_index_537196 ? add_548162 : sel_548159;
  assign add_548166 = sel_548163 + 8'h01;
  assign sel_548167 = array_index_548042 == array_index_537202 ? add_548166 : sel_548163;
  assign add_548170 = sel_548167 + 8'h01;
  assign sel_548171 = array_index_548042 == array_index_537208 ? add_548170 : sel_548167;
  assign add_548174 = sel_548171 + 8'h01;
  assign sel_548175 = array_index_548042 == array_index_537214 ? add_548174 : sel_548171;
  assign add_548178 = sel_548175 + 8'h01;
  assign sel_548179 = array_index_548042 == array_index_537220 ? add_548178 : sel_548175;
  assign add_548182 = sel_548179 + 8'h01;
  assign sel_548183 = array_index_548042 == array_index_537226 ? add_548182 : sel_548179;
  assign add_548186 = sel_548183 + 8'h01;
  assign sel_548187 = array_index_548042 == array_index_537232 ? add_548186 : sel_548183;
  assign add_548190 = sel_548187 + 8'h01;
  assign sel_548191 = array_index_548042 == array_index_537238 ? add_548190 : sel_548187;
  assign add_548194 = sel_548191 + 8'h01;
  assign sel_548195 = array_index_548042 == array_index_537244 ? add_548194 : sel_548191;
  assign add_548198 = sel_548195 + 8'h01;
  assign sel_548199 = array_index_548042 == array_index_537250 ? add_548198 : sel_548195;
  assign add_548202 = sel_548199 + 8'h01;
  assign sel_548203 = array_index_548042 == array_index_537256 ? add_548202 : sel_548199;
  assign add_548206 = sel_548203 + 8'h01;
  assign sel_548207 = array_index_548042 == array_index_537262 ? add_548206 : sel_548203;
  assign add_548210 = sel_548207 + 8'h01;
  assign sel_548211 = array_index_548042 == array_index_537268 ? add_548210 : sel_548207;
  assign add_548214 = sel_548211 + 8'h01;
  assign sel_548215 = array_index_548042 == array_index_537274 ? add_548214 : sel_548211;
  assign add_548218 = sel_548215 + 8'h01;
  assign sel_548219 = array_index_548042 == array_index_537280 ? add_548218 : sel_548215;
  assign add_548222 = sel_548219 + 8'h01;
  assign sel_548223 = array_index_548042 == array_index_537286 ? add_548222 : sel_548219;
  assign add_548226 = sel_548223 + 8'h01;
  assign sel_548227 = array_index_548042 == array_index_537292 ? add_548226 : sel_548223;
  assign add_548230 = sel_548227 + 8'h01;
  assign sel_548231 = array_index_548042 == array_index_537298 ? add_548230 : sel_548227;
  assign add_548234 = sel_548231 + 8'h01;
  assign sel_548235 = array_index_548042 == array_index_537304 ? add_548234 : sel_548231;
  assign add_548238 = sel_548235 + 8'h01;
  assign sel_548239 = array_index_548042 == array_index_537310 ? add_548238 : sel_548235;
  assign add_548242 = sel_548239 + 8'h01;
  assign sel_548243 = array_index_548042 == array_index_537316 ? add_548242 : sel_548239;
  assign add_548246 = sel_548243 + 8'h01;
  assign sel_548247 = array_index_548042 == array_index_537322 ? add_548246 : sel_548243;
  assign add_548250 = sel_548247 + 8'h01;
  assign sel_548251 = array_index_548042 == array_index_537328 ? add_548250 : sel_548247;
  assign add_548254 = sel_548251 + 8'h01;
  assign sel_548255 = array_index_548042 == array_index_537334 ? add_548254 : sel_548251;
  assign add_548258 = sel_548255 + 8'h01;
  assign sel_548259 = array_index_548042 == array_index_537340 ? add_548258 : sel_548255;
  assign add_548262 = sel_548259 + 8'h01;
  assign sel_548263 = array_index_548042 == array_index_537346 ? add_548262 : sel_548259;
  assign add_548266 = sel_548263 + 8'h01;
  assign sel_548267 = array_index_548042 == array_index_537352 ? add_548266 : sel_548263;
  assign add_548270 = sel_548267 + 8'h01;
  assign sel_548271 = array_index_548042 == array_index_537358 ? add_548270 : sel_548267;
  assign add_548274 = sel_548271 + 8'h01;
  assign sel_548275 = array_index_548042 == array_index_537364 ? add_548274 : sel_548271;
  assign add_548278 = sel_548275 + 8'h01;
  assign sel_548279 = array_index_548042 == array_index_537370 ? add_548278 : sel_548275;
  assign add_548282 = sel_548279 + 8'h01;
  assign sel_548283 = array_index_548042 == array_index_537376 ? add_548282 : sel_548279;
  assign add_548286 = sel_548283 + 8'h01;
  assign sel_548287 = array_index_548042 == array_index_537382 ? add_548286 : sel_548283;
  assign add_548290 = sel_548287 + 8'h01;
  assign sel_548291 = array_index_548042 == array_index_537388 ? add_548290 : sel_548287;
  assign add_548294 = sel_548291 + 8'h01;
  assign sel_548295 = array_index_548042 == array_index_537394 ? add_548294 : sel_548291;
  assign add_548298 = sel_548295 + 8'h01;
  assign sel_548299 = array_index_548042 == array_index_537400 ? add_548298 : sel_548295;
  assign add_548302 = sel_548299 + 8'h01;
  assign sel_548303 = array_index_548042 == array_index_537406 ? add_548302 : sel_548299;
  assign add_548306 = sel_548303 + 8'h01;
  assign sel_548307 = array_index_548042 == array_index_537412 ? add_548306 : sel_548303;
  assign add_548310 = sel_548307 + 8'h01;
  assign sel_548311 = array_index_548042 == array_index_537418 ? add_548310 : sel_548307;
  assign add_548314 = sel_548311 + 8'h01;
  assign sel_548315 = array_index_548042 == array_index_537424 ? add_548314 : sel_548311;
  assign add_548318 = sel_548315 + 8'h01;
  assign sel_548319 = array_index_548042 == array_index_537430 ? add_548318 : sel_548315;
  assign add_548322 = sel_548319 + 8'h01;
  assign sel_548323 = array_index_548042 == array_index_537436 ? add_548322 : sel_548319;
  assign add_548326 = sel_548323 + 8'h01;
  assign sel_548327 = array_index_548042 == array_index_537442 ? add_548326 : sel_548323;
  assign add_548330 = sel_548327 + 8'h01;
  assign sel_548331 = array_index_548042 == array_index_537448 ? add_548330 : sel_548327;
  assign add_548334 = sel_548331 + 8'h01;
  assign sel_548335 = array_index_548042 == array_index_537454 ? add_548334 : sel_548331;
  assign add_548338 = sel_548335 + 8'h01;
  assign sel_548339 = array_index_548042 == array_index_537460 ? add_548338 : sel_548335;
  assign add_548343 = sel_548339 + 8'h01;
  assign array_index_548344 = set1_unflattened[7'h25];
  assign sel_548345 = array_index_548042 == array_index_537466 ? add_548343 : sel_548339;
  assign add_548348 = sel_548345 + 8'h01;
  assign sel_548349 = array_index_548344 == array_index_537012 ? add_548348 : sel_548345;
  assign add_548352 = sel_548349 + 8'h01;
  assign sel_548353 = array_index_548344 == array_index_537016 ? add_548352 : sel_548349;
  assign add_548356 = sel_548353 + 8'h01;
  assign sel_548357 = array_index_548344 == array_index_537024 ? add_548356 : sel_548353;
  assign add_548360 = sel_548357 + 8'h01;
  assign sel_548361 = array_index_548344 == array_index_537032 ? add_548360 : sel_548357;
  assign add_548364 = sel_548361 + 8'h01;
  assign sel_548365 = array_index_548344 == array_index_537040 ? add_548364 : sel_548361;
  assign add_548368 = sel_548365 + 8'h01;
  assign sel_548369 = array_index_548344 == array_index_537048 ? add_548368 : sel_548365;
  assign add_548372 = sel_548369 + 8'h01;
  assign sel_548373 = array_index_548344 == array_index_537056 ? add_548372 : sel_548369;
  assign add_548376 = sel_548373 + 8'h01;
  assign sel_548377 = array_index_548344 == array_index_537064 ? add_548376 : sel_548373;
  assign add_548380 = sel_548377 + 8'h01;
  assign sel_548381 = array_index_548344 == array_index_537070 ? add_548380 : sel_548377;
  assign add_548384 = sel_548381 + 8'h01;
  assign sel_548385 = array_index_548344 == array_index_537076 ? add_548384 : sel_548381;
  assign add_548388 = sel_548385 + 8'h01;
  assign sel_548389 = array_index_548344 == array_index_537082 ? add_548388 : sel_548385;
  assign add_548392 = sel_548389 + 8'h01;
  assign sel_548393 = array_index_548344 == array_index_537088 ? add_548392 : sel_548389;
  assign add_548396 = sel_548393 + 8'h01;
  assign sel_548397 = array_index_548344 == array_index_537094 ? add_548396 : sel_548393;
  assign add_548400 = sel_548397 + 8'h01;
  assign sel_548401 = array_index_548344 == array_index_537100 ? add_548400 : sel_548397;
  assign add_548404 = sel_548401 + 8'h01;
  assign sel_548405 = array_index_548344 == array_index_537106 ? add_548404 : sel_548401;
  assign add_548408 = sel_548405 + 8'h01;
  assign sel_548409 = array_index_548344 == array_index_537112 ? add_548408 : sel_548405;
  assign add_548412 = sel_548409 + 8'h01;
  assign sel_548413 = array_index_548344 == array_index_537118 ? add_548412 : sel_548409;
  assign add_548416 = sel_548413 + 8'h01;
  assign sel_548417 = array_index_548344 == array_index_537124 ? add_548416 : sel_548413;
  assign add_548420 = sel_548417 + 8'h01;
  assign sel_548421 = array_index_548344 == array_index_537130 ? add_548420 : sel_548417;
  assign add_548424 = sel_548421 + 8'h01;
  assign sel_548425 = array_index_548344 == array_index_537136 ? add_548424 : sel_548421;
  assign add_548428 = sel_548425 + 8'h01;
  assign sel_548429 = array_index_548344 == array_index_537142 ? add_548428 : sel_548425;
  assign add_548432 = sel_548429 + 8'h01;
  assign sel_548433 = array_index_548344 == array_index_537148 ? add_548432 : sel_548429;
  assign add_548436 = sel_548433 + 8'h01;
  assign sel_548437 = array_index_548344 == array_index_537154 ? add_548436 : sel_548433;
  assign add_548440 = sel_548437 + 8'h01;
  assign sel_548441 = array_index_548344 == array_index_537160 ? add_548440 : sel_548437;
  assign add_548444 = sel_548441 + 8'h01;
  assign sel_548445 = array_index_548344 == array_index_537166 ? add_548444 : sel_548441;
  assign add_548448 = sel_548445 + 8'h01;
  assign sel_548449 = array_index_548344 == array_index_537172 ? add_548448 : sel_548445;
  assign add_548452 = sel_548449 + 8'h01;
  assign sel_548453 = array_index_548344 == array_index_537178 ? add_548452 : sel_548449;
  assign add_548456 = sel_548453 + 8'h01;
  assign sel_548457 = array_index_548344 == array_index_537184 ? add_548456 : sel_548453;
  assign add_548460 = sel_548457 + 8'h01;
  assign sel_548461 = array_index_548344 == array_index_537190 ? add_548460 : sel_548457;
  assign add_548464 = sel_548461 + 8'h01;
  assign sel_548465 = array_index_548344 == array_index_537196 ? add_548464 : sel_548461;
  assign add_548468 = sel_548465 + 8'h01;
  assign sel_548469 = array_index_548344 == array_index_537202 ? add_548468 : sel_548465;
  assign add_548472 = sel_548469 + 8'h01;
  assign sel_548473 = array_index_548344 == array_index_537208 ? add_548472 : sel_548469;
  assign add_548476 = sel_548473 + 8'h01;
  assign sel_548477 = array_index_548344 == array_index_537214 ? add_548476 : sel_548473;
  assign add_548480 = sel_548477 + 8'h01;
  assign sel_548481 = array_index_548344 == array_index_537220 ? add_548480 : sel_548477;
  assign add_548484 = sel_548481 + 8'h01;
  assign sel_548485 = array_index_548344 == array_index_537226 ? add_548484 : sel_548481;
  assign add_548488 = sel_548485 + 8'h01;
  assign sel_548489 = array_index_548344 == array_index_537232 ? add_548488 : sel_548485;
  assign add_548492 = sel_548489 + 8'h01;
  assign sel_548493 = array_index_548344 == array_index_537238 ? add_548492 : sel_548489;
  assign add_548496 = sel_548493 + 8'h01;
  assign sel_548497 = array_index_548344 == array_index_537244 ? add_548496 : sel_548493;
  assign add_548500 = sel_548497 + 8'h01;
  assign sel_548501 = array_index_548344 == array_index_537250 ? add_548500 : sel_548497;
  assign add_548504 = sel_548501 + 8'h01;
  assign sel_548505 = array_index_548344 == array_index_537256 ? add_548504 : sel_548501;
  assign add_548508 = sel_548505 + 8'h01;
  assign sel_548509 = array_index_548344 == array_index_537262 ? add_548508 : sel_548505;
  assign add_548512 = sel_548509 + 8'h01;
  assign sel_548513 = array_index_548344 == array_index_537268 ? add_548512 : sel_548509;
  assign add_548516 = sel_548513 + 8'h01;
  assign sel_548517 = array_index_548344 == array_index_537274 ? add_548516 : sel_548513;
  assign add_548520 = sel_548517 + 8'h01;
  assign sel_548521 = array_index_548344 == array_index_537280 ? add_548520 : sel_548517;
  assign add_548524 = sel_548521 + 8'h01;
  assign sel_548525 = array_index_548344 == array_index_537286 ? add_548524 : sel_548521;
  assign add_548528 = sel_548525 + 8'h01;
  assign sel_548529 = array_index_548344 == array_index_537292 ? add_548528 : sel_548525;
  assign add_548532 = sel_548529 + 8'h01;
  assign sel_548533 = array_index_548344 == array_index_537298 ? add_548532 : sel_548529;
  assign add_548536 = sel_548533 + 8'h01;
  assign sel_548537 = array_index_548344 == array_index_537304 ? add_548536 : sel_548533;
  assign add_548540 = sel_548537 + 8'h01;
  assign sel_548541 = array_index_548344 == array_index_537310 ? add_548540 : sel_548537;
  assign add_548544 = sel_548541 + 8'h01;
  assign sel_548545 = array_index_548344 == array_index_537316 ? add_548544 : sel_548541;
  assign add_548548 = sel_548545 + 8'h01;
  assign sel_548549 = array_index_548344 == array_index_537322 ? add_548548 : sel_548545;
  assign add_548552 = sel_548549 + 8'h01;
  assign sel_548553 = array_index_548344 == array_index_537328 ? add_548552 : sel_548549;
  assign add_548556 = sel_548553 + 8'h01;
  assign sel_548557 = array_index_548344 == array_index_537334 ? add_548556 : sel_548553;
  assign add_548560 = sel_548557 + 8'h01;
  assign sel_548561 = array_index_548344 == array_index_537340 ? add_548560 : sel_548557;
  assign add_548564 = sel_548561 + 8'h01;
  assign sel_548565 = array_index_548344 == array_index_537346 ? add_548564 : sel_548561;
  assign add_548568 = sel_548565 + 8'h01;
  assign sel_548569 = array_index_548344 == array_index_537352 ? add_548568 : sel_548565;
  assign add_548572 = sel_548569 + 8'h01;
  assign sel_548573 = array_index_548344 == array_index_537358 ? add_548572 : sel_548569;
  assign add_548576 = sel_548573 + 8'h01;
  assign sel_548577 = array_index_548344 == array_index_537364 ? add_548576 : sel_548573;
  assign add_548580 = sel_548577 + 8'h01;
  assign sel_548581 = array_index_548344 == array_index_537370 ? add_548580 : sel_548577;
  assign add_548584 = sel_548581 + 8'h01;
  assign sel_548585 = array_index_548344 == array_index_537376 ? add_548584 : sel_548581;
  assign add_548588 = sel_548585 + 8'h01;
  assign sel_548589 = array_index_548344 == array_index_537382 ? add_548588 : sel_548585;
  assign add_548592 = sel_548589 + 8'h01;
  assign sel_548593 = array_index_548344 == array_index_537388 ? add_548592 : sel_548589;
  assign add_548596 = sel_548593 + 8'h01;
  assign sel_548597 = array_index_548344 == array_index_537394 ? add_548596 : sel_548593;
  assign add_548600 = sel_548597 + 8'h01;
  assign sel_548601 = array_index_548344 == array_index_537400 ? add_548600 : sel_548597;
  assign add_548604 = sel_548601 + 8'h01;
  assign sel_548605 = array_index_548344 == array_index_537406 ? add_548604 : sel_548601;
  assign add_548608 = sel_548605 + 8'h01;
  assign sel_548609 = array_index_548344 == array_index_537412 ? add_548608 : sel_548605;
  assign add_548612 = sel_548609 + 8'h01;
  assign sel_548613 = array_index_548344 == array_index_537418 ? add_548612 : sel_548609;
  assign add_548616 = sel_548613 + 8'h01;
  assign sel_548617 = array_index_548344 == array_index_537424 ? add_548616 : sel_548613;
  assign add_548620 = sel_548617 + 8'h01;
  assign sel_548621 = array_index_548344 == array_index_537430 ? add_548620 : sel_548617;
  assign add_548624 = sel_548621 + 8'h01;
  assign sel_548625 = array_index_548344 == array_index_537436 ? add_548624 : sel_548621;
  assign add_548628 = sel_548625 + 8'h01;
  assign sel_548629 = array_index_548344 == array_index_537442 ? add_548628 : sel_548625;
  assign add_548632 = sel_548629 + 8'h01;
  assign sel_548633 = array_index_548344 == array_index_537448 ? add_548632 : sel_548629;
  assign add_548636 = sel_548633 + 8'h01;
  assign sel_548637 = array_index_548344 == array_index_537454 ? add_548636 : sel_548633;
  assign add_548640 = sel_548637 + 8'h01;
  assign sel_548641 = array_index_548344 == array_index_537460 ? add_548640 : sel_548637;
  assign add_548645 = sel_548641 + 8'h01;
  assign array_index_548646 = set1_unflattened[7'h26];
  assign sel_548647 = array_index_548344 == array_index_537466 ? add_548645 : sel_548641;
  assign add_548650 = sel_548647 + 8'h01;
  assign sel_548651 = array_index_548646 == array_index_537012 ? add_548650 : sel_548647;
  assign add_548654 = sel_548651 + 8'h01;
  assign sel_548655 = array_index_548646 == array_index_537016 ? add_548654 : sel_548651;
  assign add_548658 = sel_548655 + 8'h01;
  assign sel_548659 = array_index_548646 == array_index_537024 ? add_548658 : sel_548655;
  assign add_548662 = sel_548659 + 8'h01;
  assign sel_548663 = array_index_548646 == array_index_537032 ? add_548662 : sel_548659;
  assign add_548666 = sel_548663 + 8'h01;
  assign sel_548667 = array_index_548646 == array_index_537040 ? add_548666 : sel_548663;
  assign add_548670 = sel_548667 + 8'h01;
  assign sel_548671 = array_index_548646 == array_index_537048 ? add_548670 : sel_548667;
  assign add_548674 = sel_548671 + 8'h01;
  assign sel_548675 = array_index_548646 == array_index_537056 ? add_548674 : sel_548671;
  assign add_548678 = sel_548675 + 8'h01;
  assign sel_548679 = array_index_548646 == array_index_537064 ? add_548678 : sel_548675;
  assign add_548682 = sel_548679 + 8'h01;
  assign sel_548683 = array_index_548646 == array_index_537070 ? add_548682 : sel_548679;
  assign add_548686 = sel_548683 + 8'h01;
  assign sel_548687 = array_index_548646 == array_index_537076 ? add_548686 : sel_548683;
  assign add_548690 = sel_548687 + 8'h01;
  assign sel_548691 = array_index_548646 == array_index_537082 ? add_548690 : sel_548687;
  assign add_548694 = sel_548691 + 8'h01;
  assign sel_548695 = array_index_548646 == array_index_537088 ? add_548694 : sel_548691;
  assign add_548698 = sel_548695 + 8'h01;
  assign sel_548699 = array_index_548646 == array_index_537094 ? add_548698 : sel_548695;
  assign add_548702 = sel_548699 + 8'h01;
  assign sel_548703 = array_index_548646 == array_index_537100 ? add_548702 : sel_548699;
  assign add_548706 = sel_548703 + 8'h01;
  assign sel_548707 = array_index_548646 == array_index_537106 ? add_548706 : sel_548703;
  assign add_548710 = sel_548707 + 8'h01;
  assign sel_548711 = array_index_548646 == array_index_537112 ? add_548710 : sel_548707;
  assign add_548714 = sel_548711 + 8'h01;
  assign sel_548715 = array_index_548646 == array_index_537118 ? add_548714 : sel_548711;
  assign add_548718 = sel_548715 + 8'h01;
  assign sel_548719 = array_index_548646 == array_index_537124 ? add_548718 : sel_548715;
  assign add_548722 = sel_548719 + 8'h01;
  assign sel_548723 = array_index_548646 == array_index_537130 ? add_548722 : sel_548719;
  assign add_548726 = sel_548723 + 8'h01;
  assign sel_548727 = array_index_548646 == array_index_537136 ? add_548726 : sel_548723;
  assign add_548730 = sel_548727 + 8'h01;
  assign sel_548731 = array_index_548646 == array_index_537142 ? add_548730 : sel_548727;
  assign add_548734 = sel_548731 + 8'h01;
  assign sel_548735 = array_index_548646 == array_index_537148 ? add_548734 : sel_548731;
  assign add_548738 = sel_548735 + 8'h01;
  assign sel_548739 = array_index_548646 == array_index_537154 ? add_548738 : sel_548735;
  assign add_548742 = sel_548739 + 8'h01;
  assign sel_548743 = array_index_548646 == array_index_537160 ? add_548742 : sel_548739;
  assign add_548746 = sel_548743 + 8'h01;
  assign sel_548747 = array_index_548646 == array_index_537166 ? add_548746 : sel_548743;
  assign add_548750 = sel_548747 + 8'h01;
  assign sel_548751 = array_index_548646 == array_index_537172 ? add_548750 : sel_548747;
  assign add_548754 = sel_548751 + 8'h01;
  assign sel_548755 = array_index_548646 == array_index_537178 ? add_548754 : sel_548751;
  assign add_548758 = sel_548755 + 8'h01;
  assign sel_548759 = array_index_548646 == array_index_537184 ? add_548758 : sel_548755;
  assign add_548762 = sel_548759 + 8'h01;
  assign sel_548763 = array_index_548646 == array_index_537190 ? add_548762 : sel_548759;
  assign add_548766 = sel_548763 + 8'h01;
  assign sel_548767 = array_index_548646 == array_index_537196 ? add_548766 : sel_548763;
  assign add_548770 = sel_548767 + 8'h01;
  assign sel_548771 = array_index_548646 == array_index_537202 ? add_548770 : sel_548767;
  assign add_548774 = sel_548771 + 8'h01;
  assign sel_548775 = array_index_548646 == array_index_537208 ? add_548774 : sel_548771;
  assign add_548778 = sel_548775 + 8'h01;
  assign sel_548779 = array_index_548646 == array_index_537214 ? add_548778 : sel_548775;
  assign add_548782 = sel_548779 + 8'h01;
  assign sel_548783 = array_index_548646 == array_index_537220 ? add_548782 : sel_548779;
  assign add_548786 = sel_548783 + 8'h01;
  assign sel_548787 = array_index_548646 == array_index_537226 ? add_548786 : sel_548783;
  assign add_548790 = sel_548787 + 8'h01;
  assign sel_548791 = array_index_548646 == array_index_537232 ? add_548790 : sel_548787;
  assign add_548794 = sel_548791 + 8'h01;
  assign sel_548795 = array_index_548646 == array_index_537238 ? add_548794 : sel_548791;
  assign add_548798 = sel_548795 + 8'h01;
  assign sel_548799 = array_index_548646 == array_index_537244 ? add_548798 : sel_548795;
  assign add_548802 = sel_548799 + 8'h01;
  assign sel_548803 = array_index_548646 == array_index_537250 ? add_548802 : sel_548799;
  assign add_548806 = sel_548803 + 8'h01;
  assign sel_548807 = array_index_548646 == array_index_537256 ? add_548806 : sel_548803;
  assign add_548810 = sel_548807 + 8'h01;
  assign sel_548811 = array_index_548646 == array_index_537262 ? add_548810 : sel_548807;
  assign add_548814 = sel_548811 + 8'h01;
  assign sel_548815 = array_index_548646 == array_index_537268 ? add_548814 : sel_548811;
  assign add_548818 = sel_548815 + 8'h01;
  assign sel_548819 = array_index_548646 == array_index_537274 ? add_548818 : sel_548815;
  assign add_548822 = sel_548819 + 8'h01;
  assign sel_548823 = array_index_548646 == array_index_537280 ? add_548822 : sel_548819;
  assign add_548826 = sel_548823 + 8'h01;
  assign sel_548827 = array_index_548646 == array_index_537286 ? add_548826 : sel_548823;
  assign add_548830 = sel_548827 + 8'h01;
  assign sel_548831 = array_index_548646 == array_index_537292 ? add_548830 : sel_548827;
  assign add_548834 = sel_548831 + 8'h01;
  assign sel_548835 = array_index_548646 == array_index_537298 ? add_548834 : sel_548831;
  assign add_548838 = sel_548835 + 8'h01;
  assign sel_548839 = array_index_548646 == array_index_537304 ? add_548838 : sel_548835;
  assign add_548842 = sel_548839 + 8'h01;
  assign sel_548843 = array_index_548646 == array_index_537310 ? add_548842 : sel_548839;
  assign add_548846 = sel_548843 + 8'h01;
  assign sel_548847 = array_index_548646 == array_index_537316 ? add_548846 : sel_548843;
  assign add_548850 = sel_548847 + 8'h01;
  assign sel_548851 = array_index_548646 == array_index_537322 ? add_548850 : sel_548847;
  assign add_548854 = sel_548851 + 8'h01;
  assign sel_548855 = array_index_548646 == array_index_537328 ? add_548854 : sel_548851;
  assign add_548858 = sel_548855 + 8'h01;
  assign sel_548859 = array_index_548646 == array_index_537334 ? add_548858 : sel_548855;
  assign add_548862 = sel_548859 + 8'h01;
  assign sel_548863 = array_index_548646 == array_index_537340 ? add_548862 : sel_548859;
  assign add_548866 = sel_548863 + 8'h01;
  assign sel_548867 = array_index_548646 == array_index_537346 ? add_548866 : sel_548863;
  assign add_548870 = sel_548867 + 8'h01;
  assign sel_548871 = array_index_548646 == array_index_537352 ? add_548870 : sel_548867;
  assign add_548874 = sel_548871 + 8'h01;
  assign sel_548875 = array_index_548646 == array_index_537358 ? add_548874 : sel_548871;
  assign add_548878 = sel_548875 + 8'h01;
  assign sel_548879 = array_index_548646 == array_index_537364 ? add_548878 : sel_548875;
  assign add_548882 = sel_548879 + 8'h01;
  assign sel_548883 = array_index_548646 == array_index_537370 ? add_548882 : sel_548879;
  assign add_548886 = sel_548883 + 8'h01;
  assign sel_548887 = array_index_548646 == array_index_537376 ? add_548886 : sel_548883;
  assign add_548890 = sel_548887 + 8'h01;
  assign sel_548891 = array_index_548646 == array_index_537382 ? add_548890 : sel_548887;
  assign add_548894 = sel_548891 + 8'h01;
  assign sel_548895 = array_index_548646 == array_index_537388 ? add_548894 : sel_548891;
  assign add_548898 = sel_548895 + 8'h01;
  assign sel_548899 = array_index_548646 == array_index_537394 ? add_548898 : sel_548895;
  assign add_548902 = sel_548899 + 8'h01;
  assign sel_548903 = array_index_548646 == array_index_537400 ? add_548902 : sel_548899;
  assign add_548906 = sel_548903 + 8'h01;
  assign sel_548907 = array_index_548646 == array_index_537406 ? add_548906 : sel_548903;
  assign add_548910 = sel_548907 + 8'h01;
  assign sel_548911 = array_index_548646 == array_index_537412 ? add_548910 : sel_548907;
  assign add_548914 = sel_548911 + 8'h01;
  assign sel_548915 = array_index_548646 == array_index_537418 ? add_548914 : sel_548911;
  assign add_548918 = sel_548915 + 8'h01;
  assign sel_548919 = array_index_548646 == array_index_537424 ? add_548918 : sel_548915;
  assign add_548922 = sel_548919 + 8'h01;
  assign sel_548923 = array_index_548646 == array_index_537430 ? add_548922 : sel_548919;
  assign add_548926 = sel_548923 + 8'h01;
  assign sel_548927 = array_index_548646 == array_index_537436 ? add_548926 : sel_548923;
  assign add_548930 = sel_548927 + 8'h01;
  assign sel_548931 = array_index_548646 == array_index_537442 ? add_548930 : sel_548927;
  assign add_548934 = sel_548931 + 8'h01;
  assign sel_548935 = array_index_548646 == array_index_537448 ? add_548934 : sel_548931;
  assign add_548938 = sel_548935 + 8'h01;
  assign sel_548939 = array_index_548646 == array_index_537454 ? add_548938 : sel_548935;
  assign add_548942 = sel_548939 + 8'h01;
  assign sel_548943 = array_index_548646 == array_index_537460 ? add_548942 : sel_548939;
  assign add_548947 = sel_548943 + 8'h01;
  assign array_index_548948 = set1_unflattened[7'h27];
  assign sel_548949 = array_index_548646 == array_index_537466 ? add_548947 : sel_548943;
  assign add_548952 = sel_548949 + 8'h01;
  assign sel_548953 = array_index_548948 == array_index_537012 ? add_548952 : sel_548949;
  assign add_548956 = sel_548953 + 8'h01;
  assign sel_548957 = array_index_548948 == array_index_537016 ? add_548956 : sel_548953;
  assign add_548960 = sel_548957 + 8'h01;
  assign sel_548961 = array_index_548948 == array_index_537024 ? add_548960 : sel_548957;
  assign add_548964 = sel_548961 + 8'h01;
  assign sel_548965 = array_index_548948 == array_index_537032 ? add_548964 : sel_548961;
  assign add_548968 = sel_548965 + 8'h01;
  assign sel_548969 = array_index_548948 == array_index_537040 ? add_548968 : sel_548965;
  assign add_548972 = sel_548969 + 8'h01;
  assign sel_548973 = array_index_548948 == array_index_537048 ? add_548972 : sel_548969;
  assign add_548976 = sel_548973 + 8'h01;
  assign sel_548977 = array_index_548948 == array_index_537056 ? add_548976 : sel_548973;
  assign add_548980 = sel_548977 + 8'h01;
  assign sel_548981 = array_index_548948 == array_index_537064 ? add_548980 : sel_548977;
  assign add_548984 = sel_548981 + 8'h01;
  assign sel_548985 = array_index_548948 == array_index_537070 ? add_548984 : sel_548981;
  assign add_548988 = sel_548985 + 8'h01;
  assign sel_548989 = array_index_548948 == array_index_537076 ? add_548988 : sel_548985;
  assign add_548992 = sel_548989 + 8'h01;
  assign sel_548993 = array_index_548948 == array_index_537082 ? add_548992 : sel_548989;
  assign add_548996 = sel_548993 + 8'h01;
  assign sel_548997 = array_index_548948 == array_index_537088 ? add_548996 : sel_548993;
  assign add_549000 = sel_548997 + 8'h01;
  assign sel_549001 = array_index_548948 == array_index_537094 ? add_549000 : sel_548997;
  assign add_549004 = sel_549001 + 8'h01;
  assign sel_549005 = array_index_548948 == array_index_537100 ? add_549004 : sel_549001;
  assign add_549008 = sel_549005 + 8'h01;
  assign sel_549009 = array_index_548948 == array_index_537106 ? add_549008 : sel_549005;
  assign add_549012 = sel_549009 + 8'h01;
  assign sel_549013 = array_index_548948 == array_index_537112 ? add_549012 : sel_549009;
  assign add_549016 = sel_549013 + 8'h01;
  assign sel_549017 = array_index_548948 == array_index_537118 ? add_549016 : sel_549013;
  assign add_549020 = sel_549017 + 8'h01;
  assign sel_549021 = array_index_548948 == array_index_537124 ? add_549020 : sel_549017;
  assign add_549024 = sel_549021 + 8'h01;
  assign sel_549025 = array_index_548948 == array_index_537130 ? add_549024 : sel_549021;
  assign add_549028 = sel_549025 + 8'h01;
  assign sel_549029 = array_index_548948 == array_index_537136 ? add_549028 : sel_549025;
  assign add_549032 = sel_549029 + 8'h01;
  assign sel_549033 = array_index_548948 == array_index_537142 ? add_549032 : sel_549029;
  assign add_549036 = sel_549033 + 8'h01;
  assign sel_549037 = array_index_548948 == array_index_537148 ? add_549036 : sel_549033;
  assign add_549040 = sel_549037 + 8'h01;
  assign sel_549041 = array_index_548948 == array_index_537154 ? add_549040 : sel_549037;
  assign add_549044 = sel_549041 + 8'h01;
  assign sel_549045 = array_index_548948 == array_index_537160 ? add_549044 : sel_549041;
  assign add_549048 = sel_549045 + 8'h01;
  assign sel_549049 = array_index_548948 == array_index_537166 ? add_549048 : sel_549045;
  assign add_549052 = sel_549049 + 8'h01;
  assign sel_549053 = array_index_548948 == array_index_537172 ? add_549052 : sel_549049;
  assign add_549056 = sel_549053 + 8'h01;
  assign sel_549057 = array_index_548948 == array_index_537178 ? add_549056 : sel_549053;
  assign add_549060 = sel_549057 + 8'h01;
  assign sel_549061 = array_index_548948 == array_index_537184 ? add_549060 : sel_549057;
  assign add_549064 = sel_549061 + 8'h01;
  assign sel_549065 = array_index_548948 == array_index_537190 ? add_549064 : sel_549061;
  assign add_549068 = sel_549065 + 8'h01;
  assign sel_549069 = array_index_548948 == array_index_537196 ? add_549068 : sel_549065;
  assign add_549072 = sel_549069 + 8'h01;
  assign sel_549073 = array_index_548948 == array_index_537202 ? add_549072 : sel_549069;
  assign add_549076 = sel_549073 + 8'h01;
  assign sel_549077 = array_index_548948 == array_index_537208 ? add_549076 : sel_549073;
  assign add_549080 = sel_549077 + 8'h01;
  assign sel_549081 = array_index_548948 == array_index_537214 ? add_549080 : sel_549077;
  assign add_549084 = sel_549081 + 8'h01;
  assign sel_549085 = array_index_548948 == array_index_537220 ? add_549084 : sel_549081;
  assign add_549088 = sel_549085 + 8'h01;
  assign sel_549089 = array_index_548948 == array_index_537226 ? add_549088 : sel_549085;
  assign add_549092 = sel_549089 + 8'h01;
  assign sel_549093 = array_index_548948 == array_index_537232 ? add_549092 : sel_549089;
  assign add_549096 = sel_549093 + 8'h01;
  assign sel_549097 = array_index_548948 == array_index_537238 ? add_549096 : sel_549093;
  assign add_549100 = sel_549097 + 8'h01;
  assign sel_549101 = array_index_548948 == array_index_537244 ? add_549100 : sel_549097;
  assign add_549104 = sel_549101 + 8'h01;
  assign sel_549105 = array_index_548948 == array_index_537250 ? add_549104 : sel_549101;
  assign add_549108 = sel_549105 + 8'h01;
  assign sel_549109 = array_index_548948 == array_index_537256 ? add_549108 : sel_549105;
  assign add_549112 = sel_549109 + 8'h01;
  assign sel_549113 = array_index_548948 == array_index_537262 ? add_549112 : sel_549109;
  assign add_549116 = sel_549113 + 8'h01;
  assign sel_549117 = array_index_548948 == array_index_537268 ? add_549116 : sel_549113;
  assign add_549120 = sel_549117 + 8'h01;
  assign sel_549121 = array_index_548948 == array_index_537274 ? add_549120 : sel_549117;
  assign add_549124 = sel_549121 + 8'h01;
  assign sel_549125 = array_index_548948 == array_index_537280 ? add_549124 : sel_549121;
  assign add_549128 = sel_549125 + 8'h01;
  assign sel_549129 = array_index_548948 == array_index_537286 ? add_549128 : sel_549125;
  assign add_549132 = sel_549129 + 8'h01;
  assign sel_549133 = array_index_548948 == array_index_537292 ? add_549132 : sel_549129;
  assign add_549136 = sel_549133 + 8'h01;
  assign sel_549137 = array_index_548948 == array_index_537298 ? add_549136 : sel_549133;
  assign add_549140 = sel_549137 + 8'h01;
  assign sel_549141 = array_index_548948 == array_index_537304 ? add_549140 : sel_549137;
  assign add_549144 = sel_549141 + 8'h01;
  assign sel_549145 = array_index_548948 == array_index_537310 ? add_549144 : sel_549141;
  assign add_549148 = sel_549145 + 8'h01;
  assign sel_549149 = array_index_548948 == array_index_537316 ? add_549148 : sel_549145;
  assign add_549152 = sel_549149 + 8'h01;
  assign sel_549153 = array_index_548948 == array_index_537322 ? add_549152 : sel_549149;
  assign add_549156 = sel_549153 + 8'h01;
  assign sel_549157 = array_index_548948 == array_index_537328 ? add_549156 : sel_549153;
  assign add_549160 = sel_549157 + 8'h01;
  assign sel_549161 = array_index_548948 == array_index_537334 ? add_549160 : sel_549157;
  assign add_549164 = sel_549161 + 8'h01;
  assign sel_549165 = array_index_548948 == array_index_537340 ? add_549164 : sel_549161;
  assign add_549168 = sel_549165 + 8'h01;
  assign sel_549169 = array_index_548948 == array_index_537346 ? add_549168 : sel_549165;
  assign add_549172 = sel_549169 + 8'h01;
  assign sel_549173 = array_index_548948 == array_index_537352 ? add_549172 : sel_549169;
  assign add_549176 = sel_549173 + 8'h01;
  assign sel_549177 = array_index_548948 == array_index_537358 ? add_549176 : sel_549173;
  assign add_549180 = sel_549177 + 8'h01;
  assign sel_549181 = array_index_548948 == array_index_537364 ? add_549180 : sel_549177;
  assign add_549184 = sel_549181 + 8'h01;
  assign sel_549185 = array_index_548948 == array_index_537370 ? add_549184 : sel_549181;
  assign add_549188 = sel_549185 + 8'h01;
  assign sel_549189 = array_index_548948 == array_index_537376 ? add_549188 : sel_549185;
  assign add_549192 = sel_549189 + 8'h01;
  assign sel_549193 = array_index_548948 == array_index_537382 ? add_549192 : sel_549189;
  assign add_549196 = sel_549193 + 8'h01;
  assign sel_549197 = array_index_548948 == array_index_537388 ? add_549196 : sel_549193;
  assign add_549200 = sel_549197 + 8'h01;
  assign sel_549201 = array_index_548948 == array_index_537394 ? add_549200 : sel_549197;
  assign add_549204 = sel_549201 + 8'h01;
  assign sel_549205 = array_index_548948 == array_index_537400 ? add_549204 : sel_549201;
  assign add_549208 = sel_549205 + 8'h01;
  assign sel_549209 = array_index_548948 == array_index_537406 ? add_549208 : sel_549205;
  assign add_549212 = sel_549209 + 8'h01;
  assign sel_549213 = array_index_548948 == array_index_537412 ? add_549212 : sel_549209;
  assign add_549216 = sel_549213 + 8'h01;
  assign sel_549217 = array_index_548948 == array_index_537418 ? add_549216 : sel_549213;
  assign add_549220 = sel_549217 + 8'h01;
  assign sel_549221 = array_index_548948 == array_index_537424 ? add_549220 : sel_549217;
  assign add_549224 = sel_549221 + 8'h01;
  assign sel_549225 = array_index_548948 == array_index_537430 ? add_549224 : sel_549221;
  assign add_549228 = sel_549225 + 8'h01;
  assign sel_549229 = array_index_548948 == array_index_537436 ? add_549228 : sel_549225;
  assign add_549232 = sel_549229 + 8'h01;
  assign sel_549233 = array_index_548948 == array_index_537442 ? add_549232 : sel_549229;
  assign add_549236 = sel_549233 + 8'h01;
  assign sel_549237 = array_index_548948 == array_index_537448 ? add_549236 : sel_549233;
  assign add_549240 = sel_549237 + 8'h01;
  assign sel_549241 = array_index_548948 == array_index_537454 ? add_549240 : sel_549237;
  assign add_549244 = sel_549241 + 8'h01;
  assign sel_549245 = array_index_548948 == array_index_537460 ? add_549244 : sel_549241;
  assign add_549249 = sel_549245 + 8'h01;
  assign array_index_549250 = set1_unflattened[7'h28];
  assign sel_549251 = array_index_548948 == array_index_537466 ? add_549249 : sel_549245;
  assign add_549254 = sel_549251 + 8'h01;
  assign sel_549255 = array_index_549250 == array_index_537012 ? add_549254 : sel_549251;
  assign add_549258 = sel_549255 + 8'h01;
  assign sel_549259 = array_index_549250 == array_index_537016 ? add_549258 : sel_549255;
  assign add_549262 = sel_549259 + 8'h01;
  assign sel_549263 = array_index_549250 == array_index_537024 ? add_549262 : sel_549259;
  assign add_549266 = sel_549263 + 8'h01;
  assign sel_549267 = array_index_549250 == array_index_537032 ? add_549266 : sel_549263;
  assign add_549270 = sel_549267 + 8'h01;
  assign sel_549271 = array_index_549250 == array_index_537040 ? add_549270 : sel_549267;
  assign add_549274 = sel_549271 + 8'h01;
  assign sel_549275 = array_index_549250 == array_index_537048 ? add_549274 : sel_549271;
  assign add_549278 = sel_549275 + 8'h01;
  assign sel_549279 = array_index_549250 == array_index_537056 ? add_549278 : sel_549275;
  assign add_549282 = sel_549279 + 8'h01;
  assign sel_549283 = array_index_549250 == array_index_537064 ? add_549282 : sel_549279;
  assign add_549286 = sel_549283 + 8'h01;
  assign sel_549287 = array_index_549250 == array_index_537070 ? add_549286 : sel_549283;
  assign add_549290 = sel_549287 + 8'h01;
  assign sel_549291 = array_index_549250 == array_index_537076 ? add_549290 : sel_549287;
  assign add_549294 = sel_549291 + 8'h01;
  assign sel_549295 = array_index_549250 == array_index_537082 ? add_549294 : sel_549291;
  assign add_549298 = sel_549295 + 8'h01;
  assign sel_549299 = array_index_549250 == array_index_537088 ? add_549298 : sel_549295;
  assign add_549302 = sel_549299 + 8'h01;
  assign sel_549303 = array_index_549250 == array_index_537094 ? add_549302 : sel_549299;
  assign add_549306 = sel_549303 + 8'h01;
  assign sel_549307 = array_index_549250 == array_index_537100 ? add_549306 : sel_549303;
  assign add_549310 = sel_549307 + 8'h01;
  assign sel_549311 = array_index_549250 == array_index_537106 ? add_549310 : sel_549307;
  assign add_549314 = sel_549311 + 8'h01;
  assign sel_549315 = array_index_549250 == array_index_537112 ? add_549314 : sel_549311;
  assign add_549318 = sel_549315 + 8'h01;
  assign sel_549319 = array_index_549250 == array_index_537118 ? add_549318 : sel_549315;
  assign add_549322 = sel_549319 + 8'h01;
  assign sel_549323 = array_index_549250 == array_index_537124 ? add_549322 : sel_549319;
  assign add_549326 = sel_549323 + 8'h01;
  assign sel_549327 = array_index_549250 == array_index_537130 ? add_549326 : sel_549323;
  assign add_549330 = sel_549327 + 8'h01;
  assign sel_549331 = array_index_549250 == array_index_537136 ? add_549330 : sel_549327;
  assign add_549334 = sel_549331 + 8'h01;
  assign sel_549335 = array_index_549250 == array_index_537142 ? add_549334 : sel_549331;
  assign add_549338 = sel_549335 + 8'h01;
  assign sel_549339 = array_index_549250 == array_index_537148 ? add_549338 : sel_549335;
  assign add_549342 = sel_549339 + 8'h01;
  assign sel_549343 = array_index_549250 == array_index_537154 ? add_549342 : sel_549339;
  assign add_549346 = sel_549343 + 8'h01;
  assign sel_549347 = array_index_549250 == array_index_537160 ? add_549346 : sel_549343;
  assign add_549350 = sel_549347 + 8'h01;
  assign sel_549351 = array_index_549250 == array_index_537166 ? add_549350 : sel_549347;
  assign add_549354 = sel_549351 + 8'h01;
  assign sel_549355 = array_index_549250 == array_index_537172 ? add_549354 : sel_549351;
  assign add_549358 = sel_549355 + 8'h01;
  assign sel_549359 = array_index_549250 == array_index_537178 ? add_549358 : sel_549355;
  assign add_549362 = sel_549359 + 8'h01;
  assign sel_549363 = array_index_549250 == array_index_537184 ? add_549362 : sel_549359;
  assign add_549366 = sel_549363 + 8'h01;
  assign sel_549367 = array_index_549250 == array_index_537190 ? add_549366 : sel_549363;
  assign add_549370 = sel_549367 + 8'h01;
  assign sel_549371 = array_index_549250 == array_index_537196 ? add_549370 : sel_549367;
  assign add_549374 = sel_549371 + 8'h01;
  assign sel_549375 = array_index_549250 == array_index_537202 ? add_549374 : sel_549371;
  assign add_549378 = sel_549375 + 8'h01;
  assign sel_549379 = array_index_549250 == array_index_537208 ? add_549378 : sel_549375;
  assign add_549382 = sel_549379 + 8'h01;
  assign sel_549383 = array_index_549250 == array_index_537214 ? add_549382 : sel_549379;
  assign add_549386 = sel_549383 + 8'h01;
  assign sel_549387 = array_index_549250 == array_index_537220 ? add_549386 : sel_549383;
  assign add_549390 = sel_549387 + 8'h01;
  assign sel_549391 = array_index_549250 == array_index_537226 ? add_549390 : sel_549387;
  assign add_549394 = sel_549391 + 8'h01;
  assign sel_549395 = array_index_549250 == array_index_537232 ? add_549394 : sel_549391;
  assign add_549398 = sel_549395 + 8'h01;
  assign sel_549399 = array_index_549250 == array_index_537238 ? add_549398 : sel_549395;
  assign add_549402 = sel_549399 + 8'h01;
  assign sel_549403 = array_index_549250 == array_index_537244 ? add_549402 : sel_549399;
  assign add_549406 = sel_549403 + 8'h01;
  assign sel_549407 = array_index_549250 == array_index_537250 ? add_549406 : sel_549403;
  assign add_549410 = sel_549407 + 8'h01;
  assign sel_549411 = array_index_549250 == array_index_537256 ? add_549410 : sel_549407;
  assign add_549414 = sel_549411 + 8'h01;
  assign sel_549415 = array_index_549250 == array_index_537262 ? add_549414 : sel_549411;
  assign add_549418 = sel_549415 + 8'h01;
  assign sel_549419 = array_index_549250 == array_index_537268 ? add_549418 : sel_549415;
  assign add_549422 = sel_549419 + 8'h01;
  assign sel_549423 = array_index_549250 == array_index_537274 ? add_549422 : sel_549419;
  assign add_549426 = sel_549423 + 8'h01;
  assign sel_549427 = array_index_549250 == array_index_537280 ? add_549426 : sel_549423;
  assign add_549430 = sel_549427 + 8'h01;
  assign sel_549431 = array_index_549250 == array_index_537286 ? add_549430 : sel_549427;
  assign add_549434 = sel_549431 + 8'h01;
  assign sel_549435 = array_index_549250 == array_index_537292 ? add_549434 : sel_549431;
  assign add_549438 = sel_549435 + 8'h01;
  assign sel_549439 = array_index_549250 == array_index_537298 ? add_549438 : sel_549435;
  assign add_549442 = sel_549439 + 8'h01;
  assign sel_549443 = array_index_549250 == array_index_537304 ? add_549442 : sel_549439;
  assign add_549446 = sel_549443 + 8'h01;
  assign sel_549447 = array_index_549250 == array_index_537310 ? add_549446 : sel_549443;
  assign add_549450 = sel_549447 + 8'h01;
  assign sel_549451 = array_index_549250 == array_index_537316 ? add_549450 : sel_549447;
  assign add_549454 = sel_549451 + 8'h01;
  assign sel_549455 = array_index_549250 == array_index_537322 ? add_549454 : sel_549451;
  assign add_549458 = sel_549455 + 8'h01;
  assign sel_549459 = array_index_549250 == array_index_537328 ? add_549458 : sel_549455;
  assign add_549462 = sel_549459 + 8'h01;
  assign sel_549463 = array_index_549250 == array_index_537334 ? add_549462 : sel_549459;
  assign add_549466 = sel_549463 + 8'h01;
  assign sel_549467 = array_index_549250 == array_index_537340 ? add_549466 : sel_549463;
  assign add_549470 = sel_549467 + 8'h01;
  assign sel_549471 = array_index_549250 == array_index_537346 ? add_549470 : sel_549467;
  assign add_549474 = sel_549471 + 8'h01;
  assign sel_549475 = array_index_549250 == array_index_537352 ? add_549474 : sel_549471;
  assign add_549478 = sel_549475 + 8'h01;
  assign sel_549479 = array_index_549250 == array_index_537358 ? add_549478 : sel_549475;
  assign add_549482 = sel_549479 + 8'h01;
  assign sel_549483 = array_index_549250 == array_index_537364 ? add_549482 : sel_549479;
  assign add_549486 = sel_549483 + 8'h01;
  assign sel_549487 = array_index_549250 == array_index_537370 ? add_549486 : sel_549483;
  assign add_549490 = sel_549487 + 8'h01;
  assign sel_549491 = array_index_549250 == array_index_537376 ? add_549490 : sel_549487;
  assign add_549494 = sel_549491 + 8'h01;
  assign sel_549495 = array_index_549250 == array_index_537382 ? add_549494 : sel_549491;
  assign add_549498 = sel_549495 + 8'h01;
  assign sel_549499 = array_index_549250 == array_index_537388 ? add_549498 : sel_549495;
  assign add_549502 = sel_549499 + 8'h01;
  assign sel_549503 = array_index_549250 == array_index_537394 ? add_549502 : sel_549499;
  assign add_549506 = sel_549503 + 8'h01;
  assign sel_549507 = array_index_549250 == array_index_537400 ? add_549506 : sel_549503;
  assign add_549510 = sel_549507 + 8'h01;
  assign sel_549511 = array_index_549250 == array_index_537406 ? add_549510 : sel_549507;
  assign add_549514 = sel_549511 + 8'h01;
  assign sel_549515 = array_index_549250 == array_index_537412 ? add_549514 : sel_549511;
  assign add_549518 = sel_549515 + 8'h01;
  assign sel_549519 = array_index_549250 == array_index_537418 ? add_549518 : sel_549515;
  assign add_549522 = sel_549519 + 8'h01;
  assign sel_549523 = array_index_549250 == array_index_537424 ? add_549522 : sel_549519;
  assign add_549526 = sel_549523 + 8'h01;
  assign sel_549527 = array_index_549250 == array_index_537430 ? add_549526 : sel_549523;
  assign add_549530 = sel_549527 + 8'h01;
  assign sel_549531 = array_index_549250 == array_index_537436 ? add_549530 : sel_549527;
  assign add_549534 = sel_549531 + 8'h01;
  assign sel_549535 = array_index_549250 == array_index_537442 ? add_549534 : sel_549531;
  assign add_549538 = sel_549535 + 8'h01;
  assign sel_549539 = array_index_549250 == array_index_537448 ? add_549538 : sel_549535;
  assign add_549542 = sel_549539 + 8'h01;
  assign sel_549543 = array_index_549250 == array_index_537454 ? add_549542 : sel_549539;
  assign add_549546 = sel_549543 + 8'h01;
  assign sel_549547 = array_index_549250 == array_index_537460 ? add_549546 : sel_549543;
  assign add_549551 = sel_549547 + 8'h01;
  assign array_index_549552 = set1_unflattened[7'h29];
  assign sel_549553 = array_index_549250 == array_index_537466 ? add_549551 : sel_549547;
  assign add_549556 = sel_549553 + 8'h01;
  assign sel_549557 = array_index_549552 == array_index_537012 ? add_549556 : sel_549553;
  assign add_549560 = sel_549557 + 8'h01;
  assign sel_549561 = array_index_549552 == array_index_537016 ? add_549560 : sel_549557;
  assign add_549564 = sel_549561 + 8'h01;
  assign sel_549565 = array_index_549552 == array_index_537024 ? add_549564 : sel_549561;
  assign add_549568 = sel_549565 + 8'h01;
  assign sel_549569 = array_index_549552 == array_index_537032 ? add_549568 : sel_549565;
  assign add_549572 = sel_549569 + 8'h01;
  assign sel_549573 = array_index_549552 == array_index_537040 ? add_549572 : sel_549569;
  assign add_549576 = sel_549573 + 8'h01;
  assign sel_549577 = array_index_549552 == array_index_537048 ? add_549576 : sel_549573;
  assign add_549580 = sel_549577 + 8'h01;
  assign sel_549581 = array_index_549552 == array_index_537056 ? add_549580 : sel_549577;
  assign add_549584 = sel_549581 + 8'h01;
  assign sel_549585 = array_index_549552 == array_index_537064 ? add_549584 : sel_549581;
  assign add_549588 = sel_549585 + 8'h01;
  assign sel_549589 = array_index_549552 == array_index_537070 ? add_549588 : sel_549585;
  assign add_549592 = sel_549589 + 8'h01;
  assign sel_549593 = array_index_549552 == array_index_537076 ? add_549592 : sel_549589;
  assign add_549596 = sel_549593 + 8'h01;
  assign sel_549597 = array_index_549552 == array_index_537082 ? add_549596 : sel_549593;
  assign add_549600 = sel_549597 + 8'h01;
  assign sel_549601 = array_index_549552 == array_index_537088 ? add_549600 : sel_549597;
  assign add_549604 = sel_549601 + 8'h01;
  assign sel_549605 = array_index_549552 == array_index_537094 ? add_549604 : sel_549601;
  assign add_549608 = sel_549605 + 8'h01;
  assign sel_549609 = array_index_549552 == array_index_537100 ? add_549608 : sel_549605;
  assign add_549612 = sel_549609 + 8'h01;
  assign sel_549613 = array_index_549552 == array_index_537106 ? add_549612 : sel_549609;
  assign add_549616 = sel_549613 + 8'h01;
  assign sel_549617 = array_index_549552 == array_index_537112 ? add_549616 : sel_549613;
  assign add_549620 = sel_549617 + 8'h01;
  assign sel_549621 = array_index_549552 == array_index_537118 ? add_549620 : sel_549617;
  assign add_549624 = sel_549621 + 8'h01;
  assign sel_549625 = array_index_549552 == array_index_537124 ? add_549624 : sel_549621;
  assign add_549628 = sel_549625 + 8'h01;
  assign sel_549629 = array_index_549552 == array_index_537130 ? add_549628 : sel_549625;
  assign add_549632 = sel_549629 + 8'h01;
  assign sel_549633 = array_index_549552 == array_index_537136 ? add_549632 : sel_549629;
  assign add_549636 = sel_549633 + 8'h01;
  assign sel_549637 = array_index_549552 == array_index_537142 ? add_549636 : sel_549633;
  assign add_549640 = sel_549637 + 8'h01;
  assign sel_549641 = array_index_549552 == array_index_537148 ? add_549640 : sel_549637;
  assign add_549644 = sel_549641 + 8'h01;
  assign sel_549645 = array_index_549552 == array_index_537154 ? add_549644 : sel_549641;
  assign add_549648 = sel_549645 + 8'h01;
  assign sel_549649 = array_index_549552 == array_index_537160 ? add_549648 : sel_549645;
  assign add_549652 = sel_549649 + 8'h01;
  assign sel_549653 = array_index_549552 == array_index_537166 ? add_549652 : sel_549649;
  assign add_549656 = sel_549653 + 8'h01;
  assign sel_549657 = array_index_549552 == array_index_537172 ? add_549656 : sel_549653;
  assign add_549660 = sel_549657 + 8'h01;
  assign sel_549661 = array_index_549552 == array_index_537178 ? add_549660 : sel_549657;
  assign add_549664 = sel_549661 + 8'h01;
  assign sel_549665 = array_index_549552 == array_index_537184 ? add_549664 : sel_549661;
  assign add_549668 = sel_549665 + 8'h01;
  assign sel_549669 = array_index_549552 == array_index_537190 ? add_549668 : sel_549665;
  assign add_549672 = sel_549669 + 8'h01;
  assign sel_549673 = array_index_549552 == array_index_537196 ? add_549672 : sel_549669;
  assign add_549676 = sel_549673 + 8'h01;
  assign sel_549677 = array_index_549552 == array_index_537202 ? add_549676 : sel_549673;
  assign add_549680 = sel_549677 + 8'h01;
  assign sel_549681 = array_index_549552 == array_index_537208 ? add_549680 : sel_549677;
  assign add_549684 = sel_549681 + 8'h01;
  assign sel_549685 = array_index_549552 == array_index_537214 ? add_549684 : sel_549681;
  assign add_549688 = sel_549685 + 8'h01;
  assign sel_549689 = array_index_549552 == array_index_537220 ? add_549688 : sel_549685;
  assign add_549692 = sel_549689 + 8'h01;
  assign sel_549693 = array_index_549552 == array_index_537226 ? add_549692 : sel_549689;
  assign add_549696 = sel_549693 + 8'h01;
  assign sel_549697 = array_index_549552 == array_index_537232 ? add_549696 : sel_549693;
  assign add_549700 = sel_549697 + 8'h01;
  assign sel_549701 = array_index_549552 == array_index_537238 ? add_549700 : sel_549697;
  assign add_549704 = sel_549701 + 8'h01;
  assign sel_549705 = array_index_549552 == array_index_537244 ? add_549704 : sel_549701;
  assign add_549708 = sel_549705 + 8'h01;
  assign sel_549709 = array_index_549552 == array_index_537250 ? add_549708 : sel_549705;
  assign add_549712 = sel_549709 + 8'h01;
  assign sel_549713 = array_index_549552 == array_index_537256 ? add_549712 : sel_549709;
  assign add_549716 = sel_549713 + 8'h01;
  assign sel_549717 = array_index_549552 == array_index_537262 ? add_549716 : sel_549713;
  assign add_549720 = sel_549717 + 8'h01;
  assign sel_549721 = array_index_549552 == array_index_537268 ? add_549720 : sel_549717;
  assign add_549724 = sel_549721 + 8'h01;
  assign sel_549725 = array_index_549552 == array_index_537274 ? add_549724 : sel_549721;
  assign add_549728 = sel_549725 + 8'h01;
  assign sel_549729 = array_index_549552 == array_index_537280 ? add_549728 : sel_549725;
  assign add_549732 = sel_549729 + 8'h01;
  assign sel_549733 = array_index_549552 == array_index_537286 ? add_549732 : sel_549729;
  assign add_549736 = sel_549733 + 8'h01;
  assign sel_549737 = array_index_549552 == array_index_537292 ? add_549736 : sel_549733;
  assign add_549740 = sel_549737 + 8'h01;
  assign sel_549741 = array_index_549552 == array_index_537298 ? add_549740 : sel_549737;
  assign add_549744 = sel_549741 + 8'h01;
  assign sel_549745 = array_index_549552 == array_index_537304 ? add_549744 : sel_549741;
  assign add_549748 = sel_549745 + 8'h01;
  assign sel_549749 = array_index_549552 == array_index_537310 ? add_549748 : sel_549745;
  assign add_549752 = sel_549749 + 8'h01;
  assign sel_549753 = array_index_549552 == array_index_537316 ? add_549752 : sel_549749;
  assign add_549756 = sel_549753 + 8'h01;
  assign sel_549757 = array_index_549552 == array_index_537322 ? add_549756 : sel_549753;
  assign add_549760 = sel_549757 + 8'h01;
  assign sel_549761 = array_index_549552 == array_index_537328 ? add_549760 : sel_549757;
  assign add_549764 = sel_549761 + 8'h01;
  assign sel_549765 = array_index_549552 == array_index_537334 ? add_549764 : sel_549761;
  assign add_549768 = sel_549765 + 8'h01;
  assign sel_549769 = array_index_549552 == array_index_537340 ? add_549768 : sel_549765;
  assign add_549772 = sel_549769 + 8'h01;
  assign sel_549773 = array_index_549552 == array_index_537346 ? add_549772 : sel_549769;
  assign add_549776 = sel_549773 + 8'h01;
  assign sel_549777 = array_index_549552 == array_index_537352 ? add_549776 : sel_549773;
  assign add_549780 = sel_549777 + 8'h01;
  assign sel_549781 = array_index_549552 == array_index_537358 ? add_549780 : sel_549777;
  assign add_549784 = sel_549781 + 8'h01;
  assign sel_549785 = array_index_549552 == array_index_537364 ? add_549784 : sel_549781;
  assign add_549788 = sel_549785 + 8'h01;
  assign sel_549789 = array_index_549552 == array_index_537370 ? add_549788 : sel_549785;
  assign add_549792 = sel_549789 + 8'h01;
  assign sel_549793 = array_index_549552 == array_index_537376 ? add_549792 : sel_549789;
  assign add_549796 = sel_549793 + 8'h01;
  assign sel_549797 = array_index_549552 == array_index_537382 ? add_549796 : sel_549793;
  assign add_549800 = sel_549797 + 8'h01;
  assign sel_549801 = array_index_549552 == array_index_537388 ? add_549800 : sel_549797;
  assign add_549804 = sel_549801 + 8'h01;
  assign sel_549805 = array_index_549552 == array_index_537394 ? add_549804 : sel_549801;
  assign add_549808 = sel_549805 + 8'h01;
  assign sel_549809 = array_index_549552 == array_index_537400 ? add_549808 : sel_549805;
  assign add_549812 = sel_549809 + 8'h01;
  assign sel_549813 = array_index_549552 == array_index_537406 ? add_549812 : sel_549809;
  assign add_549816 = sel_549813 + 8'h01;
  assign sel_549817 = array_index_549552 == array_index_537412 ? add_549816 : sel_549813;
  assign add_549820 = sel_549817 + 8'h01;
  assign sel_549821 = array_index_549552 == array_index_537418 ? add_549820 : sel_549817;
  assign add_549824 = sel_549821 + 8'h01;
  assign sel_549825 = array_index_549552 == array_index_537424 ? add_549824 : sel_549821;
  assign add_549828 = sel_549825 + 8'h01;
  assign sel_549829 = array_index_549552 == array_index_537430 ? add_549828 : sel_549825;
  assign add_549832 = sel_549829 + 8'h01;
  assign sel_549833 = array_index_549552 == array_index_537436 ? add_549832 : sel_549829;
  assign add_549836 = sel_549833 + 8'h01;
  assign sel_549837 = array_index_549552 == array_index_537442 ? add_549836 : sel_549833;
  assign add_549840 = sel_549837 + 8'h01;
  assign sel_549841 = array_index_549552 == array_index_537448 ? add_549840 : sel_549837;
  assign add_549844 = sel_549841 + 8'h01;
  assign sel_549845 = array_index_549552 == array_index_537454 ? add_549844 : sel_549841;
  assign add_549848 = sel_549845 + 8'h01;
  assign sel_549849 = array_index_549552 == array_index_537460 ? add_549848 : sel_549845;
  assign add_549853 = sel_549849 + 8'h01;
  assign array_index_549854 = set1_unflattened[7'h2a];
  assign sel_549855 = array_index_549552 == array_index_537466 ? add_549853 : sel_549849;
  assign add_549858 = sel_549855 + 8'h01;
  assign sel_549859 = array_index_549854 == array_index_537012 ? add_549858 : sel_549855;
  assign add_549862 = sel_549859 + 8'h01;
  assign sel_549863 = array_index_549854 == array_index_537016 ? add_549862 : sel_549859;
  assign add_549866 = sel_549863 + 8'h01;
  assign sel_549867 = array_index_549854 == array_index_537024 ? add_549866 : sel_549863;
  assign add_549870 = sel_549867 + 8'h01;
  assign sel_549871 = array_index_549854 == array_index_537032 ? add_549870 : sel_549867;
  assign add_549874 = sel_549871 + 8'h01;
  assign sel_549875 = array_index_549854 == array_index_537040 ? add_549874 : sel_549871;
  assign add_549878 = sel_549875 + 8'h01;
  assign sel_549879 = array_index_549854 == array_index_537048 ? add_549878 : sel_549875;
  assign add_549882 = sel_549879 + 8'h01;
  assign sel_549883 = array_index_549854 == array_index_537056 ? add_549882 : sel_549879;
  assign add_549886 = sel_549883 + 8'h01;
  assign sel_549887 = array_index_549854 == array_index_537064 ? add_549886 : sel_549883;
  assign add_549890 = sel_549887 + 8'h01;
  assign sel_549891 = array_index_549854 == array_index_537070 ? add_549890 : sel_549887;
  assign add_549894 = sel_549891 + 8'h01;
  assign sel_549895 = array_index_549854 == array_index_537076 ? add_549894 : sel_549891;
  assign add_549898 = sel_549895 + 8'h01;
  assign sel_549899 = array_index_549854 == array_index_537082 ? add_549898 : sel_549895;
  assign add_549902 = sel_549899 + 8'h01;
  assign sel_549903 = array_index_549854 == array_index_537088 ? add_549902 : sel_549899;
  assign add_549906 = sel_549903 + 8'h01;
  assign sel_549907 = array_index_549854 == array_index_537094 ? add_549906 : sel_549903;
  assign add_549910 = sel_549907 + 8'h01;
  assign sel_549911 = array_index_549854 == array_index_537100 ? add_549910 : sel_549907;
  assign add_549914 = sel_549911 + 8'h01;
  assign sel_549915 = array_index_549854 == array_index_537106 ? add_549914 : sel_549911;
  assign add_549918 = sel_549915 + 8'h01;
  assign sel_549919 = array_index_549854 == array_index_537112 ? add_549918 : sel_549915;
  assign add_549922 = sel_549919 + 8'h01;
  assign sel_549923 = array_index_549854 == array_index_537118 ? add_549922 : sel_549919;
  assign add_549926 = sel_549923 + 8'h01;
  assign sel_549927 = array_index_549854 == array_index_537124 ? add_549926 : sel_549923;
  assign add_549930 = sel_549927 + 8'h01;
  assign sel_549931 = array_index_549854 == array_index_537130 ? add_549930 : sel_549927;
  assign add_549934 = sel_549931 + 8'h01;
  assign sel_549935 = array_index_549854 == array_index_537136 ? add_549934 : sel_549931;
  assign add_549938 = sel_549935 + 8'h01;
  assign sel_549939 = array_index_549854 == array_index_537142 ? add_549938 : sel_549935;
  assign add_549942 = sel_549939 + 8'h01;
  assign sel_549943 = array_index_549854 == array_index_537148 ? add_549942 : sel_549939;
  assign add_549946 = sel_549943 + 8'h01;
  assign sel_549947 = array_index_549854 == array_index_537154 ? add_549946 : sel_549943;
  assign add_549950 = sel_549947 + 8'h01;
  assign sel_549951 = array_index_549854 == array_index_537160 ? add_549950 : sel_549947;
  assign add_549954 = sel_549951 + 8'h01;
  assign sel_549955 = array_index_549854 == array_index_537166 ? add_549954 : sel_549951;
  assign add_549958 = sel_549955 + 8'h01;
  assign sel_549959 = array_index_549854 == array_index_537172 ? add_549958 : sel_549955;
  assign add_549962 = sel_549959 + 8'h01;
  assign sel_549963 = array_index_549854 == array_index_537178 ? add_549962 : sel_549959;
  assign add_549966 = sel_549963 + 8'h01;
  assign sel_549967 = array_index_549854 == array_index_537184 ? add_549966 : sel_549963;
  assign add_549970 = sel_549967 + 8'h01;
  assign sel_549971 = array_index_549854 == array_index_537190 ? add_549970 : sel_549967;
  assign add_549974 = sel_549971 + 8'h01;
  assign sel_549975 = array_index_549854 == array_index_537196 ? add_549974 : sel_549971;
  assign add_549978 = sel_549975 + 8'h01;
  assign sel_549979 = array_index_549854 == array_index_537202 ? add_549978 : sel_549975;
  assign add_549982 = sel_549979 + 8'h01;
  assign sel_549983 = array_index_549854 == array_index_537208 ? add_549982 : sel_549979;
  assign add_549986 = sel_549983 + 8'h01;
  assign sel_549987 = array_index_549854 == array_index_537214 ? add_549986 : sel_549983;
  assign add_549990 = sel_549987 + 8'h01;
  assign sel_549991 = array_index_549854 == array_index_537220 ? add_549990 : sel_549987;
  assign add_549994 = sel_549991 + 8'h01;
  assign sel_549995 = array_index_549854 == array_index_537226 ? add_549994 : sel_549991;
  assign add_549998 = sel_549995 + 8'h01;
  assign sel_549999 = array_index_549854 == array_index_537232 ? add_549998 : sel_549995;
  assign add_550002 = sel_549999 + 8'h01;
  assign sel_550003 = array_index_549854 == array_index_537238 ? add_550002 : sel_549999;
  assign add_550006 = sel_550003 + 8'h01;
  assign sel_550007 = array_index_549854 == array_index_537244 ? add_550006 : sel_550003;
  assign add_550010 = sel_550007 + 8'h01;
  assign sel_550011 = array_index_549854 == array_index_537250 ? add_550010 : sel_550007;
  assign add_550014 = sel_550011 + 8'h01;
  assign sel_550015 = array_index_549854 == array_index_537256 ? add_550014 : sel_550011;
  assign add_550018 = sel_550015 + 8'h01;
  assign sel_550019 = array_index_549854 == array_index_537262 ? add_550018 : sel_550015;
  assign add_550022 = sel_550019 + 8'h01;
  assign sel_550023 = array_index_549854 == array_index_537268 ? add_550022 : sel_550019;
  assign add_550026 = sel_550023 + 8'h01;
  assign sel_550027 = array_index_549854 == array_index_537274 ? add_550026 : sel_550023;
  assign add_550030 = sel_550027 + 8'h01;
  assign sel_550031 = array_index_549854 == array_index_537280 ? add_550030 : sel_550027;
  assign add_550034 = sel_550031 + 8'h01;
  assign sel_550035 = array_index_549854 == array_index_537286 ? add_550034 : sel_550031;
  assign add_550038 = sel_550035 + 8'h01;
  assign sel_550039 = array_index_549854 == array_index_537292 ? add_550038 : sel_550035;
  assign add_550042 = sel_550039 + 8'h01;
  assign sel_550043 = array_index_549854 == array_index_537298 ? add_550042 : sel_550039;
  assign add_550046 = sel_550043 + 8'h01;
  assign sel_550047 = array_index_549854 == array_index_537304 ? add_550046 : sel_550043;
  assign add_550050 = sel_550047 + 8'h01;
  assign sel_550051 = array_index_549854 == array_index_537310 ? add_550050 : sel_550047;
  assign add_550054 = sel_550051 + 8'h01;
  assign sel_550055 = array_index_549854 == array_index_537316 ? add_550054 : sel_550051;
  assign add_550058 = sel_550055 + 8'h01;
  assign sel_550059 = array_index_549854 == array_index_537322 ? add_550058 : sel_550055;
  assign add_550062 = sel_550059 + 8'h01;
  assign sel_550063 = array_index_549854 == array_index_537328 ? add_550062 : sel_550059;
  assign add_550066 = sel_550063 + 8'h01;
  assign sel_550067 = array_index_549854 == array_index_537334 ? add_550066 : sel_550063;
  assign add_550070 = sel_550067 + 8'h01;
  assign sel_550071 = array_index_549854 == array_index_537340 ? add_550070 : sel_550067;
  assign add_550074 = sel_550071 + 8'h01;
  assign sel_550075 = array_index_549854 == array_index_537346 ? add_550074 : sel_550071;
  assign add_550078 = sel_550075 + 8'h01;
  assign sel_550079 = array_index_549854 == array_index_537352 ? add_550078 : sel_550075;
  assign add_550082 = sel_550079 + 8'h01;
  assign sel_550083 = array_index_549854 == array_index_537358 ? add_550082 : sel_550079;
  assign add_550086 = sel_550083 + 8'h01;
  assign sel_550087 = array_index_549854 == array_index_537364 ? add_550086 : sel_550083;
  assign add_550090 = sel_550087 + 8'h01;
  assign sel_550091 = array_index_549854 == array_index_537370 ? add_550090 : sel_550087;
  assign add_550094 = sel_550091 + 8'h01;
  assign sel_550095 = array_index_549854 == array_index_537376 ? add_550094 : sel_550091;
  assign add_550098 = sel_550095 + 8'h01;
  assign sel_550099 = array_index_549854 == array_index_537382 ? add_550098 : sel_550095;
  assign add_550102 = sel_550099 + 8'h01;
  assign sel_550103 = array_index_549854 == array_index_537388 ? add_550102 : sel_550099;
  assign add_550106 = sel_550103 + 8'h01;
  assign sel_550107 = array_index_549854 == array_index_537394 ? add_550106 : sel_550103;
  assign add_550110 = sel_550107 + 8'h01;
  assign sel_550111 = array_index_549854 == array_index_537400 ? add_550110 : sel_550107;
  assign add_550114 = sel_550111 + 8'h01;
  assign sel_550115 = array_index_549854 == array_index_537406 ? add_550114 : sel_550111;
  assign add_550118 = sel_550115 + 8'h01;
  assign sel_550119 = array_index_549854 == array_index_537412 ? add_550118 : sel_550115;
  assign add_550122 = sel_550119 + 8'h01;
  assign sel_550123 = array_index_549854 == array_index_537418 ? add_550122 : sel_550119;
  assign add_550126 = sel_550123 + 8'h01;
  assign sel_550127 = array_index_549854 == array_index_537424 ? add_550126 : sel_550123;
  assign add_550130 = sel_550127 + 8'h01;
  assign sel_550131 = array_index_549854 == array_index_537430 ? add_550130 : sel_550127;
  assign add_550134 = sel_550131 + 8'h01;
  assign sel_550135 = array_index_549854 == array_index_537436 ? add_550134 : sel_550131;
  assign add_550138 = sel_550135 + 8'h01;
  assign sel_550139 = array_index_549854 == array_index_537442 ? add_550138 : sel_550135;
  assign add_550142 = sel_550139 + 8'h01;
  assign sel_550143 = array_index_549854 == array_index_537448 ? add_550142 : sel_550139;
  assign add_550146 = sel_550143 + 8'h01;
  assign sel_550147 = array_index_549854 == array_index_537454 ? add_550146 : sel_550143;
  assign add_550150 = sel_550147 + 8'h01;
  assign sel_550151 = array_index_549854 == array_index_537460 ? add_550150 : sel_550147;
  assign add_550155 = sel_550151 + 8'h01;
  assign array_index_550156 = set1_unflattened[7'h2b];
  assign sel_550157 = array_index_549854 == array_index_537466 ? add_550155 : sel_550151;
  assign add_550160 = sel_550157 + 8'h01;
  assign sel_550161 = array_index_550156 == array_index_537012 ? add_550160 : sel_550157;
  assign add_550164 = sel_550161 + 8'h01;
  assign sel_550165 = array_index_550156 == array_index_537016 ? add_550164 : sel_550161;
  assign add_550168 = sel_550165 + 8'h01;
  assign sel_550169 = array_index_550156 == array_index_537024 ? add_550168 : sel_550165;
  assign add_550172 = sel_550169 + 8'h01;
  assign sel_550173 = array_index_550156 == array_index_537032 ? add_550172 : sel_550169;
  assign add_550176 = sel_550173 + 8'h01;
  assign sel_550177 = array_index_550156 == array_index_537040 ? add_550176 : sel_550173;
  assign add_550180 = sel_550177 + 8'h01;
  assign sel_550181 = array_index_550156 == array_index_537048 ? add_550180 : sel_550177;
  assign add_550184 = sel_550181 + 8'h01;
  assign sel_550185 = array_index_550156 == array_index_537056 ? add_550184 : sel_550181;
  assign add_550188 = sel_550185 + 8'h01;
  assign sel_550189 = array_index_550156 == array_index_537064 ? add_550188 : sel_550185;
  assign add_550192 = sel_550189 + 8'h01;
  assign sel_550193 = array_index_550156 == array_index_537070 ? add_550192 : sel_550189;
  assign add_550196 = sel_550193 + 8'h01;
  assign sel_550197 = array_index_550156 == array_index_537076 ? add_550196 : sel_550193;
  assign add_550200 = sel_550197 + 8'h01;
  assign sel_550201 = array_index_550156 == array_index_537082 ? add_550200 : sel_550197;
  assign add_550204 = sel_550201 + 8'h01;
  assign sel_550205 = array_index_550156 == array_index_537088 ? add_550204 : sel_550201;
  assign add_550208 = sel_550205 + 8'h01;
  assign sel_550209 = array_index_550156 == array_index_537094 ? add_550208 : sel_550205;
  assign add_550212 = sel_550209 + 8'h01;
  assign sel_550213 = array_index_550156 == array_index_537100 ? add_550212 : sel_550209;
  assign add_550216 = sel_550213 + 8'h01;
  assign sel_550217 = array_index_550156 == array_index_537106 ? add_550216 : sel_550213;
  assign add_550220 = sel_550217 + 8'h01;
  assign sel_550221 = array_index_550156 == array_index_537112 ? add_550220 : sel_550217;
  assign add_550224 = sel_550221 + 8'h01;
  assign sel_550225 = array_index_550156 == array_index_537118 ? add_550224 : sel_550221;
  assign add_550228 = sel_550225 + 8'h01;
  assign sel_550229 = array_index_550156 == array_index_537124 ? add_550228 : sel_550225;
  assign add_550232 = sel_550229 + 8'h01;
  assign sel_550233 = array_index_550156 == array_index_537130 ? add_550232 : sel_550229;
  assign add_550236 = sel_550233 + 8'h01;
  assign sel_550237 = array_index_550156 == array_index_537136 ? add_550236 : sel_550233;
  assign add_550240 = sel_550237 + 8'h01;
  assign sel_550241 = array_index_550156 == array_index_537142 ? add_550240 : sel_550237;
  assign add_550244 = sel_550241 + 8'h01;
  assign sel_550245 = array_index_550156 == array_index_537148 ? add_550244 : sel_550241;
  assign add_550248 = sel_550245 + 8'h01;
  assign sel_550249 = array_index_550156 == array_index_537154 ? add_550248 : sel_550245;
  assign add_550252 = sel_550249 + 8'h01;
  assign sel_550253 = array_index_550156 == array_index_537160 ? add_550252 : sel_550249;
  assign add_550256 = sel_550253 + 8'h01;
  assign sel_550257 = array_index_550156 == array_index_537166 ? add_550256 : sel_550253;
  assign add_550260 = sel_550257 + 8'h01;
  assign sel_550261 = array_index_550156 == array_index_537172 ? add_550260 : sel_550257;
  assign add_550264 = sel_550261 + 8'h01;
  assign sel_550265 = array_index_550156 == array_index_537178 ? add_550264 : sel_550261;
  assign add_550268 = sel_550265 + 8'h01;
  assign sel_550269 = array_index_550156 == array_index_537184 ? add_550268 : sel_550265;
  assign add_550272 = sel_550269 + 8'h01;
  assign sel_550273 = array_index_550156 == array_index_537190 ? add_550272 : sel_550269;
  assign add_550276 = sel_550273 + 8'h01;
  assign sel_550277 = array_index_550156 == array_index_537196 ? add_550276 : sel_550273;
  assign add_550280 = sel_550277 + 8'h01;
  assign sel_550281 = array_index_550156 == array_index_537202 ? add_550280 : sel_550277;
  assign add_550284 = sel_550281 + 8'h01;
  assign sel_550285 = array_index_550156 == array_index_537208 ? add_550284 : sel_550281;
  assign add_550288 = sel_550285 + 8'h01;
  assign sel_550289 = array_index_550156 == array_index_537214 ? add_550288 : sel_550285;
  assign add_550292 = sel_550289 + 8'h01;
  assign sel_550293 = array_index_550156 == array_index_537220 ? add_550292 : sel_550289;
  assign add_550296 = sel_550293 + 8'h01;
  assign sel_550297 = array_index_550156 == array_index_537226 ? add_550296 : sel_550293;
  assign add_550300 = sel_550297 + 8'h01;
  assign sel_550301 = array_index_550156 == array_index_537232 ? add_550300 : sel_550297;
  assign add_550304 = sel_550301 + 8'h01;
  assign sel_550305 = array_index_550156 == array_index_537238 ? add_550304 : sel_550301;
  assign add_550308 = sel_550305 + 8'h01;
  assign sel_550309 = array_index_550156 == array_index_537244 ? add_550308 : sel_550305;
  assign add_550312 = sel_550309 + 8'h01;
  assign sel_550313 = array_index_550156 == array_index_537250 ? add_550312 : sel_550309;
  assign add_550316 = sel_550313 + 8'h01;
  assign sel_550317 = array_index_550156 == array_index_537256 ? add_550316 : sel_550313;
  assign add_550320 = sel_550317 + 8'h01;
  assign sel_550321 = array_index_550156 == array_index_537262 ? add_550320 : sel_550317;
  assign add_550324 = sel_550321 + 8'h01;
  assign sel_550325 = array_index_550156 == array_index_537268 ? add_550324 : sel_550321;
  assign add_550328 = sel_550325 + 8'h01;
  assign sel_550329 = array_index_550156 == array_index_537274 ? add_550328 : sel_550325;
  assign add_550332 = sel_550329 + 8'h01;
  assign sel_550333 = array_index_550156 == array_index_537280 ? add_550332 : sel_550329;
  assign add_550336 = sel_550333 + 8'h01;
  assign sel_550337 = array_index_550156 == array_index_537286 ? add_550336 : sel_550333;
  assign add_550340 = sel_550337 + 8'h01;
  assign sel_550341 = array_index_550156 == array_index_537292 ? add_550340 : sel_550337;
  assign add_550344 = sel_550341 + 8'h01;
  assign sel_550345 = array_index_550156 == array_index_537298 ? add_550344 : sel_550341;
  assign add_550348 = sel_550345 + 8'h01;
  assign sel_550349 = array_index_550156 == array_index_537304 ? add_550348 : sel_550345;
  assign add_550352 = sel_550349 + 8'h01;
  assign sel_550353 = array_index_550156 == array_index_537310 ? add_550352 : sel_550349;
  assign add_550356 = sel_550353 + 8'h01;
  assign sel_550357 = array_index_550156 == array_index_537316 ? add_550356 : sel_550353;
  assign add_550360 = sel_550357 + 8'h01;
  assign sel_550361 = array_index_550156 == array_index_537322 ? add_550360 : sel_550357;
  assign add_550364 = sel_550361 + 8'h01;
  assign sel_550365 = array_index_550156 == array_index_537328 ? add_550364 : sel_550361;
  assign add_550368 = sel_550365 + 8'h01;
  assign sel_550369 = array_index_550156 == array_index_537334 ? add_550368 : sel_550365;
  assign add_550372 = sel_550369 + 8'h01;
  assign sel_550373 = array_index_550156 == array_index_537340 ? add_550372 : sel_550369;
  assign add_550376 = sel_550373 + 8'h01;
  assign sel_550377 = array_index_550156 == array_index_537346 ? add_550376 : sel_550373;
  assign add_550380 = sel_550377 + 8'h01;
  assign sel_550381 = array_index_550156 == array_index_537352 ? add_550380 : sel_550377;
  assign add_550384 = sel_550381 + 8'h01;
  assign sel_550385 = array_index_550156 == array_index_537358 ? add_550384 : sel_550381;
  assign add_550388 = sel_550385 + 8'h01;
  assign sel_550389 = array_index_550156 == array_index_537364 ? add_550388 : sel_550385;
  assign add_550392 = sel_550389 + 8'h01;
  assign sel_550393 = array_index_550156 == array_index_537370 ? add_550392 : sel_550389;
  assign add_550396 = sel_550393 + 8'h01;
  assign sel_550397 = array_index_550156 == array_index_537376 ? add_550396 : sel_550393;
  assign add_550400 = sel_550397 + 8'h01;
  assign sel_550401 = array_index_550156 == array_index_537382 ? add_550400 : sel_550397;
  assign add_550404 = sel_550401 + 8'h01;
  assign sel_550405 = array_index_550156 == array_index_537388 ? add_550404 : sel_550401;
  assign add_550408 = sel_550405 + 8'h01;
  assign sel_550409 = array_index_550156 == array_index_537394 ? add_550408 : sel_550405;
  assign add_550412 = sel_550409 + 8'h01;
  assign sel_550413 = array_index_550156 == array_index_537400 ? add_550412 : sel_550409;
  assign add_550416 = sel_550413 + 8'h01;
  assign sel_550417 = array_index_550156 == array_index_537406 ? add_550416 : sel_550413;
  assign add_550420 = sel_550417 + 8'h01;
  assign sel_550421 = array_index_550156 == array_index_537412 ? add_550420 : sel_550417;
  assign add_550424 = sel_550421 + 8'h01;
  assign sel_550425 = array_index_550156 == array_index_537418 ? add_550424 : sel_550421;
  assign add_550428 = sel_550425 + 8'h01;
  assign sel_550429 = array_index_550156 == array_index_537424 ? add_550428 : sel_550425;
  assign add_550432 = sel_550429 + 8'h01;
  assign sel_550433 = array_index_550156 == array_index_537430 ? add_550432 : sel_550429;
  assign add_550436 = sel_550433 + 8'h01;
  assign sel_550437 = array_index_550156 == array_index_537436 ? add_550436 : sel_550433;
  assign add_550440 = sel_550437 + 8'h01;
  assign sel_550441 = array_index_550156 == array_index_537442 ? add_550440 : sel_550437;
  assign add_550444 = sel_550441 + 8'h01;
  assign sel_550445 = array_index_550156 == array_index_537448 ? add_550444 : sel_550441;
  assign add_550448 = sel_550445 + 8'h01;
  assign sel_550449 = array_index_550156 == array_index_537454 ? add_550448 : sel_550445;
  assign add_550452 = sel_550449 + 8'h01;
  assign sel_550453 = array_index_550156 == array_index_537460 ? add_550452 : sel_550449;
  assign add_550457 = sel_550453 + 8'h01;
  assign array_index_550458 = set1_unflattened[7'h2c];
  assign sel_550459 = array_index_550156 == array_index_537466 ? add_550457 : sel_550453;
  assign add_550462 = sel_550459 + 8'h01;
  assign sel_550463 = array_index_550458 == array_index_537012 ? add_550462 : sel_550459;
  assign add_550466 = sel_550463 + 8'h01;
  assign sel_550467 = array_index_550458 == array_index_537016 ? add_550466 : sel_550463;
  assign add_550470 = sel_550467 + 8'h01;
  assign sel_550471 = array_index_550458 == array_index_537024 ? add_550470 : sel_550467;
  assign add_550474 = sel_550471 + 8'h01;
  assign sel_550475 = array_index_550458 == array_index_537032 ? add_550474 : sel_550471;
  assign add_550478 = sel_550475 + 8'h01;
  assign sel_550479 = array_index_550458 == array_index_537040 ? add_550478 : sel_550475;
  assign add_550482 = sel_550479 + 8'h01;
  assign sel_550483 = array_index_550458 == array_index_537048 ? add_550482 : sel_550479;
  assign add_550486 = sel_550483 + 8'h01;
  assign sel_550487 = array_index_550458 == array_index_537056 ? add_550486 : sel_550483;
  assign add_550490 = sel_550487 + 8'h01;
  assign sel_550491 = array_index_550458 == array_index_537064 ? add_550490 : sel_550487;
  assign add_550494 = sel_550491 + 8'h01;
  assign sel_550495 = array_index_550458 == array_index_537070 ? add_550494 : sel_550491;
  assign add_550498 = sel_550495 + 8'h01;
  assign sel_550499 = array_index_550458 == array_index_537076 ? add_550498 : sel_550495;
  assign add_550502 = sel_550499 + 8'h01;
  assign sel_550503 = array_index_550458 == array_index_537082 ? add_550502 : sel_550499;
  assign add_550506 = sel_550503 + 8'h01;
  assign sel_550507 = array_index_550458 == array_index_537088 ? add_550506 : sel_550503;
  assign add_550510 = sel_550507 + 8'h01;
  assign sel_550511 = array_index_550458 == array_index_537094 ? add_550510 : sel_550507;
  assign add_550514 = sel_550511 + 8'h01;
  assign sel_550515 = array_index_550458 == array_index_537100 ? add_550514 : sel_550511;
  assign add_550518 = sel_550515 + 8'h01;
  assign sel_550519 = array_index_550458 == array_index_537106 ? add_550518 : sel_550515;
  assign add_550522 = sel_550519 + 8'h01;
  assign sel_550523 = array_index_550458 == array_index_537112 ? add_550522 : sel_550519;
  assign add_550526 = sel_550523 + 8'h01;
  assign sel_550527 = array_index_550458 == array_index_537118 ? add_550526 : sel_550523;
  assign add_550530 = sel_550527 + 8'h01;
  assign sel_550531 = array_index_550458 == array_index_537124 ? add_550530 : sel_550527;
  assign add_550534 = sel_550531 + 8'h01;
  assign sel_550535 = array_index_550458 == array_index_537130 ? add_550534 : sel_550531;
  assign add_550538 = sel_550535 + 8'h01;
  assign sel_550539 = array_index_550458 == array_index_537136 ? add_550538 : sel_550535;
  assign add_550542 = sel_550539 + 8'h01;
  assign sel_550543 = array_index_550458 == array_index_537142 ? add_550542 : sel_550539;
  assign add_550546 = sel_550543 + 8'h01;
  assign sel_550547 = array_index_550458 == array_index_537148 ? add_550546 : sel_550543;
  assign add_550550 = sel_550547 + 8'h01;
  assign sel_550551 = array_index_550458 == array_index_537154 ? add_550550 : sel_550547;
  assign add_550554 = sel_550551 + 8'h01;
  assign sel_550555 = array_index_550458 == array_index_537160 ? add_550554 : sel_550551;
  assign add_550558 = sel_550555 + 8'h01;
  assign sel_550559 = array_index_550458 == array_index_537166 ? add_550558 : sel_550555;
  assign add_550562 = sel_550559 + 8'h01;
  assign sel_550563 = array_index_550458 == array_index_537172 ? add_550562 : sel_550559;
  assign add_550566 = sel_550563 + 8'h01;
  assign sel_550567 = array_index_550458 == array_index_537178 ? add_550566 : sel_550563;
  assign add_550570 = sel_550567 + 8'h01;
  assign sel_550571 = array_index_550458 == array_index_537184 ? add_550570 : sel_550567;
  assign add_550574 = sel_550571 + 8'h01;
  assign sel_550575 = array_index_550458 == array_index_537190 ? add_550574 : sel_550571;
  assign add_550578 = sel_550575 + 8'h01;
  assign sel_550579 = array_index_550458 == array_index_537196 ? add_550578 : sel_550575;
  assign add_550582 = sel_550579 + 8'h01;
  assign sel_550583 = array_index_550458 == array_index_537202 ? add_550582 : sel_550579;
  assign add_550586 = sel_550583 + 8'h01;
  assign sel_550587 = array_index_550458 == array_index_537208 ? add_550586 : sel_550583;
  assign add_550590 = sel_550587 + 8'h01;
  assign sel_550591 = array_index_550458 == array_index_537214 ? add_550590 : sel_550587;
  assign add_550594 = sel_550591 + 8'h01;
  assign sel_550595 = array_index_550458 == array_index_537220 ? add_550594 : sel_550591;
  assign add_550598 = sel_550595 + 8'h01;
  assign sel_550599 = array_index_550458 == array_index_537226 ? add_550598 : sel_550595;
  assign add_550602 = sel_550599 + 8'h01;
  assign sel_550603 = array_index_550458 == array_index_537232 ? add_550602 : sel_550599;
  assign add_550606 = sel_550603 + 8'h01;
  assign sel_550607 = array_index_550458 == array_index_537238 ? add_550606 : sel_550603;
  assign add_550610 = sel_550607 + 8'h01;
  assign sel_550611 = array_index_550458 == array_index_537244 ? add_550610 : sel_550607;
  assign add_550614 = sel_550611 + 8'h01;
  assign sel_550615 = array_index_550458 == array_index_537250 ? add_550614 : sel_550611;
  assign add_550618 = sel_550615 + 8'h01;
  assign sel_550619 = array_index_550458 == array_index_537256 ? add_550618 : sel_550615;
  assign add_550622 = sel_550619 + 8'h01;
  assign sel_550623 = array_index_550458 == array_index_537262 ? add_550622 : sel_550619;
  assign add_550626 = sel_550623 + 8'h01;
  assign sel_550627 = array_index_550458 == array_index_537268 ? add_550626 : sel_550623;
  assign add_550630 = sel_550627 + 8'h01;
  assign sel_550631 = array_index_550458 == array_index_537274 ? add_550630 : sel_550627;
  assign add_550634 = sel_550631 + 8'h01;
  assign sel_550635 = array_index_550458 == array_index_537280 ? add_550634 : sel_550631;
  assign add_550638 = sel_550635 + 8'h01;
  assign sel_550639 = array_index_550458 == array_index_537286 ? add_550638 : sel_550635;
  assign add_550642 = sel_550639 + 8'h01;
  assign sel_550643 = array_index_550458 == array_index_537292 ? add_550642 : sel_550639;
  assign add_550646 = sel_550643 + 8'h01;
  assign sel_550647 = array_index_550458 == array_index_537298 ? add_550646 : sel_550643;
  assign add_550650 = sel_550647 + 8'h01;
  assign sel_550651 = array_index_550458 == array_index_537304 ? add_550650 : sel_550647;
  assign add_550654 = sel_550651 + 8'h01;
  assign sel_550655 = array_index_550458 == array_index_537310 ? add_550654 : sel_550651;
  assign add_550658 = sel_550655 + 8'h01;
  assign sel_550659 = array_index_550458 == array_index_537316 ? add_550658 : sel_550655;
  assign add_550662 = sel_550659 + 8'h01;
  assign sel_550663 = array_index_550458 == array_index_537322 ? add_550662 : sel_550659;
  assign add_550666 = sel_550663 + 8'h01;
  assign sel_550667 = array_index_550458 == array_index_537328 ? add_550666 : sel_550663;
  assign add_550670 = sel_550667 + 8'h01;
  assign sel_550671 = array_index_550458 == array_index_537334 ? add_550670 : sel_550667;
  assign add_550674 = sel_550671 + 8'h01;
  assign sel_550675 = array_index_550458 == array_index_537340 ? add_550674 : sel_550671;
  assign add_550678 = sel_550675 + 8'h01;
  assign sel_550679 = array_index_550458 == array_index_537346 ? add_550678 : sel_550675;
  assign add_550682 = sel_550679 + 8'h01;
  assign sel_550683 = array_index_550458 == array_index_537352 ? add_550682 : sel_550679;
  assign add_550686 = sel_550683 + 8'h01;
  assign sel_550687 = array_index_550458 == array_index_537358 ? add_550686 : sel_550683;
  assign add_550690 = sel_550687 + 8'h01;
  assign sel_550691 = array_index_550458 == array_index_537364 ? add_550690 : sel_550687;
  assign add_550694 = sel_550691 + 8'h01;
  assign sel_550695 = array_index_550458 == array_index_537370 ? add_550694 : sel_550691;
  assign add_550698 = sel_550695 + 8'h01;
  assign sel_550699 = array_index_550458 == array_index_537376 ? add_550698 : sel_550695;
  assign add_550702 = sel_550699 + 8'h01;
  assign sel_550703 = array_index_550458 == array_index_537382 ? add_550702 : sel_550699;
  assign add_550706 = sel_550703 + 8'h01;
  assign sel_550707 = array_index_550458 == array_index_537388 ? add_550706 : sel_550703;
  assign add_550710 = sel_550707 + 8'h01;
  assign sel_550711 = array_index_550458 == array_index_537394 ? add_550710 : sel_550707;
  assign add_550714 = sel_550711 + 8'h01;
  assign sel_550715 = array_index_550458 == array_index_537400 ? add_550714 : sel_550711;
  assign add_550718 = sel_550715 + 8'h01;
  assign sel_550719 = array_index_550458 == array_index_537406 ? add_550718 : sel_550715;
  assign add_550722 = sel_550719 + 8'h01;
  assign sel_550723 = array_index_550458 == array_index_537412 ? add_550722 : sel_550719;
  assign add_550726 = sel_550723 + 8'h01;
  assign sel_550727 = array_index_550458 == array_index_537418 ? add_550726 : sel_550723;
  assign add_550730 = sel_550727 + 8'h01;
  assign sel_550731 = array_index_550458 == array_index_537424 ? add_550730 : sel_550727;
  assign add_550734 = sel_550731 + 8'h01;
  assign sel_550735 = array_index_550458 == array_index_537430 ? add_550734 : sel_550731;
  assign add_550738 = sel_550735 + 8'h01;
  assign sel_550739 = array_index_550458 == array_index_537436 ? add_550738 : sel_550735;
  assign add_550742 = sel_550739 + 8'h01;
  assign sel_550743 = array_index_550458 == array_index_537442 ? add_550742 : sel_550739;
  assign add_550746 = sel_550743 + 8'h01;
  assign sel_550747 = array_index_550458 == array_index_537448 ? add_550746 : sel_550743;
  assign add_550750 = sel_550747 + 8'h01;
  assign sel_550751 = array_index_550458 == array_index_537454 ? add_550750 : sel_550747;
  assign add_550754 = sel_550751 + 8'h01;
  assign sel_550755 = array_index_550458 == array_index_537460 ? add_550754 : sel_550751;
  assign add_550759 = sel_550755 + 8'h01;
  assign array_index_550760 = set1_unflattened[7'h2d];
  assign sel_550761 = array_index_550458 == array_index_537466 ? add_550759 : sel_550755;
  assign add_550764 = sel_550761 + 8'h01;
  assign sel_550765 = array_index_550760 == array_index_537012 ? add_550764 : sel_550761;
  assign add_550768 = sel_550765 + 8'h01;
  assign sel_550769 = array_index_550760 == array_index_537016 ? add_550768 : sel_550765;
  assign add_550772 = sel_550769 + 8'h01;
  assign sel_550773 = array_index_550760 == array_index_537024 ? add_550772 : sel_550769;
  assign add_550776 = sel_550773 + 8'h01;
  assign sel_550777 = array_index_550760 == array_index_537032 ? add_550776 : sel_550773;
  assign add_550780 = sel_550777 + 8'h01;
  assign sel_550781 = array_index_550760 == array_index_537040 ? add_550780 : sel_550777;
  assign add_550784 = sel_550781 + 8'h01;
  assign sel_550785 = array_index_550760 == array_index_537048 ? add_550784 : sel_550781;
  assign add_550788 = sel_550785 + 8'h01;
  assign sel_550789 = array_index_550760 == array_index_537056 ? add_550788 : sel_550785;
  assign add_550792 = sel_550789 + 8'h01;
  assign sel_550793 = array_index_550760 == array_index_537064 ? add_550792 : sel_550789;
  assign add_550796 = sel_550793 + 8'h01;
  assign sel_550797 = array_index_550760 == array_index_537070 ? add_550796 : sel_550793;
  assign add_550800 = sel_550797 + 8'h01;
  assign sel_550801 = array_index_550760 == array_index_537076 ? add_550800 : sel_550797;
  assign add_550804 = sel_550801 + 8'h01;
  assign sel_550805 = array_index_550760 == array_index_537082 ? add_550804 : sel_550801;
  assign add_550808 = sel_550805 + 8'h01;
  assign sel_550809 = array_index_550760 == array_index_537088 ? add_550808 : sel_550805;
  assign add_550812 = sel_550809 + 8'h01;
  assign sel_550813 = array_index_550760 == array_index_537094 ? add_550812 : sel_550809;
  assign add_550816 = sel_550813 + 8'h01;
  assign sel_550817 = array_index_550760 == array_index_537100 ? add_550816 : sel_550813;
  assign add_550820 = sel_550817 + 8'h01;
  assign sel_550821 = array_index_550760 == array_index_537106 ? add_550820 : sel_550817;
  assign add_550824 = sel_550821 + 8'h01;
  assign sel_550825 = array_index_550760 == array_index_537112 ? add_550824 : sel_550821;
  assign add_550828 = sel_550825 + 8'h01;
  assign sel_550829 = array_index_550760 == array_index_537118 ? add_550828 : sel_550825;
  assign add_550832 = sel_550829 + 8'h01;
  assign sel_550833 = array_index_550760 == array_index_537124 ? add_550832 : sel_550829;
  assign add_550836 = sel_550833 + 8'h01;
  assign sel_550837 = array_index_550760 == array_index_537130 ? add_550836 : sel_550833;
  assign add_550840 = sel_550837 + 8'h01;
  assign sel_550841 = array_index_550760 == array_index_537136 ? add_550840 : sel_550837;
  assign add_550844 = sel_550841 + 8'h01;
  assign sel_550845 = array_index_550760 == array_index_537142 ? add_550844 : sel_550841;
  assign add_550848 = sel_550845 + 8'h01;
  assign sel_550849 = array_index_550760 == array_index_537148 ? add_550848 : sel_550845;
  assign add_550852 = sel_550849 + 8'h01;
  assign sel_550853 = array_index_550760 == array_index_537154 ? add_550852 : sel_550849;
  assign add_550856 = sel_550853 + 8'h01;
  assign sel_550857 = array_index_550760 == array_index_537160 ? add_550856 : sel_550853;
  assign add_550860 = sel_550857 + 8'h01;
  assign sel_550861 = array_index_550760 == array_index_537166 ? add_550860 : sel_550857;
  assign add_550864 = sel_550861 + 8'h01;
  assign sel_550865 = array_index_550760 == array_index_537172 ? add_550864 : sel_550861;
  assign add_550868 = sel_550865 + 8'h01;
  assign sel_550869 = array_index_550760 == array_index_537178 ? add_550868 : sel_550865;
  assign add_550872 = sel_550869 + 8'h01;
  assign sel_550873 = array_index_550760 == array_index_537184 ? add_550872 : sel_550869;
  assign add_550876 = sel_550873 + 8'h01;
  assign sel_550877 = array_index_550760 == array_index_537190 ? add_550876 : sel_550873;
  assign add_550880 = sel_550877 + 8'h01;
  assign sel_550881 = array_index_550760 == array_index_537196 ? add_550880 : sel_550877;
  assign add_550884 = sel_550881 + 8'h01;
  assign sel_550885 = array_index_550760 == array_index_537202 ? add_550884 : sel_550881;
  assign add_550888 = sel_550885 + 8'h01;
  assign sel_550889 = array_index_550760 == array_index_537208 ? add_550888 : sel_550885;
  assign add_550892 = sel_550889 + 8'h01;
  assign sel_550893 = array_index_550760 == array_index_537214 ? add_550892 : sel_550889;
  assign add_550896 = sel_550893 + 8'h01;
  assign sel_550897 = array_index_550760 == array_index_537220 ? add_550896 : sel_550893;
  assign add_550900 = sel_550897 + 8'h01;
  assign sel_550901 = array_index_550760 == array_index_537226 ? add_550900 : sel_550897;
  assign add_550904 = sel_550901 + 8'h01;
  assign sel_550905 = array_index_550760 == array_index_537232 ? add_550904 : sel_550901;
  assign add_550908 = sel_550905 + 8'h01;
  assign sel_550909 = array_index_550760 == array_index_537238 ? add_550908 : sel_550905;
  assign add_550912 = sel_550909 + 8'h01;
  assign sel_550913 = array_index_550760 == array_index_537244 ? add_550912 : sel_550909;
  assign add_550916 = sel_550913 + 8'h01;
  assign sel_550917 = array_index_550760 == array_index_537250 ? add_550916 : sel_550913;
  assign add_550920 = sel_550917 + 8'h01;
  assign sel_550921 = array_index_550760 == array_index_537256 ? add_550920 : sel_550917;
  assign add_550924 = sel_550921 + 8'h01;
  assign sel_550925 = array_index_550760 == array_index_537262 ? add_550924 : sel_550921;
  assign add_550928 = sel_550925 + 8'h01;
  assign sel_550929 = array_index_550760 == array_index_537268 ? add_550928 : sel_550925;
  assign add_550932 = sel_550929 + 8'h01;
  assign sel_550933 = array_index_550760 == array_index_537274 ? add_550932 : sel_550929;
  assign add_550936 = sel_550933 + 8'h01;
  assign sel_550937 = array_index_550760 == array_index_537280 ? add_550936 : sel_550933;
  assign add_550940 = sel_550937 + 8'h01;
  assign sel_550941 = array_index_550760 == array_index_537286 ? add_550940 : sel_550937;
  assign add_550944 = sel_550941 + 8'h01;
  assign sel_550945 = array_index_550760 == array_index_537292 ? add_550944 : sel_550941;
  assign add_550948 = sel_550945 + 8'h01;
  assign sel_550949 = array_index_550760 == array_index_537298 ? add_550948 : sel_550945;
  assign add_550952 = sel_550949 + 8'h01;
  assign sel_550953 = array_index_550760 == array_index_537304 ? add_550952 : sel_550949;
  assign add_550956 = sel_550953 + 8'h01;
  assign sel_550957 = array_index_550760 == array_index_537310 ? add_550956 : sel_550953;
  assign add_550960 = sel_550957 + 8'h01;
  assign sel_550961 = array_index_550760 == array_index_537316 ? add_550960 : sel_550957;
  assign add_550964 = sel_550961 + 8'h01;
  assign sel_550965 = array_index_550760 == array_index_537322 ? add_550964 : sel_550961;
  assign add_550968 = sel_550965 + 8'h01;
  assign sel_550969 = array_index_550760 == array_index_537328 ? add_550968 : sel_550965;
  assign add_550972 = sel_550969 + 8'h01;
  assign sel_550973 = array_index_550760 == array_index_537334 ? add_550972 : sel_550969;
  assign add_550976 = sel_550973 + 8'h01;
  assign sel_550977 = array_index_550760 == array_index_537340 ? add_550976 : sel_550973;
  assign add_550980 = sel_550977 + 8'h01;
  assign sel_550981 = array_index_550760 == array_index_537346 ? add_550980 : sel_550977;
  assign add_550984 = sel_550981 + 8'h01;
  assign sel_550985 = array_index_550760 == array_index_537352 ? add_550984 : sel_550981;
  assign add_550988 = sel_550985 + 8'h01;
  assign sel_550989 = array_index_550760 == array_index_537358 ? add_550988 : sel_550985;
  assign add_550992 = sel_550989 + 8'h01;
  assign sel_550993 = array_index_550760 == array_index_537364 ? add_550992 : sel_550989;
  assign add_550996 = sel_550993 + 8'h01;
  assign sel_550997 = array_index_550760 == array_index_537370 ? add_550996 : sel_550993;
  assign add_551000 = sel_550997 + 8'h01;
  assign sel_551001 = array_index_550760 == array_index_537376 ? add_551000 : sel_550997;
  assign add_551004 = sel_551001 + 8'h01;
  assign sel_551005 = array_index_550760 == array_index_537382 ? add_551004 : sel_551001;
  assign add_551008 = sel_551005 + 8'h01;
  assign sel_551009 = array_index_550760 == array_index_537388 ? add_551008 : sel_551005;
  assign add_551012 = sel_551009 + 8'h01;
  assign sel_551013 = array_index_550760 == array_index_537394 ? add_551012 : sel_551009;
  assign add_551016 = sel_551013 + 8'h01;
  assign sel_551017 = array_index_550760 == array_index_537400 ? add_551016 : sel_551013;
  assign add_551020 = sel_551017 + 8'h01;
  assign sel_551021 = array_index_550760 == array_index_537406 ? add_551020 : sel_551017;
  assign add_551024 = sel_551021 + 8'h01;
  assign sel_551025 = array_index_550760 == array_index_537412 ? add_551024 : sel_551021;
  assign add_551028 = sel_551025 + 8'h01;
  assign sel_551029 = array_index_550760 == array_index_537418 ? add_551028 : sel_551025;
  assign add_551032 = sel_551029 + 8'h01;
  assign sel_551033 = array_index_550760 == array_index_537424 ? add_551032 : sel_551029;
  assign add_551036 = sel_551033 + 8'h01;
  assign sel_551037 = array_index_550760 == array_index_537430 ? add_551036 : sel_551033;
  assign add_551040 = sel_551037 + 8'h01;
  assign sel_551041 = array_index_550760 == array_index_537436 ? add_551040 : sel_551037;
  assign add_551044 = sel_551041 + 8'h01;
  assign sel_551045 = array_index_550760 == array_index_537442 ? add_551044 : sel_551041;
  assign add_551048 = sel_551045 + 8'h01;
  assign sel_551049 = array_index_550760 == array_index_537448 ? add_551048 : sel_551045;
  assign add_551052 = sel_551049 + 8'h01;
  assign sel_551053 = array_index_550760 == array_index_537454 ? add_551052 : sel_551049;
  assign add_551056 = sel_551053 + 8'h01;
  assign sel_551057 = array_index_550760 == array_index_537460 ? add_551056 : sel_551053;
  assign add_551061 = sel_551057 + 8'h01;
  assign array_index_551062 = set1_unflattened[7'h2e];
  assign sel_551063 = array_index_550760 == array_index_537466 ? add_551061 : sel_551057;
  assign add_551066 = sel_551063 + 8'h01;
  assign sel_551067 = array_index_551062 == array_index_537012 ? add_551066 : sel_551063;
  assign add_551070 = sel_551067 + 8'h01;
  assign sel_551071 = array_index_551062 == array_index_537016 ? add_551070 : sel_551067;
  assign add_551074 = sel_551071 + 8'h01;
  assign sel_551075 = array_index_551062 == array_index_537024 ? add_551074 : sel_551071;
  assign add_551078 = sel_551075 + 8'h01;
  assign sel_551079 = array_index_551062 == array_index_537032 ? add_551078 : sel_551075;
  assign add_551082 = sel_551079 + 8'h01;
  assign sel_551083 = array_index_551062 == array_index_537040 ? add_551082 : sel_551079;
  assign add_551086 = sel_551083 + 8'h01;
  assign sel_551087 = array_index_551062 == array_index_537048 ? add_551086 : sel_551083;
  assign add_551090 = sel_551087 + 8'h01;
  assign sel_551091 = array_index_551062 == array_index_537056 ? add_551090 : sel_551087;
  assign add_551094 = sel_551091 + 8'h01;
  assign sel_551095 = array_index_551062 == array_index_537064 ? add_551094 : sel_551091;
  assign add_551098 = sel_551095 + 8'h01;
  assign sel_551099 = array_index_551062 == array_index_537070 ? add_551098 : sel_551095;
  assign add_551102 = sel_551099 + 8'h01;
  assign sel_551103 = array_index_551062 == array_index_537076 ? add_551102 : sel_551099;
  assign add_551106 = sel_551103 + 8'h01;
  assign sel_551107 = array_index_551062 == array_index_537082 ? add_551106 : sel_551103;
  assign add_551110 = sel_551107 + 8'h01;
  assign sel_551111 = array_index_551062 == array_index_537088 ? add_551110 : sel_551107;
  assign add_551114 = sel_551111 + 8'h01;
  assign sel_551115 = array_index_551062 == array_index_537094 ? add_551114 : sel_551111;
  assign add_551118 = sel_551115 + 8'h01;
  assign sel_551119 = array_index_551062 == array_index_537100 ? add_551118 : sel_551115;
  assign add_551122 = sel_551119 + 8'h01;
  assign sel_551123 = array_index_551062 == array_index_537106 ? add_551122 : sel_551119;
  assign add_551126 = sel_551123 + 8'h01;
  assign sel_551127 = array_index_551062 == array_index_537112 ? add_551126 : sel_551123;
  assign add_551130 = sel_551127 + 8'h01;
  assign sel_551131 = array_index_551062 == array_index_537118 ? add_551130 : sel_551127;
  assign add_551134 = sel_551131 + 8'h01;
  assign sel_551135 = array_index_551062 == array_index_537124 ? add_551134 : sel_551131;
  assign add_551138 = sel_551135 + 8'h01;
  assign sel_551139 = array_index_551062 == array_index_537130 ? add_551138 : sel_551135;
  assign add_551142 = sel_551139 + 8'h01;
  assign sel_551143 = array_index_551062 == array_index_537136 ? add_551142 : sel_551139;
  assign add_551146 = sel_551143 + 8'h01;
  assign sel_551147 = array_index_551062 == array_index_537142 ? add_551146 : sel_551143;
  assign add_551150 = sel_551147 + 8'h01;
  assign sel_551151 = array_index_551062 == array_index_537148 ? add_551150 : sel_551147;
  assign add_551154 = sel_551151 + 8'h01;
  assign sel_551155 = array_index_551062 == array_index_537154 ? add_551154 : sel_551151;
  assign add_551158 = sel_551155 + 8'h01;
  assign sel_551159 = array_index_551062 == array_index_537160 ? add_551158 : sel_551155;
  assign add_551162 = sel_551159 + 8'h01;
  assign sel_551163 = array_index_551062 == array_index_537166 ? add_551162 : sel_551159;
  assign add_551166 = sel_551163 + 8'h01;
  assign sel_551167 = array_index_551062 == array_index_537172 ? add_551166 : sel_551163;
  assign add_551170 = sel_551167 + 8'h01;
  assign sel_551171 = array_index_551062 == array_index_537178 ? add_551170 : sel_551167;
  assign add_551174 = sel_551171 + 8'h01;
  assign sel_551175 = array_index_551062 == array_index_537184 ? add_551174 : sel_551171;
  assign add_551178 = sel_551175 + 8'h01;
  assign sel_551179 = array_index_551062 == array_index_537190 ? add_551178 : sel_551175;
  assign add_551182 = sel_551179 + 8'h01;
  assign sel_551183 = array_index_551062 == array_index_537196 ? add_551182 : sel_551179;
  assign add_551186 = sel_551183 + 8'h01;
  assign sel_551187 = array_index_551062 == array_index_537202 ? add_551186 : sel_551183;
  assign add_551190 = sel_551187 + 8'h01;
  assign sel_551191 = array_index_551062 == array_index_537208 ? add_551190 : sel_551187;
  assign add_551194 = sel_551191 + 8'h01;
  assign sel_551195 = array_index_551062 == array_index_537214 ? add_551194 : sel_551191;
  assign add_551198 = sel_551195 + 8'h01;
  assign sel_551199 = array_index_551062 == array_index_537220 ? add_551198 : sel_551195;
  assign add_551202 = sel_551199 + 8'h01;
  assign sel_551203 = array_index_551062 == array_index_537226 ? add_551202 : sel_551199;
  assign add_551206 = sel_551203 + 8'h01;
  assign sel_551207 = array_index_551062 == array_index_537232 ? add_551206 : sel_551203;
  assign add_551210 = sel_551207 + 8'h01;
  assign sel_551211 = array_index_551062 == array_index_537238 ? add_551210 : sel_551207;
  assign add_551214 = sel_551211 + 8'h01;
  assign sel_551215 = array_index_551062 == array_index_537244 ? add_551214 : sel_551211;
  assign add_551218 = sel_551215 + 8'h01;
  assign sel_551219 = array_index_551062 == array_index_537250 ? add_551218 : sel_551215;
  assign add_551222 = sel_551219 + 8'h01;
  assign sel_551223 = array_index_551062 == array_index_537256 ? add_551222 : sel_551219;
  assign add_551226 = sel_551223 + 8'h01;
  assign sel_551227 = array_index_551062 == array_index_537262 ? add_551226 : sel_551223;
  assign add_551230 = sel_551227 + 8'h01;
  assign sel_551231 = array_index_551062 == array_index_537268 ? add_551230 : sel_551227;
  assign add_551234 = sel_551231 + 8'h01;
  assign sel_551235 = array_index_551062 == array_index_537274 ? add_551234 : sel_551231;
  assign add_551238 = sel_551235 + 8'h01;
  assign sel_551239 = array_index_551062 == array_index_537280 ? add_551238 : sel_551235;
  assign add_551242 = sel_551239 + 8'h01;
  assign sel_551243 = array_index_551062 == array_index_537286 ? add_551242 : sel_551239;
  assign add_551246 = sel_551243 + 8'h01;
  assign sel_551247 = array_index_551062 == array_index_537292 ? add_551246 : sel_551243;
  assign add_551250 = sel_551247 + 8'h01;
  assign sel_551251 = array_index_551062 == array_index_537298 ? add_551250 : sel_551247;
  assign add_551254 = sel_551251 + 8'h01;
  assign sel_551255 = array_index_551062 == array_index_537304 ? add_551254 : sel_551251;
  assign add_551258 = sel_551255 + 8'h01;
  assign sel_551259 = array_index_551062 == array_index_537310 ? add_551258 : sel_551255;
  assign add_551262 = sel_551259 + 8'h01;
  assign sel_551263 = array_index_551062 == array_index_537316 ? add_551262 : sel_551259;
  assign add_551266 = sel_551263 + 8'h01;
  assign sel_551267 = array_index_551062 == array_index_537322 ? add_551266 : sel_551263;
  assign add_551270 = sel_551267 + 8'h01;
  assign sel_551271 = array_index_551062 == array_index_537328 ? add_551270 : sel_551267;
  assign add_551274 = sel_551271 + 8'h01;
  assign sel_551275 = array_index_551062 == array_index_537334 ? add_551274 : sel_551271;
  assign add_551278 = sel_551275 + 8'h01;
  assign sel_551279 = array_index_551062 == array_index_537340 ? add_551278 : sel_551275;
  assign add_551282 = sel_551279 + 8'h01;
  assign sel_551283 = array_index_551062 == array_index_537346 ? add_551282 : sel_551279;
  assign add_551286 = sel_551283 + 8'h01;
  assign sel_551287 = array_index_551062 == array_index_537352 ? add_551286 : sel_551283;
  assign add_551290 = sel_551287 + 8'h01;
  assign sel_551291 = array_index_551062 == array_index_537358 ? add_551290 : sel_551287;
  assign add_551294 = sel_551291 + 8'h01;
  assign sel_551295 = array_index_551062 == array_index_537364 ? add_551294 : sel_551291;
  assign add_551298 = sel_551295 + 8'h01;
  assign sel_551299 = array_index_551062 == array_index_537370 ? add_551298 : sel_551295;
  assign add_551302 = sel_551299 + 8'h01;
  assign sel_551303 = array_index_551062 == array_index_537376 ? add_551302 : sel_551299;
  assign add_551306 = sel_551303 + 8'h01;
  assign sel_551307 = array_index_551062 == array_index_537382 ? add_551306 : sel_551303;
  assign add_551310 = sel_551307 + 8'h01;
  assign sel_551311 = array_index_551062 == array_index_537388 ? add_551310 : sel_551307;
  assign add_551314 = sel_551311 + 8'h01;
  assign sel_551315 = array_index_551062 == array_index_537394 ? add_551314 : sel_551311;
  assign add_551318 = sel_551315 + 8'h01;
  assign sel_551319 = array_index_551062 == array_index_537400 ? add_551318 : sel_551315;
  assign add_551322 = sel_551319 + 8'h01;
  assign sel_551323 = array_index_551062 == array_index_537406 ? add_551322 : sel_551319;
  assign add_551326 = sel_551323 + 8'h01;
  assign sel_551327 = array_index_551062 == array_index_537412 ? add_551326 : sel_551323;
  assign add_551330 = sel_551327 + 8'h01;
  assign sel_551331 = array_index_551062 == array_index_537418 ? add_551330 : sel_551327;
  assign add_551334 = sel_551331 + 8'h01;
  assign sel_551335 = array_index_551062 == array_index_537424 ? add_551334 : sel_551331;
  assign add_551338 = sel_551335 + 8'h01;
  assign sel_551339 = array_index_551062 == array_index_537430 ? add_551338 : sel_551335;
  assign add_551342 = sel_551339 + 8'h01;
  assign sel_551343 = array_index_551062 == array_index_537436 ? add_551342 : sel_551339;
  assign add_551346 = sel_551343 + 8'h01;
  assign sel_551347 = array_index_551062 == array_index_537442 ? add_551346 : sel_551343;
  assign add_551350 = sel_551347 + 8'h01;
  assign sel_551351 = array_index_551062 == array_index_537448 ? add_551350 : sel_551347;
  assign add_551354 = sel_551351 + 8'h01;
  assign sel_551355 = array_index_551062 == array_index_537454 ? add_551354 : sel_551351;
  assign add_551358 = sel_551355 + 8'h01;
  assign sel_551359 = array_index_551062 == array_index_537460 ? add_551358 : sel_551355;
  assign add_551363 = sel_551359 + 8'h01;
  assign array_index_551364 = set1_unflattened[7'h2f];
  assign sel_551365 = array_index_551062 == array_index_537466 ? add_551363 : sel_551359;
  assign add_551368 = sel_551365 + 8'h01;
  assign sel_551369 = array_index_551364 == array_index_537012 ? add_551368 : sel_551365;
  assign add_551372 = sel_551369 + 8'h01;
  assign sel_551373 = array_index_551364 == array_index_537016 ? add_551372 : sel_551369;
  assign add_551376 = sel_551373 + 8'h01;
  assign sel_551377 = array_index_551364 == array_index_537024 ? add_551376 : sel_551373;
  assign add_551380 = sel_551377 + 8'h01;
  assign sel_551381 = array_index_551364 == array_index_537032 ? add_551380 : sel_551377;
  assign add_551384 = sel_551381 + 8'h01;
  assign sel_551385 = array_index_551364 == array_index_537040 ? add_551384 : sel_551381;
  assign add_551388 = sel_551385 + 8'h01;
  assign sel_551389 = array_index_551364 == array_index_537048 ? add_551388 : sel_551385;
  assign add_551392 = sel_551389 + 8'h01;
  assign sel_551393 = array_index_551364 == array_index_537056 ? add_551392 : sel_551389;
  assign add_551396 = sel_551393 + 8'h01;
  assign sel_551397 = array_index_551364 == array_index_537064 ? add_551396 : sel_551393;
  assign add_551400 = sel_551397 + 8'h01;
  assign sel_551401 = array_index_551364 == array_index_537070 ? add_551400 : sel_551397;
  assign add_551404 = sel_551401 + 8'h01;
  assign sel_551405 = array_index_551364 == array_index_537076 ? add_551404 : sel_551401;
  assign add_551408 = sel_551405 + 8'h01;
  assign sel_551409 = array_index_551364 == array_index_537082 ? add_551408 : sel_551405;
  assign add_551412 = sel_551409 + 8'h01;
  assign sel_551413 = array_index_551364 == array_index_537088 ? add_551412 : sel_551409;
  assign add_551416 = sel_551413 + 8'h01;
  assign sel_551417 = array_index_551364 == array_index_537094 ? add_551416 : sel_551413;
  assign add_551420 = sel_551417 + 8'h01;
  assign sel_551421 = array_index_551364 == array_index_537100 ? add_551420 : sel_551417;
  assign add_551424 = sel_551421 + 8'h01;
  assign sel_551425 = array_index_551364 == array_index_537106 ? add_551424 : sel_551421;
  assign add_551428 = sel_551425 + 8'h01;
  assign sel_551429 = array_index_551364 == array_index_537112 ? add_551428 : sel_551425;
  assign add_551432 = sel_551429 + 8'h01;
  assign sel_551433 = array_index_551364 == array_index_537118 ? add_551432 : sel_551429;
  assign add_551436 = sel_551433 + 8'h01;
  assign sel_551437 = array_index_551364 == array_index_537124 ? add_551436 : sel_551433;
  assign add_551440 = sel_551437 + 8'h01;
  assign sel_551441 = array_index_551364 == array_index_537130 ? add_551440 : sel_551437;
  assign add_551444 = sel_551441 + 8'h01;
  assign sel_551445 = array_index_551364 == array_index_537136 ? add_551444 : sel_551441;
  assign add_551448 = sel_551445 + 8'h01;
  assign sel_551449 = array_index_551364 == array_index_537142 ? add_551448 : sel_551445;
  assign add_551452 = sel_551449 + 8'h01;
  assign sel_551453 = array_index_551364 == array_index_537148 ? add_551452 : sel_551449;
  assign add_551456 = sel_551453 + 8'h01;
  assign sel_551457 = array_index_551364 == array_index_537154 ? add_551456 : sel_551453;
  assign add_551460 = sel_551457 + 8'h01;
  assign sel_551461 = array_index_551364 == array_index_537160 ? add_551460 : sel_551457;
  assign add_551464 = sel_551461 + 8'h01;
  assign sel_551465 = array_index_551364 == array_index_537166 ? add_551464 : sel_551461;
  assign add_551468 = sel_551465 + 8'h01;
  assign sel_551469 = array_index_551364 == array_index_537172 ? add_551468 : sel_551465;
  assign add_551472 = sel_551469 + 8'h01;
  assign sel_551473 = array_index_551364 == array_index_537178 ? add_551472 : sel_551469;
  assign add_551476 = sel_551473 + 8'h01;
  assign sel_551477 = array_index_551364 == array_index_537184 ? add_551476 : sel_551473;
  assign add_551480 = sel_551477 + 8'h01;
  assign sel_551481 = array_index_551364 == array_index_537190 ? add_551480 : sel_551477;
  assign add_551484 = sel_551481 + 8'h01;
  assign sel_551485 = array_index_551364 == array_index_537196 ? add_551484 : sel_551481;
  assign add_551488 = sel_551485 + 8'h01;
  assign sel_551489 = array_index_551364 == array_index_537202 ? add_551488 : sel_551485;
  assign add_551492 = sel_551489 + 8'h01;
  assign sel_551493 = array_index_551364 == array_index_537208 ? add_551492 : sel_551489;
  assign add_551496 = sel_551493 + 8'h01;
  assign sel_551497 = array_index_551364 == array_index_537214 ? add_551496 : sel_551493;
  assign add_551500 = sel_551497 + 8'h01;
  assign sel_551501 = array_index_551364 == array_index_537220 ? add_551500 : sel_551497;
  assign add_551504 = sel_551501 + 8'h01;
  assign sel_551505 = array_index_551364 == array_index_537226 ? add_551504 : sel_551501;
  assign add_551508 = sel_551505 + 8'h01;
  assign sel_551509 = array_index_551364 == array_index_537232 ? add_551508 : sel_551505;
  assign add_551512 = sel_551509 + 8'h01;
  assign sel_551513 = array_index_551364 == array_index_537238 ? add_551512 : sel_551509;
  assign add_551516 = sel_551513 + 8'h01;
  assign sel_551517 = array_index_551364 == array_index_537244 ? add_551516 : sel_551513;
  assign add_551520 = sel_551517 + 8'h01;
  assign sel_551521 = array_index_551364 == array_index_537250 ? add_551520 : sel_551517;
  assign add_551524 = sel_551521 + 8'h01;
  assign sel_551525 = array_index_551364 == array_index_537256 ? add_551524 : sel_551521;
  assign add_551528 = sel_551525 + 8'h01;
  assign sel_551529 = array_index_551364 == array_index_537262 ? add_551528 : sel_551525;
  assign add_551532 = sel_551529 + 8'h01;
  assign sel_551533 = array_index_551364 == array_index_537268 ? add_551532 : sel_551529;
  assign add_551536 = sel_551533 + 8'h01;
  assign sel_551537 = array_index_551364 == array_index_537274 ? add_551536 : sel_551533;
  assign add_551540 = sel_551537 + 8'h01;
  assign sel_551541 = array_index_551364 == array_index_537280 ? add_551540 : sel_551537;
  assign add_551544 = sel_551541 + 8'h01;
  assign sel_551545 = array_index_551364 == array_index_537286 ? add_551544 : sel_551541;
  assign add_551548 = sel_551545 + 8'h01;
  assign sel_551549 = array_index_551364 == array_index_537292 ? add_551548 : sel_551545;
  assign add_551552 = sel_551549 + 8'h01;
  assign sel_551553 = array_index_551364 == array_index_537298 ? add_551552 : sel_551549;
  assign add_551556 = sel_551553 + 8'h01;
  assign sel_551557 = array_index_551364 == array_index_537304 ? add_551556 : sel_551553;
  assign add_551560 = sel_551557 + 8'h01;
  assign sel_551561 = array_index_551364 == array_index_537310 ? add_551560 : sel_551557;
  assign add_551564 = sel_551561 + 8'h01;
  assign sel_551565 = array_index_551364 == array_index_537316 ? add_551564 : sel_551561;
  assign add_551568 = sel_551565 + 8'h01;
  assign sel_551569 = array_index_551364 == array_index_537322 ? add_551568 : sel_551565;
  assign add_551572 = sel_551569 + 8'h01;
  assign sel_551573 = array_index_551364 == array_index_537328 ? add_551572 : sel_551569;
  assign add_551576 = sel_551573 + 8'h01;
  assign sel_551577 = array_index_551364 == array_index_537334 ? add_551576 : sel_551573;
  assign add_551580 = sel_551577 + 8'h01;
  assign sel_551581 = array_index_551364 == array_index_537340 ? add_551580 : sel_551577;
  assign add_551584 = sel_551581 + 8'h01;
  assign sel_551585 = array_index_551364 == array_index_537346 ? add_551584 : sel_551581;
  assign add_551588 = sel_551585 + 8'h01;
  assign sel_551589 = array_index_551364 == array_index_537352 ? add_551588 : sel_551585;
  assign add_551592 = sel_551589 + 8'h01;
  assign sel_551593 = array_index_551364 == array_index_537358 ? add_551592 : sel_551589;
  assign add_551596 = sel_551593 + 8'h01;
  assign sel_551597 = array_index_551364 == array_index_537364 ? add_551596 : sel_551593;
  assign add_551600 = sel_551597 + 8'h01;
  assign sel_551601 = array_index_551364 == array_index_537370 ? add_551600 : sel_551597;
  assign add_551604 = sel_551601 + 8'h01;
  assign sel_551605 = array_index_551364 == array_index_537376 ? add_551604 : sel_551601;
  assign add_551608 = sel_551605 + 8'h01;
  assign sel_551609 = array_index_551364 == array_index_537382 ? add_551608 : sel_551605;
  assign add_551612 = sel_551609 + 8'h01;
  assign sel_551613 = array_index_551364 == array_index_537388 ? add_551612 : sel_551609;
  assign add_551616 = sel_551613 + 8'h01;
  assign sel_551617 = array_index_551364 == array_index_537394 ? add_551616 : sel_551613;
  assign add_551620 = sel_551617 + 8'h01;
  assign sel_551621 = array_index_551364 == array_index_537400 ? add_551620 : sel_551617;
  assign add_551624 = sel_551621 + 8'h01;
  assign sel_551625 = array_index_551364 == array_index_537406 ? add_551624 : sel_551621;
  assign add_551628 = sel_551625 + 8'h01;
  assign sel_551629 = array_index_551364 == array_index_537412 ? add_551628 : sel_551625;
  assign add_551632 = sel_551629 + 8'h01;
  assign sel_551633 = array_index_551364 == array_index_537418 ? add_551632 : sel_551629;
  assign add_551636 = sel_551633 + 8'h01;
  assign sel_551637 = array_index_551364 == array_index_537424 ? add_551636 : sel_551633;
  assign add_551640 = sel_551637 + 8'h01;
  assign sel_551641 = array_index_551364 == array_index_537430 ? add_551640 : sel_551637;
  assign add_551644 = sel_551641 + 8'h01;
  assign sel_551645 = array_index_551364 == array_index_537436 ? add_551644 : sel_551641;
  assign add_551648 = sel_551645 + 8'h01;
  assign sel_551649 = array_index_551364 == array_index_537442 ? add_551648 : sel_551645;
  assign add_551652 = sel_551649 + 8'h01;
  assign sel_551653 = array_index_551364 == array_index_537448 ? add_551652 : sel_551649;
  assign add_551656 = sel_551653 + 8'h01;
  assign sel_551657 = array_index_551364 == array_index_537454 ? add_551656 : sel_551653;
  assign add_551660 = sel_551657 + 8'h01;
  assign sel_551661 = array_index_551364 == array_index_537460 ? add_551660 : sel_551657;
  assign add_551665 = sel_551661 + 8'h01;
  assign array_index_551666 = set1_unflattened[7'h30];
  assign sel_551667 = array_index_551364 == array_index_537466 ? add_551665 : sel_551661;
  assign add_551670 = sel_551667 + 8'h01;
  assign sel_551671 = array_index_551666 == array_index_537012 ? add_551670 : sel_551667;
  assign add_551674 = sel_551671 + 8'h01;
  assign sel_551675 = array_index_551666 == array_index_537016 ? add_551674 : sel_551671;
  assign add_551678 = sel_551675 + 8'h01;
  assign sel_551679 = array_index_551666 == array_index_537024 ? add_551678 : sel_551675;
  assign add_551682 = sel_551679 + 8'h01;
  assign sel_551683 = array_index_551666 == array_index_537032 ? add_551682 : sel_551679;
  assign add_551686 = sel_551683 + 8'h01;
  assign sel_551687 = array_index_551666 == array_index_537040 ? add_551686 : sel_551683;
  assign add_551690 = sel_551687 + 8'h01;
  assign sel_551691 = array_index_551666 == array_index_537048 ? add_551690 : sel_551687;
  assign add_551694 = sel_551691 + 8'h01;
  assign sel_551695 = array_index_551666 == array_index_537056 ? add_551694 : sel_551691;
  assign add_551698 = sel_551695 + 8'h01;
  assign sel_551699 = array_index_551666 == array_index_537064 ? add_551698 : sel_551695;
  assign add_551702 = sel_551699 + 8'h01;
  assign sel_551703 = array_index_551666 == array_index_537070 ? add_551702 : sel_551699;
  assign add_551706 = sel_551703 + 8'h01;
  assign sel_551707 = array_index_551666 == array_index_537076 ? add_551706 : sel_551703;
  assign add_551710 = sel_551707 + 8'h01;
  assign sel_551711 = array_index_551666 == array_index_537082 ? add_551710 : sel_551707;
  assign add_551714 = sel_551711 + 8'h01;
  assign sel_551715 = array_index_551666 == array_index_537088 ? add_551714 : sel_551711;
  assign add_551718 = sel_551715 + 8'h01;
  assign sel_551719 = array_index_551666 == array_index_537094 ? add_551718 : sel_551715;
  assign add_551722 = sel_551719 + 8'h01;
  assign sel_551723 = array_index_551666 == array_index_537100 ? add_551722 : sel_551719;
  assign add_551726 = sel_551723 + 8'h01;
  assign sel_551727 = array_index_551666 == array_index_537106 ? add_551726 : sel_551723;
  assign add_551730 = sel_551727 + 8'h01;
  assign sel_551731 = array_index_551666 == array_index_537112 ? add_551730 : sel_551727;
  assign add_551734 = sel_551731 + 8'h01;
  assign sel_551735 = array_index_551666 == array_index_537118 ? add_551734 : sel_551731;
  assign add_551738 = sel_551735 + 8'h01;
  assign sel_551739 = array_index_551666 == array_index_537124 ? add_551738 : sel_551735;
  assign add_551742 = sel_551739 + 8'h01;
  assign sel_551743 = array_index_551666 == array_index_537130 ? add_551742 : sel_551739;
  assign add_551746 = sel_551743 + 8'h01;
  assign sel_551747 = array_index_551666 == array_index_537136 ? add_551746 : sel_551743;
  assign add_551750 = sel_551747 + 8'h01;
  assign sel_551751 = array_index_551666 == array_index_537142 ? add_551750 : sel_551747;
  assign add_551754 = sel_551751 + 8'h01;
  assign sel_551755 = array_index_551666 == array_index_537148 ? add_551754 : sel_551751;
  assign add_551758 = sel_551755 + 8'h01;
  assign sel_551759 = array_index_551666 == array_index_537154 ? add_551758 : sel_551755;
  assign add_551762 = sel_551759 + 8'h01;
  assign sel_551763 = array_index_551666 == array_index_537160 ? add_551762 : sel_551759;
  assign add_551766 = sel_551763 + 8'h01;
  assign sel_551767 = array_index_551666 == array_index_537166 ? add_551766 : sel_551763;
  assign add_551770 = sel_551767 + 8'h01;
  assign sel_551771 = array_index_551666 == array_index_537172 ? add_551770 : sel_551767;
  assign add_551774 = sel_551771 + 8'h01;
  assign sel_551775 = array_index_551666 == array_index_537178 ? add_551774 : sel_551771;
  assign add_551778 = sel_551775 + 8'h01;
  assign sel_551779 = array_index_551666 == array_index_537184 ? add_551778 : sel_551775;
  assign add_551782 = sel_551779 + 8'h01;
  assign sel_551783 = array_index_551666 == array_index_537190 ? add_551782 : sel_551779;
  assign add_551786 = sel_551783 + 8'h01;
  assign sel_551787 = array_index_551666 == array_index_537196 ? add_551786 : sel_551783;
  assign add_551790 = sel_551787 + 8'h01;
  assign sel_551791 = array_index_551666 == array_index_537202 ? add_551790 : sel_551787;
  assign add_551794 = sel_551791 + 8'h01;
  assign sel_551795 = array_index_551666 == array_index_537208 ? add_551794 : sel_551791;
  assign add_551798 = sel_551795 + 8'h01;
  assign sel_551799 = array_index_551666 == array_index_537214 ? add_551798 : sel_551795;
  assign add_551802 = sel_551799 + 8'h01;
  assign sel_551803 = array_index_551666 == array_index_537220 ? add_551802 : sel_551799;
  assign add_551806 = sel_551803 + 8'h01;
  assign sel_551807 = array_index_551666 == array_index_537226 ? add_551806 : sel_551803;
  assign add_551810 = sel_551807 + 8'h01;
  assign sel_551811 = array_index_551666 == array_index_537232 ? add_551810 : sel_551807;
  assign add_551814 = sel_551811 + 8'h01;
  assign sel_551815 = array_index_551666 == array_index_537238 ? add_551814 : sel_551811;
  assign add_551818 = sel_551815 + 8'h01;
  assign sel_551819 = array_index_551666 == array_index_537244 ? add_551818 : sel_551815;
  assign add_551822 = sel_551819 + 8'h01;
  assign sel_551823 = array_index_551666 == array_index_537250 ? add_551822 : sel_551819;
  assign add_551826 = sel_551823 + 8'h01;
  assign sel_551827 = array_index_551666 == array_index_537256 ? add_551826 : sel_551823;
  assign add_551830 = sel_551827 + 8'h01;
  assign sel_551831 = array_index_551666 == array_index_537262 ? add_551830 : sel_551827;
  assign add_551834 = sel_551831 + 8'h01;
  assign sel_551835 = array_index_551666 == array_index_537268 ? add_551834 : sel_551831;
  assign add_551838 = sel_551835 + 8'h01;
  assign sel_551839 = array_index_551666 == array_index_537274 ? add_551838 : sel_551835;
  assign add_551842 = sel_551839 + 8'h01;
  assign sel_551843 = array_index_551666 == array_index_537280 ? add_551842 : sel_551839;
  assign add_551846 = sel_551843 + 8'h01;
  assign sel_551847 = array_index_551666 == array_index_537286 ? add_551846 : sel_551843;
  assign add_551850 = sel_551847 + 8'h01;
  assign sel_551851 = array_index_551666 == array_index_537292 ? add_551850 : sel_551847;
  assign add_551854 = sel_551851 + 8'h01;
  assign sel_551855 = array_index_551666 == array_index_537298 ? add_551854 : sel_551851;
  assign add_551858 = sel_551855 + 8'h01;
  assign sel_551859 = array_index_551666 == array_index_537304 ? add_551858 : sel_551855;
  assign add_551862 = sel_551859 + 8'h01;
  assign sel_551863 = array_index_551666 == array_index_537310 ? add_551862 : sel_551859;
  assign add_551866 = sel_551863 + 8'h01;
  assign sel_551867 = array_index_551666 == array_index_537316 ? add_551866 : sel_551863;
  assign add_551870 = sel_551867 + 8'h01;
  assign sel_551871 = array_index_551666 == array_index_537322 ? add_551870 : sel_551867;
  assign add_551874 = sel_551871 + 8'h01;
  assign sel_551875 = array_index_551666 == array_index_537328 ? add_551874 : sel_551871;
  assign add_551878 = sel_551875 + 8'h01;
  assign sel_551879 = array_index_551666 == array_index_537334 ? add_551878 : sel_551875;
  assign add_551882 = sel_551879 + 8'h01;
  assign sel_551883 = array_index_551666 == array_index_537340 ? add_551882 : sel_551879;
  assign add_551886 = sel_551883 + 8'h01;
  assign sel_551887 = array_index_551666 == array_index_537346 ? add_551886 : sel_551883;
  assign add_551890 = sel_551887 + 8'h01;
  assign sel_551891 = array_index_551666 == array_index_537352 ? add_551890 : sel_551887;
  assign add_551894 = sel_551891 + 8'h01;
  assign sel_551895 = array_index_551666 == array_index_537358 ? add_551894 : sel_551891;
  assign add_551898 = sel_551895 + 8'h01;
  assign sel_551899 = array_index_551666 == array_index_537364 ? add_551898 : sel_551895;
  assign add_551902 = sel_551899 + 8'h01;
  assign sel_551903 = array_index_551666 == array_index_537370 ? add_551902 : sel_551899;
  assign add_551906 = sel_551903 + 8'h01;
  assign sel_551907 = array_index_551666 == array_index_537376 ? add_551906 : sel_551903;
  assign add_551910 = sel_551907 + 8'h01;
  assign sel_551911 = array_index_551666 == array_index_537382 ? add_551910 : sel_551907;
  assign add_551914 = sel_551911 + 8'h01;
  assign sel_551915 = array_index_551666 == array_index_537388 ? add_551914 : sel_551911;
  assign add_551918 = sel_551915 + 8'h01;
  assign sel_551919 = array_index_551666 == array_index_537394 ? add_551918 : sel_551915;
  assign add_551922 = sel_551919 + 8'h01;
  assign sel_551923 = array_index_551666 == array_index_537400 ? add_551922 : sel_551919;
  assign add_551926 = sel_551923 + 8'h01;
  assign sel_551927 = array_index_551666 == array_index_537406 ? add_551926 : sel_551923;
  assign add_551930 = sel_551927 + 8'h01;
  assign sel_551931 = array_index_551666 == array_index_537412 ? add_551930 : sel_551927;
  assign add_551934 = sel_551931 + 8'h01;
  assign sel_551935 = array_index_551666 == array_index_537418 ? add_551934 : sel_551931;
  assign add_551938 = sel_551935 + 8'h01;
  assign sel_551939 = array_index_551666 == array_index_537424 ? add_551938 : sel_551935;
  assign add_551942 = sel_551939 + 8'h01;
  assign sel_551943 = array_index_551666 == array_index_537430 ? add_551942 : sel_551939;
  assign add_551946 = sel_551943 + 8'h01;
  assign sel_551947 = array_index_551666 == array_index_537436 ? add_551946 : sel_551943;
  assign add_551950 = sel_551947 + 8'h01;
  assign sel_551951 = array_index_551666 == array_index_537442 ? add_551950 : sel_551947;
  assign add_551954 = sel_551951 + 8'h01;
  assign sel_551955 = array_index_551666 == array_index_537448 ? add_551954 : sel_551951;
  assign add_551958 = sel_551955 + 8'h01;
  assign sel_551959 = array_index_551666 == array_index_537454 ? add_551958 : sel_551955;
  assign add_551962 = sel_551959 + 8'h01;
  assign sel_551963 = array_index_551666 == array_index_537460 ? add_551962 : sel_551959;
  assign add_551967 = sel_551963 + 8'h01;
  assign array_index_551968 = set1_unflattened[7'h31];
  assign sel_551969 = array_index_551666 == array_index_537466 ? add_551967 : sel_551963;
  assign add_551972 = sel_551969 + 8'h01;
  assign sel_551973 = array_index_551968 == array_index_537012 ? add_551972 : sel_551969;
  assign add_551976 = sel_551973 + 8'h01;
  assign sel_551977 = array_index_551968 == array_index_537016 ? add_551976 : sel_551973;
  assign add_551980 = sel_551977 + 8'h01;
  assign sel_551981 = array_index_551968 == array_index_537024 ? add_551980 : sel_551977;
  assign add_551984 = sel_551981 + 8'h01;
  assign sel_551985 = array_index_551968 == array_index_537032 ? add_551984 : sel_551981;
  assign add_551988 = sel_551985 + 8'h01;
  assign sel_551989 = array_index_551968 == array_index_537040 ? add_551988 : sel_551985;
  assign add_551992 = sel_551989 + 8'h01;
  assign sel_551993 = array_index_551968 == array_index_537048 ? add_551992 : sel_551989;
  assign add_551996 = sel_551993 + 8'h01;
  assign sel_551997 = array_index_551968 == array_index_537056 ? add_551996 : sel_551993;
  assign add_552000 = sel_551997 + 8'h01;
  assign sel_552001 = array_index_551968 == array_index_537064 ? add_552000 : sel_551997;
  assign add_552004 = sel_552001 + 8'h01;
  assign sel_552005 = array_index_551968 == array_index_537070 ? add_552004 : sel_552001;
  assign add_552008 = sel_552005 + 8'h01;
  assign sel_552009 = array_index_551968 == array_index_537076 ? add_552008 : sel_552005;
  assign add_552012 = sel_552009 + 8'h01;
  assign sel_552013 = array_index_551968 == array_index_537082 ? add_552012 : sel_552009;
  assign add_552016 = sel_552013 + 8'h01;
  assign sel_552017 = array_index_551968 == array_index_537088 ? add_552016 : sel_552013;
  assign add_552020 = sel_552017 + 8'h01;
  assign sel_552021 = array_index_551968 == array_index_537094 ? add_552020 : sel_552017;
  assign add_552024 = sel_552021 + 8'h01;
  assign sel_552025 = array_index_551968 == array_index_537100 ? add_552024 : sel_552021;
  assign add_552028 = sel_552025 + 8'h01;
  assign sel_552029 = array_index_551968 == array_index_537106 ? add_552028 : sel_552025;
  assign add_552032 = sel_552029 + 8'h01;
  assign sel_552033 = array_index_551968 == array_index_537112 ? add_552032 : sel_552029;
  assign add_552036 = sel_552033 + 8'h01;
  assign sel_552037 = array_index_551968 == array_index_537118 ? add_552036 : sel_552033;
  assign add_552040 = sel_552037 + 8'h01;
  assign sel_552041 = array_index_551968 == array_index_537124 ? add_552040 : sel_552037;
  assign add_552044 = sel_552041 + 8'h01;
  assign sel_552045 = array_index_551968 == array_index_537130 ? add_552044 : sel_552041;
  assign add_552048 = sel_552045 + 8'h01;
  assign sel_552049 = array_index_551968 == array_index_537136 ? add_552048 : sel_552045;
  assign add_552052 = sel_552049 + 8'h01;
  assign sel_552053 = array_index_551968 == array_index_537142 ? add_552052 : sel_552049;
  assign add_552056 = sel_552053 + 8'h01;
  assign sel_552057 = array_index_551968 == array_index_537148 ? add_552056 : sel_552053;
  assign add_552060 = sel_552057 + 8'h01;
  assign sel_552061 = array_index_551968 == array_index_537154 ? add_552060 : sel_552057;
  assign add_552064 = sel_552061 + 8'h01;
  assign sel_552065 = array_index_551968 == array_index_537160 ? add_552064 : sel_552061;
  assign add_552068 = sel_552065 + 8'h01;
  assign sel_552069 = array_index_551968 == array_index_537166 ? add_552068 : sel_552065;
  assign add_552072 = sel_552069 + 8'h01;
  assign sel_552073 = array_index_551968 == array_index_537172 ? add_552072 : sel_552069;
  assign add_552076 = sel_552073 + 8'h01;
  assign sel_552077 = array_index_551968 == array_index_537178 ? add_552076 : sel_552073;
  assign add_552080 = sel_552077 + 8'h01;
  assign sel_552081 = array_index_551968 == array_index_537184 ? add_552080 : sel_552077;
  assign add_552084 = sel_552081 + 8'h01;
  assign sel_552085 = array_index_551968 == array_index_537190 ? add_552084 : sel_552081;
  assign add_552088 = sel_552085 + 8'h01;
  assign sel_552089 = array_index_551968 == array_index_537196 ? add_552088 : sel_552085;
  assign add_552092 = sel_552089 + 8'h01;
  assign sel_552093 = array_index_551968 == array_index_537202 ? add_552092 : sel_552089;
  assign add_552096 = sel_552093 + 8'h01;
  assign sel_552097 = array_index_551968 == array_index_537208 ? add_552096 : sel_552093;
  assign add_552100 = sel_552097 + 8'h01;
  assign sel_552101 = array_index_551968 == array_index_537214 ? add_552100 : sel_552097;
  assign add_552104 = sel_552101 + 8'h01;
  assign sel_552105 = array_index_551968 == array_index_537220 ? add_552104 : sel_552101;
  assign add_552108 = sel_552105 + 8'h01;
  assign sel_552109 = array_index_551968 == array_index_537226 ? add_552108 : sel_552105;
  assign add_552112 = sel_552109 + 8'h01;
  assign sel_552113 = array_index_551968 == array_index_537232 ? add_552112 : sel_552109;
  assign add_552116 = sel_552113 + 8'h01;
  assign sel_552117 = array_index_551968 == array_index_537238 ? add_552116 : sel_552113;
  assign add_552120 = sel_552117 + 8'h01;
  assign sel_552121 = array_index_551968 == array_index_537244 ? add_552120 : sel_552117;
  assign add_552124 = sel_552121 + 8'h01;
  assign sel_552125 = array_index_551968 == array_index_537250 ? add_552124 : sel_552121;
  assign add_552128 = sel_552125 + 8'h01;
  assign sel_552129 = array_index_551968 == array_index_537256 ? add_552128 : sel_552125;
  assign add_552132 = sel_552129 + 8'h01;
  assign sel_552133 = array_index_551968 == array_index_537262 ? add_552132 : sel_552129;
  assign add_552136 = sel_552133 + 8'h01;
  assign sel_552137 = array_index_551968 == array_index_537268 ? add_552136 : sel_552133;
  assign add_552140 = sel_552137 + 8'h01;
  assign sel_552141 = array_index_551968 == array_index_537274 ? add_552140 : sel_552137;
  assign add_552144 = sel_552141 + 8'h01;
  assign sel_552145 = array_index_551968 == array_index_537280 ? add_552144 : sel_552141;
  assign add_552148 = sel_552145 + 8'h01;
  assign sel_552149 = array_index_551968 == array_index_537286 ? add_552148 : sel_552145;
  assign add_552152 = sel_552149 + 8'h01;
  assign sel_552153 = array_index_551968 == array_index_537292 ? add_552152 : sel_552149;
  assign add_552156 = sel_552153 + 8'h01;
  assign sel_552157 = array_index_551968 == array_index_537298 ? add_552156 : sel_552153;
  assign add_552160 = sel_552157 + 8'h01;
  assign sel_552161 = array_index_551968 == array_index_537304 ? add_552160 : sel_552157;
  assign add_552164 = sel_552161 + 8'h01;
  assign sel_552165 = array_index_551968 == array_index_537310 ? add_552164 : sel_552161;
  assign add_552168 = sel_552165 + 8'h01;
  assign sel_552169 = array_index_551968 == array_index_537316 ? add_552168 : sel_552165;
  assign add_552172 = sel_552169 + 8'h01;
  assign sel_552173 = array_index_551968 == array_index_537322 ? add_552172 : sel_552169;
  assign add_552176 = sel_552173 + 8'h01;
  assign sel_552177 = array_index_551968 == array_index_537328 ? add_552176 : sel_552173;
  assign add_552180 = sel_552177 + 8'h01;
  assign sel_552181 = array_index_551968 == array_index_537334 ? add_552180 : sel_552177;
  assign add_552184 = sel_552181 + 8'h01;
  assign sel_552185 = array_index_551968 == array_index_537340 ? add_552184 : sel_552181;
  assign add_552188 = sel_552185 + 8'h01;
  assign sel_552189 = array_index_551968 == array_index_537346 ? add_552188 : sel_552185;
  assign add_552192 = sel_552189 + 8'h01;
  assign sel_552193 = array_index_551968 == array_index_537352 ? add_552192 : sel_552189;
  assign add_552196 = sel_552193 + 8'h01;
  assign sel_552197 = array_index_551968 == array_index_537358 ? add_552196 : sel_552193;
  assign add_552200 = sel_552197 + 8'h01;
  assign sel_552201 = array_index_551968 == array_index_537364 ? add_552200 : sel_552197;
  assign add_552204 = sel_552201 + 8'h01;
  assign sel_552205 = array_index_551968 == array_index_537370 ? add_552204 : sel_552201;
  assign add_552208 = sel_552205 + 8'h01;
  assign sel_552209 = array_index_551968 == array_index_537376 ? add_552208 : sel_552205;
  assign add_552212 = sel_552209 + 8'h01;
  assign sel_552213 = array_index_551968 == array_index_537382 ? add_552212 : sel_552209;
  assign add_552216 = sel_552213 + 8'h01;
  assign sel_552217 = array_index_551968 == array_index_537388 ? add_552216 : sel_552213;
  assign add_552220 = sel_552217 + 8'h01;
  assign sel_552221 = array_index_551968 == array_index_537394 ? add_552220 : sel_552217;
  assign add_552224 = sel_552221 + 8'h01;
  assign sel_552225 = array_index_551968 == array_index_537400 ? add_552224 : sel_552221;
  assign add_552228 = sel_552225 + 8'h01;
  assign sel_552229 = array_index_551968 == array_index_537406 ? add_552228 : sel_552225;
  assign add_552232 = sel_552229 + 8'h01;
  assign sel_552233 = array_index_551968 == array_index_537412 ? add_552232 : sel_552229;
  assign add_552236 = sel_552233 + 8'h01;
  assign sel_552237 = array_index_551968 == array_index_537418 ? add_552236 : sel_552233;
  assign add_552240 = sel_552237 + 8'h01;
  assign sel_552241 = array_index_551968 == array_index_537424 ? add_552240 : sel_552237;
  assign add_552244 = sel_552241 + 8'h01;
  assign sel_552245 = array_index_551968 == array_index_537430 ? add_552244 : sel_552241;
  assign add_552248 = sel_552245 + 8'h01;
  assign sel_552249 = array_index_551968 == array_index_537436 ? add_552248 : sel_552245;
  assign add_552252 = sel_552249 + 8'h01;
  assign sel_552253 = array_index_551968 == array_index_537442 ? add_552252 : sel_552249;
  assign add_552256 = sel_552253 + 8'h01;
  assign sel_552257 = array_index_551968 == array_index_537448 ? add_552256 : sel_552253;
  assign add_552260 = sel_552257 + 8'h01;
  assign sel_552261 = array_index_551968 == array_index_537454 ? add_552260 : sel_552257;
  assign add_552264 = sel_552261 + 8'h01;
  assign sel_552265 = array_index_551968 == array_index_537460 ? add_552264 : sel_552261;
  assign add_552269 = sel_552265 + 8'h01;
  assign array_index_552270 = set1_unflattened[7'h32];
  assign sel_552271 = array_index_551968 == array_index_537466 ? add_552269 : sel_552265;
  assign add_552274 = sel_552271 + 8'h01;
  assign sel_552275 = array_index_552270 == array_index_537012 ? add_552274 : sel_552271;
  assign add_552278 = sel_552275 + 8'h01;
  assign sel_552279 = array_index_552270 == array_index_537016 ? add_552278 : sel_552275;
  assign add_552282 = sel_552279 + 8'h01;
  assign sel_552283 = array_index_552270 == array_index_537024 ? add_552282 : sel_552279;
  assign add_552286 = sel_552283 + 8'h01;
  assign sel_552287 = array_index_552270 == array_index_537032 ? add_552286 : sel_552283;
  assign add_552290 = sel_552287 + 8'h01;
  assign sel_552291 = array_index_552270 == array_index_537040 ? add_552290 : sel_552287;
  assign add_552294 = sel_552291 + 8'h01;
  assign sel_552295 = array_index_552270 == array_index_537048 ? add_552294 : sel_552291;
  assign add_552298 = sel_552295 + 8'h01;
  assign sel_552299 = array_index_552270 == array_index_537056 ? add_552298 : sel_552295;
  assign add_552302 = sel_552299 + 8'h01;
  assign sel_552303 = array_index_552270 == array_index_537064 ? add_552302 : sel_552299;
  assign add_552306 = sel_552303 + 8'h01;
  assign sel_552307 = array_index_552270 == array_index_537070 ? add_552306 : sel_552303;
  assign add_552310 = sel_552307 + 8'h01;
  assign sel_552311 = array_index_552270 == array_index_537076 ? add_552310 : sel_552307;
  assign add_552314 = sel_552311 + 8'h01;
  assign sel_552315 = array_index_552270 == array_index_537082 ? add_552314 : sel_552311;
  assign add_552318 = sel_552315 + 8'h01;
  assign sel_552319 = array_index_552270 == array_index_537088 ? add_552318 : sel_552315;
  assign add_552322 = sel_552319 + 8'h01;
  assign sel_552323 = array_index_552270 == array_index_537094 ? add_552322 : sel_552319;
  assign add_552326 = sel_552323 + 8'h01;
  assign sel_552327 = array_index_552270 == array_index_537100 ? add_552326 : sel_552323;
  assign add_552330 = sel_552327 + 8'h01;
  assign sel_552331 = array_index_552270 == array_index_537106 ? add_552330 : sel_552327;
  assign add_552334 = sel_552331 + 8'h01;
  assign sel_552335 = array_index_552270 == array_index_537112 ? add_552334 : sel_552331;
  assign add_552338 = sel_552335 + 8'h01;
  assign sel_552339 = array_index_552270 == array_index_537118 ? add_552338 : sel_552335;
  assign add_552342 = sel_552339 + 8'h01;
  assign sel_552343 = array_index_552270 == array_index_537124 ? add_552342 : sel_552339;
  assign add_552346 = sel_552343 + 8'h01;
  assign sel_552347 = array_index_552270 == array_index_537130 ? add_552346 : sel_552343;
  assign add_552350 = sel_552347 + 8'h01;
  assign sel_552351 = array_index_552270 == array_index_537136 ? add_552350 : sel_552347;
  assign add_552354 = sel_552351 + 8'h01;
  assign sel_552355 = array_index_552270 == array_index_537142 ? add_552354 : sel_552351;
  assign add_552358 = sel_552355 + 8'h01;
  assign sel_552359 = array_index_552270 == array_index_537148 ? add_552358 : sel_552355;
  assign add_552362 = sel_552359 + 8'h01;
  assign sel_552363 = array_index_552270 == array_index_537154 ? add_552362 : sel_552359;
  assign add_552366 = sel_552363 + 8'h01;
  assign sel_552367 = array_index_552270 == array_index_537160 ? add_552366 : sel_552363;
  assign add_552370 = sel_552367 + 8'h01;
  assign sel_552371 = array_index_552270 == array_index_537166 ? add_552370 : sel_552367;
  assign add_552374 = sel_552371 + 8'h01;
  assign sel_552375 = array_index_552270 == array_index_537172 ? add_552374 : sel_552371;
  assign add_552378 = sel_552375 + 8'h01;
  assign sel_552379 = array_index_552270 == array_index_537178 ? add_552378 : sel_552375;
  assign add_552382 = sel_552379 + 8'h01;
  assign sel_552383 = array_index_552270 == array_index_537184 ? add_552382 : sel_552379;
  assign add_552386 = sel_552383 + 8'h01;
  assign sel_552387 = array_index_552270 == array_index_537190 ? add_552386 : sel_552383;
  assign add_552390 = sel_552387 + 8'h01;
  assign sel_552391 = array_index_552270 == array_index_537196 ? add_552390 : sel_552387;
  assign add_552394 = sel_552391 + 8'h01;
  assign sel_552395 = array_index_552270 == array_index_537202 ? add_552394 : sel_552391;
  assign add_552398 = sel_552395 + 8'h01;
  assign sel_552399 = array_index_552270 == array_index_537208 ? add_552398 : sel_552395;
  assign add_552402 = sel_552399 + 8'h01;
  assign sel_552403 = array_index_552270 == array_index_537214 ? add_552402 : sel_552399;
  assign add_552406 = sel_552403 + 8'h01;
  assign sel_552407 = array_index_552270 == array_index_537220 ? add_552406 : sel_552403;
  assign add_552410 = sel_552407 + 8'h01;
  assign sel_552411 = array_index_552270 == array_index_537226 ? add_552410 : sel_552407;
  assign add_552414 = sel_552411 + 8'h01;
  assign sel_552415 = array_index_552270 == array_index_537232 ? add_552414 : sel_552411;
  assign add_552418 = sel_552415 + 8'h01;
  assign sel_552419 = array_index_552270 == array_index_537238 ? add_552418 : sel_552415;
  assign add_552422 = sel_552419 + 8'h01;
  assign sel_552423 = array_index_552270 == array_index_537244 ? add_552422 : sel_552419;
  assign add_552426 = sel_552423 + 8'h01;
  assign sel_552427 = array_index_552270 == array_index_537250 ? add_552426 : sel_552423;
  assign add_552430 = sel_552427 + 8'h01;
  assign sel_552431 = array_index_552270 == array_index_537256 ? add_552430 : sel_552427;
  assign add_552434 = sel_552431 + 8'h01;
  assign sel_552435 = array_index_552270 == array_index_537262 ? add_552434 : sel_552431;
  assign add_552438 = sel_552435 + 8'h01;
  assign sel_552439 = array_index_552270 == array_index_537268 ? add_552438 : sel_552435;
  assign add_552442 = sel_552439 + 8'h01;
  assign sel_552443 = array_index_552270 == array_index_537274 ? add_552442 : sel_552439;
  assign add_552446 = sel_552443 + 8'h01;
  assign sel_552447 = array_index_552270 == array_index_537280 ? add_552446 : sel_552443;
  assign add_552450 = sel_552447 + 8'h01;
  assign sel_552451 = array_index_552270 == array_index_537286 ? add_552450 : sel_552447;
  assign add_552454 = sel_552451 + 8'h01;
  assign sel_552455 = array_index_552270 == array_index_537292 ? add_552454 : sel_552451;
  assign add_552458 = sel_552455 + 8'h01;
  assign sel_552459 = array_index_552270 == array_index_537298 ? add_552458 : sel_552455;
  assign add_552462 = sel_552459 + 8'h01;
  assign sel_552463 = array_index_552270 == array_index_537304 ? add_552462 : sel_552459;
  assign add_552466 = sel_552463 + 8'h01;
  assign sel_552467 = array_index_552270 == array_index_537310 ? add_552466 : sel_552463;
  assign add_552470 = sel_552467 + 8'h01;
  assign sel_552471 = array_index_552270 == array_index_537316 ? add_552470 : sel_552467;
  assign add_552474 = sel_552471 + 8'h01;
  assign sel_552475 = array_index_552270 == array_index_537322 ? add_552474 : sel_552471;
  assign add_552478 = sel_552475 + 8'h01;
  assign sel_552479 = array_index_552270 == array_index_537328 ? add_552478 : sel_552475;
  assign add_552482 = sel_552479 + 8'h01;
  assign sel_552483 = array_index_552270 == array_index_537334 ? add_552482 : sel_552479;
  assign add_552486 = sel_552483 + 8'h01;
  assign sel_552487 = array_index_552270 == array_index_537340 ? add_552486 : sel_552483;
  assign add_552490 = sel_552487 + 8'h01;
  assign sel_552491 = array_index_552270 == array_index_537346 ? add_552490 : sel_552487;
  assign add_552494 = sel_552491 + 8'h01;
  assign sel_552495 = array_index_552270 == array_index_537352 ? add_552494 : sel_552491;
  assign add_552498 = sel_552495 + 8'h01;
  assign sel_552499 = array_index_552270 == array_index_537358 ? add_552498 : sel_552495;
  assign add_552502 = sel_552499 + 8'h01;
  assign sel_552503 = array_index_552270 == array_index_537364 ? add_552502 : sel_552499;
  assign add_552506 = sel_552503 + 8'h01;
  assign sel_552507 = array_index_552270 == array_index_537370 ? add_552506 : sel_552503;
  assign add_552510 = sel_552507 + 8'h01;
  assign sel_552511 = array_index_552270 == array_index_537376 ? add_552510 : sel_552507;
  assign add_552514 = sel_552511 + 8'h01;
  assign sel_552515 = array_index_552270 == array_index_537382 ? add_552514 : sel_552511;
  assign add_552518 = sel_552515 + 8'h01;
  assign sel_552519 = array_index_552270 == array_index_537388 ? add_552518 : sel_552515;
  assign add_552522 = sel_552519 + 8'h01;
  assign sel_552523 = array_index_552270 == array_index_537394 ? add_552522 : sel_552519;
  assign add_552526 = sel_552523 + 8'h01;
  assign sel_552527 = array_index_552270 == array_index_537400 ? add_552526 : sel_552523;
  assign add_552530 = sel_552527 + 8'h01;
  assign sel_552531 = array_index_552270 == array_index_537406 ? add_552530 : sel_552527;
  assign add_552534 = sel_552531 + 8'h01;
  assign sel_552535 = array_index_552270 == array_index_537412 ? add_552534 : sel_552531;
  assign add_552538 = sel_552535 + 8'h01;
  assign sel_552539 = array_index_552270 == array_index_537418 ? add_552538 : sel_552535;
  assign add_552542 = sel_552539 + 8'h01;
  assign sel_552543 = array_index_552270 == array_index_537424 ? add_552542 : sel_552539;
  assign add_552546 = sel_552543 + 8'h01;
  assign sel_552547 = array_index_552270 == array_index_537430 ? add_552546 : sel_552543;
  assign add_552550 = sel_552547 + 8'h01;
  assign sel_552551 = array_index_552270 == array_index_537436 ? add_552550 : sel_552547;
  assign add_552554 = sel_552551 + 8'h01;
  assign sel_552555 = array_index_552270 == array_index_537442 ? add_552554 : sel_552551;
  assign add_552558 = sel_552555 + 8'h01;
  assign sel_552559 = array_index_552270 == array_index_537448 ? add_552558 : sel_552555;
  assign add_552562 = sel_552559 + 8'h01;
  assign sel_552563 = array_index_552270 == array_index_537454 ? add_552562 : sel_552559;
  assign add_552566 = sel_552563 + 8'h01;
  assign sel_552567 = array_index_552270 == array_index_537460 ? add_552566 : sel_552563;
  assign add_552571 = sel_552567 + 8'h01;
  assign array_index_552572 = set1_unflattened[7'h33];
  assign sel_552573 = array_index_552270 == array_index_537466 ? add_552571 : sel_552567;
  assign add_552576 = sel_552573 + 8'h01;
  assign sel_552577 = array_index_552572 == array_index_537012 ? add_552576 : sel_552573;
  assign add_552580 = sel_552577 + 8'h01;
  assign sel_552581 = array_index_552572 == array_index_537016 ? add_552580 : sel_552577;
  assign add_552584 = sel_552581 + 8'h01;
  assign sel_552585 = array_index_552572 == array_index_537024 ? add_552584 : sel_552581;
  assign add_552588 = sel_552585 + 8'h01;
  assign sel_552589 = array_index_552572 == array_index_537032 ? add_552588 : sel_552585;
  assign add_552592 = sel_552589 + 8'h01;
  assign sel_552593 = array_index_552572 == array_index_537040 ? add_552592 : sel_552589;
  assign add_552596 = sel_552593 + 8'h01;
  assign sel_552597 = array_index_552572 == array_index_537048 ? add_552596 : sel_552593;
  assign add_552600 = sel_552597 + 8'h01;
  assign sel_552601 = array_index_552572 == array_index_537056 ? add_552600 : sel_552597;
  assign add_552604 = sel_552601 + 8'h01;
  assign sel_552605 = array_index_552572 == array_index_537064 ? add_552604 : sel_552601;
  assign add_552608 = sel_552605 + 8'h01;
  assign sel_552609 = array_index_552572 == array_index_537070 ? add_552608 : sel_552605;
  assign add_552612 = sel_552609 + 8'h01;
  assign sel_552613 = array_index_552572 == array_index_537076 ? add_552612 : sel_552609;
  assign add_552616 = sel_552613 + 8'h01;
  assign sel_552617 = array_index_552572 == array_index_537082 ? add_552616 : sel_552613;
  assign add_552620 = sel_552617 + 8'h01;
  assign sel_552621 = array_index_552572 == array_index_537088 ? add_552620 : sel_552617;
  assign add_552624 = sel_552621 + 8'h01;
  assign sel_552625 = array_index_552572 == array_index_537094 ? add_552624 : sel_552621;
  assign add_552628 = sel_552625 + 8'h01;
  assign sel_552629 = array_index_552572 == array_index_537100 ? add_552628 : sel_552625;
  assign add_552632 = sel_552629 + 8'h01;
  assign sel_552633 = array_index_552572 == array_index_537106 ? add_552632 : sel_552629;
  assign add_552636 = sel_552633 + 8'h01;
  assign sel_552637 = array_index_552572 == array_index_537112 ? add_552636 : sel_552633;
  assign add_552640 = sel_552637 + 8'h01;
  assign sel_552641 = array_index_552572 == array_index_537118 ? add_552640 : sel_552637;
  assign add_552644 = sel_552641 + 8'h01;
  assign sel_552645 = array_index_552572 == array_index_537124 ? add_552644 : sel_552641;
  assign add_552648 = sel_552645 + 8'h01;
  assign sel_552649 = array_index_552572 == array_index_537130 ? add_552648 : sel_552645;
  assign add_552652 = sel_552649 + 8'h01;
  assign sel_552653 = array_index_552572 == array_index_537136 ? add_552652 : sel_552649;
  assign add_552656 = sel_552653 + 8'h01;
  assign sel_552657 = array_index_552572 == array_index_537142 ? add_552656 : sel_552653;
  assign add_552660 = sel_552657 + 8'h01;
  assign sel_552661 = array_index_552572 == array_index_537148 ? add_552660 : sel_552657;
  assign add_552664 = sel_552661 + 8'h01;
  assign sel_552665 = array_index_552572 == array_index_537154 ? add_552664 : sel_552661;
  assign add_552668 = sel_552665 + 8'h01;
  assign sel_552669 = array_index_552572 == array_index_537160 ? add_552668 : sel_552665;
  assign add_552672 = sel_552669 + 8'h01;
  assign sel_552673 = array_index_552572 == array_index_537166 ? add_552672 : sel_552669;
  assign add_552676 = sel_552673 + 8'h01;
  assign sel_552677 = array_index_552572 == array_index_537172 ? add_552676 : sel_552673;
  assign add_552680 = sel_552677 + 8'h01;
  assign sel_552681 = array_index_552572 == array_index_537178 ? add_552680 : sel_552677;
  assign add_552684 = sel_552681 + 8'h01;
  assign sel_552685 = array_index_552572 == array_index_537184 ? add_552684 : sel_552681;
  assign add_552688 = sel_552685 + 8'h01;
  assign sel_552689 = array_index_552572 == array_index_537190 ? add_552688 : sel_552685;
  assign add_552692 = sel_552689 + 8'h01;
  assign sel_552693 = array_index_552572 == array_index_537196 ? add_552692 : sel_552689;
  assign add_552696 = sel_552693 + 8'h01;
  assign sel_552697 = array_index_552572 == array_index_537202 ? add_552696 : sel_552693;
  assign add_552700 = sel_552697 + 8'h01;
  assign sel_552701 = array_index_552572 == array_index_537208 ? add_552700 : sel_552697;
  assign add_552704 = sel_552701 + 8'h01;
  assign sel_552705 = array_index_552572 == array_index_537214 ? add_552704 : sel_552701;
  assign add_552708 = sel_552705 + 8'h01;
  assign sel_552709 = array_index_552572 == array_index_537220 ? add_552708 : sel_552705;
  assign add_552712 = sel_552709 + 8'h01;
  assign sel_552713 = array_index_552572 == array_index_537226 ? add_552712 : sel_552709;
  assign add_552716 = sel_552713 + 8'h01;
  assign sel_552717 = array_index_552572 == array_index_537232 ? add_552716 : sel_552713;
  assign add_552720 = sel_552717 + 8'h01;
  assign sel_552721 = array_index_552572 == array_index_537238 ? add_552720 : sel_552717;
  assign add_552724 = sel_552721 + 8'h01;
  assign sel_552725 = array_index_552572 == array_index_537244 ? add_552724 : sel_552721;
  assign add_552728 = sel_552725 + 8'h01;
  assign sel_552729 = array_index_552572 == array_index_537250 ? add_552728 : sel_552725;
  assign add_552732 = sel_552729 + 8'h01;
  assign sel_552733 = array_index_552572 == array_index_537256 ? add_552732 : sel_552729;
  assign add_552736 = sel_552733 + 8'h01;
  assign sel_552737 = array_index_552572 == array_index_537262 ? add_552736 : sel_552733;
  assign add_552740 = sel_552737 + 8'h01;
  assign sel_552741 = array_index_552572 == array_index_537268 ? add_552740 : sel_552737;
  assign add_552744 = sel_552741 + 8'h01;
  assign sel_552745 = array_index_552572 == array_index_537274 ? add_552744 : sel_552741;
  assign add_552748 = sel_552745 + 8'h01;
  assign sel_552749 = array_index_552572 == array_index_537280 ? add_552748 : sel_552745;
  assign add_552752 = sel_552749 + 8'h01;
  assign sel_552753 = array_index_552572 == array_index_537286 ? add_552752 : sel_552749;
  assign add_552756 = sel_552753 + 8'h01;
  assign sel_552757 = array_index_552572 == array_index_537292 ? add_552756 : sel_552753;
  assign add_552760 = sel_552757 + 8'h01;
  assign sel_552761 = array_index_552572 == array_index_537298 ? add_552760 : sel_552757;
  assign add_552764 = sel_552761 + 8'h01;
  assign sel_552765 = array_index_552572 == array_index_537304 ? add_552764 : sel_552761;
  assign add_552768 = sel_552765 + 8'h01;
  assign sel_552769 = array_index_552572 == array_index_537310 ? add_552768 : sel_552765;
  assign add_552772 = sel_552769 + 8'h01;
  assign sel_552773 = array_index_552572 == array_index_537316 ? add_552772 : sel_552769;
  assign add_552776 = sel_552773 + 8'h01;
  assign sel_552777 = array_index_552572 == array_index_537322 ? add_552776 : sel_552773;
  assign add_552780 = sel_552777 + 8'h01;
  assign sel_552781 = array_index_552572 == array_index_537328 ? add_552780 : sel_552777;
  assign add_552784 = sel_552781 + 8'h01;
  assign sel_552785 = array_index_552572 == array_index_537334 ? add_552784 : sel_552781;
  assign add_552788 = sel_552785 + 8'h01;
  assign sel_552789 = array_index_552572 == array_index_537340 ? add_552788 : sel_552785;
  assign add_552792 = sel_552789 + 8'h01;
  assign sel_552793 = array_index_552572 == array_index_537346 ? add_552792 : sel_552789;
  assign add_552796 = sel_552793 + 8'h01;
  assign sel_552797 = array_index_552572 == array_index_537352 ? add_552796 : sel_552793;
  assign add_552800 = sel_552797 + 8'h01;
  assign sel_552801 = array_index_552572 == array_index_537358 ? add_552800 : sel_552797;
  assign add_552804 = sel_552801 + 8'h01;
  assign sel_552805 = array_index_552572 == array_index_537364 ? add_552804 : sel_552801;
  assign add_552808 = sel_552805 + 8'h01;
  assign sel_552809 = array_index_552572 == array_index_537370 ? add_552808 : sel_552805;
  assign add_552812 = sel_552809 + 8'h01;
  assign sel_552813 = array_index_552572 == array_index_537376 ? add_552812 : sel_552809;
  assign add_552816 = sel_552813 + 8'h01;
  assign sel_552817 = array_index_552572 == array_index_537382 ? add_552816 : sel_552813;
  assign add_552820 = sel_552817 + 8'h01;
  assign sel_552821 = array_index_552572 == array_index_537388 ? add_552820 : sel_552817;
  assign add_552824 = sel_552821 + 8'h01;
  assign sel_552825 = array_index_552572 == array_index_537394 ? add_552824 : sel_552821;
  assign add_552828 = sel_552825 + 8'h01;
  assign sel_552829 = array_index_552572 == array_index_537400 ? add_552828 : sel_552825;
  assign add_552832 = sel_552829 + 8'h01;
  assign sel_552833 = array_index_552572 == array_index_537406 ? add_552832 : sel_552829;
  assign add_552836 = sel_552833 + 8'h01;
  assign sel_552837 = array_index_552572 == array_index_537412 ? add_552836 : sel_552833;
  assign add_552840 = sel_552837 + 8'h01;
  assign sel_552841 = array_index_552572 == array_index_537418 ? add_552840 : sel_552837;
  assign add_552844 = sel_552841 + 8'h01;
  assign sel_552845 = array_index_552572 == array_index_537424 ? add_552844 : sel_552841;
  assign add_552848 = sel_552845 + 8'h01;
  assign sel_552849 = array_index_552572 == array_index_537430 ? add_552848 : sel_552845;
  assign add_552852 = sel_552849 + 8'h01;
  assign sel_552853 = array_index_552572 == array_index_537436 ? add_552852 : sel_552849;
  assign add_552856 = sel_552853 + 8'h01;
  assign sel_552857 = array_index_552572 == array_index_537442 ? add_552856 : sel_552853;
  assign add_552860 = sel_552857 + 8'h01;
  assign sel_552861 = array_index_552572 == array_index_537448 ? add_552860 : sel_552857;
  assign add_552864 = sel_552861 + 8'h01;
  assign sel_552865 = array_index_552572 == array_index_537454 ? add_552864 : sel_552861;
  assign add_552868 = sel_552865 + 8'h01;
  assign sel_552869 = array_index_552572 == array_index_537460 ? add_552868 : sel_552865;
  assign add_552873 = sel_552869 + 8'h01;
  assign array_index_552874 = set1_unflattened[7'h34];
  assign sel_552875 = array_index_552572 == array_index_537466 ? add_552873 : sel_552869;
  assign add_552878 = sel_552875 + 8'h01;
  assign sel_552879 = array_index_552874 == array_index_537012 ? add_552878 : sel_552875;
  assign add_552882 = sel_552879 + 8'h01;
  assign sel_552883 = array_index_552874 == array_index_537016 ? add_552882 : sel_552879;
  assign add_552886 = sel_552883 + 8'h01;
  assign sel_552887 = array_index_552874 == array_index_537024 ? add_552886 : sel_552883;
  assign add_552890 = sel_552887 + 8'h01;
  assign sel_552891 = array_index_552874 == array_index_537032 ? add_552890 : sel_552887;
  assign add_552894 = sel_552891 + 8'h01;
  assign sel_552895 = array_index_552874 == array_index_537040 ? add_552894 : sel_552891;
  assign add_552898 = sel_552895 + 8'h01;
  assign sel_552899 = array_index_552874 == array_index_537048 ? add_552898 : sel_552895;
  assign add_552902 = sel_552899 + 8'h01;
  assign sel_552903 = array_index_552874 == array_index_537056 ? add_552902 : sel_552899;
  assign add_552906 = sel_552903 + 8'h01;
  assign sel_552907 = array_index_552874 == array_index_537064 ? add_552906 : sel_552903;
  assign add_552910 = sel_552907 + 8'h01;
  assign sel_552911 = array_index_552874 == array_index_537070 ? add_552910 : sel_552907;
  assign add_552914 = sel_552911 + 8'h01;
  assign sel_552915 = array_index_552874 == array_index_537076 ? add_552914 : sel_552911;
  assign add_552918 = sel_552915 + 8'h01;
  assign sel_552919 = array_index_552874 == array_index_537082 ? add_552918 : sel_552915;
  assign add_552922 = sel_552919 + 8'h01;
  assign sel_552923 = array_index_552874 == array_index_537088 ? add_552922 : sel_552919;
  assign add_552926 = sel_552923 + 8'h01;
  assign sel_552927 = array_index_552874 == array_index_537094 ? add_552926 : sel_552923;
  assign add_552930 = sel_552927 + 8'h01;
  assign sel_552931 = array_index_552874 == array_index_537100 ? add_552930 : sel_552927;
  assign add_552934 = sel_552931 + 8'h01;
  assign sel_552935 = array_index_552874 == array_index_537106 ? add_552934 : sel_552931;
  assign add_552938 = sel_552935 + 8'h01;
  assign sel_552939 = array_index_552874 == array_index_537112 ? add_552938 : sel_552935;
  assign add_552942 = sel_552939 + 8'h01;
  assign sel_552943 = array_index_552874 == array_index_537118 ? add_552942 : sel_552939;
  assign add_552946 = sel_552943 + 8'h01;
  assign sel_552947 = array_index_552874 == array_index_537124 ? add_552946 : sel_552943;
  assign add_552950 = sel_552947 + 8'h01;
  assign sel_552951 = array_index_552874 == array_index_537130 ? add_552950 : sel_552947;
  assign add_552954 = sel_552951 + 8'h01;
  assign sel_552955 = array_index_552874 == array_index_537136 ? add_552954 : sel_552951;
  assign add_552958 = sel_552955 + 8'h01;
  assign sel_552959 = array_index_552874 == array_index_537142 ? add_552958 : sel_552955;
  assign add_552962 = sel_552959 + 8'h01;
  assign sel_552963 = array_index_552874 == array_index_537148 ? add_552962 : sel_552959;
  assign add_552966 = sel_552963 + 8'h01;
  assign sel_552967 = array_index_552874 == array_index_537154 ? add_552966 : sel_552963;
  assign add_552970 = sel_552967 + 8'h01;
  assign sel_552971 = array_index_552874 == array_index_537160 ? add_552970 : sel_552967;
  assign add_552974 = sel_552971 + 8'h01;
  assign sel_552975 = array_index_552874 == array_index_537166 ? add_552974 : sel_552971;
  assign add_552978 = sel_552975 + 8'h01;
  assign sel_552979 = array_index_552874 == array_index_537172 ? add_552978 : sel_552975;
  assign add_552982 = sel_552979 + 8'h01;
  assign sel_552983 = array_index_552874 == array_index_537178 ? add_552982 : sel_552979;
  assign add_552986 = sel_552983 + 8'h01;
  assign sel_552987 = array_index_552874 == array_index_537184 ? add_552986 : sel_552983;
  assign add_552990 = sel_552987 + 8'h01;
  assign sel_552991 = array_index_552874 == array_index_537190 ? add_552990 : sel_552987;
  assign add_552994 = sel_552991 + 8'h01;
  assign sel_552995 = array_index_552874 == array_index_537196 ? add_552994 : sel_552991;
  assign add_552998 = sel_552995 + 8'h01;
  assign sel_552999 = array_index_552874 == array_index_537202 ? add_552998 : sel_552995;
  assign add_553002 = sel_552999 + 8'h01;
  assign sel_553003 = array_index_552874 == array_index_537208 ? add_553002 : sel_552999;
  assign add_553006 = sel_553003 + 8'h01;
  assign sel_553007 = array_index_552874 == array_index_537214 ? add_553006 : sel_553003;
  assign add_553010 = sel_553007 + 8'h01;
  assign sel_553011 = array_index_552874 == array_index_537220 ? add_553010 : sel_553007;
  assign add_553014 = sel_553011 + 8'h01;
  assign sel_553015 = array_index_552874 == array_index_537226 ? add_553014 : sel_553011;
  assign add_553018 = sel_553015 + 8'h01;
  assign sel_553019 = array_index_552874 == array_index_537232 ? add_553018 : sel_553015;
  assign add_553022 = sel_553019 + 8'h01;
  assign sel_553023 = array_index_552874 == array_index_537238 ? add_553022 : sel_553019;
  assign add_553026 = sel_553023 + 8'h01;
  assign sel_553027 = array_index_552874 == array_index_537244 ? add_553026 : sel_553023;
  assign add_553030 = sel_553027 + 8'h01;
  assign sel_553031 = array_index_552874 == array_index_537250 ? add_553030 : sel_553027;
  assign add_553034 = sel_553031 + 8'h01;
  assign sel_553035 = array_index_552874 == array_index_537256 ? add_553034 : sel_553031;
  assign add_553038 = sel_553035 + 8'h01;
  assign sel_553039 = array_index_552874 == array_index_537262 ? add_553038 : sel_553035;
  assign add_553042 = sel_553039 + 8'h01;
  assign sel_553043 = array_index_552874 == array_index_537268 ? add_553042 : sel_553039;
  assign add_553046 = sel_553043 + 8'h01;
  assign sel_553047 = array_index_552874 == array_index_537274 ? add_553046 : sel_553043;
  assign add_553050 = sel_553047 + 8'h01;
  assign sel_553051 = array_index_552874 == array_index_537280 ? add_553050 : sel_553047;
  assign add_553054 = sel_553051 + 8'h01;
  assign sel_553055 = array_index_552874 == array_index_537286 ? add_553054 : sel_553051;
  assign add_553058 = sel_553055 + 8'h01;
  assign sel_553059 = array_index_552874 == array_index_537292 ? add_553058 : sel_553055;
  assign add_553062 = sel_553059 + 8'h01;
  assign sel_553063 = array_index_552874 == array_index_537298 ? add_553062 : sel_553059;
  assign add_553066 = sel_553063 + 8'h01;
  assign sel_553067 = array_index_552874 == array_index_537304 ? add_553066 : sel_553063;
  assign add_553070 = sel_553067 + 8'h01;
  assign sel_553071 = array_index_552874 == array_index_537310 ? add_553070 : sel_553067;
  assign add_553074 = sel_553071 + 8'h01;
  assign sel_553075 = array_index_552874 == array_index_537316 ? add_553074 : sel_553071;
  assign add_553078 = sel_553075 + 8'h01;
  assign sel_553079 = array_index_552874 == array_index_537322 ? add_553078 : sel_553075;
  assign add_553082 = sel_553079 + 8'h01;
  assign sel_553083 = array_index_552874 == array_index_537328 ? add_553082 : sel_553079;
  assign add_553086 = sel_553083 + 8'h01;
  assign sel_553087 = array_index_552874 == array_index_537334 ? add_553086 : sel_553083;
  assign add_553090 = sel_553087 + 8'h01;
  assign sel_553091 = array_index_552874 == array_index_537340 ? add_553090 : sel_553087;
  assign add_553094 = sel_553091 + 8'h01;
  assign sel_553095 = array_index_552874 == array_index_537346 ? add_553094 : sel_553091;
  assign add_553098 = sel_553095 + 8'h01;
  assign sel_553099 = array_index_552874 == array_index_537352 ? add_553098 : sel_553095;
  assign add_553102 = sel_553099 + 8'h01;
  assign sel_553103 = array_index_552874 == array_index_537358 ? add_553102 : sel_553099;
  assign add_553106 = sel_553103 + 8'h01;
  assign sel_553107 = array_index_552874 == array_index_537364 ? add_553106 : sel_553103;
  assign add_553110 = sel_553107 + 8'h01;
  assign sel_553111 = array_index_552874 == array_index_537370 ? add_553110 : sel_553107;
  assign add_553114 = sel_553111 + 8'h01;
  assign sel_553115 = array_index_552874 == array_index_537376 ? add_553114 : sel_553111;
  assign add_553118 = sel_553115 + 8'h01;
  assign sel_553119 = array_index_552874 == array_index_537382 ? add_553118 : sel_553115;
  assign add_553122 = sel_553119 + 8'h01;
  assign sel_553123 = array_index_552874 == array_index_537388 ? add_553122 : sel_553119;
  assign add_553126 = sel_553123 + 8'h01;
  assign sel_553127 = array_index_552874 == array_index_537394 ? add_553126 : sel_553123;
  assign add_553130 = sel_553127 + 8'h01;
  assign sel_553131 = array_index_552874 == array_index_537400 ? add_553130 : sel_553127;
  assign add_553134 = sel_553131 + 8'h01;
  assign sel_553135 = array_index_552874 == array_index_537406 ? add_553134 : sel_553131;
  assign add_553138 = sel_553135 + 8'h01;
  assign sel_553139 = array_index_552874 == array_index_537412 ? add_553138 : sel_553135;
  assign add_553142 = sel_553139 + 8'h01;
  assign sel_553143 = array_index_552874 == array_index_537418 ? add_553142 : sel_553139;
  assign add_553146 = sel_553143 + 8'h01;
  assign sel_553147 = array_index_552874 == array_index_537424 ? add_553146 : sel_553143;
  assign add_553150 = sel_553147 + 8'h01;
  assign sel_553151 = array_index_552874 == array_index_537430 ? add_553150 : sel_553147;
  assign add_553154 = sel_553151 + 8'h01;
  assign sel_553155 = array_index_552874 == array_index_537436 ? add_553154 : sel_553151;
  assign add_553158 = sel_553155 + 8'h01;
  assign sel_553159 = array_index_552874 == array_index_537442 ? add_553158 : sel_553155;
  assign add_553162 = sel_553159 + 8'h01;
  assign sel_553163 = array_index_552874 == array_index_537448 ? add_553162 : sel_553159;
  assign add_553166 = sel_553163 + 8'h01;
  assign sel_553167 = array_index_552874 == array_index_537454 ? add_553166 : sel_553163;
  assign add_553170 = sel_553167 + 8'h01;
  assign sel_553171 = array_index_552874 == array_index_537460 ? add_553170 : sel_553167;
  assign add_553175 = sel_553171 + 8'h01;
  assign array_index_553176 = set1_unflattened[7'h35];
  assign sel_553177 = array_index_552874 == array_index_537466 ? add_553175 : sel_553171;
  assign add_553180 = sel_553177 + 8'h01;
  assign sel_553181 = array_index_553176 == array_index_537012 ? add_553180 : sel_553177;
  assign add_553184 = sel_553181 + 8'h01;
  assign sel_553185 = array_index_553176 == array_index_537016 ? add_553184 : sel_553181;
  assign add_553188 = sel_553185 + 8'h01;
  assign sel_553189 = array_index_553176 == array_index_537024 ? add_553188 : sel_553185;
  assign add_553192 = sel_553189 + 8'h01;
  assign sel_553193 = array_index_553176 == array_index_537032 ? add_553192 : sel_553189;
  assign add_553196 = sel_553193 + 8'h01;
  assign sel_553197 = array_index_553176 == array_index_537040 ? add_553196 : sel_553193;
  assign add_553200 = sel_553197 + 8'h01;
  assign sel_553201 = array_index_553176 == array_index_537048 ? add_553200 : sel_553197;
  assign add_553204 = sel_553201 + 8'h01;
  assign sel_553205 = array_index_553176 == array_index_537056 ? add_553204 : sel_553201;
  assign add_553208 = sel_553205 + 8'h01;
  assign sel_553209 = array_index_553176 == array_index_537064 ? add_553208 : sel_553205;
  assign add_553212 = sel_553209 + 8'h01;
  assign sel_553213 = array_index_553176 == array_index_537070 ? add_553212 : sel_553209;
  assign add_553216 = sel_553213 + 8'h01;
  assign sel_553217 = array_index_553176 == array_index_537076 ? add_553216 : sel_553213;
  assign add_553220 = sel_553217 + 8'h01;
  assign sel_553221 = array_index_553176 == array_index_537082 ? add_553220 : sel_553217;
  assign add_553224 = sel_553221 + 8'h01;
  assign sel_553225 = array_index_553176 == array_index_537088 ? add_553224 : sel_553221;
  assign add_553228 = sel_553225 + 8'h01;
  assign sel_553229 = array_index_553176 == array_index_537094 ? add_553228 : sel_553225;
  assign add_553232 = sel_553229 + 8'h01;
  assign sel_553233 = array_index_553176 == array_index_537100 ? add_553232 : sel_553229;
  assign add_553236 = sel_553233 + 8'h01;
  assign sel_553237 = array_index_553176 == array_index_537106 ? add_553236 : sel_553233;
  assign add_553240 = sel_553237 + 8'h01;
  assign sel_553241 = array_index_553176 == array_index_537112 ? add_553240 : sel_553237;
  assign add_553244 = sel_553241 + 8'h01;
  assign sel_553245 = array_index_553176 == array_index_537118 ? add_553244 : sel_553241;
  assign add_553248 = sel_553245 + 8'h01;
  assign sel_553249 = array_index_553176 == array_index_537124 ? add_553248 : sel_553245;
  assign add_553252 = sel_553249 + 8'h01;
  assign sel_553253 = array_index_553176 == array_index_537130 ? add_553252 : sel_553249;
  assign add_553256 = sel_553253 + 8'h01;
  assign sel_553257 = array_index_553176 == array_index_537136 ? add_553256 : sel_553253;
  assign add_553260 = sel_553257 + 8'h01;
  assign sel_553261 = array_index_553176 == array_index_537142 ? add_553260 : sel_553257;
  assign add_553264 = sel_553261 + 8'h01;
  assign sel_553265 = array_index_553176 == array_index_537148 ? add_553264 : sel_553261;
  assign add_553268 = sel_553265 + 8'h01;
  assign sel_553269 = array_index_553176 == array_index_537154 ? add_553268 : sel_553265;
  assign add_553272 = sel_553269 + 8'h01;
  assign sel_553273 = array_index_553176 == array_index_537160 ? add_553272 : sel_553269;
  assign add_553276 = sel_553273 + 8'h01;
  assign sel_553277 = array_index_553176 == array_index_537166 ? add_553276 : sel_553273;
  assign add_553280 = sel_553277 + 8'h01;
  assign sel_553281 = array_index_553176 == array_index_537172 ? add_553280 : sel_553277;
  assign add_553284 = sel_553281 + 8'h01;
  assign sel_553285 = array_index_553176 == array_index_537178 ? add_553284 : sel_553281;
  assign add_553288 = sel_553285 + 8'h01;
  assign sel_553289 = array_index_553176 == array_index_537184 ? add_553288 : sel_553285;
  assign add_553292 = sel_553289 + 8'h01;
  assign sel_553293 = array_index_553176 == array_index_537190 ? add_553292 : sel_553289;
  assign add_553296 = sel_553293 + 8'h01;
  assign sel_553297 = array_index_553176 == array_index_537196 ? add_553296 : sel_553293;
  assign add_553300 = sel_553297 + 8'h01;
  assign sel_553301 = array_index_553176 == array_index_537202 ? add_553300 : sel_553297;
  assign add_553304 = sel_553301 + 8'h01;
  assign sel_553305 = array_index_553176 == array_index_537208 ? add_553304 : sel_553301;
  assign add_553308 = sel_553305 + 8'h01;
  assign sel_553309 = array_index_553176 == array_index_537214 ? add_553308 : sel_553305;
  assign add_553312 = sel_553309 + 8'h01;
  assign sel_553313 = array_index_553176 == array_index_537220 ? add_553312 : sel_553309;
  assign add_553316 = sel_553313 + 8'h01;
  assign sel_553317 = array_index_553176 == array_index_537226 ? add_553316 : sel_553313;
  assign add_553320 = sel_553317 + 8'h01;
  assign sel_553321 = array_index_553176 == array_index_537232 ? add_553320 : sel_553317;
  assign add_553324 = sel_553321 + 8'h01;
  assign sel_553325 = array_index_553176 == array_index_537238 ? add_553324 : sel_553321;
  assign add_553328 = sel_553325 + 8'h01;
  assign sel_553329 = array_index_553176 == array_index_537244 ? add_553328 : sel_553325;
  assign add_553332 = sel_553329 + 8'h01;
  assign sel_553333 = array_index_553176 == array_index_537250 ? add_553332 : sel_553329;
  assign add_553336 = sel_553333 + 8'h01;
  assign sel_553337 = array_index_553176 == array_index_537256 ? add_553336 : sel_553333;
  assign add_553340 = sel_553337 + 8'h01;
  assign sel_553341 = array_index_553176 == array_index_537262 ? add_553340 : sel_553337;
  assign add_553344 = sel_553341 + 8'h01;
  assign sel_553345 = array_index_553176 == array_index_537268 ? add_553344 : sel_553341;
  assign add_553348 = sel_553345 + 8'h01;
  assign sel_553349 = array_index_553176 == array_index_537274 ? add_553348 : sel_553345;
  assign add_553352 = sel_553349 + 8'h01;
  assign sel_553353 = array_index_553176 == array_index_537280 ? add_553352 : sel_553349;
  assign add_553356 = sel_553353 + 8'h01;
  assign sel_553357 = array_index_553176 == array_index_537286 ? add_553356 : sel_553353;
  assign add_553360 = sel_553357 + 8'h01;
  assign sel_553361 = array_index_553176 == array_index_537292 ? add_553360 : sel_553357;
  assign add_553364 = sel_553361 + 8'h01;
  assign sel_553365 = array_index_553176 == array_index_537298 ? add_553364 : sel_553361;
  assign add_553368 = sel_553365 + 8'h01;
  assign sel_553369 = array_index_553176 == array_index_537304 ? add_553368 : sel_553365;
  assign add_553372 = sel_553369 + 8'h01;
  assign sel_553373 = array_index_553176 == array_index_537310 ? add_553372 : sel_553369;
  assign add_553376 = sel_553373 + 8'h01;
  assign sel_553377 = array_index_553176 == array_index_537316 ? add_553376 : sel_553373;
  assign add_553380 = sel_553377 + 8'h01;
  assign sel_553381 = array_index_553176 == array_index_537322 ? add_553380 : sel_553377;
  assign add_553384 = sel_553381 + 8'h01;
  assign sel_553385 = array_index_553176 == array_index_537328 ? add_553384 : sel_553381;
  assign add_553388 = sel_553385 + 8'h01;
  assign sel_553389 = array_index_553176 == array_index_537334 ? add_553388 : sel_553385;
  assign add_553392 = sel_553389 + 8'h01;
  assign sel_553393 = array_index_553176 == array_index_537340 ? add_553392 : sel_553389;
  assign add_553396 = sel_553393 + 8'h01;
  assign sel_553397 = array_index_553176 == array_index_537346 ? add_553396 : sel_553393;
  assign add_553400 = sel_553397 + 8'h01;
  assign sel_553401 = array_index_553176 == array_index_537352 ? add_553400 : sel_553397;
  assign add_553404 = sel_553401 + 8'h01;
  assign sel_553405 = array_index_553176 == array_index_537358 ? add_553404 : sel_553401;
  assign add_553408 = sel_553405 + 8'h01;
  assign sel_553409 = array_index_553176 == array_index_537364 ? add_553408 : sel_553405;
  assign add_553412 = sel_553409 + 8'h01;
  assign sel_553413 = array_index_553176 == array_index_537370 ? add_553412 : sel_553409;
  assign add_553416 = sel_553413 + 8'h01;
  assign sel_553417 = array_index_553176 == array_index_537376 ? add_553416 : sel_553413;
  assign add_553420 = sel_553417 + 8'h01;
  assign sel_553421 = array_index_553176 == array_index_537382 ? add_553420 : sel_553417;
  assign add_553424 = sel_553421 + 8'h01;
  assign sel_553425 = array_index_553176 == array_index_537388 ? add_553424 : sel_553421;
  assign add_553428 = sel_553425 + 8'h01;
  assign sel_553429 = array_index_553176 == array_index_537394 ? add_553428 : sel_553425;
  assign add_553432 = sel_553429 + 8'h01;
  assign sel_553433 = array_index_553176 == array_index_537400 ? add_553432 : sel_553429;
  assign add_553436 = sel_553433 + 8'h01;
  assign sel_553437 = array_index_553176 == array_index_537406 ? add_553436 : sel_553433;
  assign add_553440 = sel_553437 + 8'h01;
  assign sel_553441 = array_index_553176 == array_index_537412 ? add_553440 : sel_553437;
  assign add_553444 = sel_553441 + 8'h01;
  assign sel_553445 = array_index_553176 == array_index_537418 ? add_553444 : sel_553441;
  assign add_553448 = sel_553445 + 8'h01;
  assign sel_553449 = array_index_553176 == array_index_537424 ? add_553448 : sel_553445;
  assign add_553452 = sel_553449 + 8'h01;
  assign sel_553453 = array_index_553176 == array_index_537430 ? add_553452 : sel_553449;
  assign add_553456 = sel_553453 + 8'h01;
  assign sel_553457 = array_index_553176 == array_index_537436 ? add_553456 : sel_553453;
  assign add_553460 = sel_553457 + 8'h01;
  assign sel_553461 = array_index_553176 == array_index_537442 ? add_553460 : sel_553457;
  assign add_553464 = sel_553461 + 8'h01;
  assign sel_553465 = array_index_553176 == array_index_537448 ? add_553464 : sel_553461;
  assign add_553468 = sel_553465 + 8'h01;
  assign sel_553469 = array_index_553176 == array_index_537454 ? add_553468 : sel_553465;
  assign add_553472 = sel_553469 + 8'h01;
  assign sel_553473 = array_index_553176 == array_index_537460 ? add_553472 : sel_553469;
  assign add_553477 = sel_553473 + 8'h01;
  assign array_index_553478 = set1_unflattened[7'h36];
  assign sel_553479 = array_index_553176 == array_index_537466 ? add_553477 : sel_553473;
  assign add_553482 = sel_553479 + 8'h01;
  assign sel_553483 = array_index_553478 == array_index_537012 ? add_553482 : sel_553479;
  assign add_553486 = sel_553483 + 8'h01;
  assign sel_553487 = array_index_553478 == array_index_537016 ? add_553486 : sel_553483;
  assign add_553490 = sel_553487 + 8'h01;
  assign sel_553491 = array_index_553478 == array_index_537024 ? add_553490 : sel_553487;
  assign add_553494 = sel_553491 + 8'h01;
  assign sel_553495 = array_index_553478 == array_index_537032 ? add_553494 : sel_553491;
  assign add_553498 = sel_553495 + 8'h01;
  assign sel_553499 = array_index_553478 == array_index_537040 ? add_553498 : sel_553495;
  assign add_553502 = sel_553499 + 8'h01;
  assign sel_553503 = array_index_553478 == array_index_537048 ? add_553502 : sel_553499;
  assign add_553506 = sel_553503 + 8'h01;
  assign sel_553507 = array_index_553478 == array_index_537056 ? add_553506 : sel_553503;
  assign add_553510 = sel_553507 + 8'h01;
  assign sel_553511 = array_index_553478 == array_index_537064 ? add_553510 : sel_553507;
  assign add_553514 = sel_553511 + 8'h01;
  assign sel_553515 = array_index_553478 == array_index_537070 ? add_553514 : sel_553511;
  assign add_553518 = sel_553515 + 8'h01;
  assign sel_553519 = array_index_553478 == array_index_537076 ? add_553518 : sel_553515;
  assign add_553522 = sel_553519 + 8'h01;
  assign sel_553523 = array_index_553478 == array_index_537082 ? add_553522 : sel_553519;
  assign add_553526 = sel_553523 + 8'h01;
  assign sel_553527 = array_index_553478 == array_index_537088 ? add_553526 : sel_553523;
  assign add_553530 = sel_553527 + 8'h01;
  assign sel_553531 = array_index_553478 == array_index_537094 ? add_553530 : sel_553527;
  assign add_553534 = sel_553531 + 8'h01;
  assign sel_553535 = array_index_553478 == array_index_537100 ? add_553534 : sel_553531;
  assign add_553538 = sel_553535 + 8'h01;
  assign sel_553539 = array_index_553478 == array_index_537106 ? add_553538 : sel_553535;
  assign add_553542 = sel_553539 + 8'h01;
  assign sel_553543 = array_index_553478 == array_index_537112 ? add_553542 : sel_553539;
  assign add_553546 = sel_553543 + 8'h01;
  assign sel_553547 = array_index_553478 == array_index_537118 ? add_553546 : sel_553543;
  assign add_553550 = sel_553547 + 8'h01;
  assign sel_553551 = array_index_553478 == array_index_537124 ? add_553550 : sel_553547;
  assign add_553554 = sel_553551 + 8'h01;
  assign sel_553555 = array_index_553478 == array_index_537130 ? add_553554 : sel_553551;
  assign add_553558 = sel_553555 + 8'h01;
  assign sel_553559 = array_index_553478 == array_index_537136 ? add_553558 : sel_553555;
  assign add_553562 = sel_553559 + 8'h01;
  assign sel_553563 = array_index_553478 == array_index_537142 ? add_553562 : sel_553559;
  assign add_553566 = sel_553563 + 8'h01;
  assign sel_553567 = array_index_553478 == array_index_537148 ? add_553566 : sel_553563;
  assign add_553570 = sel_553567 + 8'h01;
  assign sel_553571 = array_index_553478 == array_index_537154 ? add_553570 : sel_553567;
  assign add_553574 = sel_553571 + 8'h01;
  assign sel_553575 = array_index_553478 == array_index_537160 ? add_553574 : sel_553571;
  assign add_553578 = sel_553575 + 8'h01;
  assign sel_553579 = array_index_553478 == array_index_537166 ? add_553578 : sel_553575;
  assign add_553582 = sel_553579 + 8'h01;
  assign sel_553583 = array_index_553478 == array_index_537172 ? add_553582 : sel_553579;
  assign add_553586 = sel_553583 + 8'h01;
  assign sel_553587 = array_index_553478 == array_index_537178 ? add_553586 : sel_553583;
  assign add_553590 = sel_553587 + 8'h01;
  assign sel_553591 = array_index_553478 == array_index_537184 ? add_553590 : sel_553587;
  assign add_553594 = sel_553591 + 8'h01;
  assign sel_553595 = array_index_553478 == array_index_537190 ? add_553594 : sel_553591;
  assign add_553598 = sel_553595 + 8'h01;
  assign sel_553599 = array_index_553478 == array_index_537196 ? add_553598 : sel_553595;
  assign add_553602 = sel_553599 + 8'h01;
  assign sel_553603 = array_index_553478 == array_index_537202 ? add_553602 : sel_553599;
  assign add_553606 = sel_553603 + 8'h01;
  assign sel_553607 = array_index_553478 == array_index_537208 ? add_553606 : sel_553603;
  assign add_553610 = sel_553607 + 8'h01;
  assign sel_553611 = array_index_553478 == array_index_537214 ? add_553610 : sel_553607;
  assign add_553614 = sel_553611 + 8'h01;
  assign sel_553615 = array_index_553478 == array_index_537220 ? add_553614 : sel_553611;
  assign add_553618 = sel_553615 + 8'h01;
  assign sel_553619 = array_index_553478 == array_index_537226 ? add_553618 : sel_553615;
  assign add_553622 = sel_553619 + 8'h01;
  assign sel_553623 = array_index_553478 == array_index_537232 ? add_553622 : sel_553619;
  assign add_553626 = sel_553623 + 8'h01;
  assign sel_553627 = array_index_553478 == array_index_537238 ? add_553626 : sel_553623;
  assign add_553630 = sel_553627 + 8'h01;
  assign sel_553631 = array_index_553478 == array_index_537244 ? add_553630 : sel_553627;
  assign add_553634 = sel_553631 + 8'h01;
  assign sel_553635 = array_index_553478 == array_index_537250 ? add_553634 : sel_553631;
  assign add_553638 = sel_553635 + 8'h01;
  assign sel_553639 = array_index_553478 == array_index_537256 ? add_553638 : sel_553635;
  assign add_553642 = sel_553639 + 8'h01;
  assign sel_553643 = array_index_553478 == array_index_537262 ? add_553642 : sel_553639;
  assign add_553646 = sel_553643 + 8'h01;
  assign sel_553647 = array_index_553478 == array_index_537268 ? add_553646 : sel_553643;
  assign add_553650 = sel_553647 + 8'h01;
  assign sel_553651 = array_index_553478 == array_index_537274 ? add_553650 : sel_553647;
  assign add_553654 = sel_553651 + 8'h01;
  assign sel_553655 = array_index_553478 == array_index_537280 ? add_553654 : sel_553651;
  assign add_553658 = sel_553655 + 8'h01;
  assign sel_553659 = array_index_553478 == array_index_537286 ? add_553658 : sel_553655;
  assign add_553662 = sel_553659 + 8'h01;
  assign sel_553663 = array_index_553478 == array_index_537292 ? add_553662 : sel_553659;
  assign add_553666 = sel_553663 + 8'h01;
  assign sel_553667 = array_index_553478 == array_index_537298 ? add_553666 : sel_553663;
  assign add_553670 = sel_553667 + 8'h01;
  assign sel_553671 = array_index_553478 == array_index_537304 ? add_553670 : sel_553667;
  assign add_553674 = sel_553671 + 8'h01;
  assign sel_553675 = array_index_553478 == array_index_537310 ? add_553674 : sel_553671;
  assign add_553678 = sel_553675 + 8'h01;
  assign sel_553679 = array_index_553478 == array_index_537316 ? add_553678 : sel_553675;
  assign add_553682 = sel_553679 + 8'h01;
  assign sel_553683 = array_index_553478 == array_index_537322 ? add_553682 : sel_553679;
  assign add_553686 = sel_553683 + 8'h01;
  assign sel_553687 = array_index_553478 == array_index_537328 ? add_553686 : sel_553683;
  assign add_553690 = sel_553687 + 8'h01;
  assign sel_553691 = array_index_553478 == array_index_537334 ? add_553690 : sel_553687;
  assign add_553694 = sel_553691 + 8'h01;
  assign sel_553695 = array_index_553478 == array_index_537340 ? add_553694 : sel_553691;
  assign add_553698 = sel_553695 + 8'h01;
  assign sel_553699 = array_index_553478 == array_index_537346 ? add_553698 : sel_553695;
  assign add_553702 = sel_553699 + 8'h01;
  assign sel_553703 = array_index_553478 == array_index_537352 ? add_553702 : sel_553699;
  assign add_553706 = sel_553703 + 8'h01;
  assign sel_553707 = array_index_553478 == array_index_537358 ? add_553706 : sel_553703;
  assign add_553710 = sel_553707 + 8'h01;
  assign sel_553711 = array_index_553478 == array_index_537364 ? add_553710 : sel_553707;
  assign add_553714 = sel_553711 + 8'h01;
  assign sel_553715 = array_index_553478 == array_index_537370 ? add_553714 : sel_553711;
  assign add_553718 = sel_553715 + 8'h01;
  assign sel_553719 = array_index_553478 == array_index_537376 ? add_553718 : sel_553715;
  assign add_553722 = sel_553719 + 8'h01;
  assign sel_553723 = array_index_553478 == array_index_537382 ? add_553722 : sel_553719;
  assign add_553726 = sel_553723 + 8'h01;
  assign sel_553727 = array_index_553478 == array_index_537388 ? add_553726 : sel_553723;
  assign add_553730 = sel_553727 + 8'h01;
  assign sel_553731 = array_index_553478 == array_index_537394 ? add_553730 : sel_553727;
  assign add_553734 = sel_553731 + 8'h01;
  assign sel_553735 = array_index_553478 == array_index_537400 ? add_553734 : sel_553731;
  assign add_553738 = sel_553735 + 8'h01;
  assign sel_553739 = array_index_553478 == array_index_537406 ? add_553738 : sel_553735;
  assign add_553742 = sel_553739 + 8'h01;
  assign sel_553743 = array_index_553478 == array_index_537412 ? add_553742 : sel_553739;
  assign add_553746 = sel_553743 + 8'h01;
  assign sel_553747 = array_index_553478 == array_index_537418 ? add_553746 : sel_553743;
  assign add_553750 = sel_553747 + 8'h01;
  assign sel_553751 = array_index_553478 == array_index_537424 ? add_553750 : sel_553747;
  assign add_553754 = sel_553751 + 8'h01;
  assign sel_553755 = array_index_553478 == array_index_537430 ? add_553754 : sel_553751;
  assign add_553758 = sel_553755 + 8'h01;
  assign sel_553759 = array_index_553478 == array_index_537436 ? add_553758 : sel_553755;
  assign add_553762 = sel_553759 + 8'h01;
  assign sel_553763 = array_index_553478 == array_index_537442 ? add_553762 : sel_553759;
  assign add_553766 = sel_553763 + 8'h01;
  assign sel_553767 = array_index_553478 == array_index_537448 ? add_553766 : sel_553763;
  assign add_553770 = sel_553767 + 8'h01;
  assign sel_553771 = array_index_553478 == array_index_537454 ? add_553770 : sel_553767;
  assign add_553774 = sel_553771 + 8'h01;
  assign sel_553775 = array_index_553478 == array_index_537460 ? add_553774 : sel_553771;
  assign add_553779 = sel_553775 + 8'h01;
  assign array_index_553780 = set1_unflattened[7'h37];
  assign sel_553781 = array_index_553478 == array_index_537466 ? add_553779 : sel_553775;
  assign add_553784 = sel_553781 + 8'h01;
  assign sel_553785 = array_index_553780 == array_index_537012 ? add_553784 : sel_553781;
  assign add_553788 = sel_553785 + 8'h01;
  assign sel_553789 = array_index_553780 == array_index_537016 ? add_553788 : sel_553785;
  assign add_553792 = sel_553789 + 8'h01;
  assign sel_553793 = array_index_553780 == array_index_537024 ? add_553792 : sel_553789;
  assign add_553796 = sel_553793 + 8'h01;
  assign sel_553797 = array_index_553780 == array_index_537032 ? add_553796 : sel_553793;
  assign add_553800 = sel_553797 + 8'h01;
  assign sel_553801 = array_index_553780 == array_index_537040 ? add_553800 : sel_553797;
  assign add_553804 = sel_553801 + 8'h01;
  assign sel_553805 = array_index_553780 == array_index_537048 ? add_553804 : sel_553801;
  assign add_553808 = sel_553805 + 8'h01;
  assign sel_553809 = array_index_553780 == array_index_537056 ? add_553808 : sel_553805;
  assign add_553812 = sel_553809 + 8'h01;
  assign sel_553813 = array_index_553780 == array_index_537064 ? add_553812 : sel_553809;
  assign add_553816 = sel_553813 + 8'h01;
  assign sel_553817 = array_index_553780 == array_index_537070 ? add_553816 : sel_553813;
  assign add_553820 = sel_553817 + 8'h01;
  assign sel_553821 = array_index_553780 == array_index_537076 ? add_553820 : sel_553817;
  assign add_553824 = sel_553821 + 8'h01;
  assign sel_553825 = array_index_553780 == array_index_537082 ? add_553824 : sel_553821;
  assign add_553828 = sel_553825 + 8'h01;
  assign sel_553829 = array_index_553780 == array_index_537088 ? add_553828 : sel_553825;
  assign add_553832 = sel_553829 + 8'h01;
  assign sel_553833 = array_index_553780 == array_index_537094 ? add_553832 : sel_553829;
  assign add_553836 = sel_553833 + 8'h01;
  assign sel_553837 = array_index_553780 == array_index_537100 ? add_553836 : sel_553833;
  assign add_553840 = sel_553837 + 8'h01;
  assign sel_553841 = array_index_553780 == array_index_537106 ? add_553840 : sel_553837;
  assign add_553844 = sel_553841 + 8'h01;
  assign sel_553845 = array_index_553780 == array_index_537112 ? add_553844 : sel_553841;
  assign add_553848 = sel_553845 + 8'h01;
  assign sel_553849 = array_index_553780 == array_index_537118 ? add_553848 : sel_553845;
  assign add_553852 = sel_553849 + 8'h01;
  assign sel_553853 = array_index_553780 == array_index_537124 ? add_553852 : sel_553849;
  assign add_553856 = sel_553853 + 8'h01;
  assign sel_553857 = array_index_553780 == array_index_537130 ? add_553856 : sel_553853;
  assign add_553860 = sel_553857 + 8'h01;
  assign sel_553861 = array_index_553780 == array_index_537136 ? add_553860 : sel_553857;
  assign add_553864 = sel_553861 + 8'h01;
  assign sel_553865 = array_index_553780 == array_index_537142 ? add_553864 : sel_553861;
  assign add_553868 = sel_553865 + 8'h01;
  assign sel_553869 = array_index_553780 == array_index_537148 ? add_553868 : sel_553865;
  assign add_553872 = sel_553869 + 8'h01;
  assign sel_553873 = array_index_553780 == array_index_537154 ? add_553872 : sel_553869;
  assign add_553876 = sel_553873 + 8'h01;
  assign sel_553877 = array_index_553780 == array_index_537160 ? add_553876 : sel_553873;
  assign add_553880 = sel_553877 + 8'h01;
  assign sel_553881 = array_index_553780 == array_index_537166 ? add_553880 : sel_553877;
  assign add_553884 = sel_553881 + 8'h01;
  assign sel_553885 = array_index_553780 == array_index_537172 ? add_553884 : sel_553881;
  assign add_553888 = sel_553885 + 8'h01;
  assign sel_553889 = array_index_553780 == array_index_537178 ? add_553888 : sel_553885;
  assign add_553892 = sel_553889 + 8'h01;
  assign sel_553893 = array_index_553780 == array_index_537184 ? add_553892 : sel_553889;
  assign add_553896 = sel_553893 + 8'h01;
  assign sel_553897 = array_index_553780 == array_index_537190 ? add_553896 : sel_553893;
  assign add_553900 = sel_553897 + 8'h01;
  assign sel_553901 = array_index_553780 == array_index_537196 ? add_553900 : sel_553897;
  assign add_553904 = sel_553901 + 8'h01;
  assign sel_553905 = array_index_553780 == array_index_537202 ? add_553904 : sel_553901;
  assign add_553908 = sel_553905 + 8'h01;
  assign sel_553909 = array_index_553780 == array_index_537208 ? add_553908 : sel_553905;
  assign add_553912 = sel_553909 + 8'h01;
  assign sel_553913 = array_index_553780 == array_index_537214 ? add_553912 : sel_553909;
  assign add_553916 = sel_553913 + 8'h01;
  assign sel_553917 = array_index_553780 == array_index_537220 ? add_553916 : sel_553913;
  assign add_553920 = sel_553917 + 8'h01;
  assign sel_553921 = array_index_553780 == array_index_537226 ? add_553920 : sel_553917;
  assign add_553924 = sel_553921 + 8'h01;
  assign sel_553925 = array_index_553780 == array_index_537232 ? add_553924 : sel_553921;
  assign add_553928 = sel_553925 + 8'h01;
  assign sel_553929 = array_index_553780 == array_index_537238 ? add_553928 : sel_553925;
  assign add_553932 = sel_553929 + 8'h01;
  assign sel_553933 = array_index_553780 == array_index_537244 ? add_553932 : sel_553929;
  assign add_553936 = sel_553933 + 8'h01;
  assign sel_553937 = array_index_553780 == array_index_537250 ? add_553936 : sel_553933;
  assign add_553940 = sel_553937 + 8'h01;
  assign sel_553941 = array_index_553780 == array_index_537256 ? add_553940 : sel_553937;
  assign add_553944 = sel_553941 + 8'h01;
  assign sel_553945 = array_index_553780 == array_index_537262 ? add_553944 : sel_553941;
  assign add_553948 = sel_553945 + 8'h01;
  assign sel_553949 = array_index_553780 == array_index_537268 ? add_553948 : sel_553945;
  assign add_553952 = sel_553949 + 8'h01;
  assign sel_553953 = array_index_553780 == array_index_537274 ? add_553952 : sel_553949;
  assign add_553956 = sel_553953 + 8'h01;
  assign sel_553957 = array_index_553780 == array_index_537280 ? add_553956 : sel_553953;
  assign add_553960 = sel_553957 + 8'h01;
  assign sel_553961 = array_index_553780 == array_index_537286 ? add_553960 : sel_553957;
  assign add_553964 = sel_553961 + 8'h01;
  assign sel_553965 = array_index_553780 == array_index_537292 ? add_553964 : sel_553961;
  assign add_553968 = sel_553965 + 8'h01;
  assign sel_553969 = array_index_553780 == array_index_537298 ? add_553968 : sel_553965;
  assign add_553972 = sel_553969 + 8'h01;
  assign sel_553973 = array_index_553780 == array_index_537304 ? add_553972 : sel_553969;
  assign add_553976 = sel_553973 + 8'h01;
  assign sel_553977 = array_index_553780 == array_index_537310 ? add_553976 : sel_553973;
  assign add_553980 = sel_553977 + 8'h01;
  assign sel_553981 = array_index_553780 == array_index_537316 ? add_553980 : sel_553977;
  assign add_553984 = sel_553981 + 8'h01;
  assign sel_553985 = array_index_553780 == array_index_537322 ? add_553984 : sel_553981;
  assign add_553988 = sel_553985 + 8'h01;
  assign sel_553989 = array_index_553780 == array_index_537328 ? add_553988 : sel_553985;
  assign add_553992 = sel_553989 + 8'h01;
  assign sel_553993 = array_index_553780 == array_index_537334 ? add_553992 : sel_553989;
  assign add_553996 = sel_553993 + 8'h01;
  assign sel_553997 = array_index_553780 == array_index_537340 ? add_553996 : sel_553993;
  assign add_554000 = sel_553997 + 8'h01;
  assign sel_554001 = array_index_553780 == array_index_537346 ? add_554000 : sel_553997;
  assign add_554004 = sel_554001 + 8'h01;
  assign sel_554005 = array_index_553780 == array_index_537352 ? add_554004 : sel_554001;
  assign add_554008 = sel_554005 + 8'h01;
  assign sel_554009 = array_index_553780 == array_index_537358 ? add_554008 : sel_554005;
  assign add_554012 = sel_554009 + 8'h01;
  assign sel_554013 = array_index_553780 == array_index_537364 ? add_554012 : sel_554009;
  assign add_554016 = sel_554013 + 8'h01;
  assign sel_554017 = array_index_553780 == array_index_537370 ? add_554016 : sel_554013;
  assign add_554020 = sel_554017 + 8'h01;
  assign sel_554021 = array_index_553780 == array_index_537376 ? add_554020 : sel_554017;
  assign add_554024 = sel_554021 + 8'h01;
  assign sel_554025 = array_index_553780 == array_index_537382 ? add_554024 : sel_554021;
  assign add_554028 = sel_554025 + 8'h01;
  assign sel_554029 = array_index_553780 == array_index_537388 ? add_554028 : sel_554025;
  assign add_554032 = sel_554029 + 8'h01;
  assign sel_554033 = array_index_553780 == array_index_537394 ? add_554032 : sel_554029;
  assign add_554036 = sel_554033 + 8'h01;
  assign sel_554037 = array_index_553780 == array_index_537400 ? add_554036 : sel_554033;
  assign add_554040 = sel_554037 + 8'h01;
  assign sel_554041 = array_index_553780 == array_index_537406 ? add_554040 : sel_554037;
  assign add_554044 = sel_554041 + 8'h01;
  assign sel_554045 = array_index_553780 == array_index_537412 ? add_554044 : sel_554041;
  assign add_554048 = sel_554045 + 8'h01;
  assign sel_554049 = array_index_553780 == array_index_537418 ? add_554048 : sel_554045;
  assign add_554052 = sel_554049 + 8'h01;
  assign sel_554053 = array_index_553780 == array_index_537424 ? add_554052 : sel_554049;
  assign add_554056 = sel_554053 + 8'h01;
  assign sel_554057 = array_index_553780 == array_index_537430 ? add_554056 : sel_554053;
  assign add_554060 = sel_554057 + 8'h01;
  assign sel_554061 = array_index_553780 == array_index_537436 ? add_554060 : sel_554057;
  assign add_554064 = sel_554061 + 8'h01;
  assign sel_554065 = array_index_553780 == array_index_537442 ? add_554064 : sel_554061;
  assign add_554068 = sel_554065 + 8'h01;
  assign sel_554069 = array_index_553780 == array_index_537448 ? add_554068 : sel_554065;
  assign add_554072 = sel_554069 + 8'h01;
  assign sel_554073 = array_index_553780 == array_index_537454 ? add_554072 : sel_554069;
  assign add_554076 = sel_554073 + 8'h01;
  assign sel_554077 = array_index_553780 == array_index_537460 ? add_554076 : sel_554073;
  assign add_554081 = sel_554077 + 8'h01;
  assign array_index_554082 = set1_unflattened[7'h38];
  assign sel_554083 = array_index_553780 == array_index_537466 ? add_554081 : sel_554077;
  assign add_554086 = sel_554083 + 8'h01;
  assign sel_554087 = array_index_554082 == array_index_537012 ? add_554086 : sel_554083;
  assign add_554090 = sel_554087 + 8'h01;
  assign sel_554091 = array_index_554082 == array_index_537016 ? add_554090 : sel_554087;
  assign add_554094 = sel_554091 + 8'h01;
  assign sel_554095 = array_index_554082 == array_index_537024 ? add_554094 : sel_554091;
  assign add_554098 = sel_554095 + 8'h01;
  assign sel_554099 = array_index_554082 == array_index_537032 ? add_554098 : sel_554095;
  assign add_554102 = sel_554099 + 8'h01;
  assign sel_554103 = array_index_554082 == array_index_537040 ? add_554102 : sel_554099;
  assign add_554106 = sel_554103 + 8'h01;
  assign sel_554107 = array_index_554082 == array_index_537048 ? add_554106 : sel_554103;
  assign add_554110 = sel_554107 + 8'h01;
  assign sel_554111 = array_index_554082 == array_index_537056 ? add_554110 : sel_554107;
  assign add_554114 = sel_554111 + 8'h01;
  assign sel_554115 = array_index_554082 == array_index_537064 ? add_554114 : sel_554111;
  assign add_554118 = sel_554115 + 8'h01;
  assign sel_554119 = array_index_554082 == array_index_537070 ? add_554118 : sel_554115;
  assign add_554122 = sel_554119 + 8'h01;
  assign sel_554123 = array_index_554082 == array_index_537076 ? add_554122 : sel_554119;
  assign add_554126 = sel_554123 + 8'h01;
  assign sel_554127 = array_index_554082 == array_index_537082 ? add_554126 : sel_554123;
  assign add_554130 = sel_554127 + 8'h01;
  assign sel_554131 = array_index_554082 == array_index_537088 ? add_554130 : sel_554127;
  assign add_554134 = sel_554131 + 8'h01;
  assign sel_554135 = array_index_554082 == array_index_537094 ? add_554134 : sel_554131;
  assign add_554138 = sel_554135 + 8'h01;
  assign sel_554139 = array_index_554082 == array_index_537100 ? add_554138 : sel_554135;
  assign add_554142 = sel_554139 + 8'h01;
  assign sel_554143 = array_index_554082 == array_index_537106 ? add_554142 : sel_554139;
  assign add_554146 = sel_554143 + 8'h01;
  assign sel_554147 = array_index_554082 == array_index_537112 ? add_554146 : sel_554143;
  assign add_554150 = sel_554147 + 8'h01;
  assign sel_554151 = array_index_554082 == array_index_537118 ? add_554150 : sel_554147;
  assign add_554154 = sel_554151 + 8'h01;
  assign sel_554155 = array_index_554082 == array_index_537124 ? add_554154 : sel_554151;
  assign add_554158 = sel_554155 + 8'h01;
  assign sel_554159 = array_index_554082 == array_index_537130 ? add_554158 : sel_554155;
  assign add_554162 = sel_554159 + 8'h01;
  assign sel_554163 = array_index_554082 == array_index_537136 ? add_554162 : sel_554159;
  assign add_554166 = sel_554163 + 8'h01;
  assign sel_554167 = array_index_554082 == array_index_537142 ? add_554166 : sel_554163;
  assign add_554170 = sel_554167 + 8'h01;
  assign sel_554171 = array_index_554082 == array_index_537148 ? add_554170 : sel_554167;
  assign add_554174 = sel_554171 + 8'h01;
  assign sel_554175 = array_index_554082 == array_index_537154 ? add_554174 : sel_554171;
  assign add_554178 = sel_554175 + 8'h01;
  assign sel_554179 = array_index_554082 == array_index_537160 ? add_554178 : sel_554175;
  assign add_554182 = sel_554179 + 8'h01;
  assign sel_554183 = array_index_554082 == array_index_537166 ? add_554182 : sel_554179;
  assign add_554186 = sel_554183 + 8'h01;
  assign sel_554187 = array_index_554082 == array_index_537172 ? add_554186 : sel_554183;
  assign add_554190 = sel_554187 + 8'h01;
  assign sel_554191 = array_index_554082 == array_index_537178 ? add_554190 : sel_554187;
  assign add_554194 = sel_554191 + 8'h01;
  assign sel_554195 = array_index_554082 == array_index_537184 ? add_554194 : sel_554191;
  assign add_554198 = sel_554195 + 8'h01;
  assign sel_554199 = array_index_554082 == array_index_537190 ? add_554198 : sel_554195;
  assign add_554202 = sel_554199 + 8'h01;
  assign sel_554203 = array_index_554082 == array_index_537196 ? add_554202 : sel_554199;
  assign add_554206 = sel_554203 + 8'h01;
  assign sel_554207 = array_index_554082 == array_index_537202 ? add_554206 : sel_554203;
  assign add_554210 = sel_554207 + 8'h01;
  assign sel_554211 = array_index_554082 == array_index_537208 ? add_554210 : sel_554207;
  assign add_554214 = sel_554211 + 8'h01;
  assign sel_554215 = array_index_554082 == array_index_537214 ? add_554214 : sel_554211;
  assign add_554218 = sel_554215 + 8'h01;
  assign sel_554219 = array_index_554082 == array_index_537220 ? add_554218 : sel_554215;
  assign add_554222 = sel_554219 + 8'h01;
  assign sel_554223 = array_index_554082 == array_index_537226 ? add_554222 : sel_554219;
  assign add_554226 = sel_554223 + 8'h01;
  assign sel_554227 = array_index_554082 == array_index_537232 ? add_554226 : sel_554223;
  assign add_554230 = sel_554227 + 8'h01;
  assign sel_554231 = array_index_554082 == array_index_537238 ? add_554230 : sel_554227;
  assign add_554234 = sel_554231 + 8'h01;
  assign sel_554235 = array_index_554082 == array_index_537244 ? add_554234 : sel_554231;
  assign add_554238 = sel_554235 + 8'h01;
  assign sel_554239 = array_index_554082 == array_index_537250 ? add_554238 : sel_554235;
  assign add_554242 = sel_554239 + 8'h01;
  assign sel_554243 = array_index_554082 == array_index_537256 ? add_554242 : sel_554239;
  assign add_554246 = sel_554243 + 8'h01;
  assign sel_554247 = array_index_554082 == array_index_537262 ? add_554246 : sel_554243;
  assign add_554250 = sel_554247 + 8'h01;
  assign sel_554251 = array_index_554082 == array_index_537268 ? add_554250 : sel_554247;
  assign add_554254 = sel_554251 + 8'h01;
  assign sel_554255 = array_index_554082 == array_index_537274 ? add_554254 : sel_554251;
  assign add_554258 = sel_554255 + 8'h01;
  assign sel_554259 = array_index_554082 == array_index_537280 ? add_554258 : sel_554255;
  assign add_554262 = sel_554259 + 8'h01;
  assign sel_554263 = array_index_554082 == array_index_537286 ? add_554262 : sel_554259;
  assign add_554266 = sel_554263 + 8'h01;
  assign sel_554267 = array_index_554082 == array_index_537292 ? add_554266 : sel_554263;
  assign add_554270 = sel_554267 + 8'h01;
  assign sel_554271 = array_index_554082 == array_index_537298 ? add_554270 : sel_554267;
  assign add_554274 = sel_554271 + 8'h01;
  assign sel_554275 = array_index_554082 == array_index_537304 ? add_554274 : sel_554271;
  assign add_554278 = sel_554275 + 8'h01;
  assign sel_554279 = array_index_554082 == array_index_537310 ? add_554278 : sel_554275;
  assign add_554282 = sel_554279 + 8'h01;
  assign sel_554283 = array_index_554082 == array_index_537316 ? add_554282 : sel_554279;
  assign add_554286 = sel_554283 + 8'h01;
  assign sel_554287 = array_index_554082 == array_index_537322 ? add_554286 : sel_554283;
  assign add_554290 = sel_554287 + 8'h01;
  assign sel_554291 = array_index_554082 == array_index_537328 ? add_554290 : sel_554287;
  assign add_554294 = sel_554291 + 8'h01;
  assign sel_554295 = array_index_554082 == array_index_537334 ? add_554294 : sel_554291;
  assign add_554298 = sel_554295 + 8'h01;
  assign sel_554299 = array_index_554082 == array_index_537340 ? add_554298 : sel_554295;
  assign add_554302 = sel_554299 + 8'h01;
  assign sel_554303 = array_index_554082 == array_index_537346 ? add_554302 : sel_554299;
  assign add_554306 = sel_554303 + 8'h01;
  assign sel_554307 = array_index_554082 == array_index_537352 ? add_554306 : sel_554303;
  assign add_554310 = sel_554307 + 8'h01;
  assign sel_554311 = array_index_554082 == array_index_537358 ? add_554310 : sel_554307;
  assign add_554314 = sel_554311 + 8'h01;
  assign sel_554315 = array_index_554082 == array_index_537364 ? add_554314 : sel_554311;
  assign add_554318 = sel_554315 + 8'h01;
  assign sel_554319 = array_index_554082 == array_index_537370 ? add_554318 : sel_554315;
  assign add_554322 = sel_554319 + 8'h01;
  assign sel_554323 = array_index_554082 == array_index_537376 ? add_554322 : sel_554319;
  assign add_554326 = sel_554323 + 8'h01;
  assign sel_554327 = array_index_554082 == array_index_537382 ? add_554326 : sel_554323;
  assign add_554330 = sel_554327 + 8'h01;
  assign sel_554331 = array_index_554082 == array_index_537388 ? add_554330 : sel_554327;
  assign add_554334 = sel_554331 + 8'h01;
  assign sel_554335 = array_index_554082 == array_index_537394 ? add_554334 : sel_554331;
  assign add_554338 = sel_554335 + 8'h01;
  assign sel_554339 = array_index_554082 == array_index_537400 ? add_554338 : sel_554335;
  assign add_554342 = sel_554339 + 8'h01;
  assign sel_554343 = array_index_554082 == array_index_537406 ? add_554342 : sel_554339;
  assign add_554346 = sel_554343 + 8'h01;
  assign sel_554347 = array_index_554082 == array_index_537412 ? add_554346 : sel_554343;
  assign add_554350 = sel_554347 + 8'h01;
  assign sel_554351 = array_index_554082 == array_index_537418 ? add_554350 : sel_554347;
  assign add_554354 = sel_554351 + 8'h01;
  assign sel_554355 = array_index_554082 == array_index_537424 ? add_554354 : sel_554351;
  assign add_554358 = sel_554355 + 8'h01;
  assign sel_554359 = array_index_554082 == array_index_537430 ? add_554358 : sel_554355;
  assign add_554362 = sel_554359 + 8'h01;
  assign sel_554363 = array_index_554082 == array_index_537436 ? add_554362 : sel_554359;
  assign add_554366 = sel_554363 + 8'h01;
  assign sel_554367 = array_index_554082 == array_index_537442 ? add_554366 : sel_554363;
  assign add_554370 = sel_554367 + 8'h01;
  assign sel_554371 = array_index_554082 == array_index_537448 ? add_554370 : sel_554367;
  assign add_554374 = sel_554371 + 8'h01;
  assign sel_554375 = array_index_554082 == array_index_537454 ? add_554374 : sel_554371;
  assign add_554378 = sel_554375 + 8'h01;
  assign sel_554379 = array_index_554082 == array_index_537460 ? add_554378 : sel_554375;
  assign add_554383 = sel_554379 + 8'h01;
  assign array_index_554384 = set1_unflattened[7'h39];
  assign sel_554385 = array_index_554082 == array_index_537466 ? add_554383 : sel_554379;
  assign add_554388 = sel_554385 + 8'h01;
  assign sel_554389 = array_index_554384 == array_index_537012 ? add_554388 : sel_554385;
  assign add_554392 = sel_554389 + 8'h01;
  assign sel_554393 = array_index_554384 == array_index_537016 ? add_554392 : sel_554389;
  assign add_554396 = sel_554393 + 8'h01;
  assign sel_554397 = array_index_554384 == array_index_537024 ? add_554396 : sel_554393;
  assign add_554400 = sel_554397 + 8'h01;
  assign sel_554401 = array_index_554384 == array_index_537032 ? add_554400 : sel_554397;
  assign add_554404 = sel_554401 + 8'h01;
  assign sel_554405 = array_index_554384 == array_index_537040 ? add_554404 : sel_554401;
  assign add_554408 = sel_554405 + 8'h01;
  assign sel_554409 = array_index_554384 == array_index_537048 ? add_554408 : sel_554405;
  assign add_554412 = sel_554409 + 8'h01;
  assign sel_554413 = array_index_554384 == array_index_537056 ? add_554412 : sel_554409;
  assign add_554416 = sel_554413 + 8'h01;
  assign sel_554417 = array_index_554384 == array_index_537064 ? add_554416 : sel_554413;
  assign add_554420 = sel_554417 + 8'h01;
  assign sel_554421 = array_index_554384 == array_index_537070 ? add_554420 : sel_554417;
  assign add_554424 = sel_554421 + 8'h01;
  assign sel_554425 = array_index_554384 == array_index_537076 ? add_554424 : sel_554421;
  assign add_554428 = sel_554425 + 8'h01;
  assign sel_554429 = array_index_554384 == array_index_537082 ? add_554428 : sel_554425;
  assign add_554432 = sel_554429 + 8'h01;
  assign sel_554433 = array_index_554384 == array_index_537088 ? add_554432 : sel_554429;
  assign add_554436 = sel_554433 + 8'h01;
  assign sel_554437 = array_index_554384 == array_index_537094 ? add_554436 : sel_554433;
  assign add_554440 = sel_554437 + 8'h01;
  assign sel_554441 = array_index_554384 == array_index_537100 ? add_554440 : sel_554437;
  assign add_554444 = sel_554441 + 8'h01;
  assign sel_554445 = array_index_554384 == array_index_537106 ? add_554444 : sel_554441;
  assign add_554448 = sel_554445 + 8'h01;
  assign sel_554449 = array_index_554384 == array_index_537112 ? add_554448 : sel_554445;
  assign add_554452 = sel_554449 + 8'h01;
  assign sel_554453 = array_index_554384 == array_index_537118 ? add_554452 : sel_554449;
  assign add_554456 = sel_554453 + 8'h01;
  assign sel_554457 = array_index_554384 == array_index_537124 ? add_554456 : sel_554453;
  assign add_554460 = sel_554457 + 8'h01;
  assign sel_554461 = array_index_554384 == array_index_537130 ? add_554460 : sel_554457;
  assign add_554464 = sel_554461 + 8'h01;
  assign sel_554465 = array_index_554384 == array_index_537136 ? add_554464 : sel_554461;
  assign add_554468 = sel_554465 + 8'h01;
  assign sel_554469 = array_index_554384 == array_index_537142 ? add_554468 : sel_554465;
  assign add_554472 = sel_554469 + 8'h01;
  assign sel_554473 = array_index_554384 == array_index_537148 ? add_554472 : sel_554469;
  assign add_554476 = sel_554473 + 8'h01;
  assign sel_554477 = array_index_554384 == array_index_537154 ? add_554476 : sel_554473;
  assign add_554480 = sel_554477 + 8'h01;
  assign sel_554481 = array_index_554384 == array_index_537160 ? add_554480 : sel_554477;
  assign add_554484 = sel_554481 + 8'h01;
  assign sel_554485 = array_index_554384 == array_index_537166 ? add_554484 : sel_554481;
  assign add_554488 = sel_554485 + 8'h01;
  assign sel_554489 = array_index_554384 == array_index_537172 ? add_554488 : sel_554485;
  assign add_554492 = sel_554489 + 8'h01;
  assign sel_554493 = array_index_554384 == array_index_537178 ? add_554492 : sel_554489;
  assign add_554496 = sel_554493 + 8'h01;
  assign sel_554497 = array_index_554384 == array_index_537184 ? add_554496 : sel_554493;
  assign add_554500 = sel_554497 + 8'h01;
  assign sel_554501 = array_index_554384 == array_index_537190 ? add_554500 : sel_554497;
  assign add_554504 = sel_554501 + 8'h01;
  assign sel_554505 = array_index_554384 == array_index_537196 ? add_554504 : sel_554501;
  assign add_554508 = sel_554505 + 8'h01;
  assign sel_554509 = array_index_554384 == array_index_537202 ? add_554508 : sel_554505;
  assign add_554512 = sel_554509 + 8'h01;
  assign sel_554513 = array_index_554384 == array_index_537208 ? add_554512 : sel_554509;
  assign add_554516 = sel_554513 + 8'h01;
  assign sel_554517 = array_index_554384 == array_index_537214 ? add_554516 : sel_554513;
  assign add_554520 = sel_554517 + 8'h01;
  assign sel_554521 = array_index_554384 == array_index_537220 ? add_554520 : sel_554517;
  assign add_554524 = sel_554521 + 8'h01;
  assign sel_554525 = array_index_554384 == array_index_537226 ? add_554524 : sel_554521;
  assign add_554528 = sel_554525 + 8'h01;
  assign sel_554529 = array_index_554384 == array_index_537232 ? add_554528 : sel_554525;
  assign add_554532 = sel_554529 + 8'h01;
  assign sel_554533 = array_index_554384 == array_index_537238 ? add_554532 : sel_554529;
  assign add_554536 = sel_554533 + 8'h01;
  assign sel_554537 = array_index_554384 == array_index_537244 ? add_554536 : sel_554533;
  assign add_554540 = sel_554537 + 8'h01;
  assign sel_554541 = array_index_554384 == array_index_537250 ? add_554540 : sel_554537;
  assign add_554544 = sel_554541 + 8'h01;
  assign sel_554545 = array_index_554384 == array_index_537256 ? add_554544 : sel_554541;
  assign add_554548 = sel_554545 + 8'h01;
  assign sel_554549 = array_index_554384 == array_index_537262 ? add_554548 : sel_554545;
  assign add_554552 = sel_554549 + 8'h01;
  assign sel_554553 = array_index_554384 == array_index_537268 ? add_554552 : sel_554549;
  assign add_554556 = sel_554553 + 8'h01;
  assign sel_554557 = array_index_554384 == array_index_537274 ? add_554556 : sel_554553;
  assign add_554560 = sel_554557 + 8'h01;
  assign sel_554561 = array_index_554384 == array_index_537280 ? add_554560 : sel_554557;
  assign add_554564 = sel_554561 + 8'h01;
  assign sel_554565 = array_index_554384 == array_index_537286 ? add_554564 : sel_554561;
  assign add_554568 = sel_554565 + 8'h01;
  assign sel_554569 = array_index_554384 == array_index_537292 ? add_554568 : sel_554565;
  assign add_554572 = sel_554569 + 8'h01;
  assign sel_554573 = array_index_554384 == array_index_537298 ? add_554572 : sel_554569;
  assign add_554576 = sel_554573 + 8'h01;
  assign sel_554577 = array_index_554384 == array_index_537304 ? add_554576 : sel_554573;
  assign add_554580 = sel_554577 + 8'h01;
  assign sel_554581 = array_index_554384 == array_index_537310 ? add_554580 : sel_554577;
  assign add_554584 = sel_554581 + 8'h01;
  assign sel_554585 = array_index_554384 == array_index_537316 ? add_554584 : sel_554581;
  assign add_554588 = sel_554585 + 8'h01;
  assign sel_554589 = array_index_554384 == array_index_537322 ? add_554588 : sel_554585;
  assign add_554592 = sel_554589 + 8'h01;
  assign sel_554593 = array_index_554384 == array_index_537328 ? add_554592 : sel_554589;
  assign add_554596 = sel_554593 + 8'h01;
  assign sel_554597 = array_index_554384 == array_index_537334 ? add_554596 : sel_554593;
  assign add_554600 = sel_554597 + 8'h01;
  assign sel_554601 = array_index_554384 == array_index_537340 ? add_554600 : sel_554597;
  assign add_554604 = sel_554601 + 8'h01;
  assign sel_554605 = array_index_554384 == array_index_537346 ? add_554604 : sel_554601;
  assign add_554608 = sel_554605 + 8'h01;
  assign sel_554609 = array_index_554384 == array_index_537352 ? add_554608 : sel_554605;
  assign add_554612 = sel_554609 + 8'h01;
  assign sel_554613 = array_index_554384 == array_index_537358 ? add_554612 : sel_554609;
  assign add_554616 = sel_554613 + 8'h01;
  assign sel_554617 = array_index_554384 == array_index_537364 ? add_554616 : sel_554613;
  assign add_554620 = sel_554617 + 8'h01;
  assign sel_554621 = array_index_554384 == array_index_537370 ? add_554620 : sel_554617;
  assign add_554624 = sel_554621 + 8'h01;
  assign sel_554625 = array_index_554384 == array_index_537376 ? add_554624 : sel_554621;
  assign add_554628 = sel_554625 + 8'h01;
  assign sel_554629 = array_index_554384 == array_index_537382 ? add_554628 : sel_554625;
  assign add_554632 = sel_554629 + 8'h01;
  assign sel_554633 = array_index_554384 == array_index_537388 ? add_554632 : sel_554629;
  assign add_554636 = sel_554633 + 8'h01;
  assign sel_554637 = array_index_554384 == array_index_537394 ? add_554636 : sel_554633;
  assign add_554640 = sel_554637 + 8'h01;
  assign sel_554641 = array_index_554384 == array_index_537400 ? add_554640 : sel_554637;
  assign add_554644 = sel_554641 + 8'h01;
  assign sel_554645 = array_index_554384 == array_index_537406 ? add_554644 : sel_554641;
  assign add_554648 = sel_554645 + 8'h01;
  assign sel_554649 = array_index_554384 == array_index_537412 ? add_554648 : sel_554645;
  assign add_554652 = sel_554649 + 8'h01;
  assign sel_554653 = array_index_554384 == array_index_537418 ? add_554652 : sel_554649;
  assign add_554656 = sel_554653 + 8'h01;
  assign sel_554657 = array_index_554384 == array_index_537424 ? add_554656 : sel_554653;
  assign add_554660 = sel_554657 + 8'h01;
  assign sel_554661 = array_index_554384 == array_index_537430 ? add_554660 : sel_554657;
  assign add_554664 = sel_554661 + 8'h01;
  assign sel_554665 = array_index_554384 == array_index_537436 ? add_554664 : sel_554661;
  assign add_554668 = sel_554665 + 8'h01;
  assign sel_554669 = array_index_554384 == array_index_537442 ? add_554668 : sel_554665;
  assign add_554672 = sel_554669 + 8'h01;
  assign sel_554673 = array_index_554384 == array_index_537448 ? add_554672 : sel_554669;
  assign add_554676 = sel_554673 + 8'h01;
  assign sel_554677 = array_index_554384 == array_index_537454 ? add_554676 : sel_554673;
  assign add_554680 = sel_554677 + 8'h01;
  assign sel_554681 = array_index_554384 == array_index_537460 ? add_554680 : sel_554677;
  assign add_554685 = sel_554681 + 8'h01;
  assign array_index_554686 = set1_unflattened[7'h3a];
  assign sel_554687 = array_index_554384 == array_index_537466 ? add_554685 : sel_554681;
  assign add_554690 = sel_554687 + 8'h01;
  assign sel_554691 = array_index_554686 == array_index_537012 ? add_554690 : sel_554687;
  assign add_554694 = sel_554691 + 8'h01;
  assign sel_554695 = array_index_554686 == array_index_537016 ? add_554694 : sel_554691;
  assign add_554698 = sel_554695 + 8'h01;
  assign sel_554699 = array_index_554686 == array_index_537024 ? add_554698 : sel_554695;
  assign add_554702 = sel_554699 + 8'h01;
  assign sel_554703 = array_index_554686 == array_index_537032 ? add_554702 : sel_554699;
  assign add_554706 = sel_554703 + 8'h01;
  assign sel_554707 = array_index_554686 == array_index_537040 ? add_554706 : sel_554703;
  assign add_554710 = sel_554707 + 8'h01;
  assign sel_554711 = array_index_554686 == array_index_537048 ? add_554710 : sel_554707;
  assign add_554714 = sel_554711 + 8'h01;
  assign sel_554715 = array_index_554686 == array_index_537056 ? add_554714 : sel_554711;
  assign add_554718 = sel_554715 + 8'h01;
  assign sel_554719 = array_index_554686 == array_index_537064 ? add_554718 : sel_554715;
  assign add_554722 = sel_554719 + 8'h01;
  assign sel_554723 = array_index_554686 == array_index_537070 ? add_554722 : sel_554719;
  assign add_554726 = sel_554723 + 8'h01;
  assign sel_554727 = array_index_554686 == array_index_537076 ? add_554726 : sel_554723;
  assign add_554730 = sel_554727 + 8'h01;
  assign sel_554731 = array_index_554686 == array_index_537082 ? add_554730 : sel_554727;
  assign add_554734 = sel_554731 + 8'h01;
  assign sel_554735 = array_index_554686 == array_index_537088 ? add_554734 : sel_554731;
  assign add_554738 = sel_554735 + 8'h01;
  assign sel_554739 = array_index_554686 == array_index_537094 ? add_554738 : sel_554735;
  assign add_554742 = sel_554739 + 8'h01;
  assign sel_554743 = array_index_554686 == array_index_537100 ? add_554742 : sel_554739;
  assign add_554746 = sel_554743 + 8'h01;
  assign sel_554747 = array_index_554686 == array_index_537106 ? add_554746 : sel_554743;
  assign add_554750 = sel_554747 + 8'h01;
  assign sel_554751 = array_index_554686 == array_index_537112 ? add_554750 : sel_554747;
  assign add_554754 = sel_554751 + 8'h01;
  assign sel_554755 = array_index_554686 == array_index_537118 ? add_554754 : sel_554751;
  assign add_554758 = sel_554755 + 8'h01;
  assign sel_554759 = array_index_554686 == array_index_537124 ? add_554758 : sel_554755;
  assign add_554762 = sel_554759 + 8'h01;
  assign sel_554763 = array_index_554686 == array_index_537130 ? add_554762 : sel_554759;
  assign add_554766 = sel_554763 + 8'h01;
  assign sel_554767 = array_index_554686 == array_index_537136 ? add_554766 : sel_554763;
  assign add_554770 = sel_554767 + 8'h01;
  assign sel_554771 = array_index_554686 == array_index_537142 ? add_554770 : sel_554767;
  assign add_554774 = sel_554771 + 8'h01;
  assign sel_554775 = array_index_554686 == array_index_537148 ? add_554774 : sel_554771;
  assign add_554778 = sel_554775 + 8'h01;
  assign sel_554779 = array_index_554686 == array_index_537154 ? add_554778 : sel_554775;
  assign add_554782 = sel_554779 + 8'h01;
  assign sel_554783 = array_index_554686 == array_index_537160 ? add_554782 : sel_554779;
  assign add_554786 = sel_554783 + 8'h01;
  assign sel_554787 = array_index_554686 == array_index_537166 ? add_554786 : sel_554783;
  assign add_554790 = sel_554787 + 8'h01;
  assign sel_554791 = array_index_554686 == array_index_537172 ? add_554790 : sel_554787;
  assign add_554794 = sel_554791 + 8'h01;
  assign sel_554795 = array_index_554686 == array_index_537178 ? add_554794 : sel_554791;
  assign add_554798 = sel_554795 + 8'h01;
  assign sel_554799 = array_index_554686 == array_index_537184 ? add_554798 : sel_554795;
  assign add_554802 = sel_554799 + 8'h01;
  assign sel_554803 = array_index_554686 == array_index_537190 ? add_554802 : sel_554799;
  assign add_554806 = sel_554803 + 8'h01;
  assign sel_554807 = array_index_554686 == array_index_537196 ? add_554806 : sel_554803;
  assign add_554810 = sel_554807 + 8'h01;
  assign sel_554811 = array_index_554686 == array_index_537202 ? add_554810 : sel_554807;
  assign add_554814 = sel_554811 + 8'h01;
  assign sel_554815 = array_index_554686 == array_index_537208 ? add_554814 : sel_554811;
  assign add_554818 = sel_554815 + 8'h01;
  assign sel_554819 = array_index_554686 == array_index_537214 ? add_554818 : sel_554815;
  assign add_554822 = sel_554819 + 8'h01;
  assign sel_554823 = array_index_554686 == array_index_537220 ? add_554822 : sel_554819;
  assign add_554826 = sel_554823 + 8'h01;
  assign sel_554827 = array_index_554686 == array_index_537226 ? add_554826 : sel_554823;
  assign add_554830 = sel_554827 + 8'h01;
  assign sel_554831 = array_index_554686 == array_index_537232 ? add_554830 : sel_554827;
  assign add_554834 = sel_554831 + 8'h01;
  assign sel_554835 = array_index_554686 == array_index_537238 ? add_554834 : sel_554831;
  assign add_554838 = sel_554835 + 8'h01;
  assign sel_554839 = array_index_554686 == array_index_537244 ? add_554838 : sel_554835;
  assign add_554842 = sel_554839 + 8'h01;
  assign sel_554843 = array_index_554686 == array_index_537250 ? add_554842 : sel_554839;
  assign add_554846 = sel_554843 + 8'h01;
  assign sel_554847 = array_index_554686 == array_index_537256 ? add_554846 : sel_554843;
  assign add_554850 = sel_554847 + 8'h01;
  assign sel_554851 = array_index_554686 == array_index_537262 ? add_554850 : sel_554847;
  assign add_554854 = sel_554851 + 8'h01;
  assign sel_554855 = array_index_554686 == array_index_537268 ? add_554854 : sel_554851;
  assign add_554858 = sel_554855 + 8'h01;
  assign sel_554859 = array_index_554686 == array_index_537274 ? add_554858 : sel_554855;
  assign add_554862 = sel_554859 + 8'h01;
  assign sel_554863 = array_index_554686 == array_index_537280 ? add_554862 : sel_554859;
  assign add_554866 = sel_554863 + 8'h01;
  assign sel_554867 = array_index_554686 == array_index_537286 ? add_554866 : sel_554863;
  assign add_554870 = sel_554867 + 8'h01;
  assign sel_554871 = array_index_554686 == array_index_537292 ? add_554870 : sel_554867;
  assign add_554874 = sel_554871 + 8'h01;
  assign sel_554875 = array_index_554686 == array_index_537298 ? add_554874 : sel_554871;
  assign add_554878 = sel_554875 + 8'h01;
  assign sel_554879 = array_index_554686 == array_index_537304 ? add_554878 : sel_554875;
  assign add_554882 = sel_554879 + 8'h01;
  assign sel_554883 = array_index_554686 == array_index_537310 ? add_554882 : sel_554879;
  assign add_554886 = sel_554883 + 8'h01;
  assign sel_554887 = array_index_554686 == array_index_537316 ? add_554886 : sel_554883;
  assign add_554890 = sel_554887 + 8'h01;
  assign sel_554891 = array_index_554686 == array_index_537322 ? add_554890 : sel_554887;
  assign add_554894 = sel_554891 + 8'h01;
  assign sel_554895 = array_index_554686 == array_index_537328 ? add_554894 : sel_554891;
  assign add_554898 = sel_554895 + 8'h01;
  assign sel_554899 = array_index_554686 == array_index_537334 ? add_554898 : sel_554895;
  assign add_554902 = sel_554899 + 8'h01;
  assign sel_554903 = array_index_554686 == array_index_537340 ? add_554902 : sel_554899;
  assign add_554906 = sel_554903 + 8'h01;
  assign sel_554907 = array_index_554686 == array_index_537346 ? add_554906 : sel_554903;
  assign add_554910 = sel_554907 + 8'h01;
  assign sel_554911 = array_index_554686 == array_index_537352 ? add_554910 : sel_554907;
  assign add_554914 = sel_554911 + 8'h01;
  assign sel_554915 = array_index_554686 == array_index_537358 ? add_554914 : sel_554911;
  assign add_554918 = sel_554915 + 8'h01;
  assign sel_554919 = array_index_554686 == array_index_537364 ? add_554918 : sel_554915;
  assign add_554922 = sel_554919 + 8'h01;
  assign sel_554923 = array_index_554686 == array_index_537370 ? add_554922 : sel_554919;
  assign add_554926 = sel_554923 + 8'h01;
  assign sel_554927 = array_index_554686 == array_index_537376 ? add_554926 : sel_554923;
  assign add_554930 = sel_554927 + 8'h01;
  assign sel_554931 = array_index_554686 == array_index_537382 ? add_554930 : sel_554927;
  assign add_554934 = sel_554931 + 8'h01;
  assign sel_554935 = array_index_554686 == array_index_537388 ? add_554934 : sel_554931;
  assign add_554938 = sel_554935 + 8'h01;
  assign sel_554939 = array_index_554686 == array_index_537394 ? add_554938 : sel_554935;
  assign add_554942 = sel_554939 + 8'h01;
  assign sel_554943 = array_index_554686 == array_index_537400 ? add_554942 : sel_554939;
  assign add_554946 = sel_554943 + 8'h01;
  assign sel_554947 = array_index_554686 == array_index_537406 ? add_554946 : sel_554943;
  assign add_554950 = sel_554947 + 8'h01;
  assign sel_554951 = array_index_554686 == array_index_537412 ? add_554950 : sel_554947;
  assign add_554954 = sel_554951 + 8'h01;
  assign sel_554955 = array_index_554686 == array_index_537418 ? add_554954 : sel_554951;
  assign add_554958 = sel_554955 + 8'h01;
  assign sel_554959 = array_index_554686 == array_index_537424 ? add_554958 : sel_554955;
  assign add_554962 = sel_554959 + 8'h01;
  assign sel_554963 = array_index_554686 == array_index_537430 ? add_554962 : sel_554959;
  assign add_554966 = sel_554963 + 8'h01;
  assign sel_554967 = array_index_554686 == array_index_537436 ? add_554966 : sel_554963;
  assign add_554970 = sel_554967 + 8'h01;
  assign sel_554971 = array_index_554686 == array_index_537442 ? add_554970 : sel_554967;
  assign add_554974 = sel_554971 + 8'h01;
  assign sel_554975 = array_index_554686 == array_index_537448 ? add_554974 : sel_554971;
  assign add_554978 = sel_554975 + 8'h01;
  assign sel_554979 = array_index_554686 == array_index_537454 ? add_554978 : sel_554975;
  assign add_554982 = sel_554979 + 8'h01;
  assign sel_554983 = array_index_554686 == array_index_537460 ? add_554982 : sel_554979;
  assign add_554987 = sel_554983 + 8'h01;
  assign array_index_554988 = set1_unflattened[7'h3b];
  assign sel_554989 = array_index_554686 == array_index_537466 ? add_554987 : sel_554983;
  assign add_554992 = sel_554989 + 8'h01;
  assign sel_554993 = array_index_554988 == array_index_537012 ? add_554992 : sel_554989;
  assign add_554996 = sel_554993 + 8'h01;
  assign sel_554997 = array_index_554988 == array_index_537016 ? add_554996 : sel_554993;
  assign add_555000 = sel_554997 + 8'h01;
  assign sel_555001 = array_index_554988 == array_index_537024 ? add_555000 : sel_554997;
  assign add_555004 = sel_555001 + 8'h01;
  assign sel_555005 = array_index_554988 == array_index_537032 ? add_555004 : sel_555001;
  assign add_555008 = sel_555005 + 8'h01;
  assign sel_555009 = array_index_554988 == array_index_537040 ? add_555008 : sel_555005;
  assign add_555012 = sel_555009 + 8'h01;
  assign sel_555013 = array_index_554988 == array_index_537048 ? add_555012 : sel_555009;
  assign add_555016 = sel_555013 + 8'h01;
  assign sel_555017 = array_index_554988 == array_index_537056 ? add_555016 : sel_555013;
  assign add_555020 = sel_555017 + 8'h01;
  assign sel_555021 = array_index_554988 == array_index_537064 ? add_555020 : sel_555017;
  assign add_555024 = sel_555021 + 8'h01;
  assign sel_555025 = array_index_554988 == array_index_537070 ? add_555024 : sel_555021;
  assign add_555028 = sel_555025 + 8'h01;
  assign sel_555029 = array_index_554988 == array_index_537076 ? add_555028 : sel_555025;
  assign add_555032 = sel_555029 + 8'h01;
  assign sel_555033 = array_index_554988 == array_index_537082 ? add_555032 : sel_555029;
  assign add_555036 = sel_555033 + 8'h01;
  assign sel_555037 = array_index_554988 == array_index_537088 ? add_555036 : sel_555033;
  assign add_555040 = sel_555037 + 8'h01;
  assign sel_555041 = array_index_554988 == array_index_537094 ? add_555040 : sel_555037;
  assign add_555044 = sel_555041 + 8'h01;
  assign sel_555045 = array_index_554988 == array_index_537100 ? add_555044 : sel_555041;
  assign add_555048 = sel_555045 + 8'h01;
  assign sel_555049 = array_index_554988 == array_index_537106 ? add_555048 : sel_555045;
  assign add_555052 = sel_555049 + 8'h01;
  assign sel_555053 = array_index_554988 == array_index_537112 ? add_555052 : sel_555049;
  assign add_555056 = sel_555053 + 8'h01;
  assign sel_555057 = array_index_554988 == array_index_537118 ? add_555056 : sel_555053;
  assign add_555060 = sel_555057 + 8'h01;
  assign sel_555061 = array_index_554988 == array_index_537124 ? add_555060 : sel_555057;
  assign add_555064 = sel_555061 + 8'h01;
  assign sel_555065 = array_index_554988 == array_index_537130 ? add_555064 : sel_555061;
  assign add_555068 = sel_555065 + 8'h01;
  assign sel_555069 = array_index_554988 == array_index_537136 ? add_555068 : sel_555065;
  assign add_555072 = sel_555069 + 8'h01;
  assign sel_555073 = array_index_554988 == array_index_537142 ? add_555072 : sel_555069;
  assign add_555076 = sel_555073 + 8'h01;
  assign sel_555077 = array_index_554988 == array_index_537148 ? add_555076 : sel_555073;
  assign add_555080 = sel_555077 + 8'h01;
  assign sel_555081 = array_index_554988 == array_index_537154 ? add_555080 : sel_555077;
  assign add_555084 = sel_555081 + 8'h01;
  assign sel_555085 = array_index_554988 == array_index_537160 ? add_555084 : sel_555081;
  assign add_555088 = sel_555085 + 8'h01;
  assign sel_555089 = array_index_554988 == array_index_537166 ? add_555088 : sel_555085;
  assign add_555092 = sel_555089 + 8'h01;
  assign sel_555093 = array_index_554988 == array_index_537172 ? add_555092 : sel_555089;
  assign add_555096 = sel_555093 + 8'h01;
  assign sel_555097 = array_index_554988 == array_index_537178 ? add_555096 : sel_555093;
  assign add_555100 = sel_555097 + 8'h01;
  assign sel_555101 = array_index_554988 == array_index_537184 ? add_555100 : sel_555097;
  assign add_555104 = sel_555101 + 8'h01;
  assign sel_555105 = array_index_554988 == array_index_537190 ? add_555104 : sel_555101;
  assign add_555108 = sel_555105 + 8'h01;
  assign sel_555109 = array_index_554988 == array_index_537196 ? add_555108 : sel_555105;
  assign add_555112 = sel_555109 + 8'h01;
  assign sel_555113 = array_index_554988 == array_index_537202 ? add_555112 : sel_555109;
  assign add_555116 = sel_555113 + 8'h01;
  assign sel_555117 = array_index_554988 == array_index_537208 ? add_555116 : sel_555113;
  assign add_555120 = sel_555117 + 8'h01;
  assign sel_555121 = array_index_554988 == array_index_537214 ? add_555120 : sel_555117;
  assign add_555124 = sel_555121 + 8'h01;
  assign sel_555125 = array_index_554988 == array_index_537220 ? add_555124 : sel_555121;
  assign add_555128 = sel_555125 + 8'h01;
  assign sel_555129 = array_index_554988 == array_index_537226 ? add_555128 : sel_555125;
  assign add_555132 = sel_555129 + 8'h01;
  assign sel_555133 = array_index_554988 == array_index_537232 ? add_555132 : sel_555129;
  assign add_555136 = sel_555133 + 8'h01;
  assign sel_555137 = array_index_554988 == array_index_537238 ? add_555136 : sel_555133;
  assign add_555140 = sel_555137 + 8'h01;
  assign sel_555141 = array_index_554988 == array_index_537244 ? add_555140 : sel_555137;
  assign add_555144 = sel_555141 + 8'h01;
  assign sel_555145 = array_index_554988 == array_index_537250 ? add_555144 : sel_555141;
  assign add_555148 = sel_555145 + 8'h01;
  assign sel_555149 = array_index_554988 == array_index_537256 ? add_555148 : sel_555145;
  assign add_555152 = sel_555149 + 8'h01;
  assign sel_555153 = array_index_554988 == array_index_537262 ? add_555152 : sel_555149;
  assign add_555156 = sel_555153 + 8'h01;
  assign sel_555157 = array_index_554988 == array_index_537268 ? add_555156 : sel_555153;
  assign add_555160 = sel_555157 + 8'h01;
  assign sel_555161 = array_index_554988 == array_index_537274 ? add_555160 : sel_555157;
  assign add_555164 = sel_555161 + 8'h01;
  assign sel_555165 = array_index_554988 == array_index_537280 ? add_555164 : sel_555161;
  assign add_555168 = sel_555165 + 8'h01;
  assign sel_555169 = array_index_554988 == array_index_537286 ? add_555168 : sel_555165;
  assign add_555172 = sel_555169 + 8'h01;
  assign sel_555173 = array_index_554988 == array_index_537292 ? add_555172 : sel_555169;
  assign add_555176 = sel_555173 + 8'h01;
  assign sel_555177 = array_index_554988 == array_index_537298 ? add_555176 : sel_555173;
  assign add_555180 = sel_555177 + 8'h01;
  assign sel_555181 = array_index_554988 == array_index_537304 ? add_555180 : sel_555177;
  assign add_555184 = sel_555181 + 8'h01;
  assign sel_555185 = array_index_554988 == array_index_537310 ? add_555184 : sel_555181;
  assign add_555188 = sel_555185 + 8'h01;
  assign sel_555189 = array_index_554988 == array_index_537316 ? add_555188 : sel_555185;
  assign add_555192 = sel_555189 + 8'h01;
  assign sel_555193 = array_index_554988 == array_index_537322 ? add_555192 : sel_555189;
  assign add_555196 = sel_555193 + 8'h01;
  assign sel_555197 = array_index_554988 == array_index_537328 ? add_555196 : sel_555193;
  assign add_555200 = sel_555197 + 8'h01;
  assign sel_555201 = array_index_554988 == array_index_537334 ? add_555200 : sel_555197;
  assign add_555204 = sel_555201 + 8'h01;
  assign sel_555205 = array_index_554988 == array_index_537340 ? add_555204 : sel_555201;
  assign add_555208 = sel_555205 + 8'h01;
  assign sel_555209 = array_index_554988 == array_index_537346 ? add_555208 : sel_555205;
  assign add_555212 = sel_555209 + 8'h01;
  assign sel_555213 = array_index_554988 == array_index_537352 ? add_555212 : sel_555209;
  assign add_555216 = sel_555213 + 8'h01;
  assign sel_555217 = array_index_554988 == array_index_537358 ? add_555216 : sel_555213;
  assign add_555220 = sel_555217 + 8'h01;
  assign sel_555221 = array_index_554988 == array_index_537364 ? add_555220 : sel_555217;
  assign add_555224 = sel_555221 + 8'h01;
  assign sel_555225 = array_index_554988 == array_index_537370 ? add_555224 : sel_555221;
  assign add_555228 = sel_555225 + 8'h01;
  assign sel_555229 = array_index_554988 == array_index_537376 ? add_555228 : sel_555225;
  assign add_555232 = sel_555229 + 8'h01;
  assign sel_555233 = array_index_554988 == array_index_537382 ? add_555232 : sel_555229;
  assign add_555236 = sel_555233 + 8'h01;
  assign sel_555237 = array_index_554988 == array_index_537388 ? add_555236 : sel_555233;
  assign add_555240 = sel_555237 + 8'h01;
  assign sel_555241 = array_index_554988 == array_index_537394 ? add_555240 : sel_555237;
  assign add_555244 = sel_555241 + 8'h01;
  assign sel_555245 = array_index_554988 == array_index_537400 ? add_555244 : sel_555241;
  assign add_555248 = sel_555245 + 8'h01;
  assign sel_555249 = array_index_554988 == array_index_537406 ? add_555248 : sel_555245;
  assign add_555252 = sel_555249 + 8'h01;
  assign sel_555253 = array_index_554988 == array_index_537412 ? add_555252 : sel_555249;
  assign add_555256 = sel_555253 + 8'h01;
  assign sel_555257 = array_index_554988 == array_index_537418 ? add_555256 : sel_555253;
  assign add_555260 = sel_555257 + 8'h01;
  assign sel_555261 = array_index_554988 == array_index_537424 ? add_555260 : sel_555257;
  assign add_555264 = sel_555261 + 8'h01;
  assign sel_555265 = array_index_554988 == array_index_537430 ? add_555264 : sel_555261;
  assign add_555268 = sel_555265 + 8'h01;
  assign sel_555269 = array_index_554988 == array_index_537436 ? add_555268 : sel_555265;
  assign add_555272 = sel_555269 + 8'h01;
  assign sel_555273 = array_index_554988 == array_index_537442 ? add_555272 : sel_555269;
  assign add_555276 = sel_555273 + 8'h01;
  assign sel_555277 = array_index_554988 == array_index_537448 ? add_555276 : sel_555273;
  assign add_555280 = sel_555277 + 8'h01;
  assign sel_555281 = array_index_554988 == array_index_537454 ? add_555280 : sel_555277;
  assign add_555284 = sel_555281 + 8'h01;
  assign sel_555285 = array_index_554988 == array_index_537460 ? add_555284 : sel_555281;
  assign add_555289 = sel_555285 + 8'h01;
  assign array_index_555290 = set1_unflattened[7'h3c];
  assign sel_555291 = array_index_554988 == array_index_537466 ? add_555289 : sel_555285;
  assign add_555294 = sel_555291 + 8'h01;
  assign sel_555295 = array_index_555290 == array_index_537012 ? add_555294 : sel_555291;
  assign add_555298 = sel_555295 + 8'h01;
  assign sel_555299 = array_index_555290 == array_index_537016 ? add_555298 : sel_555295;
  assign add_555302 = sel_555299 + 8'h01;
  assign sel_555303 = array_index_555290 == array_index_537024 ? add_555302 : sel_555299;
  assign add_555306 = sel_555303 + 8'h01;
  assign sel_555307 = array_index_555290 == array_index_537032 ? add_555306 : sel_555303;
  assign add_555310 = sel_555307 + 8'h01;
  assign sel_555311 = array_index_555290 == array_index_537040 ? add_555310 : sel_555307;
  assign add_555314 = sel_555311 + 8'h01;
  assign sel_555315 = array_index_555290 == array_index_537048 ? add_555314 : sel_555311;
  assign add_555318 = sel_555315 + 8'h01;
  assign sel_555319 = array_index_555290 == array_index_537056 ? add_555318 : sel_555315;
  assign add_555322 = sel_555319 + 8'h01;
  assign sel_555323 = array_index_555290 == array_index_537064 ? add_555322 : sel_555319;
  assign add_555326 = sel_555323 + 8'h01;
  assign sel_555327 = array_index_555290 == array_index_537070 ? add_555326 : sel_555323;
  assign add_555330 = sel_555327 + 8'h01;
  assign sel_555331 = array_index_555290 == array_index_537076 ? add_555330 : sel_555327;
  assign add_555334 = sel_555331 + 8'h01;
  assign sel_555335 = array_index_555290 == array_index_537082 ? add_555334 : sel_555331;
  assign add_555338 = sel_555335 + 8'h01;
  assign sel_555339 = array_index_555290 == array_index_537088 ? add_555338 : sel_555335;
  assign add_555342 = sel_555339 + 8'h01;
  assign sel_555343 = array_index_555290 == array_index_537094 ? add_555342 : sel_555339;
  assign add_555346 = sel_555343 + 8'h01;
  assign sel_555347 = array_index_555290 == array_index_537100 ? add_555346 : sel_555343;
  assign add_555350 = sel_555347 + 8'h01;
  assign sel_555351 = array_index_555290 == array_index_537106 ? add_555350 : sel_555347;
  assign add_555354 = sel_555351 + 8'h01;
  assign sel_555355 = array_index_555290 == array_index_537112 ? add_555354 : sel_555351;
  assign add_555358 = sel_555355 + 8'h01;
  assign sel_555359 = array_index_555290 == array_index_537118 ? add_555358 : sel_555355;
  assign add_555362 = sel_555359 + 8'h01;
  assign sel_555363 = array_index_555290 == array_index_537124 ? add_555362 : sel_555359;
  assign add_555366 = sel_555363 + 8'h01;
  assign sel_555367 = array_index_555290 == array_index_537130 ? add_555366 : sel_555363;
  assign add_555370 = sel_555367 + 8'h01;
  assign sel_555371 = array_index_555290 == array_index_537136 ? add_555370 : sel_555367;
  assign add_555374 = sel_555371 + 8'h01;
  assign sel_555375 = array_index_555290 == array_index_537142 ? add_555374 : sel_555371;
  assign add_555378 = sel_555375 + 8'h01;
  assign sel_555379 = array_index_555290 == array_index_537148 ? add_555378 : sel_555375;
  assign add_555382 = sel_555379 + 8'h01;
  assign sel_555383 = array_index_555290 == array_index_537154 ? add_555382 : sel_555379;
  assign add_555386 = sel_555383 + 8'h01;
  assign sel_555387 = array_index_555290 == array_index_537160 ? add_555386 : sel_555383;
  assign add_555390 = sel_555387 + 8'h01;
  assign sel_555391 = array_index_555290 == array_index_537166 ? add_555390 : sel_555387;
  assign add_555394 = sel_555391 + 8'h01;
  assign sel_555395 = array_index_555290 == array_index_537172 ? add_555394 : sel_555391;
  assign add_555398 = sel_555395 + 8'h01;
  assign sel_555399 = array_index_555290 == array_index_537178 ? add_555398 : sel_555395;
  assign add_555402 = sel_555399 + 8'h01;
  assign sel_555403 = array_index_555290 == array_index_537184 ? add_555402 : sel_555399;
  assign add_555406 = sel_555403 + 8'h01;
  assign sel_555407 = array_index_555290 == array_index_537190 ? add_555406 : sel_555403;
  assign add_555410 = sel_555407 + 8'h01;
  assign sel_555411 = array_index_555290 == array_index_537196 ? add_555410 : sel_555407;
  assign add_555414 = sel_555411 + 8'h01;
  assign sel_555415 = array_index_555290 == array_index_537202 ? add_555414 : sel_555411;
  assign add_555418 = sel_555415 + 8'h01;
  assign sel_555419 = array_index_555290 == array_index_537208 ? add_555418 : sel_555415;
  assign add_555422 = sel_555419 + 8'h01;
  assign sel_555423 = array_index_555290 == array_index_537214 ? add_555422 : sel_555419;
  assign add_555426 = sel_555423 + 8'h01;
  assign sel_555427 = array_index_555290 == array_index_537220 ? add_555426 : sel_555423;
  assign add_555430 = sel_555427 + 8'h01;
  assign sel_555431 = array_index_555290 == array_index_537226 ? add_555430 : sel_555427;
  assign add_555434 = sel_555431 + 8'h01;
  assign sel_555435 = array_index_555290 == array_index_537232 ? add_555434 : sel_555431;
  assign add_555438 = sel_555435 + 8'h01;
  assign sel_555439 = array_index_555290 == array_index_537238 ? add_555438 : sel_555435;
  assign add_555442 = sel_555439 + 8'h01;
  assign sel_555443 = array_index_555290 == array_index_537244 ? add_555442 : sel_555439;
  assign add_555446 = sel_555443 + 8'h01;
  assign sel_555447 = array_index_555290 == array_index_537250 ? add_555446 : sel_555443;
  assign add_555450 = sel_555447 + 8'h01;
  assign sel_555451 = array_index_555290 == array_index_537256 ? add_555450 : sel_555447;
  assign add_555454 = sel_555451 + 8'h01;
  assign sel_555455 = array_index_555290 == array_index_537262 ? add_555454 : sel_555451;
  assign add_555458 = sel_555455 + 8'h01;
  assign sel_555459 = array_index_555290 == array_index_537268 ? add_555458 : sel_555455;
  assign add_555462 = sel_555459 + 8'h01;
  assign sel_555463 = array_index_555290 == array_index_537274 ? add_555462 : sel_555459;
  assign add_555466 = sel_555463 + 8'h01;
  assign sel_555467 = array_index_555290 == array_index_537280 ? add_555466 : sel_555463;
  assign add_555470 = sel_555467 + 8'h01;
  assign sel_555471 = array_index_555290 == array_index_537286 ? add_555470 : sel_555467;
  assign add_555474 = sel_555471 + 8'h01;
  assign sel_555475 = array_index_555290 == array_index_537292 ? add_555474 : sel_555471;
  assign add_555478 = sel_555475 + 8'h01;
  assign sel_555479 = array_index_555290 == array_index_537298 ? add_555478 : sel_555475;
  assign add_555482 = sel_555479 + 8'h01;
  assign sel_555483 = array_index_555290 == array_index_537304 ? add_555482 : sel_555479;
  assign add_555486 = sel_555483 + 8'h01;
  assign sel_555487 = array_index_555290 == array_index_537310 ? add_555486 : sel_555483;
  assign add_555490 = sel_555487 + 8'h01;
  assign sel_555491 = array_index_555290 == array_index_537316 ? add_555490 : sel_555487;
  assign add_555494 = sel_555491 + 8'h01;
  assign sel_555495 = array_index_555290 == array_index_537322 ? add_555494 : sel_555491;
  assign add_555498 = sel_555495 + 8'h01;
  assign sel_555499 = array_index_555290 == array_index_537328 ? add_555498 : sel_555495;
  assign add_555502 = sel_555499 + 8'h01;
  assign sel_555503 = array_index_555290 == array_index_537334 ? add_555502 : sel_555499;
  assign add_555506 = sel_555503 + 8'h01;
  assign sel_555507 = array_index_555290 == array_index_537340 ? add_555506 : sel_555503;
  assign add_555510 = sel_555507 + 8'h01;
  assign sel_555511 = array_index_555290 == array_index_537346 ? add_555510 : sel_555507;
  assign add_555514 = sel_555511 + 8'h01;
  assign sel_555515 = array_index_555290 == array_index_537352 ? add_555514 : sel_555511;
  assign add_555518 = sel_555515 + 8'h01;
  assign sel_555519 = array_index_555290 == array_index_537358 ? add_555518 : sel_555515;
  assign add_555522 = sel_555519 + 8'h01;
  assign sel_555523 = array_index_555290 == array_index_537364 ? add_555522 : sel_555519;
  assign add_555526 = sel_555523 + 8'h01;
  assign sel_555527 = array_index_555290 == array_index_537370 ? add_555526 : sel_555523;
  assign add_555530 = sel_555527 + 8'h01;
  assign sel_555531 = array_index_555290 == array_index_537376 ? add_555530 : sel_555527;
  assign add_555534 = sel_555531 + 8'h01;
  assign sel_555535 = array_index_555290 == array_index_537382 ? add_555534 : sel_555531;
  assign add_555538 = sel_555535 + 8'h01;
  assign sel_555539 = array_index_555290 == array_index_537388 ? add_555538 : sel_555535;
  assign add_555542 = sel_555539 + 8'h01;
  assign sel_555543 = array_index_555290 == array_index_537394 ? add_555542 : sel_555539;
  assign add_555546 = sel_555543 + 8'h01;
  assign sel_555547 = array_index_555290 == array_index_537400 ? add_555546 : sel_555543;
  assign add_555550 = sel_555547 + 8'h01;
  assign sel_555551 = array_index_555290 == array_index_537406 ? add_555550 : sel_555547;
  assign add_555554 = sel_555551 + 8'h01;
  assign sel_555555 = array_index_555290 == array_index_537412 ? add_555554 : sel_555551;
  assign add_555558 = sel_555555 + 8'h01;
  assign sel_555559 = array_index_555290 == array_index_537418 ? add_555558 : sel_555555;
  assign add_555562 = sel_555559 + 8'h01;
  assign sel_555563 = array_index_555290 == array_index_537424 ? add_555562 : sel_555559;
  assign add_555566 = sel_555563 + 8'h01;
  assign sel_555567 = array_index_555290 == array_index_537430 ? add_555566 : sel_555563;
  assign add_555570 = sel_555567 + 8'h01;
  assign sel_555571 = array_index_555290 == array_index_537436 ? add_555570 : sel_555567;
  assign add_555574 = sel_555571 + 8'h01;
  assign sel_555575 = array_index_555290 == array_index_537442 ? add_555574 : sel_555571;
  assign add_555578 = sel_555575 + 8'h01;
  assign sel_555579 = array_index_555290 == array_index_537448 ? add_555578 : sel_555575;
  assign add_555582 = sel_555579 + 8'h01;
  assign sel_555583 = array_index_555290 == array_index_537454 ? add_555582 : sel_555579;
  assign add_555586 = sel_555583 + 8'h01;
  assign sel_555587 = array_index_555290 == array_index_537460 ? add_555586 : sel_555583;
  assign add_555591 = sel_555587 + 8'h01;
  assign array_index_555592 = set1_unflattened[7'h3d];
  assign sel_555593 = array_index_555290 == array_index_537466 ? add_555591 : sel_555587;
  assign add_555596 = sel_555593 + 8'h01;
  assign sel_555597 = array_index_555592 == array_index_537012 ? add_555596 : sel_555593;
  assign add_555600 = sel_555597 + 8'h01;
  assign sel_555601 = array_index_555592 == array_index_537016 ? add_555600 : sel_555597;
  assign add_555604 = sel_555601 + 8'h01;
  assign sel_555605 = array_index_555592 == array_index_537024 ? add_555604 : sel_555601;
  assign add_555608 = sel_555605 + 8'h01;
  assign sel_555609 = array_index_555592 == array_index_537032 ? add_555608 : sel_555605;
  assign add_555612 = sel_555609 + 8'h01;
  assign sel_555613 = array_index_555592 == array_index_537040 ? add_555612 : sel_555609;
  assign add_555616 = sel_555613 + 8'h01;
  assign sel_555617 = array_index_555592 == array_index_537048 ? add_555616 : sel_555613;
  assign add_555620 = sel_555617 + 8'h01;
  assign sel_555621 = array_index_555592 == array_index_537056 ? add_555620 : sel_555617;
  assign add_555624 = sel_555621 + 8'h01;
  assign sel_555625 = array_index_555592 == array_index_537064 ? add_555624 : sel_555621;
  assign add_555628 = sel_555625 + 8'h01;
  assign sel_555629 = array_index_555592 == array_index_537070 ? add_555628 : sel_555625;
  assign add_555632 = sel_555629 + 8'h01;
  assign sel_555633 = array_index_555592 == array_index_537076 ? add_555632 : sel_555629;
  assign add_555636 = sel_555633 + 8'h01;
  assign sel_555637 = array_index_555592 == array_index_537082 ? add_555636 : sel_555633;
  assign add_555640 = sel_555637 + 8'h01;
  assign sel_555641 = array_index_555592 == array_index_537088 ? add_555640 : sel_555637;
  assign add_555644 = sel_555641 + 8'h01;
  assign sel_555645 = array_index_555592 == array_index_537094 ? add_555644 : sel_555641;
  assign add_555648 = sel_555645 + 8'h01;
  assign sel_555649 = array_index_555592 == array_index_537100 ? add_555648 : sel_555645;
  assign add_555652 = sel_555649 + 8'h01;
  assign sel_555653 = array_index_555592 == array_index_537106 ? add_555652 : sel_555649;
  assign add_555656 = sel_555653 + 8'h01;
  assign sel_555657 = array_index_555592 == array_index_537112 ? add_555656 : sel_555653;
  assign add_555660 = sel_555657 + 8'h01;
  assign sel_555661 = array_index_555592 == array_index_537118 ? add_555660 : sel_555657;
  assign add_555664 = sel_555661 + 8'h01;
  assign sel_555665 = array_index_555592 == array_index_537124 ? add_555664 : sel_555661;
  assign add_555668 = sel_555665 + 8'h01;
  assign sel_555669 = array_index_555592 == array_index_537130 ? add_555668 : sel_555665;
  assign add_555672 = sel_555669 + 8'h01;
  assign sel_555673 = array_index_555592 == array_index_537136 ? add_555672 : sel_555669;
  assign add_555676 = sel_555673 + 8'h01;
  assign sel_555677 = array_index_555592 == array_index_537142 ? add_555676 : sel_555673;
  assign add_555680 = sel_555677 + 8'h01;
  assign sel_555681 = array_index_555592 == array_index_537148 ? add_555680 : sel_555677;
  assign add_555684 = sel_555681 + 8'h01;
  assign sel_555685 = array_index_555592 == array_index_537154 ? add_555684 : sel_555681;
  assign add_555688 = sel_555685 + 8'h01;
  assign sel_555689 = array_index_555592 == array_index_537160 ? add_555688 : sel_555685;
  assign add_555692 = sel_555689 + 8'h01;
  assign sel_555693 = array_index_555592 == array_index_537166 ? add_555692 : sel_555689;
  assign add_555696 = sel_555693 + 8'h01;
  assign sel_555697 = array_index_555592 == array_index_537172 ? add_555696 : sel_555693;
  assign add_555700 = sel_555697 + 8'h01;
  assign sel_555701 = array_index_555592 == array_index_537178 ? add_555700 : sel_555697;
  assign add_555704 = sel_555701 + 8'h01;
  assign sel_555705 = array_index_555592 == array_index_537184 ? add_555704 : sel_555701;
  assign add_555708 = sel_555705 + 8'h01;
  assign sel_555709 = array_index_555592 == array_index_537190 ? add_555708 : sel_555705;
  assign add_555712 = sel_555709 + 8'h01;
  assign sel_555713 = array_index_555592 == array_index_537196 ? add_555712 : sel_555709;
  assign add_555716 = sel_555713 + 8'h01;
  assign sel_555717 = array_index_555592 == array_index_537202 ? add_555716 : sel_555713;
  assign add_555720 = sel_555717 + 8'h01;
  assign sel_555721 = array_index_555592 == array_index_537208 ? add_555720 : sel_555717;
  assign add_555724 = sel_555721 + 8'h01;
  assign sel_555725 = array_index_555592 == array_index_537214 ? add_555724 : sel_555721;
  assign add_555728 = sel_555725 + 8'h01;
  assign sel_555729 = array_index_555592 == array_index_537220 ? add_555728 : sel_555725;
  assign add_555732 = sel_555729 + 8'h01;
  assign sel_555733 = array_index_555592 == array_index_537226 ? add_555732 : sel_555729;
  assign add_555736 = sel_555733 + 8'h01;
  assign sel_555737 = array_index_555592 == array_index_537232 ? add_555736 : sel_555733;
  assign add_555740 = sel_555737 + 8'h01;
  assign sel_555741 = array_index_555592 == array_index_537238 ? add_555740 : sel_555737;
  assign add_555744 = sel_555741 + 8'h01;
  assign sel_555745 = array_index_555592 == array_index_537244 ? add_555744 : sel_555741;
  assign add_555748 = sel_555745 + 8'h01;
  assign sel_555749 = array_index_555592 == array_index_537250 ? add_555748 : sel_555745;
  assign add_555752 = sel_555749 + 8'h01;
  assign sel_555753 = array_index_555592 == array_index_537256 ? add_555752 : sel_555749;
  assign add_555756 = sel_555753 + 8'h01;
  assign sel_555757 = array_index_555592 == array_index_537262 ? add_555756 : sel_555753;
  assign add_555760 = sel_555757 + 8'h01;
  assign sel_555761 = array_index_555592 == array_index_537268 ? add_555760 : sel_555757;
  assign add_555764 = sel_555761 + 8'h01;
  assign sel_555765 = array_index_555592 == array_index_537274 ? add_555764 : sel_555761;
  assign add_555768 = sel_555765 + 8'h01;
  assign sel_555769 = array_index_555592 == array_index_537280 ? add_555768 : sel_555765;
  assign add_555772 = sel_555769 + 8'h01;
  assign sel_555773 = array_index_555592 == array_index_537286 ? add_555772 : sel_555769;
  assign add_555776 = sel_555773 + 8'h01;
  assign sel_555777 = array_index_555592 == array_index_537292 ? add_555776 : sel_555773;
  assign add_555780 = sel_555777 + 8'h01;
  assign sel_555781 = array_index_555592 == array_index_537298 ? add_555780 : sel_555777;
  assign add_555784 = sel_555781 + 8'h01;
  assign sel_555785 = array_index_555592 == array_index_537304 ? add_555784 : sel_555781;
  assign add_555788 = sel_555785 + 8'h01;
  assign sel_555789 = array_index_555592 == array_index_537310 ? add_555788 : sel_555785;
  assign add_555792 = sel_555789 + 8'h01;
  assign sel_555793 = array_index_555592 == array_index_537316 ? add_555792 : sel_555789;
  assign add_555796 = sel_555793 + 8'h01;
  assign sel_555797 = array_index_555592 == array_index_537322 ? add_555796 : sel_555793;
  assign add_555800 = sel_555797 + 8'h01;
  assign sel_555801 = array_index_555592 == array_index_537328 ? add_555800 : sel_555797;
  assign add_555804 = sel_555801 + 8'h01;
  assign sel_555805 = array_index_555592 == array_index_537334 ? add_555804 : sel_555801;
  assign add_555808 = sel_555805 + 8'h01;
  assign sel_555809 = array_index_555592 == array_index_537340 ? add_555808 : sel_555805;
  assign add_555812 = sel_555809 + 8'h01;
  assign sel_555813 = array_index_555592 == array_index_537346 ? add_555812 : sel_555809;
  assign add_555816 = sel_555813 + 8'h01;
  assign sel_555817 = array_index_555592 == array_index_537352 ? add_555816 : sel_555813;
  assign add_555820 = sel_555817 + 8'h01;
  assign sel_555821 = array_index_555592 == array_index_537358 ? add_555820 : sel_555817;
  assign add_555824 = sel_555821 + 8'h01;
  assign sel_555825 = array_index_555592 == array_index_537364 ? add_555824 : sel_555821;
  assign add_555828 = sel_555825 + 8'h01;
  assign sel_555829 = array_index_555592 == array_index_537370 ? add_555828 : sel_555825;
  assign add_555832 = sel_555829 + 8'h01;
  assign sel_555833 = array_index_555592 == array_index_537376 ? add_555832 : sel_555829;
  assign add_555836 = sel_555833 + 8'h01;
  assign sel_555837 = array_index_555592 == array_index_537382 ? add_555836 : sel_555833;
  assign add_555840 = sel_555837 + 8'h01;
  assign sel_555841 = array_index_555592 == array_index_537388 ? add_555840 : sel_555837;
  assign add_555844 = sel_555841 + 8'h01;
  assign sel_555845 = array_index_555592 == array_index_537394 ? add_555844 : sel_555841;
  assign add_555848 = sel_555845 + 8'h01;
  assign sel_555849 = array_index_555592 == array_index_537400 ? add_555848 : sel_555845;
  assign add_555852 = sel_555849 + 8'h01;
  assign sel_555853 = array_index_555592 == array_index_537406 ? add_555852 : sel_555849;
  assign add_555856 = sel_555853 + 8'h01;
  assign sel_555857 = array_index_555592 == array_index_537412 ? add_555856 : sel_555853;
  assign add_555860 = sel_555857 + 8'h01;
  assign sel_555861 = array_index_555592 == array_index_537418 ? add_555860 : sel_555857;
  assign add_555864 = sel_555861 + 8'h01;
  assign sel_555865 = array_index_555592 == array_index_537424 ? add_555864 : sel_555861;
  assign add_555868 = sel_555865 + 8'h01;
  assign sel_555869 = array_index_555592 == array_index_537430 ? add_555868 : sel_555865;
  assign add_555872 = sel_555869 + 8'h01;
  assign sel_555873 = array_index_555592 == array_index_537436 ? add_555872 : sel_555869;
  assign add_555876 = sel_555873 + 8'h01;
  assign sel_555877 = array_index_555592 == array_index_537442 ? add_555876 : sel_555873;
  assign add_555880 = sel_555877 + 8'h01;
  assign sel_555881 = array_index_555592 == array_index_537448 ? add_555880 : sel_555877;
  assign add_555884 = sel_555881 + 8'h01;
  assign sel_555885 = array_index_555592 == array_index_537454 ? add_555884 : sel_555881;
  assign add_555888 = sel_555885 + 8'h01;
  assign sel_555889 = array_index_555592 == array_index_537460 ? add_555888 : sel_555885;
  assign add_555893 = sel_555889 + 8'h01;
  assign array_index_555894 = set1_unflattened[7'h3e];
  assign sel_555895 = array_index_555592 == array_index_537466 ? add_555893 : sel_555889;
  assign add_555898 = sel_555895 + 8'h01;
  assign sel_555899 = array_index_555894 == array_index_537012 ? add_555898 : sel_555895;
  assign add_555902 = sel_555899 + 8'h01;
  assign sel_555903 = array_index_555894 == array_index_537016 ? add_555902 : sel_555899;
  assign add_555906 = sel_555903 + 8'h01;
  assign sel_555907 = array_index_555894 == array_index_537024 ? add_555906 : sel_555903;
  assign add_555910 = sel_555907 + 8'h01;
  assign sel_555911 = array_index_555894 == array_index_537032 ? add_555910 : sel_555907;
  assign add_555914 = sel_555911 + 8'h01;
  assign sel_555915 = array_index_555894 == array_index_537040 ? add_555914 : sel_555911;
  assign add_555918 = sel_555915 + 8'h01;
  assign sel_555919 = array_index_555894 == array_index_537048 ? add_555918 : sel_555915;
  assign add_555922 = sel_555919 + 8'h01;
  assign sel_555923 = array_index_555894 == array_index_537056 ? add_555922 : sel_555919;
  assign add_555926 = sel_555923 + 8'h01;
  assign sel_555927 = array_index_555894 == array_index_537064 ? add_555926 : sel_555923;
  assign add_555930 = sel_555927 + 8'h01;
  assign sel_555931 = array_index_555894 == array_index_537070 ? add_555930 : sel_555927;
  assign add_555934 = sel_555931 + 8'h01;
  assign sel_555935 = array_index_555894 == array_index_537076 ? add_555934 : sel_555931;
  assign add_555938 = sel_555935 + 8'h01;
  assign sel_555939 = array_index_555894 == array_index_537082 ? add_555938 : sel_555935;
  assign add_555942 = sel_555939 + 8'h01;
  assign sel_555943 = array_index_555894 == array_index_537088 ? add_555942 : sel_555939;
  assign add_555946 = sel_555943 + 8'h01;
  assign sel_555947 = array_index_555894 == array_index_537094 ? add_555946 : sel_555943;
  assign add_555950 = sel_555947 + 8'h01;
  assign sel_555951 = array_index_555894 == array_index_537100 ? add_555950 : sel_555947;
  assign add_555954 = sel_555951 + 8'h01;
  assign sel_555955 = array_index_555894 == array_index_537106 ? add_555954 : sel_555951;
  assign add_555958 = sel_555955 + 8'h01;
  assign sel_555959 = array_index_555894 == array_index_537112 ? add_555958 : sel_555955;
  assign add_555962 = sel_555959 + 8'h01;
  assign sel_555963 = array_index_555894 == array_index_537118 ? add_555962 : sel_555959;
  assign add_555966 = sel_555963 + 8'h01;
  assign sel_555967 = array_index_555894 == array_index_537124 ? add_555966 : sel_555963;
  assign add_555970 = sel_555967 + 8'h01;
  assign sel_555971 = array_index_555894 == array_index_537130 ? add_555970 : sel_555967;
  assign add_555974 = sel_555971 + 8'h01;
  assign sel_555975 = array_index_555894 == array_index_537136 ? add_555974 : sel_555971;
  assign add_555978 = sel_555975 + 8'h01;
  assign sel_555979 = array_index_555894 == array_index_537142 ? add_555978 : sel_555975;
  assign add_555982 = sel_555979 + 8'h01;
  assign sel_555983 = array_index_555894 == array_index_537148 ? add_555982 : sel_555979;
  assign add_555986 = sel_555983 + 8'h01;
  assign sel_555987 = array_index_555894 == array_index_537154 ? add_555986 : sel_555983;
  assign add_555990 = sel_555987 + 8'h01;
  assign sel_555991 = array_index_555894 == array_index_537160 ? add_555990 : sel_555987;
  assign add_555994 = sel_555991 + 8'h01;
  assign sel_555995 = array_index_555894 == array_index_537166 ? add_555994 : sel_555991;
  assign add_555998 = sel_555995 + 8'h01;
  assign sel_555999 = array_index_555894 == array_index_537172 ? add_555998 : sel_555995;
  assign add_556002 = sel_555999 + 8'h01;
  assign sel_556003 = array_index_555894 == array_index_537178 ? add_556002 : sel_555999;
  assign add_556006 = sel_556003 + 8'h01;
  assign sel_556007 = array_index_555894 == array_index_537184 ? add_556006 : sel_556003;
  assign add_556010 = sel_556007 + 8'h01;
  assign sel_556011 = array_index_555894 == array_index_537190 ? add_556010 : sel_556007;
  assign add_556014 = sel_556011 + 8'h01;
  assign sel_556015 = array_index_555894 == array_index_537196 ? add_556014 : sel_556011;
  assign add_556018 = sel_556015 + 8'h01;
  assign sel_556019 = array_index_555894 == array_index_537202 ? add_556018 : sel_556015;
  assign add_556022 = sel_556019 + 8'h01;
  assign sel_556023 = array_index_555894 == array_index_537208 ? add_556022 : sel_556019;
  assign add_556026 = sel_556023 + 8'h01;
  assign sel_556027 = array_index_555894 == array_index_537214 ? add_556026 : sel_556023;
  assign add_556030 = sel_556027 + 8'h01;
  assign sel_556031 = array_index_555894 == array_index_537220 ? add_556030 : sel_556027;
  assign add_556034 = sel_556031 + 8'h01;
  assign sel_556035 = array_index_555894 == array_index_537226 ? add_556034 : sel_556031;
  assign add_556038 = sel_556035 + 8'h01;
  assign sel_556039 = array_index_555894 == array_index_537232 ? add_556038 : sel_556035;
  assign add_556042 = sel_556039 + 8'h01;
  assign sel_556043 = array_index_555894 == array_index_537238 ? add_556042 : sel_556039;
  assign add_556046 = sel_556043 + 8'h01;
  assign sel_556047 = array_index_555894 == array_index_537244 ? add_556046 : sel_556043;
  assign add_556050 = sel_556047 + 8'h01;
  assign sel_556051 = array_index_555894 == array_index_537250 ? add_556050 : sel_556047;
  assign add_556054 = sel_556051 + 8'h01;
  assign sel_556055 = array_index_555894 == array_index_537256 ? add_556054 : sel_556051;
  assign add_556058 = sel_556055 + 8'h01;
  assign sel_556059 = array_index_555894 == array_index_537262 ? add_556058 : sel_556055;
  assign add_556062 = sel_556059 + 8'h01;
  assign sel_556063 = array_index_555894 == array_index_537268 ? add_556062 : sel_556059;
  assign add_556066 = sel_556063 + 8'h01;
  assign sel_556067 = array_index_555894 == array_index_537274 ? add_556066 : sel_556063;
  assign add_556070 = sel_556067 + 8'h01;
  assign sel_556071 = array_index_555894 == array_index_537280 ? add_556070 : sel_556067;
  assign add_556074 = sel_556071 + 8'h01;
  assign sel_556075 = array_index_555894 == array_index_537286 ? add_556074 : sel_556071;
  assign add_556078 = sel_556075 + 8'h01;
  assign sel_556079 = array_index_555894 == array_index_537292 ? add_556078 : sel_556075;
  assign add_556082 = sel_556079 + 8'h01;
  assign sel_556083 = array_index_555894 == array_index_537298 ? add_556082 : sel_556079;
  assign add_556086 = sel_556083 + 8'h01;
  assign sel_556087 = array_index_555894 == array_index_537304 ? add_556086 : sel_556083;
  assign add_556090 = sel_556087 + 8'h01;
  assign sel_556091 = array_index_555894 == array_index_537310 ? add_556090 : sel_556087;
  assign add_556094 = sel_556091 + 8'h01;
  assign sel_556095 = array_index_555894 == array_index_537316 ? add_556094 : sel_556091;
  assign add_556098 = sel_556095 + 8'h01;
  assign sel_556099 = array_index_555894 == array_index_537322 ? add_556098 : sel_556095;
  assign add_556102 = sel_556099 + 8'h01;
  assign sel_556103 = array_index_555894 == array_index_537328 ? add_556102 : sel_556099;
  assign add_556106 = sel_556103 + 8'h01;
  assign sel_556107 = array_index_555894 == array_index_537334 ? add_556106 : sel_556103;
  assign add_556110 = sel_556107 + 8'h01;
  assign sel_556111 = array_index_555894 == array_index_537340 ? add_556110 : sel_556107;
  assign add_556114 = sel_556111 + 8'h01;
  assign sel_556115 = array_index_555894 == array_index_537346 ? add_556114 : sel_556111;
  assign add_556118 = sel_556115 + 8'h01;
  assign sel_556119 = array_index_555894 == array_index_537352 ? add_556118 : sel_556115;
  assign add_556122 = sel_556119 + 8'h01;
  assign sel_556123 = array_index_555894 == array_index_537358 ? add_556122 : sel_556119;
  assign add_556126 = sel_556123 + 8'h01;
  assign sel_556127 = array_index_555894 == array_index_537364 ? add_556126 : sel_556123;
  assign add_556130 = sel_556127 + 8'h01;
  assign sel_556131 = array_index_555894 == array_index_537370 ? add_556130 : sel_556127;
  assign add_556134 = sel_556131 + 8'h01;
  assign sel_556135 = array_index_555894 == array_index_537376 ? add_556134 : sel_556131;
  assign add_556138 = sel_556135 + 8'h01;
  assign sel_556139 = array_index_555894 == array_index_537382 ? add_556138 : sel_556135;
  assign add_556142 = sel_556139 + 8'h01;
  assign sel_556143 = array_index_555894 == array_index_537388 ? add_556142 : sel_556139;
  assign add_556146 = sel_556143 + 8'h01;
  assign sel_556147 = array_index_555894 == array_index_537394 ? add_556146 : sel_556143;
  assign add_556150 = sel_556147 + 8'h01;
  assign sel_556151 = array_index_555894 == array_index_537400 ? add_556150 : sel_556147;
  assign add_556154 = sel_556151 + 8'h01;
  assign sel_556155 = array_index_555894 == array_index_537406 ? add_556154 : sel_556151;
  assign add_556158 = sel_556155 + 8'h01;
  assign sel_556159 = array_index_555894 == array_index_537412 ? add_556158 : sel_556155;
  assign add_556162 = sel_556159 + 8'h01;
  assign sel_556163 = array_index_555894 == array_index_537418 ? add_556162 : sel_556159;
  assign add_556166 = sel_556163 + 8'h01;
  assign sel_556167 = array_index_555894 == array_index_537424 ? add_556166 : sel_556163;
  assign add_556170 = sel_556167 + 8'h01;
  assign sel_556171 = array_index_555894 == array_index_537430 ? add_556170 : sel_556167;
  assign add_556174 = sel_556171 + 8'h01;
  assign sel_556175 = array_index_555894 == array_index_537436 ? add_556174 : sel_556171;
  assign add_556178 = sel_556175 + 8'h01;
  assign sel_556179 = array_index_555894 == array_index_537442 ? add_556178 : sel_556175;
  assign add_556182 = sel_556179 + 8'h01;
  assign sel_556183 = array_index_555894 == array_index_537448 ? add_556182 : sel_556179;
  assign add_556186 = sel_556183 + 8'h01;
  assign sel_556187 = array_index_555894 == array_index_537454 ? add_556186 : sel_556183;
  assign add_556190 = sel_556187 + 8'h01;
  assign sel_556191 = array_index_555894 == array_index_537460 ? add_556190 : sel_556187;
  assign add_556195 = sel_556191 + 8'h01;
  assign array_index_556196 = set1_unflattened[7'h3f];
  assign sel_556197 = array_index_555894 == array_index_537466 ? add_556195 : sel_556191;
  assign add_556200 = sel_556197 + 8'h01;
  assign sel_556201 = array_index_556196 == array_index_537012 ? add_556200 : sel_556197;
  assign add_556204 = sel_556201 + 8'h01;
  assign sel_556205 = array_index_556196 == array_index_537016 ? add_556204 : sel_556201;
  assign add_556208 = sel_556205 + 8'h01;
  assign sel_556209 = array_index_556196 == array_index_537024 ? add_556208 : sel_556205;
  assign add_556212 = sel_556209 + 8'h01;
  assign sel_556213 = array_index_556196 == array_index_537032 ? add_556212 : sel_556209;
  assign add_556216 = sel_556213 + 8'h01;
  assign sel_556217 = array_index_556196 == array_index_537040 ? add_556216 : sel_556213;
  assign add_556220 = sel_556217 + 8'h01;
  assign sel_556221 = array_index_556196 == array_index_537048 ? add_556220 : sel_556217;
  assign add_556224 = sel_556221 + 8'h01;
  assign sel_556225 = array_index_556196 == array_index_537056 ? add_556224 : sel_556221;
  assign add_556228 = sel_556225 + 8'h01;
  assign sel_556229 = array_index_556196 == array_index_537064 ? add_556228 : sel_556225;
  assign add_556232 = sel_556229 + 8'h01;
  assign sel_556233 = array_index_556196 == array_index_537070 ? add_556232 : sel_556229;
  assign add_556236 = sel_556233 + 8'h01;
  assign sel_556237 = array_index_556196 == array_index_537076 ? add_556236 : sel_556233;
  assign add_556240 = sel_556237 + 8'h01;
  assign sel_556241 = array_index_556196 == array_index_537082 ? add_556240 : sel_556237;
  assign add_556244 = sel_556241 + 8'h01;
  assign sel_556245 = array_index_556196 == array_index_537088 ? add_556244 : sel_556241;
  assign add_556248 = sel_556245 + 8'h01;
  assign sel_556249 = array_index_556196 == array_index_537094 ? add_556248 : sel_556245;
  assign add_556252 = sel_556249 + 8'h01;
  assign sel_556253 = array_index_556196 == array_index_537100 ? add_556252 : sel_556249;
  assign add_556256 = sel_556253 + 8'h01;
  assign sel_556257 = array_index_556196 == array_index_537106 ? add_556256 : sel_556253;
  assign add_556260 = sel_556257 + 8'h01;
  assign sel_556261 = array_index_556196 == array_index_537112 ? add_556260 : sel_556257;
  assign add_556264 = sel_556261 + 8'h01;
  assign sel_556265 = array_index_556196 == array_index_537118 ? add_556264 : sel_556261;
  assign add_556268 = sel_556265 + 8'h01;
  assign sel_556269 = array_index_556196 == array_index_537124 ? add_556268 : sel_556265;
  assign add_556272 = sel_556269 + 8'h01;
  assign sel_556273 = array_index_556196 == array_index_537130 ? add_556272 : sel_556269;
  assign add_556276 = sel_556273 + 8'h01;
  assign sel_556277 = array_index_556196 == array_index_537136 ? add_556276 : sel_556273;
  assign add_556280 = sel_556277 + 8'h01;
  assign sel_556281 = array_index_556196 == array_index_537142 ? add_556280 : sel_556277;
  assign add_556284 = sel_556281 + 8'h01;
  assign sel_556285 = array_index_556196 == array_index_537148 ? add_556284 : sel_556281;
  assign add_556288 = sel_556285 + 8'h01;
  assign sel_556289 = array_index_556196 == array_index_537154 ? add_556288 : sel_556285;
  assign add_556292 = sel_556289 + 8'h01;
  assign sel_556293 = array_index_556196 == array_index_537160 ? add_556292 : sel_556289;
  assign add_556296 = sel_556293 + 8'h01;
  assign sel_556297 = array_index_556196 == array_index_537166 ? add_556296 : sel_556293;
  assign add_556300 = sel_556297 + 8'h01;
  assign sel_556301 = array_index_556196 == array_index_537172 ? add_556300 : sel_556297;
  assign add_556304 = sel_556301 + 8'h01;
  assign sel_556305 = array_index_556196 == array_index_537178 ? add_556304 : sel_556301;
  assign add_556308 = sel_556305 + 8'h01;
  assign sel_556309 = array_index_556196 == array_index_537184 ? add_556308 : sel_556305;
  assign add_556312 = sel_556309 + 8'h01;
  assign sel_556313 = array_index_556196 == array_index_537190 ? add_556312 : sel_556309;
  assign add_556316 = sel_556313 + 8'h01;
  assign sel_556317 = array_index_556196 == array_index_537196 ? add_556316 : sel_556313;
  assign add_556320 = sel_556317 + 8'h01;
  assign sel_556321 = array_index_556196 == array_index_537202 ? add_556320 : sel_556317;
  assign add_556324 = sel_556321 + 8'h01;
  assign sel_556325 = array_index_556196 == array_index_537208 ? add_556324 : sel_556321;
  assign add_556328 = sel_556325 + 8'h01;
  assign sel_556329 = array_index_556196 == array_index_537214 ? add_556328 : sel_556325;
  assign add_556332 = sel_556329 + 8'h01;
  assign sel_556333 = array_index_556196 == array_index_537220 ? add_556332 : sel_556329;
  assign add_556336 = sel_556333 + 8'h01;
  assign sel_556337 = array_index_556196 == array_index_537226 ? add_556336 : sel_556333;
  assign add_556340 = sel_556337 + 8'h01;
  assign sel_556341 = array_index_556196 == array_index_537232 ? add_556340 : sel_556337;
  assign add_556344 = sel_556341 + 8'h01;
  assign sel_556345 = array_index_556196 == array_index_537238 ? add_556344 : sel_556341;
  assign add_556348 = sel_556345 + 8'h01;
  assign sel_556349 = array_index_556196 == array_index_537244 ? add_556348 : sel_556345;
  assign add_556352 = sel_556349 + 8'h01;
  assign sel_556353 = array_index_556196 == array_index_537250 ? add_556352 : sel_556349;
  assign add_556356 = sel_556353 + 8'h01;
  assign sel_556357 = array_index_556196 == array_index_537256 ? add_556356 : sel_556353;
  assign add_556360 = sel_556357 + 8'h01;
  assign sel_556361 = array_index_556196 == array_index_537262 ? add_556360 : sel_556357;
  assign add_556364 = sel_556361 + 8'h01;
  assign sel_556365 = array_index_556196 == array_index_537268 ? add_556364 : sel_556361;
  assign add_556368 = sel_556365 + 8'h01;
  assign sel_556369 = array_index_556196 == array_index_537274 ? add_556368 : sel_556365;
  assign add_556372 = sel_556369 + 8'h01;
  assign sel_556373 = array_index_556196 == array_index_537280 ? add_556372 : sel_556369;
  assign add_556376 = sel_556373 + 8'h01;
  assign sel_556377 = array_index_556196 == array_index_537286 ? add_556376 : sel_556373;
  assign add_556380 = sel_556377 + 8'h01;
  assign sel_556381 = array_index_556196 == array_index_537292 ? add_556380 : sel_556377;
  assign add_556384 = sel_556381 + 8'h01;
  assign sel_556385 = array_index_556196 == array_index_537298 ? add_556384 : sel_556381;
  assign add_556388 = sel_556385 + 8'h01;
  assign sel_556389 = array_index_556196 == array_index_537304 ? add_556388 : sel_556385;
  assign add_556392 = sel_556389 + 8'h01;
  assign sel_556393 = array_index_556196 == array_index_537310 ? add_556392 : sel_556389;
  assign add_556396 = sel_556393 + 8'h01;
  assign sel_556397 = array_index_556196 == array_index_537316 ? add_556396 : sel_556393;
  assign add_556400 = sel_556397 + 8'h01;
  assign sel_556401 = array_index_556196 == array_index_537322 ? add_556400 : sel_556397;
  assign add_556404 = sel_556401 + 8'h01;
  assign sel_556405 = array_index_556196 == array_index_537328 ? add_556404 : sel_556401;
  assign add_556408 = sel_556405 + 8'h01;
  assign sel_556409 = array_index_556196 == array_index_537334 ? add_556408 : sel_556405;
  assign add_556412 = sel_556409 + 8'h01;
  assign sel_556413 = array_index_556196 == array_index_537340 ? add_556412 : sel_556409;
  assign add_556416 = sel_556413 + 8'h01;
  assign sel_556417 = array_index_556196 == array_index_537346 ? add_556416 : sel_556413;
  assign add_556420 = sel_556417 + 8'h01;
  assign sel_556421 = array_index_556196 == array_index_537352 ? add_556420 : sel_556417;
  assign add_556424 = sel_556421 + 8'h01;
  assign sel_556425 = array_index_556196 == array_index_537358 ? add_556424 : sel_556421;
  assign add_556428 = sel_556425 + 8'h01;
  assign sel_556429 = array_index_556196 == array_index_537364 ? add_556428 : sel_556425;
  assign add_556432 = sel_556429 + 8'h01;
  assign sel_556433 = array_index_556196 == array_index_537370 ? add_556432 : sel_556429;
  assign add_556436 = sel_556433 + 8'h01;
  assign sel_556437 = array_index_556196 == array_index_537376 ? add_556436 : sel_556433;
  assign add_556440 = sel_556437 + 8'h01;
  assign sel_556441 = array_index_556196 == array_index_537382 ? add_556440 : sel_556437;
  assign add_556444 = sel_556441 + 8'h01;
  assign sel_556445 = array_index_556196 == array_index_537388 ? add_556444 : sel_556441;
  assign add_556448 = sel_556445 + 8'h01;
  assign sel_556449 = array_index_556196 == array_index_537394 ? add_556448 : sel_556445;
  assign add_556452 = sel_556449 + 8'h01;
  assign sel_556453 = array_index_556196 == array_index_537400 ? add_556452 : sel_556449;
  assign add_556456 = sel_556453 + 8'h01;
  assign sel_556457 = array_index_556196 == array_index_537406 ? add_556456 : sel_556453;
  assign add_556460 = sel_556457 + 8'h01;
  assign sel_556461 = array_index_556196 == array_index_537412 ? add_556460 : sel_556457;
  assign add_556464 = sel_556461 + 8'h01;
  assign sel_556465 = array_index_556196 == array_index_537418 ? add_556464 : sel_556461;
  assign add_556468 = sel_556465 + 8'h01;
  assign sel_556469 = array_index_556196 == array_index_537424 ? add_556468 : sel_556465;
  assign add_556472 = sel_556469 + 8'h01;
  assign sel_556473 = array_index_556196 == array_index_537430 ? add_556472 : sel_556469;
  assign add_556476 = sel_556473 + 8'h01;
  assign sel_556477 = array_index_556196 == array_index_537436 ? add_556476 : sel_556473;
  assign add_556480 = sel_556477 + 8'h01;
  assign sel_556481 = array_index_556196 == array_index_537442 ? add_556480 : sel_556477;
  assign add_556484 = sel_556481 + 8'h01;
  assign sel_556485 = array_index_556196 == array_index_537448 ? add_556484 : sel_556481;
  assign add_556488 = sel_556485 + 8'h01;
  assign sel_556489 = array_index_556196 == array_index_537454 ? add_556488 : sel_556485;
  assign add_556492 = sel_556489 + 8'h01;
  assign sel_556493 = array_index_556196 == array_index_537460 ? add_556492 : sel_556489;
  assign add_556497 = sel_556493 + 8'h01;
  assign array_index_556498 = set1_unflattened[7'h40];
  assign sel_556499 = array_index_556196 == array_index_537466 ? add_556497 : sel_556493;
  assign add_556502 = sel_556499 + 8'h01;
  assign sel_556503 = array_index_556498 == array_index_537012 ? add_556502 : sel_556499;
  assign add_556506 = sel_556503 + 8'h01;
  assign sel_556507 = array_index_556498 == array_index_537016 ? add_556506 : sel_556503;
  assign add_556510 = sel_556507 + 8'h01;
  assign sel_556511 = array_index_556498 == array_index_537024 ? add_556510 : sel_556507;
  assign add_556514 = sel_556511 + 8'h01;
  assign sel_556515 = array_index_556498 == array_index_537032 ? add_556514 : sel_556511;
  assign add_556518 = sel_556515 + 8'h01;
  assign sel_556519 = array_index_556498 == array_index_537040 ? add_556518 : sel_556515;
  assign add_556522 = sel_556519 + 8'h01;
  assign sel_556523 = array_index_556498 == array_index_537048 ? add_556522 : sel_556519;
  assign add_556526 = sel_556523 + 8'h01;
  assign sel_556527 = array_index_556498 == array_index_537056 ? add_556526 : sel_556523;
  assign add_556530 = sel_556527 + 8'h01;
  assign sel_556531 = array_index_556498 == array_index_537064 ? add_556530 : sel_556527;
  assign add_556534 = sel_556531 + 8'h01;
  assign sel_556535 = array_index_556498 == array_index_537070 ? add_556534 : sel_556531;
  assign add_556538 = sel_556535 + 8'h01;
  assign sel_556539 = array_index_556498 == array_index_537076 ? add_556538 : sel_556535;
  assign add_556542 = sel_556539 + 8'h01;
  assign sel_556543 = array_index_556498 == array_index_537082 ? add_556542 : sel_556539;
  assign add_556546 = sel_556543 + 8'h01;
  assign sel_556547 = array_index_556498 == array_index_537088 ? add_556546 : sel_556543;
  assign add_556550 = sel_556547 + 8'h01;
  assign sel_556551 = array_index_556498 == array_index_537094 ? add_556550 : sel_556547;
  assign add_556554 = sel_556551 + 8'h01;
  assign sel_556555 = array_index_556498 == array_index_537100 ? add_556554 : sel_556551;
  assign add_556558 = sel_556555 + 8'h01;
  assign sel_556559 = array_index_556498 == array_index_537106 ? add_556558 : sel_556555;
  assign add_556562 = sel_556559 + 8'h01;
  assign sel_556563 = array_index_556498 == array_index_537112 ? add_556562 : sel_556559;
  assign add_556566 = sel_556563 + 8'h01;
  assign sel_556567 = array_index_556498 == array_index_537118 ? add_556566 : sel_556563;
  assign add_556570 = sel_556567 + 8'h01;
  assign sel_556571 = array_index_556498 == array_index_537124 ? add_556570 : sel_556567;
  assign add_556574 = sel_556571 + 8'h01;
  assign sel_556575 = array_index_556498 == array_index_537130 ? add_556574 : sel_556571;
  assign add_556578 = sel_556575 + 8'h01;
  assign sel_556579 = array_index_556498 == array_index_537136 ? add_556578 : sel_556575;
  assign add_556582 = sel_556579 + 8'h01;
  assign sel_556583 = array_index_556498 == array_index_537142 ? add_556582 : sel_556579;
  assign add_556586 = sel_556583 + 8'h01;
  assign sel_556587 = array_index_556498 == array_index_537148 ? add_556586 : sel_556583;
  assign add_556590 = sel_556587 + 8'h01;
  assign sel_556591 = array_index_556498 == array_index_537154 ? add_556590 : sel_556587;
  assign add_556594 = sel_556591 + 8'h01;
  assign sel_556595 = array_index_556498 == array_index_537160 ? add_556594 : sel_556591;
  assign add_556598 = sel_556595 + 8'h01;
  assign sel_556599 = array_index_556498 == array_index_537166 ? add_556598 : sel_556595;
  assign add_556602 = sel_556599 + 8'h01;
  assign sel_556603 = array_index_556498 == array_index_537172 ? add_556602 : sel_556599;
  assign add_556606 = sel_556603 + 8'h01;
  assign sel_556607 = array_index_556498 == array_index_537178 ? add_556606 : sel_556603;
  assign add_556610 = sel_556607 + 8'h01;
  assign sel_556611 = array_index_556498 == array_index_537184 ? add_556610 : sel_556607;
  assign add_556614 = sel_556611 + 8'h01;
  assign sel_556615 = array_index_556498 == array_index_537190 ? add_556614 : sel_556611;
  assign add_556618 = sel_556615 + 8'h01;
  assign sel_556619 = array_index_556498 == array_index_537196 ? add_556618 : sel_556615;
  assign add_556622 = sel_556619 + 8'h01;
  assign sel_556623 = array_index_556498 == array_index_537202 ? add_556622 : sel_556619;
  assign add_556626 = sel_556623 + 8'h01;
  assign sel_556627 = array_index_556498 == array_index_537208 ? add_556626 : sel_556623;
  assign add_556630 = sel_556627 + 8'h01;
  assign sel_556631 = array_index_556498 == array_index_537214 ? add_556630 : sel_556627;
  assign add_556634 = sel_556631 + 8'h01;
  assign sel_556635 = array_index_556498 == array_index_537220 ? add_556634 : sel_556631;
  assign add_556638 = sel_556635 + 8'h01;
  assign sel_556639 = array_index_556498 == array_index_537226 ? add_556638 : sel_556635;
  assign add_556642 = sel_556639 + 8'h01;
  assign sel_556643 = array_index_556498 == array_index_537232 ? add_556642 : sel_556639;
  assign add_556646 = sel_556643 + 8'h01;
  assign sel_556647 = array_index_556498 == array_index_537238 ? add_556646 : sel_556643;
  assign add_556650 = sel_556647 + 8'h01;
  assign sel_556651 = array_index_556498 == array_index_537244 ? add_556650 : sel_556647;
  assign add_556654 = sel_556651 + 8'h01;
  assign sel_556655 = array_index_556498 == array_index_537250 ? add_556654 : sel_556651;
  assign add_556658 = sel_556655 + 8'h01;
  assign sel_556659 = array_index_556498 == array_index_537256 ? add_556658 : sel_556655;
  assign add_556662 = sel_556659 + 8'h01;
  assign sel_556663 = array_index_556498 == array_index_537262 ? add_556662 : sel_556659;
  assign add_556666 = sel_556663 + 8'h01;
  assign sel_556667 = array_index_556498 == array_index_537268 ? add_556666 : sel_556663;
  assign add_556670 = sel_556667 + 8'h01;
  assign sel_556671 = array_index_556498 == array_index_537274 ? add_556670 : sel_556667;
  assign add_556674 = sel_556671 + 8'h01;
  assign sel_556675 = array_index_556498 == array_index_537280 ? add_556674 : sel_556671;
  assign add_556678 = sel_556675 + 8'h01;
  assign sel_556679 = array_index_556498 == array_index_537286 ? add_556678 : sel_556675;
  assign add_556682 = sel_556679 + 8'h01;
  assign sel_556683 = array_index_556498 == array_index_537292 ? add_556682 : sel_556679;
  assign add_556686 = sel_556683 + 8'h01;
  assign sel_556687 = array_index_556498 == array_index_537298 ? add_556686 : sel_556683;
  assign add_556690 = sel_556687 + 8'h01;
  assign sel_556691 = array_index_556498 == array_index_537304 ? add_556690 : sel_556687;
  assign add_556694 = sel_556691 + 8'h01;
  assign sel_556695 = array_index_556498 == array_index_537310 ? add_556694 : sel_556691;
  assign add_556698 = sel_556695 + 8'h01;
  assign sel_556699 = array_index_556498 == array_index_537316 ? add_556698 : sel_556695;
  assign add_556702 = sel_556699 + 8'h01;
  assign sel_556703 = array_index_556498 == array_index_537322 ? add_556702 : sel_556699;
  assign add_556706 = sel_556703 + 8'h01;
  assign sel_556707 = array_index_556498 == array_index_537328 ? add_556706 : sel_556703;
  assign add_556710 = sel_556707 + 8'h01;
  assign sel_556711 = array_index_556498 == array_index_537334 ? add_556710 : sel_556707;
  assign add_556714 = sel_556711 + 8'h01;
  assign sel_556715 = array_index_556498 == array_index_537340 ? add_556714 : sel_556711;
  assign add_556718 = sel_556715 + 8'h01;
  assign sel_556719 = array_index_556498 == array_index_537346 ? add_556718 : sel_556715;
  assign add_556722 = sel_556719 + 8'h01;
  assign sel_556723 = array_index_556498 == array_index_537352 ? add_556722 : sel_556719;
  assign add_556726 = sel_556723 + 8'h01;
  assign sel_556727 = array_index_556498 == array_index_537358 ? add_556726 : sel_556723;
  assign add_556730 = sel_556727 + 8'h01;
  assign sel_556731 = array_index_556498 == array_index_537364 ? add_556730 : sel_556727;
  assign add_556734 = sel_556731 + 8'h01;
  assign sel_556735 = array_index_556498 == array_index_537370 ? add_556734 : sel_556731;
  assign add_556738 = sel_556735 + 8'h01;
  assign sel_556739 = array_index_556498 == array_index_537376 ? add_556738 : sel_556735;
  assign add_556742 = sel_556739 + 8'h01;
  assign sel_556743 = array_index_556498 == array_index_537382 ? add_556742 : sel_556739;
  assign add_556746 = sel_556743 + 8'h01;
  assign sel_556747 = array_index_556498 == array_index_537388 ? add_556746 : sel_556743;
  assign add_556750 = sel_556747 + 8'h01;
  assign sel_556751 = array_index_556498 == array_index_537394 ? add_556750 : sel_556747;
  assign add_556754 = sel_556751 + 8'h01;
  assign sel_556755 = array_index_556498 == array_index_537400 ? add_556754 : sel_556751;
  assign add_556758 = sel_556755 + 8'h01;
  assign sel_556759 = array_index_556498 == array_index_537406 ? add_556758 : sel_556755;
  assign add_556762 = sel_556759 + 8'h01;
  assign sel_556763 = array_index_556498 == array_index_537412 ? add_556762 : sel_556759;
  assign add_556766 = sel_556763 + 8'h01;
  assign sel_556767 = array_index_556498 == array_index_537418 ? add_556766 : sel_556763;
  assign add_556770 = sel_556767 + 8'h01;
  assign sel_556771 = array_index_556498 == array_index_537424 ? add_556770 : sel_556767;
  assign add_556774 = sel_556771 + 8'h01;
  assign sel_556775 = array_index_556498 == array_index_537430 ? add_556774 : sel_556771;
  assign add_556778 = sel_556775 + 8'h01;
  assign sel_556779 = array_index_556498 == array_index_537436 ? add_556778 : sel_556775;
  assign add_556782 = sel_556779 + 8'h01;
  assign sel_556783 = array_index_556498 == array_index_537442 ? add_556782 : sel_556779;
  assign add_556786 = sel_556783 + 8'h01;
  assign sel_556787 = array_index_556498 == array_index_537448 ? add_556786 : sel_556783;
  assign add_556790 = sel_556787 + 8'h01;
  assign sel_556791 = array_index_556498 == array_index_537454 ? add_556790 : sel_556787;
  assign add_556794 = sel_556791 + 8'h01;
  assign sel_556795 = array_index_556498 == array_index_537460 ? add_556794 : sel_556791;
  assign add_556799 = sel_556795 + 8'h01;
  assign array_index_556800 = set1_unflattened[7'h41];
  assign sel_556801 = array_index_556498 == array_index_537466 ? add_556799 : sel_556795;
  assign add_556804 = sel_556801 + 8'h01;
  assign sel_556805 = array_index_556800 == array_index_537012 ? add_556804 : sel_556801;
  assign add_556808 = sel_556805 + 8'h01;
  assign sel_556809 = array_index_556800 == array_index_537016 ? add_556808 : sel_556805;
  assign add_556812 = sel_556809 + 8'h01;
  assign sel_556813 = array_index_556800 == array_index_537024 ? add_556812 : sel_556809;
  assign add_556816 = sel_556813 + 8'h01;
  assign sel_556817 = array_index_556800 == array_index_537032 ? add_556816 : sel_556813;
  assign add_556820 = sel_556817 + 8'h01;
  assign sel_556821 = array_index_556800 == array_index_537040 ? add_556820 : sel_556817;
  assign add_556824 = sel_556821 + 8'h01;
  assign sel_556825 = array_index_556800 == array_index_537048 ? add_556824 : sel_556821;
  assign add_556828 = sel_556825 + 8'h01;
  assign sel_556829 = array_index_556800 == array_index_537056 ? add_556828 : sel_556825;
  assign add_556832 = sel_556829 + 8'h01;
  assign sel_556833 = array_index_556800 == array_index_537064 ? add_556832 : sel_556829;
  assign add_556836 = sel_556833 + 8'h01;
  assign sel_556837 = array_index_556800 == array_index_537070 ? add_556836 : sel_556833;
  assign add_556840 = sel_556837 + 8'h01;
  assign sel_556841 = array_index_556800 == array_index_537076 ? add_556840 : sel_556837;
  assign add_556844 = sel_556841 + 8'h01;
  assign sel_556845 = array_index_556800 == array_index_537082 ? add_556844 : sel_556841;
  assign add_556848 = sel_556845 + 8'h01;
  assign sel_556849 = array_index_556800 == array_index_537088 ? add_556848 : sel_556845;
  assign add_556852 = sel_556849 + 8'h01;
  assign sel_556853 = array_index_556800 == array_index_537094 ? add_556852 : sel_556849;
  assign add_556856 = sel_556853 + 8'h01;
  assign sel_556857 = array_index_556800 == array_index_537100 ? add_556856 : sel_556853;
  assign add_556860 = sel_556857 + 8'h01;
  assign sel_556861 = array_index_556800 == array_index_537106 ? add_556860 : sel_556857;
  assign add_556864 = sel_556861 + 8'h01;
  assign sel_556865 = array_index_556800 == array_index_537112 ? add_556864 : sel_556861;
  assign add_556868 = sel_556865 + 8'h01;
  assign sel_556869 = array_index_556800 == array_index_537118 ? add_556868 : sel_556865;
  assign add_556872 = sel_556869 + 8'h01;
  assign sel_556873 = array_index_556800 == array_index_537124 ? add_556872 : sel_556869;
  assign add_556876 = sel_556873 + 8'h01;
  assign sel_556877 = array_index_556800 == array_index_537130 ? add_556876 : sel_556873;
  assign add_556880 = sel_556877 + 8'h01;
  assign sel_556881 = array_index_556800 == array_index_537136 ? add_556880 : sel_556877;
  assign add_556884 = sel_556881 + 8'h01;
  assign sel_556885 = array_index_556800 == array_index_537142 ? add_556884 : sel_556881;
  assign add_556888 = sel_556885 + 8'h01;
  assign sel_556889 = array_index_556800 == array_index_537148 ? add_556888 : sel_556885;
  assign add_556892 = sel_556889 + 8'h01;
  assign sel_556893 = array_index_556800 == array_index_537154 ? add_556892 : sel_556889;
  assign add_556896 = sel_556893 + 8'h01;
  assign sel_556897 = array_index_556800 == array_index_537160 ? add_556896 : sel_556893;
  assign add_556900 = sel_556897 + 8'h01;
  assign sel_556901 = array_index_556800 == array_index_537166 ? add_556900 : sel_556897;
  assign add_556904 = sel_556901 + 8'h01;
  assign sel_556905 = array_index_556800 == array_index_537172 ? add_556904 : sel_556901;
  assign add_556908 = sel_556905 + 8'h01;
  assign sel_556909 = array_index_556800 == array_index_537178 ? add_556908 : sel_556905;
  assign add_556912 = sel_556909 + 8'h01;
  assign sel_556913 = array_index_556800 == array_index_537184 ? add_556912 : sel_556909;
  assign add_556916 = sel_556913 + 8'h01;
  assign sel_556917 = array_index_556800 == array_index_537190 ? add_556916 : sel_556913;
  assign add_556920 = sel_556917 + 8'h01;
  assign sel_556921 = array_index_556800 == array_index_537196 ? add_556920 : sel_556917;
  assign add_556924 = sel_556921 + 8'h01;
  assign sel_556925 = array_index_556800 == array_index_537202 ? add_556924 : sel_556921;
  assign add_556928 = sel_556925 + 8'h01;
  assign sel_556929 = array_index_556800 == array_index_537208 ? add_556928 : sel_556925;
  assign add_556932 = sel_556929 + 8'h01;
  assign sel_556933 = array_index_556800 == array_index_537214 ? add_556932 : sel_556929;
  assign add_556936 = sel_556933 + 8'h01;
  assign sel_556937 = array_index_556800 == array_index_537220 ? add_556936 : sel_556933;
  assign add_556940 = sel_556937 + 8'h01;
  assign sel_556941 = array_index_556800 == array_index_537226 ? add_556940 : sel_556937;
  assign add_556944 = sel_556941 + 8'h01;
  assign sel_556945 = array_index_556800 == array_index_537232 ? add_556944 : sel_556941;
  assign add_556948 = sel_556945 + 8'h01;
  assign sel_556949 = array_index_556800 == array_index_537238 ? add_556948 : sel_556945;
  assign add_556952 = sel_556949 + 8'h01;
  assign sel_556953 = array_index_556800 == array_index_537244 ? add_556952 : sel_556949;
  assign add_556956 = sel_556953 + 8'h01;
  assign sel_556957 = array_index_556800 == array_index_537250 ? add_556956 : sel_556953;
  assign add_556960 = sel_556957 + 8'h01;
  assign sel_556961 = array_index_556800 == array_index_537256 ? add_556960 : sel_556957;
  assign add_556964 = sel_556961 + 8'h01;
  assign sel_556965 = array_index_556800 == array_index_537262 ? add_556964 : sel_556961;
  assign add_556968 = sel_556965 + 8'h01;
  assign sel_556969 = array_index_556800 == array_index_537268 ? add_556968 : sel_556965;
  assign add_556972 = sel_556969 + 8'h01;
  assign sel_556973 = array_index_556800 == array_index_537274 ? add_556972 : sel_556969;
  assign add_556976 = sel_556973 + 8'h01;
  assign sel_556977 = array_index_556800 == array_index_537280 ? add_556976 : sel_556973;
  assign add_556980 = sel_556977 + 8'h01;
  assign sel_556981 = array_index_556800 == array_index_537286 ? add_556980 : sel_556977;
  assign add_556984 = sel_556981 + 8'h01;
  assign sel_556985 = array_index_556800 == array_index_537292 ? add_556984 : sel_556981;
  assign add_556988 = sel_556985 + 8'h01;
  assign sel_556989 = array_index_556800 == array_index_537298 ? add_556988 : sel_556985;
  assign add_556992 = sel_556989 + 8'h01;
  assign sel_556993 = array_index_556800 == array_index_537304 ? add_556992 : sel_556989;
  assign add_556996 = sel_556993 + 8'h01;
  assign sel_556997 = array_index_556800 == array_index_537310 ? add_556996 : sel_556993;
  assign add_557000 = sel_556997 + 8'h01;
  assign sel_557001 = array_index_556800 == array_index_537316 ? add_557000 : sel_556997;
  assign add_557004 = sel_557001 + 8'h01;
  assign sel_557005 = array_index_556800 == array_index_537322 ? add_557004 : sel_557001;
  assign add_557008 = sel_557005 + 8'h01;
  assign sel_557009 = array_index_556800 == array_index_537328 ? add_557008 : sel_557005;
  assign add_557012 = sel_557009 + 8'h01;
  assign sel_557013 = array_index_556800 == array_index_537334 ? add_557012 : sel_557009;
  assign add_557016 = sel_557013 + 8'h01;
  assign sel_557017 = array_index_556800 == array_index_537340 ? add_557016 : sel_557013;
  assign add_557020 = sel_557017 + 8'h01;
  assign sel_557021 = array_index_556800 == array_index_537346 ? add_557020 : sel_557017;
  assign add_557024 = sel_557021 + 8'h01;
  assign sel_557025 = array_index_556800 == array_index_537352 ? add_557024 : sel_557021;
  assign add_557028 = sel_557025 + 8'h01;
  assign sel_557029 = array_index_556800 == array_index_537358 ? add_557028 : sel_557025;
  assign add_557032 = sel_557029 + 8'h01;
  assign sel_557033 = array_index_556800 == array_index_537364 ? add_557032 : sel_557029;
  assign add_557036 = sel_557033 + 8'h01;
  assign sel_557037 = array_index_556800 == array_index_537370 ? add_557036 : sel_557033;
  assign add_557040 = sel_557037 + 8'h01;
  assign sel_557041 = array_index_556800 == array_index_537376 ? add_557040 : sel_557037;
  assign add_557044 = sel_557041 + 8'h01;
  assign sel_557045 = array_index_556800 == array_index_537382 ? add_557044 : sel_557041;
  assign add_557048 = sel_557045 + 8'h01;
  assign sel_557049 = array_index_556800 == array_index_537388 ? add_557048 : sel_557045;
  assign add_557052 = sel_557049 + 8'h01;
  assign sel_557053 = array_index_556800 == array_index_537394 ? add_557052 : sel_557049;
  assign add_557056 = sel_557053 + 8'h01;
  assign sel_557057 = array_index_556800 == array_index_537400 ? add_557056 : sel_557053;
  assign add_557060 = sel_557057 + 8'h01;
  assign sel_557061 = array_index_556800 == array_index_537406 ? add_557060 : sel_557057;
  assign add_557064 = sel_557061 + 8'h01;
  assign sel_557065 = array_index_556800 == array_index_537412 ? add_557064 : sel_557061;
  assign add_557068 = sel_557065 + 8'h01;
  assign sel_557069 = array_index_556800 == array_index_537418 ? add_557068 : sel_557065;
  assign add_557072 = sel_557069 + 8'h01;
  assign sel_557073 = array_index_556800 == array_index_537424 ? add_557072 : sel_557069;
  assign add_557076 = sel_557073 + 8'h01;
  assign sel_557077 = array_index_556800 == array_index_537430 ? add_557076 : sel_557073;
  assign add_557080 = sel_557077 + 8'h01;
  assign sel_557081 = array_index_556800 == array_index_537436 ? add_557080 : sel_557077;
  assign add_557084 = sel_557081 + 8'h01;
  assign sel_557085 = array_index_556800 == array_index_537442 ? add_557084 : sel_557081;
  assign add_557088 = sel_557085 + 8'h01;
  assign sel_557089 = array_index_556800 == array_index_537448 ? add_557088 : sel_557085;
  assign add_557092 = sel_557089 + 8'h01;
  assign sel_557093 = array_index_556800 == array_index_537454 ? add_557092 : sel_557089;
  assign add_557096 = sel_557093 + 8'h01;
  assign sel_557097 = array_index_556800 == array_index_537460 ? add_557096 : sel_557093;
  assign add_557101 = sel_557097 + 8'h01;
  assign array_index_557102 = set1_unflattened[7'h42];
  assign sel_557103 = array_index_556800 == array_index_537466 ? add_557101 : sel_557097;
  assign add_557106 = sel_557103 + 8'h01;
  assign sel_557107 = array_index_557102 == array_index_537012 ? add_557106 : sel_557103;
  assign add_557110 = sel_557107 + 8'h01;
  assign sel_557111 = array_index_557102 == array_index_537016 ? add_557110 : sel_557107;
  assign add_557114 = sel_557111 + 8'h01;
  assign sel_557115 = array_index_557102 == array_index_537024 ? add_557114 : sel_557111;
  assign add_557118 = sel_557115 + 8'h01;
  assign sel_557119 = array_index_557102 == array_index_537032 ? add_557118 : sel_557115;
  assign add_557122 = sel_557119 + 8'h01;
  assign sel_557123 = array_index_557102 == array_index_537040 ? add_557122 : sel_557119;
  assign add_557126 = sel_557123 + 8'h01;
  assign sel_557127 = array_index_557102 == array_index_537048 ? add_557126 : sel_557123;
  assign add_557130 = sel_557127 + 8'h01;
  assign sel_557131 = array_index_557102 == array_index_537056 ? add_557130 : sel_557127;
  assign add_557134 = sel_557131 + 8'h01;
  assign sel_557135 = array_index_557102 == array_index_537064 ? add_557134 : sel_557131;
  assign add_557138 = sel_557135 + 8'h01;
  assign sel_557139 = array_index_557102 == array_index_537070 ? add_557138 : sel_557135;
  assign add_557142 = sel_557139 + 8'h01;
  assign sel_557143 = array_index_557102 == array_index_537076 ? add_557142 : sel_557139;
  assign add_557146 = sel_557143 + 8'h01;
  assign sel_557147 = array_index_557102 == array_index_537082 ? add_557146 : sel_557143;
  assign add_557150 = sel_557147 + 8'h01;
  assign sel_557151 = array_index_557102 == array_index_537088 ? add_557150 : sel_557147;
  assign add_557154 = sel_557151 + 8'h01;
  assign sel_557155 = array_index_557102 == array_index_537094 ? add_557154 : sel_557151;
  assign add_557158 = sel_557155 + 8'h01;
  assign sel_557159 = array_index_557102 == array_index_537100 ? add_557158 : sel_557155;
  assign add_557162 = sel_557159 + 8'h01;
  assign sel_557163 = array_index_557102 == array_index_537106 ? add_557162 : sel_557159;
  assign add_557166 = sel_557163 + 8'h01;
  assign sel_557167 = array_index_557102 == array_index_537112 ? add_557166 : sel_557163;
  assign add_557170 = sel_557167 + 8'h01;
  assign sel_557171 = array_index_557102 == array_index_537118 ? add_557170 : sel_557167;
  assign add_557174 = sel_557171 + 8'h01;
  assign sel_557175 = array_index_557102 == array_index_537124 ? add_557174 : sel_557171;
  assign add_557178 = sel_557175 + 8'h01;
  assign sel_557179 = array_index_557102 == array_index_537130 ? add_557178 : sel_557175;
  assign add_557182 = sel_557179 + 8'h01;
  assign sel_557183 = array_index_557102 == array_index_537136 ? add_557182 : sel_557179;
  assign add_557186 = sel_557183 + 8'h01;
  assign sel_557187 = array_index_557102 == array_index_537142 ? add_557186 : sel_557183;
  assign add_557190 = sel_557187 + 8'h01;
  assign sel_557191 = array_index_557102 == array_index_537148 ? add_557190 : sel_557187;
  assign add_557194 = sel_557191 + 8'h01;
  assign sel_557195 = array_index_557102 == array_index_537154 ? add_557194 : sel_557191;
  assign add_557198 = sel_557195 + 8'h01;
  assign sel_557199 = array_index_557102 == array_index_537160 ? add_557198 : sel_557195;
  assign add_557202 = sel_557199 + 8'h01;
  assign sel_557203 = array_index_557102 == array_index_537166 ? add_557202 : sel_557199;
  assign add_557206 = sel_557203 + 8'h01;
  assign sel_557207 = array_index_557102 == array_index_537172 ? add_557206 : sel_557203;
  assign add_557210 = sel_557207 + 8'h01;
  assign sel_557211 = array_index_557102 == array_index_537178 ? add_557210 : sel_557207;
  assign add_557214 = sel_557211 + 8'h01;
  assign sel_557215 = array_index_557102 == array_index_537184 ? add_557214 : sel_557211;
  assign add_557218 = sel_557215 + 8'h01;
  assign sel_557219 = array_index_557102 == array_index_537190 ? add_557218 : sel_557215;
  assign add_557222 = sel_557219 + 8'h01;
  assign sel_557223 = array_index_557102 == array_index_537196 ? add_557222 : sel_557219;
  assign add_557226 = sel_557223 + 8'h01;
  assign sel_557227 = array_index_557102 == array_index_537202 ? add_557226 : sel_557223;
  assign add_557230 = sel_557227 + 8'h01;
  assign sel_557231 = array_index_557102 == array_index_537208 ? add_557230 : sel_557227;
  assign add_557234 = sel_557231 + 8'h01;
  assign sel_557235 = array_index_557102 == array_index_537214 ? add_557234 : sel_557231;
  assign add_557238 = sel_557235 + 8'h01;
  assign sel_557239 = array_index_557102 == array_index_537220 ? add_557238 : sel_557235;
  assign add_557242 = sel_557239 + 8'h01;
  assign sel_557243 = array_index_557102 == array_index_537226 ? add_557242 : sel_557239;
  assign add_557246 = sel_557243 + 8'h01;
  assign sel_557247 = array_index_557102 == array_index_537232 ? add_557246 : sel_557243;
  assign add_557250 = sel_557247 + 8'h01;
  assign sel_557251 = array_index_557102 == array_index_537238 ? add_557250 : sel_557247;
  assign add_557254 = sel_557251 + 8'h01;
  assign sel_557255 = array_index_557102 == array_index_537244 ? add_557254 : sel_557251;
  assign add_557258 = sel_557255 + 8'h01;
  assign sel_557259 = array_index_557102 == array_index_537250 ? add_557258 : sel_557255;
  assign add_557262 = sel_557259 + 8'h01;
  assign sel_557263 = array_index_557102 == array_index_537256 ? add_557262 : sel_557259;
  assign add_557266 = sel_557263 + 8'h01;
  assign sel_557267 = array_index_557102 == array_index_537262 ? add_557266 : sel_557263;
  assign add_557270 = sel_557267 + 8'h01;
  assign sel_557271 = array_index_557102 == array_index_537268 ? add_557270 : sel_557267;
  assign add_557274 = sel_557271 + 8'h01;
  assign sel_557275 = array_index_557102 == array_index_537274 ? add_557274 : sel_557271;
  assign add_557278 = sel_557275 + 8'h01;
  assign sel_557279 = array_index_557102 == array_index_537280 ? add_557278 : sel_557275;
  assign add_557282 = sel_557279 + 8'h01;
  assign sel_557283 = array_index_557102 == array_index_537286 ? add_557282 : sel_557279;
  assign add_557286 = sel_557283 + 8'h01;
  assign sel_557287 = array_index_557102 == array_index_537292 ? add_557286 : sel_557283;
  assign add_557290 = sel_557287 + 8'h01;
  assign sel_557291 = array_index_557102 == array_index_537298 ? add_557290 : sel_557287;
  assign add_557294 = sel_557291 + 8'h01;
  assign sel_557295 = array_index_557102 == array_index_537304 ? add_557294 : sel_557291;
  assign add_557298 = sel_557295 + 8'h01;
  assign sel_557299 = array_index_557102 == array_index_537310 ? add_557298 : sel_557295;
  assign add_557302 = sel_557299 + 8'h01;
  assign sel_557303 = array_index_557102 == array_index_537316 ? add_557302 : sel_557299;
  assign add_557306 = sel_557303 + 8'h01;
  assign sel_557307 = array_index_557102 == array_index_537322 ? add_557306 : sel_557303;
  assign add_557310 = sel_557307 + 8'h01;
  assign sel_557311 = array_index_557102 == array_index_537328 ? add_557310 : sel_557307;
  assign add_557314 = sel_557311 + 8'h01;
  assign sel_557315 = array_index_557102 == array_index_537334 ? add_557314 : sel_557311;
  assign add_557318 = sel_557315 + 8'h01;
  assign sel_557319 = array_index_557102 == array_index_537340 ? add_557318 : sel_557315;
  assign add_557322 = sel_557319 + 8'h01;
  assign sel_557323 = array_index_557102 == array_index_537346 ? add_557322 : sel_557319;
  assign add_557326 = sel_557323 + 8'h01;
  assign sel_557327 = array_index_557102 == array_index_537352 ? add_557326 : sel_557323;
  assign add_557330 = sel_557327 + 8'h01;
  assign sel_557331 = array_index_557102 == array_index_537358 ? add_557330 : sel_557327;
  assign add_557334 = sel_557331 + 8'h01;
  assign sel_557335 = array_index_557102 == array_index_537364 ? add_557334 : sel_557331;
  assign add_557338 = sel_557335 + 8'h01;
  assign sel_557339 = array_index_557102 == array_index_537370 ? add_557338 : sel_557335;
  assign add_557342 = sel_557339 + 8'h01;
  assign sel_557343 = array_index_557102 == array_index_537376 ? add_557342 : sel_557339;
  assign add_557346 = sel_557343 + 8'h01;
  assign sel_557347 = array_index_557102 == array_index_537382 ? add_557346 : sel_557343;
  assign add_557350 = sel_557347 + 8'h01;
  assign sel_557351 = array_index_557102 == array_index_537388 ? add_557350 : sel_557347;
  assign add_557354 = sel_557351 + 8'h01;
  assign sel_557355 = array_index_557102 == array_index_537394 ? add_557354 : sel_557351;
  assign add_557358 = sel_557355 + 8'h01;
  assign sel_557359 = array_index_557102 == array_index_537400 ? add_557358 : sel_557355;
  assign add_557362 = sel_557359 + 8'h01;
  assign sel_557363 = array_index_557102 == array_index_537406 ? add_557362 : sel_557359;
  assign add_557366 = sel_557363 + 8'h01;
  assign sel_557367 = array_index_557102 == array_index_537412 ? add_557366 : sel_557363;
  assign add_557370 = sel_557367 + 8'h01;
  assign sel_557371 = array_index_557102 == array_index_537418 ? add_557370 : sel_557367;
  assign add_557374 = sel_557371 + 8'h01;
  assign sel_557375 = array_index_557102 == array_index_537424 ? add_557374 : sel_557371;
  assign add_557378 = sel_557375 + 8'h01;
  assign sel_557379 = array_index_557102 == array_index_537430 ? add_557378 : sel_557375;
  assign add_557382 = sel_557379 + 8'h01;
  assign sel_557383 = array_index_557102 == array_index_537436 ? add_557382 : sel_557379;
  assign add_557386 = sel_557383 + 8'h01;
  assign sel_557387 = array_index_557102 == array_index_537442 ? add_557386 : sel_557383;
  assign add_557390 = sel_557387 + 8'h01;
  assign sel_557391 = array_index_557102 == array_index_537448 ? add_557390 : sel_557387;
  assign add_557394 = sel_557391 + 8'h01;
  assign sel_557395 = array_index_557102 == array_index_537454 ? add_557394 : sel_557391;
  assign add_557398 = sel_557395 + 8'h01;
  assign sel_557399 = array_index_557102 == array_index_537460 ? add_557398 : sel_557395;
  assign add_557403 = sel_557399 + 8'h01;
  assign array_index_557404 = set1_unflattened[7'h43];
  assign sel_557405 = array_index_557102 == array_index_537466 ? add_557403 : sel_557399;
  assign add_557408 = sel_557405 + 8'h01;
  assign sel_557409 = array_index_557404 == array_index_537012 ? add_557408 : sel_557405;
  assign add_557412 = sel_557409 + 8'h01;
  assign sel_557413 = array_index_557404 == array_index_537016 ? add_557412 : sel_557409;
  assign add_557416 = sel_557413 + 8'h01;
  assign sel_557417 = array_index_557404 == array_index_537024 ? add_557416 : sel_557413;
  assign add_557420 = sel_557417 + 8'h01;
  assign sel_557421 = array_index_557404 == array_index_537032 ? add_557420 : sel_557417;
  assign add_557424 = sel_557421 + 8'h01;
  assign sel_557425 = array_index_557404 == array_index_537040 ? add_557424 : sel_557421;
  assign add_557428 = sel_557425 + 8'h01;
  assign sel_557429 = array_index_557404 == array_index_537048 ? add_557428 : sel_557425;
  assign add_557432 = sel_557429 + 8'h01;
  assign sel_557433 = array_index_557404 == array_index_537056 ? add_557432 : sel_557429;
  assign add_557436 = sel_557433 + 8'h01;
  assign sel_557437 = array_index_557404 == array_index_537064 ? add_557436 : sel_557433;
  assign add_557440 = sel_557437 + 8'h01;
  assign sel_557441 = array_index_557404 == array_index_537070 ? add_557440 : sel_557437;
  assign add_557444 = sel_557441 + 8'h01;
  assign sel_557445 = array_index_557404 == array_index_537076 ? add_557444 : sel_557441;
  assign add_557448 = sel_557445 + 8'h01;
  assign sel_557449 = array_index_557404 == array_index_537082 ? add_557448 : sel_557445;
  assign add_557452 = sel_557449 + 8'h01;
  assign sel_557453 = array_index_557404 == array_index_537088 ? add_557452 : sel_557449;
  assign add_557456 = sel_557453 + 8'h01;
  assign sel_557457 = array_index_557404 == array_index_537094 ? add_557456 : sel_557453;
  assign add_557460 = sel_557457 + 8'h01;
  assign sel_557461 = array_index_557404 == array_index_537100 ? add_557460 : sel_557457;
  assign add_557464 = sel_557461 + 8'h01;
  assign sel_557465 = array_index_557404 == array_index_537106 ? add_557464 : sel_557461;
  assign add_557468 = sel_557465 + 8'h01;
  assign sel_557469 = array_index_557404 == array_index_537112 ? add_557468 : sel_557465;
  assign add_557472 = sel_557469 + 8'h01;
  assign sel_557473 = array_index_557404 == array_index_537118 ? add_557472 : sel_557469;
  assign add_557476 = sel_557473 + 8'h01;
  assign sel_557477 = array_index_557404 == array_index_537124 ? add_557476 : sel_557473;
  assign add_557480 = sel_557477 + 8'h01;
  assign sel_557481 = array_index_557404 == array_index_537130 ? add_557480 : sel_557477;
  assign add_557484 = sel_557481 + 8'h01;
  assign sel_557485 = array_index_557404 == array_index_537136 ? add_557484 : sel_557481;
  assign add_557488 = sel_557485 + 8'h01;
  assign sel_557489 = array_index_557404 == array_index_537142 ? add_557488 : sel_557485;
  assign add_557492 = sel_557489 + 8'h01;
  assign sel_557493 = array_index_557404 == array_index_537148 ? add_557492 : sel_557489;
  assign add_557496 = sel_557493 + 8'h01;
  assign sel_557497 = array_index_557404 == array_index_537154 ? add_557496 : sel_557493;
  assign add_557500 = sel_557497 + 8'h01;
  assign sel_557501 = array_index_557404 == array_index_537160 ? add_557500 : sel_557497;
  assign add_557504 = sel_557501 + 8'h01;
  assign sel_557505 = array_index_557404 == array_index_537166 ? add_557504 : sel_557501;
  assign add_557508 = sel_557505 + 8'h01;
  assign sel_557509 = array_index_557404 == array_index_537172 ? add_557508 : sel_557505;
  assign add_557512 = sel_557509 + 8'h01;
  assign sel_557513 = array_index_557404 == array_index_537178 ? add_557512 : sel_557509;
  assign add_557516 = sel_557513 + 8'h01;
  assign sel_557517 = array_index_557404 == array_index_537184 ? add_557516 : sel_557513;
  assign add_557520 = sel_557517 + 8'h01;
  assign sel_557521 = array_index_557404 == array_index_537190 ? add_557520 : sel_557517;
  assign add_557524 = sel_557521 + 8'h01;
  assign sel_557525 = array_index_557404 == array_index_537196 ? add_557524 : sel_557521;
  assign add_557528 = sel_557525 + 8'h01;
  assign sel_557529 = array_index_557404 == array_index_537202 ? add_557528 : sel_557525;
  assign add_557532 = sel_557529 + 8'h01;
  assign sel_557533 = array_index_557404 == array_index_537208 ? add_557532 : sel_557529;
  assign add_557536 = sel_557533 + 8'h01;
  assign sel_557537 = array_index_557404 == array_index_537214 ? add_557536 : sel_557533;
  assign add_557540 = sel_557537 + 8'h01;
  assign sel_557541 = array_index_557404 == array_index_537220 ? add_557540 : sel_557537;
  assign add_557544 = sel_557541 + 8'h01;
  assign sel_557545 = array_index_557404 == array_index_537226 ? add_557544 : sel_557541;
  assign add_557548 = sel_557545 + 8'h01;
  assign sel_557549 = array_index_557404 == array_index_537232 ? add_557548 : sel_557545;
  assign add_557552 = sel_557549 + 8'h01;
  assign sel_557553 = array_index_557404 == array_index_537238 ? add_557552 : sel_557549;
  assign add_557556 = sel_557553 + 8'h01;
  assign sel_557557 = array_index_557404 == array_index_537244 ? add_557556 : sel_557553;
  assign add_557560 = sel_557557 + 8'h01;
  assign sel_557561 = array_index_557404 == array_index_537250 ? add_557560 : sel_557557;
  assign add_557564 = sel_557561 + 8'h01;
  assign sel_557565 = array_index_557404 == array_index_537256 ? add_557564 : sel_557561;
  assign add_557568 = sel_557565 + 8'h01;
  assign sel_557569 = array_index_557404 == array_index_537262 ? add_557568 : sel_557565;
  assign add_557572 = sel_557569 + 8'h01;
  assign sel_557573 = array_index_557404 == array_index_537268 ? add_557572 : sel_557569;
  assign add_557576 = sel_557573 + 8'h01;
  assign sel_557577 = array_index_557404 == array_index_537274 ? add_557576 : sel_557573;
  assign add_557580 = sel_557577 + 8'h01;
  assign sel_557581 = array_index_557404 == array_index_537280 ? add_557580 : sel_557577;
  assign add_557584 = sel_557581 + 8'h01;
  assign sel_557585 = array_index_557404 == array_index_537286 ? add_557584 : sel_557581;
  assign add_557588 = sel_557585 + 8'h01;
  assign sel_557589 = array_index_557404 == array_index_537292 ? add_557588 : sel_557585;
  assign add_557592 = sel_557589 + 8'h01;
  assign sel_557593 = array_index_557404 == array_index_537298 ? add_557592 : sel_557589;
  assign add_557596 = sel_557593 + 8'h01;
  assign sel_557597 = array_index_557404 == array_index_537304 ? add_557596 : sel_557593;
  assign add_557600 = sel_557597 + 8'h01;
  assign sel_557601 = array_index_557404 == array_index_537310 ? add_557600 : sel_557597;
  assign add_557604 = sel_557601 + 8'h01;
  assign sel_557605 = array_index_557404 == array_index_537316 ? add_557604 : sel_557601;
  assign add_557608 = sel_557605 + 8'h01;
  assign sel_557609 = array_index_557404 == array_index_537322 ? add_557608 : sel_557605;
  assign add_557612 = sel_557609 + 8'h01;
  assign sel_557613 = array_index_557404 == array_index_537328 ? add_557612 : sel_557609;
  assign add_557616 = sel_557613 + 8'h01;
  assign sel_557617 = array_index_557404 == array_index_537334 ? add_557616 : sel_557613;
  assign add_557620 = sel_557617 + 8'h01;
  assign sel_557621 = array_index_557404 == array_index_537340 ? add_557620 : sel_557617;
  assign add_557624 = sel_557621 + 8'h01;
  assign sel_557625 = array_index_557404 == array_index_537346 ? add_557624 : sel_557621;
  assign add_557628 = sel_557625 + 8'h01;
  assign sel_557629 = array_index_557404 == array_index_537352 ? add_557628 : sel_557625;
  assign add_557632 = sel_557629 + 8'h01;
  assign sel_557633 = array_index_557404 == array_index_537358 ? add_557632 : sel_557629;
  assign add_557636 = sel_557633 + 8'h01;
  assign sel_557637 = array_index_557404 == array_index_537364 ? add_557636 : sel_557633;
  assign add_557640 = sel_557637 + 8'h01;
  assign sel_557641 = array_index_557404 == array_index_537370 ? add_557640 : sel_557637;
  assign add_557644 = sel_557641 + 8'h01;
  assign sel_557645 = array_index_557404 == array_index_537376 ? add_557644 : sel_557641;
  assign add_557648 = sel_557645 + 8'h01;
  assign sel_557649 = array_index_557404 == array_index_537382 ? add_557648 : sel_557645;
  assign add_557652 = sel_557649 + 8'h01;
  assign sel_557653 = array_index_557404 == array_index_537388 ? add_557652 : sel_557649;
  assign add_557656 = sel_557653 + 8'h01;
  assign sel_557657 = array_index_557404 == array_index_537394 ? add_557656 : sel_557653;
  assign add_557660 = sel_557657 + 8'h01;
  assign sel_557661 = array_index_557404 == array_index_537400 ? add_557660 : sel_557657;
  assign add_557664 = sel_557661 + 8'h01;
  assign sel_557665 = array_index_557404 == array_index_537406 ? add_557664 : sel_557661;
  assign add_557668 = sel_557665 + 8'h01;
  assign sel_557669 = array_index_557404 == array_index_537412 ? add_557668 : sel_557665;
  assign add_557672 = sel_557669 + 8'h01;
  assign sel_557673 = array_index_557404 == array_index_537418 ? add_557672 : sel_557669;
  assign add_557676 = sel_557673 + 8'h01;
  assign sel_557677 = array_index_557404 == array_index_537424 ? add_557676 : sel_557673;
  assign add_557680 = sel_557677 + 8'h01;
  assign sel_557681 = array_index_557404 == array_index_537430 ? add_557680 : sel_557677;
  assign add_557684 = sel_557681 + 8'h01;
  assign sel_557685 = array_index_557404 == array_index_537436 ? add_557684 : sel_557681;
  assign add_557688 = sel_557685 + 8'h01;
  assign sel_557689 = array_index_557404 == array_index_537442 ? add_557688 : sel_557685;
  assign add_557692 = sel_557689 + 8'h01;
  assign sel_557693 = array_index_557404 == array_index_537448 ? add_557692 : sel_557689;
  assign add_557696 = sel_557693 + 8'h01;
  assign sel_557697 = array_index_557404 == array_index_537454 ? add_557696 : sel_557693;
  assign add_557700 = sel_557697 + 8'h01;
  assign sel_557701 = array_index_557404 == array_index_537460 ? add_557700 : sel_557697;
  assign add_557705 = sel_557701 + 8'h01;
  assign array_index_557706 = set1_unflattened[7'h44];
  assign sel_557707 = array_index_557404 == array_index_537466 ? add_557705 : sel_557701;
  assign add_557710 = sel_557707 + 8'h01;
  assign sel_557711 = array_index_557706 == array_index_537012 ? add_557710 : sel_557707;
  assign add_557714 = sel_557711 + 8'h01;
  assign sel_557715 = array_index_557706 == array_index_537016 ? add_557714 : sel_557711;
  assign add_557718 = sel_557715 + 8'h01;
  assign sel_557719 = array_index_557706 == array_index_537024 ? add_557718 : sel_557715;
  assign add_557722 = sel_557719 + 8'h01;
  assign sel_557723 = array_index_557706 == array_index_537032 ? add_557722 : sel_557719;
  assign add_557726 = sel_557723 + 8'h01;
  assign sel_557727 = array_index_557706 == array_index_537040 ? add_557726 : sel_557723;
  assign add_557730 = sel_557727 + 8'h01;
  assign sel_557731 = array_index_557706 == array_index_537048 ? add_557730 : sel_557727;
  assign add_557734 = sel_557731 + 8'h01;
  assign sel_557735 = array_index_557706 == array_index_537056 ? add_557734 : sel_557731;
  assign add_557738 = sel_557735 + 8'h01;
  assign sel_557739 = array_index_557706 == array_index_537064 ? add_557738 : sel_557735;
  assign add_557742 = sel_557739 + 8'h01;
  assign sel_557743 = array_index_557706 == array_index_537070 ? add_557742 : sel_557739;
  assign add_557746 = sel_557743 + 8'h01;
  assign sel_557747 = array_index_557706 == array_index_537076 ? add_557746 : sel_557743;
  assign add_557750 = sel_557747 + 8'h01;
  assign sel_557751 = array_index_557706 == array_index_537082 ? add_557750 : sel_557747;
  assign add_557754 = sel_557751 + 8'h01;
  assign sel_557755 = array_index_557706 == array_index_537088 ? add_557754 : sel_557751;
  assign add_557758 = sel_557755 + 8'h01;
  assign sel_557759 = array_index_557706 == array_index_537094 ? add_557758 : sel_557755;
  assign add_557762 = sel_557759 + 8'h01;
  assign sel_557763 = array_index_557706 == array_index_537100 ? add_557762 : sel_557759;
  assign add_557766 = sel_557763 + 8'h01;
  assign sel_557767 = array_index_557706 == array_index_537106 ? add_557766 : sel_557763;
  assign add_557770 = sel_557767 + 8'h01;
  assign sel_557771 = array_index_557706 == array_index_537112 ? add_557770 : sel_557767;
  assign add_557774 = sel_557771 + 8'h01;
  assign sel_557775 = array_index_557706 == array_index_537118 ? add_557774 : sel_557771;
  assign add_557778 = sel_557775 + 8'h01;
  assign sel_557779 = array_index_557706 == array_index_537124 ? add_557778 : sel_557775;
  assign add_557782 = sel_557779 + 8'h01;
  assign sel_557783 = array_index_557706 == array_index_537130 ? add_557782 : sel_557779;
  assign add_557786 = sel_557783 + 8'h01;
  assign sel_557787 = array_index_557706 == array_index_537136 ? add_557786 : sel_557783;
  assign add_557790 = sel_557787 + 8'h01;
  assign sel_557791 = array_index_557706 == array_index_537142 ? add_557790 : sel_557787;
  assign add_557794 = sel_557791 + 8'h01;
  assign sel_557795 = array_index_557706 == array_index_537148 ? add_557794 : sel_557791;
  assign add_557798 = sel_557795 + 8'h01;
  assign sel_557799 = array_index_557706 == array_index_537154 ? add_557798 : sel_557795;
  assign add_557802 = sel_557799 + 8'h01;
  assign sel_557803 = array_index_557706 == array_index_537160 ? add_557802 : sel_557799;
  assign add_557806 = sel_557803 + 8'h01;
  assign sel_557807 = array_index_557706 == array_index_537166 ? add_557806 : sel_557803;
  assign add_557810 = sel_557807 + 8'h01;
  assign sel_557811 = array_index_557706 == array_index_537172 ? add_557810 : sel_557807;
  assign add_557814 = sel_557811 + 8'h01;
  assign sel_557815 = array_index_557706 == array_index_537178 ? add_557814 : sel_557811;
  assign add_557818 = sel_557815 + 8'h01;
  assign sel_557819 = array_index_557706 == array_index_537184 ? add_557818 : sel_557815;
  assign add_557822 = sel_557819 + 8'h01;
  assign sel_557823 = array_index_557706 == array_index_537190 ? add_557822 : sel_557819;
  assign add_557826 = sel_557823 + 8'h01;
  assign sel_557827 = array_index_557706 == array_index_537196 ? add_557826 : sel_557823;
  assign add_557830 = sel_557827 + 8'h01;
  assign sel_557831 = array_index_557706 == array_index_537202 ? add_557830 : sel_557827;
  assign add_557834 = sel_557831 + 8'h01;
  assign sel_557835 = array_index_557706 == array_index_537208 ? add_557834 : sel_557831;
  assign add_557838 = sel_557835 + 8'h01;
  assign sel_557839 = array_index_557706 == array_index_537214 ? add_557838 : sel_557835;
  assign add_557842 = sel_557839 + 8'h01;
  assign sel_557843 = array_index_557706 == array_index_537220 ? add_557842 : sel_557839;
  assign add_557846 = sel_557843 + 8'h01;
  assign sel_557847 = array_index_557706 == array_index_537226 ? add_557846 : sel_557843;
  assign add_557850 = sel_557847 + 8'h01;
  assign sel_557851 = array_index_557706 == array_index_537232 ? add_557850 : sel_557847;
  assign add_557854 = sel_557851 + 8'h01;
  assign sel_557855 = array_index_557706 == array_index_537238 ? add_557854 : sel_557851;
  assign add_557858 = sel_557855 + 8'h01;
  assign sel_557859 = array_index_557706 == array_index_537244 ? add_557858 : sel_557855;
  assign add_557862 = sel_557859 + 8'h01;
  assign sel_557863 = array_index_557706 == array_index_537250 ? add_557862 : sel_557859;
  assign add_557866 = sel_557863 + 8'h01;
  assign sel_557867 = array_index_557706 == array_index_537256 ? add_557866 : sel_557863;
  assign add_557870 = sel_557867 + 8'h01;
  assign sel_557871 = array_index_557706 == array_index_537262 ? add_557870 : sel_557867;
  assign add_557874 = sel_557871 + 8'h01;
  assign sel_557875 = array_index_557706 == array_index_537268 ? add_557874 : sel_557871;
  assign add_557878 = sel_557875 + 8'h01;
  assign sel_557879 = array_index_557706 == array_index_537274 ? add_557878 : sel_557875;
  assign add_557882 = sel_557879 + 8'h01;
  assign sel_557883 = array_index_557706 == array_index_537280 ? add_557882 : sel_557879;
  assign add_557886 = sel_557883 + 8'h01;
  assign sel_557887 = array_index_557706 == array_index_537286 ? add_557886 : sel_557883;
  assign add_557890 = sel_557887 + 8'h01;
  assign sel_557891 = array_index_557706 == array_index_537292 ? add_557890 : sel_557887;
  assign add_557894 = sel_557891 + 8'h01;
  assign sel_557895 = array_index_557706 == array_index_537298 ? add_557894 : sel_557891;
  assign add_557898 = sel_557895 + 8'h01;
  assign sel_557899 = array_index_557706 == array_index_537304 ? add_557898 : sel_557895;
  assign add_557902 = sel_557899 + 8'h01;
  assign sel_557903 = array_index_557706 == array_index_537310 ? add_557902 : sel_557899;
  assign add_557906 = sel_557903 + 8'h01;
  assign sel_557907 = array_index_557706 == array_index_537316 ? add_557906 : sel_557903;
  assign add_557910 = sel_557907 + 8'h01;
  assign sel_557911 = array_index_557706 == array_index_537322 ? add_557910 : sel_557907;
  assign add_557914 = sel_557911 + 8'h01;
  assign sel_557915 = array_index_557706 == array_index_537328 ? add_557914 : sel_557911;
  assign add_557918 = sel_557915 + 8'h01;
  assign sel_557919 = array_index_557706 == array_index_537334 ? add_557918 : sel_557915;
  assign add_557922 = sel_557919 + 8'h01;
  assign sel_557923 = array_index_557706 == array_index_537340 ? add_557922 : sel_557919;
  assign add_557926 = sel_557923 + 8'h01;
  assign sel_557927 = array_index_557706 == array_index_537346 ? add_557926 : sel_557923;
  assign add_557930 = sel_557927 + 8'h01;
  assign sel_557931 = array_index_557706 == array_index_537352 ? add_557930 : sel_557927;
  assign add_557934 = sel_557931 + 8'h01;
  assign sel_557935 = array_index_557706 == array_index_537358 ? add_557934 : sel_557931;
  assign add_557938 = sel_557935 + 8'h01;
  assign sel_557939 = array_index_557706 == array_index_537364 ? add_557938 : sel_557935;
  assign add_557942 = sel_557939 + 8'h01;
  assign sel_557943 = array_index_557706 == array_index_537370 ? add_557942 : sel_557939;
  assign add_557946 = sel_557943 + 8'h01;
  assign sel_557947 = array_index_557706 == array_index_537376 ? add_557946 : sel_557943;
  assign add_557950 = sel_557947 + 8'h01;
  assign sel_557951 = array_index_557706 == array_index_537382 ? add_557950 : sel_557947;
  assign add_557954 = sel_557951 + 8'h01;
  assign sel_557955 = array_index_557706 == array_index_537388 ? add_557954 : sel_557951;
  assign add_557958 = sel_557955 + 8'h01;
  assign sel_557959 = array_index_557706 == array_index_537394 ? add_557958 : sel_557955;
  assign add_557962 = sel_557959 + 8'h01;
  assign sel_557963 = array_index_557706 == array_index_537400 ? add_557962 : sel_557959;
  assign add_557966 = sel_557963 + 8'h01;
  assign sel_557967 = array_index_557706 == array_index_537406 ? add_557966 : sel_557963;
  assign add_557970 = sel_557967 + 8'h01;
  assign sel_557971 = array_index_557706 == array_index_537412 ? add_557970 : sel_557967;
  assign add_557974 = sel_557971 + 8'h01;
  assign sel_557975 = array_index_557706 == array_index_537418 ? add_557974 : sel_557971;
  assign add_557978 = sel_557975 + 8'h01;
  assign sel_557979 = array_index_557706 == array_index_537424 ? add_557978 : sel_557975;
  assign add_557982 = sel_557979 + 8'h01;
  assign sel_557983 = array_index_557706 == array_index_537430 ? add_557982 : sel_557979;
  assign add_557986 = sel_557983 + 8'h01;
  assign sel_557987 = array_index_557706 == array_index_537436 ? add_557986 : sel_557983;
  assign add_557990 = sel_557987 + 8'h01;
  assign sel_557991 = array_index_557706 == array_index_537442 ? add_557990 : sel_557987;
  assign add_557994 = sel_557991 + 8'h01;
  assign sel_557995 = array_index_557706 == array_index_537448 ? add_557994 : sel_557991;
  assign add_557998 = sel_557995 + 8'h01;
  assign sel_557999 = array_index_557706 == array_index_537454 ? add_557998 : sel_557995;
  assign add_558002 = sel_557999 + 8'h01;
  assign sel_558003 = array_index_557706 == array_index_537460 ? add_558002 : sel_557999;
  assign add_558007 = sel_558003 + 8'h01;
  assign array_index_558008 = set1_unflattened[7'h45];
  assign sel_558009 = array_index_557706 == array_index_537466 ? add_558007 : sel_558003;
  assign add_558012 = sel_558009 + 8'h01;
  assign sel_558013 = array_index_558008 == array_index_537012 ? add_558012 : sel_558009;
  assign add_558016 = sel_558013 + 8'h01;
  assign sel_558017 = array_index_558008 == array_index_537016 ? add_558016 : sel_558013;
  assign add_558020 = sel_558017 + 8'h01;
  assign sel_558021 = array_index_558008 == array_index_537024 ? add_558020 : sel_558017;
  assign add_558024 = sel_558021 + 8'h01;
  assign sel_558025 = array_index_558008 == array_index_537032 ? add_558024 : sel_558021;
  assign add_558028 = sel_558025 + 8'h01;
  assign sel_558029 = array_index_558008 == array_index_537040 ? add_558028 : sel_558025;
  assign add_558032 = sel_558029 + 8'h01;
  assign sel_558033 = array_index_558008 == array_index_537048 ? add_558032 : sel_558029;
  assign add_558036 = sel_558033 + 8'h01;
  assign sel_558037 = array_index_558008 == array_index_537056 ? add_558036 : sel_558033;
  assign add_558040 = sel_558037 + 8'h01;
  assign sel_558041 = array_index_558008 == array_index_537064 ? add_558040 : sel_558037;
  assign add_558044 = sel_558041 + 8'h01;
  assign sel_558045 = array_index_558008 == array_index_537070 ? add_558044 : sel_558041;
  assign add_558048 = sel_558045 + 8'h01;
  assign sel_558049 = array_index_558008 == array_index_537076 ? add_558048 : sel_558045;
  assign add_558052 = sel_558049 + 8'h01;
  assign sel_558053 = array_index_558008 == array_index_537082 ? add_558052 : sel_558049;
  assign add_558056 = sel_558053 + 8'h01;
  assign sel_558057 = array_index_558008 == array_index_537088 ? add_558056 : sel_558053;
  assign add_558060 = sel_558057 + 8'h01;
  assign sel_558061 = array_index_558008 == array_index_537094 ? add_558060 : sel_558057;
  assign add_558064 = sel_558061 + 8'h01;
  assign sel_558065 = array_index_558008 == array_index_537100 ? add_558064 : sel_558061;
  assign add_558068 = sel_558065 + 8'h01;
  assign sel_558069 = array_index_558008 == array_index_537106 ? add_558068 : sel_558065;
  assign add_558072 = sel_558069 + 8'h01;
  assign sel_558073 = array_index_558008 == array_index_537112 ? add_558072 : sel_558069;
  assign add_558076 = sel_558073 + 8'h01;
  assign sel_558077 = array_index_558008 == array_index_537118 ? add_558076 : sel_558073;
  assign add_558080 = sel_558077 + 8'h01;
  assign sel_558081 = array_index_558008 == array_index_537124 ? add_558080 : sel_558077;
  assign add_558084 = sel_558081 + 8'h01;
  assign sel_558085 = array_index_558008 == array_index_537130 ? add_558084 : sel_558081;
  assign add_558088 = sel_558085 + 8'h01;
  assign sel_558089 = array_index_558008 == array_index_537136 ? add_558088 : sel_558085;
  assign add_558092 = sel_558089 + 8'h01;
  assign sel_558093 = array_index_558008 == array_index_537142 ? add_558092 : sel_558089;
  assign add_558096 = sel_558093 + 8'h01;
  assign sel_558097 = array_index_558008 == array_index_537148 ? add_558096 : sel_558093;
  assign add_558100 = sel_558097 + 8'h01;
  assign sel_558101 = array_index_558008 == array_index_537154 ? add_558100 : sel_558097;
  assign add_558104 = sel_558101 + 8'h01;
  assign sel_558105 = array_index_558008 == array_index_537160 ? add_558104 : sel_558101;
  assign add_558108 = sel_558105 + 8'h01;
  assign sel_558109 = array_index_558008 == array_index_537166 ? add_558108 : sel_558105;
  assign add_558112 = sel_558109 + 8'h01;
  assign sel_558113 = array_index_558008 == array_index_537172 ? add_558112 : sel_558109;
  assign add_558116 = sel_558113 + 8'h01;
  assign sel_558117 = array_index_558008 == array_index_537178 ? add_558116 : sel_558113;
  assign add_558120 = sel_558117 + 8'h01;
  assign sel_558121 = array_index_558008 == array_index_537184 ? add_558120 : sel_558117;
  assign add_558124 = sel_558121 + 8'h01;
  assign sel_558125 = array_index_558008 == array_index_537190 ? add_558124 : sel_558121;
  assign add_558128 = sel_558125 + 8'h01;
  assign sel_558129 = array_index_558008 == array_index_537196 ? add_558128 : sel_558125;
  assign add_558132 = sel_558129 + 8'h01;
  assign sel_558133 = array_index_558008 == array_index_537202 ? add_558132 : sel_558129;
  assign add_558136 = sel_558133 + 8'h01;
  assign sel_558137 = array_index_558008 == array_index_537208 ? add_558136 : sel_558133;
  assign add_558140 = sel_558137 + 8'h01;
  assign sel_558141 = array_index_558008 == array_index_537214 ? add_558140 : sel_558137;
  assign add_558144 = sel_558141 + 8'h01;
  assign sel_558145 = array_index_558008 == array_index_537220 ? add_558144 : sel_558141;
  assign add_558148 = sel_558145 + 8'h01;
  assign sel_558149 = array_index_558008 == array_index_537226 ? add_558148 : sel_558145;
  assign add_558152 = sel_558149 + 8'h01;
  assign sel_558153 = array_index_558008 == array_index_537232 ? add_558152 : sel_558149;
  assign add_558156 = sel_558153 + 8'h01;
  assign sel_558157 = array_index_558008 == array_index_537238 ? add_558156 : sel_558153;
  assign add_558160 = sel_558157 + 8'h01;
  assign sel_558161 = array_index_558008 == array_index_537244 ? add_558160 : sel_558157;
  assign add_558164 = sel_558161 + 8'h01;
  assign sel_558165 = array_index_558008 == array_index_537250 ? add_558164 : sel_558161;
  assign add_558168 = sel_558165 + 8'h01;
  assign sel_558169 = array_index_558008 == array_index_537256 ? add_558168 : sel_558165;
  assign add_558172 = sel_558169 + 8'h01;
  assign sel_558173 = array_index_558008 == array_index_537262 ? add_558172 : sel_558169;
  assign add_558176 = sel_558173 + 8'h01;
  assign sel_558177 = array_index_558008 == array_index_537268 ? add_558176 : sel_558173;
  assign add_558180 = sel_558177 + 8'h01;
  assign sel_558181 = array_index_558008 == array_index_537274 ? add_558180 : sel_558177;
  assign add_558184 = sel_558181 + 8'h01;
  assign sel_558185 = array_index_558008 == array_index_537280 ? add_558184 : sel_558181;
  assign add_558188 = sel_558185 + 8'h01;
  assign sel_558189 = array_index_558008 == array_index_537286 ? add_558188 : sel_558185;
  assign add_558192 = sel_558189 + 8'h01;
  assign sel_558193 = array_index_558008 == array_index_537292 ? add_558192 : sel_558189;
  assign add_558196 = sel_558193 + 8'h01;
  assign sel_558197 = array_index_558008 == array_index_537298 ? add_558196 : sel_558193;
  assign add_558200 = sel_558197 + 8'h01;
  assign sel_558201 = array_index_558008 == array_index_537304 ? add_558200 : sel_558197;
  assign add_558204 = sel_558201 + 8'h01;
  assign sel_558205 = array_index_558008 == array_index_537310 ? add_558204 : sel_558201;
  assign add_558208 = sel_558205 + 8'h01;
  assign sel_558209 = array_index_558008 == array_index_537316 ? add_558208 : sel_558205;
  assign add_558212 = sel_558209 + 8'h01;
  assign sel_558213 = array_index_558008 == array_index_537322 ? add_558212 : sel_558209;
  assign add_558216 = sel_558213 + 8'h01;
  assign sel_558217 = array_index_558008 == array_index_537328 ? add_558216 : sel_558213;
  assign add_558220 = sel_558217 + 8'h01;
  assign sel_558221 = array_index_558008 == array_index_537334 ? add_558220 : sel_558217;
  assign add_558224 = sel_558221 + 8'h01;
  assign sel_558225 = array_index_558008 == array_index_537340 ? add_558224 : sel_558221;
  assign add_558228 = sel_558225 + 8'h01;
  assign sel_558229 = array_index_558008 == array_index_537346 ? add_558228 : sel_558225;
  assign add_558232 = sel_558229 + 8'h01;
  assign sel_558233 = array_index_558008 == array_index_537352 ? add_558232 : sel_558229;
  assign add_558236 = sel_558233 + 8'h01;
  assign sel_558237 = array_index_558008 == array_index_537358 ? add_558236 : sel_558233;
  assign add_558240 = sel_558237 + 8'h01;
  assign sel_558241 = array_index_558008 == array_index_537364 ? add_558240 : sel_558237;
  assign add_558244 = sel_558241 + 8'h01;
  assign sel_558245 = array_index_558008 == array_index_537370 ? add_558244 : sel_558241;
  assign add_558248 = sel_558245 + 8'h01;
  assign sel_558249 = array_index_558008 == array_index_537376 ? add_558248 : sel_558245;
  assign add_558252 = sel_558249 + 8'h01;
  assign sel_558253 = array_index_558008 == array_index_537382 ? add_558252 : sel_558249;
  assign add_558256 = sel_558253 + 8'h01;
  assign sel_558257 = array_index_558008 == array_index_537388 ? add_558256 : sel_558253;
  assign add_558260 = sel_558257 + 8'h01;
  assign sel_558261 = array_index_558008 == array_index_537394 ? add_558260 : sel_558257;
  assign add_558264 = sel_558261 + 8'h01;
  assign sel_558265 = array_index_558008 == array_index_537400 ? add_558264 : sel_558261;
  assign add_558268 = sel_558265 + 8'h01;
  assign sel_558269 = array_index_558008 == array_index_537406 ? add_558268 : sel_558265;
  assign add_558272 = sel_558269 + 8'h01;
  assign sel_558273 = array_index_558008 == array_index_537412 ? add_558272 : sel_558269;
  assign add_558276 = sel_558273 + 8'h01;
  assign sel_558277 = array_index_558008 == array_index_537418 ? add_558276 : sel_558273;
  assign add_558280 = sel_558277 + 8'h01;
  assign sel_558281 = array_index_558008 == array_index_537424 ? add_558280 : sel_558277;
  assign add_558284 = sel_558281 + 8'h01;
  assign sel_558285 = array_index_558008 == array_index_537430 ? add_558284 : sel_558281;
  assign add_558288 = sel_558285 + 8'h01;
  assign sel_558289 = array_index_558008 == array_index_537436 ? add_558288 : sel_558285;
  assign add_558292 = sel_558289 + 8'h01;
  assign sel_558293 = array_index_558008 == array_index_537442 ? add_558292 : sel_558289;
  assign add_558296 = sel_558293 + 8'h01;
  assign sel_558297 = array_index_558008 == array_index_537448 ? add_558296 : sel_558293;
  assign add_558300 = sel_558297 + 8'h01;
  assign sel_558301 = array_index_558008 == array_index_537454 ? add_558300 : sel_558297;
  assign add_558304 = sel_558301 + 8'h01;
  assign sel_558305 = array_index_558008 == array_index_537460 ? add_558304 : sel_558301;
  assign add_558309 = sel_558305 + 8'h01;
  assign array_index_558310 = set1_unflattened[7'h46];
  assign sel_558311 = array_index_558008 == array_index_537466 ? add_558309 : sel_558305;
  assign add_558314 = sel_558311 + 8'h01;
  assign sel_558315 = array_index_558310 == array_index_537012 ? add_558314 : sel_558311;
  assign add_558318 = sel_558315 + 8'h01;
  assign sel_558319 = array_index_558310 == array_index_537016 ? add_558318 : sel_558315;
  assign add_558322 = sel_558319 + 8'h01;
  assign sel_558323 = array_index_558310 == array_index_537024 ? add_558322 : sel_558319;
  assign add_558326 = sel_558323 + 8'h01;
  assign sel_558327 = array_index_558310 == array_index_537032 ? add_558326 : sel_558323;
  assign add_558330 = sel_558327 + 8'h01;
  assign sel_558331 = array_index_558310 == array_index_537040 ? add_558330 : sel_558327;
  assign add_558334 = sel_558331 + 8'h01;
  assign sel_558335 = array_index_558310 == array_index_537048 ? add_558334 : sel_558331;
  assign add_558338 = sel_558335 + 8'h01;
  assign sel_558339 = array_index_558310 == array_index_537056 ? add_558338 : sel_558335;
  assign add_558342 = sel_558339 + 8'h01;
  assign sel_558343 = array_index_558310 == array_index_537064 ? add_558342 : sel_558339;
  assign add_558346 = sel_558343 + 8'h01;
  assign sel_558347 = array_index_558310 == array_index_537070 ? add_558346 : sel_558343;
  assign add_558350 = sel_558347 + 8'h01;
  assign sel_558351 = array_index_558310 == array_index_537076 ? add_558350 : sel_558347;
  assign add_558354 = sel_558351 + 8'h01;
  assign sel_558355 = array_index_558310 == array_index_537082 ? add_558354 : sel_558351;
  assign add_558358 = sel_558355 + 8'h01;
  assign sel_558359 = array_index_558310 == array_index_537088 ? add_558358 : sel_558355;
  assign add_558362 = sel_558359 + 8'h01;
  assign sel_558363 = array_index_558310 == array_index_537094 ? add_558362 : sel_558359;
  assign add_558366 = sel_558363 + 8'h01;
  assign sel_558367 = array_index_558310 == array_index_537100 ? add_558366 : sel_558363;
  assign add_558370 = sel_558367 + 8'h01;
  assign sel_558371 = array_index_558310 == array_index_537106 ? add_558370 : sel_558367;
  assign add_558374 = sel_558371 + 8'h01;
  assign sel_558375 = array_index_558310 == array_index_537112 ? add_558374 : sel_558371;
  assign add_558378 = sel_558375 + 8'h01;
  assign sel_558379 = array_index_558310 == array_index_537118 ? add_558378 : sel_558375;
  assign add_558382 = sel_558379 + 8'h01;
  assign sel_558383 = array_index_558310 == array_index_537124 ? add_558382 : sel_558379;
  assign add_558386 = sel_558383 + 8'h01;
  assign sel_558387 = array_index_558310 == array_index_537130 ? add_558386 : sel_558383;
  assign add_558390 = sel_558387 + 8'h01;
  assign sel_558391 = array_index_558310 == array_index_537136 ? add_558390 : sel_558387;
  assign add_558394 = sel_558391 + 8'h01;
  assign sel_558395 = array_index_558310 == array_index_537142 ? add_558394 : sel_558391;
  assign add_558398 = sel_558395 + 8'h01;
  assign sel_558399 = array_index_558310 == array_index_537148 ? add_558398 : sel_558395;
  assign add_558402 = sel_558399 + 8'h01;
  assign sel_558403 = array_index_558310 == array_index_537154 ? add_558402 : sel_558399;
  assign add_558406 = sel_558403 + 8'h01;
  assign sel_558407 = array_index_558310 == array_index_537160 ? add_558406 : sel_558403;
  assign add_558410 = sel_558407 + 8'h01;
  assign sel_558411 = array_index_558310 == array_index_537166 ? add_558410 : sel_558407;
  assign add_558414 = sel_558411 + 8'h01;
  assign sel_558415 = array_index_558310 == array_index_537172 ? add_558414 : sel_558411;
  assign add_558418 = sel_558415 + 8'h01;
  assign sel_558419 = array_index_558310 == array_index_537178 ? add_558418 : sel_558415;
  assign add_558422 = sel_558419 + 8'h01;
  assign sel_558423 = array_index_558310 == array_index_537184 ? add_558422 : sel_558419;
  assign add_558426 = sel_558423 + 8'h01;
  assign sel_558427 = array_index_558310 == array_index_537190 ? add_558426 : sel_558423;
  assign add_558430 = sel_558427 + 8'h01;
  assign sel_558431 = array_index_558310 == array_index_537196 ? add_558430 : sel_558427;
  assign add_558434 = sel_558431 + 8'h01;
  assign sel_558435 = array_index_558310 == array_index_537202 ? add_558434 : sel_558431;
  assign add_558438 = sel_558435 + 8'h01;
  assign sel_558439 = array_index_558310 == array_index_537208 ? add_558438 : sel_558435;
  assign add_558442 = sel_558439 + 8'h01;
  assign sel_558443 = array_index_558310 == array_index_537214 ? add_558442 : sel_558439;
  assign add_558446 = sel_558443 + 8'h01;
  assign sel_558447 = array_index_558310 == array_index_537220 ? add_558446 : sel_558443;
  assign add_558450 = sel_558447 + 8'h01;
  assign sel_558451 = array_index_558310 == array_index_537226 ? add_558450 : sel_558447;
  assign add_558454 = sel_558451 + 8'h01;
  assign sel_558455 = array_index_558310 == array_index_537232 ? add_558454 : sel_558451;
  assign add_558458 = sel_558455 + 8'h01;
  assign sel_558459 = array_index_558310 == array_index_537238 ? add_558458 : sel_558455;
  assign add_558462 = sel_558459 + 8'h01;
  assign sel_558463 = array_index_558310 == array_index_537244 ? add_558462 : sel_558459;
  assign add_558466 = sel_558463 + 8'h01;
  assign sel_558467 = array_index_558310 == array_index_537250 ? add_558466 : sel_558463;
  assign add_558470 = sel_558467 + 8'h01;
  assign sel_558471 = array_index_558310 == array_index_537256 ? add_558470 : sel_558467;
  assign add_558474 = sel_558471 + 8'h01;
  assign sel_558475 = array_index_558310 == array_index_537262 ? add_558474 : sel_558471;
  assign add_558478 = sel_558475 + 8'h01;
  assign sel_558479 = array_index_558310 == array_index_537268 ? add_558478 : sel_558475;
  assign add_558482 = sel_558479 + 8'h01;
  assign sel_558483 = array_index_558310 == array_index_537274 ? add_558482 : sel_558479;
  assign add_558486 = sel_558483 + 8'h01;
  assign sel_558487 = array_index_558310 == array_index_537280 ? add_558486 : sel_558483;
  assign add_558490 = sel_558487 + 8'h01;
  assign sel_558491 = array_index_558310 == array_index_537286 ? add_558490 : sel_558487;
  assign add_558494 = sel_558491 + 8'h01;
  assign sel_558495 = array_index_558310 == array_index_537292 ? add_558494 : sel_558491;
  assign add_558498 = sel_558495 + 8'h01;
  assign sel_558499 = array_index_558310 == array_index_537298 ? add_558498 : sel_558495;
  assign add_558502 = sel_558499 + 8'h01;
  assign sel_558503 = array_index_558310 == array_index_537304 ? add_558502 : sel_558499;
  assign add_558506 = sel_558503 + 8'h01;
  assign sel_558507 = array_index_558310 == array_index_537310 ? add_558506 : sel_558503;
  assign add_558510 = sel_558507 + 8'h01;
  assign sel_558511 = array_index_558310 == array_index_537316 ? add_558510 : sel_558507;
  assign add_558514 = sel_558511 + 8'h01;
  assign sel_558515 = array_index_558310 == array_index_537322 ? add_558514 : sel_558511;
  assign add_558518 = sel_558515 + 8'h01;
  assign sel_558519 = array_index_558310 == array_index_537328 ? add_558518 : sel_558515;
  assign add_558522 = sel_558519 + 8'h01;
  assign sel_558523 = array_index_558310 == array_index_537334 ? add_558522 : sel_558519;
  assign add_558526 = sel_558523 + 8'h01;
  assign sel_558527 = array_index_558310 == array_index_537340 ? add_558526 : sel_558523;
  assign add_558530 = sel_558527 + 8'h01;
  assign sel_558531 = array_index_558310 == array_index_537346 ? add_558530 : sel_558527;
  assign add_558534 = sel_558531 + 8'h01;
  assign sel_558535 = array_index_558310 == array_index_537352 ? add_558534 : sel_558531;
  assign add_558538 = sel_558535 + 8'h01;
  assign sel_558539 = array_index_558310 == array_index_537358 ? add_558538 : sel_558535;
  assign add_558542 = sel_558539 + 8'h01;
  assign sel_558543 = array_index_558310 == array_index_537364 ? add_558542 : sel_558539;
  assign add_558546 = sel_558543 + 8'h01;
  assign sel_558547 = array_index_558310 == array_index_537370 ? add_558546 : sel_558543;
  assign add_558550 = sel_558547 + 8'h01;
  assign sel_558551 = array_index_558310 == array_index_537376 ? add_558550 : sel_558547;
  assign add_558554 = sel_558551 + 8'h01;
  assign sel_558555 = array_index_558310 == array_index_537382 ? add_558554 : sel_558551;
  assign add_558558 = sel_558555 + 8'h01;
  assign sel_558559 = array_index_558310 == array_index_537388 ? add_558558 : sel_558555;
  assign add_558562 = sel_558559 + 8'h01;
  assign sel_558563 = array_index_558310 == array_index_537394 ? add_558562 : sel_558559;
  assign add_558566 = sel_558563 + 8'h01;
  assign sel_558567 = array_index_558310 == array_index_537400 ? add_558566 : sel_558563;
  assign add_558570 = sel_558567 + 8'h01;
  assign sel_558571 = array_index_558310 == array_index_537406 ? add_558570 : sel_558567;
  assign add_558574 = sel_558571 + 8'h01;
  assign sel_558575 = array_index_558310 == array_index_537412 ? add_558574 : sel_558571;
  assign add_558578 = sel_558575 + 8'h01;
  assign sel_558579 = array_index_558310 == array_index_537418 ? add_558578 : sel_558575;
  assign add_558582 = sel_558579 + 8'h01;
  assign sel_558583 = array_index_558310 == array_index_537424 ? add_558582 : sel_558579;
  assign add_558586 = sel_558583 + 8'h01;
  assign sel_558587 = array_index_558310 == array_index_537430 ? add_558586 : sel_558583;
  assign add_558590 = sel_558587 + 8'h01;
  assign sel_558591 = array_index_558310 == array_index_537436 ? add_558590 : sel_558587;
  assign add_558594 = sel_558591 + 8'h01;
  assign sel_558595 = array_index_558310 == array_index_537442 ? add_558594 : sel_558591;
  assign add_558598 = sel_558595 + 8'h01;
  assign sel_558599 = array_index_558310 == array_index_537448 ? add_558598 : sel_558595;
  assign add_558602 = sel_558599 + 8'h01;
  assign sel_558603 = array_index_558310 == array_index_537454 ? add_558602 : sel_558599;
  assign add_558606 = sel_558603 + 8'h01;
  assign sel_558607 = array_index_558310 == array_index_537460 ? add_558606 : sel_558603;
  assign add_558611 = sel_558607 + 8'h01;
  assign array_index_558612 = set1_unflattened[7'h47];
  assign sel_558613 = array_index_558310 == array_index_537466 ? add_558611 : sel_558607;
  assign add_558616 = sel_558613 + 8'h01;
  assign sel_558617 = array_index_558612 == array_index_537012 ? add_558616 : sel_558613;
  assign add_558620 = sel_558617 + 8'h01;
  assign sel_558621 = array_index_558612 == array_index_537016 ? add_558620 : sel_558617;
  assign add_558624 = sel_558621 + 8'h01;
  assign sel_558625 = array_index_558612 == array_index_537024 ? add_558624 : sel_558621;
  assign add_558628 = sel_558625 + 8'h01;
  assign sel_558629 = array_index_558612 == array_index_537032 ? add_558628 : sel_558625;
  assign add_558632 = sel_558629 + 8'h01;
  assign sel_558633 = array_index_558612 == array_index_537040 ? add_558632 : sel_558629;
  assign add_558636 = sel_558633 + 8'h01;
  assign sel_558637 = array_index_558612 == array_index_537048 ? add_558636 : sel_558633;
  assign add_558640 = sel_558637 + 8'h01;
  assign sel_558641 = array_index_558612 == array_index_537056 ? add_558640 : sel_558637;
  assign add_558644 = sel_558641 + 8'h01;
  assign sel_558645 = array_index_558612 == array_index_537064 ? add_558644 : sel_558641;
  assign add_558648 = sel_558645 + 8'h01;
  assign sel_558649 = array_index_558612 == array_index_537070 ? add_558648 : sel_558645;
  assign add_558652 = sel_558649 + 8'h01;
  assign sel_558653 = array_index_558612 == array_index_537076 ? add_558652 : sel_558649;
  assign add_558656 = sel_558653 + 8'h01;
  assign sel_558657 = array_index_558612 == array_index_537082 ? add_558656 : sel_558653;
  assign add_558660 = sel_558657 + 8'h01;
  assign sel_558661 = array_index_558612 == array_index_537088 ? add_558660 : sel_558657;
  assign add_558664 = sel_558661 + 8'h01;
  assign sel_558665 = array_index_558612 == array_index_537094 ? add_558664 : sel_558661;
  assign add_558668 = sel_558665 + 8'h01;
  assign sel_558669 = array_index_558612 == array_index_537100 ? add_558668 : sel_558665;
  assign add_558672 = sel_558669 + 8'h01;
  assign sel_558673 = array_index_558612 == array_index_537106 ? add_558672 : sel_558669;
  assign add_558676 = sel_558673 + 8'h01;
  assign sel_558677 = array_index_558612 == array_index_537112 ? add_558676 : sel_558673;
  assign add_558680 = sel_558677 + 8'h01;
  assign sel_558681 = array_index_558612 == array_index_537118 ? add_558680 : sel_558677;
  assign add_558684 = sel_558681 + 8'h01;
  assign sel_558685 = array_index_558612 == array_index_537124 ? add_558684 : sel_558681;
  assign add_558688 = sel_558685 + 8'h01;
  assign sel_558689 = array_index_558612 == array_index_537130 ? add_558688 : sel_558685;
  assign add_558692 = sel_558689 + 8'h01;
  assign sel_558693 = array_index_558612 == array_index_537136 ? add_558692 : sel_558689;
  assign add_558696 = sel_558693 + 8'h01;
  assign sel_558697 = array_index_558612 == array_index_537142 ? add_558696 : sel_558693;
  assign add_558700 = sel_558697 + 8'h01;
  assign sel_558701 = array_index_558612 == array_index_537148 ? add_558700 : sel_558697;
  assign add_558704 = sel_558701 + 8'h01;
  assign sel_558705 = array_index_558612 == array_index_537154 ? add_558704 : sel_558701;
  assign add_558708 = sel_558705 + 8'h01;
  assign sel_558709 = array_index_558612 == array_index_537160 ? add_558708 : sel_558705;
  assign add_558712 = sel_558709 + 8'h01;
  assign sel_558713 = array_index_558612 == array_index_537166 ? add_558712 : sel_558709;
  assign add_558716 = sel_558713 + 8'h01;
  assign sel_558717 = array_index_558612 == array_index_537172 ? add_558716 : sel_558713;
  assign add_558720 = sel_558717 + 8'h01;
  assign sel_558721 = array_index_558612 == array_index_537178 ? add_558720 : sel_558717;
  assign add_558724 = sel_558721 + 8'h01;
  assign sel_558725 = array_index_558612 == array_index_537184 ? add_558724 : sel_558721;
  assign add_558728 = sel_558725 + 8'h01;
  assign sel_558729 = array_index_558612 == array_index_537190 ? add_558728 : sel_558725;
  assign add_558732 = sel_558729 + 8'h01;
  assign sel_558733 = array_index_558612 == array_index_537196 ? add_558732 : sel_558729;
  assign add_558736 = sel_558733 + 8'h01;
  assign sel_558737 = array_index_558612 == array_index_537202 ? add_558736 : sel_558733;
  assign add_558740 = sel_558737 + 8'h01;
  assign sel_558741 = array_index_558612 == array_index_537208 ? add_558740 : sel_558737;
  assign add_558744 = sel_558741 + 8'h01;
  assign sel_558745 = array_index_558612 == array_index_537214 ? add_558744 : sel_558741;
  assign add_558748 = sel_558745 + 8'h01;
  assign sel_558749 = array_index_558612 == array_index_537220 ? add_558748 : sel_558745;
  assign add_558752 = sel_558749 + 8'h01;
  assign sel_558753 = array_index_558612 == array_index_537226 ? add_558752 : sel_558749;
  assign add_558756 = sel_558753 + 8'h01;
  assign sel_558757 = array_index_558612 == array_index_537232 ? add_558756 : sel_558753;
  assign add_558760 = sel_558757 + 8'h01;
  assign sel_558761 = array_index_558612 == array_index_537238 ? add_558760 : sel_558757;
  assign add_558764 = sel_558761 + 8'h01;
  assign sel_558765 = array_index_558612 == array_index_537244 ? add_558764 : sel_558761;
  assign add_558768 = sel_558765 + 8'h01;
  assign sel_558769 = array_index_558612 == array_index_537250 ? add_558768 : sel_558765;
  assign add_558772 = sel_558769 + 8'h01;
  assign sel_558773 = array_index_558612 == array_index_537256 ? add_558772 : sel_558769;
  assign add_558776 = sel_558773 + 8'h01;
  assign sel_558777 = array_index_558612 == array_index_537262 ? add_558776 : sel_558773;
  assign add_558780 = sel_558777 + 8'h01;
  assign sel_558781 = array_index_558612 == array_index_537268 ? add_558780 : sel_558777;
  assign add_558784 = sel_558781 + 8'h01;
  assign sel_558785 = array_index_558612 == array_index_537274 ? add_558784 : sel_558781;
  assign add_558788 = sel_558785 + 8'h01;
  assign sel_558789 = array_index_558612 == array_index_537280 ? add_558788 : sel_558785;
  assign add_558792 = sel_558789 + 8'h01;
  assign sel_558793 = array_index_558612 == array_index_537286 ? add_558792 : sel_558789;
  assign add_558796 = sel_558793 + 8'h01;
  assign sel_558797 = array_index_558612 == array_index_537292 ? add_558796 : sel_558793;
  assign add_558800 = sel_558797 + 8'h01;
  assign sel_558801 = array_index_558612 == array_index_537298 ? add_558800 : sel_558797;
  assign add_558804 = sel_558801 + 8'h01;
  assign sel_558805 = array_index_558612 == array_index_537304 ? add_558804 : sel_558801;
  assign add_558808 = sel_558805 + 8'h01;
  assign sel_558809 = array_index_558612 == array_index_537310 ? add_558808 : sel_558805;
  assign add_558812 = sel_558809 + 8'h01;
  assign sel_558813 = array_index_558612 == array_index_537316 ? add_558812 : sel_558809;
  assign add_558816 = sel_558813 + 8'h01;
  assign sel_558817 = array_index_558612 == array_index_537322 ? add_558816 : sel_558813;
  assign add_558820 = sel_558817 + 8'h01;
  assign sel_558821 = array_index_558612 == array_index_537328 ? add_558820 : sel_558817;
  assign add_558824 = sel_558821 + 8'h01;
  assign sel_558825 = array_index_558612 == array_index_537334 ? add_558824 : sel_558821;
  assign add_558828 = sel_558825 + 8'h01;
  assign sel_558829 = array_index_558612 == array_index_537340 ? add_558828 : sel_558825;
  assign add_558832 = sel_558829 + 8'h01;
  assign sel_558833 = array_index_558612 == array_index_537346 ? add_558832 : sel_558829;
  assign add_558836 = sel_558833 + 8'h01;
  assign sel_558837 = array_index_558612 == array_index_537352 ? add_558836 : sel_558833;
  assign add_558840 = sel_558837 + 8'h01;
  assign sel_558841 = array_index_558612 == array_index_537358 ? add_558840 : sel_558837;
  assign add_558844 = sel_558841 + 8'h01;
  assign sel_558845 = array_index_558612 == array_index_537364 ? add_558844 : sel_558841;
  assign add_558848 = sel_558845 + 8'h01;
  assign sel_558849 = array_index_558612 == array_index_537370 ? add_558848 : sel_558845;
  assign add_558852 = sel_558849 + 8'h01;
  assign sel_558853 = array_index_558612 == array_index_537376 ? add_558852 : sel_558849;
  assign add_558856 = sel_558853 + 8'h01;
  assign sel_558857 = array_index_558612 == array_index_537382 ? add_558856 : sel_558853;
  assign add_558860 = sel_558857 + 8'h01;
  assign sel_558861 = array_index_558612 == array_index_537388 ? add_558860 : sel_558857;
  assign add_558864 = sel_558861 + 8'h01;
  assign sel_558865 = array_index_558612 == array_index_537394 ? add_558864 : sel_558861;
  assign add_558868 = sel_558865 + 8'h01;
  assign sel_558869 = array_index_558612 == array_index_537400 ? add_558868 : sel_558865;
  assign add_558872 = sel_558869 + 8'h01;
  assign sel_558873 = array_index_558612 == array_index_537406 ? add_558872 : sel_558869;
  assign add_558876 = sel_558873 + 8'h01;
  assign sel_558877 = array_index_558612 == array_index_537412 ? add_558876 : sel_558873;
  assign add_558880 = sel_558877 + 8'h01;
  assign sel_558881 = array_index_558612 == array_index_537418 ? add_558880 : sel_558877;
  assign add_558884 = sel_558881 + 8'h01;
  assign sel_558885 = array_index_558612 == array_index_537424 ? add_558884 : sel_558881;
  assign add_558888 = sel_558885 + 8'h01;
  assign sel_558889 = array_index_558612 == array_index_537430 ? add_558888 : sel_558885;
  assign add_558892 = sel_558889 + 8'h01;
  assign sel_558893 = array_index_558612 == array_index_537436 ? add_558892 : sel_558889;
  assign add_558896 = sel_558893 + 8'h01;
  assign sel_558897 = array_index_558612 == array_index_537442 ? add_558896 : sel_558893;
  assign add_558900 = sel_558897 + 8'h01;
  assign sel_558901 = array_index_558612 == array_index_537448 ? add_558900 : sel_558897;
  assign add_558904 = sel_558901 + 8'h01;
  assign sel_558905 = array_index_558612 == array_index_537454 ? add_558904 : sel_558901;
  assign add_558908 = sel_558905 + 8'h01;
  assign sel_558909 = array_index_558612 == array_index_537460 ? add_558908 : sel_558905;
  assign add_558913 = sel_558909 + 8'h01;
  assign array_index_558914 = set1_unflattened[7'h48];
  assign sel_558915 = array_index_558612 == array_index_537466 ? add_558913 : sel_558909;
  assign add_558918 = sel_558915 + 8'h01;
  assign sel_558919 = array_index_558914 == array_index_537012 ? add_558918 : sel_558915;
  assign add_558922 = sel_558919 + 8'h01;
  assign sel_558923 = array_index_558914 == array_index_537016 ? add_558922 : sel_558919;
  assign add_558926 = sel_558923 + 8'h01;
  assign sel_558927 = array_index_558914 == array_index_537024 ? add_558926 : sel_558923;
  assign add_558930 = sel_558927 + 8'h01;
  assign sel_558931 = array_index_558914 == array_index_537032 ? add_558930 : sel_558927;
  assign add_558934 = sel_558931 + 8'h01;
  assign sel_558935 = array_index_558914 == array_index_537040 ? add_558934 : sel_558931;
  assign add_558938 = sel_558935 + 8'h01;
  assign sel_558939 = array_index_558914 == array_index_537048 ? add_558938 : sel_558935;
  assign add_558942 = sel_558939 + 8'h01;
  assign sel_558943 = array_index_558914 == array_index_537056 ? add_558942 : sel_558939;
  assign add_558946 = sel_558943 + 8'h01;
  assign sel_558947 = array_index_558914 == array_index_537064 ? add_558946 : sel_558943;
  assign add_558950 = sel_558947 + 8'h01;
  assign sel_558951 = array_index_558914 == array_index_537070 ? add_558950 : sel_558947;
  assign add_558954 = sel_558951 + 8'h01;
  assign sel_558955 = array_index_558914 == array_index_537076 ? add_558954 : sel_558951;
  assign add_558958 = sel_558955 + 8'h01;
  assign sel_558959 = array_index_558914 == array_index_537082 ? add_558958 : sel_558955;
  assign add_558962 = sel_558959 + 8'h01;
  assign sel_558963 = array_index_558914 == array_index_537088 ? add_558962 : sel_558959;
  assign add_558966 = sel_558963 + 8'h01;
  assign sel_558967 = array_index_558914 == array_index_537094 ? add_558966 : sel_558963;
  assign add_558970 = sel_558967 + 8'h01;
  assign sel_558971 = array_index_558914 == array_index_537100 ? add_558970 : sel_558967;
  assign add_558974 = sel_558971 + 8'h01;
  assign sel_558975 = array_index_558914 == array_index_537106 ? add_558974 : sel_558971;
  assign add_558978 = sel_558975 + 8'h01;
  assign sel_558979 = array_index_558914 == array_index_537112 ? add_558978 : sel_558975;
  assign add_558982 = sel_558979 + 8'h01;
  assign sel_558983 = array_index_558914 == array_index_537118 ? add_558982 : sel_558979;
  assign add_558986 = sel_558983 + 8'h01;
  assign sel_558987 = array_index_558914 == array_index_537124 ? add_558986 : sel_558983;
  assign add_558990 = sel_558987 + 8'h01;
  assign sel_558991 = array_index_558914 == array_index_537130 ? add_558990 : sel_558987;
  assign add_558994 = sel_558991 + 8'h01;
  assign sel_558995 = array_index_558914 == array_index_537136 ? add_558994 : sel_558991;
  assign add_558998 = sel_558995 + 8'h01;
  assign sel_558999 = array_index_558914 == array_index_537142 ? add_558998 : sel_558995;
  assign add_559002 = sel_558999 + 8'h01;
  assign sel_559003 = array_index_558914 == array_index_537148 ? add_559002 : sel_558999;
  assign add_559006 = sel_559003 + 8'h01;
  assign sel_559007 = array_index_558914 == array_index_537154 ? add_559006 : sel_559003;
  assign add_559010 = sel_559007 + 8'h01;
  assign sel_559011 = array_index_558914 == array_index_537160 ? add_559010 : sel_559007;
  assign add_559014 = sel_559011 + 8'h01;
  assign sel_559015 = array_index_558914 == array_index_537166 ? add_559014 : sel_559011;
  assign add_559018 = sel_559015 + 8'h01;
  assign sel_559019 = array_index_558914 == array_index_537172 ? add_559018 : sel_559015;
  assign add_559022 = sel_559019 + 8'h01;
  assign sel_559023 = array_index_558914 == array_index_537178 ? add_559022 : sel_559019;
  assign add_559026 = sel_559023 + 8'h01;
  assign sel_559027 = array_index_558914 == array_index_537184 ? add_559026 : sel_559023;
  assign add_559030 = sel_559027 + 8'h01;
  assign sel_559031 = array_index_558914 == array_index_537190 ? add_559030 : sel_559027;
  assign add_559034 = sel_559031 + 8'h01;
  assign sel_559035 = array_index_558914 == array_index_537196 ? add_559034 : sel_559031;
  assign add_559038 = sel_559035 + 8'h01;
  assign sel_559039 = array_index_558914 == array_index_537202 ? add_559038 : sel_559035;
  assign add_559042 = sel_559039 + 8'h01;
  assign sel_559043 = array_index_558914 == array_index_537208 ? add_559042 : sel_559039;
  assign add_559046 = sel_559043 + 8'h01;
  assign sel_559047 = array_index_558914 == array_index_537214 ? add_559046 : sel_559043;
  assign add_559050 = sel_559047 + 8'h01;
  assign sel_559051 = array_index_558914 == array_index_537220 ? add_559050 : sel_559047;
  assign add_559054 = sel_559051 + 8'h01;
  assign sel_559055 = array_index_558914 == array_index_537226 ? add_559054 : sel_559051;
  assign add_559058 = sel_559055 + 8'h01;
  assign sel_559059 = array_index_558914 == array_index_537232 ? add_559058 : sel_559055;
  assign add_559062 = sel_559059 + 8'h01;
  assign sel_559063 = array_index_558914 == array_index_537238 ? add_559062 : sel_559059;
  assign add_559066 = sel_559063 + 8'h01;
  assign sel_559067 = array_index_558914 == array_index_537244 ? add_559066 : sel_559063;
  assign add_559070 = sel_559067 + 8'h01;
  assign sel_559071 = array_index_558914 == array_index_537250 ? add_559070 : sel_559067;
  assign add_559074 = sel_559071 + 8'h01;
  assign sel_559075 = array_index_558914 == array_index_537256 ? add_559074 : sel_559071;
  assign add_559078 = sel_559075 + 8'h01;
  assign sel_559079 = array_index_558914 == array_index_537262 ? add_559078 : sel_559075;
  assign add_559082 = sel_559079 + 8'h01;
  assign sel_559083 = array_index_558914 == array_index_537268 ? add_559082 : sel_559079;
  assign add_559086 = sel_559083 + 8'h01;
  assign sel_559087 = array_index_558914 == array_index_537274 ? add_559086 : sel_559083;
  assign add_559090 = sel_559087 + 8'h01;
  assign sel_559091 = array_index_558914 == array_index_537280 ? add_559090 : sel_559087;
  assign add_559094 = sel_559091 + 8'h01;
  assign sel_559095 = array_index_558914 == array_index_537286 ? add_559094 : sel_559091;
  assign add_559098 = sel_559095 + 8'h01;
  assign sel_559099 = array_index_558914 == array_index_537292 ? add_559098 : sel_559095;
  assign add_559102 = sel_559099 + 8'h01;
  assign sel_559103 = array_index_558914 == array_index_537298 ? add_559102 : sel_559099;
  assign add_559106 = sel_559103 + 8'h01;
  assign sel_559107 = array_index_558914 == array_index_537304 ? add_559106 : sel_559103;
  assign add_559110 = sel_559107 + 8'h01;
  assign sel_559111 = array_index_558914 == array_index_537310 ? add_559110 : sel_559107;
  assign add_559114 = sel_559111 + 8'h01;
  assign sel_559115 = array_index_558914 == array_index_537316 ? add_559114 : sel_559111;
  assign add_559118 = sel_559115 + 8'h01;
  assign sel_559119 = array_index_558914 == array_index_537322 ? add_559118 : sel_559115;
  assign add_559122 = sel_559119 + 8'h01;
  assign sel_559123 = array_index_558914 == array_index_537328 ? add_559122 : sel_559119;
  assign add_559126 = sel_559123 + 8'h01;
  assign sel_559127 = array_index_558914 == array_index_537334 ? add_559126 : sel_559123;
  assign add_559130 = sel_559127 + 8'h01;
  assign sel_559131 = array_index_558914 == array_index_537340 ? add_559130 : sel_559127;
  assign add_559134 = sel_559131 + 8'h01;
  assign sel_559135 = array_index_558914 == array_index_537346 ? add_559134 : sel_559131;
  assign add_559138 = sel_559135 + 8'h01;
  assign sel_559139 = array_index_558914 == array_index_537352 ? add_559138 : sel_559135;
  assign add_559142 = sel_559139 + 8'h01;
  assign sel_559143 = array_index_558914 == array_index_537358 ? add_559142 : sel_559139;
  assign add_559146 = sel_559143 + 8'h01;
  assign sel_559147 = array_index_558914 == array_index_537364 ? add_559146 : sel_559143;
  assign add_559150 = sel_559147 + 8'h01;
  assign sel_559151 = array_index_558914 == array_index_537370 ? add_559150 : sel_559147;
  assign add_559154 = sel_559151 + 8'h01;
  assign sel_559155 = array_index_558914 == array_index_537376 ? add_559154 : sel_559151;
  assign add_559158 = sel_559155 + 8'h01;
  assign sel_559159 = array_index_558914 == array_index_537382 ? add_559158 : sel_559155;
  assign add_559162 = sel_559159 + 8'h01;
  assign sel_559163 = array_index_558914 == array_index_537388 ? add_559162 : sel_559159;
  assign add_559166 = sel_559163 + 8'h01;
  assign sel_559167 = array_index_558914 == array_index_537394 ? add_559166 : sel_559163;
  assign add_559170 = sel_559167 + 8'h01;
  assign sel_559171 = array_index_558914 == array_index_537400 ? add_559170 : sel_559167;
  assign add_559174 = sel_559171 + 8'h01;
  assign sel_559175 = array_index_558914 == array_index_537406 ? add_559174 : sel_559171;
  assign add_559178 = sel_559175 + 8'h01;
  assign sel_559179 = array_index_558914 == array_index_537412 ? add_559178 : sel_559175;
  assign add_559182 = sel_559179 + 8'h01;
  assign sel_559183 = array_index_558914 == array_index_537418 ? add_559182 : sel_559179;
  assign add_559186 = sel_559183 + 8'h01;
  assign sel_559187 = array_index_558914 == array_index_537424 ? add_559186 : sel_559183;
  assign add_559190 = sel_559187 + 8'h01;
  assign sel_559191 = array_index_558914 == array_index_537430 ? add_559190 : sel_559187;
  assign add_559194 = sel_559191 + 8'h01;
  assign sel_559195 = array_index_558914 == array_index_537436 ? add_559194 : sel_559191;
  assign add_559198 = sel_559195 + 8'h01;
  assign sel_559199 = array_index_558914 == array_index_537442 ? add_559198 : sel_559195;
  assign add_559202 = sel_559199 + 8'h01;
  assign sel_559203 = array_index_558914 == array_index_537448 ? add_559202 : sel_559199;
  assign add_559206 = sel_559203 + 8'h01;
  assign sel_559207 = array_index_558914 == array_index_537454 ? add_559206 : sel_559203;
  assign add_559210 = sel_559207 + 8'h01;
  assign sel_559211 = array_index_558914 == array_index_537460 ? add_559210 : sel_559207;
  assign add_559215 = sel_559211 + 8'h01;
  assign array_index_559216 = set1_unflattened[7'h49];
  assign sel_559217 = array_index_558914 == array_index_537466 ? add_559215 : sel_559211;
  assign add_559220 = sel_559217 + 8'h01;
  assign sel_559221 = array_index_559216 == array_index_537012 ? add_559220 : sel_559217;
  assign add_559224 = sel_559221 + 8'h01;
  assign sel_559225 = array_index_559216 == array_index_537016 ? add_559224 : sel_559221;
  assign add_559228 = sel_559225 + 8'h01;
  assign sel_559229 = array_index_559216 == array_index_537024 ? add_559228 : sel_559225;
  assign add_559232 = sel_559229 + 8'h01;
  assign sel_559233 = array_index_559216 == array_index_537032 ? add_559232 : sel_559229;
  assign add_559236 = sel_559233 + 8'h01;
  assign sel_559237 = array_index_559216 == array_index_537040 ? add_559236 : sel_559233;
  assign add_559240 = sel_559237 + 8'h01;
  assign sel_559241 = array_index_559216 == array_index_537048 ? add_559240 : sel_559237;
  assign add_559244 = sel_559241 + 8'h01;
  assign sel_559245 = array_index_559216 == array_index_537056 ? add_559244 : sel_559241;
  assign add_559248 = sel_559245 + 8'h01;
  assign sel_559249 = array_index_559216 == array_index_537064 ? add_559248 : sel_559245;
  assign add_559252 = sel_559249 + 8'h01;
  assign sel_559253 = array_index_559216 == array_index_537070 ? add_559252 : sel_559249;
  assign add_559256 = sel_559253 + 8'h01;
  assign sel_559257 = array_index_559216 == array_index_537076 ? add_559256 : sel_559253;
  assign add_559260 = sel_559257 + 8'h01;
  assign sel_559261 = array_index_559216 == array_index_537082 ? add_559260 : sel_559257;
  assign add_559264 = sel_559261 + 8'h01;
  assign sel_559265 = array_index_559216 == array_index_537088 ? add_559264 : sel_559261;
  assign add_559268 = sel_559265 + 8'h01;
  assign sel_559269 = array_index_559216 == array_index_537094 ? add_559268 : sel_559265;
  assign add_559272 = sel_559269 + 8'h01;
  assign sel_559273 = array_index_559216 == array_index_537100 ? add_559272 : sel_559269;
  assign add_559276 = sel_559273 + 8'h01;
  assign sel_559277 = array_index_559216 == array_index_537106 ? add_559276 : sel_559273;
  assign add_559280 = sel_559277 + 8'h01;
  assign sel_559281 = array_index_559216 == array_index_537112 ? add_559280 : sel_559277;
  assign add_559284 = sel_559281 + 8'h01;
  assign sel_559285 = array_index_559216 == array_index_537118 ? add_559284 : sel_559281;
  assign add_559288 = sel_559285 + 8'h01;
  assign sel_559289 = array_index_559216 == array_index_537124 ? add_559288 : sel_559285;
  assign add_559292 = sel_559289 + 8'h01;
  assign sel_559293 = array_index_559216 == array_index_537130 ? add_559292 : sel_559289;
  assign add_559296 = sel_559293 + 8'h01;
  assign sel_559297 = array_index_559216 == array_index_537136 ? add_559296 : sel_559293;
  assign add_559300 = sel_559297 + 8'h01;
  assign sel_559301 = array_index_559216 == array_index_537142 ? add_559300 : sel_559297;
  assign add_559304 = sel_559301 + 8'h01;
  assign sel_559305 = array_index_559216 == array_index_537148 ? add_559304 : sel_559301;
  assign add_559308 = sel_559305 + 8'h01;
  assign sel_559309 = array_index_559216 == array_index_537154 ? add_559308 : sel_559305;
  assign add_559312 = sel_559309 + 8'h01;
  assign sel_559313 = array_index_559216 == array_index_537160 ? add_559312 : sel_559309;
  assign add_559316 = sel_559313 + 8'h01;
  assign sel_559317 = array_index_559216 == array_index_537166 ? add_559316 : sel_559313;
  assign add_559320 = sel_559317 + 8'h01;
  assign sel_559321 = array_index_559216 == array_index_537172 ? add_559320 : sel_559317;
  assign add_559324 = sel_559321 + 8'h01;
  assign sel_559325 = array_index_559216 == array_index_537178 ? add_559324 : sel_559321;
  assign add_559328 = sel_559325 + 8'h01;
  assign sel_559329 = array_index_559216 == array_index_537184 ? add_559328 : sel_559325;
  assign add_559332 = sel_559329 + 8'h01;
  assign sel_559333 = array_index_559216 == array_index_537190 ? add_559332 : sel_559329;
  assign add_559336 = sel_559333 + 8'h01;
  assign sel_559337 = array_index_559216 == array_index_537196 ? add_559336 : sel_559333;
  assign add_559340 = sel_559337 + 8'h01;
  assign sel_559341 = array_index_559216 == array_index_537202 ? add_559340 : sel_559337;
  assign add_559344 = sel_559341 + 8'h01;
  assign sel_559345 = array_index_559216 == array_index_537208 ? add_559344 : sel_559341;
  assign add_559348 = sel_559345 + 8'h01;
  assign sel_559349 = array_index_559216 == array_index_537214 ? add_559348 : sel_559345;
  assign add_559352 = sel_559349 + 8'h01;
  assign sel_559353 = array_index_559216 == array_index_537220 ? add_559352 : sel_559349;
  assign add_559356 = sel_559353 + 8'h01;
  assign sel_559357 = array_index_559216 == array_index_537226 ? add_559356 : sel_559353;
  assign add_559360 = sel_559357 + 8'h01;
  assign sel_559361 = array_index_559216 == array_index_537232 ? add_559360 : sel_559357;
  assign add_559364 = sel_559361 + 8'h01;
  assign sel_559365 = array_index_559216 == array_index_537238 ? add_559364 : sel_559361;
  assign add_559368 = sel_559365 + 8'h01;
  assign sel_559369 = array_index_559216 == array_index_537244 ? add_559368 : sel_559365;
  assign add_559372 = sel_559369 + 8'h01;
  assign sel_559373 = array_index_559216 == array_index_537250 ? add_559372 : sel_559369;
  assign add_559376 = sel_559373 + 8'h01;
  assign sel_559377 = array_index_559216 == array_index_537256 ? add_559376 : sel_559373;
  assign add_559380 = sel_559377 + 8'h01;
  assign sel_559381 = array_index_559216 == array_index_537262 ? add_559380 : sel_559377;
  assign add_559384 = sel_559381 + 8'h01;
  assign sel_559385 = array_index_559216 == array_index_537268 ? add_559384 : sel_559381;
  assign add_559388 = sel_559385 + 8'h01;
  assign sel_559389 = array_index_559216 == array_index_537274 ? add_559388 : sel_559385;
  assign add_559392 = sel_559389 + 8'h01;
  assign sel_559393 = array_index_559216 == array_index_537280 ? add_559392 : sel_559389;
  assign add_559396 = sel_559393 + 8'h01;
  assign sel_559397 = array_index_559216 == array_index_537286 ? add_559396 : sel_559393;
  assign add_559400 = sel_559397 + 8'h01;
  assign sel_559401 = array_index_559216 == array_index_537292 ? add_559400 : sel_559397;
  assign add_559404 = sel_559401 + 8'h01;
  assign sel_559405 = array_index_559216 == array_index_537298 ? add_559404 : sel_559401;
  assign add_559408 = sel_559405 + 8'h01;
  assign sel_559409 = array_index_559216 == array_index_537304 ? add_559408 : sel_559405;
  assign add_559412 = sel_559409 + 8'h01;
  assign sel_559413 = array_index_559216 == array_index_537310 ? add_559412 : sel_559409;
  assign add_559416 = sel_559413 + 8'h01;
  assign sel_559417 = array_index_559216 == array_index_537316 ? add_559416 : sel_559413;
  assign add_559420 = sel_559417 + 8'h01;
  assign sel_559421 = array_index_559216 == array_index_537322 ? add_559420 : sel_559417;
  assign add_559424 = sel_559421 + 8'h01;
  assign sel_559425 = array_index_559216 == array_index_537328 ? add_559424 : sel_559421;
  assign add_559428 = sel_559425 + 8'h01;
  assign sel_559429 = array_index_559216 == array_index_537334 ? add_559428 : sel_559425;
  assign add_559432 = sel_559429 + 8'h01;
  assign sel_559433 = array_index_559216 == array_index_537340 ? add_559432 : sel_559429;
  assign add_559436 = sel_559433 + 8'h01;
  assign sel_559437 = array_index_559216 == array_index_537346 ? add_559436 : sel_559433;
  assign add_559440 = sel_559437 + 8'h01;
  assign sel_559441 = array_index_559216 == array_index_537352 ? add_559440 : sel_559437;
  assign add_559444 = sel_559441 + 8'h01;
  assign sel_559445 = array_index_559216 == array_index_537358 ? add_559444 : sel_559441;
  assign add_559448 = sel_559445 + 8'h01;
  assign sel_559449 = array_index_559216 == array_index_537364 ? add_559448 : sel_559445;
  assign add_559452 = sel_559449 + 8'h01;
  assign sel_559453 = array_index_559216 == array_index_537370 ? add_559452 : sel_559449;
  assign add_559456 = sel_559453 + 8'h01;
  assign sel_559457 = array_index_559216 == array_index_537376 ? add_559456 : sel_559453;
  assign add_559460 = sel_559457 + 8'h01;
  assign sel_559461 = array_index_559216 == array_index_537382 ? add_559460 : sel_559457;
  assign add_559464 = sel_559461 + 8'h01;
  assign sel_559465 = array_index_559216 == array_index_537388 ? add_559464 : sel_559461;
  assign add_559468 = sel_559465 + 8'h01;
  assign sel_559469 = array_index_559216 == array_index_537394 ? add_559468 : sel_559465;
  assign add_559472 = sel_559469 + 8'h01;
  assign sel_559473 = array_index_559216 == array_index_537400 ? add_559472 : sel_559469;
  assign add_559476 = sel_559473 + 8'h01;
  assign sel_559477 = array_index_559216 == array_index_537406 ? add_559476 : sel_559473;
  assign add_559480 = sel_559477 + 8'h01;
  assign sel_559481 = array_index_559216 == array_index_537412 ? add_559480 : sel_559477;
  assign add_559484 = sel_559481 + 8'h01;
  assign sel_559485 = array_index_559216 == array_index_537418 ? add_559484 : sel_559481;
  assign add_559488 = sel_559485 + 8'h01;
  assign sel_559489 = array_index_559216 == array_index_537424 ? add_559488 : sel_559485;
  assign add_559492 = sel_559489 + 8'h01;
  assign sel_559493 = array_index_559216 == array_index_537430 ? add_559492 : sel_559489;
  assign add_559496 = sel_559493 + 8'h01;
  assign sel_559497 = array_index_559216 == array_index_537436 ? add_559496 : sel_559493;
  assign add_559500 = sel_559497 + 8'h01;
  assign sel_559501 = array_index_559216 == array_index_537442 ? add_559500 : sel_559497;
  assign add_559504 = sel_559501 + 8'h01;
  assign sel_559505 = array_index_559216 == array_index_537448 ? add_559504 : sel_559501;
  assign add_559508 = sel_559505 + 8'h01;
  assign sel_559509 = array_index_559216 == array_index_537454 ? add_559508 : sel_559505;
  assign add_559512 = sel_559509 + 8'h01;
  assign sel_559513 = array_index_559216 == array_index_537460 ? add_559512 : sel_559509;
  assign add_559517 = sel_559513 + 8'h01;
  assign array_index_559518 = set1_unflattened[7'h4a];
  assign sel_559519 = array_index_559216 == array_index_537466 ? add_559517 : sel_559513;
  assign add_559522 = sel_559519 + 8'h01;
  assign sel_559523 = array_index_559518 == array_index_537012 ? add_559522 : sel_559519;
  assign add_559526 = sel_559523 + 8'h01;
  assign sel_559527 = array_index_559518 == array_index_537016 ? add_559526 : sel_559523;
  assign add_559530 = sel_559527 + 8'h01;
  assign sel_559531 = array_index_559518 == array_index_537024 ? add_559530 : sel_559527;
  assign add_559534 = sel_559531 + 8'h01;
  assign sel_559535 = array_index_559518 == array_index_537032 ? add_559534 : sel_559531;
  assign add_559538 = sel_559535 + 8'h01;
  assign sel_559539 = array_index_559518 == array_index_537040 ? add_559538 : sel_559535;
  assign add_559542 = sel_559539 + 8'h01;
  assign sel_559543 = array_index_559518 == array_index_537048 ? add_559542 : sel_559539;
  assign add_559546 = sel_559543 + 8'h01;
  assign sel_559547 = array_index_559518 == array_index_537056 ? add_559546 : sel_559543;
  assign add_559550 = sel_559547 + 8'h01;
  assign sel_559551 = array_index_559518 == array_index_537064 ? add_559550 : sel_559547;
  assign add_559554 = sel_559551 + 8'h01;
  assign sel_559555 = array_index_559518 == array_index_537070 ? add_559554 : sel_559551;
  assign add_559558 = sel_559555 + 8'h01;
  assign sel_559559 = array_index_559518 == array_index_537076 ? add_559558 : sel_559555;
  assign add_559562 = sel_559559 + 8'h01;
  assign sel_559563 = array_index_559518 == array_index_537082 ? add_559562 : sel_559559;
  assign add_559566 = sel_559563 + 8'h01;
  assign sel_559567 = array_index_559518 == array_index_537088 ? add_559566 : sel_559563;
  assign add_559570 = sel_559567 + 8'h01;
  assign sel_559571 = array_index_559518 == array_index_537094 ? add_559570 : sel_559567;
  assign add_559574 = sel_559571 + 8'h01;
  assign sel_559575 = array_index_559518 == array_index_537100 ? add_559574 : sel_559571;
  assign add_559578 = sel_559575 + 8'h01;
  assign sel_559579 = array_index_559518 == array_index_537106 ? add_559578 : sel_559575;
  assign add_559582 = sel_559579 + 8'h01;
  assign sel_559583 = array_index_559518 == array_index_537112 ? add_559582 : sel_559579;
  assign add_559586 = sel_559583 + 8'h01;
  assign sel_559587 = array_index_559518 == array_index_537118 ? add_559586 : sel_559583;
  assign add_559590 = sel_559587 + 8'h01;
  assign sel_559591 = array_index_559518 == array_index_537124 ? add_559590 : sel_559587;
  assign add_559594 = sel_559591 + 8'h01;
  assign sel_559595 = array_index_559518 == array_index_537130 ? add_559594 : sel_559591;
  assign add_559598 = sel_559595 + 8'h01;
  assign sel_559599 = array_index_559518 == array_index_537136 ? add_559598 : sel_559595;
  assign add_559602 = sel_559599 + 8'h01;
  assign sel_559603 = array_index_559518 == array_index_537142 ? add_559602 : sel_559599;
  assign add_559606 = sel_559603 + 8'h01;
  assign sel_559607 = array_index_559518 == array_index_537148 ? add_559606 : sel_559603;
  assign add_559610 = sel_559607 + 8'h01;
  assign sel_559611 = array_index_559518 == array_index_537154 ? add_559610 : sel_559607;
  assign add_559614 = sel_559611 + 8'h01;
  assign sel_559615 = array_index_559518 == array_index_537160 ? add_559614 : sel_559611;
  assign add_559618 = sel_559615 + 8'h01;
  assign sel_559619 = array_index_559518 == array_index_537166 ? add_559618 : sel_559615;
  assign add_559622 = sel_559619 + 8'h01;
  assign sel_559623 = array_index_559518 == array_index_537172 ? add_559622 : sel_559619;
  assign add_559626 = sel_559623 + 8'h01;
  assign sel_559627 = array_index_559518 == array_index_537178 ? add_559626 : sel_559623;
  assign add_559630 = sel_559627 + 8'h01;
  assign sel_559631 = array_index_559518 == array_index_537184 ? add_559630 : sel_559627;
  assign add_559634 = sel_559631 + 8'h01;
  assign sel_559635 = array_index_559518 == array_index_537190 ? add_559634 : sel_559631;
  assign add_559638 = sel_559635 + 8'h01;
  assign sel_559639 = array_index_559518 == array_index_537196 ? add_559638 : sel_559635;
  assign add_559642 = sel_559639 + 8'h01;
  assign sel_559643 = array_index_559518 == array_index_537202 ? add_559642 : sel_559639;
  assign add_559646 = sel_559643 + 8'h01;
  assign sel_559647 = array_index_559518 == array_index_537208 ? add_559646 : sel_559643;
  assign add_559650 = sel_559647 + 8'h01;
  assign sel_559651 = array_index_559518 == array_index_537214 ? add_559650 : sel_559647;
  assign add_559654 = sel_559651 + 8'h01;
  assign sel_559655 = array_index_559518 == array_index_537220 ? add_559654 : sel_559651;
  assign add_559658 = sel_559655 + 8'h01;
  assign sel_559659 = array_index_559518 == array_index_537226 ? add_559658 : sel_559655;
  assign add_559662 = sel_559659 + 8'h01;
  assign sel_559663 = array_index_559518 == array_index_537232 ? add_559662 : sel_559659;
  assign add_559666 = sel_559663 + 8'h01;
  assign sel_559667 = array_index_559518 == array_index_537238 ? add_559666 : sel_559663;
  assign add_559670 = sel_559667 + 8'h01;
  assign sel_559671 = array_index_559518 == array_index_537244 ? add_559670 : sel_559667;
  assign add_559674 = sel_559671 + 8'h01;
  assign sel_559675 = array_index_559518 == array_index_537250 ? add_559674 : sel_559671;
  assign add_559678 = sel_559675 + 8'h01;
  assign sel_559679 = array_index_559518 == array_index_537256 ? add_559678 : sel_559675;
  assign add_559682 = sel_559679 + 8'h01;
  assign sel_559683 = array_index_559518 == array_index_537262 ? add_559682 : sel_559679;
  assign add_559686 = sel_559683 + 8'h01;
  assign sel_559687 = array_index_559518 == array_index_537268 ? add_559686 : sel_559683;
  assign add_559690 = sel_559687 + 8'h01;
  assign sel_559691 = array_index_559518 == array_index_537274 ? add_559690 : sel_559687;
  assign add_559694 = sel_559691 + 8'h01;
  assign sel_559695 = array_index_559518 == array_index_537280 ? add_559694 : sel_559691;
  assign add_559698 = sel_559695 + 8'h01;
  assign sel_559699 = array_index_559518 == array_index_537286 ? add_559698 : sel_559695;
  assign add_559702 = sel_559699 + 8'h01;
  assign sel_559703 = array_index_559518 == array_index_537292 ? add_559702 : sel_559699;
  assign add_559706 = sel_559703 + 8'h01;
  assign sel_559707 = array_index_559518 == array_index_537298 ? add_559706 : sel_559703;
  assign add_559710 = sel_559707 + 8'h01;
  assign sel_559711 = array_index_559518 == array_index_537304 ? add_559710 : sel_559707;
  assign add_559714 = sel_559711 + 8'h01;
  assign sel_559715 = array_index_559518 == array_index_537310 ? add_559714 : sel_559711;
  assign add_559718 = sel_559715 + 8'h01;
  assign sel_559719 = array_index_559518 == array_index_537316 ? add_559718 : sel_559715;
  assign add_559722 = sel_559719 + 8'h01;
  assign sel_559723 = array_index_559518 == array_index_537322 ? add_559722 : sel_559719;
  assign add_559726 = sel_559723 + 8'h01;
  assign sel_559727 = array_index_559518 == array_index_537328 ? add_559726 : sel_559723;
  assign add_559730 = sel_559727 + 8'h01;
  assign sel_559731 = array_index_559518 == array_index_537334 ? add_559730 : sel_559727;
  assign add_559734 = sel_559731 + 8'h01;
  assign sel_559735 = array_index_559518 == array_index_537340 ? add_559734 : sel_559731;
  assign add_559738 = sel_559735 + 8'h01;
  assign sel_559739 = array_index_559518 == array_index_537346 ? add_559738 : sel_559735;
  assign add_559742 = sel_559739 + 8'h01;
  assign sel_559743 = array_index_559518 == array_index_537352 ? add_559742 : sel_559739;
  assign add_559746 = sel_559743 + 8'h01;
  assign sel_559747 = array_index_559518 == array_index_537358 ? add_559746 : sel_559743;
  assign add_559750 = sel_559747 + 8'h01;
  assign sel_559751 = array_index_559518 == array_index_537364 ? add_559750 : sel_559747;
  assign add_559754 = sel_559751 + 8'h01;
  assign sel_559755 = array_index_559518 == array_index_537370 ? add_559754 : sel_559751;
  assign add_559758 = sel_559755 + 8'h01;
  assign sel_559759 = array_index_559518 == array_index_537376 ? add_559758 : sel_559755;
  assign add_559762 = sel_559759 + 8'h01;
  assign sel_559763 = array_index_559518 == array_index_537382 ? add_559762 : sel_559759;
  assign add_559766 = sel_559763 + 8'h01;
  assign sel_559767 = array_index_559518 == array_index_537388 ? add_559766 : sel_559763;
  assign add_559770 = sel_559767 + 8'h01;
  assign sel_559771 = array_index_559518 == array_index_537394 ? add_559770 : sel_559767;
  assign add_559774 = sel_559771 + 8'h01;
  assign sel_559775 = array_index_559518 == array_index_537400 ? add_559774 : sel_559771;
  assign add_559778 = sel_559775 + 8'h01;
  assign sel_559779 = array_index_559518 == array_index_537406 ? add_559778 : sel_559775;
  assign add_559782 = sel_559779 + 8'h01;
  assign sel_559783 = array_index_559518 == array_index_537412 ? add_559782 : sel_559779;
  assign add_559786 = sel_559783 + 8'h01;
  assign sel_559787 = array_index_559518 == array_index_537418 ? add_559786 : sel_559783;
  assign add_559790 = sel_559787 + 8'h01;
  assign sel_559791 = array_index_559518 == array_index_537424 ? add_559790 : sel_559787;
  assign add_559794 = sel_559791 + 8'h01;
  assign sel_559795 = array_index_559518 == array_index_537430 ? add_559794 : sel_559791;
  assign add_559798 = sel_559795 + 8'h01;
  assign sel_559799 = array_index_559518 == array_index_537436 ? add_559798 : sel_559795;
  assign add_559802 = sel_559799 + 8'h01;
  assign sel_559803 = array_index_559518 == array_index_537442 ? add_559802 : sel_559799;
  assign add_559806 = sel_559803 + 8'h01;
  assign sel_559807 = array_index_559518 == array_index_537448 ? add_559806 : sel_559803;
  assign add_559810 = sel_559807 + 8'h01;
  assign sel_559811 = array_index_559518 == array_index_537454 ? add_559810 : sel_559807;
  assign add_559814 = sel_559811 + 8'h01;
  assign sel_559815 = array_index_559518 == array_index_537460 ? add_559814 : sel_559811;
  assign add_559818 = sel_559815 + 8'h01;
  assign out = {array_index_559518 == array_index_537466 ? add_559818 : sel_559815, {set1_unflattened[74], set1_unflattened[73], set1_unflattened[72], set1_unflattened[71], set1_unflattened[70], set1_unflattened[69], set1_unflattened[68], set1_unflattened[67], set1_unflattened[66], set1_unflattened[65], set1_unflattened[64], set1_unflattened[63], set1_unflattened[62], set1_unflattened[61], set1_unflattened[60], set1_unflattened[59], set1_unflattened[58], set1_unflattened[57], set1_unflattened[56], set1_unflattened[55], set1_unflattened[54], set1_unflattened[53], set1_unflattened[52], set1_unflattened[51], set1_unflattened[50], set1_unflattened[49], set1_unflattened[48], set1_unflattened[47], set1_unflattened[46], set1_unflattened[45], set1_unflattened[44], set1_unflattened[43], set1_unflattened[42], set1_unflattened[41], set1_unflattened[40], set1_unflattened[39], set1_unflattened[38], set1_unflattened[37], set1_unflattened[36], set1_unflattened[35], set1_unflattened[34], set1_unflattened[33], set1_unflattened[32], set1_unflattened[31], set1_unflattened[30], set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[74], set2_unflattened[73], set2_unflattened[72], set2_unflattened[71], set2_unflattened[70], set2_unflattened[69], set2_unflattened[68], set2_unflattened[67], set2_unflattened[66], set2_unflattened[65], set2_unflattened[64], set2_unflattened[63], set2_unflattened[62], set2_unflattened[61], set2_unflattened[60], set2_unflattened[59], set2_unflattened[58], set2_unflattened[57], set2_unflattened[56], set2_unflattened[55], set2_unflattened[54], set2_unflattened[53], set2_unflattened[52], set2_unflattened[51], set2_unflattened[50], set2_unflattened[49], set2_unflattened[48], set2_unflattened[47], set2_unflattened[46], set2_unflattened[45], set2_unflattened[44], set2_unflattened[43], set2_unflattened[42], set2_unflattened[41], set2_unflattened[40], set2_unflattened[39], set2_unflattened[38], set2_unflattened[37], set2_unflattened[36], set2_unflattened[35], set2_unflattened[34], set2_unflattened[33], set2_unflattened[32], set2_unflattened[31], set2_unflattened[30], set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
