module min_hash(
  input wire [799:0] set1,
  input wire [799:0] set2,
  output wire [1607:0] out
);
  wire [15:0] set1_unflattened[50];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  assign set1_unflattened[30] = set1[495:480];
  assign set1_unflattened[31] = set1[511:496];
  assign set1_unflattened[32] = set1[527:512];
  assign set1_unflattened[33] = set1[543:528];
  assign set1_unflattened[34] = set1[559:544];
  assign set1_unflattened[35] = set1[575:560];
  assign set1_unflattened[36] = set1[591:576];
  assign set1_unflattened[37] = set1[607:592];
  assign set1_unflattened[38] = set1[623:608];
  assign set1_unflattened[39] = set1[639:624];
  assign set1_unflattened[40] = set1[655:640];
  assign set1_unflattened[41] = set1[671:656];
  assign set1_unflattened[42] = set1[687:672];
  assign set1_unflattened[43] = set1[703:688];
  assign set1_unflattened[44] = set1[719:704];
  assign set1_unflattened[45] = set1[735:720];
  assign set1_unflattened[46] = set1[751:736];
  assign set1_unflattened[47] = set1[767:752];
  assign set1_unflattened[48] = set1[783:768];
  assign set1_unflattened[49] = set1[799:784];
  wire [15:0] set2_unflattened[50];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  assign set2_unflattened[30] = set2[495:480];
  assign set2_unflattened[31] = set2[511:496];
  assign set2_unflattened[32] = set2[527:512];
  assign set2_unflattened[33] = set2[543:528];
  assign set2_unflattened[34] = set2[559:544];
  assign set2_unflattened[35] = set2[575:560];
  assign set2_unflattened[36] = set2[591:576];
  assign set2_unflattened[37] = set2[607:592];
  assign set2_unflattened[38] = set2[623:608];
  assign set2_unflattened[39] = set2[639:624];
  assign set2_unflattened[40] = set2[655:640];
  assign set2_unflattened[41] = set2[671:656];
  assign set2_unflattened[42] = set2[687:672];
  assign set2_unflattened[43] = set2[703:688];
  assign set2_unflattened[44] = set2[719:704];
  assign set2_unflattened[45] = set2[735:720];
  assign set2_unflattened[46] = set2[751:736];
  assign set2_unflattened[47] = set2[767:752];
  assign set2_unflattened[48] = set2[783:768];
  assign set2_unflattened[49] = set2[799:784];
  wire [15:0] array_index_239311;
  wire [15:0] array_index_239312;
  wire [15:0] array_index_239316;
  wire [1:0] concat_239317;
  wire [1:0] add_239320;
  wire [15:0] array_index_239324;
  wire [2:0] concat_239325;
  wire [2:0] add_239328;
  wire [15:0] array_index_239332;
  wire [3:0] concat_239333;
  wire [3:0] add_239336;
  wire [15:0] array_index_239340;
  wire [4:0] concat_239341;
  wire [4:0] add_239344;
  wire [15:0] array_index_239348;
  wire [5:0] concat_239349;
  wire [5:0] add_239352;
  wire [15:0] array_index_239356;
  wire [6:0] concat_239357;
  wire [6:0] add_239360;
  wire [15:0] array_index_239364;
  wire [7:0] concat_239365;
  wire [7:0] add_239369;
  wire [15:0] array_index_239370;
  wire [7:0] sel_239371;
  wire [7:0] add_239375;
  wire [15:0] array_index_239376;
  wire [7:0] sel_239377;
  wire [7:0] add_239381;
  wire [15:0] array_index_239382;
  wire [7:0] sel_239383;
  wire [7:0] add_239387;
  wire [15:0] array_index_239388;
  wire [7:0] sel_239389;
  wire [7:0] add_239393;
  wire [15:0] array_index_239394;
  wire [7:0] sel_239395;
  wire [7:0] add_239399;
  wire [15:0] array_index_239400;
  wire [7:0] sel_239401;
  wire [7:0] add_239405;
  wire [15:0] array_index_239406;
  wire [7:0] sel_239407;
  wire [7:0] add_239411;
  wire [15:0] array_index_239412;
  wire [7:0] sel_239413;
  wire [7:0] add_239417;
  wire [15:0] array_index_239418;
  wire [7:0] sel_239419;
  wire [7:0] add_239423;
  wire [15:0] array_index_239424;
  wire [7:0] sel_239425;
  wire [7:0] add_239429;
  wire [15:0] array_index_239430;
  wire [7:0] sel_239431;
  wire [7:0] add_239435;
  wire [15:0] array_index_239436;
  wire [7:0] sel_239437;
  wire [7:0] add_239441;
  wire [15:0] array_index_239442;
  wire [7:0] sel_239443;
  wire [7:0] add_239447;
  wire [15:0] array_index_239448;
  wire [7:0] sel_239449;
  wire [7:0] add_239453;
  wire [15:0] array_index_239454;
  wire [7:0] sel_239455;
  wire [7:0] add_239459;
  wire [15:0] array_index_239460;
  wire [7:0] sel_239461;
  wire [7:0] add_239465;
  wire [15:0] array_index_239466;
  wire [7:0] sel_239467;
  wire [7:0] add_239471;
  wire [15:0] array_index_239472;
  wire [7:0] sel_239473;
  wire [7:0] add_239477;
  wire [15:0] array_index_239478;
  wire [7:0] sel_239479;
  wire [7:0] add_239483;
  wire [15:0] array_index_239484;
  wire [7:0] sel_239485;
  wire [7:0] add_239489;
  wire [15:0] array_index_239490;
  wire [7:0] sel_239491;
  wire [7:0] add_239495;
  wire [15:0] array_index_239496;
  wire [7:0] sel_239497;
  wire [7:0] add_239501;
  wire [15:0] array_index_239502;
  wire [7:0] sel_239503;
  wire [7:0] add_239507;
  wire [15:0] array_index_239508;
  wire [7:0] sel_239509;
  wire [7:0] add_239513;
  wire [15:0] array_index_239514;
  wire [7:0] sel_239515;
  wire [7:0] add_239519;
  wire [15:0] array_index_239520;
  wire [7:0] sel_239521;
  wire [7:0] add_239525;
  wire [15:0] array_index_239526;
  wire [7:0] sel_239527;
  wire [7:0] add_239531;
  wire [15:0] array_index_239532;
  wire [7:0] sel_239533;
  wire [7:0] add_239537;
  wire [15:0] array_index_239538;
  wire [7:0] sel_239539;
  wire [7:0] add_239543;
  wire [15:0] array_index_239544;
  wire [7:0] sel_239545;
  wire [7:0] add_239549;
  wire [15:0] array_index_239550;
  wire [7:0] sel_239551;
  wire [7:0] add_239555;
  wire [15:0] array_index_239556;
  wire [7:0] sel_239557;
  wire [7:0] add_239561;
  wire [15:0] array_index_239562;
  wire [7:0] sel_239563;
  wire [7:0] add_239567;
  wire [15:0] array_index_239568;
  wire [7:0] sel_239569;
  wire [7:0] add_239573;
  wire [15:0] array_index_239574;
  wire [7:0] sel_239575;
  wire [7:0] add_239579;
  wire [15:0] array_index_239580;
  wire [7:0] sel_239581;
  wire [7:0] add_239585;
  wire [15:0] array_index_239586;
  wire [7:0] sel_239587;
  wire [7:0] add_239591;
  wire [15:0] array_index_239592;
  wire [7:0] sel_239593;
  wire [7:0] add_239597;
  wire [15:0] array_index_239598;
  wire [7:0] sel_239599;
  wire [7:0] add_239603;
  wire [15:0] array_index_239604;
  wire [7:0] sel_239605;
  wire [7:0] add_239609;
  wire [15:0] array_index_239610;
  wire [7:0] sel_239611;
  wire [7:0] add_239615;
  wire [15:0] array_index_239616;
  wire [7:0] sel_239617;
  wire [7:0] add_239621;
  wire [15:0] array_index_239622;
  wire [7:0] sel_239623;
  wire [7:0] add_239626;
  wire [7:0] sel_239627;
  wire [7:0] add_239630;
  wire [7:0] sel_239631;
  wire [7:0] add_239634;
  wire [7:0] sel_239635;
  wire [7:0] add_239638;
  wire [7:0] sel_239639;
  wire [7:0] add_239642;
  wire [7:0] sel_239643;
  wire [7:0] add_239646;
  wire [7:0] sel_239647;
  wire [7:0] add_239650;
  wire [7:0] sel_239651;
  wire [7:0] add_239654;
  wire [7:0] sel_239655;
  wire [7:0] add_239658;
  wire [7:0] sel_239659;
  wire [7:0] add_239662;
  wire [7:0] sel_239663;
  wire [7:0] add_239666;
  wire [7:0] sel_239667;
  wire [7:0] add_239670;
  wire [7:0] sel_239671;
  wire [7:0] add_239674;
  wire [7:0] sel_239675;
  wire [7:0] add_239678;
  wire [7:0] sel_239679;
  wire [7:0] add_239682;
  wire [7:0] sel_239683;
  wire [7:0] add_239686;
  wire [7:0] sel_239687;
  wire [7:0] add_239690;
  wire [7:0] sel_239691;
  wire [7:0] add_239694;
  wire [7:0] sel_239695;
  wire [7:0] add_239698;
  wire [7:0] sel_239699;
  wire [7:0] add_239702;
  wire [7:0] sel_239703;
  wire [7:0] add_239706;
  wire [7:0] sel_239707;
  wire [7:0] add_239710;
  wire [7:0] sel_239711;
  wire [7:0] add_239714;
  wire [7:0] sel_239715;
  wire [7:0] add_239718;
  wire [7:0] sel_239719;
  wire [7:0] add_239722;
  wire [7:0] sel_239723;
  wire [7:0] add_239726;
  wire [7:0] sel_239727;
  wire [7:0] add_239730;
  wire [7:0] sel_239731;
  wire [7:0] add_239734;
  wire [7:0] sel_239735;
  wire [7:0] add_239738;
  wire [7:0] sel_239739;
  wire [7:0] add_239742;
  wire [7:0] sel_239743;
  wire [7:0] add_239746;
  wire [7:0] sel_239747;
  wire [7:0] add_239750;
  wire [7:0] sel_239751;
  wire [7:0] add_239754;
  wire [7:0] sel_239755;
  wire [7:0] add_239758;
  wire [7:0] sel_239759;
  wire [7:0] add_239762;
  wire [7:0] sel_239763;
  wire [7:0] add_239766;
  wire [7:0] sel_239767;
  wire [7:0] add_239770;
  wire [7:0] sel_239771;
  wire [7:0] add_239774;
  wire [7:0] sel_239775;
  wire [7:0] add_239778;
  wire [7:0] sel_239779;
  wire [7:0] add_239782;
  wire [7:0] sel_239783;
  wire [7:0] add_239786;
  wire [7:0] sel_239787;
  wire [7:0] add_239790;
  wire [7:0] sel_239791;
  wire [7:0] add_239794;
  wire [7:0] sel_239795;
  wire [7:0] add_239798;
  wire [7:0] sel_239799;
  wire [7:0] add_239802;
  wire [7:0] sel_239803;
  wire [7:0] add_239806;
  wire [7:0] sel_239807;
  wire [7:0] add_239810;
  wire [7:0] sel_239811;
  wire [7:0] add_239814;
  wire [7:0] sel_239815;
  wire [7:0] add_239818;
  wire [7:0] sel_239819;
  wire [7:0] add_239823;
  wire [15:0] array_index_239824;
  wire [7:0] sel_239825;
  wire [7:0] add_239828;
  wire [7:0] sel_239829;
  wire [7:0] add_239832;
  wire [7:0] sel_239833;
  wire [7:0] add_239836;
  wire [7:0] sel_239837;
  wire [7:0] add_239840;
  wire [7:0] sel_239841;
  wire [7:0] add_239844;
  wire [7:0] sel_239845;
  wire [7:0] add_239848;
  wire [7:0] sel_239849;
  wire [7:0] add_239852;
  wire [7:0] sel_239853;
  wire [7:0] add_239856;
  wire [7:0] sel_239857;
  wire [7:0] add_239860;
  wire [7:0] sel_239861;
  wire [7:0] add_239864;
  wire [7:0] sel_239865;
  wire [7:0] add_239868;
  wire [7:0] sel_239869;
  wire [7:0] add_239872;
  wire [7:0] sel_239873;
  wire [7:0] add_239876;
  wire [7:0] sel_239877;
  wire [7:0] add_239880;
  wire [7:0] sel_239881;
  wire [7:0] add_239884;
  wire [7:0] sel_239885;
  wire [7:0] add_239888;
  wire [7:0] sel_239889;
  wire [7:0] add_239892;
  wire [7:0] sel_239893;
  wire [7:0] add_239896;
  wire [7:0] sel_239897;
  wire [7:0] add_239900;
  wire [7:0] sel_239901;
  wire [7:0] add_239904;
  wire [7:0] sel_239905;
  wire [7:0] add_239908;
  wire [7:0] sel_239909;
  wire [7:0] add_239912;
  wire [7:0] sel_239913;
  wire [7:0] add_239916;
  wire [7:0] sel_239917;
  wire [7:0] add_239920;
  wire [7:0] sel_239921;
  wire [7:0] add_239924;
  wire [7:0] sel_239925;
  wire [7:0] add_239928;
  wire [7:0] sel_239929;
  wire [7:0] add_239932;
  wire [7:0] sel_239933;
  wire [7:0] add_239936;
  wire [7:0] sel_239937;
  wire [7:0] add_239940;
  wire [7:0] sel_239941;
  wire [7:0] add_239944;
  wire [7:0] sel_239945;
  wire [7:0] add_239948;
  wire [7:0] sel_239949;
  wire [7:0] add_239952;
  wire [7:0] sel_239953;
  wire [7:0] add_239956;
  wire [7:0] sel_239957;
  wire [7:0] add_239960;
  wire [7:0] sel_239961;
  wire [7:0] add_239964;
  wire [7:0] sel_239965;
  wire [7:0] add_239968;
  wire [7:0] sel_239969;
  wire [7:0] add_239972;
  wire [7:0] sel_239973;
  wire [7:0] add_239976;
  wire [7:0] sel_239977;
  wire [7:0] add_239980;
  wire [7:0] sel_239981;
  wire [7:0] add_239984;
  wire [7:0] sel_239985;
  wire [7:0] add_239988;
  wire [7:0] sel_239989;
  wire [7:0] add_239992;
  wire [7:0] sel_239993;
  wire [7:0] add_239996;
  wire [7:0] sel_239997;
  wire [7:0] add_240000;
  wire [7:0] sel_240001;
  wire [7:0] add_240004;
  wire [7:0] sel_240005;
  wire [7:0] add_240008;
  wire [7:0] sel_240009;
  wire [7:0] add_240012;
  wire [7:0] sel_240013;
  wire [7:0] add_240016;
  wire [7:0] sel_240017;
  wire [7:0] add_240020;
  wire [7:0] sel_240021;
  wire [7:0] add_240025;
  wire [15:0] array_index_240026;
  wire [7:0] sel_240027;
  wire [7:0] add_240030;
  wire [7:0] sel_240031;
  wire [7:0] add_240034;
  wire [7:0] sel_240035;
  wire [7:0] add_240038;
  wire [7:0] sel_240039;
  wire [7:0] add_240042;
  wire [7:0] sel_240043;
  wire [7:0] add_240046;
  wire [7:0] sel_240047;
  wire [7:0] add_240050;
  wire [7:0] sel_240051;
  wire [7:0] add_240054;
  wire [7:0] sel_240055;
  wire [7:0] add_240058;
  wire [7:0] sel_240059;
  wire [7:0] add_240062;
  wire [7:0] sel_240063;
  wire [7:0] add_240066;
  wire [7:0] sel_240067;
  wire [7:0] add_240070;
  wire [7:0] sel_240071;
  wire [7:0] add_240074;
  wire [7:0] sel_240075;
  wire [7:0] add_240078;
  wire [7:0] sel_240079;
  wire [7:0] add_240082;
  wire [7:0] sel_240083;
  wire [7:0] add_240086;
  wire [7:0] sel_240087;
  wire [7:0] add_240090;
  wire [7:0] sel_240091;
  wire [7:0] add_240094;
  wire [7:0] sel_240095;
  wire [7:0] add_240098;
  wire [7:0] sel_240099;
  wire [7:0] add_240102;
  wire [7:0] sel_240103;
  wire [7:0] add_240106;
  wire [7:0] sel_240107;
  wire [7:0] add_240110;
  wire [7:0] sel_240111;
  wire [7:0] add_240114;
  wire [7:0] sel_240115;
  wire [7:0] add_240118;
  wire [7:0] sel_240119;
  wire [7:0] add_240122;
  wire [7:0] sel_240123;
  wire [7:0] add_240126;
  wire [7:0] sel_240127;
  wire [7:0] add_240130;
  wire [7:0] sel_240131;
  wire [7:0] add_240134;
  wire [7:0] sel_240135;
  wire [7:0] add_240138;
  wire [7:0] sel_240139;
  wire [7:0] add_240142;
  wire [7:0] sel_240143;
  wire [7:0] add_240146;
  wire [7:0] sel_240147;
  wire [7:0] add_240150;
  wire [7:0] sel_240151;
  wire [7:0] add_240154;
  wire [7:0] sel_240155;
  wire [7:0] add_240158;
  wire [7:0] sel_240159;
  wire [7:0] add_240162;
  wire [7:0] sel_240163;
  wire [7:0] add_240166;
  wire [7:0] sel_240167;
  wire [7:0] add_240170;
  wire [7:0] sel_240171;
  wire [7:0] add_240174;
  wire [7:0] sel_240175;
  wire [7:0] add_240178;
  wire [7:0] sel_240179;
  wire [7:0] add_240182;
  wire [7:0] sel_240183;
  wire [7:0] add_240186;
  wire [7:0] sel_240187;
  wire [7:0] add_240190;
  wire [7:0] sel_240191;
  wire [7:0] add_240194;
  wire [7:0] sel_240195;
  wire [7:0] add_240198;
  wire [7:0] sel_240199;
  wire [7:0] add_240202;
  wire [7:0] sel_240203;
  wire [7:0] add_240206;
  wire [7:0] sel_240207;
  wire [7:0] add_240210;
  wire [7:0] sel_240211;
  wire [7:0] add_240214;
  wire [7:0] sel_240215;
  wire [7:0] add_240218;
  wire [7:0] sel_240219;
  wire [7:0] add_240222;
  wire [7:0] sel_240223;
  wire [7:0] add_240227;
  wire [15:0] array_index_240228;
  wire [7:0] sel_240229;
  wire [7:0] add_240232;
  wire [7:0] sel_240233;
  wire [7:0] add_240236;
  wire [7:0] sel_240237;
  wire [7:0] add_240240;
  wire [7:0] sel_240241;
  wire [7:0] add_240244;
  wire [7:0] sel_240245;
  wire [7:0] add_240248;
  wire [7:0] sel_240249;
  wire [7:0] add_240252;
  wire [7:0] sel_240253;
  wire [7:0] add_240256;
  wire [7:0] sel_240257;
  wire [7:0] add_240260;
  wire [7:0] sel_240261;
  wire [7:0] add_240264;
  wire [7:0] sel_240265;
  wire [7:0] add_240268;
  wire [7:0] sel_240269;
  wire [7:0] add_240272;
  wire [7:0] sel_240273;
  wire [7:0] add_240276;
  wire [7:0] sel_240277;
  wire [7:0] add_240280;
  wire [7:0] sel_240281;
  wire [7:0] add_240284;
  wire [7:0] sel_240285;
  wire [7:0] add_240288;
  wire [7:0] sel_240289;
  wire [7:0] add_240292;
  wire [7:0] sel_240293;
  wire [7:0] add_240296;
  wire [7:0] sel_240297;
  wire [7:0] add_240300;
  wire [7:0] sel_240301;
  wire [7:0] add_240304;
  wire [7:0] sel_240305;
  wire [7:0] add_240308;
  wire [7:0] sel_240309;
  wire [7:0] add_240312;
  wire [7:0] sel_240313;
  wire [7:0] add_240316;
  wire [7:0] sel_240317;
  wire [7:0] add_240320;
  wire [7:0] sel_240321;
  wire [7:0] add_240324;
  wire [7:0] sel_240325;
  wire [7:0] add_240328;
  wire [7:0] sel_240329;
  wire [7:0] add_240332;
  wire [7:0] sel_240333;
  wire [7:0] add_240336;
  wire [7:0] sel_240337;
  wire [7:0] add_240340;
  wire [7:0] sel_240341;
  wire [7:0] add_240344;
  wire [7:0] sel_240345;
  wire [7:0] add_240348;
  wire [7:0] sel_240349;
  wire [7:0] add_240352;
  wire [7:0] sel_240353;
  wire [7:0] add_240356;
  wire [7:0] sel_240357;
  wire [7:0] add_240360;
  wire [7:0] sel_240361;
  wire [7:0] add_240364;
  wire [7:0] sel_240365;
  wire [7:0] add_240368;
  wire [7:0] sel_240369;
  wire [7:0] add_240372;
  wire [7:0] sel_240373;
  wire [7:0] add_240376;
  wire [7:0] sel_240377;
  wire [7:0] add_240380;
  wire [7:0] sel_240381;
  wire [7:0] add_240384;
  wire [7:0] sel_240385;
  wire [7:0] add_240388;
  wire [7:0] sel_240389;
  wire [7:0] add_240392;
  wire [7:0] sel_240393;
  wire [7:0] add_240396;
  wire [7:0] sel_240397;
  wire [7:0] add_240400;
  wire [7:0] sel_240401;
  wire [7:0] add_240404;
  wire [7:0] sel_240405;
  wire [7:0] add_240408;
  wire [7:0] sel_240409;
  wire [7:0] add_240412;
  wire [7:0] sel_240413;
  wire [7:0] add_240416;
  wire [7:0] sel_240417;
  wire [7:0] add_240420;
  wire [7:0] sel_240421;
  wire [7:0] add_240424;
  wire [7:0] sel_240425;
  wire [7:0] add_240429;
  wire [15:0] array_index_240430;
  wire [7:0] sel_240431;
  wire [7:0] add_240434;
  wire [7:0] sel_240435;
  wire [7:0] add_240438;
  wire [7:0] sel_240439;
  wire [7:0] add_240442;
  wire [7:0] sel_240443;
  wire [7:0] add_240446;
  wire [7:0] sel_240447;
  wire [7:0] add_240450;
  wire [7:0] sel_240451;
  wire [7:0] add_240454;
  wire [7:0] sel_240455;
  wire [7:0] add_240458;
  wire [7:0] sel_240459;
  wire [7:0] add_240462;
  wire [7:0] sel_240463;
  wire [7:0] add_240466;
  wire [7:0] sel_240467;
  wire [7:0] add_240470;
  wire [7:0] sel_240471;
  wire [7:0] add_240474;
  wire [7:0] sel_240475;
  wire [7:0] add_240478;
  wire [7:0] sel_240479;
  wire [7:0] add_240482;
  wire [7:0] sel_240483;
  wire [7:0] add_240486;
  wire [7:0] sel_240487;
  wire [7:0] add_240490;
  wire [7:0] sel_240491;
  wire [7:0] add_240494;
  wire [7:0] sel_240495;
  wire [7:0] add_240498;
  wire [7:0] sel_240499;
  wire [7:0] add_240502;
  wire [7:0] sel_240503;
  wire [7:0] add_240506;
  wire [7:0] sel_240507;
  wire [7:0] add_240510;
  wire [7:0] sel_240511;
  wire [7:0] add_240514;
  wire [7:0] sel_240515;
  wire [7:0] add_240518;
  wire [7:0] sel_240519;
  wire [7:0] add_240522;
  wire [7:0] sel_240523;
  wire [7:0] add_240526;
  wire [7:0] sel_240527;
  wire [7:0] add_240530;
  wire [7:0] sel_240531;
  wire [7:0] add_240534;
  wire [7:0] sel_240535;
  wire [7:0] add_240538;
  wire [7:0] sel_240539;
  wire [7:0] add_240542;
  wire [7:0] sel_240543;
  wire [7:0] add_240546;
  wire [7:0] sel_240547;
  wire [7:0] add_240550;
  wire [7:0] sel_240551;
  wire [7:0] add_240554;
  wire [7:0] sel_240555;
  wire [7:0] add_240558;
  wire [7:0] sel_240559;
  wire [7:0] add_240562;
  wire [7:0] sel_240563;
  wire [7:0] add_240566;
  wire [7:0] sel_240567;
  wire [7:0] add_240570;
  wire [7:0] sel_240571;
  wire [7:0] add_240574;
  wire [7:0] sel_240575;
  wire [7:0] add_240578;
  wire [7:0] sel_240579;
  wire [7:0] add_240582;
  wire [7:0] sel_240583;
  wire [7:0] add_240586;
  wire [7:0] sel_240587;
  wire [7:0] add_240590;
  wire [7:0] sel_240591;
  wire [7:0] add_240594;
  wire [7:0] sel_240595;
  wire [7:0] add_240598;
  wire [7:0] sel_240599;
  wire [7:0] add_240602;
  wire [7:0] sel_240603;
  wire [7:0] add_240606;
  wire [7:0] sel_240607;
  wire [7:0] add_240610;
  wire [7:0] sel_240611;
  wire [7:0] add_240614;
  wire [7:0] sel_240615;
  wire [7:0] add_240618;
  wire [7:0] sel_240619;
  wire [7:0] add_240622;
  wire [7:0] sel_240623;
  wire [7:0] add_240626;
  wire [7:0] sel_240627;
  wire [7:0] add_240631;
  wire [15:0] array_index_240632;
  wire [7:0] sel_240633;
  wire [7:0] add_240636;
  wire [7:0] sel_240637;
  wire [7:0] add_240640;
  wire [7:0] sel_240641;
  wire [7:0] add_240644;
  wire [7:0] sel_240645;
  wire [7:0] add_240648;
  wire [7:0] sel_240649;
  wire [7:0] add_240652;
  wire [7:0] sel_240653;
  wire [7:0] add_240656;
  wire [7:0] sel_240657;
  wire [7:0] add_240660;
  wire [7:0] sel_240661;
  wire [7:0] add_240664;
  wire [7:0] sel_240665;
  wire [7:0] add_240668;
  wire [7:0] sel_240669;
  wire [7:0] add_240672;
  wire [7:0] sel_240673;
  wire [7:0] add_240676;
  wire [7:0] sel_240677;
  wire [7:0] add_240680;
  wire [7:0] sel_240681;
  wire [7:0] add_240684;
  wire [7:0] sel_240685;
  wire [7:0] add_240688;
  wire [7:0] sel_240689;
  wire [7:0] add_240692;
  wire [7:0] sel_240693;
  wire [7:0] add_240696;
  wire [7:0] sel_240697;
  wire [7:0] add_240700;
  wire [7:0] sel_240701;
  wire [7:0] add_240704;
  wire [7:0] sel_240705;
  wire [7:0] add_240708;
  wire [7:0] sel_240709;
  wire [7:0] add_240712;
  wire [7:0] sel_240713;
  wire [7:0] add_240716;
  wire [7:0] sel_240717;
  wire [7:0] add_240720;
  wire [7:0] sel_240721;
  wire [7:0] add_240724;
  wire [7:0] sel_240725;
  wire [7:0] add_240728;
  wire [7:0] sel_240729;
  wire [7:0] add_240732;
  wire [7:0] sel_240733;
  wire [7:0] add_240736;
  wire [7:0] sel_240737;
  wire [7:0] add_240740;
  wire [7:0] sel_240741;
  wire [7:0] add_240744;
  wire [7:0] sel_240745;
  wire [7:0] add_240748;
  wire [7:0] sel_240749;
  wire [7:0] add_240752;
  wire [7:0] sel_240753;
  wire [7:0] add_240756;
  wire [7:0] sel_240757;
  wire [7:0] add_240760;
  wire [7:0] sel_240761;
  wire [7:0] add_240764;
  wire [7:0] sel_240765;
  wire [7:0] add_240768;
  wire [7:0] sel_240769;
  wire [7:0] add_240772;
  wire [7:0] sel_240773;
  wire [7:0] add_240776;
  wire [7:0] sel_240777;
  wire [7:0] add_240780;
  wire [7:0] sel_240781;
  wire [7:0] add_240784;
  wire [7:0] sel_240785;
  wire [7:0] add_240788;
  wire [7:0] sel_240789;
  wire [7:0] add_240792;
  wire [7:0] sel_240793;
  wire [7:0] add_240796;
  wire [7:0] sel_240797;
  wire [7:0] add_240800;
  wire [7:0] sel_240801;
  wire [7:0] add_240804;
  wire [7:0] sel_240805;
  wire [7:0] add_240808;
  wire [7:0] sel_240809;
  wire [7:0] add_240812;
  wire [7:0] sel_240813;
  wire [7:0] add_240816;
  wire [7:0] sel_240817;
  wire [7:0] add_240820;
  wire [7:0] sel_240821;
  wire [7:0] add_240824;
  wire [7:0] sel_240825;
  wire [7:0] add_240828;
  wire [7:0] sel_240829;
  wire [7:0] add_240833;
  wire [15:0] array_index_240834;
  wire [7:0] sel_240835;
  wire [7:0] add_240838;
  wire [7:0] sel_240839;
  wire [7:0] add_240842;
  wire [7:0] sel_240843;
  wire [7:0] add_240846;
  wire [7:0] sel_240847;
  wire [7:0] add_240850;
  wire [7:0] sel_240851;
  wire [7:0] add_240854;
  wire [7:0] sel_240855;
  wire [7:0] add_240858;
  wire [7:0] sel_240859;
  wire [7:0] add_240862;
  wire [7:0] sel_240863;
  wire [7:0] add_240866;
  wire [7:0] sel_240867;
  wire [7:0] add_240870;
  wire [7:0] sel_240871;
  wire [7:0] add_240874;
  wire [7:0] sel_240875;
  wire [7:0] add_240878;
  wire [7:0] sel_240879;
  wire [7:0] add_240882;
  wire [7:0] sel_240883;
  wire [7:0] add_240886;
  wire [7:0] sel_240887;
  wire [7:0] add_240890;
  wire [7:0] sel_240891;
  wire [7:0] add_240894;
  wire [7:0] sel_240895;
  wire [7:0] add_240898;
  wire [7:0] sel_240899;
  wire [7:0] add_240902;
  wire [7:0] sel_240903;
  wire [7:0] add_240906;
  wire [7:0] sel_240907;
  wire [7:0] add_240910;
  wire [7:0] sel_240911;
  wire [7:0] add_240914;
  wire [7:0] sel_240915;
  wire [7:0] add_240918;
  wire [7:0] sel_240919;
  wire [7:0] add_240922;
  wire [7:0] sel_240923;
  wire [7:0] add_240926;
  wire [7:0] sel_240927;
  wire [7:0] add_240930;
  wire [7:0] sel_240931;
  wire [7:0] add_240934;
  wire [7:0] sel_240935;
  wire [7:0] add_240938;
  wire [7:0] sel_240939;
  wire [7:0] add_240942;
  wire [7:0] sel_240943;
  wire [7:0] add_240946;
  wire [7:0] sel_240947;
  wire [7:0] add_240950;
  wire [7:0] sel_240951;
  wire [7:0] add_240954;
  wire [7:0] sel_240955;
  wire [7:0] add_240958;
  wire [7:0] sel_240959;
  wire [7:0] add_240962;
  wire [7:0] sel_240963;
  wire [7:0] add_240966;
  wire [7:0] sel_240967;
  wire [7:0] add_240970;
  wire [7:0] sel_240971;
  wire [7:0] add_240974;
  wire [7:0] sel_240975;
  wire [7:0] add_240978;
  wire [7:0] sel_240979;
  wire [7:0] add_240982;
  wire [7:0] sel_240983;
  wire [7:0] add_240986;
  wire [7:0] sel_240987;
  wire [7:0] add_240990;
  wire [7:0] sel_240991;
  wire [7:0] add_240994;
  wire [7:0] sel_240995;
  wire [7:0] add_240998;
  wire [7:0] sel_240999;
  wire [7:0] add_241002;
  wire [7:0] sel_241003;
  wire [7:0] add_241006;
  wire [7:0] sel_241007;
  wire [7:0] add_241010;
  wire [7:0] sel_241011;
  wire [7:0] add_241014;
  wire [7:0] sel_241015;
  wire [7:0] add_241018;
  wire [7:0] sel_241019;
  wire [7:0] add_241022;
  wire [7:0] sel_241023;
  wire [7:0] add_241026;
  wire [7:0] sel_241027;
  wire [7:0] add_241030;
  wire [7:0] sel_241031;
  wire [7:0] add_241035;
  wire [15:0] array_index_241036;
  wire [7:0] sel_241037;
  wire [7:0] add_241040;
  wire [7:0] sel_241041;
  wire [7:0] add_241044;
  wire [7:0] sel_241045;
  wire [7:0] add_241048;
  wire [7:0] sel_241049;
  wire [7:0] add_241052;
  wire [7:0] sel_241053;
  wire [7:0] add_241056;
  wire [7:0] sel_241057;
  wire [7:0] add_241060;
  wire [7:0] sel_241061;
  wire [7:0] add_241064;
  wire [7:0] sel_241065;
  wire [7:0] add_241068;
  wire [7:0] sel_241069;
  wire [7:0] add_241072;
  wire [7:0] sel_241073;
  wire [7:0] add_241076;
  wire [7:0] sel_241077;
  wire [7:0] add_241080;
  wire [7:0] sel_241081;
  wire [7:0] add_241084;
  wire [7:0] sel_241085;
  wire [7:0] add_241088;
  wire [7:0] sel_241089;
  wire [7:0] add_241092;
  wire [7:0] sel_241093;
  wire [7:0] add_241096;
  wire [7:0] sel_241097;
  wire [7:0] add_241100;
  wire [7:0] sel_241101;
  wire [7:0] add_241104;
  wire [7:0] sel_241105;
  wire [7:0] add_241108;
  wire [7:0] sel_241109;
  wire [7:0] add_241112;
  wire [7:0] sel_241113;
  wire [7:0] add_241116;
  wire [7:0] sel_241117;
  wire [7:0] add_241120;
  wire [7:0] sel_241121;
  wire [7:0] add_241124;
  wire [7:0] sel_241125;
  wire [7:0] add_241128;
  wire [7:0] sel_241129;
  wire [7:0] add_241132;
  wire [7:0] sel_241133;
  wire [7:0] add_241136;
  wire [7:0] sel_241137;
  wire [7:0] add_241140;
  wire [7:0] sel_241141;
  wire [7:0] add_241144;
  wire [7:0] sel_241145;
  wire [7:0] add_241148;
  wire [7:0] sel_241149;
  wire [7:0] add_241152;
  wire [7:0] sel_241153;
  wire [7:0] add_241156;
  wire [7:0] sel_241157;
  wire [7:0] add_241160;
  wire [7:0] sel_241161;
  wire [7:0] add_241164;
  wire [7:0] sel_241165;
  wire [7:0] add_241168;
  wire [7:0] sel_241169;
  wire [7:0] add_241172;
  wire [7:0] sel_241173;
  wire [7:0] add_241176;
  wire [7:0] sel_241177;
  wire [7:0] add_241180;
  wire [7:0] sel_241181;
  wire [7:0] add_241184;
  wire [7:0] sel_241185;
  wire [7:0] add_241188;
  wire [7:0] sel_241189;
  wire [7:0] add_241192;
  wire [7:0] sel_241193;
  wire [7:0] add_241196;
  wire [7:0] sel_241197;
  wire [7:0] add_241200;
  wire [7:0] sel_241201;
  wire [7:0] add_241204;
  wire [7:0] sel_241205;
  wire [7:0] add_241208;
  wire [7:0] sel_241209;
  wire [7:0] add_241212;
  wire [7:0] sel_241213;
  wire [7:0] add_241216;
  wire [7:0] sel_241217;
  wire [7:0] add_241220;
  wire [7:0] sel_241221;
  wire [7:0] add_241224;
  wire [7:0] sel_241225;
  wire [7:0] add_241228;
  wire [7:0] sel_241229;
  wire [7:0] add_241232;
  wire [7:0] sel_241233;
  wire [7:0] add_241237;
  wire [15:0] array_index_241238;
  wire [7:0] sel_241239;
  wire [7:0] add_241242;
  wire [7:0] sel_241243;
  wire [7:0] add_241246;
  wire [7:0] sel_241247;
  wire [7:0] add_241250;
  wire [7:0] sel_241251;
  wire [7:0] add_241254;
  wire [7:0] sel_241255;
  wire [7:0] add_241258;
  wire [7:0] sel_241259;
  wire [7:0] add_241262;
  wire [7:0] sel_241263;
  wire [7:0] add_241266;
  wire [7:0] sel_241267;
  wire [7:0] add_241270;
  wire [7:0] sel_241271;
  wire [7:0] add_241274;
  wire [7:0] sel_241275;
  wire [7:0] add_241278;
  wire [7:0] sel_241279;
  wire [7:0] add_241282;
  wire [7:0] sel_241283;
  wire [7:0] add_241286;
  wire [7:0] sel_241287;
  wire [7:0] add_241290;
  wire [7:0] sel_241291;
  wire [7:0] add_241294;
  wire [7:0] sel_241295;
  wire [7:0] add_241298;
  wire [7:0] sel_241299;
  wire [7:0] add_241302;
  wire [7:0] sel_241303;
  wire [7:0] add_241306;
  wire [7:0] sel_241307;
  wire [7:0] add_241310;
  wire [7:0] sel_241311;
  wire [7:0] add_241314;
  wire [7:0] sel_241315;
  wire [7:0] add_241318;
  wire [7:0] sel_241319;
  wire [7:0] add_241322;
  wire [7:0] sel_241323;
  wire [7:0] add_241326;
  wire [7:0] sel_241327;
  wire [7:0] add_241330;
  wire [7:0] sel_241331;
  wire [7:0] add_241334;
  wire [7:0] sel_241335;
  wire [7:0] add_241338;
  wire [7:0] sel_241339;
  wire [7:0] add_241342;
  wire [7:0] sel_241343;
  wire [7:0] add_241346;
  wire [7:0] sel_241347;
  wire [7:0] add_241350;
  wire [7:0] sel_241351;
  wire [7:0] add_241354;
  wire [7:0] sel_241355;
  wire [7:0] add_241358;
  wire [7:0] sel_241359;
  wire [7:0] add_241362;
  wire [7:0] sel_241363;
  wire [7:0] add_241366;
  wire [7:0] sel_241367;
  wire [7:0] add_241370;
  wire [7:0] sel_241371;
  wire [7:0] add_241374;
  wire [7:0] sel_241375;
  wire [7:0] add_241378;
  wire [7:0] sel_241379;
  wire [7:0] add_241382;
  wire [7:0] sel_241383;
  wire [7:0] add_241386;
  wire [7:0] sel_241387;
  wire [7:0] add_241390;
  wire [7:0] sel_241391;
  wire [7:0] add_241394;
  wire [7:0] sel_241395;
  wire [7:0] add_241398;
  wire [7:0] sel_241399;
  wire [7:0] add_241402;
  wire [7:0] sel_241403;
  wire [7:0] add_241406;
  wire [7:0] sel_241407;
  wire [7:0] add_241410;
  wire [7:0] sel_241411;
  wire [7:0] add_241414;
  wire [7:0] sel_241415;
  wire [7:0] add_241418;
  wire [7:0] sel_241419;
  wire [7:0] add_241422;
  wire [7:0] sel_241423;
  wire [7:0] add_241426;
  wire [7:0] sel_241427;
  wire [7:0] add_241430;
  wire [7:0] sel_241431;
  wire [7:0] add_241434;
  wire [7:0] sel_241435;
  wire [7:0] add_241439;
  wire [15:0] array_index_241440;
  wire [7:0] sel_241441;
  wire [7:0] add_241444;
  wire [7:0] sel_241445;
  wire [7:0] add_241448;
  wire [7:0] sel_241449;
  wire [7:0] add_241452;
  wire [7:0] sel_241453;
  wire [7:0] add_241456;
  wire [7:0] sel_241457;
  wire [7:0] add_241460;
  wire [7:0] sel_241461;
  wire [7:0] add_241464;
  wire [7:0] sel_241465;
  wire [7:0] add_241468;
  wire [7:0] sel_241469;
  wire [7:0] add_241472;
  wire [7:0] sel_241473;
  wire [7:0] add_241476;
  wire [7:0] sel_241477;
  wire [7:0] add_241480;
  wire [7:0] sel_241481;
  wire [7:0] add_241484;
  wire [7:0] sel_241485;
  wire [7:0] add_241488;
  wire [7:0] sel_241489;
  wire [7:0] add_241492;
  wire [7:0] sel_241493;
  wire [7:0] add_241496;
  wire [7:0] sel_241497;
  wire [7:0] add_241500;
  wire [7:0] sel_241501;
  wire [7:0] add_241504;
  wire [7:0] sel_241505;
  wire [7:0] add_241508;
  wire [7:0] sel_241509;
  wire [7:0] add_241512;
  wire [7:0] sel_241513;
  wire [7:0] add_241516;
  wire [7:0] sel_241517;
  wire [7:0] add_241520;
  wire [7:0] sel_241521;
  wire [7:0] add_241524;
  wire [7:0] sel_241525;
  wire [7:0] add_241528;
  wire [7:0] sel_241529;
  wire [7:0] add_241532;
  wire [7:0] sel_241533;
  wire [7:0] add_241536;
  wire [7:0] sel_241537;
  wire [7:0] add_241540;
  wire [7:0] sel_241541;
  wire [7:0] add_241544;
  wire [7:0] sel_241545;
  wire [7:0] add_241548;
  wire [7:0] sel_241549;
  wire [7:0] add_241552;
  wire [7:0] sel_241553;
  wire [7:0] add_241556;
  wire [7:0] sel_241557;
  wire [7:0] add_241560;
  wire [7:0] sel_241561;
  wire [7:0] add_241564;
  wire [7:0] sel_241565;
  wire [7:0] add_241568;
  wire [7:0] sel_241569;
  wire [7:0] add_241572;
  wire [7:0] sel_241573;
  wire [7:0] add_241576;
  wire [7:0] sel_241577;
  wire [7:0] add_241580;
  wire [7:0] sel_241581;
  wire [7:0] add_241584;
  wire [7:0] sel_241585;
  wire [7:0] add_241588;
  wire [7:0] sel_241589;
  wire [7:0] add_241592;
  wire [7:0] sel_241593;
  wire [7:0] add_241596;
  wire [7:0] sel_241597;
  wire [7:0] add_241600;
  wire [7:0] sel_241601;
  wire [7:0] add_241604;
  wire [7:0] sel_241605;
  wire [7:0] add_241608;
  wire [7:0] sel_241609;
  wire [7:0] add_241612;
  wire [7:0] sel_241613;
  wire [7:0] add_241616;
  wire [7:0] sel_241617;
  wire [7:0] add_241620;
  wire [7:0] sel_241621;
  wire [7:0] add_241624;
  wire [7:0] sel_241625;
  wire [7:0] add_241628;
  wire [7:0] sel_241629;
  wire [7:0] add_241632;
  wire [7:0] sel_241633;
  wire [7:0] add_241636;
  wire [7:0] sel_241637;
  wire [7:0] add_241641;
  wire [15:0] array_index_241642;
  wire [7:0] sel_241643;
  wire [7:0] add_241646;
  wire [7:0] sel_241647;
  wire [7:0] add_241650;
  wire [7:0] sel_241651;
  wire [7:0] add_241654;
  wire [7:0] sel_241655;
  wire [7:0] add_241658;
  wire [7:0] sel_241659;
  wire [7:0] add_241662;
  wire [7:0] sel_241663;
  wire [7:0] add_241666;
  wire [7:0] sel_241667;
  wire [7:0] add_241670;
  wire [7:0] sel_241671;
  wire [7:0] add_241674;
  wire [7:0] sel_241675;
  wire [7:0] add_241678;
  wire [7:0] sel_241679;
  wire [7:0] add_241682;
  wire [7:0] sel_241683;
  wire [7:0] add_241686;
  wire [7:0] sel_241687;
  wire [7:0] add_241690;
  wire [7:0] sel_241691;
  wire [7:0] add_241694;
  wire [7:0] sel_241695;
  wire [7:0] add_241698;
  wire [7:0] sel_241699;
  wire [7:0] add_241702;
  wire [7:0] sel_241703;
  wire [7:0] add_241706;
  wire [7:0] sel_241707;
  wire [7:0] add_241710;
  wire [7:0] sel_241711;
  wire [7:0] add_241714;
  wire [7:0] sel_241715;
  wire [7:0] add_241718;
  wire [7:0] sel_241719;
  wire [7:0] add_241722;
  wire [7:0] sel_241723;
  wire [7:0] add_241726;
  wire [7:0] sel_241727;
  wire [7:0] add_241730;
  wire [7:0] sel_241731;
  wire [7:0] add_241734;
  wire [7:0] sel_241735;
  wire [7:0] add_241738;
  wire [7:0] sel_241739;
  wire [7:0] add_241742;
  wire [7:0] sel_241743;
  wire [7:0] add_241746;
  wire [7:0] sel_241747;
  wire [7:0] add_241750;
  wire [7:0] sel_241751;
  wire [7:0] add_241754;
  wire [7:0] sel_241755;
  wire [7:0] add_241758;
  wire [7:0] sel_241759;
  wire [7:0] add_241762;
  wire [7:0] sel_241763;
  wire [7:0] add_241766;
  wire [7:0] sel_241767;
  wire [7:0] add_241770;
  wire [7:0] sel_241771;
  wire [7:0] add_241774;
  wire [7:0] sel_241775;
  wire [7:0] add_241778;
  wire [7:0] sel_241779;
  wire [7:0] add_241782;
  wire [7:0] sel_241783;
  wire [7:0] add_241786;
  wire [7:0] sel_241787;
  wire [7:0] add_241790;
  wire [7:0] sel_241791;
  wire [7:0] add_241794;
  wire [7:0] sel_241795;
  wire [7:0] add_241798;
  wire [7:0] sel_241799;
  wire [7:0] add_241802;
  wire [7:0] sel_241803;
  wire [7:0] add_241806;
  wire [7:0] sel_241807;
  wire [7:0] add_241810;
  wire [7:0] sel_241811;
  wire [7:0] add_241814;
  wire [7:0] sel_241815;
  wire [7:0] add_241818;
  wire [7:0] sel_241819;
  wire [7:0] add_241822;
  wire [7:0] sel_241823;
  wire [7:0] add_241826;
  wire [7:0] sel_241827;
  wire [7:0] add_241830;
  wire [7:0] sel_241831;
  wire [7:0] add_241834;
  wire [7:0] sel_241835;
  wire [7:0] add_241838;
  wire [7:0] sel_241839;
  wire [7:0] add_241843;
  wire [15:0] array_index_241844;
  wire [7:0] sel_241845;
  wire [7:0] add_241848;
  wire [7:0] sel_241849;
  wire [7:0] add_241852;
  wire [7:0] sel_241853;
  wire [7:0] add_241856;
  wire [7:0] sel_241857;
  wire [7:0] add_241860;
  wire [7:0] sel_241861;
  wire [7:0] add_241864;
  wire [7:0] sel_241865;
  wire [7:0] add_241868;
  wire [7:0] sel_241869;
  wire [7:0] add_241872;
  wire [7:0] sel_241873;
  wire [7:0] add_241876;
  wire [7:0] sel_241877;
  wire [7:0] add_241880;
  wire [7:0] sel_241881;
  wire [7:0] add_241884;
  wire [7:0] sel_241885;
  wire [7:0] add_241888;
  wire [7:0] sel_241889;
  wire [7:0] add_241892;
  wire [7:0] sel_241893;
  wire [7:0] add_241896;
  wire [7:0] sel_241897;
  wire [7:0] add_241900;
  wire [7:0] sel_241901;
  wire [7:0] add_241904;
  wire [7:0] sel_241905;
  wire [7:0] add_241908;
  wire [7:0] sel_241909;
  wire [7:0] add_241912;
  wire [7:0] sel_241913;
  wire [7:0] add_241916;
  wire [7:0] sel_241917;
  wire [7:0] add_241920;
  wire [7:0] sel_241921;
  wire [7:0] add_241924;
  wire [7:0] sel_241925;
  wire [7:0] add_241928;
  wire [7:0] sel_241929;
  wire [7:0] add_241932;
  wire [7:0] sel_241933;
  wire [7:0] add_241936;
  wire [7:0] sel_241937;
  wire [7:0] add_241940;
  wire [7:0] sel_241941;
  wire [7:0] add_241944;
  wire [7:0] sel_241945;
  wire [7:0] add_241948;
  wire [7:0] sel_241949;
  wire [7:0] add_241952;
  wire [7:0] sel_241953;
  wire [7:0] add_241956;
  wire [7:0] sel_241957;
  wire [7:0] add_241960;
  wire [7:0] sel_241961;
  wire [7:0] add_241964;
  wire [7:0] sel_241965;
  wire [7:0] add_241968;
  wire [7:0] sel_241969;
  wire [7:0] add_241972;
  wire [7:0] sel_241973;
  wire [7:0] add_241976;
  wire [7:0] sel_241977;
  wire [7:0] add_241980;
  wire [7:0] sel_241981;
  wire [7:0] add_241984;
  wire [7:0] sel_241985;
  wire [7:0] add_241988;
  wire [7:0] sel_241989;
  wire [7:0] add_241992;
  wire [7:0] sel_241993;
  wire [7:0] add_241996;
  wire [7:0] sel_241997;
  wire [7:0] add_242000;
  wire [7:0] sel_242001;
  wire [7:0] add_242004;
  wire [7:0] sel_242005;
  wire [7:0] add_242008;
  wire [7:0] sel_242009;
  wire [7:0] add_242012;
  wire [7:0] sel_242013;
  wire [7:0] add_242016;
  wire [7:0] sel_242017;
  wire [7:0] add_242020;
  wire [7:0] sel_242021;
  wire [7:0] add_242024;
  wire [7:0] sel_242025;
  wire [7:0] add_242028;
  wire [7:0] sel_242029;
  wire [7:0] add_242032;
  wire [7:0] sel_242033;
  wire [7:0] add_242036;
  wire [7:0] sel_242037;
  wire [7:0] add_242040;
  wire [7:0] sel_242041;
  wire [7:0] add_242045;
  wire [15:0] array_index_242046;
  wire [7:0] sel_242047;
  wire [7:0] add_242050;
  wire [7:0] sel_242051;
  wire [7:0] add_242054;
  wire [7:0] sel_242055;
  wire [7:0] add_242058;
  wire [7:0] sel_242059;
  wire [7:0] add_242062;
  wire [7:0] sel_242063;
  wire [7:0] add_242066;
  wire [7:0] sel_242067;
  wire [7:0] add_242070;
  wire [7:0] sel_242071;
  wire [7:0] add_242074;
  wire [7:0] sel_242075;
  wire [7:0] add_242078;
  wire [7:0] sel_242079;
  wire [7:0] add_242082;
  wire [7:0] sel_242083;
  wire [7:0] add_242086;
  wire [7:0] sel_242087;
  wire [7:0] add_242090;
  wire [7:0] sel_242091;
  wire [7:0] add_242094;
  wire [7:0] sel_242095;
  wire [7:0] add_242098;
  wire [7:0] sel_242099;
  wire [7:0] add_242102;
  wire [7:0] sel_242103;
  wire [7:0] add_242106;
  wire [7:0] sel_242107;
  wire [7:0] add_242110;
  wire [7:0] sel_242111;
  wire [7:0] add_242114;
  wire [7:0] sel_242115;
  wire [7:0] add_242118;
  wire [7:0] sel_242119;
  wire [7:0] add_242122;
  wire [7:0] sel_242123;
  wire [7:0] add_242126;
  wire [7:0] sel_242127;
  wire [7:0] add_242130;
  wire [7:0] sel_242131;
  wire [7:0] add_242134;
  wire [7:0] sel_242135;
  wire [7:0] add_242138;
  wire [7:0] sel_242139;
  wire [7:0] add_242142;
  wire [7:0] sel_242143;
  wire [7:0] add_242146;
  wire [7:0] sel_242147;
  wire [7:0] add_242150;
  wire [7:0] sel_242151;
  wire [7:0] add_242154;
  wire [7:0] sel_242155;
  wire [7:0] add_242158;
  wire [7:0] sel_242159;
  wire [7:0] add_242162;
  wire [7:0] sel_242163;
  wire [7:0] add_242166;
  wire [7:0] sel_242167;
  wire [7:0] add_242170;
  wire [7:0] sel_242171;
  wire [7:0] add_242174;
  wire [7:0] sel_242175;
  wire [7:0] add_242178;
  wire [7:0] sel_242179;
  wire [7:0] add_242182;
  wire [7:0] sel_242183;
  wire [7:0] add_242186;
  wire [7:0] sel_242187;
  wire [7:0] add_242190;
  wire [7:0] sel_242191;
  wire [7:0] add_242194;
  wire [7:0] sel_242195;
  wire [7:0] add_242198;
  wire [7:0] sel_242199;
  wire [7:0] add_242202;
  wire [7:0] sel_242203;
  wire [7:0] add_242206;
  wire [7:0] sel_242207;
  wire [7:0] add_242210;
  wire [7:0] sel_242211;
  wire [7:0] add_242214;
  wire [7:0] sel_242215;
  wire [7:0] add_242218;
  wire [7:0] sel_242219;
  wire [7:0] add_242222;
  wire [7:0] sel_242223;
  wire [7:0] add_242226;
  wire [7:0] sel_242227;
  wire [7:0] add_242230;
  wire [7:0] sel_242231;
  wire [7:0] add_242234;
  wire [7:0] sel_242235;
  wire [7:0] add_242238;
  wire [7:0] sel_242239;
  wire [7:0] add_242242;
  wire [7:0] sel_242243;
  wire [7:0] add_242247;
  wire [15:0] array_index_242248;
  wire [7:0] sel_242249;
  wire [7:0] add_242252;
  wire [7:0] sel_242253;
  wire [7:0] add_242256;
  wire [7:0] sel_242257;
  wire [7:0] add_242260;
  wire [7:0] sel_242261;
  wire [7:0] add_242264;
  wire [7:0] sel_242265;
  wire [7:0] add_242268;
  wire [7:0] sel_242269;
  wire [7:0] add_242272;
  wire [7:0] sel_242273;
  wire [7:0] add_242276;
  wire [7:0] sel_242277;
  wire [7:0] add_242280;
  wire [7:0] sel_242281;
  wire [7:0] add_242284;
  wire [7:0] sel_242285;
  wire [7:0] add_242288;
  wire [7:0] sel_242289;
  wire [7:0] add_242292;
  wire [7:0] sel_242293;
  wire [7:0] add_242296;
  wire [7:0] sel_242297;
  wire [7:0] add_242300;
  wire [7:0] sel_242301;
  wire [7:0] add_242304;
  wire [7:0] sel_242305;
  wire [7:0] add_242308;
  wire [7:0] sel_242309;
  wire [7:0] add_242312;
  wire [7:0] sel_242313;
  wire [7:0] add_242316;
  wire [7:0] sel_242317;
  wire [7:0] add_242320;
  wire [7:0] sel_242321;
  wire [7:0] add_242324;
  wire [7:0] sel_242325;
  wire [7:0] add_242328;
  wire [7:0] sel_242329;
  wire [7:0] add_242332;
  wire [7:0] sel_242333;
  wire [7:0] add_242336;
  wire [7:0] sel_242337;
  wire [7:0] add_242340;
  wire [7:0] sel_242341;
  wire [7:0] add_242344;
  wire [7:0] sel_242345;
  wire [7:0] add_242348;
  wire [7:0] sel_242349;
  wire [7:0] add_242352;
  wire [7:0] sel_242353;
  wire [7:0] add_242356;
  wire [7:0] sel_242357;
  wire [7:0] add_242360;
  wire [7:0] sel_242361;
  wire [7:0] add_242364;
  wire [7:0] sel_242365;
  wire [7:0] add_242368;
  wire [7:0] sel_242369;
  wire [7:0] add_242372;
  wire [7:0] sel_242373;
  wire [7:0] add_242376;
  wire [7:0] sel_242377;
  wire [7:0] add_242380;
  wire [7:0] sel_242381;
  wire [7:0] add_242384;
  wire [7:0] sel_242385;
  wire [7:0] add_242388;
  wire [7:0] sel_242389;
  wire [7:0] add_242392;
  wire [7:0] sel_242393;
  wire [7:0] add_242396;
  wire [7:0] sel_242397;
  wire [7:0] add_242400;
  wire [7:0] sel_242401;
  wire [7:0] add_242404;
  wire [7:0] sel_242405;
  wire [7:0] add_242408;
  wire [7:0] sel_242409;
  wire [7:0] add_242412;
  wire [7:0] sel_242413;
  wire [7:0] add_242416;
  wire [7:0] sel_242417;
  wire [7:0] add_242420;
  wire [7:0] sel_242421;
  wire [7:0] add_242424;
  wire [7:0] sel_242425;
  wire [7:0] add_242428;
  wire [7:0] sel_242429;
  wire [7:0] add_242432;
  wire [7:0] sel_242433;
  wire [7:0] add_242436;
  wire [7:0] sel_242437;
  wire [7:0] add_242440;
  wire [7:0] sel_242441;
  wire [7:0] add_242444;
  wire [7:0] sel_242445;
  wire [7:0] add_242449;
  wire [15:0] array_index_242450;
  wire [7:0] sel_242451;
  wire [7:0] add_242454;
  wire [7:0] sel_242455;
  wire [7:0] add_242458;
  wire [7:0] sel_242459;
  wire [7:0] add_242462;
  wire [7:0] sel_242463;
  wire [7:0] add_242466;
  wire [7:0] sel_242467;
  wire [7:0] add_242470;
  wire [7:0] sel_242471;
  wire [7:0] add_242474;
  wire [7:0] sel_242475;
  wire [7:0] add_242478;
  wire [7:0] sel_242479;
  wire [7:0] add_242482;
  wire [7:0] sel_242483;
  wire [7:0] add_242486;
  wire [7:0] sel_242487;
  wire [7:0] add_242490;
  wire [7:0] sel_242491;
  wire [7:0] add_242494;
  wire [7:0] sel_242495;
  wire [7:0] add_242498;
  wire [7:0] sel_242499;
  wire [7:0] add_242502;
  wire [7:0] sel_242503;
  wire [7:0] add_242506;
  wire [7:0] sel_242507;
  wire [7:0] add_242510;
  wire [7:0] sel_242511;
  wire [7:0] add_242514;
  wire [7:0] sel_242515;
  wire [7:0] add_242518;
  wire [7:0] sel_242519;
  wire [7:0] add_242522;
  wire [7:0] sel_242523;
  wire [7:0] add_242526;
  wire [7:0] sel_242527;
  wire [7:0] add_242530;
  wire [7:0] sel_242531;
  wire [7:0] add_242534;
  wire [7:0] sel_242535;
  wire [7:0] add_242538;
  wire [7:0] sel_242539;
  wire [7:0] add_242542;
  wire [7:0] sel_242543;
  wire [7:0] add_242546;
  wire [7:0] sel_242547;
  wire [7:0] add_242550;
  wire [7:0] sel_242551;
  wire [7:0] add_242554;
  wire [7:0] sel_242555;
  wire [7:0] add_242558;
  wire [7:0] sel_242559;
  wire [7:0] add_242562;
  wire [7:0] sel_242563;
  wire [7:0] add_242566;
  wire [7:0] sel_242567;
  wire [7:0] add_242570;
  wire [7:0] sel_242571;
  wire [7:0] add_242574;
  wire [7:0] sel_242575;
  wire [7:0] add_242578;
  wire [7:0] sel_242579;
  wire [7:0] add_242582;
  wire [7:0] sel_242583;
  wire [7:0] add_242586;
  wire [7:0] sel_242587;
  wire [7:0] add_242590;
  wire [7:0] sel_242591;
  wire [7:0] add_242594;
  wire [7:0] sel_242595;
  wire [7:0] add_242598;
  wire [7:0] sel_242599;
  wire [7:0] add_242602;
  wire [7:0] sel_242603;
  wire [7:0] add_242606;
  wire [7:0] sel_242607;
  wire [7:0] add_242610;
  wire [7:0] sel_242611;
  wire [7:0] add_242614;
  wire [7:0] sel_242615;
  wire [7:0] add_242618;
  wire [7:0] sel_242619;
  wire [7:0] add_242622;
  wire [7:0] sel_242623;
  wire [7:0] add_242626;
  wire [7:0] sel_242627;
  wire [7:0] add_242630;
  wire [7:0] sel_242631;
  wire [7:0] add_242634;
  wire [7:0] sel_242635;
  wire [7:0] add_242638;
  wire [7:0] sel_242639;
  wire [7:0] add_242642;
  wire [7:0] sel_242643;
  wire [7:0] add_242646;
  wire [7:0] sel_242647;
  wire [7:0] add_242651;
  wire [15:0] array_index_242652;
  wire [7:0] sel_242653;
  wire [7:0] add_242656;
  wire [7:0] sel_242657;
  wire [7:0] add_242660;
  wire [7:0] sel_242661;
  wire [7:0] add_242664;
  wire [7:0] sel_242665;
  wire [7:0] add_242668;
  wire [7:0] sel_242669;
  wire [7:0] add_242672;
  wire [7:0] sel_242673;
  wire [7:0] add_242676;
  wire [7:0] sel_242677;
  wire [7:0] add_242680;
  wire [7:0] sel_242681;
  wire [7:0] add_242684;
  wire [7:0] sel_242685;
  wire [7:0] add_242688;
  wire [7:0] sel_242689;
  wire [7:0] add_242692;
  wire [7:0] sel_242693;
  wire [7:0] add_242696;
  wire [7:0] sel_242697;
  wire [7:0] add_242700;
  wire [7:0] sel_242701;
  wire [7:0] add_242704;
  wire [7:0] sel_242705;
  wire [7:0] add_242708;
  wire [7:0] sel_242709;
  wire [7:0] add_242712;
  wire [7:0] sel_242713;
  wire [7:0] add_242716;
  wire [7:0] sel_242717;
  wire [7:0] add_242720;
  wire [7:0] sel_242721;
  wire [7:0] add_242724;
  wire [7:0] sel_242725;
  wire [7:0] add_242728;
  wire [7:0] sel_242729;
  wire [7:0] add_242732;
  wire [7:0] sel_242733;
  wire [7:0] add_242736;
  wire [7:0] sel_242737;
  wire [7:0] add_242740;
  wire [7:0] sel_242741;
  wire [7:0] add_242744;
  wire [7:0] sel_242745;
  wire [7:0] add_242748;
  wire [7:0] sel_242749;
  wire [7:0] add_242752;
  wire [7:0] sel_242753;
  wire [7:0] add_242756;
  wire [7:0] sel_242757;
  wire [7:0] add_242760;
  wire [7:0] sel_242761;
  wire [7:0] add_242764;
  wire [7:0] sel_242765;
  wire [7:0] add_242768;
  wire [7:0] sel_242769;
  wire [7:0] add_242772;
  wire [7:0] sel_242773;
  wire [7:0] add_242776;
  wire [7:0] sel_242777;
  wire [7:0] add_242780;
  wire [7:0] sel_242781;
  wire [7:0] add_242784;
  wire [7:0] sel_242785;
  wire [7:0] add_242788;
  wire [7:0] sel_242789;
  wire [7:0] add_242792;
  wire [7:0] sel_242793;
  wire [7:0] add_242796;
  wire [7:0] sel_242797;
  wire [7:0] add_242800;
  wire [7:0] sel_242801;
  wire [7:0] add_242804;
  wire [7:0] sel_242805;
  wire [7:0] add_242808;
  wire [7:0] sel_242809;
  wire [7:0] add_242812;
  wire [7:0] sel_242813;
  wire [7:0] add_242816;
  wire [7:0] sel_242817;
  wire [7:0] add_242820;
  wire [7:0] sel_242821;
  wire [7:0] add_242824;
  wire [7:0] sel_242825;
  wire [7:0] add_242828;
  wire [7:0] sel_242829;
  wire [7:0] add_242832;
  wire [7:0] sel_242833;
  wire [7:0] add_242836;
  wire [7:0] sel_242837;
  wire [7:0] add_242840;
  wire [7:0] sel_242841;
  wire [7:0] add_242844;
  wire [7:0] sel_242845;
  wire [7:0] add_242848;
  wire [7:0] sel_242849;
  wire [7:0] add_242853;
  wire [15:0] array_index_242854;
  wire [7:0] sel_242855;
  wire [7:0] add_242858;
  wire [7:0] sel_242859;
  wire [7:0] add_242862;
  wire [7:0] sel_242863;
  wire [7:0] add_242866;
  wire [7:0] sel_242867;
  wire [7:0] add_242870;
  wire [7:0] sel_242871;
  wire [7:0] add_242874;
  wire [7:0] sel_242875;
  wire [7:0] add_242878;
  wire [7:0] sel_242879;
  wire [7:0] add_242882;
  wire [7:0] sel_242883;
  wire [7:0] add_242886;
  wire [7:0] sel_242887;
  wire [7:0] add_242890;
  wire [7:0] sel_242891;
  wire [7:0] add_242894;
  wire [7:0] sel_242895;
  wire [7:0] add_242898;
  wire [7:0] sel_242899;
  wire [7:0] add_242902;
  wire [7:0] sel_242903;
  wire [7:0] add_242906;
  wire [7:0] sel_242907;
  wire [7:0] add_242910;
  wire [7:0] sel_242911;
  wire [7:0] add_242914;
  wire [7:0] sel_242915;
  wire [7:0] add_242918;
  wire [7:0] sel_242919;
  wire [7:0] add_242922;
  wire [7:0] sel_242923;
  wire [7:0] add_242926;
  wire [7:0] sel_242927;
  wire [7:0] add_242930;
  wire [7:0] sel_242931;
  wire [7:0] add_242934;
  wire [7:0] sel_242935;
  wire [7:0] add_242938;
  wire [7:0] sel_242939;
  wire [7:0] add_242942;
  wire [7:0] sel_242943;
  wire [7:0] add_242946;
  wire [7:0] sel_242947;
  wire [7:0] add_242950;
  wire [7:0] sel_242951;
  wire [7:0] add_242954;
  wire [7:0] sel_242955;
  wire [7:0] add_242958;
  wire [7:0] sel_242959;
  wire [7:0] add_242962;
  wire [7:0] sel_242963;
  wire [7:0] add_242966;
  wire [7:0] sel_242967;
  wire [7:0] add_242970;
  wire [7:0] sel_242971;
  wire [7:0] add_242974;
  wire [7:0] sel_242975;
  wire [7:0] add_242978;
  wire [7:0] sel_242979;
  wire [7:0] add_242982;
  wire [7:0] sel_242983;
  wire [7:0] add_242986;
  wire [7:0] sel_242987;
  wire [7:0] add_242990;
  wire [7:0] sel_242991;
  wire [7:0] add_242994;
  wire [7:0] sel_242995;
  wire [7:0] add_242998;
  wire [7:0] sel_242999;
  wire [7:0] add_243002;
  wire [7:0] sel_243003;
  wire [7:0] add_243006;
  wire [7:0] sel_243007;
  wire [7:0] add_243010;
  wire [7:0] sel_243011;
  wire [7:0] add_243014;
  wire [7:0] sel_243015;
  wire [7:0] add_243018;
  wire [7:0] sel_243019;
  wire [7:0] add_243022;
  wire [7:0] sel_243023;
  wire [7:0] add_243026;
  wire [7:0] sel_243027;
  wire [7:0] add_243030;
  wire [7:0] sel_243031;
  wire [7:0] add_243034;
  wire [7:0] sel_243035;
  wire [7:0] add_243038;
  wire [7:0] sel_243039;
  wire [7:0] add_243042;
  wire [7:0] sel_243043;
  wire [7:0] add_243046;
  wire [7:0] sel_243047;
  wire [7:0] add_243050;
  wire [7:0] sel_243051;
  wire [7:0] add_243055;
  wire [15:0] array_index_243056;
  wire [7:0] sel_243057;
  wire [7:0] add_243060;
  wire [7:0] sel_243061;
  wire [7:0] add_243064;
  wire [7:0] sel_243065;
  wire [7:0] add_243068;
  wire [7:0] sel_243069;
  wire [7:0] add_243072;
  wire [7:0] sel_243073;
  wire [7:0] add_243076;
  wire [7:0] sel_243077;
  wire [7:0] add_243080;
  wire [7:0] sel_243081;
  wire [7:0] add_243084;
  wire [7:0] sel_243085;
  wire [7:0] add_243088;
  wire [7:0] sel_243089;
  wire [7:0] add_243092;
  wire [7:0] sel_243093;
  wire [7:0] add_243096;
  wire [7:0] sel_243097;
  wire [7:0] add_243100;
  wire [7:0] sel_243101;
  wire [7:0] add_243104;
  wire [7:0] sel_243105;
  wire [7:0] add_243108;
  wire [7:0] sel_243109;
  wire [7:0] add_243112;
  wire [7:0] sel_243113;
  wire [7:0] add_243116;
  wire [7:0] sel_243117;
  wire [7:0] add_243120;
  wire [7:0] sel_243121;
  wire [7:0] add_243124;
  wire [7:0] sel_243125;
  wire [7:0] add_243128;
  wire [7:0] sel_243129;
  wire [7:0] add_243132;
  wire [7:0] sel_243133;
  wire [7:0] add_243136;
  wire [7:0] sel_243137;
  wire [7:0] add_243140;
  wire [7:0] sel_243141;
  wire [7:0] add_243144;
  wire [7:0] sel_243145;
  wire [7:0] add_243148;
  wire [7:0] sel_243149;
  wire [7:0] add_243152;
  wire [7:0] sel_243153;
  wire [7:0] add_243156;
  wire [7:0] sel_243157;
  wire [7:0] add_243160;
  wire [7:0] sel_243161;
  wire [7:0] add_243164;
  wire [7:0] sel_243165;
  wire [7:0] add_243168;
  wire [7:0] sel_243169;
  wire [7:0] add_243172;
  wire [7:0] sel_243173;
  wire [7:0] add_243176;
  wire [7:0] sel_243177;
  wire [7:0] add_243180;
  wire [7:0] sel_243181;
  wire [7:0] add_243184;
  wire [7:0] sel_243185;
  wire [7:0] add_243188;
  wire [7:0] sel_243189;
  wire [7:0] add_243192;
  wire [7:0] sel_243193;
  wire [7:0] add_243196;
  wire [7:0] sel_243197;
  wire [7:0] add_243200;
  wire [7:0] sel_243201;
  wire [7:0] add_243204;
  wire [7:0] sel_243205;
  wire [7:0] add_243208;
  wire [7:0] sel_243209;
  wire [7:0] add_243212;
  wire [7:0] sel_243213;
  wire [7:0] add_243216;
  wire [7:0] sel_243217;
  wire [7:0] add_243220;
  wire [7:0] sel_243221;
  wire [7:0] add_243224;
  wire [7:0] sel_243225;
  wire [7:0] add_243228;
  wire [7:0] sel_243229;
  wire [7:0] add_243232;
  wire [7:0] sel_243233;
  wire [7:0] add_243236;
  wire [7:0] sel_243237;
  wire [7:0] add_243240;
  wire [7:0] sel_243241;
  wire [7:0] add_243244;
  wire [7:0] sel_243245;
  wire [7:0] add_243248;
  wire [7:0] sel_243249;
  wire [7:0] add_243252;
  wire [7:0] sel_243253;
  wire [7:0] add_243257;
  wire [15:0] array_index_243258;
  wire [7:0] sel_243259;
  wire [7:0] add_243262;
  wire [7:0] sel_243263;
  wire [7:0] add_243266;
  wire [7:0] sel_243267;
  wire [7:0] add_243270;
  wire [7:0] sel_243271;
  wire [7:0] add_243274;
  wire [7:0] sel_243275;
  wire [7:0] add_243278;
  wire [7:0] sel_243279;
  wire [7:0] add_243282;
  wire [7:0] sel_243283;
  wire [7:0] add_243286;
  wire [7:0] sel_243287;
  wire [7:0] add_243290;
  wire [7:0] sel_243291;
  wire [7:0] add_243294;
  wire [7:0] sel_243295;
  wire [7:0] add_243298;
  wire [7:0] sel_243299;
  wire [7:0] add_243302;
  wire [7:0] sel_243303;
  wire [7:0] add_243306;
  wire [7:0] sel_243307;
  wire [7:0] add_243310;
  wire [7:0] sel_243311;
  wire [7:0] add_243314;
  wire [7:0] sel_243315;
  wire [7:0] add_243318;
  wire [7:0] sel_243319;
  wire [7:0] add_243322;
  wire [7:0] sel_243323;
  wire [7:0] add_243326;
  wire [7:0] sel_243327;
  wire [7:0] add_243330;
  wire [7:0] sel_243331;
  wire [7:0] add_243334;
  wire [7:0] sel_243335;
  wire [7:0] add_243338;
  wire [7:0] sel_243339;
  wire [7:0] add_243342;
  wire [7:0] sel_243343;
  wire [7:0] add_243346;
  wire [7:0] sel_243347;
  wire [7:0] add_243350;
  wire [7:0] sel_243351;
  wire [7:0] add_243354;
  wire [7:0] sel_243355;
  wire [7:0] add_243358;
  wire [7:0] sel_243359;
  wire [7:0] add_243362;
  wire [7:0] sel_243363;
  wire [7:0] add_243366;
  wire [7:0] sel_243367;
  wire [7:0] add_243370;
  wire [7:0] sel_243371;
  wire [7:0] add_243374;
  wire [7:0] sel_243375;
  wire [7:0] add_243378;
  wire [7:0] sel_243379;
  wire [7:0] add_243382;
  wire [7:0] sel_243383;
  wire [7:0] add_243386;
  wire [7:0] sel_243387;
  wire [7:0] add_243390;
  wire [7:0] sel_243391;
  wire [7:0] add_243394;
  wire [7:0] sel_243395;
  wire [7:0] add_243398;
  wire [7:0] sel_243399;
  wire [7:0] add_243402;
  wire [7:0] sel_243403;
  wire [7:0] add_243406;
  wire [7:0] sel_243407;
  wire [7:0] add_243410;
  wire [7:0] sel_243411;
  wire [7:0] add_243414;
  wire [7:0] sel_243415;
  wire [7:0] add_243418;
  wire [7:0] sel_243419;
  wire [7:0] add_243422;
  wire [7:0] sel_243423;
  wire [7:0] add_243426;
  wire [7:0] sel_243427;
  wire [7:0] add_243430;
  wire [7:0] sel_243431;
  wire [7:0] add_243434;
  wire [7:0] sel_243435;
  wire [7:0] add_243438;
  wire [7:0] sel_243439;
  wire [7:0] add_243442;
  wire [7:0] sel_243443;
  wire [7:0] add_243446;
  wire [7:0] sel_243447;
  wire [7:0] add_243450;
  wire [7:0] sel_243451;
  wire [7:0] add_243454;
  wire [7:0] sel_243455;
  wire [7:0] add_243459;
  wire [15:0] array_index_243460;
  wire [7:0] sel_243461;
  wire [7:0] add_243464;
  wire [7:0] sel_243465;
  wire [7:0] add_243468;
  wire [7:0] sel_243469;
  wire [7:0] add_243472;
  wire [7:0] sel_243473;
  wire [7:0] add_243476;
  wire [7:0] sel_243477;
  wire [7:0] add_243480;
  wire [7:0] sel_243481;
  wire [7:0] add_243484;
  wire [7:0] sel_243485;
  wire [7:0] add_243488;
  wire [7:0] sel_243489;
  wire [7:0] add_243492;
  wire [7:0] sel_243493;
  wire [7:0] add_243496;
  wire [7:0] sel_243497;
  wire [7:0] add_243500;
  wire [7:0] sel_243501;
  wire [7:0] add_243504;
  wire [7:0] sel_243505;
  wire [7:0] add_243508;
  wire [7:0] sel_243509;
  wire [7:0] add_243512;
  wire [7:0] sel_243513;
  wire [7:0] add_243516;
  wire [7:0] sel_243517;
  wire [7:0] add_243520;
  wire [7:0] sel_243521;
  wire [7:0] add_243524;
  wire [7:0] sel_243525;
  wire [7:0] add_243528;
  wire [7:0] sel_243529;
  wire [7:0] add_243532;
  wire [7:0] sel_243533;
  wire [7:0] add_243536;
  wire [7:0] sel_243537;
  wire [7:0] add_243540;
  wire [7:0] sel_243541;
  wire [7:0] add_243544;
  wire [7:0] sel_243545;
  wire [7:0] add_243548;
  wire [7:0] sel_243549;
  wire [7:0] add_243552;
  wire [7:0] sel_243553;
  wire [7:0] add_243556;
  wire [7:0] sel_243557;
  wire [7:0] add_243560;
  wire [7:0] sel_243561;
  wire [7:0] add_243564;
  wire [7:0] sel_243565;
  wire [7:0] add_243568;
  wire [7:0] sel_243569;
  wire [7:0] add_243572;
  wire [7:0] sel_243573;
  wire [7:0] add_243576;
  wire [7:0] sel_243577;
  wire [7:0] add_243580;
  wire [7:0] sel_243581;
  wire [7:0] add_243584;
  wire [7:0] sel_243585;
  wire [7:0] add_243588;
  wire [7:0] sel_243589;
  wire [7:0] add_243592;
  wire [7:0] sel_243593;
  wire [7:0] add_243596;
  wire [7:0] sel_243597;
  wire [7:0] add_243600;
  wire [7:0] sel_243601;
  wire [7:0] add_243604;
  wire [7:0] sel_243605;
  wire [7:0] add_243608;
  wire [7:0] sel_243609;
  wire [7:0] add_243612;
  wire [7:0] sel_243613;
  wire [7:0] add_243616;
  wire [7:0] sel_243617;
  wire [7:0] add_243620;
  wire [7:0] sel_243621;
  wire [7:0] add_243624;
  wire [7:0] sel_243625;
  wire [7:0] add_243628;
  wire [7:0] sel_243629;
  wire [7:0] add_243632;
  wire [7:0] sel_243633;
  wire [7:0] add_243636;
  wire [7:0] sel_243637;
  wire [7:0] add_243640;
  wire [7:0] sel_243641;
  wire [7:0] add_243644;
  wire [7:0] sel_243645;
  wire [7:0] add_243648;
  wire [7:0] sel_243649;
  wire [7:0] add_243652;
  wire [7:0] sel_243653;
  wire [7:0] add_243656;
  wire [7:0] sel_243657;
  wire [7:0] add_243661;
  wire [15:0] array_index_243662;
  wire [7:0] sel_243663;
  wire [7:0] add_243666;
  wire [7:0] sel_243667;
  wire [7:0] add_243670;
  wire [7:0] sel_243671;
  wire [7:0] add_243674;
  wire [7:0] sel_243675;
  wire [7:0] add_243678;
  wire [7:0] sel_243679;
  wire [7:0] add_243682;
  wire [7:0] sel_243683;
  wire [7:0] add_243686;
  wire [7:0] sel_243687;
  wire [7:0] add_243690;
  wire [7:0] sel_243691;
  wire [7:0] add_243694;
  wire [7:0] sel_243695;
  wire [7:0] add_243698;
  wire [7:0] sel_243699;
  wire [7:0] add_243702;
  wire [7:0] sel_243703;
  wire [7:0] add_243706;
  wire [7:0] sel_243707;
  wire [7:0] add_243710;
  wire [7:0] sel_243711;
  wire [7:0] add_243714;
  wire [7:0] sel_243715;
  wire [7:0] add_243718;
  wire [7:0] sel_243719;
  wire [7:0] add_243722;
  wire [7:0] sel_243723;
  wire [7:0] add_243726;
  wire [7:0] sel_243727;
  wire [7:0] add_243730;
  wire [7:0] sel_243731;
  wire [7:0] add_243734;
  wire [7:0] sel_243735;
  wire [7:0] add_243738;
  wire [7:0] sel_243739;
  wire [7:0] add_243742;
  wire [7:0] sel_243743;
  wire [7:0] add_243746;
  wire [7:0] sel_243747;
  wire [7:0] add_243750;
  wire [7:0] sel_243751;
  wire [7:0] add_243754;
  wire [7:0] sel_243755;
  wire [7:0] add_243758;
  wire [7:0] sel_243759;
  wire [7:0] add_243762;
  wire [7:0] sel_243763;
  wire [7:0] add_243766;
  wire [7:0] sel_243767;
  wire [7:0] add_243770;
  wire [7:0] sel_243771;
  wire [7:0] add_243774;
  wire [7:0] sel_243775;
  wire [7:0] add_243778;
  wire [7:0] sel_243779;
  wire [7:0] add_243782;
  wire [7:0] sel_243783;
  wire [7:0] add_243786;
  wire [7:0] sel_243787;
  wire [7:0] add_243790;
  wire [7:0] sel_243791;
  wire [7:0] add_243794;
  wire [7:0] sel_243795;
  wire [7:0] add_243798;
  wire [7:0] sel_243799;
  wire [7:0] add_243802;
  wire [7:0] sel_243803;
  wire [7:0] add_243806;
  wire [7:0] sel_243807;
  wire [7:0] add_243810;
  wire [7:0] sel_243811;
  wire [7:0] add_243814;
  wire [7:0] sel_243815;
  wire [7:0] add_243818;
  wire [7:0] sel_243819;
  wire [7:0] add_243822;
  wire [7:0] sel_243823;
  wire [7:0] add_243826;
  wire [7:0] sel_243827;
  wire [7:0] add_243830;
  wire [7:0] sel_243831;
  wire [7:0] add_243834;
  wire [7:0] sel_243835;
  wire [7:0] add_243838;
  wire [7:0] sel_243839;
  wire [7:0] add_243842;
  wire [7:0] sel_243843;
  wire [7:0] add_243846;
  wire [7:0] sel_243847;
  wire [7:0] add_243850;
  wire [7:0] sel_243851;
  wire [7:0] add_243854;
  wire [7:0] sel_243855;
  wire [7:0] add_243858;
  wire [7:0] sel_243859;
  wire [7:0] add_243863;
  wire [15:0] array_index_243864;
  wire [7:0] sel_243865;
  wire [7:0] add_243868;
  wire [7:0] sel_243869;
  wire [7:0] add_243872;
  wire [7:0] sel_243873;
  wire [7:0] add_243876;
  wire [7:0] sel_243877;
  wire [7:0] add_243880;
  wire [7:0] sel_243881;
  wire [7:0] add_243884;
  wire [7:0] sel_243885;
  wire [7:0] add_243888;
  wire [7:0] sel_243889;
  wire [7:0] add_243892;
  wire [7:0] sel_243893;
  wire [7:0] add_243896;
  wire [7:0] sel_243897;
  wire [7:0] add_243900;
  wire [7:0] sel_243901;
  wire [7:0] add_243904;
  wire [7:0] sel_243905;
  wire [7:0] add_243908;
  wire [7:0] sel_243909;
  wire [7:0] add_243912;
  wire [7:0] sel_243913;
  wire [7:0] add_243916;
  wire [7:0] sel_243917;
  wire [7:0] add_243920;
  wire [7:0] sel_243921;
  wire [7:0] add_243924;
  wire [7:0] sel_243925;
  wire [7:0] add_243928;
  wire [7:0] sel_243929;
  wire [7:0] add_243932;
  wire [7:0] sel_243933;
  wire [7:0] add_243936;
  wire [7:0] sel_243937;
  wire [7:0] add_243940;
  wire [7:0] sel_243941;
  wire [7:0] add_243944;
  wire [7:0] sel_243945;
  wire [7:0] add_243948;
  wire [7:0] sel_243949;
  wire [7:0] add_243952;
  wire [7:0] sel_243953;
  wire [7:0] add_243956;
  wire [7:0] sel_243957;
  wire [7:0] add_243960;
  wire [7:0] sel_243961;
  wire [7:0] add_243964;
  wire [7:0] sel_243965;
  wire [7:0] add_243968;
  wire [7:0] sel_243969;
  wire [7:0] add_243972;
  wire [7:0] sel_243973;
  wire [7:0] add_243976;
  wire [7:0] sel_243977;
  wire [7:0] add_243980;
  wire [7:0] sel_243981;
  wire [7:0] add_243984;
  wire [7:0] sel_243985;
  wire [7:0] add_243988;
  wire [7:0] sel_243989;
  wire [7:0] add_243992;
  wire [7:0] sel_243993;
  wire [7:0] add_243996;
  wire [7:0] sel_243997;
  wire [7:0] add_244000;
  wire [7:0] sel_244001;
  wire [7:0] add_244004;
  wire [7:0] sel_244005;
  wire [7:0] add_244008;
  wire [7:0] sel_244009;
  wire [7:0] add_244012;
  wire [7:0] sel_244013;
  wire [7:0] add_244016;
  wire [7:0] sel_244017;
  wire [7:0] add_244020;
  wire [7:0] sel_244021;
  wire [7:0] add_244024;
  wire [7:0] sel_244025;
  wire [7:0] add_244028;
  wire [7:0] sel_244029;
  wire [7:0] add_244032;
  wire [7:0] sel_244033;
  wire [7:0] add_244036;
  wire [7:0] sel_244037;
  wire [7:0] add_244040;
  wire [7:0] sel_244041;
  wire [7:0] add_244044;
  wire [7:0] sel_244045;
  wire [7:0] add_244048;
  wire [7:0] sel_244049;
  wire [7:0] add_244052;
  wire [7:0] sel_244053;
  wire [7:0] add_244056;
  wire [7:0] sel_244057;
  wire [7:0] add_244060;
  wire [7:0] sel_244061;
  wire [7:0] add_244065;
  wire [15:0] array_index_244066;
  wire [7:0] sel_244067;
  wire [7:0] add_244070;
  wire [7:0] sel_244071;
  wire [7:0] add_244074;
  wire [7:0] sel_244075;
  wire [7:0] add_244078;
  wire [7:0] sel_244079;
  wire [7:0] add_244082;
  wire [7:0] sel_244083;
  wire [7:0] add_244086;
  wire [7:0] sel_244087;
  wire [7:0] add_244090;
  wire [7:0] sel_244091;
  wire [7:0] add_244094;
  wire [7:0] sel_244095;
  wire [7:0] add_244098;
  wire [7:0] sel_244099;
  wire [7:0] add_244102;
  wire [7:0] sel_244103;
  wire [7:0] add_244106;
  wire [7:0] sel_244107;
  wire [7:0] add_244110;
  wire [7:0] sel_244111;
  wire [7:0] add_244114;
  wire [7:0] sel_244115;
  wire [7:0] add_244118;
  wire [7:0] sel_244119;
  wire [7:0] add_244122;
  wire [7:0] sel_244123;
  wire [7:0] add_244126;
  wire [7:0] sel_244127;
  wire [7:0] add_244130;
  wire [7:0] sel_244131;
  wire [7:0] add_244134;
  wire [7:0] sel_244135;
  wire [7:0] add_244138;
  wire [7:0] sel_244139;
  wire [7:0] add_244142;
  wire [7:0] sel_244143;
  wire [7:0] add_244146;
  wire [7:0] sel_244147;
  wire [7:0] add_244150;
  wire [7:0] sel_244151;
  wire [7:0] add_244154;
  wire [7:0] sel_244155;
  wire [7:0] add_244158;
  wire [7:0] sel_244159;
  wire [7:0] add_244162;
  wire [7:0] sel_244163;
  wire [7:0] add_244166;
  wire [7:0] sel_244167;
  wire [7:0] add_244170;
  wire [7:0] sel_244171;
  wire [7:0] add_244174;
  wire [7:0] sel_244175;
  wire [7:0] add_244178;
  wire [7:0] sel_244179;
  wire [7:0] add_244182;
  wire [7:0] sel_244183;
  wire [7:0] add_244186;
  wire [7:0] sel_244187;
  wire [7:0] add_244190;
  wire [7:0] sel_244191;
  wire [7:0] add_244194;
  wire [7:0] sel_244195;
  wire [7:0] add_244198;
  wire [7:0] sel_244199;
  wire [7:0] add_244202;
  wire [7:0] sel_244203;
  wire [7:0] add_244206;
  wire [7:0] sel_244207;
  wire [7:0] add_244210;
  wire [7:0] sel_244211;
  wire [7:0] add_244214;
  wire [7:0] sel_244215;
  wire [7:0] add_244218;
  wire [7:0] sel_244219;
  wire [7:0] add_244222;
  wire [7:0] sel_244223;
  wire [7:0] add_244226;
  wire [7:0] sel_244227;
  wire [7:0] add_244230;
  wire [7:0] sel_244231;
  wire [7:0] add_244234;
  wire [7:0] sel_244235;
  wire [7:0] add_244238;
  wire [7:0] sel_244239;
  wire [7:0] add_244242;
  wire [7:0] sel_244243;
  wire [7:0] add_244246;
  wire [7:0] sel_244247;
  wire [7:0] add_244250;
  wire [7:0] sel_244251;
  wire [7:0] add_244254;
  wire [7:0] sel_244255;
  wire [7:0] add_244258;
  wire [7:0] sel_244259;
  wire [7:0] add_244262;
  wire [7:0] sel_244263;
  wire [7:0] add_244267;
  wire [15:0] array_index_244268;
  wire [7:0] sel_244269;
  wire [7:0] add_244272;
  wire [7:0] sel_244273;
  wire [7:0] add_244276;
  wire [7:0] sel_244277;
  wire [7:0] add_244280;
  wire [7:0] sel_244281;
  wire [7:0] add_244284;
  wire [7:0] sel_244285;
  wire [7:0] add_244288;
  wire [7:0] sel_244289;
  wire [7:0] add_244292;
  wire [7:0] sel_244293;
  wire [7:0] add_244296;
  wire [7:0] sel_244297;
  wire [7:0] add_244300;
  wire [7:0] sel_244301;
  wire [7:0] add_244304;
  wire [7:0] sel_244305;
  wire [7:0] add_244308;
  wire [7:0] sel_244309;
  wire [7:0] add_244312;
  wire [7:0] sel_244313;
  wire [7:0] add_244316;
  wire [7:0] sel_244317;
  wire [7:0] add_244320;
  wire [7:0] sel_244321;
  wire [7:0] add_244324;
  wire [7:0] sel_244325;
  wire [7:0] add_244328;
  wire [7:0] sel_244329;
  wire [7:0] add_244332;
  wire [7:0] sel_244333;
  wire [7:0] add_244336;
  wire [7:0] sel_244337;
  wire [7:0] add_244340;
  wire [7:0] sel_244341;
  wire [7:0] add_244344;
  wire [7:0] sel_244345;
  wire [7:0] add_244348;
  wire [7:0] sel_244349;
  wire [7:0] add_244352;
  wire [7:0] sel_244353;
  wire [7:0] add_244356;
  wire [7:0] sel_244357;
  wire [7:0] add_244360;
  wire [7:0] sel_244361;
  wire [7:0] add_244364;
  wire [7:0] sel_244365;
  wire [7:0] add_244368;
  wire [7:0] sel_244369;
  wire [7:0] add_244372;
  wire [7:0] sel_244373;
  wire [7:0] add_244376;
  wire [7:0] sel_244377;
  wire [7:0] add_244380;
  wire [7:0] sel_244381;
  wire [7:0] add_244384;
  wire [7:0] sel_244385;
  wire [7:0] add_244388;
  wire [7:0] sel_244389;
  wire [7:0] add_244392;
  wire [7:0] sel_244393;
  wire [7:0] add_244396;
  wire [7:0] sel_244397;
  wire [7:0] add_244400;
  wire [7:0] sel_244401;
  wire [7:0] add_244404;
  wire [7:0] sel_244405;
  wire [7:0] add_244408;
  wire [7:0] sel_244409;
  wire [7:0] add_244412;
  wire [7:0] sel_244413;
  wire [7:0] add_244416;
  wire [7:0] sel_244417;
  wire [7:0] add_244420;
  wire [7:0] sel_244421;
  wire [7:0] add_244424;
  wire [7:0] sel_244425;
  wire [7:0] add_244428;
  wire [7:0] sel_244429;
  wire [7:0] add_244432;
  wire [7:0] sel_244433;
  wire [7:0] add_244436;
  wire [7:0] sel_244437;
  wire [7:0] add_244440;
  wire [7:0] sel_244441;
  wire [7:0] add_244444;
  wire [7:0] sel_244445;
  wire [7:0] add_244448;
  wire [7:0] sel_244449;
  wire [7:0] add_244452;
  wire [7:0] sel_244453;
  wire [7:0] add_244456;
  wire [7:0] sel_244457;
  wire [7:0] add_244460;
  wire [7:0] sel_244461;
  wire [7:0] add_244464;
  wire [7:0] sel_244465;
  wire [7:0] add_244469;
  wire [15:0] array_index_244470;
  wire [7:0] sel_244471;
  wire [7:0] add_244474;
  wire [7:0] sel_244475;
  wire [7:0] add_244478;
  wire [7:0] sel_244479;
  wire [7:0] add_244482;
  wire [7:0] sel_244483;
  wire [7:0] add_244486;
  wire [7:0] sel_244487;
  wire [7:0] add_244490;
  wire [7:0] sel_244491;
  wire [7:0] add_244494;
  wire [7:0] sel_244495;
  wire [7:0] add_244498;
  wire [7:0] sel_244499;
  wire [7:0] add_244502;
  wire [7:0] sel_244503;
  wire [7:0] add_244506;
  wire [7:0] sel_244507;
  wire [7:0] add_244510;
  wire [7:0] sel_244511;
  wire [7:0] add_244514;
  wire [7:0] sel_244515;
  wire [7:0] add_244518;
  wire [7:0] sel_244519;
  wire [7:0] add_244522;
  wire [7:0] sel_244523;
  wire [7:0] add_244526;
  wire [7:0] sel_244527;
  wire [7:0] add_244530;
  wire [7:0] sel_244531;
  wire [7:0] add_244534;
  wire [7:0] sel_244535;
  wire [7:0] add_244538;
  wire [7:0] sel_244539;
  wire [7:0] add_244542;
  wire [7:0] sel_244543;
  wire [7:0] add_244546;
  wire [7:0] sel_244547;
  wire [7:0] add_244550;
  wire [7:0] sel_244551;
  wire [7:0] add_244554;
  wire [7:0] sel_244555;
  wire [7:0] add_244558;
  wire [7:0] sel_244559;
  wire [7:0] add_244562;
  wire [7:0] sel_244563;
  wire [7:0] add_244566;
  wire [7:0] sel_244567;
  wire [7:0] add_244570;
  wire [7:0] sel_244571;
  wire [7:0] add_244574;
  wire [7:0] sel_244575;
  wire [7:0] add_244578;
  wire [7:0] sel_244579;
  wire [7:0] add_244582;
  wire [7:0] sel_244583;
  wire [7:0] add_244586;
  wire [7:0] sel_244587;
  wire [7:0] add_244590;
  wire [7:0] sel_244591;
  wire [7:0] add_244594;
  wire [7:0] sel_244595;
  wire [7:0] add_244598;
  wire [7:0] sel_244599;
  wire [7:0] add_244602;
  wire [7:0] sel_244603;
  wire [7:0] add_244606;
  wire [7:0] sel_244607;
  wire [7:0] add_244610;
  wire [7:0] sel_244611;
  wire [7:0] add_244614;
  wire [7:0] sel_244615;
  wire [7:0] add_244618;
  wire [7:0] sel_244619;
  wire [7:0] add_244622;
  wire [7:0] sel_244623;
  wire [7:0] add_244626;
  wire [7:0] sel_244627;
  wire [7:0] add_244630;
  wire [7:0] sel_244631;
  wire [7:0] add_244634;
  wire [7:0] sel_244635;
  wire [7:0] add_244638;
  wire [7:0] sel_244639;
  wire [7:0] add_244642;
  wire [7:0] sel_244643;
  wire [7:0] add_244646;
  wire [7:0] sel_244647;
  wire [7:0] add_244650;
  wire [7:0] sel_244651;
  wire [7:0] add_244654;
  wire [7:0] sel_244655;
  wire [7:0] add_244658;
  wire [7:0] sel_244659;
  wire [7:0] add_244662;
  wire [7:0] sel_244663;
  wire [7:0] add_244666;
  wire [7:0] sel_244667;
  wire [7:0] add_244671;
  wire [15:0] array_index_244672;
  wire [7:0] sel_244673;
  wire [7:0] add_244676;
  wire [7:0] sel_244677;
  wire [7:0] add_244680;
  wire [7:0] sel_244681;
  wire [7:0] add_244684;
  wire [7:0] sel_244685;
  wire [7:0] add_244688;
  wire [7:0] sel_244689;
  wire [7:0] add_244692;
  wire [7:0] sel_244693;
  wire [7:0] add_244696;
  wire [7:0] sel_244697;
  wire [7:0] add_244700;
  wire [7:0] sel_244701;
  wire [7:0] add_244704;
  wire [7:0] sel_244705;
  wire [7:0] add_244708;
  wire [7:0] sel_244709;
  wire [7:0] add_244712;
  wire [7:0] sel_244713;
  wire [7:0] add_244716;
  wire [7:0] sel_244717;
  wire [7:0] add_244720;
  wire [7:0] sel_244721;
  wire [7:0] add_244724;
  wire [7:0] sel_244725;
  wire [7:0] add_244728;
  wire [7:0] sel_244729;
  wire [7:0] add_244732;
  wire [7:0] sel_244733;
  wire [7:0] add_244736;
  wire [7:0] sel_244737;
  wire [7:0] add_244740;
  wire [7:0] sel_244741;
  wire [7:0] add_244744;
  wire [7:0] sel_244745;
  wire [7:0] add_244748;
  wire [7:0] sel_244749;
  wire [7:0] add_244752;
  wire [7:0] sel_244753;
  wire [7:0] add_244756;
  wire [7:0] sel_244757;
  wire [7:0] add_244760;
  wire [7:0] sel_244761;
  wire [7:0] add_244764;
  wire [7:0] sel_244765;
  wire [7:0] add_244768;
  wire [7:0] sel_244769;
  wire [7:0] add_244772;
  wire [7:0] sel_244773;
  wire [7:0] add_244776;
  wire [7:0] sel_244777;
  wire [7:0] add_244780;
  wire [7:0] sel_244781;
  wire [7:0] add_244784;
  wire [7:0] sel_244785;
  wire [7:0] add_244788;
  wire [7:0] sel_244789;
  wire [7:0] add_244792;
  wire [7:0] sel_244793;
  wire [7:0] add_244796;
  wire [7:0] sel_244797;
  wire [7:0] add_244800;
  wire [7:0] sel_244801;
  wire [7:0] add_244804;
  wire [7:0] sel_244805;
  wire [7:0] add_244808;
  wire [7:0] sel_244809;
  wire [7:0] add_244812;
  wire [7:0] sel_244813;
  wire [7:0] add_244816;
  wire [7:0] sel_244817;
  wire [7:0] add_244820;
  wire [7:0] sel_244821;
  wire [7:0] add_244824;
  wire [7:0] sel_244825;
  wire [7:0] add_244828;
  wire [7:0] sel_244829;
  wire [7:0] add_244832;
  wire [7:0] sel_244833;
  wire [7:0] add_244836;
  wire [7:0] sel_244837;
  wire [7:0] add_244840;
  wire [7:0] sel_244841;
  wire [7:0] add_244844;
  wire [7:0] sel_244845;
  wire [7:0] add_244848;
  wire [7:0] sel_244849;
  wire [7:0] add_244852;
  wire [7:0] sel_244853;
  wire [7:0] add_244856;
  wire [7:0] sel_244857;
  wire [7:0] add_244860;
  wire [7:0] sel_244861;
  wire [7:0] add_244864;
  wire [7:0] sel_244865;
  wire [7:0] add_244868;
  wire [7:0] sel_244869;
  wire [7:0] add_244873;
  wire [15:0] array_index_244874;
  wire [7:0] sel_244875;
  wire [7:0] add_244878;
  wire [7:0] sel_244879;
  wire [7:0] add_244882;
  wire [7:0] sel_244883;
  wire [7:0] add_244886;
  wire [7:0] sel_244887;
  wire [7:0] add_244890;
  wire [7:0] sel_244891;
  wire [7:0] add_244894;
  wire [7:0] sel_244895;
  wire [7:0] add_244898;
  wire [7:0] sel_244899;
  wire [7:0] add_244902;
  wire [7:0] sel_244903;
  wire [7:0] add_244906;
  wire [7:0] sel_244907;
  wire [7:0] add_244910;
  wire [7:0] sel_244911;
  wire [7:0] add_244914;
  wire [7:0] sel_244915;
  wire [7:0] add_244918;
  wire [7:0] sel_244919;
  wire [7:0] add_244922;
  wire [7:0] sel_244923;
  wire [7:0] add_244926;
  wire [7:0] sel_244927;
  wire [7:0] add_244930;
  wire [7:0] sel_244931;
  wire [7:0] add_244934;
  wire [7:0] sel_244935;
  wire [7:0] add_244938;
  wire [7:0] sel_244939;
  wire [7:0] add_244942;
  wire [7:0] sel_244943;
  wire [7:0] add_244946;
  wire [7:0] sel_244947;
  wire [7:0] add_244950;
  wire [7:0] sel_244951;
  wire [7:0] add_244954;
  wire [7:0] sel_244955;
  wire [7:0] add_244958;
  wire [7:0] sel_244959;
  wire [7:0] add_244962;
  wire [7:0] sel_244963;
  wire [7:0] add_244966;
  wire [7:0] sel_244967;
  wire [7:0] add_244970;
  wire [7:0] sel_244971;
  wire [7:0] add_244974;
  wire [7:0] sel_244975;
  wire [7:0] add_244978;
  wire [7:0] sel_244979;
  wire [7:0] add_244982;
  wire [7:0] sel_244983;
  wire [7:0] add_244986;
  wire [7:0] sel_244987;
  wire [7:0] add_244990;
  wire [7:0] sel_244991;
  wire [7:0] add_244994;
  wire [7:0] sel_244995;
  wire [7:0] add_244998;
  wire [7:0] sel_244999;
  wire [7:0] add_245002;
  wire [7:0] sel_245003;
  wire [7:0] add_245006;
  wire [7:0] sel_245007;
  wire [7:0] add_245010;
  wire [7:0] sel_245011;
  wire [7:0] add_245014;
  wire [7:0] sel_245015;
  wire [7:0] add_245018;
  wire [7:0] sel_245019;
  wire [7:0] add_245022;
  wire [7:0] sel_245023;
  wire [7:0] add_245026;
  wire [7:0] sel_245027;
  wire [7:0] add_245030;
  wire [7:0] sel_245031;
  wire [7:0] add_245034;
  wire [7:0] sel_245035;
  wire [7:0] add_245038;
  wire [7:0] sel_245039;
  wire [7:0] add_245042;
  wire [7:0] sel_245043;
  wire [7:0] add_245046;
  wire [7:0] sel_245047;
  wire [7:0] add_245050;
  wire [7:0] sel_245051;
  wire [7:0] add_245054;
  wire [7:0] sel_245055;
  wire [7:0] add_245058;
  wire [7:0] sel_245059;
  wire [7:0] add_245062;
  wire [7:0] sel_245063;
  wire [7:0] add_245066;
  wire [7:0] sel_245067;
  wire [7:0] add_245070;
  wire [7:0] sel_245071;
  wire [7:0] add_245075;
  wire [15:0] array_index_245076;
  wire [7:0] sel_245077;
  wire [7:0] add_245080;
  wire [7:0] sel_245081;
  wire [7:0] add_245084;
  wire [7:0] sel_245085;
  wire [7:0] add_245088;
  wire [7:0] sel_245089;
  wire [7:0] add_245092;
  wire [7:0] sel_245093;
  wire [7:0] add_245096;
  wire [7:0] sel_245097;
  wire [7:0] add_245100;
  wire [7:0] sel_245101;
  wire [7:0] add_245104;
  wire [7:0] sel_245105;
  wire [7:0] add_245108;
  wire [7:0] sel_245109;
  wire [7:0] add_245112;
  wire [7:0] sel_245113;
  wire [7:0] add_245116;
  wire [7:0] sel_245117;
  wire [7:0] add_245120;
  wire [7:0] sel_245121;
  wire [7:0] add_245124;
  wire [7:0] sel_245125;
  wire [7:0] add_245128;
  wire [7:0] sel_245129;
  wire [7:0] add_245132;
  wire [7:0] sel_245133;
  wire [7:0] add_245136;
  wire [7:0] sel_245137;
  wire [7:0] add_245140;
  wire [7:0] sel_245141;
  wire [7:0] add_245144;
  wire [7:0] sel_245145;
  wire [7:0] add_245148;
  wire [7:0] sel_245149;
  wire [7:0] add_245152;
  wire [7:0] sel_245153;
  wire [7:0] add_245156;
  wire [7:0] sel_245157;
  wire [7:0] add_245160;
  wire [7:0] sel_245161;
  wire [7:0] add_245164;
  wire [7:0] sel_245165;
  wire [7:0] add_245168;
  wire [7:0] sel_245169;
  wire [7:0] add_245172;
  wire [7:0] sel_245173;
  wire [7:0] add_245176;
  wire [7:0] sel_245177;
  wire [7:0] add_245180;
  wire [7:0] sel_245181;
  wire [7:0] add_245184;
  wire [7:0] sel_245185;
  wire [7:0] add_245188;
  wire [7:0] sel_245189;
  wire [7:0] add_245192;
  wire [7:0] sel_245193;
  wire [7:0] add_245196;
  wire [7:0] sel_245197;
  wire [7:0] add_245200;
  wire [7:0] sel_245201;
  wire [7:0] add_245204;
  wire [7:0] sel_245205;
  wire [7:0] add_245208;
  wire [7:0] sel_245209;
  wire [7:0] add_245212;
  wire [7:0] sel_245213;
  wire [7:0] add_245216;
  wire [7:0] sel_245217;
  wire [7:0] add_245220;
  wire [7:0] sel_245221;
  wire [7:0] add_245224;
  wire [7:0] sel_245225;
  wire [7:0] add_245228;
  wire [7:0] sel_245229;
  wire [7:0] add_245232;
  wire [7:0] sel_245233;
  wire [7:0] add_245236;
  wire [7:0] sel_245237;
  wire [7:0] add_245240;
  wire [7:0] sel_245241;
  wire [7:0] add_245244;
  wire [7:0] sel_245245;
  wire [7:0] add_245248;
  wire [7:0] sel_245249;
  wire [7:0] add_245252;
  wire [7:0] sel_245253;
  wire [7:0] add_245256;
  wire [7:0] sel_245257;
  wire [7:0] add_245260;
  wire [7:0] sel_245261;
  wire [7:0] add_245264;
  wire [7:0] sel_245265;
  wire [7:0] add_245268;
  wire [7:0] sel_245269;
  wire [7:0] add_245272;
  wire [7:0] sel_245273;
  wire [7:0] add_245277;
  wire [15:0] array_index_245278;
  wire [7:0] sel_245279;
  wire [7:0] add_245282;
  wire [7:0] sel_245283;
  wire [7:0] add_245286;
  wire [7:0] sel_245287;
  wire [7:0] add_245290;
  wire [7:0] sel_245291;
  wire [7:0] add_245294;
  wire [7:0] sel_245295;
  wire [7:0] add_245298;
  wire [7:0] sel_245299;
  wire [7:0] add_245302;
  wire [7:0] sel_245303;
  wire [7:0] add_245306;
  wire [7:0] sel_245307;
  wire [7:0] add_245310;
  wire [7:0] sel_245311;
  wire [7:0] add_245314;
  wire [7:0] sel_245315;
  wire [7:0] add_245318;
  wire [7:0] sel_245319;
  wire [7:0] add_245322;
  wire [7:0] sel_245323;
  wire [7:0] add_245326;
  wire [7:0] sel_245327;
  wire [7:0] add_245330;
  wire [7:0] sel_245331;
  wire [7:0] add_245334;
  wire [7:0] sel_245335;
  wire [7:0] add_245338;
  wire [7:0] sel_245339;
  wire [7:0] add_245342;
  wire [7:0] sel_245343;
  wire [7:0] add_245346;
  wire [7:0] sel_245347;
  wire [7:0] add_245350;
  wire [7:0] sel_245351;
  wire [7:0] add_245354;
  wire [7:0] sel_245355;
  wire [7:0] add_245358;
  wire [7:0] sel_245359;
  wire [7:0] add_245362;
  wire [7:0] sel_245363;
  wire [7:0] add_245366;
  wire [7:0] sel_245367;
  wire [7:0] add_245370;
  wire [7:0] sel_245371;
  wire [7:0] add_245374;
  wire [7:0] sel_245375;
  wire [7:0] add_245378;
  wire [7:0] sel_245379;
  wire [7:0] add_245382;
  wire [7:0] sel_245383;
  wire [7:0] add_245386;
  wire [7:0] sel_245387;
  wire [7:0] add_245390;
  wire [7:0] sel_245391;
  wire [7:0] add_245394;
  wire [7:0] sel_245395;
  wire [7:0] add_245398;
  wire [7:0] sel_245399;
  wire [7:0] add_245402;
  wire [7:0] sel_245403;
  wire [7:0] add_245406;
  wire [7:0] sel_245407;
  wire [7:0] add_245410;
  wire [7:0] sel_245411;
  wire [7:0] add_245414;
  wire [7:0] sel_245415;
  wire [7:0] add_245418;
  wire [7:0] sel_245419;
  wire [7:0] add_245422;
  wire [7:0] sel_245423;
  wire [7:0] add_245426;
  wire [7:0] sel_245427;
  wire [7:0] add_245430;
  wire [7:0] sel_245431;
  wire [7:0] add_245434;
  wire [7:0] sel_245435;
  wire [7:0] add_245438;
  wire [7:0] sel_245439;
  wire [7:0] add_245442;
  wire [7:0] sel_245443;
  wire [7:0] add_245446;
  wire [7:0] sel_245447;
  wire [7:0] add_245450;
  wire [7:0] sel_245451;
  wire [7:0] add_245454;
  wire [7:0] sel_245455;
  wire [7:0] add_245458;
  wire [7:0] sel_245459;
  wire [7:0] add_245462;
  wire [7:0] sel_245463;
  wire [7:0] add_245466;
  wire [7:0] sel_245467;
  wire [7:0] add_245470;
  wire [7:0] sel_245471;
  wire [7:0] add_245474;
  wire [7:0] sel_245475;
  wire [7:0] add_245479;
  wire [15:0] array_index_245480;
  wire [7:0] sel_245481;
  wire [7:0] add_245484;
  wire [7:0] sel_245485;
  wire [7:0] add_245488;
  wire [7:0] sel_245489;
  wire [7:0] add_245492;
  wire [7:0] sel_245493;
  wire [7:0] add_245496;
  wire [7:0] sel_245497;
  wire [7:0] add_245500;
  wire [7:0] sel_245501;
  wire [7:0] add_245504;
  wire [7:0] sel_245505;
  wire [7:0] add_245508;
  wire [7:0] sel_245509;
  wire [7:0] add_245512;
  wire [7:0] sel_245513;
  wire [7:0] add_245516;
  wire [7:0] sel_245517;
  wire [7:0] add_245520;
  wire [7:0] sel_245521;
  wire [7:0] add_245524;
  wire [7:0] sel_245525;
  wire [7:0] add_245528;
  wire [7:0] sel_245529;
  wire [7:0] add_245532;
  wire [7:0] sel_245533;
  wire [7:0] add_245536;
  wire [7:0] sel_245537;
  wire [7:0] add_245540;
  wire [7:0] sel_245541;
  wire [7:0] add_245544;
  wire [7:0] sel_245545;
  wire [7:0] add_245548;
  wire [7:0] sel_245549;
  wire [7:0] add_245552;
  wire [7:0] sel_245553;
  wire [7:0] add_245556;
  wire [7:0] sel_245557;
  wire [7:0] add_245560;
  wire [7:0] sel_245561;
  wire [7:0] add_245564;
  wire [7:0] sel_245565;
  wire [7:0] add_245568;
  wire [7:0] sel_245569;
  wire [7:0] add_245572;
  wire [7:0] sel_245573;
  wire [7:0] add_245576;
  wire [7:0] sel_245577;
  wire [7:0] add_245580;
  wire [7:0] sel_245581;
  wire [7:0] add_245584;
  wire [7:0] sel_245585;
  wire [7:0] add_245588;
  wire [7:0] sel_245589;
  wire [7:0] add_245592;
  wire [7:0] sel_245593;
  wire [7:0] add_245596;
  wire [7:0] sel_245597;
  wire [7:0] add_245600;
  wire [7:0] sel_245601;
  wire [7:0] add_245604;
  wire [7:0] sel_245605;
  wire [7:0] add_245608;
  wire [7:0] sel_245609;
  wire [7:0] add_245612;
  wire [7:0] sel_245613;
  wire [7:0] add_245616;
  wire [7:0] sel_245617;
  wire [7:0] add_245620;
  wire [7:0] sel_245621;
  wire [7:0] add_245624;
  wire [7:0] sel_245625;
  wire [7:0] add_245628;
  wire [7:0] sel_245629;
  wire [7:0] add_245632;
  wire [7:0] sel_245633;
  wire [7:0] add_245636;
  wire [7:0] sel_245637;
  wire [7:0] add_245640;
  wire [7:0] sel_245641;
  wire [7:0] add_245644;
  wire [7:0] sel_245645;
  wire [7:0] add_245648;
  wire [7:0] sel_245649;
  wire [7:0] add_245652;
  wire [7:0] sel_245653;
  wire [7:0] add_245656;
  wire [7:0] sel_245657;
  wire [7:0] add_245660;
  wire [7:0] sel_245661;
  wire [7:0] add_245664;
  wire [7:0] sel_245665;
  wire [7:0] add_245668;
  wire [7:0] sel_245669;
  wire [7:0] add_245672;
  wire [7:0] sel_245673;
  wire [7:0] add_245676;
  wire [7:0] sel_245677;
  wire [7:0] add_245681;
  wire [15:0] array_index_245682;
  wire [7:0] sel_245683;
  wire [7:0] add_245686;
  wire [7:0] sel_245687;
  wire [7:0] add_245690;
  wire [7:0] sel_245691;
  wire [7:0] add_245694;
  wire [7:0] sel_245695;
  wire [7:0] add_245698;
  wire [7:0] sel_245699;
  wire [7:0] add_245702;
  wire [7:0] sel_245703;
  wire [7:0] add_245706;
  wire [7:0] sel_245707;
  wire [7:0] add_245710;
  wire [7:0] sel_245711;
  wire [7:0] add_245714;
  wire [7:0] sel_245715;
  wire [7:0] add_245718;
  wire [7:0] sel_245719;
  wire [7:0] add_245722;
  wire [7:0] sel_245723;
  wire [7:0] add_245726;
  wire [7:0] sel_245727;
  wire [7:0] add_245730;
  wire [7:0] sel_245731;
  wire [7:0] add_245734;
  wire [7:0] sel_245735;
  wire [7:0] add_245738;
  wire [7:0] sel_245739;
  wire [7:0] add_245742;
  wire [7:0] sel_245743;
  wire [7:0] add_245746;
  wire [7:0] sel_245747;
  wire [7:0] add_245750;
  wire [7:0] sel_245751;
  wire [7:0] add_245754;
  wire [7:0] sel_245755;
  wire [7:0] add_245758;
  wire [7:0] sel_245759;
  wire [7:0] add_245762;
  wire [7:0] sel_245763;
  wire [7:0] add_245766;
  wire [7:0] sel_245767;
  wire [7:0] add_245770;
  wire [7:0] sel_245771;
  wire [7:0] add_245774;
  wire [7:0] sel_245775;
  wire [7:0] add_245778;
  wire [7:0] sel_245779;
  wire [7:0] add_245782;
  wire [7:0] sel_245783;
  wire [7:0] add_245786;
  wire [7:0] sel_245787;
  wire [7:0] add_245790;
  wire [7:0] sel_245791;
  wire [7:0] add_245794;
  wire [7:0] sel_245795;
  wire [7:0] add_245798;
  wire [7:0] sel_245799;
  wire [7:0] add_245802;
  wire [7:0] sel_245803;
  wire [7:0] add_245806;
  wire [7:0] sel_245807;
  wire [7:0] add_245810;
  wire [7:0] sel_245811;
  wire [7:0] add_245814;
  wire [7:0] sel_245815;
  wire [7:0] add_245818;
  wire [7:0] sel_245819;
  wire [7:0] add_245822;
  wire [7:0] sel_245823;
  wire [7:0] add_245826;
  wire [7:0] sel_245827;
  wire [7:0] add_245830;
  wire [7:0] sel_245831;
  wire [7:0] add_245834;
  wire [7:0] sel_245835;
  wire [7:0] add_245838;
  wire [7:0] sel_245839;
  wire [7:0] add_245842;
  wire [7:0] sel_245843;
  wire [7:0] add_245846;
  wire [7:0] sel_245847;
  wire [7:0] add_245850;
  wire [7:0] sel_245851;
  wire [7:0] add_245854;
  wire [7:0] sel_245855;
  wire [7:0] add_245858;
  wire [7:0] sel_245859;
  wire [7:0] add_245862;
  wire [7:0] sel_245863;
  wire [7:0] add_245866;
  wire [7:0] sel_245867;
  wire [7:0] add_245870;
  wire [7:0] sel_245871;
  wire [7:0] add_245874;
  wire [7:0] sel_245875;
  wire [7:0] add_245878;
  wire [7:0] sel_245879;
  wire [7:0] add_245883;
  wire [15:0] array_index_245884;
  wire [7:0] sel_245885;
  wire [7:0] add_245888;
  wire [7:0] sel_245889;
  wire [7:0] add_245892;
  wire [7:0] sel_245893;
  wire [7:0] add_245896;
  wire [7:0] sel_245897;
  wire [7:0] add_245900;
  wire [7:0] sel_245901;
  wire [7:0] add_245904;
  wire [7:0] sel_245905;
  wire [7:0] add_245908;
  wire [7:0] sel_245909;
  wire [7:0] add_245912;
  wire [7:0] sel_245913;
  wire [7:0] add_245916;
  wire [7:0] sel_245917;
  wire [7:0] add_245920;
  wire [7:0] sel_245921;
  wire [7:0] add_245924;
  wire [7:0] sel_245925;
  wire [7:0] add_245928;
  wire [7:0] sel_245929;
  wire [7:0] add_245932;
  wire [7:0] sel_245933;
  wire [7:0] add_245936;
  wire [7:0] sel_245937;
  wire [7:0] add_245940;
  wire [7:0] sel_245941;
  wire [7:0] add_245944;
  wire [7:0] sel_245945;
  wire [7:0] add_245948;
  wire [7:0] sel_245949;
  wire [7:0] add_245952;
  wire [7:0] sel_245953;
  wire [7:0] add_245956;
  wire [7:0] sel_245957;
  wire [7:0] add_245960;
  wire [7:0] sel_245961;
  wire [7:0] add_245964;
  wire [7:0] sel_245965;
  wire [7:0] add_245968;
  wire [7:0] sel_245969;
  wire [7:0] add_245972;
  wire [7:0] sel_245973;
  wire [7:0] add_245976;
  wire [7:0] sel_245977;
  wire [7:0] add_245980;
  wire [7:0] sel_245981;
  wire [7:0] add_245984;
  wire [7:0] sel_245985;
  wire [7:0] add_245988;
  wire [7:0] sel_245989;
  wire [7:0] add_245992;
  wire [7:0] sel_245993;
  wire [7:0] add_245996;
  wire [7:0] sel_245997;
  wire [7:0] add_246000;
  wire [7:0] sel_246001;
  wire [7:0] add_246004;
  wire [7:0] sel_246005;
  wire [7:0] add_246008;
  wire [7:0] sel_246009;
  wire [7:0] add_246012;
  wire [7:0] sel_246013;
  wire [7:0] add_246016;
  wire [7:0] sel_246017;
  wire [7:0] add_246020;
  wire [7:0] sel_246021;
  wire [7:0] add_246024;
  wire [7:0] sel_246025;
  wire [7:0] add_246028;
  wire [7:0] sel_246029;
  wire [7:0] add_246032;
  wire [7:0] sel_246033;
  wire [7:0] add_246036;
  wire [7:0] sel_246037;
  wire [7:0] add_246040;
  wire [7:0] sel_246041;
  wire [7:0] add_246044;
  wire [7:0] sel_246045;
  wire [7:0] add_246048;
  wire [7:0] sel_246049;
  wire [7:0] add_246052;
  wire [7:0] sel_246053;
  wire [7:0] add_246056;
  wire [7:0] sel_246057;
  wire [7:0] add_246060;
  wire [7:0] sel_246061;
  wire [7:0] add_246064;
  wire [7:0] sel_246065;
  wire [7:0] add_246068;
  wire [7:0] sel_246069;
  wire [7:0] add_246072;
  wire [7:0] sel_246073;
  wire [7:0] add_246076;
  wire [7:0] sel_246077;
  wire [7:0] add_246080;
  wire [7:0] sel_246081;
  wire [7:0] add_246085;
  wire [15:0] array_index_246086;
  wire [7:0] sel_246087;
  wire [7:0] add_246090;
  wire [7:0] sel_246091;
  wire [7:0] add_246094;
  wire [7:0] sel_246095;
  wire [7:0] add_246098;
  wire [7:0] sel_246099;
  wire [7:0] add_246102;
  wire [7:0] sel_246103;
  wire [7:0] add_246106;
  wire [7:0] sel_246107;
  wire [7:0] add_246110;
  wire [7:0] sel_246111;
  wire [7:0] add_246114;
  wire [7:0] sel_246115;
  wire [7:0] add_246118;
  wire [7:0] sel_246119;
  wire [7:0] add_246122;
  wire [7:0] sel_246123;
  wire [7:0] add_246126;
  wire [7:0] sel_246127;
  wire [7:0] add_246130;
  wire [7:0] sel_246131;
  wire [7:0] add_246134;
  wire [7:0] sel_246135;
  wire [7:0] add_246138;
  wire [7:0] sel_246139;
  wire [7:0] add_246142;
  wire [7:0] sel_246143;
  wire [7:0] add_246146;
  wire [7:0] sel_246147;
  wire [7:0] add_246150;
  wire [7:0] sel_246151;
  wire [7:0] add_246154;
  wire [7:0] sel_246155;
  wire [7:0] add_246158;
  wire [7:0] sel_246159;
  wire [7:0] add_246162;
  wire [7:0] sel_246163;
  wire [7:0] add_246166;
  wire [7:0] sel_246167;
  wire [7:0] add_246170;
  wire [7:0] sel_246171;
  wire [7:0] add_246174;
  wire [7:0] sel_246175;
  wire [7:0] add_246178;
  wire [7:0] sel_246179;
  wire [7:0] add_246182;
  wire [7:0] sel_246183;
  wire [7:0] add_246186;
  wire [7:0] sel_246187;
  wire [7:0] add_246190;
  wire [7:0] sel_246191;
  wire [7:0] add_246194;
  wire [7:0] sel_246195;
  wire [7:0] add_246198;
  wire [7:0] sel_246199;
  wire [7:0] add_246202;
  wire [7:0] sel_246203;
  wire [7:0] add_246206;
  wire [7:0] sel_246207;
  wire [7:0] add_246210;
  wire [7:0] sel_246211;
  wire [7:0] add_246214;
  wire [7:0] sel_246215;
  wire [7:0] add_246218;
  wire [7:0] sel_246219;
  wire [7:0] add_246222;
  wire [7:0] sel_246223;
  wire [7:0] add_246226;
  wire [7:0] sel_246227;
  wire [7:0] add_246230;
  wire [7:0] sel_246231;
  wire [7:0] add_246234;
  wire [7:0] sel_246235;
  wire [7:0] add_246238;
  wire [7:0] sel_246239;
  wire [7:0] add_246242;
  wire [7:0] sel_246243;
  wire [7:0] add_246246;
  wire [7:0] sel_246247;
  wire [7:0] add_246250;
  wire [7:0] sel_246251;
  wire [7:0] add_246254;
  wire [7:0] sel_246255;
  wire [7:0] add_246258;
  wire [7:0] sel_246259;
  wire [7:0] add_246262;
  wire [7:0] sel_246263;
  wire [7:0] add_246266;
  wire [7:0] sel_246267;
  wire [7:0] add_246270;
  wire [7:0] sel_246271;
  wire [7:0] add_246274;
  wire [7:0] sel_246275;
  wire [7:0] add_246278;
  wire [7:0] sel_246279;
  wire [7:0] add_246282;
  wire [7:0] sel_246283;
  wire [7:0] add_246287;
  wire [15:0] array_index_246288;
  wire [7:0] sel_246289;
  wire [7:0] add_246292;
  wire [7:0] sel_246293;
  wire [7:0] add_246296;
  wire [7:0] sel_246297;
  wire [7:0] add_246300;
  wire [7:0] sel_246301;
  wire [7:0] add_246304;
  wire [7:0] sel_246305;
  wire [7:0] add_246308;
  wire [7:0] sel_246309;
  wire [7:0] add_246312;
  wire [7:0] sel_246313;
  wire [7:0] add_246316;
  wire [7:0] sel_246317;
  wire [7:0] add_246320;
  wire [7:0] sel_246321;
  wire [7:0] add_246324;
  wire [7:0] sel_246325;
  wire [7:0] add_246328;
  wire [7:0] sel_246329;
  wire [7:0] add_246332;
  wire [7:0] sel_246333;
  wire [7:0] add_246336;
  wire [7:0] sel_246337;
  wire [7:0] add_246340;
  wire [7:0] sel_246341;
  wire [7:0] add_246344;
  wire [7:0] sel_246345;
  wire [7:0] add_246348;
  wire [7:0] sel_246349;
  wire [7:0] add_246352;
  wire [7:0] sel_246353;
  wire [7:0] add_246356;
  wire [7:0] sel_246357;
  wire [7:0] add_246360;
  wire [7:0] sel_246361;
  wire [7:0] add_246364;
  wire [7:0] sel_246365;
  wire [7:0] add_246368;
  wire [7:0] sel_246369;
  wire [7:0] add_246372;
  wire [7:0] sel_246373;
  wire [7:0] add_246376;
  wire [7:0] sel_246377;
  wire [7:0] add_246380;
  wire [7:0] sel_246381;
  wire [7:0] add_246384;
  wire [7:0] sel_246385;
  wire [7:0] add_246388;
  wire [7:0] sel_246389;
  wire [7:0] add_246392;
  wire [7:0] sel_246393;
  wire [7:0] add_246396;
  wire [7:0] sel_246397;
  wire [7:0] add_246400;
  wire [7:0] sel_246401;
  wire [7:0] add_246404;
  wire [7:0] sel_246405;
  wire [7:0] add_246408;
  wire [7:0] sel_246409;
  wire [7:0] add_246412;
  wire [7:0] sel_246413;
  wire [7:0] add_246416;
  wire [7:0] sel_246417;
  wire [7:0] add_246420;
  wire [7:0] sel_246421;
  wire [7:0] add_246424;
  wire [7:0] sel_246425;
  wire [7:0] add_246428;
  wire [7:0] sel_246429;
  wire [7:0] add_246432;
  wire [7:0] sel_246433;
  wire [7:0] add_246436;
  wire [7:0] sel_246437;
  wire [7:0] add_246440;
  wire [7:0] sel_246441;
  wire [7:0] add_246444;
  wire [7:0] sel_246445;
  wire [7:0] add_246448;
  wire [7:0] sel_246449;
  wire [7:0] add_246452;
  wire [7:0] sel_246453;
  wire [7:0] add_246456;
  wire [7:0] sel_246457;
  wire [7:0] add_246460;
  wire [7:0] sel_246461;
  wire [7:0] add_246464;
  wire [7:0] sel_246465;
  wire [7:0] add_246468;
  wire [7:0] sel_246469;
  wire [7:0] add_246472;
  wire [7:0] sel_246473;
  wire [7:0] add_246476;
  wire [7:0] sel_246477;
  wire [7:0] add_246480;
  wire [7:0] sel_246481;
  wire [7:0] add_246484;
  wire [7:0] sel_246485;
  wire [7:0] add_246489;
  wire [15:0] array_index_246490;
  wire [7:0] sel_246491;
  wire [7:0] add_246494;
  wire [7:0] sel_246495;
  wire [7:0] add_246498;
  wire [7:0] sel_246499;
  wire [7:0] add_246502;
  wire [7:0] sel_246503;
  wire [7:0] add_246506;
  wire [7:0] sel_246507;
  wire [7:0] add_246510;
  wire [7:0] sel_246511;
  wire [7:0] add_246514;
  wire [7:0] sel_246515;
  wire [7:0] add_246518;
  wire [7:0] sel_246519;
  wire [7:0] add_246522;
  wire [7:0] sel_246523;
  wire [7:0] add_246526;
  wire [7:0] sel_246527;
  wire [7:0] add_246530;
  wire [7:0] sel_246531;
  wire [7:0] add_246534;
  wire [7:0] sel_246535;
  wire [7:0] add_246538;
  wire [7:0] sel_246539;
  wire [7:0] add_246542;
  wire [7:0] sel_246543;
  wire [7:0] add_246546;
  wire [7:0] sel_246547;
  wire [7:0] add_246550;
  wire [7:0] sel_246551;
  wire [7:0] add_246554;
  wire [7:0] sel_246555;
  wire [7:0] add_246558;
  wire [7:0] sel_246559;
  wire [7:0] add_246562;
  wire [7:0] sel_246563;
  wire [7:0] add_246566;
  wire [7:0] sel_246567;
  wire [7:0] add_246570;
  wire [7:0] sel_246571;
  wire [7:0] add_246574;
  wire [7:0] sel_246575;
  wire [7:0] add_246578;
  wire [7:0] sel_246579;
  wire [7:0] add_246582;
  wire [7:0] sel_246583;
  wire [7:0] add_246586;
  wire [7:0] sel_246587;
  wire [7:0] add_246590;
  wire [7:0] sel_246591;
  wire [7:0] add_246594;
  wire [7:0] sel_246595;
  wire [7:0] add_246598;
  wire [7:0] sel_246599;
  wire [7:0] add_246602;
  wire [7:0] sel_246603;
  wire [7:0] add_246606;
  wire [7:0] sel_246607;
  wire [7:0] add_246610;
  wire [7:0] sel_246611;
  wire [7:0] add_246614;
  wire [7:0] sel_246615;
  wire [7:0] add_246618;
  wire [7:0] sel_246619;
  wire [7:0] add_246622;
  wire [7:0] sel_246623;
  wire [7:0] add_246626;
  wire [7:0] sel_246627;
  wire [7:0] add_246630;
  wire [7:0] sel_246631;
  wire [7:0] add_246634;
  wire [7:0] sel_246635;
  wire [7:0] add_246638;
  wire [7:0] sel_246639;
  wire [7:0] add_246642;
  wire [7:0] sel_246643;
  wire [7:0] add_246646;
  wire [7:0] sel_246647;
  wire [7:0] add_246650;
  wire [7:0] sel_246651;
  wire [7:0] add_246654;
  wire [7:0] sel_246655;
  wire [7:0] add_246658;
  wire [7:0] sel_246659;
  wire [7:0] add_246662;
  wire [7:0] sel_246663;
  wire [7:0] add_246666;
  wire [7:0] sel_246667;
  wire [7:0] add_246670;
  wire [7:0] sel_246671;
  wire [7:0] add_246674;
  wire [7:0] sel_246675;
  wire [7:0] add_246678;
  wire [7:0] sel_246679;
  wire [7:0] add_246682;
  wire [7:0] sel_246683;
  wire [7:0] add_246686;
  wire [7:0] sel_246687;
  wire [7:0] add_246691;
  wire [15:0] array_index_246692;
  wire [7:0] sel_246693;
  wire [7:0] add_246696;
  wire [7:0] sel_246697;
  wire [7:0] add_246700;
  wire [7:0] sel_246701;
  wire [7:0] add_246704;
  wire [7:0] sel_246705;
  wire [7:0] add_246708;
  wire [7:0] sel_246709;
  wire [7:0] add_246712;
  wire [7:0] sel_246713;
  wire [7:0] add_246716;
  wire [7:0] sel_246717;
  wire [7:0] add_246720;
  wire [7:0] sel_246721;
  wire [7:0] add_246724;
  wire [7:0] sel_246725;
  wire [7:0] add_246728;
  wire [7:0] sel_246729;
  wire [7:0] add_246732;
  wire [7:0] sel_246733;
  wire [7:0] add_246736;
  wire [7:0] sel_246737;
  wire [7:0] add_246740;
  wire [7:0] sel_246741;
  wire [7:0] add_246744;
  wire [7:0] sel_246745;
  wire [7:0] add_246748;
  wire [7:0] sel_246749;
  wire [7:0] add_246752;
  wire [7:0] sel_246753;
  wire [7:0] add_246756;
  wire [7:0] sel_246757;
  wire [7:0] add_246760;
  wire [7:0] sel_246761;
  wire [7:0] add_246764;
  wire [7:0] sel_246765;
  wire [7:0] add_246768;
  wire [7:0] sel_246769;
  wire [7:0] add_246772;
  wire [7:0] sel_246773;
  wire [7:0] add_246776;
  wire [7:0] sel_246777;
  wire [7:0] add_246780;
  wire [7:0] sel_246781;
  wire [7:0] add_246784;
  wire [7:0] sel_246785;
  wire [7:0] add_246788;
  wire [7:0] sel_246789;
  wire [7:0] add_246792;
  wire [7:0] sel_246793;
  wire [7:0] add_246796;
  wire [7:0] sel_246797;
  wire [7:0] add_246800;
  wire [7:0] sel_246801;
  wire [7:0] add_246804;
  wire [7:0] sel_246805;
  wire [7:0] add_246808;
  wire [7:0] sel_246809;
  wire [7:0] add_246812;
  wire [7:0] sel_246813;
  wire [7:0] add_246816;
  wire [7:0] sel_246817;
  wire [7:0] add_246820;
  wire [7:0] sel_246821;
  wire [7:0] add_246824;
  wire [7:0] sel_246825;
  wire [7:0] add_246828;
  wire [7:0] sel_246829;
  wire [7:0] add_246832;
  wire [7:0] sel_246833;
  wire [7:0] add_246836;
  wire [7:0] sel_246837;
  wire [7:0] add_246840;
  wire [7:0] sel_246841;
  wire [7:0] add_246844;
  wire [7:0] sel_246845;
  wire [7:0] add_246848;
  wire [7:0] sel_246849;
  wire [7:0] add_246852;
  wire [7:0] sel_246853;
  wire [7:0] add_246856;
  wire [7:0] sel_246857;
  wire [7:0] add_246860;
  wire [7:0] sel_246861;
  wire [7:0] add_246864;
  wire [7:0] sel_246865;
  wire [7:0] add_246868;
  wire [7:0] sel_246869;
  wire [7:0] add_246872;
  wire [7:0] sel_246873;
  wire [7:0] add_246876;
  wire [7:0] sel_246877;
  wire [7:0] add_246880;
  wire [7:0] sel_246881;
  wire [7:0] add_246884;
  wire [7:0] sel_246885;
  wire [7:0] add_246888;
  wire [7:0] sel_246889;
  wire [7:0] add_246893;
  wire [15:0] array_index_246894;
  wire [7:0] sel_246895;
  wire [7:0] add_246898;
  wire [7:0] sel_246899;
  wire [7:0] add_246902;
  wire [7:0] sel_246903;
  wire [7:0] add_246906;
  wire [7:0] sel_246907;
  wire [7:0] add_246910;
  wire [7:0] sel_246911;
  wire [7:0] add_246914;
  wire [7:0] sel_246915;
  wire [7:0] add_246918;
  wire [7:0] sel_246919;
  wire [7:0] add_246922;
  wire [7:0] sel_246923;
  wire [7:0] add_246926;
  wire [7:0] sel_246927;
  wire [7:0] add_246930;
  wire [7:0] sel_246931;
  wire [7:0] add_246934;
  wire [7:0] sel_246935;
  wire [7:0] add_246938;
  wire [7:0] sel_246939;
  wire [7:0] add_246942;
  wire [7:0] sel_246943;
  wire [7:0] add_246946;
  wire [7:0] sel_246947;
  wire [7:0] add_246950;
  wire [7:0] sel_246951;
  wire [7:0] add_246954;
  wire [7:0] sel_246955;
  wire [7:0] add_246958;
  wire [7:0] sel_246959;
  wire [7:0] add_246962;
  wire [7:0] sel_246963;
  wire [7:0] add_246966;
  wire [7:0] sel_246967;
  wire [7:0] add_246970;
  wire [7:0] sel_246971;
  wire [7:0] add_246974;
  wire [7:0] sel_246975;
  wire [7:0] add_246978;
  wire [7:0] sel_246979;
  wire [7:0] add_246982;
  wire [7:0] sel_246983;
  wire [7:0] add_246986;
  wire [7:0] sel_246987;
  wire [7:0] add_246990;
  wire [7:0] sel_246991;
  wire [7:0] add_246994;
  wire [7:0] sel_246995;
  wire [7:0] add_246998;
  wire [7:0] sel_246999;
  wire [7:0] add_247002;
  wire [7:0] sel_247003;
  wire [7:0] add_247006;
  wire [7:0] sel_247007;
  wire [7:0] add_247010;
  wire [7:0] sel_247011;
  wire [7:0] add_247014;
  wire [7:0] sel_247015;
  wire [7:0] add_247018;
  wire [7:0] sel_247019;
  wire [7:0] add_247022;
  wire [7:0] sel_247023;
  wire [7:0] add_247026;
  wire [7:0] sel_247027;
  wire [7:0] add_247030;
  wire [7:0] sel_247031;
  wire [7:0] add_247034;
  wire [7:0] sel_247035;
  wire [7:0] add_247038;
  wire [7:0] sel_247039;
  wire [7:0] add_247042;
  wire [7:0] sel_247043;
  wire [7:0] add_247046;
  wire [7:0] sel_247047;
  wire [7:0] add_247050;
  wire [7:0] sel_247051;
  wire [7:0] add_247054;
  wire [7:0] sel_247055;
  wire [7:0] add_247058;
  wire [7:0] sel_247059;
  wire [7:0] add_247062;
  wire [7:0] sel_247063;
  wire [7:0] add_247066;
  wire [7:0] sel_247067;
  wire [7:0] add_247070;
  wire [7:0] sel_247071;
  wire [7:0] add_247074;
  wire [7:0] sel_247075;
  wire [7:0] add_247078;
  wire [7:0] sel_247079;
  wire [7:0] add_247082;
  wire [7:0] sel_247083;
  wire [7:0] add_247086;
  wire [7:0] sel_247087;
  wire [7:0] add_247090;
  wire [7:0] sel_247091;
  wire [7:0] add_247095;
  wire [15:0] array_index_247096;
  wire [7:0] sel_247097;
  wire [7:0] add_247100;
  wire [7:0] sel_247101;
  wire [7:0] add_247104;
  wire [7:0] sel_247105;
  wire [7:0] add_247108;
  wire [7:0] sel_247109;
  wire [7:0] add_247112;
  wire [7:0] sel_247113;
  wire [7:0] add_247116;
  wire [7:0] sel_247117;
  wire [7:0] add_247120;
  wire [7:0] sel_247121;
  wire [7:0] add_247124;
  wire [7:0] sel_247125;
  wire [7:0] add_247128;
  wire [7:0] sel_247129;
  wire [7:0] add_247132;
  wire [7:0] sel_247133;
  wire [7:0] add_247136;
  wire [7:0] sel_247137;
  wire [7:0] add_247140;
  wire [7:0] sel_247141;
  wire [7:0] add_247144;
  wire [7:0] sel_247145;
  wire [7:0] add_247148;
  wire [7:0] sel_247149;
  wire [7:0] add_247152;
  wire [7:0] sel_247153;
  wire [7:0] add_247156;
  wire [7:0] sel_247157;
  wire [7:0] add_247160;
  wire [7:0] sel_247161;
  wire [7:0] add_247164;
  wire [7:0] sel_247165;
  wire [7:0] add_247168;
  wire [7:0] sel_247169;
  wire [7:0] add_247172;
  wire [7:0] sel_247173;
  wire [7:0] add_247176;
  wire [7:0] sel_247177;
  wire [7:0] add_247180;
  wire [7:0] sel_247181;
  wire [7:0] add_247184;
  wire [7:0] sel_247185;
  wire [7:0] add_247188;
  wire [7:0] sel_247189;
  wire [7:0] add_247192;
  wire [7:0] sel_247193;
  wire [7:0] add_247196;
  wire [7:0] sel_247197;
  wire [7:0] add_247200;
  wire [7:0] sel_247201;
  wire [7:0] add_247204;
  wire [7:0] sel_247205;
  wire [7:0] add_247208;
  wire [7:0] sel_247209;
  wire [7:0] add_247212;
  wire [7:0] sel_247213;
  wire [7:0] add_247216;
  wire [7:0] sel_247217;
  wire [7:0] add_247220;
  wire [7:0] sel_247221;
  wire [7:0] add_247224;
  wire [7:0] sel_247225;
  wire [7:0] add_247228;
  wire [7:0] sel_247229;
  wire [7:0] add_247232;
  wire [7:0] sel_247233;
  wire [7:0] add_247236;
  wire [7:0] sel_247237;
  wire [7:0] add_247240;
  wire [7:0] sel_247241;
  wire [7:0] add_247244;
  wire [7:0] sel_247245;
  wire [7:0] add_247248;
  wire [7:0] sel_247249;
  wire [7:0] add_247252;
  wire [7:0] sel_247253;
  wire [7:0] add_247256;
  wire [7:0] sel_247257;
  wire [7:0] add_247260;
  wire [7:0] sel_247261;
  wire [7:0] add_247264;
  wire [7:0] sel_247265;
  wire [7:0] add_247268;
  wire [7:0] sel_247269;
  wire [7:0] add_247272;
  wire [7:0] sel_247273;
  wire [7:0] add_247276;
  wire [7:0] sel_247277;
  wire [7:0] add_247280;
  wire [7:0] sel_247281;
  wire [7:0] add_247284;
  wire [7:0] sel_247285;
  wire [7:0] add_247288;
  wire [7:0] sel_247289;
  wire [7:0] add_247292;
  wire [7:0] sel_247293;
  wire [7:0] add_247297;
  wire [15:0] array_index_247298;
  wire [7:0] sel_247299;
  wire [7:0] add_247302;
  wire [7:0] sel_247303;
  wire [7:0] add_247306;
  wire [7:0] sel_247307;
  wire [7:0] add_247310;
  wire [7:0] sel_247311;
  wire [7:0] add_247314;
  wire [7:0] sel_247315;
  wire [7:0] add_247318;
  wire [7:0] sel_247319;
  wire [7:0] add_247322;
  wire [7:0] sel_247323;
  wire [7:0] add_247326;
  wire [7:0] sel_247327;
  wire [7:0] add_247330;
  wire [7:0] sel_247331;
  wire [7:0] add_247334;
  wire [7:0] sel_247335;
  wire [7:0] add_247338;
  wire [7:0] sel_247339;
  wire [7:0] add_247342;
  wire [7:0] sel_247343;
  wire [7:0] add_247346;
  wire [7:0] sel_247347;
  wire [7:0] add_247350;
  wire [7:0] sel_247351;
  wire [7:0] add_247354;
  wire [7:0] sel_247355;
  wire [7:0] add_247358;
  wire [7:0] sel_247359;
  wire [7:0] add_247362;
  wire [7:0] sel_247363;
  wire [7:0] add_247366;
  wire [7:0] sel_247367;
  wire [7:0] add_247370;
  wire [7:0] sel_247371;
  wire [7:0] add_247374;
  wire [7:0] sel_247375;
  wire [7:0] add_247378;
  wire [7:0] sel_247379;
  wire [7:0] add_247382;
  wire [7:0] sel_247383;
  wire [7:0] add_247386;
  wire [7:0] sel_247387;
  wire [7:0] add_247390;
  wire [7:0] sel_247391;
  wire [7:0] add_247394;
  wire [7:0] sel_247395;
  wire [7:0] add_247398;
  wire [7:0] sel_247399;
  wire [7:0] add_247402;
  wire [7:0] sel_247403;
  wire [7:0] add_247406;
  wire [7:0] sel_247407;
  wire [7:0] add_247410;
  wire [7:0] sel_247411;
  wire [7:0] add_247414;
  wire [7:0] sel_247415;
  wire [7:0] add_247418;
  wire [7:0] sel_247419;
  wire [7:0] add_247422;
  wire [7:0] sel_247423;
  wire [7:0] add_247426;
  wire [7:0] sel_247427;
  wire [7:0] add_247430;
  wire [7:0] sel_247431;
  wire [7:0] add_247434;
  wire [7:0] sel_247435;
  wire [7:0] add_247438;
  wire [7:0] sel_247439;
  wire [7:0] add_247442;
  wire [7:0] sel_247443;
  wire [7:0] add_247446;
  wire [7:0] sel_247447;
  wire [7:0] add_247450;
  wire [7:0] sel_247451;
  wire [7:0] add_247454;
  wire [7:0] sel_247455;
  wire [7:0] add_247458;
  wire [7:0] sel_247459;
  wire [7:0] add_247462;
  wire [7:0] sel_247463;
  wire [7:0] add_247466;
  wire [7:0] sel_247467;
  wire [7:0] add_247470;
  wire [7:0] sel_247471;
  wire [7:0] add_247474;
  wire [7:0] sel_247475;
  wire [7:0] add_247478;
  wire [7:0] sel_247479;
  wire [7:0] add_247482;
  wire [7:0] sel_247483;
  wire [7:0] add_247486;
  wire [7:0] sel_247487;
  wire [7:0] add_247490;
  wire [7:0] sel_247491;
  wire [7:0] add_247494;
  wire [7:0] sel_247495;
  wire [7:0] add_247499;
  wire [15:0] array_index_247500;
  wire [7:0] sel_247501;
  wire [7:0] add_247504;
  wire [7:0] sel_247505;
  wire [7:0] add_247508;
  wire [7:0] sel_247509;
  wire [7:0] add_247512;
  wire [7:0] sel_247513;
  wire [7:0] add_247516;
  wire [7:0] sel_247517;
  wire [7:0] add_247520;
  wire [7:0] sel_247521;
  wire [7:0] add_247524;
  wire [7:0] sel_247525;
  wire [7:0] add_247528;
  wire [7:0] sel_247529;
  wire [7:0] add_247532;
  wire [7:0] sel_247533;
  wire [7:0] add_247536;
  wire [7:0] sel_247537;
  wire [7:0] add_247540;
  wire [7:0] sel_247541;
  wire [7:0] add_247544;
  wire [7:0] sel_247545;
  wire [7:0] add_247548;
  wire [7:0] sel_247549;
  wire [7:0] add_247552;
  wire [7:0] sel_247553;
  wire [7:0] add_247556;
  wire [7:0] sel_247557;
  wire [7:0] add_247560;
  wire [7:0] sel_247561;
  wire [7:0] add_247564;
  wire [7:0] sel_247565;
  wire [7:0] add_247568;
  wire [7:0] sel_247569;
  wire [7:0] add_247572;
  wire [7:0] sel_247573;
  wire [7:0] add_247576;
  wire [7:0] sel_247577;
  wire [7:0] add_247580;
  wire [7:0] sel_247581;
  wire [7:0] add_247584;
  wire [7:0] sel_247585;
  wire [7:0] add_247588;
  wire [7:0] sel_247589;
  wire [7:0] add_247592;
  wire [7:0] sel_247593;
  wire [7:0] add_247596;
  wire [7:0] sel_247597;
  wire [7:0] add_247600;
  wire [7:0] sel_247601;
  wire [7:0] add_247604;
  wire [7:0] sel_247605;
  wire [7:0] add_247608;
  wire [7:0] sel_247609;
  wire [7:0] add_247612;
  wire [7:0] sel_247613;
  wire [7:0] add_247616;
  wire [7:0] sel_247617;
  wire [7:0] add_247620;
  wire [7:0] sel_247621;
  wire [7:0] add_247624;
  wire [7:0] sel_247625;
  wire [7:0] add_247628;
  wire [7:0] sel_247629;
  wire [7:0] add_247632;
  wire [7:0] sel_247633;
  wire [7:0] add_247636;
  wire [7:0] sel_247637;
  wire [7:0] add_247640;
  wire [7:0] sel_247641;
  wire [7:0] add_247644;
  wire [7:0] sel_247645;
  wire [7:0] add_247648;
  wire [7:0] sel_247649;
  wire [7:0] add_247652;
  wire [7:0] sel_247653;
  wire [7:0] add_247656;
  wire [7:0] sel_247657;
  wire [7:0] add_247660;
  wire [7:0] sel_247661;
  wire [7:0] add_247664;
  wire [7:0] sel_247665;
  wire [7:0] add_247668;
  wire [7:0] sel_247669;
  wire [7:0] add_247672;
  wire [7:0] sel_247673;
  wire [7:0] add_247676;
  wire [7:0] sel_247677;
  wire [7:0] add_247680;
  wire [7:0] sel_247681;
  wire [7:0] add_247684;
  wire [7:0] sel_247685;
  wire [7:0] add_247688;
  wire [7:0] sel_247689;
  wire [7:0] add_247692;
  wire [7:0] sel_247693;
  wire [7:0] add_247696;
  wire [7:0] sel_247697;
  wire [7:0] add_247701;
  wire [15:0] array_index_247702;
  wire [7:0] sel_247703;
  wire [7:0] add_247706;
  wire [7:0] sel_247707;
  wire [7:0] add_247710;
  wire [7:0] sel_247711;
  wire [7:0] add_247714;
  wire [7:0] sel_247715;
  wire [7:0] add_247718;
  wire [7:0] sel_247719;
  wire [7:0] add_247722;
  wire [7:0] sel_247723;
  wire [7:0] add_247726;
  wire [7:0] sel_247727;
  wire [7:0] add_247730;
  wire [7:0] sel_247731;
  wire [7:0] add_247734;
  wire [7:0] sel_247735;
  wire [7:0] add_247738;
  wire [7:0] sel_247739;
  wire [7:0] add_247742;
  wire [7:0] sel_247743;
  wire [7:0] add_247746;
  wire [7:0] sel_247747;
  wire [7:0] add_247750;
  wire [7:0] sel_247751;
  wire [7:0] add_247754;
  wire [7:0] sel_247755;
  wire [7:0] add_247758;
  wire [7:0] sel_247759;
  wire [7:0] add_247762;
  wire [7:0] sel_247763;
  wire [7:0] add_247766;
  wire [7:0] sel_247767;
  wire [7:0] add_247770;
  wire [7:0] sel_247771;
  wire [7:0] add_247774;
  wire [7:0] sel_247775;
  wire [7:0] add_247778;
  wire [7:0] sel_247779;
  wire [7:0] add_247782;
  wire [7:0] sel_247783;
  wire [7:0] add_247786;
  wire [7:0] sel_247787;
  wire [7:0] add_247790;
  wire [7:0] sel_247791;
  wire [7:0] add_247794;
  wire [7:0] sel_247795;
  wire [7:0] add_247798;
  wire [7:0] sel_247799;
  wire [7:0] add_247802;
  wire [7:0] sel_247803;
  wire [7:0] add_247806;
  wire [7:0] sel_247807;
  wire [7:0] add_247810;
  wire [7:0] sel_247811;
  wire [7:0] add_247814;
  wire [7:0] sel_247815;
  wire [7:0] add_247818;
  wire [7:0] sel_247819;
  wire [7:0] add_247822;
  wire [7:0] sel_247823;
  wire [7:0] add_247826;
  wire [7:0] sel_247827;
  wire [7:0] add_247830;
  wire [7:0] sel_247831;
  wire [7:0] add_247834;
  wire [7:0] sel_247835;
  wire [7:0] add_247838;
  wire [7:0] sel_247839;
  wire [7:0] add_247842;
  wire [7:0] sel_247843;
  wire [7:0] add_247846;
  wire [7:0] sel_247847;
  wire [7:0] add_247850;
  wire [7:0] sel_247851;
  wire [7:0] add_247854;
  wire [7:0] sel_247855;
  wire [7:0] add_247858;
  wire [7:0] sel_247859;
  wire [7:0] add_247862;
  wire [7:0] sel_247863;
  wire [7:0] add_247866;
  wire [7:0] sel_247867;
  wire [7:0] add_247870;
  wire [7:0] sel_247871;
  wire [7:0] add_247874;
  wire [7:0] sel_247875;
  wire [7:0] add_247878;
  wire [7:0] sel_247879;
  wire [7:0] add_247882;
  wire [7:0] sel_247883;
  wire [7:0] add_247886;
  wire [7:0] sel_247887;
  wire [7:0] add_247890;
  wire [7:0] sel_247891;
  wire [7:0] add_247894;
  wire [7:0] sel_247895;
  wire [7:0] add_247898;
  wire [7:0] sel_247899;
  wire [7:0] add_247903;
  wire [15:0] array_index_247904;
  wire [7:0] sel_247905;
  wire [7:0] add_247908;
  wire [7:0] sel_247909;
  wire [7:0] add_247912;
  wire [7:0] sel_247913;
  wire [7:0] add_247916;
  wire [7:0] sel_247917;
  wire [7:0] add_247920;
  wire [7:0] sel_247921;
  wire [7:0] add_247924;
  wire [7:0] sel_247925;
  wire [7:0] add_247928;
  wire [7:0] sel_247929;
  wire [7:0] add_247932;
  wire [7:0] sel_247933;
  wire [7:0] add_247936;
  wire [7:0] sel_247937;
  wire [7:0] add_247940;
  wire [7:0] sel_247941;
  wire [7:0] add_247944;
  wire [7:0] sel_247945;
  wire [7:0] add_247948;
  wire [7:0] sel_247949;
  wire [7:0] add_247952;
  wire [7:0] sel_247953;
  wire [7:0] add_247956;
  wire [7:0] sel_247957;
  wire [7:0] add_247960;
  wire [7:0] sel_247961;
  wire [7:0] add_247964;
  wire [7:0] sel_247965;
  wire [7:0] add_247968;
  wire [7:0] sel_247969;
  wire [7:0] add_247972;
  wire [7:0] sel_247973;
  wire [7:0] add_247976;
  wire [7:0] sel_247977;
  wire [7:0] add_247980;
  wire [7:0] sel_247981;
  wire [7:0] add_247984;
  wire [7:0] sel_247985;
  wire [7:0] add_247988;
  wire [7:0] sel_247989;
  wire [7:0] add_247992;
  wire [7:0] sel_247993;
  wire [7:0] add_247996;
  wire [7:0] sel_247997;
  wire [7:0] add_248000;
  wire [7:0] sel_248001;
  wire [7:0] add_248004;
  wire [7:0] sel_248005;
  wire [7:0] add_248008;
  wire [7:0] sel_248009;
  wire [7:0] add_248012;
  wire [7:0] sel_248013;
  wire [7:0] add_248016;
  wire [7:0] sel_248017;
  wire [7:0] add_248020;
  wire [7:0] sel_248021;
  wire [7:0] add_248024;
  wire [7:0] sel_248025;
  wire [7:0] add_248028;
  wire [7:0] sel_248029;
  wire [7:0] add_248032;
  wire [7:0] sel_248033;
  wire [7:0] add_248036;
  wire [7:0] sel_248037;
  wire [7:0] add_248040;
  wire [7:0] sel_248041;
  wire [7:0] add_248044;
  wire [7:0] sel_248045;
  wire [7:0] add_248048;
  wire [7:0] sel_248049;
  wire [7:0] add_248052;
  wire [7:0] sel_248053;
  wire [7:0] add_248056;
  wire [7:0] sel_248057;
  wire [7:0] add_248060;
  wire [7:0] sel_248061;
  wire [7:0] add_248064;
  wire [7:0] sel_248065;
  wire [7:0] add_248068;
  wire [7:0] sel_248069;
  wire [7:0] add_248072;
  wire [7:0] sel_248073;
  wire [7:0] add_248076;
  wire [7:0] sel_248077;
  wire [7:0] add_248080;
  wire [7:0] sel_248081;
  wire [7:0] add_248084;
  wire [7:0] sel_248085;
  wire [7:0] add_248088;
  wire [7:0] sel_248089;
  wire [7:0] add_248092;
  wire [7:0] sel_248093;
  wire [7:0] add_248096;
  wire [7:0] sel_248097;
  wire [7:0] add_248100;
  wire [7:0] sel_248101;
  wire [7:0] add_248105;
  wire [15:0] array_index_248106;
  wire [7:0] sel_248107;
  wire [7:0] add_248110;
  wire [7:0] sel_248111;
  wire [7:0] add_248114;
  wire [7:0] sel_248115;
  wire [7:0] add_248118;
  wire [7:0] sel_248119;
  wire [7:0] add_248122;
  wire [7:0] sel_248123;
  wire [7:0] add_248126;
  wire [7:0] sel_248127;
  wire [7:0] add_248130;
  wire [7:0] sel_248131;
  wire [7:0] add_248134;
  wire [7:0] sel_248135;
  wire [7:0] add_248138;
  wire [7:0] sel_248139;
  wire [7:0] add_248142;
  wire [7:0] sel_248143;
  wire [7:0] add_248146;
  wire [7:0] sel_248147;
  wire [7:0] add_248150;
  wire [7:0] sel_248151;
  wire [7:0] add_248154;
  wire [7:0] sel_248155;
  wire [7:0] add_248158;
  wire [7:0] sel_248159;
  wire [7:0] add_248162;
  wire [7:0] sel_248163;
  wire [7:0] add_248166;
  wire [7:0] sel_248167;
  wire [7:0] add_248170;
  wire [7:0] sel_248171;
  wire [7:0] add_248174;
  wire [7:0] sel_248175;
  wire [7:0] add_248178;
  wire [7:0] sel_248179;
  wire [7:0] add_248182;
  wire [7:0] sel_248183;
  wire [7:0] add_248186;
  wire [7:0] sel_248187;
  wire [7:0] add_248190;
  wire [7:0] sel_248191;
  wire [7:0] add_248194;
  wire [7:0] sel_248195;
  wire [7:0] add_248198;
  wire [7:0] sel_248199;
  wire [7:0] add_248202;
  wire [7:0] sel_248203;
  wire [7:0] add_248206;
  wire [7:0] sel_248207;
  wire [7:0] add_248210;
  wire [7:0] sel_248211;
  wire [7:0] add_248214;
  wire [7:0] sel_248215;
  wire [7:0] add_248218;
  wire [7:0] sel_248219;
  wire [7:0] add_248222;
  wire [7:0] sel_248223;
  wire [7:0] add_248226;
  wire [7:0] sel_248227;
  wire [7:0] add_248230;
  wire [7:0] sel_248231;
  wire [7:0] add_248234;
  wire [7:0] sel_248235;
  wire [7:0] add_248238;
  wire [7:0] sel_248239;
  wire [7:0] add_248242;
  wire [7:0] sel_248243;
  wire [7:0] add_248246;
  wire [7:0] sel_248247;
  wire [7:0] add_248250;
  wire [7:0] sel_248251;
  wire [7:0] add_248254;
  wire [7:0] sel_248255;
  wire [7:0] add_248258;
  wire [7:0] sel_248259;
  wire [7:0] add_248262;
  wire [7:0] sel_248263;
  wire [7:0] add_248266;
  wire [7:0] sel_248267;
  wire [7:0] add_248270;
  wire [7:0] sel_248271;
  wire [7:0] add_248274;
  wire [7:0] sel_248275;
  wire [7:0] add_248278;
  wire [7:0] sel_248279;
  wire [7:0] add_248282;
  wire [7:0] sel_248283;
  wire [7:0] add_248286;
  wire [7:0] sel_248287;
  wire [7:0] add_248290;
  wire [7:0] sel_248291;
  wire [7:0] add_248294;
  wire [7:0] sel_248295;
  wire [7:0] add_248298;
  wire [7:0] sel_248299;
  wire [7:0] add_248302;
  wire [7:0] sel_248303;
  wire [7:0] add_248307;
  wire [15:0] array_index_248308;
  wire [7:0] sel_248309;
  wire [7:0] add_248312;
  wire [7:0] sel_248313;
  wire [7:0] add_248316;
  wire [7:0] sel_248317;
  wire [7:0] add_248320;
  wire [7:0] sel_248321;
  wire [7:0] add_248324;
  wire [7:0] sel_248325;
  wire [7:0] add_248328;
  wire [7:0] sel_248329;
  wire [7:0] add_248332;
  wire [7:0] sel_248333;
  wire [7:0] add_248336;
  wire [7:0] sel_248337;
  wire [7:0] add_248340;
  wire [7:0] sel_248341;
  wire [7:0] add_248344;
  wire [7:0] sel_248345;
  wire [7:0] add_248348;
  wire [7:0] sel_248349;
  wire [7:0] add_248352;
  wire [7:0] sel_248353;
  wire [7:0] add_248356;
  wire [7:0] sel_248357;
  wire [7:0] add_248360;
  wire [7:0] sel_248361;
  wire [7:0] add_248364;
  wire [7:0] sel_248365;
  wire [7:0] add_248368;
  wire [7:0] sel_248369;
  wire [7:0] add_248372;
  wire [7:0] sel_248373;
  wire [7:0] add_248376;
  wire [7:0] sel_248377;
  wire [7:0] add_248380;
  wire [7:0] sel_248381;
  wire [7:0] add_248384;
  wire [7:0] sel_248385;
  wire [7:0] add_248388;
  wire [7:0] sel_248389;
  wire [7:0] add_248392;
  wire [7:0] sel_248393;
  wire [7:0] add_248396;
  wire [7:0] sel_248397;
  wire [7:0] add_248400;
  wire [7:0] sel_248401;
  wire [7:0] add_248404;
  wire [7:0] sel_248405;
  wire [7:0] add_248408;
  wire [7:0] sel_248409;
  wire [7:0] add_248412;
  wire [7:0] sel_248413;
  wire [7:0] add_248416;
  wire [7:0] sel_248417;
  wire [7:0] add_248420;
  wire [7:0] sel_248421;
  wire [7:0] add_248424;
  wire [7:0] sel_248425;
  wire [7:0] add_248428;
  wire [7:0] sel_248429;
  wire [7:0] add_248432;
  wire [7:0] sel_248433;
  wire [7:0] add_248436;
  wire [7:0] sel_248437;
  wire [7:0] add_248440;
  wire [7:0] sel_248441;
  wire [7:0] add_248444;
  wire [7:0] sel_248445;
  wire [7:0] add_248448;
  wire [7:0] sel_248449;
  wire [7:0] add_248452;
  wire [7:0] sel_248453;
  wire [7:0] add_248456;
  wire [7:0] sel_248457;
  wire [7:0] add_248460;
  wire [7:0] sel_248461;
  wire [7:0] add_248464;
  wire [7:0] sel_248465;
  wire [7:0] add_248468;
  wire [7:0] sel_248469;
  wire [7:0] add_248472;
  wire [7:0] sel_248473;
  wire [7:0] add_248476;
  wire [7:0] sel_248477;
  wire [7:0] add_248480;
  wire [7:0] sel_248481;
  wire [7:0] add_248484;
  wire [7:0] sel_248485;
  wire [7:0] add_248488;
  wire [7:0] sel_248489;
  wire [7:0] add_248492;
  wire [7:0] sel_248493;
  wire [7:0] add_248496;
  wire [7:0] sel_248497;
  wire [7:0] add_248500;
  wire [7:0] sel_248501;
  wire [7:0] add_248504;
  wire [7:0] sel_248505;
  wire [7:0] add_248509;
  wire [15:0] array_index_248510;
  wire [7:0] sel_248511;
  wire [7:0] add_248514;
  wire [7:0] sel_248515;
  wire [7:0] add_248518;
  wire [7:0] sel_248519;
  wire [7:0] add_248522;
  wire [7:0] sel_248523;
  wire [7:0] add_248526;
  wire [7:0] sel_248527;
  wire [7:0] add_248530;
  wire [7:0] sel_248531;
  wire [7:0] add_248534;
  wire [7:0] sel_248535;
  wire [7:0] add_248538;
  wire [7:0] sel_248539;
  wire [7:0] add_248542;
  wire [7:0] sel_248543;
  wire [7:0] add_248546;
  wire [7:0] sel_248547;
  wire [7:0] add_248550;
  wire [7:0] sel_248551;
  wire [7:0] add_248554;
  wire [7:0] sel_248555;
  wire [7:0] add_248558;
  wire [7:0] sel_248559;
  wire [7:0] add_248562;
  wire [7:0] sel_248563;
  wire [7:0] add_248566;
  wire [7:0] sel_248567;
  wire [7:0] add_248570;
  wire [7:0] sel_248571;
  wire [7:0] add_248574;
  wire [7:0] sel_248575;
  wire [7:0] add_248578;
  wire [7:0] sel_248579;
  wire [7:0] add_248582;
  wire [7:0] sel_248583;
  wire [7:0] add_248586;
  wire [7:0] sel_248587;
  wire [7:0] add_248590;
  wire [7:0] sel_248591;
  wire [7:0] add_248594;
  wire [7:0] sel_248595;
  wire [7:0] add_248598;
  wire [7:0] sel_248599;
  wire [7:0] add_248602;
  wire [7:0] sel_248603;
  wire [7:0] add_248606;
  wire [7:0] sel_248607;
  wire [7:0] add_248610;
  wire [7:0] sel_248611;
  wire [7:0] add_248614;
  wire [7:0] sel_248615;
  wire [7:0] add_248618;
  wire [7:0] sel_248619;
  wire [7:0] add_248622;
  wire [7:0] sel_248623;
  wire [7:0] add_248626;
  wire [7:0] sel_248627;
  wire [7:0] add_248630;
  wire [7:0] sel_248631;
  wire [7:0] add_248634;
  wire [7:0] sel_248635;
  wire [7:0] add_248638;
  wire [7:0] sel_248639;
  wire [7:0] add_248642;
  wire [7:0] sel_248643;
  wire [7:0] add_248646;
  wire [7:0] sel_248647;
  wire [7:0] add_248650;
  wire [7:0] sel_248651;
  wire [7:0] add_248654;
  wire [7:0] sel_248655;
  wire [7:0] add_248658;
  wire [7:0] sel_248659;
  wire [7:0] add_248662;
  wire [7:0] sel_248663;
  wire [7:0] add_248666;
  wire [7:0] sel_248667;
  wire [7:0] add_248670;
  wire [7:0] sel_248671;
  wire [7:0] add_248674;
  wire [7:0] sel_248675;
  wire [7:0] add_248678;
  wire [7:0] sel_248679;
  wire [7:0] add_248682;
  wire [7:0] sel_248683;
  wire [7:0] add_248686;
  wire [7:0] sel_248687;
  wire [7:0] add_248690;
  wire [7:0] sel_248691;
  wire [7:0] add_248694;
  wire [7:0] sel_248695;
  wire [7:0] add_248698;
  wire [7:0] sel_248699;
  wire [7:0] add_248702;
  wire [7:0] sel_248703;
  wire [7:0] add_248706;
  wire [7:0] sel_248707;
  wire [7:0] add_248711;
  wire [15:0] array_index_248712;
  wire [7:0] sel_248713;
  wire [7:0] add_248716;
  wire [7:0] sel_248717;
  wire [7:0] add_248720;
  wire [7:0] sel_248721;
  wire [7:0] add_248724;
  wire [7:0] sel_248725;
  wire [7:0] add_248728;
  wire [7:0] sel_248729;
  wire [7:0] add_248732;
  wire [7:0] sel_248733;
  wire [7:0] add_248736;
  wire [7:0] sel_248737;
  wire [7:0] add_248740;
  wire [7:0] sel_248741;
  wire [7:0] add_248744;
  wire [7:0] sel_248745;
  wire [7:0] add_248748;
  wire [7:0] sel_248749;
  wire [7:0] add_248752;
  wire [7:0] sel_248753;
  wire [7:0] add_248756;
  wire [7:0] sel_248757;
  wire [7:0] add_248760;
  wire [7:0] sel_248761;
  wire [7:0] add_248764;
  wire [7:0] sel_248765;
  wire [7:0] add_248768;
  wire [7:0] sel_248769;
  wire [7:0] add_248772;
  wire [7:0] sel_248773;
  wire [7:0] add_248776;
  wire [7:0] sel_248777;
  wire [7:0] add_248780;
  wire [7:0] sel_248781;
  wire [7:0] add_248784;
  wire [7:0] sel_248785;
  wire [7:0] add_248788;
  wire [7:0] sel_248789;
  wire [7:0] add_248792;
  wire [7:0] sel_248793;
  wire [7:0] add_248796;
  wire [7:0] sel_248797;
  wire [7:0] add_248800;
  wire [7:0] sel_248801;
  wire [7:0] add_248804;
  wire [7:0] sel_248805;
  wire [7:0] add_248808;
  wire [7:0] sel_248809;
  wire [7:0] add_248812;
  wire [7:0] sel_248813;
  wire [7:0] add_248816;
  wire [7:0] sel_248817;
  wire [7:0] add_248820;
  wire [7:0] sel_248821;
  wire [7:0] add_248824;
  wire [7:0] sel_248825;
  wire [7:0] add_248828;
  wire [7:0] sel_248829;
  wire [7:0] add_248832;
  wire [7:0] sel_248833;
  wire [7:0] add_248836;
  wire [7:0] sel_248837;
  wire [7:0] add_248840;
  wire [7:0] sel_248841;
  wire [7:0] add_248844;
  wire [7:0] sel_248845;
  wire [7:0] add_248848;
  wire [7:0] sel_248849;
  wire [7:0] add_248852;
  wire [7:0] sel_248853;
  wire [7:0] add_248856;
  wire [7:0] sel_248857;
  wire [7:0] add_248860;
  wire [7:0] sel_248861;
  wire [7:0] add_248864;
  wire [7:0] sel_248865;
  wire [7:0] add_248868;
  wire [7:0] sel_248869;
  wire [7:0] add_248872;
  wire [7:0] sel_248873;
  wire [7:0] add_248876;
  wire [7:0] sel_248877;
  wire [7:0] add_248880;
  wire [7:0] sel_248881;
  wire [7:0] add_248884;
  wire [7:0] sel_248885;
  wire [7:0] add_248888;
  wire [7:0] sel_248889;
  wire [7:0] add_248892;
  wire [7:0] sel_248893;
  wire [7:0] add_248896;
  wire [7:0] sel_248897;
  wire [7:0] add_248900;
  wire [7:0] sel_248901;
  wire [7:0] add_248904;
  wire [7:0] sel_248905;
  wire [7:0] add_248908;
  wire [7:0] sel_248909;
  wire [7:0] add_248913;
  wire [15:0] array_index_248914;
  wire [7:0] sel_248915;
  wire [7:0] add_248918;
  wire [7:0] sel_248919;
  wire [7:0] add_248922;
  wire [7:0] sel_248923;
  wire [7:0] add_248926;
  wire [7:0] sel_248927;
  wire [7:0] add_248930;
  wire [7:0] sel_248931;
  wire [7:0] add_248934;
  wire [7:0] sel_248935;
  wire [7:0] add_248938;
  wire [7:0] sel_248939;
  wire [7:0] add_248942;
  wire [7:0] sel_248943;
  wire [7:0] add_248946;
  wire [7:0] sel_248947;
  wire [7:0] add_248950;
  wire [7:0] sel_248951;
  wire [7:0] add_248954;
  wire [7:0] sel_248955;
  wire [7:0] add_248958;
  wire [7:0] sel_248959;
  wire [7:0] add_248962;
  wire [7:0] sel_248963;
  wire [7:0] add_248966;
  wire [7:0] sel_248967;
  wire [7:0] add_248970;
  wire [7:0] sel_248971;
  wire [7:0] add_248974;
  wire [7:0] sel_248975;
  wire [7:0] add_248978;
  wire [7:0] sel_248979;
  wire [7:0] add_248982;
  wire [7:0] sel_248983;
  wire [7:0] add_248986;
  wire [7:0] sel_248987;
  wire [7:0] add_248990;
  wire [7:0] sel_248991;
  wire [7:0] add_248994;
  wire [7:0] sel_248995;
  wire [7:0] add_248998;
  wire [7:0] sel_248999;
  wire [7:0] add_249002;
  wire [7:0] sel_249003;
  wire [7:0] add_249006;
  wire [7:0] sel_249007;
  wire [7:0] add_249010;
  wire [7:0] sel_249011;
  wire [7:0] add_249014;
  wire [7:0] sel_249015;
  wire [7:0] add_249018;
  wire [7:0] sel_249019;
  wire [7:0] add_249022;
  wire [7:0] sel_249023;
  wire [7:0] add_249026;
  wire [7:0] sel_249027;
  wire [7:0] add_249030;
  wire [7:0] sel_249031;
  wire [7:0] add_249034;
  wire [7:0] sel_249035;
  wire [7:0] add_249038;
  wire [7:0] sel_249039;
  wire [7:0] add_249042;
  wire [7:0] sel_249043;
  wire [7:0] add_249046;
  wire [7:0] sel_249047;
  wire [7:0] add_249050;
  wire [7:0] sel_249051;
  wire [7:0] add_249054;
  wire [7:0] sel_249055;
  wire [7:0] add_249058;
  wire [7:0] sel_249059;
  wire [7:0] add_249062;
  wire [7:0] sel_249063;
  wire [7:0] add_249066;
  wire [7:0] sel_249067;
  wire [7:0] add_249070;
  wire [7:0] sel_249071;
  wire [7:0] add_249074;
  wire [7:0] sel_249075;
  wire [7:0] add_249078;
  wire [7:0] sel_249079;
  wire [7:0] add_249082;
  wire [7:0] sel_249083;
  wire [7:0] add_249086;
  wire [7:0] sel_249087;
  wire [7:0] add_249090;
  wire [7:0] sel_249091;
  wire [7:0] add_249094;
  wire [7:0] sel_249095;
  wire [7:0] add_249098;
  wire [7:0] sel_249099;
  wire [7:0] add_249102;
  wire [7:0] sel_249103;
  wire [7:0] add_249106;
  wire [7:0] sel_249107;
  wire [7:0] add_249110;
  wire [7:0] sel_249111;
  wire [7:0] add_249115;
  wire [15:0] array_index_249116;
  wire [7:0] sel_249117;
  wire [7:0] add_249120;
  wire [7:0] sel_249121;
  wire [7:0] add_249124;
  wire [7:0] sel_249125;
  wire [7:0] add_249128;
  wire [7:0] sel_249129;
  wire [7:0] add_249132;
  wire [7:0] sel_249133;
  wire [7:0] add_249136;
  wire [7:0] sel_249137;
  wire [7:0] add_249140;
  wire [7:0] sel_249141;
  wire [7:0] add_249144;
  wire [7:0] sel_249145;
  wire [7:0] add_249148;
  wire [7:0] sel_249149;
  wire [7:0] add_249152;
  wire [7:0] sel_249153;
  wire [7:0] add_249156;
  wire [7:0] sel_249157;
  wire [7:0] add_249160;
  wire [7:0] sel_249161;
  wire [7:0] add_249164;
  wire [7:0] sel_249165;
  wire [7:0] add_249168;
  wire [7:0] sel_249169;
  wire [7:0] add_249172;
  wire [7:0] sel_249173;
  wire [7:0] add_249176;
  wire [7:0] sel_249177;
  wire [7:0] add_249180;
  wire [7:0] sel_249181;
  wire [7:0] add_249184;
  wire [7:0] sel_249185;
  wire [7:0] add_249188;
  wire [7:0] sel_249189;
  wire [7:0] add_249192;
  wire [7:0] sel_249193;
  wire [7:0] add_249196;
  wire [7:0] sel_249197;
  wire [7:0] add_249200;
  wire [7:0] sel_249201;
  wire [7:0] add_249204;
  wire [7:0] sel_249205;
  wire [7:0] add_249208;
  wire [7:0] sel_249209;
  wire [7:0] add_249212;
  wire [7:0] sel_249213;
  wire [7:0] add_249216;
  wire [7:0] sel_249217;
  wire [7:0] add_249220;
  wire [7:0] sel_249221;
  wire [7:0] add_249224;
  wire [7:0] sel_249225;
  wire [7:0] add_249228;
  wire [7:0] sel_249229;
  wire [7:0] add_249232;
  wire [7:0] sel_249233;
  wire [7:0] add_249236;
  wire [7:0] sel_249237;
  wire [7:0] add_249240;
  wire [7:0] sel_249241;
  wire [7:0] add_249244;
  wire [7:0] sel_249245;
  wire [7:0] add_249248;
  wire [7:0] sel_249249;
  wire [7:0] add_249252;
  wire [7:0] sel_249253;
  wire [7:0] add_249256;
  wire [7:0] sel_249257;
  wire [7:0] add_249260;
  wire [7:0] sel_249261;
  wire [7:0] add_249264;
  wire [7:0] sel_249265;
  wire [7:0] add_249268;
  wire [7:0] sel_249269;
  wire [7:0] add_249272;
  wire [7:0] sel_249273;
  wire [7:0] add_249276;
  wire [7:0] sel_249277;
  wire [7:0] add_249280;
  wire [7:0] sel_249281;
  wire [7:0] add_249284;
  wire [7:0] sel_249285;
  wire [7:0] add_249288;
  wire [7:0] sel_249289;
  wire [7:0] add_249292;
  wire [7:0] sel_249293;
  wire [7:0] add_249296;
  wire [7:0] sel_249297;
  wire [7:0] add_249300;
  wire [7:0] sel_249301;
  wire [7:0] add_249304;
  wire [7:0] sel_249305;
  wire [7:0] add_249308;
  wire [7:0] sel_249309;
  wire [7:0] add_249312;
  wire [7:0] sel_249313;
  wire [7:0] add_249317;
  wire [15:0] array_index_249318;
  wire [7:0] sel_249319;
  wire [7:0] add_249322;
  wire [7:0] sel_249323;
  wire [7:0] add_249326;
  wire [7:0] sel_249327;
  wire [7:0] add_249330;
  wire [7:0] sel_249331;
  wire [7:0] add_249334;
  wire [7:0] sel_249335;
  wire [7:0] add_249338;
  wire [7:0] sel_249339;
  wire [7:0] add_249342;
  wire [7:0] sel_249343;
  wire [7:0] add_249346;
  wire [7:0] sel_249347;
  wire [7:0] add_249350;
  wire [7:0] sel_249351;
  wire [7:0] add_249354;
  wire [7:0] sel_249355;
  wire [7:0] add_249358;
  wire [7:0] sel_249359;
  wire [7:0] add_249362;
  wire [7:0] sel_249363;
  wire [7:0] add_249366;
  wire [7:0] sel_249367;
  wire [7:0] add_249370;
  wire [7:0] sel_249371;
  wire [7:0] add_249374;
  wire [7:0] sel_249375;
  wire [7:0] add_249378;
  wire [7:0] sel_249379;
  wire [7:0] add_249382;
  wire [7:0] sel_249383;
  wire [7:0] add_249386;
  wire [7:0] sel_249387;
  wire [7:0] add_249390;
  wire [7:0] sel_249391;
  wire [7:0] add_249394;
  wire [7:0] sel_249395;
  wire [7:0] add_249398;
  wire [7:0] sel_249399;
  wire [7:0] add_249402;
  wire [7:0] sel_249403;
  wire [7:0] add_249406;
  wire [7:0] sel_249407;
  wire [7:0] add_249410;
  wire [7:0] sel_249411;
  wire [7:0] add_249414;
  wire [7:0] sel_249415;
  wire [7:0] add_249418;
  wire [7:0] sel_249419;
  wire [7:0] add_249422;
  wire [7:0] sel_249423;
  wire [7:0] add_249426;
  wire [7:0] sel_249427;
  wire [7:0] add_249430;
  wire [7:0] sel_249431;
  wire [7:0] add_249434;
  wire [7:0] sel_249435;
  wire [7:0] add_249438;
  wire [7:0] sel_249439;
  wire [7:0] add_249442;
  wire [7:0] sel_249443;
  wire [7:0] add_249446;
  wire [7:0] sel_249447;
  wire [7:0] add_249450;
  wire [7:0] sel_249451;
  wire [7:0] add_249454;
  wire [7:0] sel_249455;
  wire [7:0] add_249458;
  wire [7:0] sel_249459;
  wire [7:0] add_249462;
  wire [7:0] sel_249463;
  wire [7:0] add_249466;
  wire [7:0] sel_249467;
  wire [7:0] add_249470;
  wire [7:0] sel_249471;
  wire [7:0] add_249474;
  wire [7:0] sel_249475;
  wire [7:0] add_249478;
  wire [7:0] sel_249479;
  wire [7:0] add_249482;
  wire [7:0] sel_249483;
  wire [7:0] add_249486;
  wire [7:0] sel_249487;
  wire [7:0] add_249490;
  wire [7:0] sel_249491;
  wire [7:0] add_249494;
  wire [7:0] sel_249495;
  wire [7:0] add_249498;
  wire [7:0] sel_249499;
  wire [7:0] add_249502;
  wire [7:0] sel_249503;
  wire [7:0] add_249506;
  wire [7:0] sel_249507;
  wire [7:0] add_249510;
  wire [7:0] sel_249511;
  wire [7:0] add_249514;
  wire [7:0] sel_249515;
  wire [7:0] add_249518;
  assign array_index_239311 = set1_unflattened[6'h00];
  assign array_index_239312 = set2_unflattened[6'h00];
  assign array_index_239316 = set2_unflattened[6'h01];
  assign concat_239317 = {1'h0, array_index_239311 == array_index_239312};
  assign add_239320 = concat_239317 + 2'h1;
  assign array_index_239324 = set2_unflattened[6'h02];
  assign concat_239325 = {1'h0, array_index_239311 == array_index_239316 ? add_239320 : concat_239317};
  assign add_239328 = concat_239325 + 3'h1;
  assign array_index_239332 = set2_unflattened[6'h03];
  assign concat_239333 = {1'h0, array_index_239311 == array_index_239324 ? add_239328 : concat_239325};
  assign add_239336 = concat_239333 + 4'h1;
  assign array_index_239340 = set2_unflattened[6'h04];
  assign concat_239341 = {1'h0, array_index_239311 == array_index_239332 ? add_239336 : concat_239333};
  assign add_239344 = concat_239341 + 5'h01;
  assign array_index_239348 = set2_unflattened[6'h05];
  assign concat_239349 = {1'h0, array_index_239311 == array_index_239340 ? add_239344 : concat_239341};
  assign add_239352 = concat_239349 + 6'h01;
  assign array_index_239356 = set2_unflattened[6'h06];
  assign concat_239357 = {1'h0, array_index_239311 == array_index_239348 ? add_239352 : concat_239349};
  assign add_239360 = concat_239357 + 7'h01;
  assign array_index_239364 = set2_unflattened[6'h07];
  assign concat_239365 = {1'h0, array_index_239311 == array_index_239356 ? add_239360 : concat_239357};
  assign add_239369 = concat_239365 + 8'h01;
  assign array_index_239370 = set2_unflattened[6'h08];
  assign sel_239371 = array_index_239311 == array_index_239364 ? add_239369 : concat_239365;
  assign add_239375 = sel_239371 + 8'h01;
  assign array_index_239376 = set2_unflattened[6'h09];
  assign sel_239377 = array_index_239311 == array_index_239370 ? add_239375 : sel_239371;
  assign add_239381 = sel_239377 + 8'h01;
  assign array_index_239382 = set2_unflattened[6'h0a];
  assign sel_239383 = array_index_239311 == array_index_239376 ? add_239381 : sel_239377;
  assign add_239387 = sel_239383 + 8'h01;
  assign array_index_239388 = set2_unflattened[6'h0b];
  assign sel_239389 = array_index_239311 == array_index_239382 ? add_239387 : sel_239383;
  assign add_239393 = sel_239389 + 8'h01;
  assign array_index_239394 = set2_unflattened[6'h0c];
  assign sel_239395 = array_index_239311 == array_index_239388 ? add_239393 : sel_239389;
  assign add_239399 = sel_239395 + 8'h01;
  assign array_index_239400 = set2_unflattened[6'h0d];
  assign sel_239401 = array_index_239311 == array_index_239394 ? add_239399 : sel_239395;
  assign add_239405 = sel_239401 + 8'h01;
  assign array_index_239406 = set2_unflattened[6'h0e];
  assign sel_239407 = array_index_239311 == array_index_239400 ? add_239405 : sel_239401;
  assign add_239411 = sel_239407 + 8'h01;
  assign array_index_239412 = set2_unflattened[6'h0f];
  assign sel_239413 = array_index_239311 == array_index_239406 ? add_239411 : sel_239407;
  assign add_239417 = sel_239413 + 8'h01;
  assign array_index_239418 = set2_unflattened[6'h10];
  assign sel_239419 = array_index_239311 == array_index_239412 ? add_239417 : sel_239413;
  assign add_239423 = sel_239419 + 8'h01;
  assign array_index_239424 = set2_unflattened[6'h11];
  assign sel_239425 = array_index_239311 == array_index_239418 ? add_239423 : sel_239419;
  assign add_239429 = sel_239425 + 8'h01;
  assign array_index_239430 = set2_unflattened[6'h12];
  assign sel_239431 = array_index_239311 == array_index_239424 ? add_239429 : sel_239425;
  assign add_239435 = sel_239431 + 8'h01;
  assign array_index_239436 = set2_unflattened[6'h13];
  assign sel_239437 = array_index_239311 == array_index_239430 ? add_239435 : sel_239431;
  assign add_239441 = sel_239437 + 8'h01;
  assign array_index_239442 = set2_unflattened[6'h14];
  assign sel_239443 = array_index_239311 == array_index_239436 ? add_239441 : sel_239437;
  assign add_239447 = sel_239443 + 8'h01;
  assign array_index_239448 = set2_unflattened[6'h15];
  assign sel_239449 = array_index_239311 == array_index_239442 ? add_239447 : sel_239443;
  assign add_239453 = sel_239449 + 8'h01;
  assign array_index_239454 = set2_unflattened[6'h16];
  assign sel_239455 = array_index_239311 == array_index_239448 ? add_239453 : sel_239449;
  assign add_239459 = sel_239455 + 8'h01;
  assign array_index_239460 = set2_unflattened[6'h17];
  assign sel_239461 = array_index_239311 == array_index_239454 ? add_239459 : sel_239455;
  assign add_239465 = sel_239461 + 8'h01;
  assign array_index_239466 = set2_unflattened[6'h18];
  assign sel_239467 = array_index_239311 == array_index_239460 ? add_239465 : sel_239461;
  assign add_239471 = sel_239467 + 8'h01;
  assign array_index_239472 = set2_unflattened[6'h19];
  assign sel_239473 = array_index_239311 == array_index_239466 ? add_239471 : sel_239467;
  assign add_239477 = sel_239473 + 8'h01;
  assign array_index_239478 = set2_unflattened[6'h1a];
  assign sel_239479 = array_index_239311 == array_index_239472 ? add_239477 : sel_239473;
  assign add_239483 = sel_239479 + 8'h01;
  assign array_index_239484 = set2_unflattened[6'h1b];
  assign sel_239485 = array_index_239311 == array_index_239478 ? add_239483 : sel_239479;
  assign add_239489 = sel_239485 + 8'h01;
  assign array_index_239490 = set2_unflattened[6'h1c];
  assign sel_239491 = array_index_239311 == array_index_239484 ? add_239489 : sel_239485;
  assign add_239495 = sel_239491 + 8'h01;
  assign array_index_239496 = set2_unflattened[6'h1d];
  assign sel_239497 = array_index_239311 == array_index_239490 ? add_239495 : sel_239491;
  assign add_239501 = sel_239497 + 8'h01;
  assign array_index_239502 = set2_unflattened[6'h1e];
  assign sel_239503 = array_index_239311 == array_index_239496 ? add_239501 : sel_239497;
  assign add_239507 = sel_239503 + 8'h01;
  assign array_index_239508 = set2_unflattened[6'h1f];
  assign sel_239509 = array_index_239311 == array_index_239502 ? add_239507 : sel_239503;
  assign add_239513 = sel_239509 + 8'h01;
  assign array_index_239514 = set2_unflattened[6'h20];
  assign sel_239515 = array_index_239311 == array_index_239508 ? add_239513 : sel_239509;
  assign add_239519 = sel_239515 + 8'h01;
  assign array_index_239520 = set2_unflattened[6'h21];
  assign sel_239521 = array_index_239311 == array_index_239514 ? add_239519 : sel_239515;
  assign add_239525 = sel_239521 + 8'h01;
  assign array_index_239526 = set2_unflattened[6'h22];
  assign sel_239527 = array_index_239311 == array_index_239520 ? add_239525 : sel_239521;
  assign add_239531 = sel_239527 + 8'h01;
  assign array_index_239532 = set2_unflattened[6'h23];
  assign sel_239533 = array_index_239311 == array_index_239526 ? add_239531 : sel_239527;
  assign add_239537 = sel_239533 + 8'h01;
  assign array_index_239538 = set2_unflattened[6'h24];
  assign sel_239539 = array_index_239311 == array_index_239532 ? add_239537 : sel_239533;
  assign add_239543 = sel_239539 + 8'h01;
  assign array_index_239544 = set2_unflattened[6'h25];
  assign sel_239545 = array_index_239311 == array_index_239538 ? add_239543 : sel_239539;
  assign add_239549 = sel_239545 + 8'h01;
  assign array_index_239550 = set2_unflattened[6'h26];
  assign sel_239551 = array_index_239311 == array_index_239544 ? add_239549 : sel_239545;
  assign add_239555 = sel_239551 + 8'h01;
  assign array_index_239556 = set2_unflattened[6'h27];
  assign sel_239557 = array_index_239311 == array_index_239550 ? add_239555 : sel_239551;
  assign add_239561 = sel_239557 + 8'h01;
  assign array_index_239562 = set2_unflattened[6'h28];
  assign sel_239563 = array_index_239311 == array_index_239556 ? add_239561 : sel_239557;
  assign add_239567 = sel_239563 + 8'h01;
  assign array_index_239568 = set2_unflattened[6'h29];
  assign sel_239569 = array_index_239311 == array_index_239562 ? add_239567 : sel_239563;
  assign add_239573 = sel_239569 + 8'h01;
  assign array_index_239574 = set2_unflattened[6'h2a];
  assign sel_239575 = array_index_239311 == array_index_239568 ? add_239573 : sel_239569;
  assign add_239579 = sel_239575 + 8'h01;
  assign array_index_239580 = set2_unflattened[6'h2b];
  assign sel_239581 = array_index_239311 == array_index_239574 ? add_239579 : sel_239575;
  assign add_239585 = sel_239581 + 8'h01;
  assign array_index_239586 = set2_unflattened[6'h2c];
  assign sel_239587 = array_index_239311 == array_index_239580 ? add_239585 : sel_239581;
  assign add_239591 = sel_239587 + 8'h01;
  assign array_index_239592 = set2_unflattened[6'h2d];
  assign sel_239593 = array_index_239311 == array_index_239586 ? add_239591 : sel_239587;
  assign add_239597 = sel_239593 + 8'h01;
  assign array_index_239598 = set2_unflattened[6'h2e];
  assign sel_239599 = array_index_239311 == array_index_239592 ? add_239597 : sel_239593;
  assign add_239603 = sel_239599 + 8'h01;
  assign array_index_239604 = set2_unflattened[6'h2f];
  assign sel_239605 = array_index_239311 == array_index_239598 ? add_239603 : sel_239599;
  assign add_239609 = sel_239605 + 8'h01;
  assign array_index_239610 = set2_unflattened[6'h30];
  assign sel_239611 = array_index_239311 == array_index_239604 ? add_239609 : sel_239605;
  assign add_239615 = sel_239611 + 8'h01;
  assign array_index_239616 = set2_unflattened[6'h31];
  assign sel_239617 = array_index_239311 == array_index_239610 ? add_239615 : sel_239611;
  assign add_239621 = sel_239617 + 8'h01;
  assign array_index_239622 = set1_unflattened[6'h01];
  assign sel_239623 = array_index_239311 == array_index_239616 ? add_239621 : sel_239617;
  assign add_239626 = sel_239623 + 8'h01;
  assign sel_239627 = array_index_239622 == array_index_239312 ? add_239626 : sel_239623;
  assign add_239630 = sel_239627 + 8'h01;
  assign sel_239631 = array_index_239622 == array_index_239316 ? add_239630 : sel_239627;
  assign add_239634 = sel_239631 + 8'h01;
  assign sel_239635 = array_index_239622 == array_index_239324 ? add_239634 : sel_239631;
  assign add_239638 = sel_239635 + 8'h01;
  assign sel_239639 = array_index_239622 == array_index_239332 ? add_239638 : sel_239635;
  assign add_239642 = sel_239639 + 8'h01;
  assign sel_239643 = array_index_239622 == array_index_239340 ? add_239642 : sel_239639;
  assign add_239646 = sel_239643 + 8'h01;
  assign sel_239647 = array_index_239622 == array_index_239348 ? add_239646 : sel_239643;
  assign add_239650 = sel_239647 + 8'h01;
  assign sel_239651 = array_index_239622 == array_index_239356 ? add_239650 : sel_239647;
  assign add_239654 = sel_239651 + 8'h01;
  assign sel_239655 = array_index_239622 == array_index_239364 ? add_239654 : sel_239651;
  assign add_239658 = sel_239655 + 8'h01;
  assign sel_239659 = array_index_239622 == array_index_239370 ? add_239658 : sel_239655;
  assign add_239662 = sel_239659 + 8'h01;
  assign sel_239663 = array_index_239622 == array_index_239376 ? add_239662 : sel_239659;
  assign add_239666 = sel_239663 + 8'h01;
  assign sel_239667 = array_index_239622 == array_index_239382 ? add_239666 : sel_239663;
  assign add_239670 = sel_239667 + 8'h01;
  assign sel_239671 = array_index_239622 == array_index_239388 ? add_239670 : sel_239667;
  assign add_239674 = sel_239671 + 8'h01;
  assign sel_239675 = array_index_239622 == array_index_239394 ? add_239674 : sel_239671;
  assign add_239678 = sel_239675 + 8'h01;
  assign sel_239679 = array_index_239622 == array_index_239400 ? add_239678 : sel_239675;
  assign add_239682 = sel_239679 + 8'h01;
  assign sel_239683 = array_index_239622 == array_index_239406 ? add_239682 : sel_239679;
  assign add_239686 = sel_239683 + 8'h01;
  assign sel_239687 = array_index_239622 == array_index_239412 ? add_239686 : sel_239683;
  assign add_239690 = sel_239687 + 8'h01;
  assign sel_239691 = array_index_239622 == array_index_239418 ? add_239690 : sel_239687;
  assign add_239694 = sel_239691 + 8'h01;
  assign sel_239695 = array_index_239622 == array_index_239424 ? add_239694 : sel_239691;
  assign add_239698 = sel_239695 + 8'h01;
  assign sel_239699 = array_index_239622 == array_index_239430 ? add_239698 : sel_239695;
  assign add_239702 = sel_239699 + 8'h01;
  assign sel_239703 = array_index_239622 == array_index_239436 ? add_239702 : sel_239699;
  assign add_239706 = sel_239703 + 8'h01;
  assign sel_239707 = array_index_239622 == array_index_239442 ? add_239706 : sel_239703;
  assign add_239710 = sel_239707 + 8'h01;
  assign sel_239711 = array_index_239622 == array_index_239448 ? add_239710 : sel_239707;
  assign add_239714 = sel_239711 + 8'h01;
  assign sel_239715 = array_index_239622 == array_index_239454 ? add_239714 : sel_239711;
  assign add_239718 = sel_239715 + 8'h01;
  assign sel_239719 = array_index_239622 == array_index_239460 ? add_239718 : sel_239715;
  assign add_239722 = sel_239719 + 8'h01;
  assign sel_239723 = array_index_239622 == array_index_239466 ? add_239722 : sel_239719;
  assign add_239726 = sel_239723 + 8'h01;
  assign sel_239727 = array_index_239622 == array_index_239472 ? add_239726 : sel_239723;
  assign add_239730 = sel_239727 + 8'h01;
  assign sel_239731 = array_index_239622 == array_index_239478 ? add_239730 : sel_239727;
  assign add_239734 = sel_239731 + 8'h01;
  assign sel_239735 = array_index_239622 == array_index_239484 ? add_239734 : sel_239731;
  assign add_239738 = sel_239735 + 8'h01;
  assign sel_239739 = array_index_239622 == array_index_239490 ? add_239738 : sel_239735;
  assign add_239742 = sel_239739 + 8'h01;
  assign sel_239743 = array_index_239622 == array_index_239496 ? add_239742 : sel_239739;
  assign add_239746 = sel_239743 + 8'h01;
  assign sel_239747 = array_index_239622 == array_index_239502 ? add_239746 : sel_239743;
  assign add_239750 = sel_239747 + 8'h01;
  assign sel_239751 = array_index_239622 == array_index_239508 ? add_239750 : sel_239747;
  assign add_239754 = sel_239751 + 8'h01;
  assign sel_239755 = array_index_239622 == array_index_239514 ? add_239754 : sel_239751;
  assign add_239758 = sel_239755 + 8'h01;
  assign sel_239759 = array_index_239622 == array_index_239520 ? add_239758 : sel_239755;
  assign add_239762 = sel_239759 + 8'h01;
  assign sel_239763 = array_index_239622 == array_index_239526 ? add_239762 : sel_239759;
  assign add_239766 = sel_239763 + 8'h01;
  assign sel_239767 = array_index_239622 == array_index_239532 ? add_239766 : sel_239763;
  assign add_239770 = sel_239767 + 8'h01;
  assign sel_239771 = array_index_239622 == array_index_239538 ? add_239770 : sel_239767;
  assign add_239774 = sel_239771 + 8'h01;
  assign sel_239775 = array_index_239622 == array_index_239544 ? add_239774 : sel_239771;
  assign add_239778 = sel_239775 + 8'h01;
  assign sel_239779 = array_index_239622 == array_index_239550 ? add_239778 : sel_239775;
  assign add_239782 = sel_239779 + 8'h01;
  assign sel_239783 = array_index_239622 == array_index_239556 ? add_239782 : sel_239779;
  assign add_239786 = sel_239783 + 8'h01;
  assign sel_239787 = array_index_239622 == array_index_239562 ? add_239786 : sel_239783;
  assign add_239790 = sel_239787 + 8'h01;
  assign sel_239791 = array_index_239622 == array_index_239568 ? add_239790 : sel_239787;
  assign add_239794 = sel_239791 + 8'h01;
  assign sel_239795 = array_index_239622 == array_index_239574 ? add_239794 : sel_239791;
  assign add_239798 = sel_239795 + 8'h01;
  assign sel_239799 = array_index_239622 == array_index_239580 ? add_239798 : sel_239795;
  assign add_239802 = sel_239799 + 8'h01;
  assign sel_239803 = array_index_239622 == array_index_239586 ? add_239802 : sel_239799;
  assign add_239806 = sel_239803 + 8'h01;
  assign sel_239807 = array_index_239622 == array_index_239592 ? add_239806 : sel_239803;
  assign add_239810 = sel_239807 + 8'h01;
  assign sel_239811 = array_index_239622 == array_index_239598 ? add_239810 : sel_239807;
  assign add_239814 = sel_239811 + 8'h01;
  assign sel_239815 = array_index_239622 == array_index_239604 ? add_239814 : sel_239811;
  assign add_239818 = sel_239815 + 8'h01;
  assign sel_239819 = array_index_239622 == array_index_239610 ? add_239818 : sel_239815;
  assign add_239823 = sel_239819 + 8'h01;
  assign array_index_239824 = set1_unflattened[6'h02];
  assign sel_239825 = array_index_239622 == array_index_239616 ? add_239823 : sel_239819;
  assign add_239828 = sel_239825 + 8'h01;
  assign sel_239829 = array_index_239824 == array_index_239312 ? add_239828 : sel_239825;
  assign add_239832 = sel_239829 + 8'h01;
  assign sel_239833 = array_index_239824 == array_index_239316 ? add_239832 : sel_239829;
  assign add_239836 = sel_239833 + 8'h01;
  assign sel_239837 = array_index_239824 == array_index_239324 ? add_239836 : sel_239833;
  assign add_239840 = sel_239837 + 8'h01;
  assign sel_239841 = array_index_239824 == array_index_239332 ? add_239840 : sel_239837;
  assign add_239844 = sel_239841 + 8'h01;
  assign sel_239845 = array_index_239824 == array_index_239340 ? add_239844 : sel_239841;
  assign add_239848 = sel_239845 + 8'h01;
  assign sel_239849 = array_index_239824 == array_index_239348 ? add_239848 : sel_239845;
  assign add_239852 = sel_239849 + 8'h01;
  assign sel_239853 = array_index_239824 == array_index_239356 ? add_239852 : sel_239849;
  assign add_239856 = sel_239853 + 8'h01;
  assign sel_239857 = array_index_239824 == array_index_239364 ? add_239856 : sel_239853;
  assign add_239860 = sel_239857 + 8'h01;
  assign sel_239861 = array_index_239824 == array_index_239370 ? add_239860 : sel_239857;
  assign add_239864 = sel_239861 + 8'h01;
  assign sel_239865 = array_index_239824 == array_index_239376 ? add_239864 : sel_239861;
  assign add_239868 = sel_239865 + 8'h01;
  assign sel_239869 = array_index_239824 == array_index_239382 ? add_239868 : sel_239865;
  assign add_239872 = sel_239869 + 8'h01;
  assign sel_239873 = array_index_239824 == array_index_239388 ? add_239872 : sel_239869;
  assign add_239876 = sel_239873 + 8'h01;
  assign sel_239877 = array_index_239824 == array_index_239394 ? add_239876 : sel_239873;
  assign add_239880 = sel_239877 + 8'h01;
  assign sel_239881 = array_index_239824 == array_index_239400 ? add_239880 : sel_239877;
  assign add_239884 = sel_239881 + 8'h01;
  assign sel_239885 = array_index_239824 == array_index_239406 ? add_239884 : sel_239881;
  assign add_239888 = sel_239885 + 8'h01;
  assign sel_239889 = array_index_239824 == array_index_239412 ? add_239888 : sel_239885;
  assign add_239892 = sel_239889 + 8'h01;
  assign sel_239893 = array_index_239824 == array_index_239418 ? add_239892 : sel_239889;
  assign add_239896 = sel_239893 + 8'h01;
  assign sel_239897 = array_index_239824 == array_index_239424 ? add_239896 : sel_239893;
  assign add_239900 = sel_239897 + 8'h01;
  assign sel_239901 = array_index_239824 == array_index_239430 ? add_239900 : sel_239897;
  assign add_239904 = sel_239901 + 8'h01;
  assign sel_239905 = array_index_239824 == array_index_239436 ? add_239904 : sel_239901;
  assign add_239908 = sel_239905 + 8'h01;
  assign sel_239909 = array_index_239824 == array_index_239442 ? add_239908 : sel_239905;
  assign add_239912 = sel_239909 + 8'h01;
  assign sel_239913 = array_index_239824 == array_index_239448 ? add_239912 : sel_239909;
  assign add_239916 = sel_239913 + 8'h01;
  assign sel_239917 = array_index_239824 == array_index_239454 ? add_239916 : sel_239913;
  assign add_239920 = sel_239917 + 8'h01;
  assign sel_239921 = array_index_239824 == array_index_239460 ? add_239920 : sel_239917;
  assign add_239924 = sel_239921 + 8'h01;
  assign sel_239925 = array_index_239824 == array_index_239466 ? add_239924 : sel_239921;
  assign add_239928 = sel_239925 + 8'h01;
  assign sel_239929 = array_index_239824 == array_index_239472 ? add_239928 : sel_239925;
  assign add_239932 = sel_239929 + 8'h01;
  assign sel_239933 = array_index_239824 == array_index_239478 ? add_239932 : sel_239929;
  assign add_239936 = sel_239933 + 8'h01;
  assign sel_239937 = array_index_239824 == array_index_239484 ? add_239936 : sel_239933;
  assign add_239940 = sel_239937 + 8'h01;
  assign sel_239941 = array_index_239824 == array_index_239490 ? add_239940 : sel_239937;
  assign add_239944 = sel_239941 + 8'h01;
  assign sel_239945 = array_index_239824 == array_index_239496 ? add_239944 : sel_239941;
  assign add_239948 = sel_239945 + 8'h01;
  assign sel_239949 = array_index_239824 == array_index_239502 ? add_239948 : sel_239945;
  assign add_239952 = sel_239949 + 8'h01;
  assign sel_239953 = array_index_239824 == array_index_239508 ? add_239952 : sel_239949;
  assign add_239956 = sel_239953 + 8'h01;
  assign sel_239957 = array_index_239824 == array_index_239514 ? add_239956 : sel_239953;
  assign add_239960 = sel_239957 + 8'h01;
  assign sel_239961 = array_index_239824 == array_index_239520 ? add_239960 : sel_239957;
  assign add_239964 = sel_239961 + 8'h01;
  assign sel_239965 = array_index_239824 == array_index_239526 ? add_239964 : sel_239961;
  assign add_239968 = sel_239965 + 8'h01;
  assign sel_239969 = array_index_239824 == array_index_239532 ? add_239968 : sel_239965;
  assign add_239972 = sel_239969 + 8'h01;
  assign sel_239973 = array_index_239824 == array_index_239538 ? add_239972 : sel_239969;
  assign add_239976 = sel_239973 + 8'h01;
  assign sel_239977 = array_index_239824 == array_index_239544 ? add_239976 : sel_239973;
  assign add_239980 = sel_239977 + 8'h01;
  assign sel_239981 = array_index_239824 == array_index_239550 ? add_239980 : sel_239977;
  assign add_239984 = sel_239981 + 8'h01;
  assign sel_239985 = array_index_239824 == array_index_239556 ? add_239984 : sel_239981;
  assign add_239988 = sel_239985 + 8'h01;
  assign sel_239989 = array_index_239824 == array_index_239562 ? add_239988 : sel_239985;
  assign add_239992 = sel_239989 + 8'h01;
  assign sel_239993 = array_index_239824 == array_index_239568 ? add_239992 : sel_239989;
  assign add_239996 = sel_239993 + 8'h01;
  assign sel_239997 = array_index_239824 == array_index_239574 ? add_239996 : sel_239993;
  assign add_240000 = sel_239997 + 8'h01;
  assign sel_240001 = array_index_239824 == array_index_239580 ? add_240000 : sel_239997;
  assign add_240004 = sel_240001 + 8'h01;
  assign sel_240005 = array_index_239824 == array_index_239586 ? add_240004 : sel_240001;
  assign add_240008 = sel_240005 + 8'h01;
  assign sel_240009 = array_index_239824 == array_index_239592 ? add_240008 : sel_240005;
  assign add_240012 = sel_240009 + 8'h01;
  assign sel_240013 = array_index_239824 == array_index_239598 ? add_240012 : sel_240009;
  assign add_240016 = sel_240013 + 8'h01;
  assign sel_240017 = array_index_239824 == array_index_239604 ? add_240016 : sel_240013;
  assign add_240020 = sel_240017 + 8'h01;
  assign sel_240021 = array_index_239824 == array_index_239610 ? add_240020 : sel_240017;
  assign add_240025 = sel_240021 + 8'h01;
  assign array_index_240026 = set1_unflattened[6'h03];
  assign sel_240027 = array_index_239824 == array_index_239616 ? add_240025 : sel_240021;
  assign add_240030 = sel_240027 + 8'h01;
  assign sel_240031 = array_index_240026 == array_index_239312 ? add_240030 : sel_240027;
  assign add_240034 = sel_240031 + 8'h01;
  assign sel_240035 = array_index_240026 == array_index_239316 ? add_240034 : sel_240031;
  assign add_240038 = sel_240035 + 8'h01;
  assign sel_240039 = array_index_240026 == array_index_239324 ? add_240038 : sel_240035;
  assign add_240042 = sel_240039 + 8'h01;
  assign sel_240043 = array_index_240026 == array_index_239332 ? add_240042 : sel_240039;
  assign add_240046 = sel_240043 + 8'h01;
  assign sel_240047 = array_index_240026 == array_index_239340 ? add_240046 : sel_240043;
  assign add_240050 = sel_240047 + 8'h01;
  assign sel_240051 = array_index_240026 == array_index_239348 ? add_240050 : sel_240047;
  assign add_240054 = sel_240051 + 8'h01;
  assign sel_240055 = array_index_240026 == array_index_239356 ? add_240054 : sel_240051;
  assign add_240058 = sel_240055 + 8'h01;
  assign sel_240059 = array_index_240026 == array_index_239364 ? add_240058 : sel_240055;
  assign add_240062 = sel_240059 + 8'h01;
  assign sel_240063 = array_index_240026 == array_index_239370 ? add_240062 : sel_240059;
  assign add_240066 = sel_240063 + 8'h01;
  assign sel_240067 = array_index_240026 == array_index_239376 ? add_240066 : sel_240063;
  assign add_240070 = sel_240067 + 8'h01;
  assign sel_240071 = array_index_240026 == array_index_239382 ? add_240070 : sel_240067;
  assign add_240074 = sel_240071 + 8'h01;
  assign sel_240075 = array_index_240026 == array_index_239388 ? add_240074 : sel_240071;
  assign add_240078 = sel_240075 + 8'h01;
  assign sel_240079 = array_index_240026 == array_index_239394 ? add_240078 : sel_240075;
  assign add_240082 = sel_240079 + 8'h01;
  assign sel_240083 = array_index_240026 == array_index_239400 ? add_240082 : sel_240079;
  assign add_240086 = sel_240083 + 8'h01;
  assign sel_240087 = array_index_240026 == array_index_239406 ? add_240086 : sel_240083;
  assign add_240090 = sel_240087 + 8'h01;
  assign sel_240091 = array_index_240026 == array_index_239412 ? add_240090 : sel_240087;
  assign add_240094 = sel_240091 + 8'h01;
  assign sel_240095 = array_index_240026 == array_index_239418 ? add_240094 : sel_240091;
  assign add_240098 = sel_240095 + 8'h01;
  assign sel_240099 = array_index_240026 == array_index_239424 ? add_240098 : sel_240095;
  assign add_240102 = sel_240099 + 8'h01;
  assign sel_240103 = array_index_240026 == array_index_239430 ? add_240102 : sel_240099;
  assign add_240106 = sel_240103 + 8'h01;
  assign sel_240107 = array_index_240026 == array_index_239436 ? add_240106 : sel_240103;
  assign add_240110 = sel_240107 + 8'h01;
  assign sel_240111 = array_index_240026 == array_index_239442 ? add_240110 : sel_240107;
  assign add_240114 = sel_240111 + 8'h01;
  assign sel_240115 = array_index_240026 == array_index_239448 ? add_240114 : sel_240111;
  assign add_240118 = sel_240115 + 8'h01;
  assign sel_240119 = array_index_240026 == array_index_239454 ? add_240118 : sel_240115;
  assign add_240122 = sel_240119 + 8'h01;
  assign sel_240123 = array_index_240026 == array_index_239460 ? add_240122 : sel_240119;
  assign add_240126 = sel_240123 + 8'h01;
  assign sel_240127 = array_index_240026 == array_index_239466 ? add_240126 : sel_240123;
  assign add_240130 = sel_240127 + 8'h01;
  assign sel_240131 = array_index_240026 == array_index_239472 ? add_240130 : sel_240127;
  assign add_240134 = sel_240131 + 8'h01;
  assign sel_240135 = array_index_240026 == array_index_239478 ? add_240134 : sel_240131;
  assign add_240138 = sel_240135 + 8'h01;
  assign sel_240139 = array_index_240026 == array_index_239484 ? add_240138 : sel_240135;
  assign add_240142 = sel_240139 + 8'h01;
  assign sel_240143 = array_index_240026 == array_index_239490 ? add_240142 : sel_240139;
  assign add_240146 = sel_240143 + 8'h01;
  assign sel_240147 = array_index_240026 == array_index_239496 ? add_240146 : sel_240143;
  assign add_240150 = sel_240147 + 8'h01;
  assign sel_240151 = array_index_240026 == array_index_239502 ? add_240150 : sel_240147;
  assign add_240154 = sel_240151 + 8'h01;
  assign sel_240155 = array_index_240026 == array_index_239508 ? add_240154 : sel_240151;
  assign add_240158 = sel_240155 + 8'h01;
  assign sel_240159 = array_index_240026 == array_index_239514 ? add_240158 : sel_240155;
  assign add_240162 = sel_240159 + 8'h01;
  assign sel_240163 = array_index_240026 == array_index_239520 ? add_240162 : sel_240159;
  assign add_240166 = sel_240163 + 8'h01;
  assign sel_240167 = array_index_240026 == array_index_239526 ? add_240166 : sel_240163;
  assign add_240170 = sel_240167 + 8'h01;
  assign sel_240171 = array_index_240026 == array_index_239532 ? add_240170 : sel_240167;
  assign add_240174 = sel_240171 + 8'h01;
  assign sel_240175 = array_index_240026 == array_index_239538 ? add_240174 : sel_240171;
  assign add_240178 = sel_240175 + 8'h01;
  assign sel_240179 = array_index_240026 == array_index_239544 ? add_240178 : sel_240175;
  assign add_240182 = sel_240179 + 8'h01;
  assign sel_240183 = array_index_240026 == array_index_239550 ? add_240182 : sel_240179;
  assign add_240186 = sel_240183 + 8'h01;
  assign sel_240187 = array_index_240026 == array_index_239556 ? add_240186 : sel_240183;
  assign add_240190 = sel_240187 + 8'h01;
  assign sel_240191 = array_index_240026 == array_index_239562 ? add_240190 : sel_240187;
  assign add_240194 = sel_240191 + 8'h01;
  assign sel_240195 = array_index_240026 == array_index_239568 ? add_240194 : sel_240191;
  assign add_240198 = sel_240195 + 8'h01;
  assign sel_240199 = array_index_240026 == array_index_239574 ? add_240198 : sel_240195;
  assign add_240202 = sel_240199 + 8'h01;
  assign sel_240203 = array_index_240026 == array_index_239580 ? add_240202 : sel_240199;
  assign add_240206 = sel_240203 + 8'h01;
  assign sel_240207 = array_index_240026 == array_index_239586 ? add_240206 : sel_240203;
  assign add_240210 = sel_240207 + 8'h01;
  assign sel_240211 = array_index_240026 == array_index_239592 ? add_240210 : sel_240207;
  assign add_240214 = sel_240211 + 8'h01;
  assign sel_240215 = array_index_240026 == array_index_239598 ? add_240214 : sel_240211;
  assign add_240218 = sel_240215 + 8'h01;
  assign sel_240219 = array_index_240026 == array_index_239604 ? add_240218 : sel_240215;
  assign add_240222 = sel_240219 + 8'h01;
  assign sel_240223 = array_index_240026 == array_index_239610 ? add_240222 : sel_240219;
  assign add_240227 = sel_240223 + 8'h01;
  assign array_index_240228 = set1_unflattened[6'h04];
  assign sel_240229 = array_index_240026 == array_index_239616 ? add_240227 : sel_240223;
  assign add_240232 = sel_240229 + 8'h01;
  assign sel_240233 = array_index_240228 == array_index_239312 ? add_240232 : sel_240229;
  assign add_240236 = sel_240233 + 8'h01;
  assign sel_240237 = array_index_240228 == array_index_239316 ? add_240236 : sel_240233;
  assign add_240240 = sel_240237 + 8'h01;
  assign sel_240241 = array_index_240228 == array_index_239324 ? add_240240 : sel_240237;
  assign add_240244 = sel_240241 + 8'h01;
  assign sel_240245 = array_index_240228 == array_index_239332 ? add_240244 : sel_240241;
  assign add_240248 = sel_240245 + 8'h01;
  assign sel_240249 = array_index_240228 == array_index_239340 ? add_240248 : sel_240245;
  assign add_240252 = sel_240249 + 8'h01;
  assign sel_240253 = array_index_240228 == array_index_239348 ? add_240252 : sel_240249;
  assign add_240256 = sel_240253 + 8'h01;
  assign sel_240257 = array_index_240228 == array_index_239356 ? add_240256 : sel_240253;
  assign add_240260 = sel_240257 + 8'h01;
  assign sel_240261 = array_index_240228 == array_index_239364 ? add_240260 : sel_240257;
  assign add_240264 = sel_240261 + 8'h01;
  assign sel_240265 = array_index_240228 == array_index_239370 ? add_240264 : sel_240261;
  assign add_240268 = sel_240265 + 8'h01;
  assign sel_240269 = array_index_240228 == array_index_239376 ? add_240268 : sel_240265;
  assign add_240272 = sel_240269 + 8'h01;
  assign sel_240273 = array_index_240228 == array_index_239382 ? add_240272 : sel_240269;
  assign add_240276 = sel_240273 + 8'h01;
  assign sel_240277 = array_index_240228 == array_index_239388 ? add_240276 : sel_240273;
  assign add_240280 = sel_240277 + 8'h01;
  assign sel_240281 = array_index_240228 == array_index_239394 ? add_240280 : sel_240277;
  assign add_240284 = sel_240281 + 8'h01;
  assign sel_240285 = array_index_240228 == array_index_239400 ? add_240284 : sel_240281;
  assign add_240288 = sel_240285 + 8'h01;
  assign sel_240289 = array_index_240228 == array_index_239406 ? add_240288 : sel_240285;
  assign add_240292 = sel_240289 + 8'h01;
  assign sel_240293 = array_index_240228 == array_index_239412 ? add_240292 : sel_240289;
  assign add_240296 = sel_240293 + 8'h01;
  assign sel_240297 = array_index_240228 == array_index_239418 ? add_240296 : sel_240293;
  assign add_240300 = sel_240297 + 8'h01;
  assign sel_240301 = array_index_240228 == array_index_239424 ? add_240300 : sel_240297;
  assign add_240304 = sel_240301 + 8'h01;
  assign sel_240305 = array_index_240228 == array_index_239430 ? add_240304 : sel_240301;
  assign add_240308 = sel_240305 + 8'h01;
  assign sel_240309 = array_index_240228 == array_index_239436 ? add_240308 : sel_240305;
  assign add_240312 = sel_240309 + 8'h01;
  assign sel_240313 = array_index_240228 == array_index_239442 ? add_240312 : sel_240309;
  assign add_240316 = sel_240313 + 8'h01;
  assign sel_240317 = array_index_240228 == array_index_239448 ? add_240316 : sel_240313;
  assign add_240320 = sel_240317 + 8'h01;
  assign sel_240321 = array_index_240228 == array_index_239454 ? add_240320 : sel_240317;
  assign add_240324 = sel_240321 + 8'h01;
  assign sel_240325 = array_index_240228 == array_index_239460 ? add_240324 : sel_240321;
  assign add_240328 = sel_240325 + 8'h01;
  assign sel_240329 = array_index_240228 == array_index_239466 ? add_240328 : sel_240325;
  assign add_240332 = sel_240329 + 8'h01;
  assign sel_240333 = array_index_240228 == array_index_239472 ? add_240332 : sel_240329;
  assign add_240336 = sel_240333 + 8'h01;
  assign sel_240337 = array_index_240228 == array_index_239478 ? add_240336 : sel_240333;
  assign add_240340 = sel_240337 + 8'h01;
  assign sel_240341 = array_index_240228 == array_index_239484 ? add_240340 : sel_240337;
  assign add_240344 = sel_240341 + 8'h01;
  assign sel_240345 = array_index_240228 == array_index_239490 ? add_240344 : sel_240341;
  assign add_240348 = sel_240345 + 8'h01;
  assign sel_240349 = array_index_240228 == array_index_239496 ? add_240348 : sel_240345;
  assign add_240352 = sel_240349 + 8'h01;
  assign sel_240353 = array_index_240228 == array_index_239502 ? add_240352 : sel_240349;
  assign add_240356 = sel_240353 + 8'h01;
  assign sel_240357 = array_index_240228 == array_index_239508 ? add_240356 : sel_240353;
  assign add_240360 = sel_240357 + 8'h01;
  assign sel_240361 = array_index_240228 == array_index_239514 ? add_240360 : sel_240357;
  assign add_240364 = sel_240361 + 8'h01;
  assign sel_240365 = array_index_240228 == array_index_239520 ? add_240364 : sel_240361;
  assign add_240368 = sel_240365 + 8'h01;
  assign sel_240369 = array_index_240228 == array_index_239526 ? add_240368 : sel_240365;
  assign add_240372 = sel_240369 + 8'h01;
  assign sel_240373 = array_index_240228 == array_index_239532 ? add_240372 : sel_240369;
  assign add_240376 = sel_240373 + 8'h01;
  assign sel_240377 = array_index_240228 == array_index_239538 ? add_240376 : sel_240373;
  assign add_240380 = sel_240377 + 8'h01;
  assign sel_240381 = array_index_240228 == array_index_239544 ? add_240380 : sel_240377;
  assign add_240384 = sel_240381 + 8'h01;
  assign sel_240385 = array_index_240228 == array_index_239550 ? add_240384 : sel_240381;
  assign add_240388 = sel_240385 + 8'h01;
  assign sel_240389 = array_index_240228 == array_index_239556 ? add_240388 : sel_240385;
  assign add_240392 = sel_240389 + 8'h01;
  assign sel_240393 = array_index_240228 == array_index_239562 ? add_240392 : sel_240389;
  assign add_240396 = sel_240393 + 8'h01;
  assign sel_240397 = array_index_240228 == array_index_239568 ? add_240396 : sel_240393;
  assign add_240400 = sel_240397 + 8'h01;
  assign sel_240401 = array_index_240228 == array_index_239574 ? add_240400 : sel_240397;
  assign add_240404 = sel_240401 + 8'h01;
  assign sel_240405 = array_index_240228 == array_index_239580 ? add_240404 : sel_240401;
  assign add_240408 = sel_240405 + 8'h01;
  assign sel_240409 = array_index_240228 == array_index_239586 ? add_240408 : sel_240405;
  assign add_240412 = sel_240409 + 8'h01;
  assign sel_240413 = array_index_240228 == array_index_239592 ? add_240412 : sel_240409;
  assign add_240416 = sel_240413 + 8'h01;
  assign sel_240417 = array_index_240228 == array_index_239598 ? add_240416 : sel_240413;
  assign add_240420 = sel_240417 + 8'h01;
  assign sel_240421 = array_index_240228 == array_index_239604 ? add_240420 : sel_240417;
  assign add_240424 = sel_240421 + 8'h01;
  assign sel_240425 = array_index_240228 == array_index_239610 ? add_240424 : sel_240421;
  assign add_240429 = sel_240425 + 8'h01;
  assign array_index_240430 = set1_unflattened[6'h05];
  assign sel_240431 = array_index_240228 == array_index_239616 ? add_240429 : sel_240425;
  assign add_240434 = sel_240431 + 8'h01;
  assign sel_240435 = array_index_240430 == array_index_239312 ? add_240434 : sel_240431;
  assign add_240438 = sel_240435 + 8'h01;
  assign sel_240439 = array_index_240430 == array_index_239316 ? add_240438 : sel_240435;
  assign add_240442 = sel_240439 + 8'h01;
  assign sel_240443 = array_index_240430 == array_index_239324 ? add_240442 : sel_240439;
  assign add_240446 = sel_240443 + 8'h01;
  assign sel_240447 = array_index_240430 == array_index_239332 ? add_240446 : sel_240443;
  assign add_240450 = sel_240447 + 8'h01;
  assign sel_240451 = array_index_240430 == array_index_239340 ? add_240450 : sel_240447;
  assign add_240454 = sel_240451 + 8'h01;
  assign sel_240455 = array_index_240430 == array_index_239348 ? add_240454 : sel_240451;
  assign add_240458 = sel_240455 + 8'h01;
  assign sel_240459 = array_index_240430 == array_index_239356 ? add_240458 : sel_240455;
  assign add_240462 = sel_240459 + 8'h01;
  assign sel_240463 = array_index_240430 == array_index_239364 ? add_240462 : sel_240459;
  assign add_240466 = sel_240463 + 8'h01;
  assign sel_240467 = array_index_240430 == array_index_239370 ? add_240466 : sel_240463;
  assign add_240470 = sel_240467 + 8'h01;
  assign sel_240471 = array_index_240430 == array_index_239376 ? add_240470 : sel_240467;
  assign add_240474 = sel_240471 + 8'h01;
  assign sel_240475 = array_index_240430 == array_index_239382 ? add_240474 : sel_240471;
  assign add_240478 = sel_240475 + 8'h01;
  assign sel_240479 = array_index_240430 == array_index_239388 ? add_240478 : sel_240475;
  assign add_240482 = sel_240479 + 8'h01;
  assign sel_240483 = array_index_240430 == array_index_239394 ? add_240482 : sel_240479;
  assign add_240486 = sel_240483 + 8'h01;
  assign sel_240487 = array_index_240430 == array_index_239400 ? add_240486 : sel_240483;
  assign add_240490 = sel_240487 + 8'h01;
  assign sel_240491 = array_index_240430 == array_index_239406 ? add_240490 : sel_240487;
  assign add_240494 = sel_240491 + 8'h01;
  assign sel_240495 = array_index_240430 == array_index_239412 ? add_240494 : sel_240491;
  assign add_240498 = sel_240495 + 8'h01;
  assign sel_240499 = array_index_240430 == array_index_239418 ? add_240498 : sel_240495;
  assign add_240502 = sel_240499 + 8'h01;
  assign sel_240503 = array_index_240430 == array_index_239424 ? add_240502 : sel_240499;
  assign add_240506 = sel_240503 + 8'h01;
  assign sel_240507 = array_index_240430 == array_index_239430 ? add_240506 : sel_240503;
  assign add_240510 = sel_240507 + 8'h01;
  assign sel_240511 = array_index_240430 == array_index_239436 ? add_240510 : sel_240507;
  assign add_240514 = sel_240511 + 8'h01;
  assign sel_240515 = array_index_240430 == array_index_239442 ? add_240514 : sel_240511;
  assign add_240518 = sel_240515 + 8'h01;
  assign sel_240519 = array_index_240430 == array_index_239448 ? add_240518 : sel_240515;
  assign add_240522 = sel_240519 + 8'h01;
  assign sel_240523 = array_index_240430 == array_index_239454 ? add_240522 : sel_240519;
  assign add_240526 = sel_240523 + 8'h01;
  assign sel_240527 = array_index_240430 == array_index_239460 ? add_240526 : sel_240523;
  assign add_240530 = sel_240527 + 8'h01;
  assign sel_240531 = array_index_240430 == array_index_239466 ? add_240530 : sel_240527;
  assign add_240534 = sel_240531 + 8'h01;
  assign sel_240535 = array_index_240430 == array_index_239472 ? add_240534 : sel_240531;
  assign add_240538 = sel_240535 + 8'h01;
  assign sel_240539 = array_index_240430 == array_index_239478 ? add_240538 : sel_240535;
  assign add_240542 = sel_240539 + 8'h01;
  assign sel_240543 = array_index_240430 == array_index_239484 ? add_240542 : sel_240539;
  assign add_240546 = sel_240543 + 8'h01;
  assign sel_240547 = array_index_240430 == array_index_239490 ? add_240546 : sel_240543;
  assign add_240550 = sel_240547 + 8'h01;
  assign sel_240551 = array_index_240430 == array_index_239496 ? add_240550 : sel_240547;
  assign add_240554 = sel_240551 + 8'h01;
  assign sel_240555 = array_index_240430 == array_index_239502 ? add_240554 : sel_240551;
  assign add_240558 = sel_240555 + 8'h01;
  assign sel_240559 = array_index_240430 == array_index_239508 ? add_240558 : sel_240555;
  assign add_240562 = sel_240559 + 8'h01;
  assign sel_240563 = array_index_240430 == array_index_239514 ? add_240562 : sel_240559;
  assign add_240566 = sel_240563 + 8'h01;
  assign sel_240567 = array_index_240430 == array_index_239520 ? add_240566 : sel_240563;
  assign add_240570 = sel_240567 + 8'h01;
  assign sel_240571 = array_index_240430 == array_index_239526 ? add_240570 : sel_240567;
  assign add_240574 = sel_240571 + 8'h01;
  assign sel_240575 = array_index_240430 == array_index_239532 ? add_240574 : sel_240571;
  assign add_240578 = sel_240575 + 8'h01;
  assign sel_240579 = array_index_240430 == array_index_239538 ? add_240578 : sel_240575;
  assign add_240582 = sel_240579 + 8'h01;
  assign sel_240583 = array_index_240430 == array_index_239544 ? add_240582 : sel_240579;
  assign add_240586 = sel_240583 + 8'h01;
  assign sel_240587 = array_index_240430 == array_index_239550 ? add_240586 : sel_240583;
  assign add_240590 = sel_240587 + 8'h01;
  assign sel_240591 = array_index_240430 == array_index_239556 ? add_240590 : sel_240587;
  assign add_240594 = sel_240591 + 8'h01;
  assign sel_240595 = array_index_240430 == array_index_239562 ? add_240594 : sel_240591;
  assign add_240598 = sel_240595 + 8'h01;
  assign sel_240599 = array_index_240430 == array_index_239568 ? add_240598 : sel_240595;
  assign add_240602 = sel_240599 + 8'h01;
  assign sel_240603 = array_index_240430 == array_index_239574 ? add_240602 : sel_240599;
  assign add_240606 = sel_240603 + 8'h01;
  assign sel_240607 = array_index_240430 == array_index_239580 ? add_240606 : sel_240603;
  assign add_240610 = sel_240607 + 8'h01;
  assign sel_240611 = array_index_240430 == array_index_239586 ? add_240610 : sel_240607;
  assign add_240614 = sel_240611 + 8'h01;
  assign sel_240615 = array_index_240430 == array_index_239592 ? add_240614 : sel_240611;
  assign add_240618 = sel_240615 + 8'h01;
  assign sel_240619 = array_index_240430 == array_index_239598 ? add_240618 : sel_240615;
  assign add_240622 = sel_240619 + 8'h01;
  assign sel_240623 = array_index_240430 == array_index_239604 ? add_240622 : sel_240619;
  assign add_240626 = sel_240623 + 8'h01;
  assign sel_240627 = array_index_240430 == array_index_239610 ? add_240626 : sel_240623;
  assign add_240631 = sel_240627 + 8'h01;
  assign array_index_240632 = set1_unflattened[6'h06];
  assign sel_240633 = array_index_240430 == array_index_239616 ? add_240631 : sel_240627;
  assign add_240636 = sel_240633 + 8'h01;
  assign sel_240637 = array_index_240632 == array_index_239312 ? add_240636 : sel_240633;
  assign add_240640 = sel_240637 + 8'h01;
  assign sel_240641 = array_index_240632 == array_index_239316 ? add_240640 : sel_240637;
  assign add_240644 = sel_240641 + 8'h01;
  assign sel_240645 = array_index_240632 == array_index_239324 ? add_240644 : sel_240641;
  assign add_240648 = sel_240645 + 8'h01;
  assign sel_240649 = array_index_240632 == array_index_239332 ? add_240648 : sel_240645;
  assign add_240652 = sel_240649 + 8'h01;
  assign sel_240653 = array_index_240632 == array_index_239340 ? add_240652 : sel_240649;
  assign add_240656 = sel_240653 + 8'h01;
  assign sel_240657 = array_index_240632 == array_index_239348 ? add_240656 : sel_240653;
  assign add_240660 = sel_240657 + 8'h01;
  assign sel_240661 = array_index_240632 == array_index_239356 ? add_240660 : sel_240657;
  assign add_240664 = sel_240661 + 8'h01;
  assign sel_240665 = array_index_240632 == array_index_239364 ? add_240664 : sel_240661;
  assign add_240668 = sel_240665 + 8'h01;
  assign sel_240669 = array_index_240632 == array_index_239370 ? add_240668 : sel_240665;
  assign add_240672 = sel_240669 + 8'h01;
  assign sel_240673 = array_index_240632 == array_index_239376 ? add_240672 : sel_240669;
  assign add_240676 = sel_240673 + 8'h01;
  assign sel_240677 = array_index_240632 == array_index_239382 ? add_240676 : sel_240673;
  assign add_240680 = sel_240677 + 8'h01;
  assign sel_240681 = array_index_240632 == array_index_239388 ? add_240680 : sel_240677;
  assign add_240684 = sel_240681 + 8'h01;
  assign sel_240685 = array_index_240632 == array_index_239394 ? add_240684 : sel_240681;
  assign add_240688 = sel_240685 + 8'h01;
  assign sel_240689 = array_index_240632 == array_index_239400 ? add_240688 : sel_240685;
  assign add_240692 = sel_240689 + 8'h01;
  assign sel_240693 = array_index_240632 == array_index_239406 ? add_240692 : sel_240689;
  assign add_240696 = sel_240693 + 8'h01;
  assign sel_240697 = array_index_240632 == array_index_239412 ? add_240696 : sel_240693;
  assign add_240700 = sel_240697 + 8'h01;
  assign sel_240701 = array_index_240632 == array_index_239418 ? add_240700 : sel_240697;
  assign add_240704 = sel_240701 + 8'h01;
  assign sel_240705 = array_index_240632 == array_index_239424 ? add_240704 : sel_240701;
  assign add_240708 = sel_240705 + 8'h01;
  assign sel_240709 = array_index_240632 == array_index_239430 ? add_240708 : sel_240705;
  assign add_240712 = sel_240709 + 8'h01;
  assign sel_240713 = array_index_240632 == array_index_239436 ? add_240712 : sel_240709;
  assign add_240716 = sel_240713 + 8'h01;
  assign sel_240717 = array_index_240632 == array_index_239442 ? add_240716 : sel_240713;
  assign add_240720 = sel_240717 + 8'h01;
  assign sel_240721 = array_index_240632 == array_index_239448 ? add_240720 : sel_240717;
  assign add_240724 = sel_240721 + 8'h01;
  assign sel_240725 = array_index_240632 == array_index_239454 ? add_240724 : sel_240721;
  assign add_240728 = sel_240725 + 8'h01;
  assign sel_240729 = array_index_240632 == array_index_239460 ? add_240728 : sel_240725;
  assign add_240732 = sel_240729 + 8'h01;
  assign sel_240733 = array_index_240632 == array_index_239466 ? add_240732 : sel_240729;
  assign add_240736 = sel_240733 + 8'h01;
  assign sel_240737 = array_index_240632 == array_index_239472 ? add_240736 : sel_240733;
  assign add_240740 = sel_240737 + 8'h01;
  assign sel_240741 = array_index_240632 == array_index_239478 ? add_240740 : sel_240737;
  assign add_240744 = sel_240741 + 8'h01;
  assign sel_240745 = array_index_240632 == array_index_239484 ? add_240744 : sel_240741;
  assign add_240748 = sel_240745 + 8'h01;
  assign sel_240749 = array_index_240632 == array_index_239490 ? add_240748 : sel_240745;
  assign add_240752 = sel_240749 + 8'h01;
  assign sel_240753 = array_index_240632 == array_index_239496 ? add_240752 : sel_240749;
  assign add_240756 = sel_240753 + 8'h01;
  assign sel_240757 = array_index_240632 == array_index_239502 ? add_240756 : sel_240753;
  assign add_240760 = sel_240757 + 8'h01;
  assign sel_240761 = array_index_240632 == array_index_239508 ? add_240760 : sel_240757;
  assign add_240764 = sel_240761 + 8'h01;
  assign sel_240765 = array_index_240632 == array_index_239514 ? add_240764 : sel_240761;
  assign add_240768 = sel_240765 + 8'h01;
  assign sel_240769 = array_index_240632 == array_index_239520 ? add_240768 : sel_240765;
  assign add_240772 = sel_240769 + 8'h01;
  assign sel_240773 = array_index_240632 == array_index_239526 ? add_240772 : sel_240769;
  assign add_240776 = sel_240773 + 8'h01;
  assign sel_240777 = array_index_240632 == array_index_239532 ? add_240776 : sel_240773;
  assign add_240780 = sel_240777 + 8'h01;
  assign sel_240781 = array_index_240632 == array_index_239538 ? add_240780 : sel_240777;
  assign add_240784 = sel_240781 + 8'h01;
  assign sel_240785 = array_index_240632 == array_index_239544 ? add_240784 : sel_240781;
  assign add_240788 = sel_240785 + 8'h01;
  assign sel_240789 = array_index_240632 == array_index_239550 ? add_240788 : sel_240785;
  assign add_240792 = sel_240789 + 8'h01;
  assign sel_240793 = array_index_240632 == array_index_239556 ? add_240792 : sel_240789;
  assign add_240796 = sel_240793 + 8'h01;
  assign sel_240797 = array_index_240632 == array_index_239562 ? add_240796 : sel_240793;
  assign add_240800 = sel_240797 + 8'h01;
  assign sel_240801 = array_index_240632 == array_index_239568 ? add_240800 : sel_240797;
  assign add_240804 = sel_240801 + 8'h01;
  assign sel_240805 = array_index_240632 == array_index_239574 ? add_240804 : sel_240801;
  assign add_240808 = sel_240805 + 8'h01;
  assign sel_240809 = array_index_240632 == array_index_239580 ? add_240808 : sel_240805;
  assign add_240812 = sel_240809 + 8'h01;
  assign sel_240813 = array_index_240632 == array_index_239586 ? add_240812 : sel_240809;
  assign add_240816 = sel_240813 + 8'h01;
  assign sel_240817 = array_index_240632 == array_index_239592 ? add_240816 : sel_240813;
  assign add_240820 = sel_240817 + 8'h01;
  assign sel_240821 = array_index_240632 == array_index_239598 ? add_240820 : sel_240817;
  assign add_240824 = sel_240821 + 8'h01;
  assign sel_240825 = array_index_240632 == array_index_239604 ? add_240824 : sel_240821;
  assign add_240828 = sel_240825 + 8'h01;
  assign sel_240829 = array_index_240632 == array_index_239610 ? add_240828 : sel_240825;
  assign add_240833 = sel_240829 + 8'h01;
  assign array_index_240834 = set1_unflattened[6'h07];
  assign sel_240835 = array_index_240632 == array_index_239616 ? add_240833 : sel_240829;
  assign add_240838 = sel_240835 + 8'h01;
  assign sel_240839 = array_index_240834 == array_index_239312 ? add_240838 : sel_240835;
  assign add_240842 = sel_240839 + 8'h01;
  assign sel_240843 = array_index_240834 == array_index_239316 ? add_240842 : sel_240839;
  assign add_240846 = sel_240843 + 8'h01;
  assign sel_240847 = array_index_240834 == array_index_239324 ? add_240846 : sel_240843;
  assign add_240850 = sel_240847 + 8'h01;
  assign sel_240851 = array_index_240834 == array_index_239332 ? add_240850 : sel_240847;
  assign add_240854 = sel_240851 + 8'h01;
  assign sel_240855 = array_index_240834 == array_index_239340 ? add_240854 : sel_240851;
  assign add_240858 = sel_240855 + 8'h01;
  assign sel_240859 = array_index_240834 == array_index_239348 ? add_240858 : sel_240855;
  assign add_240862 = sel_240859 + 8'h01;
  assign sel_240863 = array_index_240834 == array_index_239356 ? add_240862 : sel_240859;
  assign add_240866 = sel_240863 + 8'h01;
  assign sel_240867 = array_index_240834 == array_index_239364 ? add_240866 : sel_240863;
  assign add_240870 = sel_240867 + 8'h01;
  assign sel_240871 = array_index_240834 == array_index_239370 ? add_240870 : sel_240867;
  assign add_240874 = sel_240871 + 8'h01;
  assign sel_240875 = array_index_240834 == array_index_239376 ? add_240874 : sel_240871;
  assign add_240878 = sel_240875 + 8'h01;
  assign sel_240879 = array_index_240834 == array_index_239382 ? add_240878 : sel_240875;
  assign add_240882 = sel_240879 + 8'h01;
  assign sel_240883 = array_index_240834 == array_index_239388 ? add_240882 : sel_240879;
  assign add_240886 = sel_240883 + 8'h01;
  assign sel_240887 = array_index_240834 == array_index_239394 ? add_240886 : sel_240883;
  assign add_240890 = sel_240887 + 8'h01;
  assign sel_240891 = array_index_240834 == array_index_239400 ? add_240890 : sel_240887;
  assign add_240894 = sel_240891 + 8'h01;
  assign sel_240895 = array_index_240834 == array_index_239406 ? add_240894 : sel_240891;
  assign add_240898 = sel_240895 + 8'h01;
  assign sel_240899 = array_index_240834 == array_index_239412 ? add_240898 : sel_240895;
  assign add_240902 = sel_240899 + 8'h01;
  assign sel_240903 = array_index_240834 == array_index_239418 ? add_240902 : sel_240899;
  assign add_240906 = sel_240903 + 8'h01;
  assign sel_240907 = array_index_240834 == array_index_239424 ? add_240906 : sel_240903;
  assign add_240910 = sel_240907 + 8'h01;
  assign sel_240911 = array_index_240834 == array_index_239430 ? add_240910 : sel_240907;
  assign add_240914 = sel_240911 + 8'h01;
  assign sel_240915 = array_index_240834 == array_index_239436 ? add_240914 : sel_240911;
  assign add_240918 = sel_240915 + 8'h01;
  assign sel_240919 = array_index_240834 == array_index_239442 ? add_240918 : sel_240915;
  assign add_240922 = sel_240919 + 8'h01;
  assign sel_240923 = array_index_240834 == array_index_239448 ? add_240922 : sel_240919;
  assign add_240926 = sel_240923 + 8'h01;
  assign sel_240927 = array_index_240834 == array_index_239454 ? add_240926 : sel_240923;
  assign add_240930 = sel_240927 + 8'h01;
  assign sel_240931 = array_index_240834 == array_index_239460 ? add_240930 : sel_240927;
  assign add_240934 = sel_240931 + 8'h01;
  assign sel_240935 = array_index_240834 == array_index_239466 ? add_240934 : sel_240931;
  assign add_240938 = sel_240935 + 8'h01;
  assign sel_240939 = array_index_240834 == array_index_239472 ? add_240938 : sel_240935;
  assign add_240942 = sel_240939 + 8'h01;
  assign sel_240943 = array_index_240834 == array_index_239478 ? add_240942 : sel_240939;
  assign add_240946 = sel_240943 + 8'h01;
  assign sel_240947 = array_index_240834 == array_index_239484 ? add_240946 : sel_240943;
  assign add_240950 = sel_240947 + 8'h01;
  assign sel_240951 = array_index_240834 == array_index_239490 ? add_240950 : sel_240947;
  assign add_240954 = sel_240951 + 8'h01;
  assign sel_240955 = array_index_240834 == array_index_239496 ? add_240954 : sel_240951;
  assign add_240958 = sel_240955 + 8'h01;
  assign sel_240959 = array_index_240834 == array_index_239502 ? add_240958 : sel_240955;
  assign add_240962 = sel_240959 + 8'h01;
  assign sel_240963 = array_index_240834 == array_index_239508 ? add_240962 : sel_240959;
  assign add_240966 = sel_240963 + 8'h01;
  assign sel_240967 = array_index_240834 == array_index_239514 ? add_240966 : sel_240963;
  assign add_240970 = sel_240967 + 8'h01;
  assign sel_240971 = array_index_240834 == array_index_239520 ? add_240970 : sel_240967;
  assign add_240974 = sel_240971 + 8'h01;
  assign sel_240975 = array_index_240834 == array_index_239526 ? add_240974 : sel_240971;
  assign add_240978 = sel_240975 + 8'h01;
  assign sel_240979 = array_index_240834 == array_index_239532 ? add_240978 : sel_240975;
  assign add_240982 = sel_240979 + 8'h01;
  assign sel_240983 = array_index_240834 == array_index_239538 ? add_240982 : sel_240979;
  assign add_240986 = sel_240983 + 8'h01;
  assign sel_240987 = array_index_240834 == array_index_239544 ? add_240986 : sel_240983;
  assign add_240990 = sel_240987 + 8'h01;
  assign sel_240991 = array_index_240834 == array_index_239550 ? add_240990 : sel_240987;
  assign add_240994 = sel_240991 + 8'h01;
  assign sel_240995 = array_index_240834 == array_index_239556 ? add_240994 : sel_240991;
  assign add_240998 = sel_240995 + 8'h01;
  assign sel_240999 = array_index_240834 == array_index_239562 ? add_240998 : sel_240995;
  assign add_241002 = sel_240999 + 8'h01;
  assign sel_241003 = array_index_240834 == array_index_239568 ? add_241002 : sel_240999;
  assign add_241006 = sel_241003 + 8'h01;
  assign sel_241007 = array_index_240834 == array_index_239574 ? add_241006 : sel_241003;
  assign add_241010 = sel_241007 + 8'h01;
  assign sel_241011 = array_index_240834 == array_index_239580 ? add_241010 : sel_241007;
  assign add_241014 = sel_241011 + 8'h01;
  assign sel_241015 = array_index_240834 == array_index_239586 ? add_241014 : sel_241011;
  assign add_241018 = sel_241015 + 8'h01;
  assign sel_241019 = array_index_240834 == array_index_239592 ? add_241018 : sel_241015;
  assign add_241022 = sel_241019 + 8'h01;
  assign sel_241023 = array_index_240834 == array_index_239598 ? add_241022 : sel_241019;
  assign add_241026 = sel_241023 + 8'h01;
  assign sel_241027 = array_index_240834 == array_index_239604 ? add_241026 : sel_241023;
  assign add_241030 = sel_241027 + 8'h01;
  assign sel_241031 = array_index_240834 == array_index_239610 ? add_241030 : sel_241027;
  assign add_241035 = sel_241031 + 8'h01;
  assign array_index_241036 = set1_unflattened[6'h08];
  assign sel_241037 = array_index_240834 == array_index_239616 ? add_241035 : sel_241031;
  assign add_241040 = sel_241037 + 8'h01;
  assign sel_241041 = array_index_241036 == array_index_239312 ? add_241040 : sel_241037;
  assign add_241044 = sel_241041 + 8'h01;
  assign sel_241045 = array_index_241036 == array_index_239316 ? add_241044 : sel_241041;
  assign add_241048 = sel_241045 + 8'h01;
  assign sel_241049 = array_index_241036 == array_index_239324 ? add_241048 : sel_241045;
  assign add_241052 = sel_241049 + 8'h01;
  assign sel_241053 = array_index_241036 == array_index_239332 ? add_241052 : sel_241049;
  assign add_241056 = sel_241053 + 8'h01;
  assign sel_241057 = array_index_241036 == array_index_239340 ? add_241056 : sel_241053;
  assign add_241060 = sel_241057 + 8'h01;
  assign sel_241061 = array_index_241036 == array_index_239348 ? add_241060 : sel_241057;
  assign add_241064 = sel_241061 + 8'h01;
  assign sel_241065 = array_index_241036 == array_index_239356 ? add_241064 : sel_241061;
  assign add_241068 = sel_241065 + 8'h01;
  assign sel_241069 = array_index_241036 == array_index_239364 ? add_241068 : sel_241065;
  assign add_241072 = sel_241069 + 8'h01;
  assign sel_241073 = array_index_241036 == array_index_239370 ? add_241072 : sel_241069;
  assign add_241076 = sel_241073 + 8'h01;
  assign sel_241077 = array_index_241036 == array_index_239376 ? add_241076 : sel_241073;
  assign add_241080 = sel_241077 + 8'h01;
  assign sel_241081 = array_index_241036 == array_index_239382 ? add_241080 : sel_241077;
  assign add_241084 = sel_241081 + 8'h01;
  assign sel_241085 = array_index_241036 == array_index_239388 ? add_241084 : sel_241081;
  assign add_241088 = sel_241085 + 8'h01;
  assign sel_241089 = array_index_241036 == array_index_239394 ? add_241088 : sel_241085;
  assign add_241092 = sel_241089 + 8'h01;
  assign sel_241093 = array_index_241036 == array_index_239400 ? add_241092 : sel_241089;
  assign add_241096 = sel_241093 + 8'h01;
  assign sel_241097 = array_index_241036 == array_index_239406 ? add_241096 : sel_241093;
  assign add_241100 = sel_241097 + 8'h01;
  assign sel_241101 = array_index_241036 == array_index_239412 ? add_241100 : sel_241097;
  assign add_241104 = sel_241101 + 8'h01;
  assign sel_241105 = array_index_241036 == array_index_239418 ? add_241104 : sel_241101;
  assign add_241108 = sel_241105 + 8'h01;
  assign sel_241109 = array_index_241036 == array_index_239424 ? add_241108 : sel_241105;
  assign add_241112 = sel_241109 + 8'h01;
  assign sel_241113 = array_index_241036 == array_index_239430 ? add_241112 : sel_241109;
  assign add_241116 = sel_241113 + 8'h01;
  assign sel_241117 = array_index_241036 == array_index_239436 ? add_241116 : sel_241113;
  assign add_241120 = sel_241117 + 8'h01;
  assign sel_241121 = array_index_241036 == array_index_239442 ? add_241120 : sel_241117;
  assign add_241124 = sel_241121 + 8'h01;
  assign sel_241125 = array_index_241036 == array_index_239448 ? add_241124 : sel_241121;
  assign add_241128 = sel_241125 + 8'h01;
  assign sel_241129 = array_index_241036 == array_index_239454 ? add_241128 : sel_241125;
  assign add_241132 = sel_241129 + 8'h01;
  assign sel_241133 = array_index_241036 == array_index_239460 ? add_241132 : sel_241129;
  assign add_241136 = sel_241133 + 8'h01;
  assign sel_241137 = array_index_241036 == array_index_239466 ? add_241136 : sel_241133;
  assign add_241140 = sel_241137 + 8'h01;
  assign sel_241141 = array_index_241036 == array_index_239472 ? add_241140 : sel_241137;
  assign add_241144 = sel_241141 + 8'h01;
  assign sel_241145 = array_index_241036 == array_index_239478 ? add_241144 : sel_241141;
  assign add_241148 = sel_241145 + 8'h01;
  assign sel_241149 = array_index_241036 == array_index_239484 ? add_241148 : sel_241145;
  assign add_241152 = sel_241149 + 8'h01;
  assign sel_241153 = array_index_241036 == array_index_239490 ? add_241152 : sel_241149;
  assign add_241156 = sel_241153 + 8'h01;
  assign sel_241157 = array_index_241036 == array_index_239496 ? add_241156 : sel_241153;
  assign add_241160 = sel_241157 + 8'h01;
  assign sel_241161 = array_index_241036 == array_index_239502 ? add_241160 : sel_241157;
  assign add_241164 = sel_241161 + 8'h01;
  assign sel_241165 = array_index_241036 == array_index_239508 ? add_241164 : sel_241161;
  assign add_241168 = sel_241165 + 8'h01;
  assign sel_241169 = array_index_241036 == array_index_239514 ? add_241168 : sel_241165;
  assign add_241172 = sel_241169 + 8'h01;
  assign sel_241173 = array_index_241036 == array_index_239520 ? add_241172 : sel_241169;
  assign add_241176 = sel_241173 + 8'h01;
  assign sel_241177 = array_index_241036 == array_index_239526 ? add_241176 : sel_241173;
  assign add_241180 = sel_241177 + 8'h01;
  assign sel_241181 = array_index_241036 == array_index_239532 ? add_241180 : sel_241177;
  assign add_241184 = sel_241181 + 8'h01;
  assign sel_241185 = array_index_241036 == array_index_239538 ? add_241184 : sel_241181;
  assign add_241188 = sel_241185 + 8'h01;
  assign sel_241189 = array_index_241036 == array_index_239544 ? add_241188 : sel_241185;
  assign add_241192 = sel_241189 + 8'h01;
  assign sel_241193 = array_index_241036 == array_index_239550 ? add_241192 : sel_241189;
  assign add_241196 = sel_241193 + 8'h01;
  assign sel_241197 = array_index_241036 == array_index_239556 ? add_241196 : sel_241193;
  assign add_241200 = sel_241197 + 8'h01;
  assign sel_241201 = array_index_241036 == array_index_239562 ? add_241200 : sel_241197;
  assign add_241204 = sel_241201 + 8'h01;
  assign sel_241205 = array_index_241036 == array_index_239568 ? add_241204 : sel_241201;
  assign add_241208 = sel_241205 + 8'h01;
  assign sel_241209 = array_index_241036 == array_index_239574 ? add_241208 : sel_241205;
  assign add_241212 = sel_241209 + 8'h01;
  assign sel_241213 = array_index_241036 == array_index_239580 ? add_241212 : sel_241209;
  assign add_241216 = sel_241213 + 8'h01;
  assign sel_241217 = array_index_241036 == array_index_239586 ? add_241216 : sel_241213;
  assign add_241220 = sel_241217 + 8'h01;
  assign sel_241221 = array_index_241036 == array_index_239592 ? add_241220 : sel_241217;
  assign add_241224 = sel_241221 + 8'h01;
  assign sel_241225 = array_index_241036 == array_index_239598 ? add_241224 : sel_241221;
  assign add_241228 = sel_241225 + 8'h01;
  assign sel_241229 = array_index_241036 == array_index_239604 ? add_241228 : sel_241225;
  assign add_241232 = sel_241229 + 8'h01;
  assign sel_241233 = array_index_241036 == array_index_239610 ? add_241232 : sel_241229;
  assign add_241237 = sel_241233 + 8'h01;
  assign array_index_241238 = set1_unflattened[6'h09];
  assign sel_241239 = array_index_241036 == array_index_239616 ? add_241237 : sel_241233;
  assign add_241242 = sel_241239 + 8'h01;
  assign sel_241243 = array_index_241238 == array_index_239312 ? add_241242 : sel_241239;
  assign add_241246 = sel_241243 + 8'h01;
  assign sel_241247 = array_index_241238 == array_index_239316 ? add_241246 : sel_241243;
  assign add_241250 = sel_241247 + 8'h01;
  assign sel_241251 = array_index_241238 == array_index_239324 ? add_241250 : sel_241247;
  assign add_241254 = sel_241251 + 8'h01;
  assign sel_241255 = array_index_241238 == array_index_239332 ? add_241254 : sel_241251;
  assign add_241258 = sel_241255 + 8'h01;
  assign sel_241259 = array_index_241238 == array_index_239340 ? add_241258 : sel_241255;
  assign add_241262 = sel_241259 + 8'h01;
  assign sel_241263 = array_index_241238 == array_index_239348 ? add_241262 : sel_241259;
  assign add_241266 = sel_241263 + 8'h01;
  assign sel_241267 = array_index_241238 == array_index_239356 ? add_241266 : sel_241263;
  assign add_241270 = sel_241267 + 8'h01;
  assign sel_241271 = array_index_241238 == array_index_239364 ? add_241270 : sel_241267;
  assign add_241274 = sel_241271 + 8'h01;
  assign sel_241275 = array_index_241238 == array_index_239370 ? add_241274 : sel_241271;
  assign add_241278 = sel_241275 + 8'h01;
  assign sel_241279 = array_index_241238 == array_index_239376 ? add_241278 : sel_241275;
  assign add_241282 = sel_241279 + 8'h01;
  assign sel_241283 = array_index_241238 == array_index_239382 ? add_241282 : sel_241279;
  assign add_241286 = sel_241283 + 8'h01;
  assign sel_241287 = array_index_241238 == array_index_239388 ? add_241286 : sel_241283;
  assign add_241290 = sel_241287 + 8'h01;
  assign sel_241291 = array_index_241238 == array_index_239394 ? add_241290 : sel_241287;
  assign add_241294 = sel_241291 + 8'h01;
  assign sel_241295 = array_index_241238 == array_index_239400 ? add_241294 : sel_241291;
  assign add_241298 = sel_241295 + 8'h01;
  assign sel_241299 = array_index_241238 == array_index_239406 ? add_241298 : sel_241295;
  assign add_241302 = sel_241299 + 8'h01;
  assign sel_241303 = array_index_241238 == array_index_239412 ? add_241302 : sel_241299;
  assign add_241306 = sel_241303 + 8'h01;
  assign sel_241307 = array_index_241238 == array_index_239418 ? add_241306 : sel_241303;
  assign add_241310 = sel_241307 + 8'h01;
  assign sel_241311 = array_index_241238 == array_index_239424 ? add_241310 : sel_241307;
  assign add_241314 = sel_241311 + 8'h01;
  assign sel_241315 = array_index_241238 == array_index_239430 ? add_241314 : sel_241311;
  assign add_241318 = sel_241315 + 8'h01;
  assign sel_241319 = array_index_241238 == array_index_239436 ? add_241318 : sel_241315;
  assign add_241322 = sel_241319 + 8'h01;
  assign sel_241323 = array_index_241238 == array_index_239442 ? add_241322 : sel_241319;
  assign add_241326 = sel_241323 + 8'h01;
  assign sel_241327 = array_index_241238 == array_index_239448 ? add_241326 : sel_241323;
  assign add_241330 = sel_241327 + 8'h01;
  assign sel_241331 = array_index_241238 == array_index_239454 ? add_241330 : sel_241327;
  assign add_241334 = sel_241331 + 8'h01;
  assign sel_241335 = array_index_241238 == array_index_239460 ? add_241334 : sel_241331;
  assign add_241338 = sel_241335 + 8'h01;
  assign sel_241339 = array_index_241238 == array_index_239466 ? add_241338 : sel_241335;
  assign add_241342 = sel_241339 + 8'h01;
  assign sel_241343 = array_index_241238 == array_index_239472 ? add_241342 : sel_241339;
  assign add_241346 = sel_241343 + 8'h01;
  assign sel_241347 = array_index_241238 == array_index_239478 ? add_241346 : sel_241343;
  assign add_241350 = sel_241347 + 8'h01;
  assign sel_241351 = array_index_241238 == array_index_239484 ? add_241350 : sel_241347;
  assign add_241354 = sel_241351 + 8'h01;
  assign sel_241355 = array_index_241238 == array_index_239490 ? add_241354 : sel_241351;
  assign add_241358 = sel_241355 + 8'h01;
  assign sel_241359 = array_index_241238 == array_index_239496 ? add_241358 : sel_241355;
  assign add_241362 = sel_241359 + 8'h01;
  assign sel_241363 = array_index_241238 == array_index_239502 ? add_241362 : sel_241359;
  assign add_241366 = sel_241363 + 8'h01;
  assign sel_241367 = array_index_241238 == array_index_239508 ? add_241366 : sel_241363;
  assign add_241370 = sel_241367 + 8'h01;
  assign sel_241371 = array_index_241238 == array_index_239514 ? add_241370 : sel_241367;
  assign add_241374 = sel_241371 + 8'h01;
  assign sel_241375 = array_index_241238 == array_index_239520 ? add_241374 : sel_241371;
  assign add_241378 = sel_241375 + 8'h01;
  assign sel_241379 = array_index_241238 == array_index_239526 ? add_241378 : sel_241375;
  assign add_241382 = sel_241379 + 8'h01;
  assign sel_241383 = array_index_241238 == array_index_239532 ? add_241382 : sel_241379;
  assign add_241386 = sel_241383 + 8'h01;
  assign sel_241387 = array_index_241238 == array_index_239538 ? add_241386 : sel_241383;
  assign add_241390 = sel_241387 + 8'h01;
  assign sel_241391 = array_index_241238 == array_index_239544 ? add_241390 : sel_241387;
  assign add_241394 = sel_241391 + 8'h01;
  assign sel_241395 = array_index_241238 == array_index_239550 ? add_241394 : sel_241391;
  assign add_241398 = sel_241395 + 8'h01;
  assign sel_241399 = array_index_241238 == array_index_239556 ? add_241398 : sel_241395;
  assign add_241402 = sel_241399 + 8'h01;
  assign sel_241403 = array_index_241238 == array_index_239562 ? add_241402 : sel_241399;
  assign add_241406 = sel_241403 + 8'h01;
  assign sel_241407 = array_index_241238 == array_index_239568 ? add_241406 : sel_241403;
  assign add_241410 = sel_241407 + 8'h01;
  assign sel_241411 = array_index_241238 == array_index_239574 ? add_241410 : sel_241407;
  assign add_241414 = sel_241411 + 8'h01;
  assign sel_241415 = array_index_241238 == array_index_239580 ? add_241414 : sel_241411;
  assign add_241418 = sel_241415 + 8'h01;
  assign sel_241419 = array_index_241238 == array_index_239586 ? add_241418 : sel_241415;
  assign add_241422 = sel_241419 + 8'h01;
  assign sel_241423 = array_index_241238 == array_index_239592 ? add_241422 : sel_241419;
  assign add_241426 = sel_241423 + 8'h01;
  assign sel_241427 = array_index_241238 == array_index_239598 ? add_241426 : sel_241423;
  assign add_241430 = sel_241427 + 8'h01;
  assign sel_241431 = array_index_241238 == array_index_239604 ? add_241430 : sel_241427;
  assign add_241434 = sel_241431 + 8'h01;
  assign sel_241435 = array_index_241238 == array_index_239610 ? add_241434 : sel_241431;
  assign add_241439 = sel_241435 + 8'h01;
  assign array_index_241440 = set1_unflattened[6'h0a];
  assign sel_241441 = array_index_241238 == array_index_239616 ? add_241439 : sel_241435;
  assign add_241444 = sel_241441 + 8'h01;
  assign sel_241445 = array_index_241440 == array_index_239312 ? add_241444 : sel_241441;
  assign add_241448 = sel_241445 + 8'h01;
  assign sel_241449 = array_index_241440 == array_index_239316 ? add_241448 : sel_241445;
  assign add_241452 = sel_241449 + 8'h01;
  assign sel_241453 = array_index_241440 == array_index_239324 ? add_241452 : sel_241449;
  assign add_241456 = sel_241453 + 8'h01;
  assign sel_241457 = array_index_241440 == array_index_239332 ? add_241456 : sel_241453;
  assign add_241460 = sel_241457 + 8'h01;
  assign sel_241461 = array_index_241440 == array_index_239340 ? add_241460 : sel_241457;
  assign add_241464 = sel_241461 + 8'h01;
  assign sel_241465 = array_index_241440 == array_index_239348 ? add_241464 : sel_241461;
  assign add_241468 = sel_241465 + 8'h01;
  assign sel_241469 = array_index_241440 == array_index_239356 ? add_241468 : sel_241465;
  assign add_241472 = sel_241469 + 8'h01;
  assign sel_241473 = array_index_241440 == array_index_239364 ? add_241472 : sel_241469;
  assign add_241476 = sel_241473 + 8'h01;
  assign sel_241477 = array_index_241440 == array_index_239370 ? add_241476 : sel_241473;
  assign add_241480 = sel_241477 + 8'h01;
  assign sel_241481 = array_index_241440 == array_index_239376 ? add_241480 : sel_241477;
  assign add_241484 = sel_241481 + 8'h01;
  assign sel_241485 = array_index_241440 == array_index_239382 ? add_241484 : sel_241481;
  assign add_241488 = sel_241485 + 8'h01;
  assign sel_241489 = array_index_241440 == array_index_239388 ? add_241488 : sel_241485;
  assign add_241492 = sel_241489 + 8'h01;
  assign sel_241493 = array_index_241440 == array_index_239394 ? add_241492 : sel_241489;
  assign add_241496 = sel_241493 + 8'h01;
  assign sel_241497 = array_index_241440 == array_index_239400 ? add_241496 : sel_241493;
  assign add_241500 = sel_241497 + 8'h01;
  assign sel_241501 = array_index_241440 == array_index_239406 ? add_241500 : sel_241497;
  assign add_241504 = sel_241501 + 8'h01;
  assign sel_241505 = array_index_241440 == array_index_239412 ? add_241504 : sel_241501;
  assign add_241508 = sel_241505 + 8'h01;
  assign sel_241509 = array_index_241440 == array_index_239418 ? add_241508 : sel_241505;
  assign add_241512 = sel_241509 + 8'h01;
  assign sel_241513 = array_index_241440 == array_index_239424 ? add_241512 : sel_241509;
  assign add_241516 = sel_241513 + 8'h01;
  assign sel_241517 = array_index_241440 == array_index_239430 ? add_241516 : sel_241513;
  assign add_241520 = sel_241517 + 8'h01;
  assign sel_241521 = array_index_241440 == array_index_239436 ? add_241520 : sel_241517;
  assign add_241524 = sel_241521 + 8'h01;
  assign sel_241525 = array_index_241440 == array_index_239442 ? add_241524 : sel_241521;
  assign add_241528 = sel_241525 + 8'h01;
  assign sel_241529 = array_index_241440 == array_index_239448 ? add_241528 : sel_241525;
  assign add_241532 = sel_241529 + 8'h01;
  assign sel_241533 = array_index_241440 == array_index_239454 ? add_241532 : sel_241529;
  assign add_241536 = sel_241533 + 8'h01;
  assign sel_241537 = array_index_241440 == array_index_239460 ? add_241536 : sel_241533;
  assign add_241540 = sel_241537 + 8'h01;
  assign sel_241541 = array_index_241440 == array_index_239466 ? add_241540 : sel_241537;
  assign add_241544 = sel_241541 + 8'h01;
  assign sel_241545 = array_index_241440 == array_index_239472 ? add_241544 : sel_241541;
  assign add_241548 = sel_241545 + 8'h01;
  assign sel_241549 = array_index_241440 == array_index_239478 ? add_241548 : sel_241545;
  assign add_241552 = sel_241549 + 8'h01;
  assign sel_241553 = array_index_241440 == array_index_239484 ? add_241552 : sel_241549;
  assign add_241556 = sel_241553 + 8'h01;
  assign sel_241557 = array_index_241440 == array_index_239490 ? add_241556 : sel_241553;
  assign add_241560 = sel_241557 + 8'h01;
  assign sel_241561 = array_index_241440 == array_index_239496 ? add_241560 : sel_241557;
  assign add_241564 = sel_241561 + 8'h01;
  assign sel_241565 = array_index_241440 == array_index_239502 ? add_241564 : sel_241561;
  assign add_241568 = sel_241565 + 8'h01;
  assign sel_241569 = array_index_241440 == array_index_239508 ? add_241568 : sel_241565;
  assign add_241572 = sel_241569 + 8'h01;
  assign sel_241573 = array_index_241440 == array_index_239514 ? add_241572 : sel_241569;
  assign add_241576 = sel_241573 + 8'h01;
  assign sel_241577 = array_index_241440 == array_index_239520 ? add_241576 : sel_241573;
  assign add_241580 = sel_241577 + 8'h01;
  assign sel_241581 = array_index_241440 == array_index_239526 ? add_241580 : sel_241577;
  assign add_241584 = sel_241581 + 8'h01;
  assign sel_241585 = array_index_241440 == array_index_239532 ? add_241584 : sel_241581;
  assign add_241588 = sel_241585 + 8'h01;
  assign sel_241589 = array_index_241440 == array_index_239538 ? add_241588 : sel_241585;
  assign add_241592 = sel_241589 + 8'h01;
  assign sel_241593 = array_index_241440 == array_index_239544 ? add_241592 : sel_241589;
  assign add_241596 = sel_241593 + 8'h01;
  assign sel_241597 = array_index_241440 == array_index_239550 ? add_241596 : sel_241593;
  assign add_241600 = sel_241597 + 8'h01;
  assign sel_241601 = array_index_241440 == array_index_239556 ? add_241600 : sel_241597;
  assign add_241604 = sel_241601 + 8'h01;
  assign sel_241605 = array_index_241440 == array_index_239562 ? add_241604 : sel_241601;
  assign add_241608 = sel_241605 + 8'h01;
  assign sel_241609 = array_index_241440 == array_index_239568 ? add_241608 : sel_241605;
  assign add_241612 = sel_241609 + 8'h01;
  assign sel_241613 = array_index_241440 == array_index_239574 ? add_241612 : sel_241609;
  assign add_241616 = sel_241613 + 8'h01;
  assign sel_241617 = array_index_241440 == array_index_239580 ? add_241616 : sel_241613;
  assign add_241620 = sel_241617 + 8'h01;
  assign sel_241621 = array_index_241440 == array_index_239586 ? add_241620 : sel_241617;
  assign add_241624 = sel_241621 + 8'h01;
  assign sel_241625 = array_index_241440 == array_index_239592 ? add_241624 : sel_241621;
  assign add_241628 = sel_241625 + 8'h01;
  assign sel_241629 = array_index_241440 == array_index_239598 ? add_241628 : sel_241625;
  assign add_241632 = sel_241629 + 8'h01;
  assign sel_241633 = array_index_241440 == array_index_239604 ? add_241632 : sel_241629;
  assign add_241636 = sel_241633 + 8'h01;
  assign sel_241637 = array_index_241440 == array_index_239610 ? add_241636 : sel_241633;
  assign add_241641 = sel_241637 + 8'h01;
  assign array_index_241642 = set1_unflattened[6'h0b];
  assign sel_241643 = array_index_241440 == array_index_239616 ? add_241641 : sel_241637;
  assign add_241646 = sel_241643 + 8'h01;
  assign sel_241647 = array_index_241642 == array_index_239312 ? add_241646 : sel_241643;
  assign add_241650 = sel_241647 + 8'h01;
  assign sel_241651 = array_index_241642 == array_index_239316 ? add_241650 : sel_241647;
  assign add_241654 = sel_241651 + 8'h01;
  assign sel_241655 = array_index_241642 == array_index_239324 ? add_241654 : sel_241651;
  assign add_241658 = sel_241655 + 8'h01;
  assign sel_241659 = array_index_241642 == array_index_239332 ? add_241658 : sel_241655;
  assign add_241662 = sel_241659 + 8'h01;
  assign sel_241663 = array_index_241642 == array_index_239340 ? add_241662 : sel_241659;
  assign add_241666 = sel_241663 + 8'h01;
  assign sel_241667 = array_index_241642 == array_index_239348 ? add_241666 : sel_241663;
  assign add_241670 = sel_241667 + 8'h01;
  assign sel_241671 = array_index_241642 == array_index_239356 ? add_241670 : sel_241667;
  assign add_241674 = sel_241671 + 8'h01;
  assign sel_241675 = array_index_241642 == array_index_239364 ? add_241674 : sel_241671;
  assign add_241678 = sel_241675 + 8'h01;
  assign sel_241679 = array_index_241642 == array_index_239370 ? add_241678 : sel_241675;
  assign add_241682 = sel_241679 + 8'h01;
  assign sel_241683 = array_index_241642 == array_index_239376 ? add_241682 : sel_241679;
  assign add_241686 = sel_241683 + 8'h01;
  assign sel_241687 = array_index_241642 == array_index_239382 ? add_241686 : sel_241683;
  assign add_241690 = sel_241687 + 8'h01;
  assign sel_241691 = array_index_241642 == array_index_239388 ? add_241690 : sel_241687;
  assign add_241694 = sel_241691 + 8'h01;
  assign sel_241695 = array_index_241642 == array_index_239394 ? add_241694 : sel_241691;
  assign add_241698 = sel_241695 + 8'h01;
  assign sel_241699 = array_index_241642 == array_index_239400 ? add_241698 : sel_241695;
  assign add_241702 = sel_241699 + 8'h01;
  assign sel_241703 = array_index_241642 == array_index_239406 ? add_241702 : sel_241699;
  assign add_241706 = sel_241703 + 8'h01;
  assign sel_241707 = array_index_241642 == array_index_239412 ? add_241706 : sel_241703;
  assign add_241710 = sel_241707 + 8'h01;
  assign sel_241711 = array_index_241642 == array_index_239418 ? add_241710 : sel_241707;
  assign add_241714 = sel_241711 + 8'h01;
  assign sel_241715 = array_index_241642 == array_index_239424 ? add_241714 : sel_241711;
  assign add_241718 = sel_241715 + 8'h01;
  assign sel_241719 = array_index_241642 == array_index_239430 ? add_241718 : sel_241715;
  assign add_241722 = sel_241719 + 8'h01;
  assign sel_241723 = array_index_241642 == array_index_239436 ? add_241722 : sel_241719;
  assign add_241726 = sel_241723 + 8'h01;
  assign sel_241727 = array_index_241642 == array_index_239442 ? add_241726 : sel_241723;
  assign add_241730 = sel_241727 + 8'h01;
  assign sel_241731 = array_index_241642 == array_index_239448 ? add_241730 : sel_241727;
  assign add_241734 = sel_241731 + 8'h01;
  assign sel_241735 = array_index_241642 == array_index_239454 ? add_241734 : sel_241731;
  assign add_241738 = sel_241735 + 8'h01;
  assign sel_241739 = array_index_241642 == array_index_239460 ? add_241738 : sel_241735;
  assign add_241742 = sel_241739 + 8'h01;
  assign sel_241743 = array_index_241642 == array_index_239466 ? add_241742 : sel_241739;
  assign add_241746 = sel_241743 + 8'h01;
  assign sel_241747 = array_index_241642 == array_index_239472 ? add_241746 : sel_241743;
  assign add_241750 = sel_241747 + 8'h01;
  assign sel_241751 = array_index_241642 == array_index_239478 ? add_241750 : sel_241747;
  assign add_241754 = sel_241751 + 8'h01;
  assign sel_241755 = array_index_241642 == array_index_239484 ? add_241754 : sel_241751;
  assign add_241758 = sel_241755 + 8'h01;
  assign sel_241759 = array_index_241642 == array_index_239490 ? add_241758 : sel_241755;
  assign add_241762 = sel_241759 + 8'h01;
  assign sel_241763 = array_index_241642 == array_index_239496 ? add_241762 : sel_241759;
  assign add_241766 = sel_241763 + 8'h01;
  assign sel_241767 = array_index_241642 == array_index_239502 ? add_241766 : sel_241763;
  assign add_241770 = sel_241767 + 8'h01;
  assign sel_241771 = array_index_241642 == array_index_239508 ? add_241770 : sel_241767;
  assign add_241774 = sel_241771 + 8'h01;
  assign sel_241775 = array_index_241642 == array_index_239514 ? add_241774 : sel_241771;
  assign add_241778 = sel_241775 + 8'h01;
  assign sel_241779 = array_index_241642 == array_index_239520 ? add_241778 : sel_241775;
  assign add_241782 = sel_241779 + 8'h01;
  assign sel_241783 = array_index_241642 == array_index_239526 ? add_241782 : sel_241779;
  assign add_241786 = sel_241783 + 8'h01;
  assign sel_241787 = array_index_241642 == array_index_239532 ? add_241786 : sel_241783;
  assign add_241790 = sel_241787 + 8'h01;
  assign sel_241791 = array_index_241642 == array_index_239538 ? add_241790 : sel_241787;
  assign add_241794 = sel_241791 + 8'h01;
  assign sel_241795 = array_index_241642 == array_index_239544 ? add_241794 : sel_241791;
  assign add_241798 = sel_241795 + 8'h01;
  assign sel_241799 = array_index_241642 == array_index_239550 ? add_241798 : sel_241795;
  assign add_241802 = sel_241799 + 8'h01;
  assign sel_241803 = array_index_241642 == array_index_239556 ? add_241802 : sel_241799;
  assign add_241806 = sel_241803 + 8'h01;
  assign sel_241807 = array_index_241642 == array_index_239562 ? add_241806 : sel_241803;
  assign add_241810 = sel_241807 + 8'h01;
  assign sel_241811 = array_index_241642 == array_index_239568 ? add_241810 : sel_241807;
  assign add_241814 = sel_241811 + 8'h01;
  assign sel_241815 = array_index_241642 == array_index_239574 ? add_241814 : sel_241811;
  assign add_241818 = sel_241815 + 8'h01;
  assign sel_241819 = array_index_241642 == array_index_239580 ? add_241818 : sel_241815;
  assign add_241822 = sel_241819 + 8'h01;
  assign sel_241823 = array_index_241642 == array_index_239586 ? add_241822 : sel_241819;
  assign add_241826 = sel_241823 + 8'h01;
  assign sel_241827 = array_index_241642 == array_index_239592 ? add_241826 : sel_241823;
  assign add_241830 = sel_241827 + 8'h01;
  assign sel_241831 = array_index_241642 == array_index_239598 ? add_241830 : sel_241827;
  assign add_241834 = sel_241831 + 8'h01;
  assign sel_241835 = array_index_241642 == array_index_239604 ? add_241834 : sel_241831;
  assign add_241838 = sel_241835 + 8'h01;
  assign sel_241839 = array_index_241642 == array_index_239610 ? add_241838 : sel_241835;
  assign add_241843 = sel_241839 + 8'h01;
  assign array_index_241844 = set1_unflattened[6'h0c];
  assign sel_241845 = array_index_241642 == array_index_239616 ? add_241843 : sel_241839;
  assign add_241848 = sel_241845 + 8'h01;
  assign sel_241849 = array_index_241844 == array_index_239312 ? add_241848 : sel_241845;
  assign add_241852 = sel_241849 + 8'h01;
  assign sel_241853 = array_index_241844 == array_index_239316 ? add_241852 : sel_241849;
  assign add_241856 = sel_241853 + 8'h01;
  assign sel_241857 = array_index_241844 == array_index_239324 ? add_241856 : sel_241853;
  assign add_241860 = sel_241857 + 8'h01;
  assign sel_241861 = array_index_241844 == array_index_239332 ? add_241860 : sel_241857;
  assign add_241864 = sel_241861 + 8'h01;
  assign sel_241865 = array_index_241844 == array_index_239340 ? add_241864 : sel_241861;
  assign add_241868 = sel_241865 + 8'h01;
  assign sel_241869 = array_index_241844 == array_index_239348 ? add_241868 : sel_241865;
  assign add_241872 = sel_241869 + 8'h01;
  assign sel_241873 = array_index_241844 == array_index_239356 ? add_241872 : sel_241869;
  assign add_241876 = sel_241873 + 8'h01;
  assign sel_241877 = array_index_241844 == array_index_239364 ? add_241876 : sel_241873;
  assign add_241880 = sel_241877 + 8'h01;
  assign sel_241881 = array_index_241844 == array_index_239370 ? add_241880 : sel_241877;
  assign add_241884 = sel_241881 + 8'h01;
  assign sel_241885 = array_index_241844 == array_index_239376 ? add_241884 : sel_241881;
  assign add_241888 = sel_241885 + 8'h01;
  assign sel_241889 = array_index_241844 == array_index_239382 ? add_241888 : sel_241885;
  assign add_241892 = sel_241889 + 8'h01;
  assign sel_241893 = array_index_241844 == array_index_239388 ? add_241892 : sel_241889;
  assign add_241896 = sel_241893 + 8'h01;
  assign sel_241897 = array_index_241844 == array_index_239394 ? add_241896 : sel_241893;
  assign add_241900 = sel_241897 + 8'h01;
  assign sel_241901 = array_index_241844 == array_index_239400 ? add_241900 : sel_241897;
  assign add_241904 = sel_241901 + 8'h01;
  assign sel_241905 = array_index_241844 == array_index_239406 ? add_241904 : sel_241901;
  assign add_241908 = sel_241905 + 8'h01;
  assign sel_241909 = array_index_241844 == array_index_239412 ? add_241908 : sel_241905;
  assign add_241912 = sel_241909 + 8'h01;
  assign sel_241913 = array_index_241844 == array_index_239418 ? add_241912 : sel_241909;
  assign add_241916 = sel_241913 + 8'h01;
  assign sel_241917 = array_index_241844 == array_index_239424 ? add_241916 : sel_241913;
  assign add_241920 = sel_241917 + 8'h01;
  assign sel_241921 = array_index_241844 == array_index_239430 ? add_241920 : sel_241917;
  assign add_241924 = sel_241921 + 8'h01;
  assign sel_241925 = array_index_241844 == array_index_239436 ? add_241924 : sel_241921;
  assign add_241928 = sel_241925 + 8'h01;
  assign sel_241929 = array_index_241844 == array_index_239442 ? add_241928 : sel_241925;
  assign add_241932 = sel_241929 + 8'h01;
  assign sel_241933 = array_index_241844 == array_index_239448 ? add_241932 : sel_241929;
  assign add_241936 = sel_241933 + 8'h01;
  assign sel_241937 = array_index_241844 == array_index_239454 ? add_241936 : sel_241933;
  assign add_241940 = sel_241937 + 8'h01;
  assign sel_241941 = array_index_241844 == array_index_239460 ? add_241940 : sel_241937;
  assign add_241944 = sel_241941 + 8'h01;
  assign sel_241945 = array_index_241844 == array_index_239466 ? add_241944 : sel_241941;
  assign add_241948 = sel_241945 + 8'h01;
  assign sel_241949 = array_index_241844 == array_index_239472 ? add_241948 : sel_241945;
  assign add_241952 = sel_241949 + 8'h01;
  assign sel_241953 = array_index_241844 == array_index_239478 ? add_241952 : sel_241949;
  assign add_241956 = sel_241953 + 8'h01;
  assign sel_241957 = array_index_241844 == array_index_239484 ? add_241956 : sel_241953;
  assign add_241960 = sel_241957 + 8'h01;
  assign sel_241961 = array_index_241844 == array_index_239490 ? add_241960 : sel_241957;
  assign add_241964 = sel_241961 + 8'h01;
  assign sel_241965 = array_index_241844 == array_index_239496 ? add_241964 : sel_241961;
  assign add_241968 = sel_241965 + 8'h01;
  assign sel_241969 = array_index_241844 == array_index_239502 ? add_241968 : sel_241965;
  assign add_241972 = sel_241969 + 8'h01;
  assign sel_241973 = array_index_241844 == array_index_239508 ? add_241972 : sel_241969;
  assign add_241976 = sel_241973 + 8'h01;
  assign sel_241977 = array_index_241844 == array_index_239514 ? add_241976 : sel_241973;
  assign add_241980 = sel_241977 + 8'h01;
  assign sel_241981 = array_index_241844 == array_index_239520 ? add_241980 : sel_241977;
  assign add_241984 = sel_241981 + 8'h01;
  assign sel_241985 = array_index_241844 == array_index_239526 ? add_241984 : sel_241981;
  assign add_241988 = sel_241985 + 8'h01;
  assign sel_241989 = array_index_241844 == array_index_239532 ? add_241988 : sel_241985;
  assign add_241992 = sel_241989 + 8'h01;
  assign sel_241993 = array_index_241844 == array_index_239538 ? add_241992 : sel_241989;
  assign add_241996 = sel_241993 + 8'h01;
  assign sel_241997 = array_index_241844 == array_index_239544 ? add_241996 : sel_241993;
  assign add_242000 = sel_241997 + 8'h01;
  assign sel_242001 = array_index_241844 == array_index_239550 ? add_242000 : sel_241997;
  assign add_242004 = sel_242001 + 8'h01;
  assign sel_242005 = array_index_241844 == array_index_239556 ? add_242004 : sel_242001;
  assign add_242008 = sel_242005 + 8'h01;
  assign sel_242009 = array_index_241844 == array_index_239562 ? add_242008 : sel_242005;
  assign add_242012 = sel_242009 + 8'h01;
  assign sel_242013 = array_index_241844 == array_index_239568 ? add_242012 : sel_242009;
  assign add_242016 = sel_242013 + 8'h01;
  assign sel_242017 = array_index_241844 == array_index_239574 ? add_242016 : sel_242013;
  assign add_242020 = sel_242017 + 8'h01;
  assign sel_242021 = array_index_241844 == array_index_239580 ? add_242020 : sel_242017;
  assign add_242024 = sel_242021 + 8'h01;
  assign sel_242025 = array_index_241844 == array_index_239586 ? add_242024 : sel_242021;
  assign add_242028 = sel_242025 + 8'h01;
  assign sel_242029 = array_index_241844 == array_index_239592 ? add_242028 : sel_242025;
  assign add_242032 = sel_242029 + 8'h01;
  assign sel_242033 = array_index_241844 == array_index_239598 ? add_242032 : sel_242029;
  assign add_242036 = sel_242033 + 8'h01;
  assign sel_242037 = array_index_241844 == array_index_239604 ? add_242036 : sel_242033;
  assign add_242040 = sel_242037 + 8'h01;
  assign sel_242041 = array_index_241844 == array_index_239610 ? add_242040 : sel_242037;
  assign add_242045 = sel_242041 + 8'h01;
  assign array_index_242046 = set1_unflattened[6'h0d];
  assign sel_242047 = array_index_241844 == array_index_239616 ? add_242045 : sel_242041;
  assign add_242050 = sel_242047 + 8'h01;
  assign sel_242051 = array_index_242046 == array_index_239312 ? add_242050 : sel_242047;
  assign add_242054 = sel_242051 + 8'h01;
  assign sel_242055 = array_index_242046 == array_index_239316 ? add_242054 : sel_242051;
  assign add_242058 = sel_242055 + 8'h01;
  assign sel_242059 = array_index_242046 == array_index_239324 ? add_242058 : sel_242055;
  assign add_242062 = sel_242059 + 8'h01;
  assign sel_242063 = array_index_242046 == array_index_239332 ? add_242062 : sel_242059;
  assign add_242066 = sel_242063 + 8'h01;
  assign sel_242067 = array_index_242046 == array_index_239340 ? add_242066 : sel_242063;
  assign add_242070 = sel_242067 + 8'h01;
  assign sel_242071 = array_index_242046 == array_index_239348 ? add_242070 : sel_242067;
  assign add_242074 = sel_242071 + 8'h01;
  assign sel_242075 = array_index_242046 == array_index_239356 ? add_242074 : sel_242071;
  assign add_242078 = sel_242075 + 8'h01;
  assign sel_242079 = array_index_242046 == array_index_239364 ? add_242078 : sel_242075;
  assign add_242082 = sel_242079 + 8'h01;
  assign sel_242083 = array_index_242046 == array_index_239370 ? add_242082 : sel_242079;
  assign add_242086 = sel_242083 + 8'h01;
  assign sel_242087 = array_index_242046 == array_index_239376 ? add_242086 : sel_242083;
  assign add_242090 = sel_242087 + 8'h01;
  assign sel_242091 = array_index_242046 == array_index_239382 ? add_242090 : sel_242087;
  assign add_242094 = sel_242091 + 8'h01;
  assign sel_242095 = array_index_242046 == array_index_239388 ? add_242094 : sel_242091;
  assign add_242098 = sel_242095 + 8'h01;
  assign sel_242099 = array_index_242046 == array_index_239394 ? add_242098 : sel_242095;
  assign add_242102 = sel_242099 + 8'h01;
  assign sel_242103 = array_index_242046 == array_index_239400 ? add_242102 : sel_242099;
  assign add_242106 = sel_242103 + 8'h01;
  assign sel_242107 = array_index_242046 == array_index_239406 ? add_242106 : sel_242103;
  assign add_242110 = sel_242107 + 8'h01;
  assign sel_242111 = array_index_242046 == array_index_239412 ? add_242110 : sel_242107;
  assign add_242114 = sel_242111 + 8'h01;
  assign sel_242115 = array_index_242046 == array_index_239418 ? add_242114 : sel_242111;
  assign add_242118 = sel_242115 + 8'h01;
  assign sel_242119 = array_index_242046 == array_index_239424 ? add_242118 : sel_242115;
  assign add_242122 = sel_242119 + 8'h01;
  assign sel_242123 = array_index_242046 == array_index_239430 ? add_242122 : sel_242119;
  assign add_242126 = sel_242123 + 8'h01;
  assign sel_242127 = array_index_242046 == array_index_239436 ? add_242126 : sel_242123;
  assign add_242130 = sel_242127 + 8'h01;
  assign sel_242131 = array_index_242046 == array_index_239442 ? add_242130 : sel_242127;
  assign add_242134 = sel_242131 + 8'h01;
  assign sel_242135 = array_index_242046 == array_index_239448 ? add_242134 : sel_242131;
  assign add_242138 = sel_242135 + 8'h01;
  assign sel_242139 = array_index_242046 == array_index_239454 ? add_242138 : sel_242135;
  assign add_242142 = sel_242139 + 8'h01;
  assign sel_242143 = array_index_242046 == array_index_239460 ? add_242142 : sel_242139;
  assign add_242146 = sel_242143 + 8'h01;
  assign sel_242147 = array_index_242046 == array_index_239466 ? add_242146 : sel_242143;
  assign add_242150 = sel_242147 + 8'h01;
  assign sel_242151 = array_index_242046 == array_index_239472 ? add_242150 : sel_242147;
  assign add_242154 = sel_242151 + 8'h01;
  assign sel_242155 = array_index_242046 == array_index_239478 ? add_242154 : sel_242151;
  assign add_242158 = sel_242155 + 8'h01;
  assign sel_242159 = array_index_242046 == array_index_239484 ? add_242158 : sel_242155;
  assign add_242162 = sel_242159 + 8'h01;
  assign sel_242163 = array_index_242046 == array_index_239490 ? add_242162 : sel_242159;
  assign add_242166 = sel_242163 + 8'h01;
  assign sel_242167 = array_index_242046 == array_index_239496 ? add_242166 : sel_242163;
  assign add_242170 = sel_242167 + 8'h01;
  assign sel_242171 = array_index_242046 == array_index_239502 ? add_242170 : sel_242167;
  assign add_242174 = sel_242171 + 8'h01;
  assign sel_242175 = array_index_242046 == array_index_239508 ? add_242174 : sel_242171;
  assign add_242178 = sel_242175 + 8'h01;
  assign sel_242179 = array_index_242046 == array_index_239514 ? add_242178 : sel_242175;
  assign add_242182 = sel_242179 + 8'h01;
  assign sel_242183 = array_index_242046 == array_index_239520 ? add_242182 : sel_242179;
  assign add_242186 = sel_242183 + 8'h01;
  assign sel_242187 = array_index_242046 == array_index_239526 ? add_242186 : sel_242183;
  assign add_242190 = sel_242187 + 8'h01;
  assign sel_242191 = array_index_242046 == array_index_239532 ? add_242190 : sel_242187;
  assign add_242194 = sel_242191 + 8'h01;
  assign sel_242195 = array_index_242046 == array_index_239538 ? add_242194 : sel_242191;
  assign add_242198 = sel_242195 + 8'h01;
  assign sel_242199 = array_index_242046 == array_index_239544 ? add_242198 : sel_242195;
  assign add_242202 = sel_242199 + 8'h01;
  assign sel_242203 = array_index_242046 == array_index_239550 ? add_242202 : sel_242199;
  assign add_242206 = sel_242203 + 8'h01;
  assign sel_242207 = array_index_242046 == array_index_239556 ? add_242206 : sel_242203;
  assign add_242210 = sel_242207 + 8'h01;
  assign sel_242211 = array_index_242046 == array_index_239562 ? add_242210 : sel_242207;
  assign add_242214 = sel_242211 + 8'h01;
  assign sel_242215 = array_index_242046 == array_index_239568 ? add_242214 : sel_242211;
  assign add_242218 = sel_242215 + 8'h01;
  assign sel_242219 = array_index_242046 == array_index_239574 ? add_242218 : sel_242215;
  assign add_242222 = sel_242219 + 8'h01;
  assign sel_242223 = array_index_242046 == array_index_239580 ? add_242222 : sel_242219;
  assign add_242226 = sel_242223 + 8'h01;
  assign sel_242227 = array_index_242046 == array_index_239586 ? add_242226 : sel_242223;
  assign add_242230 = sel_242227 + 8'h01;
  assign sel_242231 = array_index_242046 == array_index_239592 ? add_242230 : sel_242227;
  assign add_242234 = sel_242231 + 8'h01;
  assign sel_242235 = array_index_242046 == array_index_239598 ? add_242234 : sel_242231;
  assign add_242238 = sel_242235 + 8'h01;
  assign sel_242239 = array_index_242046 == array_index_239604 ? add_242238 : sel_242235;
  assign add_242242 = sel_242239 + 8'h01;
  assign sel_242243 = array_index_242046 == array_index_239610 ? add_242242 : sel_242239;
  assign add_242247 = sel_242243 + 8'h01;
  assign array_index_242248 = set1_unflattened[6'h0e];
  assign sel_242249 = array_index_242046 == array_index_239616 ? add_242247 : sel_242243;
  assign add_242252 = sel_242249 + 8'h01;
  assign sel_242253 = array_index_242248 == array_index_239312 ? add_242252 : sel_242249;
  assign add_242256 = sel_242253 + 8'h01;
  assign sel_242257 = array_index_242248 == array_index_239316 ? add_242256 : sel_242253;
  assign add_242260 = sel_242257 + 8'h01;
  assign sel_242261 = array_index_242248 == array_index_239324 ? add_242260 : sel_242257;
  assign add_242264 = sel_242261 + 8'h01;
  assign sel_242265 = array_index_242248 == array_index_239332 ? add_242264 : sel_242261;
  assign add_242268 = sel_242265 + 8'h01;
  assign sel_242269 = array_index_242248 == array_index_239340 ? add_242268 : sel_242265;
  assign add_242272 = sel_242269 + 8'h01;
  assign sel_242273 = array_index_242248 == array_index_239348 ? add_242272 : sel_242269;
  assign add_242276 = sel_242273 + 8'h01;
  assign sel_242277 = array_index_242248 == array_index_239356 ? add_242276 : sel_242273;
  assign add_242280 = sel_242277 + 8'h01;
  assign sel_242281 = array_index_242248 == array_index_239364 ? add_242280 : sel_242277;
  assign add_242284 = sel_242281 + 8'h01;
  assign sel_242285 = array_index_242248 == array_index_239370 ? add_242284 : sel_242281;
  assign add_242288 = sel_242285 + 8'h01;
  assign sel_242289 = array_index_242248 == array_index_239376 ? add_242288 : sel_242285;
  assign add_242292 = sel_242289 + 8'h01;
  assign sel_242293 = array_index_242248 == array_index_239382 ? add_242292 : sel_242289;
  assign add_242296 = sel_242293 + 8'h01;
  assign sel_242297 = array_index_242248 == array_index_239388 ? add_242296 : sel_242293;
  assign add_242300 = sel_242297 + 8'h01;
  assign sel_242301 = array_index_242248 == array_index_239394 ? add_242300 : sel_242297;
  assign add_242304 = sel_242301 + 8'h01;
  assign sel_242305 = array_index_242248 == array_index_239400 ? add_242304 : sel_242301;
  assign add_242308 = sel_242305 + 8'h01;
  assign sel_242309 = array_index_242248 == array_index_239406 ? add_242308 : sel_242305;
  assign add_242312 = sel_242309 + 8'h01;
  assign sel_242313 = array_index_242248 == array_index_239412 ? add_242312 : sel_242309;
  assign add_242316 = sel_242313 + 8'h01;
  assign sel_242317 = array_index_242248 == array_index_239418 ? add_242316 : sel_242313;
  assign add_242320 = sel_242317 + 8'h01;
  assign sel_242321 = array_index_242248 == array_index_239424 ? add_242320 : sel_242317;
  assign add_242324 = sel_242321 + 8'h01;
  assign sel_242325 = array_index_242248 == array_index_239430 ? add_242324 : sel_242321;
  assign add_242328 = sel_242325 + 8'h01;
  assign sel_242329 = array_index_242248 == array_index_239436 ? add_242328 : sel_242325;
  assign add_242332 = sel_242329 + 8'h01;
  assign sel_242333 = array_index_242248 == array_index_239442 ? add_242332 : sel_242329;
  assign add_242336 = sel_242333 + 8'h01;
  assign sel_242337 = array_index_242248 == array_index_239448 ? add_242336 : sel_242333;
  assign add_242340 = sel_242337 + 8'h01;
  assign sel_242341 = array_index_242248 == array_index_239454 ? add_242340 : sel_242337;
  assign add_242344 = sel_242341 + 8'h01;
  assign sel_242345 = array_index_242248 == array_index_239460 ? add_242344 : sel_242341;
  assign add_242348 = sel_242345 + 8'h01;
  assign sel_242349 = array_index_242248 == array_index_239466 ? add_242348 : sel_242345;
  assign add_242352 = sel_242349 + 8'h01;
  assign sel_242353 = array_index_242248 == array_index_239472 ? add_242352 : sel_242349;
  assign add_242356 = sel_242353 + 8'h01;
  assign sel_242357 = array_index_242248 == array_index_239478 ? add_242356 : sel_242353;
  assign add_242360 = sel_242357 + 8'h01;
  assign sel_242361 = array_index_242248 == array_index_239484 ? add_242360 : sel_242357;
  assign add_242364 = sel_242361 + 8'h01;
  assign sel_242365 = array_index_242248 == array_index_239490 ? add_242364 : sel_242361;
  assign add_242368 = sel_242365 + 8'h01;
  assign sel_242369 = array_index_242248 == array_index_239496 ? add_242368 : sel_242365;
  assign add_242372 = sel_242369 + 8'h01;
  assign sel_242373 = array_index_242248 == array_index_239502 ? add_242372 : sel_242369;
  assign add_242376 = sel_242373 + 8'h01;
  assign sel_242377 = array_index_242248 == array_index_239508 ? add_242376 : sel_242373;
  assign add_242380 = sel_242377 + 8'h01;
  assign sel_242381 = array_index_242248 == array_index_239514 ? add_242380 : sel_242377;
  assign add_242384 = sel_242381 + 8'h01;
  assign sel_242385 = array_index_242248 == array_index_239520 ? add_242384 : sel_242381;
  assign add_242388 = sel_242385 + 8'h01;
  assign sel_242389 = array_index_242248 == array_index_239526 ? add_242388 : sel_242385;
  assign add_242392 = sel_242389 + 8'h01;
  assign sel_242393 = array_index_242248 == array_index_239532 ? add_242392 : sel_242389;
  assign add_242396 = sel_242393 + 8'h01;
  assign sel_242397 = array_index_242248 == array_index_239538 ? add_242396 : sel_242393;
  assign add_242400 = sel_242397 + 8'h01;
  assign sel_242401 = array_index_242248 == array_index_239544 ? add_242400 : sel_242397;
  assign add_242404 = sel_242401 + 8'h01;
  assign sel_242405 = array_index_242248 == array_index_239550 ? add_242404 : sel_242401;
  assign add_242408 = sel_242405 + 8'h01;
  assign sel_242409 = array_index_242248 == array_index_239556 ? add_242408 : sel_242405;
  assign add_242412 = sel_242409 + 8'h01;
  assign sel_242413 = array_index_242248 == array_index_239562 ? add_242412 : sel_242409;
  assign add_242416 = sel_242413 + 8'h01;
  assign sel_242417 = array_index_242248 == array_index_239568 ? add_242416 : sel_242413;
  assign add_242420 = sel_242417 + 8'h01;
  assign sel_242421 = array_index_242248 == array_index_239574 ? add_242420 : sel_242417;
  assign add_242424 = sel_242421 + 8'h01;
  assign sel_242425 = array_index_242248 == array_index_239580 ? add_242424 : sel_242421;
  assign add_242428 = sel_242425 + 8'h01;
  assign sel_242429 = array_index_242248 == array_index_239586 ? add_242428 : sel_242425;
  assign add_242432 = sel_242429 + 8'h01;
  assign sel_242433 = array_index_242248 == array_index_239592 ? add_242432 : sel_242429;
  assign add_242436 = sel_242433 + 8'h01;
  assign sel_242437 = array_index_242248 == array_index_239598 ? add_242436 : sel_242433;
  assign add_242440 = sel_242437 + 8'h01;
  assign sel_242441 = array_index_242248 == array_index_239604 ? add_242440 : sel_242437;
  assign add_242444 = sel_242441 + 8'h01;
  assign sel_242445 = array_index_242248 == array_index_239610 ? add_242444 : sel_242441;
  assign add_242449 = sel_242445 + 8'h01;
  assign array_index_242450 = set1_unflattened[6'h0f];
  assign sel_242451 = array_index_242248 == array_index_239616 ? add_242449 : sel_242445;
  assign add_242454 = sel_242451 + 8'h01;
  assign sel_242455 = array_index_242450 == array_index_239312 ? add_242454 : sel_242451;
  assign add_242458 = sel_242455 + 8'h01;
  assign sel_242459 = array_index_242450 == array_index_239316 ? add_242458 : sel_242455;
  assign add_242462 = sel_242459 + 8'h01;
  assign sel_242463 = array_index_242450 == array_index_239324 ? add_242462 : sel_242459;
  assign add_242466 = sel_242463 + 8'h01;
  assign sel_242467 = array_index_242450 == array_index_239332 ? add_242466 : sel_242463;
  assign add_242470 = sel_242467 + 8'h01;
  assign sel_242471 = array_index_242450 == array_index_239340 ? add_242470 : sel_242467;
  assign add_242474 = sel_242471 + 8'h01;
  assign sel_242475 = array_index_242450 == array_index_239348 ? add_242474 : sel_242471;
  assign add_242478 = sel_242475 + 8'h01;
  assign sel_242479 = array_index_242450 == array_index_239356 ? add_242478 : sel_242475;
  assign add_242482 = sel_242479 + 8'h01;
  assign sel_242483 = array_index_242450 == array_index_239364 ? add_242482 : sel_242479;
  assign add_242486 = sel_242483 + 8'h01;
  assign sel_242487 = array_index_242450 == array_index_239370 ? add_242486 : sel_242483;
  assign add_242490 = sel_242487 + 8'h01;
  assign sel_242491 = array_index_242450 == array_index_239376 ? add_242490 : sel_242487;
  assign add_242494 = sel_242491 + 8'h01;
  assign sel_242495 = array_index_242450 == array_index_239382 ? add_242494 : sel_242491;
  assign add_242498 = sel_242495 + 8'h01;
  assign sel_242499 = array_index_242450 == array_index_239388 ? add_242498 : sel_242495;
  assign add_242502 = sel_242499 + 8'h01;
  assign sel_242503 = array_index_242450 == array_index_239394 ? add_242502 : sel_242499;
  assign add_242506 = sel_242503 + 8'h01;
  assign sel_242507 = array_index_242450 == array_index_239400 ? add_242506 : sel_242503;
  assign add_242510 = sel_242507 + 8'h01;
  assign sel_242511 = array_index_242450 == array_index_239406 ? add_242510 : sel_242507;
  assign add_242514 = sel_242511 + 8'h01;
  assign sel_242515 = array_index_242450 == array_index_239412 ? add_242514 : sel_242511;
  assign add_242518 = sel_242515 + 8'h01;
  assign sel_242519 = array_index_242450 == array_index_239418 ? add_242518 : sel_242515;
  assign add_242522 = sel_242519 + 8'h01;
  assign sel_242523 = array_index_242450 == array_index_239424 ? add_242522 : sel_242519;
  assign add_242526 = sel_242523 + 8'h01;
  assign sel_242527 = array_index_242450 == array_index_239430 ? add_242526 : sel_242523;
  assign add_242530 = sel_242527 + 8'h01;
  assign sel_242531 = array_index_242450 == array_index_239436 ? add_242530 : sel_242527;
  assign add_242534 = sel_242531 + 8'h01;
  assign sel_242535 = array_index_242450 == array_index_239442 ? add_242534 : sel_242531;
  assign add_242538 = sel_242535 + 8'h01;
  assign sel_242539 = array_index_242450 == array_index_239448 ? add_242538 : sel_242535;
  assign add_242542 = sel_242539 + 8'h01;
  assign sel_242543 = array_index_242450 == array_index_239454 ? add_242542 : sel_242539;
  assign add_242546 = sel_242543 + 8'h01;
  assign sel_242547 = array_index_242450 == array_index_239460 ? add_242546 : sel_242543;
  assign add_242550 = sel_242547 + 8'h01;
  assign sel_242551 = array_index_242450 == array_index_239466 ? add_242550 : sel_242547;
  assign add_242554 = sel_242551 + 8'h01;
  assign sel_242555 = array_index_242450 == array_index_239472 ? add_242554 : sel_242551;
  assign add_242558 = sel_242555 + 8'h01;
  assign sel_242559 = array_index_242450 == array_index_239478 ? add_242558 : sel_242555;
  assign add_242562 = sel_242559 + 8'h01;
  assign sel_242563 = array_index_242450 == array_index_239484 ? add_242562 : sel_242559;
  assign add_242566 = sel_242563 + 8'h01;
  assign sel_242567 = array_index_242450 == array_index_239490 ? add_242566 : sel_242563;
  assign add_242570 = sel_242567 + 8'h01;
  assign sel_242571 = array_index_242450 == array_index_239496 ? add_242570 : sel_242567;
  assign add_242574 = sel_242571 + 8'h01;
  assign sel_242575 = array_index_242450 == array_index_239502 ? add_242574 : sel_242571;
  assign add_242578 = sel_242575 + 8'h01;
  assign sel_242579 = array_index_242450 == array_index_239508 ? add_242578 : sel_242575;
  assign add_242582 = sel_242579 + 8'h01;
  assign sel_242583 = array_index_242450 == array_index_239514 ? add_242582 : sel_242579;
  assign add_242586 = sel_242583 + 8'h01;
  assign sel_242587 = array_index_242450 == array_index_239520 ? add_242586 : sel_242583;
  assign add_242590 = sel_242587 + 8'h01;
  assign sel_242591 = array_index_242450 == array_index_239526 ? add_242590 : sel_242587;
  assign add_242594 = sel_242591 + 8'h01;
  assign sel_242595 = array_index_242450 == array_index_239532 ? add_242594 : sel_242591;
  assign add_242598 = sel_242595 + 8'h01;
  assign sel_242599 = array_index_242450 == array_index_239538 ? add_242598 : sel_242595;
  assign add_242602 = sel_242599 + 8'h01;
  assign sel_242603 = array_index_242450 == array_index_239544 ? add_242602 : sel_242599;
  assign add_242606 = sel_242603 + 8'h01;
  assign sel_242607 = array_index_242450 == array_index_239550 ? add_242606 : sel_242603;
  assign add_242610 = sel_242607 + 8'h01;
  assign sel_242611 = array_index_242450 == array_index_239556 ? add_242610 : sel_242607;
  assign add_242614 = sel_242611 + 8'h01;
  assign sel_242615 = array_index_242450 == array_index_239562 ? add_242614 : sel_242611;
  assign add_242618 = sel_242615 + 8'h01;
  assign sel_242619 = array_index_242450 == array_index_239568 ? add_242618 : sel_242615;
  assign add_242622 = sel_242619 + 8'h01;
  assign sel_242623 = array_index_242450 == array_index_239574 ? add_242622 : sel_242619;
  assign add_242626 = sel_242623 + 8'h01;
  assign sel_242627 = array_index_242450 == array_index_239580 ? add_242626 : sel_242623;
  assign add_242630 = sel_242627 + 8'h01;
  assign sel_242631 = array_index_242450 == array_index_239586 ? add_242630 : sel_242627;
  assign add_242634 = sel_242631 + 8'h01;
  assign sel_242635 = array_index_242450 == array_index_239592 ? add_242634 : sel_242631;
  assign add_242638 = sel_242635 + 8'h01;
  assign sel_242639 = array_index_242450 == array_index_239598 ? add_242638 : sel_242635;
  assign add_242642 = sel_242639 + 8'h01;
  assign sel_242643 = array_index_242450 == array_index_239604 ? add_242642 : sel_242639;
  assign add_242646 = sel_242643 + 8'h01;
  assign sel_242647 = array_index_242450 == array_index_239610 ? add_242646 : sel_242643;
  assign add_242651 = sel_242647 + 8'h01;
  assign array_index_242652 = set1_unflattened[6'h10];
  assign sel_242653 = array_index_242450 == array_index_239616 ? add_242651 : sel_242647;
  assign add_242656 = sel_242653 + 8'h01;
  assign sel_242657 = array_index_242652 == array_index_239312 ? add_242656 : sel_242653;
  assign add_242660 = sel_242657 + 8'h01;
  assign sel_242661 = array_index_242652 == array_index_239316 ? add_242660 : sel_242657;
  assign add_242664 = sel_242661 + 8'h01;
  assign sel_242665 = array_index_242652 == array_index_239324 ? add_242664 : sel_242661;
  assign add_242668 = sel_242665 + 8'h01;
  assign sel_242669 = array_index_242652 == array_index_239332 ? add_242668 : sel_242665;
  assign add_242672 = sel_242669 + 8'h01;
  assign sel_242673 = array_index_242652 == array_index_239340 ? add_242672 : sel_242669;
  assign add_242676 = sel_242673 + 8'h01;
  assign sel_242677 = array_index_242652 == array_index_239348 ? add_242676 : sel_242673;
  assign add_242680 = sel_242677 + 8'h01;
  assign sel_242681 = array_index_242652 == array_index_239356 ? add_242680 : sel_242677;
  assign add_242684 = sel_242681 + 8'h01;
  assign sel_242685 = array_index_242652 == array_index_239364 ? add_242684 : sel_242681;
  assign add_242688 = sel_242685 + 8'h01;
  assign sel_242689 = array_index_242652 == array_index_239370 ? add_242688 : sel_242685;
  assign add_242692 = sel_242689 + 8'h01;
  assign sel_242693 = array_index_242652 == array_index_239376 ? add_242692 : sel_242689;
  assign add_242696 = sel_242693 + 8'h01;
  assign sel_242697 = array_index_242652 == array_index_239382 ? add_242696 : sel_242693;
  assign add_242700 = sel_242697 + 8'h01;
  assign sel_242701 = array_index_242652 == array_index_239388 ? add_242700 : sel_242697;
  assign add_242704 = sel_242701 + 8'h01;
  assign sel_242705 = array_index_242652 == array_index_239394 ? add_242704 : sel_242701;
  assign add_242708 = sel_242705 + 8'h01;
  assign sel_242709 = array_index_242652 == array_index_239400 ? add_242708 : sel_242705;
  assign add_242712 = sel_242709 + 8'h01;
  assign sel_242713 = array_index_242652 == array_index_239406 ? add_242712 : sel_242709;
  assign add_242716 = sel_242713 + 8'h01;
  assign sel_242717 = array_index_242652 == array_index_239412 ? add_242716 : sel_242713;
  assign add_242720 = sel_242717 + 8'h01;
  assign sel_242721 = array_index_242652 == array_index_239418 ? add_242720 : sel_242717;
  assign add_242724 = sel_242721 + 8'h01;
  assign sel_242725 = array_index_242652 == array_index_239424 ? add_242724 : sel_242721;
  assign add_242728 = sel_242725 + 8'h01;
  assign sel_242729 = array_index_242652 == array_index_239430 ? add_242728 : sel_242725;
  assign add_242732 = sel_242729 + 8'h01;
  assign sel_242733 = array_index_242652 == array_index_239436 ? add_242732 : sel_242729;
  assign add_242736 = sel_242733 + 8'h01;
  assign sel_242737 = array_index_242652 == array_index_239442 ? add_242736 : sel_242733;
  assign add_242740 = sel_242737 + 8'h01;
  assign sel_242741 = array_index_242652 == array_index_239448 ? add_242740 : sel_242737;
  assign add_242744 = sel_242741 + 8'h01;
  assign sel_242745 = array_index_242652 == array_index_239454 ? add_242744 : sel_242741;
  assign add_242748 = sel_242745 + 8'h01;
  assign sel_242749 = array_index_242652 == array_index_239460 ? add_242748 : sel_242745;
  assign add_242752 = sel_242749 + 8'h01;
  assign sel_242753 = array_index_242652 == array_index_239466 ? add_242752 : sel_242749;
  assign add_242756 = sel_242753 + 8'h01;
  assign sel_242757 = array_index_242652 == array_index_239472 ? add_242756 : sel_242753;
  assign add_242760 = sel_242757 + 8'h01;
  assign sel_242761 = array_index_242652 == array_index_239478 ? add_242760 : sel_242757;
  assign add_242764 = sel_242761 + 8'h01;
  assign sel_242765 = array_index_242652 == array_index_239484 ? add_242764 : sel_242761;
  assign add_242768 = sel_242765 + 8'h01;
  assign sel_242769 = array_index_242652 == array_index_239490 ? add_242768 : sel_242765;
  assign add_242772 = sel_242769 + 8'h01;
  assign sel_242773 = array_index_242652 == array_index_239496 ? add_242772 : sel_242769;
  assign add_242776 = sel_242773 + 8'h01;
  assign sel_242777 = array_index_242652 == array_index_239502 ? add_242776 : sel_242773;
  assign add_242780 = sel_242777 + 8'h01;
  assign sel_242781 = array_index_242652 == array_index_239508 ? add_242780 : sel_242777;
  assign add_242784 = sel_242781 + 8'h01;
  assign sel_242785 = array_index_242652 == array_index_239514 ? add_242784 : sel_242781;
  assign add_242788 = sel_242785 + 8'h01;
  assign sel_242789 = array_index_242652 == array_index_239520 ? add_242788 : sel_242785;
  assign add_242792 = sel_242789 + 8'h01;
  assign sel_242793 = array_index_242652 == array_index_239526 ? add_242792 : sel_242789;
  assign add_242796 = sel_242793 + 8'h01;
  assign sel_242797 = array_index_242652 == array_index_239532 ? add_242796 : sel_242793;
  assign add_242800 = sel_242797 + 8'h01;
  assign sel_242801 = array_index_242652 == array_index_239538 ? add_242800 : sel_242797;
  assign add_242804 = sel_242801 + 8'h01;
  assign sel_242805 = array_index_242652 == array_index_239544 ? add_242804 : sel_242801;
  assign add_242808 = sel_242805 + 8'h01;
  assign sel_242809 = array_index_242652 == array_index_239550 ? add_242808 : sel_242805;
  assign add_242812 = sel_242809 + 8'h01;
  assign sel_242813 = array_index_242652 == array_index_239556 ? add_242812 : sel_242809;
  assign add_242816 = sel_242813 + 8'h01;
  assign sel_242817 = array_index_242652 == array_index_239562 ? add_242816 : sel_242813;
  assign add_242820 = sel_242817 + 8'h01;
  assign sel_242821 = array_index_242652 == array_index_239568 ? add_242820 : sel_242817;
  assign add_242824 = sel_242821 + 8'h01;
  assign sel_242825 = array_index_242652 == array_index_239574 ? add_242824 : sel_242821;
  assign add_242828 = sel_242825 + 8'h01;
  assign sel_242829 = array_index_242652 == array_index_239580 ? add_242828 : sel_242825;
  assign add_242832 = sel_242829 + 8'h01;
  assign sel_242833 = array_index_242652 == array_index_239586 ? add_242832 : sel_242829;
  assign add_242836 = sel_242833 + 8'h01;
  assign sel_242837 = array_index_242652 == array_index_239592 ? add_242836 : sel_242833;
  assign add_242840 = sel_242837 + 8'h01;
  assign sel_242841 = array_index_242652 == array_index_239598 ? add_242840 : sel_242837;
  assign add_242844 = sel_242841 + 8'h01;
  assign sel_242845 = array_index_242652 == array_index_239604 ? add_242844 : sel_242841;
  assign add_242848 = sel_242845 + 8'h01;
  assign sel_242849 = array_index_242652 == array_index_239610 ? add_242848 : sel_242845;
  assign add_242853 = sel_242849 + 8'h01;
  assign array_index_242854 = set1_unflattened[6'h11];
  assign sel_242855 = array_index_242652 == array_index_239616 ? add_242853 : sel_242849;
  assign add_242858 = sel_242855 + 8'h01;
  assign sel_242859 = array_index_242854 == array_index_239312 ? add_242858 : sel_242855;
  assign add_242862 = sel_242859 + 8'h01;
  assign sel_242863 = array_index_242854 == array_index_239316 ? add_242862 : sel_242859;
  assign add_242866 = sel_242863 + 8'h01;
  assign sel_242867 = array_index_242854 == array_index_239324 ? add_242866 : sel_242863;
  assign add_242870 = sel_242867 + 8'h01;
  assign sel_242871 = array_index_242854 == array_index_239332 ? add_242870 : sel_242867;
  assign add_242874 = sel_242871 + 8'h01;
  assign sel_242875 = array_index_242854 == array_index_239340 ? add_242874 : sel_242871;
  assign add_242878 = sel_242875 + 8'h01;
  assign sel_242879 = array_index_242854 == array_index_239348 ? add_242878 : sel_242875;
  assign add_242882 = sel_242879 + 8'h01;
  assign sel_242883 = array_index_242854 == array_index_239356 ? add_242882 : sel_242879;
  assign add_242886 = sel_242883 + 8'h01;
  assign sel_242887 = array_index_242854 == array_index_239364 ? add_242886 : sel_242883;
  assign add_242890 = sel_242887 + 8'h01;
  assign sel_242891 = array_index_242854 == array_index_239370 ? add_242890 : sel_242887;
  assign add_242894 = sel_242891 + 8'h01;
  assign sel_242895 = array_index_242854 == array_index_239376 ? add_242894 : sel_242891;
  assign add_242898 = sel_242895 + 8'h01;
  assign sel_242899 = array_index_242854 == array_index_239382 ? add_242898 : sel_242895;
  assign add_242902 = sel_242899 + 8'h01;
  assign sel_242903 = array_index_242854 == array_index_239388 ? add_242902 : sel_242899;
  assign add_242906 = sel_242903 + 8'h01;
  assign sel_242907 = array_index_242854 == array_index_239394 ? add_242906 : sel_242903;
  assign add_242910 = sel_242907 + 8'h01;
  assign sel_242911 = array_index_242854 == array_index_239400 ? add_242910 : sel_242907;
  assign add_242914 = sel_242911 + 8'h01;
  assign sel_242915 = array_index_242854 == array_index_239406 ? add_242914 : sel_242911;
  assign add_242918 = sel_242915 + 8'h01;
  assign sel_242919 = array_index_242854 == array_index_239412 ? add_242918 : sel_242915;
  assign add_242922 = sel_242919 + 8'h01;
  assign sel_242923 = array_index_242854 == array_index_239418 ? add_242922 : sel_242919;
  assign add_242926 = sel_242923 + 8'h01;
  assign sel_242927 = array_index_242854 == array_index_239424 ? add_242926 : sel_242923;
  assign add_242930 = sel_242927 + 8'h01;
  assign sel_242931 = array_index_242854 == array_index_239430 ? add_242930 : sel_242927;
  assign add_242934 = sel_242931 + 8'h01;
  assign sel_242935 = array_index_242854 == array_index_239436 ? add_242934 : sel_242931;
  assign add_242938 = sel_242935 + 8'h01;
  assign sel_242939 = array_index_242854 == array_index_239442 ? add_242938 : sel_242935;
  assign add_242942 = sel_242939 + 8'h01;
  assign sel_242943 = array_index_242854 == array_index_239448 ? add_242942 : sel_242939;
  assign add_242946 = sel_242943 + 8'h01;
  assign sel_242947 = array_index_242854 == array_index_239454 ? add_242946 : sel_242943;
  assign add_242950 = sel_242947 + 8'h01;
  assign sel_242951 = array_index_242854 == array_index_239460 ? add_242950 : sel_242947;
  assign add_242954 = sel_242951 + 8'h01;
  assign sel_242955 = array_index_242854 == array_index_239466 ? add_242954 : sel_242951;
  assign add_242958 = sel_242955 + 8'h01;
  assign sel_242959 = array_index_242854 == array_index_239472 ? add_242958 : sel_242955;
  assign add_242962 = sel_242959 + 8'h01;
  assign sel_242963 = array_index_242854 == array_index_239478 ? add_242962 : sel_242959;
  assign add_242966 = sel_242963 + 8'h01;
  assign sel_242967 = array_index_242854 == array_index_239484 ? add_242966 : sel_242963;
  assign add_242970 = sel_242967 + 8'h01;
  assign sel_242971 = array_index_242854 == array_index_239490 ? add_242970 : sel_242967;
  assign add_242974 = sel_242971 + 8'h01;
  assign sel_242975 = array_index_242854 == array_index_239496 ? add_242974 : sel_242971;
  assign add_242978 = sel_242975 + 8'h01;
  assign sel_242979 = array_index_242854 == array_index_239502 ? add_242978 : sel_242975;
  assign add_242982 = sel_242979 + 8'h01;
  assign sel_242983 = array_index_242854 == array_index_239508 ? add_242982 : sel_242979;
  assign add_242986 = sel_242983 + 8'h01;
  assign sel_242987 = array_index_242854 == array_index_239514 ? add_242986 : sel_242983;
  assign add_242990 = sel_242987 + 8'h01;
  assign sel_242991 = array_index_242854 == array_index_239520 ? add_242990 : sel_242987;
  assign add_242994 = sel_242991 + 8'h01;
  assign sel_242995 = array_index_242854 == array_index_239526 ? add_242994 : sel_242991;
  assign add_242998 = sel_242995 + 8'h01;
  assign sel_242999 = array_index_242854 == array_index_239532 ? add_242998 : sel_242995;
  assign add_243002 = sel_242999 + 8'h01;
  assign sel_243003 = array_index_242854 == array_index_239538 ? add_243002 : sel_242999;
  assign add_243006 = sel_243003 + 8'h01;
  assign sel_243007 = array_index_242854 == array_index_239544 ? add_243006 : sel_243003;
  assign add_243010 = sel_243007 + 8'h01;
  assign sel_243011 = array_index_242854 == array_index_239550 ? add_243010 : sel_243007;
  assign add_243014 = sel_243011 + 8'h01;
  assign sel_243015 = array_index_242854 == array_index_239556 ? add_243014 : sel_243011;
  assign add_243018 = sel_243015 + 8'h01;
  assign sel_243019 = array_index_242854 == array_index_239562 ? add_243018 : sel_243015;
  assign add_243022 = sel_243019 + 8'h01;
  assign sel_243023 = array_index_242854 == array_index_239568 ? add_243022 : sel_243019;
  assign add_243026 = sel_243023 + 8'h01;
  assign sel_243027 = array_index_242854 == array_index_239574 ? add_243026 : sel_243023;
  assign add_243030 = sel_243027 + 8'h01;
  assign sel_243031 = array_index_242854 == array_index_239580 ? add_243030 : sel_243027;
  assign add_243034 = sel_243031 + 8'h01;
  assign sel_243035 = array_index_242854 == array_index_239586 ? add_243034 : sel_243031;
  assign add_243038 = sel_243035 + 8'h01;
  assign sel_243039 = array_index_242854 == array_index_239592 ? add_243038 : sel_243035;
  assign add_243042 = sel_243039 + 8'h01;
  assign sel_243043 = array_index_242854 == array_index_239598 ? add_243042 : sel_243039;
  assign add_243046 = sel_243043 + 8'h01;
  assign sel_243047 = array_index_242854 == array_index_239604 ? add_243046 : sel_243043;
  assign add_243050 = sel_243047 + 8'h01;
  assign sel_243051 = array_index_242854 == array_index_239610 ? add_243050 : sel_243047;
  assign add_243055 = sel_243051 + 8'h01;
  assign array_index_243056 = set1_unflattened[6'h12];
  assign sel_243057 = array_index_242854 == array_index_239616 ? add_243055 : sel_243051;
  assign add_243060 = sel_243057 + 8'h01;
  assign sel_243061 = array_index_243056 == array_index_239312 ? add_243060 : sel_243057;
  assign add_243064 = sel_243061 + 8'h01;
  assign sel_243065 = array_index_243056 == array_index_239316 ? add_243064 : sel_243061;
  assign add_243068 = sel_243065 + 8'h01;
  assign sel_243069 = array_index_243056 == array_index_239324 ? add_243068 : sel_243065;
  assign add_243072 = sel_243069 + 8'h01;
  assign sel_243073 = array_index_243056 == array_index_239332 ? add_243072 : sel_243069;
  assign add_243076 = sel_243073 + 8'h01;
  assign sel_243077 = array_index_243056 == array_index_239340 ? add_243076 : sel_243073;
  assign add_243080 = sel_243077 + 8'h01;
  assign sel_243081 = array_index_243056 == array_index_239348 ? add_243080 : sel_243077;
  assign add_243084 = sel_243081 + 8'h01;
  assign sel_243085 = array_index_243056 == array_index_239356 ? add_243084 : sel_243081;
  assign add_243088 = sel_243085 + 8'h01;
  assign sel_243089 = array_index_243056 == array_index_239364 ? add_243088 : sel_243085;
  assign add_243092 = sel_243089 + 8'h01;
  assign sel_243093 = array_index_243056 == array_index_239370 ? add_243092 : sel_243089;
  assign add_243096 = sel_243093 + 8'h01;
  assign sel_243097 = array_index_243056 == array_index_239376 ? add_243096 : sel_243093;
  assign add_243100 = sel_243097 + 8'h01;
  assign sel_243101 = array_index_243056 == array_index_239382 ? add_243100 : sel_243097;
  assign add_243104 = sel_243101 + 8'h01;
  assign sel_243105 = array_index_243056 == array_index_239388 ? add_243104 : sel_243101;
  assign add_243108 = sel_243105 + 8'h01;
  assign sel_243109 = array_index_243056 == array_index_239394 ? add_243108 : sel_243105;
  assign add_243112 = sel_243109 + 8'h01;
  assign sel_243113 = array_index_243056 == array_index_239400 ? add_243112 : sel_243109;
  assign add_243116 = sel_243113 + 8'h01;
  assign sel_243117 = array_index_243056 == array_index_239406 ? add_243116 : sel_243113;
  assign add_243120 = sel_243117 + 8'h01;
  assign sel_243121 = array_index_243056 == array_index_239412 ? add_243120 : sel_243117;
  assign add_243124 = sel_243121 + 8'h01;
  assign sel_243125 = array_index_243056 == array_index_239418 ? add_243124 : sel_243121;
  assign add_243128 = sel_243125 + 8'h01;
  assign sel_243129 = array_index_243056 == array_index_239424 ? add_243128 : sel_243125;
  assign add_243132 = sel_243129 + 8'h01;
  assign sel_243133 = array_index_243056 == array_index_239430 ? add_243132 : sel_243129;
  assign add_243136 = sel_243133 + 8'h01;
  assign sel_243137 = array_index_243056 == array_index_239436 ? add_243136 : sel_243133;
  assign add_243140 = sel_243137 + 8'h01;
  assign sel_243141 = array_index_243056 == array_index_239442 ? add_243140 : sel_243137;
  assign add_243144 = sel_243141 + 8'h01;
  assign sel_243145 = array_index_243056 == array_index_239448 ? add_243144 : sel_243141;
  assign add_243148 = sel_243145 + 8'h01;
  assign sel_243149 = array_index_243056 == array_index_239454 ? add_243148 : sel_243145;
  assign add_243152 = sel_243149 + 8'h01;
  assign sel_243153 = array_index_243056 == array_index_239460 ? add_243152 : sel_243149;
  assign add_243156 = sel_243153 + 8'h01;
  assign sel_243157 = array_index_243056 == array_index_239466 ? add_243156 : sel_243153;
  assign add_243160 = sel_243157 + 8'h01;
  assign sel_243161 = array_index_243056 == array_index_239472 ? add_243160 : sel_243157;
  assign add_243164 = sel_243161 + 8'h01;
  assign sel_243165 = array_index_243056 == array_index_239478 ? add_243164 : sel_243161;
  assign add_243168 = sel_243165 + 8'h01;
  assign sel_243169 = array_index_243056 == array_index_239484 ? add_243168 : sel_243165;
  assign add_243172 = sel_243169 + 8'h01;
  assign sel_243173 = array_index_243056 == array_index_239490 ? add_243172 : sel_243169;
  assign add_243176 = sel_243173 + 8'h01;
  assign sel_243177 = array_index_243056 == array_index_239496 ? add_243176 : sel_243173;
  assign add_243180 = sel_243177 + 8'h01;
  assign sel_243181 = array_index_243056 == array_index_239502 ? add_243180 : sel_243177;
  assign add_243184 = sel_243181 + 8'h01;
  assign sel_243185 = array_index_243056 == array_index_239508 ? add_243184 : sel_243181;
  assign add_243188 = sel_243185 + 8'h01;
  assign sel_243189 = array_index_243056 == array_index_239514 ? add_243188 : sel_243185;
  assign add_243192 = sel_243189 + 8'h01;
  assign sel_243193 = array_index_243056 == array_index_239520 ? add_243192 : sel_243189;
  assign add_243196 = sel_243193 + 8'h01;
  assign sel_243197 = array_index_243056 == array_index_239526 ? add_243196 : sel_243193;
  assign add_243200 = sel_243197 + 8'h01;
  assign sel_243201 = array_index_243056 == array_index_239532 ? add_243200 : sel_243197;
  assign add_243204 = sel_243201 + 8'h01;
  assign sel_243205 = array_index_243056 == array_index_239538 ? add_243204 : sel_243201;
  assign add_243208 = sel_243205 + 8'h01;
  assign sel_243209 = array_index_243056 == array_index_239544 ? add_243208 : sel_243205;
  assign add_243212 = sel_243209 + 8'h01;
  assign sel_243213 = array_index_243056 == array_index_239550 ? add_243212 : sel_243209;
  assign add_243216 = sel_243213 + 8'h01;
  assign sel_243217 = array_index_243056 == array_index_239556 ? add_243216 : sel_243213;
  assign add_243220 = sel_243217 + 8'h01;
  assign sel_243221 = array_index_243056 == array_index_239562 ? add_243220 : sel_243217;
  assign add_243224 = sel_243221 + 8'h01;
  assign sel_243225 = array_index_243056 == array_index_239568 ? add_243224 : sel_243221;
  assign add_243228 = sel_243225 + 8'h01;
  assign sel_243229 = array_index_243056 == array_index_239574 ? add_243228 : sel_243225;
  assign add_243232 = sel_243229 + 8'h01;
  assign sel_243233 = array_index_243056 == array_index_239580 ? add_243232 : sel_243229;
  assign add_243236 = sel_243233 + 8'h01;
  assign sel_243237 = array_index_243056 == array_index_239586 ? add_243236 : sel_243233;
  assign add_243240 = sel_243237 + 8'h01;
  assign sel_243241 = array_index_243056 == array_index_239592 ? add_243240 : sel_243237;
  assign add_243244 = sel_243241 + 8'h01;
  assign sel_243245 = array_index_243056 == array_index_239598 ? add_243244 : sel_243241;
  assign add_243248 = sel_243245 + 8'h01;
  assign sel_243249 = array_index_243056 == array_index_239604 ? add_243248 : sel_243245;
  assign add_243252 = sel_243249 + 8'h01;
  assign sel_243253 = array_index_243056 == array_index_239610 ? add_243252 : sel_243249;
  assign add_243257 = sel_243253 + 8'h01;
  assign array_index_243258 = set1_unflattened[6'h13];
  assign sel_243259 = array_index_243056 == array_index_239616 ? add_243257 : sel_243253;
  assign add_243262 = sel_243259 + 8'h01;
  assign sel_243263 = array_index_243258 == array_index_239312 ? add_243262 : sel_243259;
  assign add_243266 = sel_243263 + 8'h01;
  assign sel_243267 = array_index_243258 == array_index_239316 ? add_243266 : sel_243263;
  assign add_243270 = sel_243267 + 8'h01;
  assign sel_243271 = array_index_243258 == array_index_239324 ? add_243270 : sel_243267;
  assign add_243274 = sel_243271 + 8'h01;
  assign sel_243275 = array_index_243258 == array_index_239332 ? add_243274 : sel_243271;
  assign add_243278 = sel_243275 + 8'h01;
  assign sel_243279 = array_index_243258 == array_index_239340 ? add_243278 : sel_243275;
  assign add_243282 = sel_243279 + 8'h01;
  assign sel_243283 = array_index_243258 == array_index_239348 ? add_243282 : sel_243279;
  assign add_243286 = sel_243283 + 8'h01;
  assign sel_243287 = array_index_243258 == array_index_239356 ? add_243286 : sel_243283;
  assign add_243290 = sel_243287 + 8'h01;
  assign sel_243291 = array_index_243258 == array_index_239364 ? add_243290 : sel_243287;
  assign add_243294 = sel_243291 + 8'h01;
  assign sel_243295 = array_index_243258 == array_index_239370 ? add_243294 : sel_243291;
  assign add_243298 = sel_243295 + 8'h01;
  assign sel_243299 = array_index_243258 == array_index_239376 ? add_243298 : sel_243295;
  assign add_243302 = sel_243299 + 8'h01;
  assign sel_243303 = array_index_243258 == array_index_239382 ? add_243302 : sel_243299;
  assign add_243306 = sel_243303 + 8'h01;
  assign sel_243307 = array_index_243258 == array_index_239388 ? add_243306 : sel_243303;
  assign add_243310 = sel_243307 + 8'h01;
  assign sel_243311 = array_index_243258 == array_index_239394 ? add_243310 : sel_243307;
  assign add_243314 = sel_243311 + 8'h01;
  assign sel_243315 = array_index_243258 == array_index_239400 ? add_243314 : sel_243311;
  assign add_243318 = sel_243315 + 8'h01;
  assign sel_243319 = array_index_243258 == array_index_239406 ? add_243318 : sel_243315;
  assign add_243322 = sel_243319 + 8'h01;
  assign sel_243323 = array_index_243258 == array_index_239412 ? add_243322 : sel_243319;
  assign add_243326 = sel_243323 + 8'h01;
  assign sel_243327 = array_index_243258 == array_index_239418 ? add_243326 : sel_243323;
  assign add_243330 = sel_243327 + 8'h01;
  assign sel_243331 = array_index_243258 == array_index_239424 ? add_243330 : sel_243327;
  assign add_243334 = sel_243331 + 8'h01;
  assign sel_243335 = array_index_243258 == array_index_239430 ? add_243334 : sel_243331;
  assign add_243338 = sel_243335 + 8'h01;
  assign sel_243339 = array_index_243258 == array_index_239436 ? add_243338 : sel_243335;
  assign add_243342 = sel_243339 + 8'h01;
  assign sel_243343 = array_index_243258 == array_index_239442 ? add_243342 : sel_243339;
  assign add_243346 = sel_243343 + 8'h01;
  assign sel_243347 = array_index_243258 == array_index_239448 ? add_243346 : sel_243343;
  assign add_243350 = sel_243347 + 8'h01;
  assign sel_243351 = array_index_243258 == array_index_239454 ? add_243350 : sel_243347;
  assign add_243354 = sel_243351 + 8'h01;
  assign sel_243355 = array_index_243258 == array_index_239460 ? add_243354 : sel_243351;
  assign add_243358 = sel_243355 + 8'h01;
  assign sel_243359 = array_index_243258 == array_index_239466 ? add_243358 : sel_243355;
  assign add_243362 = sel_243359 + 8'h01;
  assign sel_243363 = array_index_243258 == array_index_239472 ? add_243362 : sel_243359;
  assign add_243366 = sel_243363 + 8'h01;
  assign sel_243367 = array_index_243258 == array_index_239478 ? add_243366 : sel_243363;
  assign add_243370 = sel_243367 + 8'h01;
  assign sel_243371 = array_index_243258 == array_index_239484 ? add_243370 : sel_243367;
  assign add_243374 = sel_243371 + 8'h01;
  assign sel_243375 = array_index_243258 == array_index_239490 ? add_243374 : sel_243371;
  assign add_243378 = sel_243375 + 8'h01;
  assign sel_243379 = array_index_243258 == array_index_239496 ? add_243378 : sel_243375;
  assign add_243382 = sel_243379 + 8'h01;
  assign sel_243383 = array_index_243258 == array_index_239502 ? add_243382 : sel_243379;
  assign add_243386 = sel_243383 + 8'h01;
  assign sel_243387 = array_index_243258 == array_index_239508 ? add_243386 : sel_243383;
  assign add_243390 = sel_243387 + 8'h01;
  assign sel_243391 = array_index_243258 == array_index_239514 ? add_243390 : sel_243387;
  assign add_243394 = sel_243391 + 8'h01;
  assign sel_243395 = array_index_243258 == array_index_239520 ? add_243394 : sel_243391;
  assign add_243398 = sel_243395 + 8'h01;
  assign sel_243399 = array_index_243258 == array_index_239526 ? add_243398 : sel_243395;
  assign add_243402 = sel_243399 + 8'h01;
  assign sel_243403 = array_index_243258 == array_index_239532 ? add_243402 : sel_243399;
  assign add_243406 = sel_243403 + 8'h01;
  assign sel_243407 = array_index_243258 == array_index_239538 ? add_243406 : sel_243403;
  assign add_243410 = sel_243407 + 8'h01;
  assign sel_243411 = array_index_243258 == array_index_239544 ? add_243410 : sel_243407;
  assign add_243414 = sel_243411 + 8'h01;
  assign sel_243415 = array_index_243258 == array_index_239550 ? add_243414 : sel_243411;
  assign add_243418 = sel_243415 + 8'h01;
  assign sel_243419 = array_index_243258 == array_index_239556 ? add_243418 : sel_243415;
  assign add_243422 = sel_243419 + 8'h01;
  assign sel_243423 = array_index_243258 == array_index_239562 ? add_243422 : sel_243419;
  assign add_243426 = sel_243423 + 8'h01;
  assign sel_243427 = array_index_243258 == array_index_239568 ? add_243426 : sel_243423;
  assign add_243430 = sel_243427 + 8'h01;
  assign sel_243431 = array_index_243258 == array_index_239574 ? add_243430 : sel_243427;
  assign add_243434 = sel_243431 + 8'h01;
  assign sel_243435 = array_index_243258 == array_index_239580 ? add_243434 : sel_243431;
  assign add_243438 = sel_243435 + 8'h01;
  assign sel_243439 = array_index_243258 == array_index_239586 ? add_243438 : sel_243435;
  assign add_243442 = sel_243439 + 8'h01;
  assign sel_243443 = array_index_243258 == array_index_239592 ? add_243442 : sel_243439;
  assign add_243446 = sel_243443 + 8'h01;
  assign sel_243447 = array_index_243258 == array_index_239598 ? add_243446 : sel_243443;
  assign add_243450 = sel_243447 + 8'h01;
  assign sel_243451 = array_index_243258 == array_index_239604 ? add_243450 : sel_243447;
  assign add_243454 = sel_243451 + 8'h01;
  assign sel_243455 = array_index_243258 == array_index_239610 ? add_243454 : sel_243451;
  assign add_243459 = sel_243455 + 8'h01;
  assign array_index_243460 = set1_unflattened[6'h14];
  assign sel_243461 = array_index_243258 == array_index_239616 ? add_243459 : sel_243455;
  assign add_243464 = sel_243461 + 8'h01;
  assign sel_243465 = array_index_243460 == array_index_239312 ? add_243464 : sel_243461;
  assign add_243468 = sel_243465 + 8'h01;
  assign sel_243469 = array_index_243460 == array_index_239316 ? add_243468 : sel_243465;
  assign add_243472 = sel_243469 + 8'h01;
  assign sel_243473 = array_index_243460 == array_index_239324 ? add_243472 : sel_243469;
  assign add_243476 = sel_243473 + 8'h01;
  assign sel_243477 = array_index_243460 == array_index_239332 ? add_243476 : sel_243473;
  assign add_243480 = sel_243477 + 8'h01;
  assign sel_243481 = array_index_243460 == array_index_239340 ? add_243480 : sel_243477;
  assign add_243484 = sel_243481 + 8'h01;
  assign sel_243485 = array_index_243460 == array_index_239348 ? add_243484 : sel_243481;
  assign add_243488 = sel_243485 + 8'h01;
  assign sel_243489 = array_index_243460 == array_index_239356 ? add_243488 : sel_243485;
  assign add_243492 = sel_243489 + 8'h01;
  assign sel_243493 = array_index_243460 == array_index_239364 ? add_243492 : sel_243489;
  assign add_243496 = sel_243493 + 8'h01;
  assign sel_243497 = array_index_243460 == array_index_239370 ? add_243496 : sel_243493;
  assign add_243500 = sel_243497 + 8'h01;
  assign sel_243501 = array_index_243460 == array_index_239376 ? add_243500 : sel_243497;
  assign add_243504 = sel_243501 + 8'h01;
  assign sel_243505 = array_index_243460 == array_index_239382 ? add_243504 : sel_243501;
  assign add_243508 = sel_243505 + 8'h01;
  assign sel_243509 = array_index_243460 == array_index_239388 ? add_243508 : sel_243505;
  assign add_243512 = sel_243509 + 8'h01;
  assign sel_243513 = array_index_243460 == array_index_239394 ? add_243512 : sel_243509;
  assign add_243516 = sel_243513 + 8'h01;
  assign sel_243517 = array_index_243460 == array_index_239400 ? add_243516 : sel_243513;
  assign add_243520 = sel_243517 + 8'h01;
  assign sel_243521 = array_index_243460 == array_index_239406 ? add_243520 : sel_243517;
  assign add_243524 = sel_243521 + 8'h01;
  assign sel_243525 = array_index_243460 == array_index_239412 ? add_243524 : sel_243521;
  assign add_243528 = sel_243525 + 8'h01;
  assign sel_243529 = array_index_243460 == array_index_239418 ? add_243528 : sel_243525;
  assign add_243532 = sel_243529 + 8'h01;
  assign sel_243533 = array_index_243460 == array_index_239424 ? add_243532 : sel_243529;
  assign add_243536 = sel_243533 + 8'h01;
  assign sel_243537 = array_index_243460 == array_index_239430 ? add_243536 : sel_243533;
  assign add_243540 = sel_243537 + 8'h01;
  assign sel_243541 = array_index_243460 == array_index_239436 ? add_243540 : sel_243537;
  assign add_243544 = sel_243541 + 8'h01;
  assign sel_243545 = array_index_243460 == array_index_239442 ? add_243544 : sel_243541;
  assign add_243548 = sel_243545 + 8'h01;
  assign sel_243549 = array_index_243460 == array_index_239448 ? add_243548 : sel_243545;
  assign add_243552 = sel_243549 + 8'h01;
  assign sel_243553 = array_index_243460 == array_index_239454 ? add_243552 : sel_243549;
  assign add_243556 = sel_243553 + 8'h01;
  assign sel_243557 = array_index_243460 == array_index_239460 ? add_243556 : sel_243553;
  assign add_243560 = sel_243557 + 8'h01;
  assign sel_243561 = array_index_243460 == array_index_239466 ? add_243560 : sel_243557;
  assign add_243564 = sel_243561 + 8'h01;
  assign sel_243565 = array_index_243460 == array_index_239472 ? add_243564 : sel_243561;
  assign add_243568 = sel_243565 + 8'h01;
  assign sel_243569 = array_index_243460 == array_index_239478 ? add_243568 : sel_243565;
  assign add_243572 = sel_243569 + 8'h01;
  assign sel_243573 = array_index_243460 == array_index_239484 ? add_243572 : sel_243569;
  assign add_243576 = sel_243573 + 8'h01;
  assign sel_243577 = array_index_243460 == array_index_239490 ? add_243576 : sel_243573;
  assign add_243580 = sel_243577 + 8'h01;
  assign sel_243581 = array_index_243460 == array_index_239496 ? add_243580 : sel_243577;
  assign add_243584 = sel_243581 + 8'h01;
  assign sel_243585 = array_index_243460 == array_index_239502 ? add_243584 : sel_243581;
  assign add_243588 = sel_243585 + 8'h01;
  assign sel_243589 = array_index_243460 == array_index_239508 ? add_243588 : sel_243585;
  assign add_243592 = sel_243589 + 8'h01;
  assign sel_243593 = array_index_243460 == array_index_239514 ? add_243592 : sel_243589;
  assign add_243596 = sel_243593 + 8'h01;
  assign sel_243597 = array_index_243460 == array_index_239520 ? add_243596 : sel_243593;
  assign add_243600 = sel_243597 + 8'h01;
  assign sel_243601 = array_index_243460 == array_index_239526 ? add_243600 : sel_243597;
  assign add_243604 = sel_243601 + 8'h01;
  assign sel_243605 = array_index_243460 == array_index_239532 ? add_243604 : sel_243601;
  assign add_243608 = sel_243605 + 8'h01;
  assign sel_243609 = array_index_243460 == array_index_239538 ? add_243608 : sel_243605;
  assign add_243612 = sel_243609 + 8'h01;
  assign sel_243613 = array_index_243460 == array_index_239544 ? add_243612 : sel_243609;
  assign add_243616 = sel_243613 + 8'h01;
  assign sel_243617 = array_index_243460 == array_index_239550 ? add_243616 : sel_243613;
  assign add_243620 = sel_243617 + 8'h01;
  assign sel_243621 = array_index_243460 == array_index_239556 ? add_243620 : sel_243617;
  assign add_243624 = sel_243621 + 8'h01;
  assign sel_243625 = array_index_243460 == array_index_239562 ? add_243624 : sel_243621;
  assign add_243628 = sel_243625 + 8'h01;
  assign sel_243629 = array_index_243460 == array_index_239568 ? add_243628 : sel_243625;
  assign add_243632 = sel_243629 + 8'h01;
  assign sel_243633 = array_index_243460 == array_index_239574 ? add_243632 : sel_243629;
  assign add_243636 = sel_243633 + 8'h01;
  assign sel_243637 = array_index_243460 == array_index_239580 ? add_243636 : sel_243633;
  assign add_243640 = sel_243637 + 8'h01;
  assign sel_243641 = array_index_243460 == array_index_239586 ? add_243640 : sel_243637;
  assign add_243644 = sel_243641 + 8'h01;
  assign sel_243645 = array_index_243460 == array_index_239592 ? add_243644 : sel_243641;
  assign add_243648 = sel_243645 + 8'h01;
  assign sel_243649 = array_index_243460 == array_index_239598 ? add_243648 : sel_243645;
  assign add_243652 = sel_243649 + 8'h01;
  assign sel_243653 = array_index_243460 == array_index_239604 ? add_243652 : sel_243649;
  assign add_243656 = sel_243653 + 8'h01;
  assign sel_243657 = array_index_243460 == array_index_239610 ? add_243656 : sel_243653;
  assign add_243661 = sel_243657 + 8'h01;
  assign array_index_243662 = set1_unflattened[6'h15];
  assign sel_243663 = array_index_243460 == array_index_239616 ? add_243661 : sel_243657;
  assign add_243666 = sel_243663 + 8'h01;
  assign sel_243667 = array_index_243662 == array_index_239312 ? add_243666 : sel_243663;
  assign add_243670 = sel_243667 + 8'h01;
  assign sel_243671 = array_index_243662 == array_index_239316 ? add_243670 : sel_243667;
  assign add_243674 = sel_243671 + 8'h01;
  assign sel_243675 = array_index_243662 == array_index_239324 ? add_243674 : sel_243671;
  assign add_243678 = sel_243675 + 8'h01;
  assign sel_243679 = array_index_243662 == array_index_239332 ? add_243678 : sel_243675;
  assign add_243682 = sel_243679 + 8'h01;
  assign sel_243683 = array_index_243662 == array_index_239340 ? add_243682 : sel_243679;
  assign add_243686 = sel_243683 + 8'h01;
  assign sel_243687 = array_index_243662 == array_index_239348 ? add_243686 : sel_243683;
  assign add_243690 = sel_243687 + 8'h01;
  assign sel_243691 = array_index_243662 == array_index_239356 ? add_243690 : sel_243687;
  assign add_243694 = sel_243691 + 8'h01;
  assign sel_243695 = array_index_243662 == array_index_239364 ? add_243694 : sel_243691;
  assign add_243698 = sel_243695 + 8'h01;
  assign sel_243699 = array_index_243662 == array_index_239370 ? add_243698 : sel_243695;
  assign add_243702 = sel_243699 + 8'h01;
  assign sel_243703 = array_index_243662 == array_index_239376 ? add_243702 : sel_243699;
  assign add_243706 = sel_243703 + 8'h01;
  assign sel_243707 = array_index_243662 == array_index_239382 ? add_243706 : sel_243703;
  assign add_243710 = sel_243707 + 8'h01;
  assign sel_243711 = array_index_243662 == array_index_239388 ? add_243710 : sel_243707;
  assign add_243714 = sel_243711 + 8'h01;
  assign sel_243715 = array_index_243662 == array_index_239394 ? add_243714 : sel_243711;
  assign add_243718 = sel_243715 + 8'h01;
  assign sel_243719 = array_index_243662 == array_index_239400 ? add_243718 : sel_243715;
  assign add_243722 = sel_243719 + 8'h01;
  assign sel_243723 = array_index_243662 == array_index_239406 ? add_243722 : sel_243719;
  assign add_243726 = sel_243723 + 8'h01;
  assign sel_243727 = array_index_243662 == array_index_239412 ? add_243726 : sel_243723;
  assign add_243730 = sel_243727 + 8'h01;
  assign sel_243731 = array_index_243662 == array_index_239418 ? add_243730 : sel_243727;
  assign add_243734 = sel_243731 + 8'h01;
  assign sel_243735 = array_index_243662 == array_index_239424 ? add_243734 : sel_243731;
  assign add_243738 = sel_243735 + 8'h01;
  assign sel_243739 = array_index_243662 == array_index_239430 ? add_243738 : sel_243735;
  assign add_243742 = sel_243739 + 8'h01;
  assign sel_243743 = array_index_243662 == array_index_239436 ? add_243742 : sel_243739;
  assign add_243746 = sel_243743 + 8'h01;
  assign sel_243747 = array_index_243662 == array_index_239442 ? add_243746 : sel_243743;
  assign add_243750 = sel_243747 + 8'h01;
  assign sel_243751 = array_index_243662 == array_index_239448 ? add_243750 : sel_243747;
  assign add_243754 = sel_243751 + 8'h01;
  assign sel_243755 = array_index_243662 == array_index_239454 ? add_243754 : sel_243751;
  assign add_243758 = sel_243755 + 8'h01;
  assign sel_243759 = array_index_243662 == array_index_239460 ? add_243758 : sel_243755;
  assign add_243762 = sel_243759 + 8'h01;
  assign sel_243763 = array_index_243662 == array_index_239466 ? add_243762 : sel_243759;
  assign add_243766 = sel_243763 + 8'h01;
  assign sel_243767 = array_index_243662 == array_index_239472 ? add_243766 : sel_243763;
  assign add_243770 = sel_243767 + 8'h01;
  assign sel_243771 = array_index_243662 == array_index_239478 ? add_243770 : sel_243767;
  assign add_243774 = sel_243771 + 8'h01;
  assign sel_243775 = array_index_243662 == array_index_239484 ? add_243774 : sel_243771;
  assign add_243778 = sel_243775 + 8'h01;
  assign sel_243779 = array_index_243662 == array_index_239490 ? add_243778 : sel_243775;
  assign add_243782 = sel_243779 + 8'h01;
  assign sel_243783 = array_index_243662 == array_index_239496 ? add_243782 : sel_243779;
  assign add_243786 = sel_243783 + 8'h01;
  assign sel_243787 = array_index_243662 == array_index_239502 ? add_243786 : sel_243783;
  assign add_243790 = sel_243787 + 8'h01;
  assign sel_243791 = array_index_243662 == array_index_239508 ? add_243790 : sel_243787;
  assign add_243794 = sel_243791 + 8'h01;
  assign sel_243795 = array_index_243662 == array_index_239514 ? add_243794 : sel_243791;
  assign add_243798 = sel_243795 + 8'h01;
  assign sel_243799 = array_index_243662 == array_index_239520 ? add_243798 : sel_243795;
  assign add_243802 = sel_243799 + 8'h01;
  assign sel_243803 = array_index_243662 == array_index_239526 ? add_243802 : sel_243799;
  assign add_243806 = sel_243803 + 8'h01;
  assign sel_243807 = array_index_243662 == array_index_239532 ? add_243806 : sel_243803;
  assign add_243810 = sel_243807 + 8'h01;
  assign sel_243811 = array_index_243662 == array_index_239538 ? add_243810 : sel_243807;
  assign add_243814 = sel_243811 + 8'h01;
  assign sel_243815 = array_index_243662 == array_index_239544 ? add_243814 : sel_243811;
  assign add_243818 = sel_243815 + 8'h01;
  assign sel_243819 = array_index_243662 == array_index_239550 ? add_243818 : sel_243815;
  assign add_243822 = sel_243819 + 8'h01;
  assign sel_243823 = array_index_243662 == array_index_239556 ? add_243822 : sel_243819;
  assign add_243826 = sel_243823 + 8'h01;
  assign sel_243827 = array_index_243662 == array_index_239562 ? add_243826 : sel_243823;
  assign add_243830 = sel_243827 + 8'h01;
  assign sel_243831 = array_index_243662 == array_index_239568 ? add_243830 : sel_243827;
  assign add_243834 = sel_243831 + 8'h01;
  assign sel_243835 = array_index_243662 == array_index_239574 ? add_243834 : sel_243831;
  assign add_243838 = sel_243835 + 8'h01;
  assign sel_243839 = array_index_243662 == array_index_239580 ? add_243838 : sel_243835;
  assign add_243842 = sel_243839 + 8'h01;
  assign sel_243843 = array_index_243662 == array_index_239586 ? add_243842 : sel_243839;
  assign add_243846 = sel_243843 + 8'h01;
  assign sel_243847 = array_index_243662 == array_index_239592 ? add_243846 : sel_243843;
  assign add_243850 = sel_243847 + 8'h01;
  assign sel_243851 = array_index_243662 == array_index_239598 ? add_243850 : sel_243847;
  assign add_243854 = sel_243851 + 8'h01;
  assign sel_243855 = array_index_243662 == array_index_239604 ? add_243854 : sel_243851;
  assign add_243858 = sel_243855 + 8'h01;
  assign sel_243859 = array_index_243662 == array_index_239610 ? add_243858 : sel_243855;
  assign add_243863 = sel_243859 + 8'h01;
  assign array_index_243864 = set1_unflattened[6'h16];
  assign sel_243865 = array_index_243662 == array_index_239616 ? add_243863 : sel_243859;
  assign add_243868 = sel_243865 + 8'h01;
  assign sel_243869 = array_index_243864 == array_index_239312 ? add_243868 : sel_243865;
  assign add_243872 = sel_243869 + 8'h01;
  assign sel_243873 = array_index_243864 == array_index_239316 ? add_243872 : sel_243869;
  assign add_243876 = sel_243873 + 8'h01;
  assign sel_243877 = array_index_243864 == array_index_239324 ? add_243876 : sel_243873;
  assign add_243880 = sel_243877 + 8'h01;
  assign sel_243881 = array_index_243864 == array_index_239332 ? add_243880 : sel_243877;
  assign add_243884 = sel_243881 + 8'h01;
  assign sel_243885 = array_index_243864 == array_index_239340 ? add_243884 : sel_243881;
  assign add_243888 = sel_243885 + 8'h01;
  assign sel_243889 = array_index_243864 == array_index_239348 ? add_243888 : sel_243885;
  assign add_243892 = sel_243889 + 8'h01;
  assign sel_243893 = array_index_243864 == array_index_239356 ? add_243892 : sel_243889;
  assign add_243896 = sel_243893 + 8'h01;
  assign sel_243897 = array_index_243864 == array_index_239364 ? add_243896 : sel_243893;
  assign add_243900 = sel_243897 + 8'h01;
  assign sel_243901 = array_index_243864 == array_index_239370 ? add_243900 : sel_243897;
  assign add_243904 = sel_243901 + 8'h01;
  assign sel_243905 = array_index_243864 == array_index_239376 ? add_243904 : sel_243901;
  assign add_243908 = sel_243905 + 8'h01;
  assign sel_243909 = array_index_243864 == array_index_239382 ? add_243908 : sel_243905;
  assign add_243912 = sel_243909 + 8'h01;
  assign sel_243913 = array_index_243864 == array_index_239388 ? add_243912 : sel_243909;
  assign add_243916 = sel_243913 + 8'h01;
  assign sel_243917 = array_index_243864 == array_index_239394 ? add_243916 : sel_243913;
  assign add_243920 = sel_243917 + 8'h01;
  assign sel_243921 = array_index_243864 == array_index_239400 ? add_243920 : sel_243917;
  assign add_243924 = sel_243921 + 8'h01;
  assign sel_243925 = array_index_243864 == array_index_239406 ? add_243924 : sel_243921;
  assign add_243928 = sel_243925 + 8'h01;
  assign sel_243929 = array_index_243864 == array_index_239412 ? add_243928 : sel_243925;
  assign add_243932 = sel_243929 + 8'h01;
  assign sel_243933 = array_index_243864 == array_index_239418 ? add_243932 : sel_243929;
  assign add_243936 = sel_243933 + 8'h01;
  assign sel_243937 = array_index_243864 == array_index_239424 ? add_243936 : sel_243933;
  assign add_243940 = sel_243937 + 8'h01;
  assign sel_243941 = array_index_243864 == array_index_239430 ? add_243940 : sel_243937;
  assign add_243944 = sel_243941 + 8'h01;
  assign sel_243945 = array_index_243864 == array_index_239436 ? add_243944 : sel_243941;
  assign add_243948 = sel_243945 + 8'h01;
  assign sel_243949 = array_index_243864 == array_index_239442 ? add_243948 : sel_243945;
  assign add_243952 = sel_243949 + 8'h01;
  assign sel_243953 = array_index_243864 == array_index_239448 ? add_243952 : sel_243949;
  assign add_243956 = sel_243953 + 8'h01;
  assign sel_243957 = array_index_243864 == array_index_239454 ? add_243956 : sel_243953;
  assign add_243960 = sel_243957 + 8'h01;
  assign sel_243961 = array_index_243864 == array_index_239460 ? add_243960 : sel_243957;
  assign add_243964 = sel_243961 + 8'h01;
  assign sel_243965 = array_index_243864 == array_index_239466 ? add_243964 : sel_243961;
  assign add_243968 = sel_243965 + 8'h01;
  assign sel_243969 = array_index_243864 == array_index_239472 ? add_243968 : sel_243965;
  assign add_243972 = sel_243969 + 8'h01;
  assign sel_243973 = array_index_243864 == array_index_239478 ? add_243972 : sel_243969;
  assign add_243976 = sel_243973 + 8'h01;
  assign sel_243977 = array_index_243864 == array_index_239484 ? add_243976 : sel_243973;
  assign add_243980 = sel_243977 + 8'h01;
  assign sel_243981 = array_index_243864 == array_index_239490 ? add_243980 : sel_243977;
  assign add_243984 = sel_243981 + 8'h01;
  assign sel_243985 = array_index_243864 == array_index_239496 ? add_243984 : sel_243981;
  assign add_243988 = sel_243985 + 8'h01;
  assign sel_243989 = array_index_243864 == array_index_239502 ? add_243988 : sel_243985;
  assign add_243992 = sel_243989 + 8'h01;
  assign sel_243993 = array_index_243864 == array_index_239508 ? add_243992 : sel_243989;
  assign add_243996 = sel_243993 + 8'h01;
  assign sel_243997 = array_index_243864 == array_index_239514 ? add_243996 : sel_243993;
  assign add_244000 = sel_243997 + 8'h01;
  assign sel_244001 = array_index_243864 == array_index_239520 ? add_244000 : sel_243997;
  assign add_244004 = sel_244001 + 8'h01;
  assign sel_244005 = array_index_243864 == array_index_239526 ? add_244004 : sel_244001;
  assign add_244008 = sel_244005 + 8'h01;
  assign sel_244009 = array_index_243864 == array_index_239532 ? add_244008 : sel_244005;
  assign add_244012 = sel_244009 + 8'h01;
  assign sel_244013 = array_index_243864 == array_index_239538 ? add_244012 : sel_244009;
  assign add_244016 = sel_244013 + 8'h01;
  assign sel_244017 = array_index_243864 == array_index_239544 ? add_244016 : sel_244013;
  assign add_244020 = sel_244017 + 8'h01;
  assign sel_244021 = array_index_243864 == array_index_239550 ? add_244020 : sel_244017;
  assign add_244024 = sel_244021 + 8'h01;
  assign sel_244025 = array_index_243864 == array_index_239556 ? add_244024 : sel_244021;
  assign add_244028 = sel_244025 + 8'h01;
  assign sel_244029 = array_index_243864 == array_index_239562 ? add_244028 : sel_244025;
  assign add_244032 = sel_244029 + 8'h01;
  assign sel_244033 = array_index_243864 == array_index_239568 ? add_244032 : sel_244029;
  assign add_244036 = sel_244033 + 8'h01;
  assign sel_244037 = array_index_243864 == array_index_239574 ? add_244036 : sel_244033;
  assign add_244040 = sel_244037 + 8'h01;
  assign sel_244041 = array_index_243864 == array_index_239580 ? add_244040 : sel_244037;
  assign add_244044 = sel_244041 + 8'h01;
  assign sel_244045 = array_index_243864 == array_index_239586 ? add_244044 : sel_244041;
  assign add_244048 = sel_244045 + 8'h01;
  assign sel_244049 = array_index_243864 == array_index_239592 ? add_244048 : sel_244045;
  assign add_244052 = sel_244049 + 8'h01;
  assign sel_244053 = array_index_243864 == array_index_239598 ? add_244052 : sel_244049;
  assign add_244056 = sel_244053 + 8'h01;
  assign sel_244057 = array_index_243864 == array_index_239604 ? add_244056 : sel_244053;
  assign add_244060 = sel_244057 + 8'h01;
  assign sel_244061 = array_index_243864 == array_index_239610 ? add_244060 : sel_244057;
  assign add_244065 = sel_244061 + 8'h01;
  assign array_index_244066 = set1_unflattened[6'h17];
  assign sel_244067 = array_index_243864 == array_index_239616 ? add_244065 : sel_244061;
  assign add_244070 = sel_244067 + 8'h01;
  assign sel_244071 = array_index_244066 == array_index_239312 ? add_244070 : sel_244067;
  assign add_244074 = sel_244071 + 8'h01;
  assign sel_244075 = array_index_244066 == array_index_239316 ? add_244074 : sel_244071;
  assign add_244078 = sel_244075 + 8'h01;
  assign sel_244079 = array_index_244066 == array_index_239324 ? add_244078 : sel_244075;
  assign add_244082 = sel_244079 + 8'h01;
  assign sel_244083 = array_index_244066 == array_index_239332 ? add_244082 : sel_244079;
  assign add_244086 = sel_244083 + 8'h01;
  assign sel_244087 = array_index_244066 == array_index_239340 ? add_244086 : sel_244083;
  assign add_244090 = sel_244087 + 8'h01;
  assign sel_244091 = array_index_244066 == array_index_239348 ? add_244090 : sel_244087;
  assign add_244094 = sel_244091 + 8'h01;
  assign sel_244095 = array_index_244066 == array_index_239356 ? add_244094 : sel_244091;
  assign add_244098 = sel_244095 + 8'h01;
  assign sel_244099 = array_index_244066 == array_index_239364 ? add_244098 : sel_244095;
  assign add_244102 = sel_244099 + 8'h01;
  assign sel_244103 = array_index_244066 == array_index_239370 ? add_244102 : sel_244099;
  assign add_244106 = sel_244103 + 8'h01;
  assign sel_244107 = array_index_244066 == array_index_239376 ? add_244106 : sel_244103;
  assign add_244110 = sel_244107 + 8'h01;
  assign sel_244111 = array_index_244066 == array_index_239382 ? add_244110 : sel_244107;
  assign add_244114 = sel_244111 + 8'h01;
  assign sel_244115 = array_index_244066 == array_index_239388 ? add_244114 : sel_244111;
  assign add_244118 = sel_244115 + 8'h01;
  assign sel_244119 = array_index_244066 == array_index_239394 ? add_244118 : sel_244115;
  assign add_244122 = sel_244119 + 8'h01;
  assign sel_244123 = array_index_244066 == array_index_239400 ? add_244122 : sel_244119;
  assign add_244126 = sel_244123 + 8'h01;
  assign sel_244127 = array_index_244066 == array_index_239406 ? add_244126 : sel_244123;
  assign add_244130 = sel_244127 + 8'h01;
  assign sel_244131 = array_index_244066 == array_index_239412 ? add_244130 : sel_244127;
  assign add_244134 = sel_244131 + 8'h01;
  assign sel_244135 = array_index_244066 == array_index_239418 ? add_244134 : sel_244131;
  assign add_244138 = sel_244135 + 8'h01;
  assign sel_244139 = array_index_244066 == array_index_239424 ? add_244138 : sel_244135;
  assign add_244142 = sel_244139 + 8'h01;
  assign sel_244143 = array_index_244066 == array_index_239430 ? add_244142 : sel_244139;
  assign add_244146 = sel_244143 + 8'h01;
  assign sel_244147 = array_index_244066 == array_index_239436 ? add_244146 : sel_244143;
  assign add_244150 = sel_244147 + 8'h01;
  assign sel_244151 = array_index_244066 == array_index_239442 ? add_244150 : sel_244147;
  assign add_244154 = sel_244151 + 8'h01;
  assign sel_244155 = array_index_244066 == array_index_239448 ? add_244154 : sel_244151;
  assign add_244158 = sel_244155 + 8'h01;
  assign sel_244159 = array_index_244066 == array_index_239454 ? add_244158 : sel_244155;
  assign add_244162 = sel_244159 + 8'h01;
  assign sel_244163 = array_index_244066 == array_index_239460 ? add_244162 : sel_244159;
  assign add_244166 = sel_244163 + 8'h01;
  assign sel_244167 = array_index_244066 == array_index_239466 ? add_244166 : sel_244163;
  assign add_244170 = sel_244167 + 8'h01;
  assign sel_244171 = array_index_244066 == array_index_239472 ? add_244170 : sel_244167;
  assign add_244174 = sel_244171 + 8'h01;
  assign sel_244175 = array_index_244066 == array_index_239478 ? add_244174 : sel_244171;
  assign add_244178 = sel_244175 + 8'h01;
  assign sel_244179 = array_index_244066 == array_index_239484 ? add_244178 : sel_244175;
  assign add_244182 = sel_244179 + 8'h01;
  assign sel_244183 = array_index_244066 == array_index_239490 ? add_244182 : sel_244179;
  assign add_244186 = sel_244183 + 8'h01;
  assign sel_244187 = array_index_244066 == array_index_239496 ? add_244186 : sel_244183;
  assign add_244190 = sel_244187 + 8'h01;
  assign sel_244191 = array_index_244066 == array_index_239502 ? add_244190 : sel_244187;
  assign add_244194 = sel_244191 + 8'h01;
  assign sel_244195 = array_index_244066 == array_index_239508 ? add_244194 : sel_244191;
  assign add_244198 = sel_244195 + 8'h01;
  assign sel_244199 = array_index_244066 == array_index_239514 ? add_244198 : sel_244195;
  assign add_244202 = sel_244199 + 8'h01;
  assign sel_244203 = array_index_244066 == array_index_239520 ? add_244202 : sel_244199;
  assign add_244206 = sel_244203 + 8'h01;
  assign sel_244207 = array_index_244066 == array_index_239526 ? add_244206 : sel_244203;
  assign add_244210 = sel_244207 + 8'h01;
  assign sel_244211 = array_index_244066 == array_index_239532 ? add_244210 : sel_244207;
  assign add_244214 = sel_244211 + 8'h01;
  assign sel_244215 = array_index_244066 == array_index_239538 ? add_244214 : sel_244211;
  assign add_244218 = sel_244215 + 8'h01;
  assign sel_244219 = array_index_244066 == array_index_239544 ? add_244218 : sel_244215;
  assign add_244222 = sel_244219 + 8'h01;
  assign sel_244223 = array_index_244066 == array_index_239550 ? add_244222 : sel_244219;
  assign add_244226 = sel_244223 + 8'h01;
  assign sel_244227 = array_index_244066 == array_index_239556 ? add_244226 : sel_244223;
  assign add_244230 = sel_244227 + 8'h01;
  assign sel_244231 = array_index_244066 == array_index_239562 ? add_244230 : sel_244227;
  assign add_244234 = sel_244231 + 8'h01;
  assign sel_244235 = array_index_244066 == array_index_239568 ? add_244234 : sel_244231;
  assign add_244238 = sel_244235 + 8'h01;
  assign sel_244239 = array_index_244066 == array_index_239574 ? add_244238 : sel_244235;
  assign add_244242 = sel_244239 + 8'h01;
  assign sel_244243 = array_index_244066 == array_index_239580 ? add_244242 : sel_244239;
  assign add_244246 = sel_244243 + 8'h01;
  assign sel_244247 = array_index_244066 == array_index_239586 ? add_244246 : sel_244243;
  assign add_244250 = sel_244247 + 8'h01;
  assign sel_244251 = array_index_244066 == array_index_239592 ? add_244250 : sel_244247;
  assign add_244254 = sel_244251 + 8'h01;
  assign sel_244255 = array_index_244066 == array_index_239598 ? add_244254 : sel_244251;
  assign add_244258 = sel_244255 + 8'h01;
  assign sel_244259 = array_index_244066 == array_index_239604 ? add_244258 : sel_244255;
  assign add_244262 = sel_244259 + 8'h01;
  assign sel_244263 = array_index_244066 == array_index_239610 ? add_244262 : sel_244259;
  assign add_244267 = sel_244263 + 8'h01;
  assign array_index_244268 = set1_unflattened[6'h18];
  assign sel_244269 = array_index_244066 == array_index_239616 ? add_244267 : sel_244263;
  assign add_244272 = sel_244269 + 8'h01;
  assign sel_244273 = array_index_244268 == array_index_239312 ? add_244272 : sel_244269;
  assign add_244276 = sel_244273 + 8'h01;
  assign sel_244277 = array_index_244268 == array_index_239316 ? add_244276 : sel_244273;
  assign add_244280 = sel_244277 + 8'h01;
  assign sel_244281 = array_index_244268 == array_index_239324 ? add_244280 : sel_244277;
  assign add_244284 = sel_244281 + 8'h01;
  assign sel_244285 = array_index_244268 == array_index_239332 ? add_244284 : sel_244281;
  assign add_244288 = sel_244285 + 8'h01;
  assign sel_244289 = array_index_244268 == array_index_239340 ? add_244288 : sel_244285;
  assign add_244292 = sel_244289 + 8'h01;
  assign sel_244293 = array_index_244268 == array_index_239348 ? add_244292 : sel_244289;
  assign add_244296 = sel_244293 + 8'h01;
  assign sel_244297 = array_index_244268 == array_index_239356 ? add_244296 : sel_244293;
  assign add_244300 = sel_244297 + 8'h01;
  assign sel_244301 = array_index_244268 == array_index_239364 ? add_244300 : sel_244297;
  assign add_244304 = sel_244301 + 8'h01;
  assign sel_244305 = array_index_244268 == array_index_239370 ? add_244304 : sel_244301;
  assign add_244308 = sel_244305 + 8'h01;
  assign sel_244309 = array_index_244268 == array_index_239376 ? add_244308 : sel_244305;
  assign add_244312 = sel_244309 + 8'h01;
  assign sel_244313 = array_index_244268 == array_index_239382 ? add_244312 : sel_244309;
  assign add_244316 = sel_244313 + 8'h01;
  assign sel_244317 = array_index_244268 == array_index_239388 ? add_244316 : sel_244313;
  assign add_244320 = sel_244317 + 8'h01;
  assign sel_244321 = array_index_244268 == array_index_239394 ? add_244320 : sel_244317;
  assign add_244324 = sel_244321 + 8'h01;
  assign sel_244325 = array_index_244268 == array_index_239400 ? add_244324 : sel_244321;
  assign add_244328 = sel_244325 + 8'h01;
  assign sel_244329 = array_index_244268 == array_index_239406 ? add_244328 : sel_244325;
  assign add_244332 = sel_244329 + 8'h01;
  assign sel_244333 = array_index_244268 == array_index_239412 ? add_244332 : sel_244329;
  assign add_244336 = sel_244333 + 8'h01;
  assign sel_244337 = array_index_244268 == array_index_239418 ? add_244336 : sel_244333;
  assign add_244340 = sel_244337 + 8'h01;
  assign sel_244341 = array_index_244268 == array_index_239424 ? add_244340 : sel_244337;
  assign add_244344 = sel_244341 + 8'h01;
  assign sel_244345 = array_index_244268 == array_index_239430 ? add_244344 : sel_244341;
  assign add_244348 = sel_244345 + 8'h01;
  assign sel_244349 = array_index_244268 == array_index_239436 ? add_244348 : sel_244345;
  assign add_244352 = sel_244349 + 8'h01;
  assign sel_244353 = array_index_244268 == array_index_239442 ? add_244352 : sel_244349;
  assign add_244356 = sel_244353 + 8'h01;
  assign sel_244357 = array_index_244268 == array_index_239448 ? add_244356 : sel_244353;
  assign add_244360 = sel_244357 + 8'h01;
  assign sel_244361 = array_index_244268 == array_index_239454 ? add_244360 : sel_244357;
  assign add_244364 = sel_244361 + 8'h01;
  assign sel_244365 = array_index_244268 == array_index_239460 ? add_244364 : sel_244361;
  assign add_244368 = sel_244365 + 8'h01;
  assign sel_244369 = array_index_244268 == array_index_239466 ? add_244368 : sel_244365;
  assign add_244372 = sel_244369 + 8'h01;
  assign sel_244373 = array_index_244268 == array_index_239472 ? add_244372 : sel_244369;
  assign add_244376 = sel_244373 + 8'h01;
  assign sel_244377 = array_index_244268 == array_index_239478 ? add_244376 : sel_244373;
  assign add_244380 = sel_244377 + 8'h01;
  assign sel_244381 = array_index_244268 == array_index_239484 ? add_244380 : sel_244377;
  assign add_244384 = sel_244381 + 8'h01;
  assign sel_244385 = array_index_244268 == array_index_239490 ? add_244384 : sel_244381;
  assign add_244388 = sel_244385 + 8'h01;
  assign sel_244389 = array_index_244268 == array_index_239496 ? add_244388 : sel_244385;
  assign add_244392 = sel_244389 + 8'h01;
  assign sel_244393 = array_index_244268 == array_index_239502 ? add_244392 : sel_244389;
  assign add_244396 = sel_244393 + 8'h01;
  assign sel_244397 = array_index_244268 == array_index_239508 ? add_244396 : sel_244393;
  assign add_244400 = sel_244397 + 8'h01;
  assign sel_244401 = array_index_244268 == array_index_239514 ? add_244400 : sel_244397;
  assign add_244404 = sel_244401 + 8'h01;
  assign sel_244405 = array_index_244268 == array_index_239520 ? add_244404 : sel_244401;
  assign add_244408 = sel_244405 + 8'h01;
  assign sel_244409 = array_index_244268 == array_index_239526 ? add_244408 : sel_244405;
  assign add_244412 = sel_244409 + 8'h01;
  assign sel_244413 = array_index_244268 == array_index_239532 ? add_244412 : sel_244409;
  assign add_244416 = sel_244413 + 8'h01;
  assign sel_244417 = array_index_244268 == array_index_239538 ? add_244416 : sel_244413;
  assign add_244420 = sel_244417 + 8'h01;
  assign sel_244421 = array_index_244268 == array_index_239544 ? add_244420 : sel_244417;
  assign add_244424 = sel_244421 + 8'h01;
  assign sel_244425 = array_index_244268 == array_index_239550 ? add_244424 : sel_244421;
  assign add_244428 = sel_244425 + 8'h01;
  assign sel_244429 = array_index_244268 == array_index_239556 ? add_244428 : sel_244425;
  assign add_244432 = sel_244429 + 8'h01;
  assign sel_244433 = array_index_244268 == array_index_239562 ? add_244432 : sel_244429;
  assign add_244436 = sel_244433 + 8'h01;
  assign sel_244437 = array_index_244268 == array_index_239568 ? add_244436 : sel_244433;
  assign add_244440 = sel_244437 + 8'h01;
  assign sel_244441 = array_index_244268 == array_index_239574 ? add_244440 : sel_244437;
  assign add_244444 = sel_244441 + 8'h01;
  assign sel_244445 = array_index_244268 == array_index_239580 ? add_244444 : sel_244441;
  assign add_244448 = sel_244445 + 8'h01;
  assign sel_244449 = array_index_244268 == array_index_239586 ? add_244448 : sel_244445;
  assign add_244452 = sel_244449 + 8'h01;
  assign sel_244453 = array_index_244268 == array_index_239592 ? add_244452 : sel_244449;
  assign add_244456 = sel_244453 + 8'h01;
  assign sel_244457 = array_index_244268 == array_index_239598 ? add_244456 : sel_244453;
  assign add_244460 = sel_244457 + 8'h01;
  assign sel_244461 = array_index_244268 == array_index_239604 ? add_244460 : sel_244457;
  assign add_244464 = sel_244461 + 8'h01;
  assign sel_244465 = array_index_244268 == array_index_239610 ? add_244464 : sel_244461;
  assign add_244469 = sel_244465 + 8'h01;
  assign array_index_244470 = set1_unflattened[6'h19];
  assign sel_244471 = array_index_244268 == array_index_239616 ? add_244469 : sel_244465;
  assign add_244474 = sel_244471 + 8'h01;
  assign sel_244475 = array_index_244470 == array_index_239312 ? add_244474 : sel_244471;
  assign add_244478 = sel_244475 + 8'h01;
  assign sel_244479 = array_index_244470 == array_index_239316 ? add_244478 : sel_244475;
  assign add_244482 = sel_244479 + 8'h01;
  assign sel_244483 = array_index_244470 == array_index_239324 ? add_244482 : sel_244479;
  assign add_244486 = sel_244483 + 8'h01;
  assign sel_244487 = array_index_244470 == array_index_239332 ? add_244486 : sel_244483;
  assign add_244490 = sel_244487 + 8'h01;
  assign sel_244491 = array_index_244470 == array_index_239340 ? add_244490 : sel_244487;
  assign add_244494 = sel_244491 + 8'h01;
  assign sel_244495 = array_index_244470 == array_index_239348 ? add_244494 : sel_244491;
  assign add_244498 = sel_244495 + 8'h01;
  assign sel_244499 = array_index_244470 == array_index_239356 ? add_244498 : sel_244495;
  assign add_244502 = sel_244499 + 8'h01;
  assign sel_244503 = array_index_244470 == array_index_239364 ? add_244502 : sel_244499;
  assign add_244506 = sel_244503 + 8'h01;
  assign sel_244507 = array_index_244470 == array_index_239370 ? add_244506 : sel_244503;
  assign add_244510 = sel_244507 + 8'h01;
  assign sel_244511 = array_index_244470 == array_index_239376 ? add_244510 : sel_244507;
  assign add_244514 = sel_244511 + 8'h01;
  assign sel_244515 = array_index_244470 == array_index_239382 ? add_244514 : sel_244511;
  assign add_244518 = sel_244515 + 8'h01;
  assign sel_244519 = array_index_244470 == array_index_239388 ? add_244518 : sel_244515;
  assign add_244522 = sel_244519 + 8'h01;
  assign sel_244523 = array_index_244470 == array_index_239394 ? add_244522 : sel_244519;
  assign add_244526 = sel_244523 + 8'h01;
  assign sel_244527 = array_index_244470 == array_index_239400 ? add_244526 : sel_244523;
  assign add_244530 = sel_244527 + 8'h01;
  assign sel_244531 = array_index_244470 == array_index_239406 ? add_244530 : sel_244527;
  assign add_244534 = sel_244531 + 8'h01;
  assign sel_244535 = array_index_244470 == array_index_239412 ? add_244534 : sel_244531;
  assign add_244538 = sel_244535 + 8'h01;
  assign sel_244539 = array_index_244470 == array_index_239418 ? add_244538 : sel_244535;
  assign add_244542 = sel_244539 + 8'h01;
  assign sel_244543 = array_index_244470 == array_index_239424 ? add_244542 : sel_244539;
  assign add_244546 = sel_244543 + 8'h01;
  assign sel_244547 = array_index_244470 == array_index_239430 ? add_244546 : sel_244543;
  assign add_244550 = sel_244547 + 8'h01;
  assign sel_244551 = array_index_244470 == array_index_239436 ? add_244550 : sel_244547;
  assign add_244554 = sel_244551 + 8'h01;
  assign sel_244555 = array_index_244470 == array_index_239442 ? add_244554 : sel_244551;
  assign add_244558 = sel_244555 + 8'h01;
  assign sel_244559 = array_index_244470 == array_index_239448 ? add_244558 : sel_244555;
  assign add_244562 = sel_244559 + 8'h01;
  assign sel_244563 = array_index_244470 == array_index_239454 ? add_244562 : sel_244559;
  assign add_244566 = sel_244563 + 8'h01;
  assign sel_244567 = array_index_244470 == array_index_239460 ? add_244566 : sel_244563;
  assign add_244570 = sel_244567 + 8'h01;
  assign sel_244571 = array_index_244470 == array_index_239466 ? add_244570 : sel_244567;
  assign add_244574 = sel_244571 + 8'h01;
  assign sel_244575 = array_index_244470 == array_index_239472 ? add_244574 : sel_244571;
  assign add_244578 = sel_244575 + 8'h01;
  assign sel_244579 = array_index_244470 == array_index_239478 ? add_244578 : sel_244575;
  assign add_244582 = sel_244579 + 8'h01;
  assign sel_244583 = array_index_244470 == array_index_239484 ? add_244582 : sel_244579;
  assign add_244586 = sel_244583 + 8'h01;
  assign sel_244587 = array_index_244470 == array_index_239490 ? add_244586 : sel_244583;
  assign add_244590 = sel_244587 + 8'h01;
  assign sel_244591 = array_index_244470 == array_index_239496 ? add_244590 : sel_244587;
  assign add_244594 = sel_244591 + 8'h01;
  assign sel_244595 = array_index_244470 == array_index_239502 ? add_244594 : sel_244591;
  assign add_244598 = sel_244595 + 8'h01;
  assign sel_244599 = array_index_244470 == array_index_239508 ? add_244598 : sel_244595;
  assign add_244602 = sel_244599 + 8'h01;
  assign sel_244603 = array_index_244470 == array_index_239514 ? add_244602 : sel_244599;
  assign add_244606 = sel_244603 + 8'h01;
  assign sel_244607 = array_index_244470 == array_index_239520 ? add_244606 : sel_244603;
  assign add_244610 = sel_244607 + 8'h01;
  assign sel_244611 = array_index_244470 == array_index_239526 ? add_244610 : sel_244607;
  assign add_244614 = sel_244611 + 8'h01;
  assign sel_244615 = array_index_244470 == array_index_239532 ? add_244614 : sel_244611;
  assign add_244618 = sel_244615 + 8'h01;
  assign sel_244619 = array_index_244470 == array_index_239538 ? add_244618 : sel_244615;
  assign add_244622 = sel_244619 + 8'h01;
  assign sel_244623 = array_index_244470 == array_index_239544 ? add_244622 : sel_244619;
  assign add_244626 = sel_244623 + 8'h01;
  assign sel_244627 = array_index_244470 == array_index_239550 ? add_244626 : sel_244623;
  assign add_244630 = sel_244627 + 8'h01;
  assign sel_244631 = array_index_244470 == array_index_239556 ? add_244630 : sel_244627;
  assign add_244634 = sel_244631 + 8'h01;
  assign sel_244635 = array_index_244470 == array_index_239562 ? add_244634 : sel_244631;
  assign add_244638 = sel_244635 + 8'h01;
  assign sel_244639 = array_index_244470 == array_index_239568 ? add_244638 : sel_244635;
  assign add_244642 = sel_244639 + 8'h01;
  assign sel_244643 = array_index_244470 == array_index_239574 ? add_244642 : sel_244639;
  assign add_244646 = sel_244643 + 8'h01;
  assign sel_244647 = array_index_244470 == array_index_239580 ? add_244646 : sel_244643;
  assign add_244650 = sel_244647 + 8'h01;
  assign sel_244651 = array_index_244470 == array_index_239586 ? add_244650 : sel_244647;
  assign add_244654 = sel_244651 + 8'h01;
  assign sel_244655 = array_index_244470 == array_index_239592 ? add_244654 : sel_244651;
  assign add_244658 = sel_244655 + 8'h01;
  assign sel_244659 = array_index_244470 == array_index_239598 ? add_244658 : sel_244655;
  assign add_244662 = sel_244659 + 8'h01;
  assign sel_244663 = array_index_244470 == array_index_239604 ? add_244662 : sel_244659;
  assign add_244666 = sel_244663 + 8'h01;
  assign sel_244667 = array_index_244470 == array_index_239610 ? add_244666 : sel_244663;
  assign add_244671 = sel_244667 + 8'h01;
  assign array_index_244672 = set1_unflattened[6'h1a];
  assign sel_244673 = array_index_244470 == array_index_239616 ? add_244671 : sel_244667;
  assign add_244676 = sel_244673 + 8'h01;
  assign sel_244677 = array_index_244672 == array_index_239312 ? add_244676 : sel_244673;
  assign add_244680 = sel_244677 + 8'h01;
  assign sel_244681 = array_index_244672 == array_index_239316 ? add_244680 : sel_244677;
  assign add_244684 = sel_244681 + 8'h01;
  assign sel_244685 = array_index_244672 == array_index_239324 ? add_244684 : sel_244681;
  assign add_244688 = sel_244685 + 8'h01;
  assign sel_244689 = array_index_244672 == array_index_239332 ? add_244688 : sel_244685;
  assign add_244692 = sel_244689 + 8'h01;
  assign sel_244693 = array_index_244672 == array_index_239340 ? add_244692 : sel_244689;
  assign add_244696 = sel_244693 + 8'h01;
  assign sel_244697 = array_index_244672 == array_index_239348 ? add_244696 : sel_244693;
  assign add_244700 = sel_244697 + 8'h01;
  assign sel_244701 = array_index_244672 == array_index_239356 ? add_244700 : sel_244697;
  assign add_244704 = sel_244701 + 8'h01;
  assign sel_244705 = array_index_244672 == array_index_239364 ? add_244704 : sel_244701;
  assign add_244708 = sel_244705 + 8'h01;
  assign sel_244709 = array_index_244672 == array_index_239370 ? add_244708 : sel_244705;
  assign add_244712 = sel_244709 + 8'h01;
  assign sel_244713 = array_index_244672 == array_index_239376 ? add_244712 : sel_244709;
  assign add_244716 = sel_244713 + 8'h01;
  assign sel_244717 = array_index_244672 == array_index_239382 ? add_244716 : sel_244713;
  assign add_244720 = sel_244717 + 8'h01;
  assign sel_244721 = array_index_244672 == array_index_239388 ? add_244720 : sel_244717;
  assign add_244724 = sel_244721 + 8'h01;
  assign sel_244725 = array_index_244672 == array_index_239394 ? add_244724 : sel_244721;
  assign add_244728 = sel_244725 + 8'h01;
  assign sel_244729 = array_index_244672 == array_index_239400 ? add_244728 : sel_244725;
  assign add_244732 = sel_244729 + 8'h01;
  assign sel_244733 = array_index_244672 == array_index_239406 ? add_244732 : sel_244729;
  assign add_244736 = sel_244733 + 8'h01;
  assign sel_244737 = array_index_244672 == array_index_239412 ? add_244736 : sel_244733;
  assign add_244740 = sel_244737 + 8'h01;
  assign sel_244741 = array_index_244672 == array_index_239418 ? add_244740 : sel_244737;
  assign add_244744 = sel_244741 + 8'h01;
  assign sel_244745 = array_index_244672 == array_index_239424 ? add_244744 : sel_244741;
  assign add_244748 = sel_244745 + 8'h01;
  assign sel_244749 = array_index_244672 == array_index_239430 ? add_244748 : sel_244745;
  assign add_244752 = sel_244749 + 8'h01;
  assign sel_244753 = array_index_244672 == array_index_239436 ? add_244752 : sel_244749;
  assign add_244756 = sel_244753 + 8'h01;
  assign sel_244757 = array_index_244672 == array_index_239442 ? add_244756 : sel_244753;
  assign add_244760 = sel_244757 + 8'h01;
  assign sel_244761 = array_index_244672 == array_index_239448 ? add_244760 : sel_244757;
  assign add_244764 = sel_244761 + 8'h01;
  assign sel_244765 = array_index_244672 == array_index_239454 ? add_244764 : sel_244761;
  assign add_244768 = sel_244765 + 8'h01;
  assign sel_244769 = array_index_244672 == array_index_239460 ? add_244768 : sel_244765;
  assign add_244772 = sel_244769 + 8'h01;
  assign sel_244773 = array_index_244672 == array_index_239466 ? add_244772 : sel_244769;
  assign add_244776 = sel_244773 + 8'h01;
  assign sel_244777 = array_index_244672 == array_index_239472 ? add_244776 : sel_244773;
  assign add_244780 = sel_244777 + 8'h01;
  assign sel_244781 = array_index_244672 == array_index_239478 ? add_244780 : sel_244777;
  assign add_244784 = sel_244781 + 8'h01;
  assign sel_244785 = array_index_244672 == array_index_239484 ? add_244784 : sel_244781;
  assign add_244788 = sel_244785 + 8'h01;
  assign sel_244789 = array_index_244672 == array_index_239490 ? add_244788 : sel_244785;
  assign add_244792 = sel_244789 + 8'h01;
  assign sel_244793 = array_index_244672 == array_index_239496 ? add_244792 : sel_244789;
  assign add_244796 = sel_244793 + 8'h01;
  assign sel_244797 = array_index_244672 == array_index_239502 ? add_244796 : sel_244793;
  assign add_244800 = sel_244797 + 8'h01;
  assign sel_244801 = array_index_244672 == array_index_239508 ? add_244800 : sel_244797;
  assign add_244804 = sel_244801 + 8'h01;
  assign sel_244805 = array_index_244672 == array_index_239514 ? add_244804 : sel_244801;
  assign add_244808 = sel_244805 + 8'h01;
  assign sel_244809 = array_index_244672 == array_index_239520 ? add_244808 : sel_244805;
  assign add_244812 = sel_244809 + 8'h01;
  assign sel_244813 = array_index_244672 == array_index_239526 ? add_244812 : sel_244809;
  assign add_244816 = sel_244813 + 8'h01;
  assign sel_244817 = array_index_244672 == array_index_239532 ? add_244816 : sel_244813;
  assign add_244820 = sel_244817 + 8'h01;
  assign sel_244821 = array_index_244672 == array_index_239538 ? add_244820 : sel_244817;
  assign add_244824 = sel_244821 + 8'h01;
  assign sel_244825 = array_index_244672 == array_index_239544 ? add_244824 : sel_244821;
  assign add_244828 = sel_244825 + 8'h01;
  assign sel_244829 = array_index_244672 == array_index_239550 ? add_244828 : sel_244825;
  assign add_244832 = sel_244829 + 8'h01;
  assign sel_244833 = array_index_244672 == array_index_239556 ? add_244832 : sel_244829;
  assign add_244836 = sel_244833 + 8'h01;
  assign sel_244837 = array_index_244672 == array_index_239562 ? add_244836 : sel_244833;
  assign add_244840 = sel_244837 + 8'h01;
  assign sel_244841 = array_index_244672 == array_index_239568 ? add_244840 : sel_244837;
  assign add_244844 = sel_244841 + 8'h01;
  assign sel_244845 = array_index_244672 == array_index_239574 ? add_244844 : sel_244841;
  assign add_244848 = sel_244845 + 8'h01;
  assign sel_244849 = array_index_244672 == array_index_239580 ? add_244848 : sel_244845;
  assign add_244852 = sel_244849 + 8'h01;
  assign sel_244853 = array_index_244672 == array_index_239586 ? add_244852 : sel_244849;
  assign add_244856 = sel_244853 + 8'h01;
  assign sel_244857 = array_index_244672 == array_index_239592 ? add_244856 : sel_244853;
  assign add_244860 = sel_244857 + 8'h01;
  assign sel_244861 = array_index_244672 == array_index_239598 ? add_244860 : sel_244857;
  assign add_244864 = sel_244861 + 8'h01;
  assign sel_244865 = array_index_244672 == array_index_239604 ? add_244864 : sel_244861;
  assign add_244868 = sel_244865 + 8'h01;
  assign sel_244869 = array_index_244672 == array_index_239610 ? add_244868 : sel_244865;
  assign add_244873 = sel_244869 + 8'h01;
  assign array_index_244874 = set1_unflattened[6'h1b];
  assign sel_244875 = array_index_244672 == array_index_239616 ? add_244873 : sel_244869;
  assign add_244878 = sel_244875 + 8'h01;
  assign sel_244879 = array_index_244874 == array_index_239312 ? add_244878 : sel_244875;
  assign add_244882 = sel_244879 + 8'h01;
  assign sel_244883 = array_index_244874 == array_index_239316 ? add_244882 : sel_244879;
  assign add_244886 = sel_244883 + 8'h01;
  assign sel_244887 = array_index_244874 == array_index_239324 ? add_244886 : sel_244883;
  assign add_244890 = sel_244887 + 8'h01;
  assign sel_244891 = array_index_244874 == array_index_239332 ? add_244890 : sel_244887;
  assign add_244894 = sel_244891 + 8'h01;
  assign sel_244895 = array_index_244874 == array_index_239340 ? add_244894 : sel_244891;
  assign add_244898 = sel_244895 + 8'h01;
  assign sel_244899 = array_index_244874 == array_index_239348 ? add_244898 : sel_244895;
  assign add_244902 = sel_244899 + 8'h01;
  assign sel_244903 = array_index_244874 == array_index_239356 ? add_244902 : sel_244899;
  assign add_244906 = sel_244903 + 8'h01;
  assign sel_244907 = array_index_244874 == array_index_239364 ? add_244906 : sel_244903;
  assign add_244910 = sel_244907 + 8'h01;
  assign sel_244911 = array_index_244874 == array_index_239370 ? add_244910 : sel_244907;
  assign add_244914 = sel_244911 + 8'h01;
  assign sel_244915 = array_index_244874 == array_index_239376 ? add_244914 : sel_244911;
  assign add_244918 = sel_244915 + 8'h01;
  assign sel_244919 = array_index_244874 == array_index_239382 ? add_244918 : sel_244915;
  assign add_244922 = sel_244919 + 8'h01;
  assign sel_244923 = array_index_244874 == array_index_239388 ? add_244922 : sel_244919;
  assign add_244926 = sel_244923 + 8'h01;
  assign sel_244927 = array_index_244874 == array_index_239394 ? add_244926 : sel_244923;
  assign add_244930 = sel_244927 + 8'h01;
  assign sel_244931 = array_index_244874 == array_index_239400 ? add_244930 : sel_244927;
  assign add_244934 = sel_244931 + 8'h01;
  assign sel_244935 = array_index_244874 == array_index_239406 ? add_244934 : sel_244931;
  assign add_244938 = sel_244935 + 8'h01;
  assign sel_244939 = array_index_244874 == array_index_239412 ? add_244938 : sel_244935;
  assign add_244942 = sel_244939 + 8'h01;
  assign sel_244943 = array_index_244874 == array_index_239418 ? add_244942 : sel_244939;
  assign add_244946 = sel_244943 + 8'h01;
  assign sel_244947 = array_index_244874 == array_index_239424 ? add_244946 : sel_244943;
  assign add_244950 = sel_244947 + 8'h01;
  assign sel_244951 = array_index_244874 == array_index_239430 ? add_244950 : sel_244947;
  assign add_244954 = sel_244951 + 8'h01;
  assign sel_244955 = array_index_244874 == array_index_239436 ? add_244954 : sel_244951;
  assign add_244958 = sel_244955 + 8'h01;
  assign sel_244959 = array_index_244874 == array_index_239442 ? add_244958 : sel_244955;
  assign add_244962 = sel_244959 + 8'h01;
  assign sel_244963 = array_index_244874 == array_index_239448 ? add_244962 : sel_244959;
  assign add_244966 = sel_244963 + 8'h01;
  assign sel_244967 = array_index_244874 == array_index_239454 ? add_244966 : sel_244963;
  assign add_244970 = sel_244967 + 8'h01;
  assign sel_244971 = array_index_244874 == array_index_239460 ? add_244970 : sel_244967;
  assign add_244974 = sel_244971 + 8'h01;
  assign sel_244975 = array_index_244874 == array_index_239466 ? add_244974 : sel_244971;
  assign add_244978 = sel_244975 + 8'h01;
  assign sel_244979 = array_index_244874 == array_index_239472 ? add_244978 : sel_244975;
  assign add_244982 = sel_244979 + 8'h01;
  assign sel_244983 = array_index_244874 == array_index_239478 ? add_244982 : sel_244979;
  assign add_244986 = sel_244983 + 8'h01;
  assign sel_244987 = array_index_244874 == array_index_239484 ? add_244986 : sel_244983;
  assign add_244990 = sel_244987 + 8'h01;
  assign sel_244991 = array_index_244874 == array_index_239490 ? add_244990 : sel_244987;
  assign add_244994 = sel_244991 + 8'h01;
  assign sel_244995 = array_index_244874 == array_index_239496 ? add_244994 : sel_244991;
  assign add_244998 = sel_244995 + 8'h01;
  assign sel_244999 = array_index_244874 == array_index_239502 ? add_244998 : sel_244995;
  assign add_245002 = sel_244999 + 8'h01;
  assign sel_245003 = array_index_244874 == array_index_239508 ? add_245002 : sel_244999;
  assign add_245006 = sel_245003 + 8'h01;
  assign sel_245007 = array_index_244874 == array_index_239514 ? add_245006 : sel_245003;
  assign add_245010 = sel_245007 + 8'h01;
  assign sel_245011 = array_index_244874 == array_index_239520 ? add_245010 : sel_245007;
  assign add_245014 = sel_245011 + 8'h01;
  assign sel_245015 = array_index_244874 == array_index_239526 ? add_245014 : sel_245011;
  assign add_245018 = sel_245015 + 8'h01;
  assign sel_245019 = array_index_244874 == array_index_239532 ? add_245018 : sel_245015;
  assign add_245022 = sel_245019 + 8'h01;
  assign sel_245023 = array_index_244874 == array_index_239538 ? add_245022 : sel_245019;
  assign add_245026 = sel_245023 + 8'h01;
  assign sel_245027 = array_index_244874 == array_index_239544 ? add_245026 : sel_245023;
  assign add_245030 = sel_245027 + 8'h01;
  assign sel_245031 = array_index_244874 == array_index_239550 ? add_245030 : sel_245027;
  assign add_245034 = sel_245031 + 8'h01;
  assign sel_245035 = array_index_244874 == array_index_239556 ? add_245034 : sel_245031;
  assign add_245038 = sel_245035 + 8'h01;
  assign sel_245039 = array_index_244874 == array_index_239562 ? add_245038 : sel_245035;
  assign add_245042 = sel_245039 + 8'h01;
  assign sel_245043 = array_index_244874 == array_index_239568 ? add_245042 : sel_245039;
  assign add_245046 = sel_245043 + 8'h01;
  assign sel_245047 = array_index_244874 == array_index_239574 ? add_245046 : sel_245043;
  assign add_245050 = sel_245047 + 8'h01;
  assign sel_245051 = array_index_244874 == array_index_239580 ? add_245050 : sel_245047;
  assign add_245054 = sel_245051 + 8'h01;
  assign sel_245055 = array_index_244874 == array_index_239586 ? add_245054 : sel_245051;
  assign add_245058 = sel_245055 + 8'h01;
  assign sel_245059 = array_index_244874 == array_index_239592 ? add_245058 : sel_245055;
  assign add_245062 = sel_245059 + 8'h01;
  assign sel_245063 = array_index_244874 == array_index_239598 ? add_245062 : sel_245059;
  assign add_245066 = sel_245063 + 8'h01;
  assign sel_245067 = array_index_244874 == array_index_239604 ? add_245066 : sel_245063;
  assign add_245070 = sel_245067 + 8'h01;
  assign sel_245071 = array_index_244874 == array_index_239610 ? add_245070 : sel_245067;
  assign add_245075 = sel_245071 + 8'h01;
  assign array_index_245076 = set1_unflattened[6'h1c];
  assign sel_245077 = array_index_244874 == array_index_239616 ? add_245075 : sel_245071;
  assign add_245080 = sel_245077 + 8'h01;
  assign sel_245081 = array_index_245076 == array_index_239312 ? add_245080 : sel_245077;
  assign add_245084 = sel_245081 + 8'h01;
  assign sel_245085 = array_index_245076 == array_index_239316 ? add_245084 : sel_245081;
  assign add_245088 = sel_245085 + 8'h01;
  assign sel_245089 = array_index_245076 == array_index_239324 ? add_245088 : sel_245085;
  assign add_245092 = sel_245089 + 8'h01;
  assign sel_245093 = array_index_245076 == array_index_239332 ? add_245092 : sel_245089;
  assign add_245096 = sel_245093 + 8'h01;
  assign sel_245097 = array_index_245076 == array_index_239340 ? add_245096 : sel_245093;
  assign add_245100 = sel_245097 + 8'h01;
  assign sel_245101 = array_index_245076 == array_index_239348 ? add_245100 : sel_245097;
  assign add_245104 = sel_245101 + 8'h01;
  assign sel_245105 = array_index_245076 == array_index_239356 ? add_245104 : sel_245101;
  assign add_245108 = sel_245105 + 8'h01;
  assign sel_245109 = array_index_245076 == array_index_239364 ? add_245108 : sel_245105;
  assign add_245112 = sel_245109 + 8'h01;
  assign sel_245113 = array_index_245076 == array_index_239370 ? add_245112 : sel_245109;
  assign add_245116 = sel_245113 + 8'h01;
  assign sel_245117 = array_index_245076 == array_index_239376 ? add_245116 : sel_245113;
  assign add_245120 = sel_245117 + 8'h01;
  assign sel_245121 = array_index_245076 == array_index_239382 ? add_245120 : sel_245117;
  assign add_245124 = sel_245121 + 8'h01;
  assign sel_245125 = array_index_245076 == array_index_239388 ? add_245124 : sel_245121;
  assign add_245128 = sel_245125 + 8'h01;
  assign sel_245129 = array_index_245076 == array_index_239394 ? add_245128 : sel_245125;
  assign add_245132 = sel_245129 + 8'h01;
  assign sel_245133 = array_index_245076 == array_index_239400 ? add_245132 : sel_245129;
  assign add_245136 = sel_245133 + 8'h01;
  assign sel_245137 = array_index_245076 == array_index_239406 ? add_245136 : sel_245133;
  assign add_245140 = sel_245137 + 8'h01;
  assign sel_245141 = array_index_245076 == array_index_239412 ? add_245140 : sel_245137;
  assign add_245144 = sel_245141 + 8'h01;
  assign sel_245145 = array_index_245076 == array_index_239418 ? add_245144 : sel_245141;
  assign add_245148 = sel_245145 + 8'h01;
  assign sel_245149 = array_index_245076 == array_index_239424 ? add_245148 : sel_245145;
  assign add_245152 = sel_245149 + 8'h01;
  assign sel_245153 = array_index_245076 == array_index_239430 ? add_245152 : sel_245149;
  assign add_245156 = sel_245153 + 8'h01;
  assign sel_245157 = array_index_245076 == array_index_239436 ? add_245156 : sel_245153;
  assign add_245160 = sel_245157 + 8'h01;
  assign sel_245161 = array_index_245076 == array_index_239442 ? add_245160 : sel_245157;
  assign add_245164 = sel_245161 + 8'h01;
  assign sel_245165 = array_index_245076 == array_index_239448 ? add_245164 : sel_245161;
  assign add_245168 = sel_245165 + 8'h01;
  assign sel_245169 = array_index_245076 == array_index_239454 ? add_245168 : sel_245165;
  assign add_245172 = sel_245169 + 8'h01;
  assign sel_245173 = array_index_245076 == array_index_239460 ? add_245172 : sel_245169;
  assign add_245176 = sel_245173 + 8'h01;
  assign sel_245177 = array_index_245076 == array_index_239466 ? add_245176 : sel_245173;
  assign add_245180 = sel_245177 + 8'h01;
  assign sel_245181 = array_index_245076 == array_index_239472 ? add_245180 : sel_245177;
  assign add_245184 = sel_245181 + 8'h01;
  assign sel_245185 = array_index_245076 == array_index_239478 ? add_245184 : sel_245181;
  assign add_245188 = sel_245185 + 8'h01;
  assign sel_245189 = array_index_245076 == array_index_239484 ? add_245188 : sel_245185;
  assign add_245192 = sel_245189 + 8'h01;
  assign sel_245193 = array_index_245076 == array_index_239490 ? add_245192 : sel_245189;
  assign add_245196 = sel_245193 + 8'h01;
  assign sel_245197 = array_index_245076 == array_index_239496 ? add_245196 : sel_245193;
  assign add_245200 = sel_245197 + 8'h01;
  assign sel_245201 = array_index_245076 == array_index_239502 ? add_245200 : sel_245197;
  assign add_245204 = sel_245201 + 8'h01;
  assign sel_245205 = array_index_245076 == array_index_239508 ? add_245204 : sel_245201;
  assign add_245208 = sel_245205 + 8'h01;
  assign sel_245209 = array_index_245076 == array_index_239514 ? add_245208 : sel_245205;
  assign add_245212 = sel_245209 + 8'h01;
  assign sel_245213 = array_index_245076 == array_index_239520 ? add_245212 : sel_245209;
  assign add_245216 = sel_245213 + 8'h01;
  assign sel_245217 = array_index_245076 == array_index_239526 ? add_245216 : sel_245213;
  assign add_245220 = sel_245217 + 8'h01;
  assign sel_245221 = array_index_245076 == array_index_239532 ? add_245220 : sel_245217;
  assign add_245224 = sel_245221 + 8'h01;
  assign sel_245225 = array_index_245076 == array_index_239538 ? add_245224 : sel_245221;
  assign add_245228 = sel_245225 + 8'h01;
  assign sel_245229 = array_index_245076 == array_index_239544 ? add_245228 : sel_245225;
  assign add_245232 = sel_245229 + 8'h01;
  assign sel_245233 = array_index_245076 == array_index_239550 ? add_245232 : sel_245229;
  assign add_245236 = sel_245233 + 8'h01;
  assign sel_245237 = array_index_245076 == array_index_239556 ? add_245236 : sel_245233;
  assign add_245240 = sel_245237 + 8'h01;
  assign sel_245241 = array_index_245076 == array_index_239562 ? add_245240 : sel_245237;
  assign add_245244 = sel_245241 + 8'h01;
  assign sel_245245 = array_index_245076 == array_index_239568 ? add_245244 : sel_245241;
  assign add_245248 = sel_245245 + 8'h01;
  assign sel_245249 = array_index_245076 == array_index_239574 ? add_245248 : sel_245245;
  assign add_245252 = sel_245249 + 8'h01;
  assign sel_245253 = array_index_245076 == array_index_239580 ? add_245252 : sel_245249;
  assign add_245256 = sel_245253 + 8'h01;
  assign sel_245257 = array_index_245076 == array_index_239586 ? add_245256 : sel_245253;
  assign add_245260 = sel_245257 + 8'h01;
  assign sel_245261 = array_index_245076 == array_index_239592 ? add_245260 : sel_245257;
  assign add_245264 = sel_245261 + 8'h01;
  assign sel_245265 = array_index_245076 == array_index_239598 ? add_245264 : sel_245261;
  assign add_245268 = sel_245265 + 8'h01;
  assign sel_245269 = array_index_245076 == array_index_239604 ? add_245268 : sel_245265;
  assign add_245272 = sel_245269 + 8'h01;
  assign sel_245273 = array_index_245076 == array_index_239610 ? add_245272 : sel_245269;
  assign add_245277 = sel_245273 + 8'h01;
  assign array_index_245278 = set1_unflattened[6'h1d];
  assign sel_245279 = array_index_245076 == array_index_239616 ? add_245277 : sel_245273;
  assign add_245282 = sel_245279 + 8'h01;
  assign sel_245283 = array_index_245278 == array_index_239312 ? add_245282 : sel_245279;
  assign add_245286 = sel_245283 + 8'h01;
  assign sel_245287 = array_index_245278 == array_index_239316 ? add_245286 : sel_245283;
  assign add_245290 = sel_245287 + 8'h01;
  assign sel_245291 = array_index_245278 == array_index_239324 ? add_245290 : sel_245287;
  assign add_245294 = sel_245291 + 8'h01;
  assign sel_245295 = array_index_245278 == array_index_239332 ? add_245294 : sel_245291;
  assign add_245298 = sel_245295 + 8'h01;
  assign sel_245299 = array_index_245278 == array_index_239340 ? add_245298 : sel_245295;
  assign add_245302 = sel_245299 + 8'h01;
  assign sel_245303 = array_index_245278 == array_index_239348 ? add_245302 : sel_245299;
  assign add_245306 = sel_245303 + 8'h01;
  assign sel_245307 = array_index_245278 == array_index_239356 ? add_245306 : sel_245303;
  assign add_245310 = sel_245307 + 8'h01;
  assign sel_245311 = array_index_245278 == array_index_239364 ? add_245310 : sel_245307;
  assign add_245314 = sel_245311 + 8'h01;
  assign sel_245315 = array_index_245278 == array_index_239370 ? add_245314 : sel_245311;
  assign add_245318 = sel_245315 + 8'h01;
  assign sel_245319 = array_index_245278 == array_index_239376 ? add_245318 : sel_245315;
  assign add_245322 = sel_245319 + 8'h01;
  assign sel_245323 = array_index_245278 == array_index_239382 ? add_245322 : sel_245319;
  assign add_245326 = sel_245323 + 8'h01;
  assign sel_245327 = array_index_245278 == array_index_239388 ? add_245326 : sel_245323;
  assign add_245330 = sel_245327 + 8'h01;
  assign sel_245331 = array_index_245278 == array_index_239394 ? add_245330 : sel_245327;
  assign add_245334 = sel_245331 + 8'h01;
  assign sel_245335 = array_index_245278 == array_index_239400 ? add_245334 : sel_245331;
  assign add_245338 = sel_245335 + 8'h01;
  assign sel_245339 = array_index_245278 == array_index_239406 ? add_245338 : sel_245335;
  assign add_245342 = sel_245339 + 8'h01;
  assign sel_245343 = array_index_245278 == array_index_239412 ? add_245342 : sel_245339;
  assign add_245346 = sel_245343 + 8'h01;
  assign sel_245347 = array_index_245278 == array_index_239418 ? add_245346 : sel_245343;
  assign add_245350 = sel_245347 + 8'h01;
  assign sel_245351 = array_index_245278 == array_index_239424 ? add_245350 : sel_245347;
  assign add_245354 = sel_245351 + 8'h01;
  assign sel_245355 = array_index_245278 == array_index_239430 ? add_245354 : sel_245351;
  assign add_245358 = sel_245355 + 8'h01;
  assign sel_245359 = array_index_245278 == array_index_239436 ? add_245358 : sel_245355;
  assign add_245362 = sel_245359 + 8'h01;
  assign sel_245363 = array_index_245278 == array_index_239442 ? add_245362 : sel_245359;
  assign add_245366 = sel_245363 + 8'h01;
  assign sel_245367 = array_index_245278 == array_index_239448 ? add_245366 : sel_245363;
  assign add_245370 = sel_245367 + 8'h01;
  assign sel_245371 = array_index_245278 == array_index_239454 ? add_245370 : sel_245367;
  assign add_245374 = sel_245371 + 8'h01;
  assign sel_245375 = array_index_245278 == array_index_239460 ? add_245374 : sel_245371;
  assign add_245378 = sel_245375 + 8'h01;
  assign sel_245379 = array_index_245278 == array_index_239466 ? add_245378 : sel_245375;
  assign add_245382 = sel_245379 + 8'h01;
  assign sel_245383 = array_index_245278 == array_index_239472 ? add_245382 : sel_245379;
  assign add_245386 = sel_245383 + 8'h01;
  assign sel_245387 = array_index_245278 == array_index_239478 ? add_245386 : sel_245383;
  assign add_245390 = sel_245387 + 8'h01;
  assign sel_245391 = array_index_245278 == array_index_239484 ? add_245390 : sel_245387;
  assign add_245394 = sel_245391 + 8'h01;
  assign sel_245395 = array_index_245278 == array_index_239490 ? add_245394 : sel_245391;
  assign add_245398 = sel_245395 + 8'h01;
  assign sel_245399 = array_index_245278 == array_index_239496 ? add_245398 : sel_245395;
  assign add_245402 = sel_245399 + 8'h01;
  assign sel_245403 = array_index_245278 == array_index_239502 ? add_245402 : sel_245399;
  assign add_245406 = sel_245403 + 8'h01;
  assign sel_245407 = array_index_245278 == array_index_239508 ? add_245406 : sel_245403;
  assign add_245410 = sel_245407 + 8'h01;
  assign sel_245411 = array_index_245278 == array_index_239514 ? add_245410 : sel_245407;
  assign add_245414 = sel_245411 + 8'h01;
  assign sel_245415 = array_index_245278 == array_index_239520 ? add_245414 : sel_245411;
  assign add_245418 = sel_245415 + 8'h01;
  assign sel_245419 = array_index_245278 == array_index_239526 ? add_245418 : sel_245415;
  assign add_245422 = sel_245419 + 8'h01;
  assign sel_245423 = array_index_245278 == array_index_239532 ? add_245422 : sel_245419;
  assign add_245426 = sel_245423 + 8'h01;
  assign sel_245427 = array_index_245278 == array_index_239538 ? add_245426 : sel_245423;
  assign add_245430 = sel_245427 + 8'h01;
  assign sel_245431 = array_index_245278 == array_index_239544 ? add_245430 : sel_245427;
  assign add_245434 = sel_245431 + 8'h01;
  assign sel_245435 = array_index_245278 == array_index_239550 ? add_245434 : sel_245431;
  assign add_245438 = sel_245435 + 8'h01;
  assign sel_245439 = array_index_245278 == array_index_239556 ? add_245438 : sel_245435;
  assign add_245442 = sel_245439 + 8'h01;
  assign sel_245443 = array_index_245278 == array_index_239562 ? add_245442 : sel_245439;
  assign add_245446 = sel_245443 + 8'h01;
  assign sel_245447 = array_index_245278 == array_index_239568 ? add_245446 : sel_245443;
  assign add_245450 = sel_245447 + 8'h01;
  assign sel_245451 = array_index_245278 == array_index_239574 ? add_245450 : sel_245447;
  assign add_245454 = sel_245451 + 8'h01;
  assign sel_245455 = array_index_245278 == array_index_239580 ? add_245454 : sel_245451;
  assign add_245458 = sel_245455 + 8'h01;
  assign sel_245459 = array_index_245278 == array_index_239586 ? add_245458 : sel_245455;
  assign add_245462 = sel_245459 + 8'h01;
  assign sel_245463 = array_index_245278 == array_index_239592 ? add_245462 : sel_245459;
  assign add_245466 = sel_245463 + 8'h01;
  assign sel_245467 = array_index_245278 == array_index_239598 ? add_245466 : sel_245463;
  assign add_245470 = sel_245467 + 8'h01;
  assign sel_245471 = array_index_245278 == array_index_239604 ? add_245470 : sel_245467;
  assign add_245474 = sel_245471 + 8'h01;
  assign sel_245475 = array_index_245278 == array_index_239610 ? add_245474 : sel_245471;
  assign add_245479 = sel_245475 + 8'h01;
  assign array_index_245480 = set1_unflattened[6'h1e];
  assign sel_245481 = array_index_245278 == array_index_239616 ? add_245479 : sel_245475;
  assign add_245484 = sel_245481 + 8'h01;
  assign sel_245485 = array_index_245480 == array_index_239312 ? add_245484 : sel_245481;
  assign add_245488 = sel_245485 + 8'h01;
  assign sel_245489 = array_index_245480 == array_index_239316 ? add_245488 : sel_245485;
  assign add_245492 = sel_245489 + 8'h01;
  assign sel_245493 = array_index_245480 == array_index_239324 ? add_245492 : sel_245489;
  assign add_245496 = sel_245493 + 8'h01;
  assign sel_245497 = array_index_245480 == array_index_239332 ? add_245496 : sel_245493;
  assign add_245500 = sel_245497 + 8'h01;
  assign sel_245501 = array_index_245480 == array_index_239340 ? add_245500 : sel_245497;
  assign add_245504 = sel_245501 + 8'h01;
  assign sel_245505 = array_index_245480 == array_index_239348 ? add_245504 : sel_245501;
  assign add_245508 = sel_245505 + 8'h01;
  assign sel_245509 = array_index_245480 == array_index_239356 ? add_245508 : sel_245505;
  assign add_245512 = sel_245509 + 8'h01;
  assign sel_245513 = array_index_245480 == array_index_239364 ? add_245512 : sel_245509;
  assign add_245516 = sel_245513 + 8'h01;
  assign sel_245517 = array_index_245480 == array_index_239370 ? add_245516 : sel_245513;
  assign add_245520 = sel_245517 + 8'h01;
  assign sel_245521 = array_index_245480 == array_index_239376 ? add_245520 : sel_245517;
  assign add_245524 = sel_245521 + 8'h01;
  assign sel_245525 = array_index_245480 == array_index_239382 ? add_245524 : sel_245521;
  assign add_245528 = sel_245525 + 8'h01;
  assign sel_245529 = array_index_245480 == array_index_239388 ? add_245528 : sel_245525;
  assign add_245532 = sel_245529 + 8'h01;
  assign sel_245533 = array_index_245480 == array_index_239394 ? add_245532 : sel_245529;
  assign add_245536 = sel_245533 + 8'h01;
  assign sel_245537 = array_index_245480 == array_index_239400 ? add_245536 : sel_245533;
  assign add_245540 = sel_245537 + 8'h01;
  assign sel_245541 = array_index_245480 == array_index_239406 ? add_245540 : sel_245537;
  assign add_245544 = sel_245541 + 8'h01;
  assign sel_245545 = array_index_245480 == array_index_239412 ? add_245544 : sel_245541;
  assign add_245548 = sel_245545 + 8'h01;
  assign sel_245549 = array_index_245480 == array_index_239418 ? add_245548 : sel_245545;
  assign add_245552 = sel_245549 + 8'h01;
  assign sel_245553 = array_index_245480 == array_index_239424 ? add_245552 : sel_245549;
  assign add_245556 = sel_245553 + 8'h01;
  assign sel_245557 = array_index_245480 == array_index_239430 ? add_245556 : sel_245553;
  assign add_245560 = sel_245557 + 8'h01;
  assign sel_245561 = array_index_245480 == array_index_239436 ? add_245560 : sel_245557;
  assign add_245564 = sel_245561 + 8'h01;
  assign sel_245565 = array_index_245480 == array_index_239442 ? add_245564 : sel_245561;
  assign add_245568 = sel_245565 + 8'h01;
  assign sel_245569 = array_index_245480 == array_index_239448 ? add_245568 : sel_245565;
  assign add_245572 = sel_245569 + 8'h01;
  assign sel_245573 = array_index_245480 == array_index_239454 ? add_245572 : sel_245569;
  assign add_245576 = sel_245573 + 8'h01;
  assign sel_245577 = array_index_245480 == array_index_239460 ? add_245576 : sel_245573;
  assign add_245580 = sel_245577 + 8'h01;
  assign sel_245581 = array_index_245480 == array_index_239466 ? add_245580 : sel_245577;
  assign add_245584 = sel_245581 + 8'h01;
  assign sel_245585 = array_index_245480 == array_index_239472 ? add_245584 : sel_245581;
  assign add_245588 = sel_245585 + 8'h01;
  assign sel_245589 = array_index_245480 == array_index_239478 ? add_245588 : sel_245585;
  assign add_245592 = sel_245589 + 8'h01;
  assign sel_245593 = array_index_245480 == array_index_239484 ? add_245592 : sel_245589;
  assign add_245596 = sel_245593 + 8'h01;
  assign sel_245597 = array_index_245480 == array_index_239490 ? add_245596 : sel_245593;
  assign add_245600 = sel_245597 + 8'h01;
  assign sel_245601 = array_index_245480 == array_index_239496 ? add_245600 : sel_245597;
  assign add_245604 = sel_245601 + 8'h01;
  assign sel_245605 = array_index_245480 == array_index_239502 ? add_245604 : sel_245601;
  assign add_245608 = sel_245605 + 8'h01;
  assign sel_245609 = array_index_245480 == array_index_239508 ? add_245608 : sel_245605;
  assign add_245612 = sel_245609 + 8'h01;
  assign sel_245613 = array_index_245480 == array_index_239514 ? add_245612 : sel_245609;
  assign add_245616 = sel_245613 + 8'h01;
  assign sel_245617 = array_index_245480 == array_index_239520 ? add_245616 : sel_245613;
  assign add_245620 = sel_245617 + 8'h01;
  assign sel_245621 = array_index_245480 == array_index_239526 ? add_245620 : sel_245617;
  assign add_245624 = sel_245621 + 8'h01;
  assign sel_245625 = array_index_245480 == array_index_239532 ? add_245624 : sel_245621;
  assign add_245628 = sel_245625 + 8'h01;
  assign sel_245629 = array_index_245480 == array_index_239538 ? add_245628 : sel_245625;
  assign add_245632 = sel_245629 + 8'h01;
  assign sel_245633 = array_index_245480 == array_index_239544 ? add_245632 : sel_245629;
  assign add_245636 = sel_245633 + 8'h01;
  assign sel_245637 = array_index_245480 == array_index_239550 ? add_245636 : sel_245633;
  assign add_245640 = sel_245637 + 8'h01;
  assign sel_245641 = array_index_245480 == array_index_239556 ? add_245640 : sel_245637;
  assign add_245644 = sel_245641 + 8'h01;
  assign sel_245645 = array_index_245480 == array_index_239562 ? add_245644 : sel_245641;
  assign add_245648 = sel_245645 + 8'h01;
  assign sel_245649 = array_index_245480 == array_index_239568 ? add_245648 : sel_245645;
  assign add_245652 = sel_245649 + 8'h01;
  assign sel_245653 = array_index_245480 == array_index_239574 ? add_245652 : sel_245649;
  assign add_245656 = sel_245653 + 8'h01;
  assign sel_245657 = array_index_245480 == array_index_239580 ? add_245656 : sel_245653;
  assign add_245660 = sel_245657 + 8'h01;
  assign sel_245661 = array_index_245480 == array_index_239586 ? add_245660 : sel_245657;
  assign add_245664 = sel_245661 + 8'h01;
  assign sel_245665 = array_index_245480 == array_index_239592 ? add_245664 : sel_245661;
  assign add_245668 = sel_245665 + 8'h01;
  assign sel_245669 = array_index_245480 == array_index_239598 ? add_245668 : sel_245665;
  assign add_245672 = sel_245669 + 8'h01;
  assign sel_245673 = array_index_245480 == array_index_239604 ? add_245672 : sel_245669;
  assign add_245676 = sel_245673 + 8'h01;
  assign sel_245677 = array_index_245480 == array_index_239610 ? add_245676 : sel_245673;
  assign add_245681 = sel_245677 + 8'h01;
  assign array_index_245682 = set1_unflattened[6'h1f];
  assign sel_245683 = array_index_245480 == array_index_239616 ? add_245681 : sel_245677;
  assign add_245686 = sel_245683 + 8'h01;
  assign sel_245687 = array_index_245682 == array_index_239312 ? add_245686 : sel_245683;
  assign add_245690 = sel_245687 + 8'h01;
  assign sel_245691 = array_index_245682 == array_index_239316 ? add_245690 : sel_245687;
  assign add_245694 = sel_245691 + 8'h01;
  assign sel_245695 = array_index_245682 == array_index_239324 ? add_245694 : sel_245691;
  assign add_245698 = sel_245695 + 8'h01;
  assign sel_245699 = array_index_245682 == array_index_239332 ? add_245698 : sel_245695;
  assign add_245702 = sel_245699 + 8'h01;
  assign sel_245703 = array_index_245682 == array_index_239340 ? add_245702 : sel_245699;
  assign add_245706 = sel_245703 + 8'h01;
  assign sel_245707 = array_index_245682 == array_index_239348 ? add_245706 : sel_245703;
  assign add_245710 = sel_245707 + 8'h01;
  assign sel_245711 = array_index_245682 == array_index_239356 ? add_245710 : sel_245707;
  assign add_245714 = sel_245711 + 8'h01;
  assign sel_245715 = array_index_245682 == array_index_239364 ? add_245714 : sel_245711;
  assign add_245718 = sel_245715 + 8'h01;
  assign sel_245719 = array_index_245682 == array_index_239370 ? add_245718 : sel_245715;
  assign add_245722 = sel_245719 + 8'h01;
  assign sel_245723 = array_index_245682 == array_index_239376 ? add_245722 : sel_245719;
  assign add_245726 = sel_245723 + 8'h01;
  assign sel_245727 = array_index_245682 == array_index_239382 ? add_245726 : sel_245723;
  assign add_245730 = sel_245727 + 8'h01;
  assign sel_245731 = array_index_245682 == array_index_239388 ? add_245730 : sel_245727;
  assign add_245734 = sel_245731 + 8'h01;
  assign sel_245735 = array_index_245682 == array_index_239394 ? add_245734 : sel_245731;
  assign add_245738 = sel_245735 + 8'h01;
  assign sel_245739 = array_index_245682 == array_index_239400 ? add_245738 : sel_245735;
  assign add_245742 = sel_245739 + 8'h01;
  assign sel_245743 = array_index_245682 == array_index_239406 ? add_245742 : sel_245739;
  assign add_245746 = sel_245743 + 8'h01;
  assign sel_245747 = array_index_245682 == array_index_239412 ? add_245746 : sel_245743;
  assign add_245750 = sel_245747 + 8'h01;
  assign sel_245751 = array_index_245682 == array_index_239418 ? add_245750 : sel_245747;
  assign add_245754 = sel_245751 + 8'h01;
  assign sel_245755 = array_index_245682 == array_index_239424 ? add_245754 : sel_245751;
  assign add_245758 = sel_245755 + 8'h01;
  assign sel_245759 = array_index_245682 == array_index_239430 ? add_245758 : sel_245755;
  assign add_245762 = sel_245759 + 8'h01;
  assign sel_245763 = array_index_245682 == array_index_239436 ? add_245762 : sel_245759;
  assign add_245766 = sel_245763 + 8'h01;
  assign sel_245767 = array_index_245682 == array_index_239442 ? add_245766 : sel_245763;
  assign add_245770 = sel_245767 + 8'h01;
  assign sel_245771 = array_index_245682 == array_index_239448 ? add_245770 : sel_245767;
  assign add_245774 = sel_245771 + 8'h01;
  assign sel_245775 = array_index_245682 == array_index_239454 ? add_245774 : sel_245771;
  assign add_245778 = sel_245775 + 8'h01;
  assign sel_245779 = array_index_245682 == array_index_239460 ? add_245778 : sel_245775;
  assign add_245782 = sel_245779 + 8'h01;
  assign sel_245783 = array_index_245682 == array_index_239466 ? add_245782 : sel_245779;
  assign add_245786 = sel_245783 + 8'h01;
  assign sel_245787 = array_index_245682 == array_index_239472 ? add_245786 : sel_245783;
  assign add_245790 = sel_245787 + 8'h01;
  assign sel_245791 = array_index_245682 == array_index_239478 ? add_245790 : sel_245787;
  assign add_245794 = sel_245791 + 8'h01;
  assign sel_245795 = array_index_245682 == array_index_239484 ? add_245794 : sel_245791;
  assign add_245798 = sel_245795 + 8'h01;
  assign sel_245799 = array_index_245682 == array_index_239490 ? add_245798 : sel_245795;
  assign add_245802 = sel_245799 + 8'h01;
  assign sel_245803 = array_index_245682 == array_index_239496 ? add_245802 : sel_245799;
  assign add_245806 = sel_245803 + 8'h01;
  assign sel_245807 = array_index_245682 == array_index_239502 ? add_245806 : sel_245803;
  assign add_245810 = sel_245807 + 8'h01;
  assign sel_245811 = array_index_245682 == array_index_239508 ? add_245810 : sel_245807;
  assign add_245814 = sel_245811 + 8'h01;
  assign sel_245815 = array_index_245682 == array_index_239514 ? add_245814 : sel_245811;
  assign add_245818 = sel_245815 + 8'h01;
  assign sel_245819 = array_index_245682 == array_index_239520 ? add_245818 : sel_245815;
  assign add_245822 = sel_245819 + 8'h01;
  assign sel_245823 = array_index_245682 == array_index_239526 ? add_245822 : sel_245819;
  assign add_245826 = sel_245823 + 8'h01;
  assign sel_245827 = array_index_245682 == array_index_239532 ? add_245826 : sel_245823;
  assign add_245830 = sel_245827 + 8'h01;
  assign sel_245831 = array_index_245682 == array_index_239538 ? add_245830 : sel_245827;
  assign add_245834 = sel_245831 + 8'h01;
  assign sel_245835 = array_index_245682 == array_index_239544 ? add_245834 : sel_245831;
  assign add_245838 = sel_245835 + 8'h01;
  assign sel_245839 = array_index_245682 == array_index_239550 ? add_245838 : sel_245835;
  assign add_245842 = sel_245839 + 8'h01;
  assign sel_245843 = array_index_245682 == array_index_239556 ? add_245842 : sel_245839;
  assign add_245846 = sel_245843 + 8'h01;
  assign sel_245847 = array_index_245682 == array_index_239562 ? add_245846 : sel_245843;
  assign add_245850 = sel_245847 + 8'h01;
  assign sel_245851 = array_index_245682 == array_index_239568 ? add_245850 : sel_245847;
  assign add_245854 = sel_245851 + 8'h01;
  assign sel_245855 = array_index_245682 == array_index_239574 ? add_245854 : sel_245851;
  assign add_245858 = sel_245855 + 8'h01;
  assign sel_245859 = array_index_245682 == array_index_239580 ? add_245858 : sel_245855;
  assign add_245862 = sel_245859 + 8'h01;
  assign sel_245863 = array_index_245682 == array_index_239586 ? add_245862 : sel_245859;
  assign add_245866 = sel_245863 + 8'h01;
  assign sel_245867 = array_index_245682 == array_index_239592 ? add_245866 : sel_245863;
  assign add_245870 = sel_245867 + 8'h01;
  assign sel_245871 = array_index_245682 == array_index_239598 ? add_245870 : sel_245867;
  assign add_245874 = sel_245871 + 8'h01;
  assign sel_245875 = array_index_245682 == array_index_239604 ? add_245874 : sel_245871;
  assign add_245878 = sel_245875 + 8'h01;
  assign sel_245879 = array_index_245682 == array_index_239610 ? add_245878 : sel_245875;
  assign add_245883 = sel_245879 + 8'h01;
  assign array_index_245884 = set1_unflattened[6'h20];
  assign sel_245885 = array_index_245682 == array_index_239616 ? add_245883 : sel_245879;
  assign add_245888 = sel_245885 + 8'h01;
  assign sel_245889 = array_index_245884 == array_index_239312 ? add_245888 : sel_245885;
  assign add_245892 = sel_245889 + 8'h01;
  assign sel_245893 = array_index_245884 == array_index_239316 ? add_245892 : sel_245889;
  assign add_245896 = sel_245893 + 8'h01;
  assign sel_245897 = array_index_245884 == array_index_239324 ? add_245896 : sel_245893;
  assign add_245900 = sel_245897 + 8'h01;
  assign sel_245901 = array_index_245884 == array_index_239332 ? add_245900 : sel_245897;
  assign add_245904 = sel_245901 + 8'h01;
  assign sel_245905 = array_index_245884 == array_index_239340 ? add_245904 : sel_245901;
  assign add_245908 = sel_245905 + 8'h01;
  assign sel_245909 = array_index_245884 == array_index_239348 ? add_245908 : sel_245905;
  assign add_245912 = sel_245909 + 8'h01;
  assign sel_245913 = array_index_245884 == array_index_239356 ? add_245912 : sel_245909;
  assign add_245916 = sel_245913 + 8'h01;
  assign sel_245917 = array_index_245884 == array_index_239364 ? add_245916 : sel_245913;
  assign add_245920 = sel_245917 + 8'h01;
  assign sel_245921 = array_index_245884 == array_index_239370 ? add_245920 : sel_245917;
  assign add_245924 = sel_245921 + 8'h01;
  assign sel_245925 = array_index_245884 == array_index_239376 ? add_245924 : sel_245921;
  assign add_245928 = sel_245925 + 8'h01;
  assign sel_245929 = array_index_245884 == array_index_239382 ? add_245928 : sel_245925;
  assign add_245932 = sel_245929 + 8'h01;
  assign sel_245933 = array_index_245884 == array_index_239388 ? add_245932 : sel_245929;
  assign add_245936 = sel_245933 + 8'h01;
  assign sel_245937 = array_index_245884 == array_index_239394 ? add_245936 : sel_245933;
  assign add_245940 = sel_245937 + 8'h01;
  assign sel_245941 = array_index_245884 == array_index_239400 ? add_245940 : sel_245937;
  assign add_245944 = sel_245941 + 8'h01;
  assign sel_245945 = array_index_245884 == array_index_239406 ? add_245944 : sel_245941;
  assign add_245948 = sel_245945 + 8'h01;
  assign sel_245949 = array_index_245884 == array_index_239412 ? add_245948 : sel_245945;
  assign add_245952 = sel_245949 + 8'h01;
  assign sel_245953 = array_index_245884 == array_index_239418 ? add_245952 : sel_245949;
  assign add_245956 = sel_245953 + 8'h01;
  assign sel_245957 = array_index_245884 == array_index_239424 ? add_245956 : sel_245953;
  assign add_245960 = sel_245957 + 8'h01;
  assign sel_245961 = array_index_245884 == array_index_239430 ? add_245960 : sel_245957;
  assign add_245964 = sel_245961 + 8'h01;
  assign sel_245965 = array_index_245884 == array_index_239436 ? add_245964 : sel_245961;
  assign add_245968 = sel_245965 + 8'h01;
  assign sel_245969 = array_index_245884 == array_index_239442 ? add_245968 : sel_245965;
  assign add_245972 = sel_245969 + 8'h01;
  assign sel_245973 = array_index_245884 == array_index_239448 ? add_245972 : sel_245969;
  assign add_245976 = sel_245973 + 8'h01;
  assign sel_245977 = array_index_245884 == array_index_239454 ? add_245976 : sel_245973;
  assign add_245980 = sel_245977 + 8'h01;
  assign sel_245981 = array_index_245884 == array_index_239460 ? add_245980 : sel_245977;
  assign add_245984 = sel_245981 + 8'h01;
  assign sel_245985 = array_index_245884 == array_index_239466 ? add_245984 : sel_245981;
  assign add_245988 = sel_245985 + 8'h01;
  assign sel_245989 = array_index_245884 == array_index_239472 ? add_245988 : sel_245985;
  assign add_245992 = sel_245989 + 8'h01;
  assign sel_245993 = array_index_245884 == array_index_239478 ? add_245992 : sel_245989;
  assign add_245996 = sel_245993 + 8'h01;
  assign sel_245997 = array_index_245884 == array_index_239484 ? add_245996 : sel_245993;
  assign add_246000 = sel_245997 + 8'h01;
  assign sel_246001 = array_index_245884 == array_index_239490 ? add_246000 : sel_245997;
  assign add_246004 = sel_246001 + 8'h01;
  assign sel_246005 = array_index_245884 == array_index_239496 ? add_246004 : sel_246001;
  assign add_246008 = sel_246005 + 8'h01;
  assign sel_246009 = array_index_245884 == array_index_239502 ? add_246008 : sel_246005;
  assign add_246012 = sel_246009 + 8'h01;
  assign sel_246013 = array_index_245884 == array_index_239508 ? add_246012 : sel_246009;
  assign add_246016 = sel_246013 + 8'h01;
  assign sel_246017 = array_index_245884 == array_index_239514 ? add_246016 : sel_246013;
  assign add_246020 = sel_246017 + 8'h01;
  assign sel_246021 = array_index_245884 == array_index_239520 ? add_246020 : sel_246017;
  assign add_246024 = sel_246021 + 8'h01;
  assign sel_246025 = array_index_245884 == array_index_239526 ? add_246024 : sel_246021;
  assign add_246028 = sel_246025 + 8'h01;
  assign sel_246029 = array_index_245884 == array_index_239532 ? add_246028 : sel_246025;
  assign add_246032 = sel_246029 + 8'h01;
  assign sel_246033 = array_index_245884 == array_index_239538 ? add_246032 : sel_246029;
  assign add_246036 = sel_246033 + 8'h01;
  assign sel_246037 = array_index_245884 == array_index_239544 ? add_246036 : sel_246033;
  assign add_246040 = sel_246037 + 8'h01;
  assign sel_246041 = array_index_245884 == array_index_239550 ? add_246040 : sel_246037;
  assign add_246044 = sel_246041 + 8'h01;
  assign sel_246045 = array_index_245884 == array_index_239556 ? add_246044 : sel_246041;
  assign add_246048 = sel_246045 + 8'h01;
  assign sel_246049 = array_index_245884 == array_index_239562 ? add_246048 : sel_246045;
  assign add_246052 = sel_246049 + 8'h01;
  assign sel_246053 = array_index_245884 == array_index_239568 ? add_246052 : sel_246049;
  assign add_246056 = sel_246053 + 8'h01;
  assign sel_246057 = array_index_245884 == array_index_239574 ? add_246056 : sel_246053;
  assign add_246060 = sel_246057 + 8'h01;
  assign sel_246061 = array_index_245884 == array_index_239580 ? add_246060 : sel_246057;
  assign add_246064 = sel_246061 + 8'h01;
  assign sel_246065 = array_index_245884 == array_index_239586 ? add_246064 : sel_246061;
  assign add_246068 = sel_246065 + 8'h01;
  assign sel_246069 = array_index_245884 == array_index_239592 ? add_246068 : sel_246065;
  assign add_246072 = sel_246069 + 8'h01;
  assign sel_246073 = array_index_245884 == array_index_239598 ? add_246072 : sel_246069;
  assign add_246076 = sel_246073 + 8'h01;
  assign sel_246077 = array_index_245884 == array_index_239604 ? add_246076 : sel_246073;
  assign add_246080 = sel_246077 + 8'h01;
  assign sel_246081 = array_index_245884 == array_index_239610 ? add_246080 : sel_246077;
  assign add_246085 = sel_246081 + 8'h01;
  assign array_index_246086 = set1_unflattened[6'h21];
  assign sel_246087 = array_index_245884 == array_index_239616 ? add_246085 : sel_246081;
  assign add_246090 = sel_246087 + 8'h01;
  assign sel_246091 = array_index_246086 == array_index_239312 ? add_246090 : sel_246087;
  assign add_246094 = sel_246091 + 8'h01;
  assign sel_246095 = array_index_246086 == array_index_239316 ? add_246094 : sel_246091;
  assign add_246098 = sel_246095 + 8'h01;
  assign sel_246099 = array_index_246086 == array_index_239324 ? add_246098 : sel_246095;
  assign add_246102 = sel_246099 + 8'h01;
  assign sel_246103 = array_index_246086 == array_index_239332 ? add_246102 : sel_246099;
  assign add_246106 = sel_246103 + 8'h01;
  assign sel_246107 = array_index_246086 == array_index_239340 ? add_246106 : sel_246103;
  assign add_246110 = sel_246107 + 8'h01;
  assign sel_246111 = array_index_246086 == array_index_239348 ? add_246110 : sel_246107;
  assign add_246114 = sel_246111 + 8'h01;
  assign sel_246115 = array_index_246086 == array_index_239356 ? add_246114 : sel_246111;
  assign add_246118 = sel_246115 + 8'h01;
  assign sel_246119 = array_index_246086 == array_index_239364 ? add_246118 : sel_246115;
  assign add_246122 = sel_246119 + 8'h01;
  assign sel_246123 = array_index_246086 == array_index_239370 ? add_246122 : sel_246119;
  assign add_246126 = sel_246123 + 8'h01;
  assign sel_246127 = array_index_246086 == array_index_239376 ? add_246126 : sel_246123;
  assign add_246130 = sel_246127 + 8'h01;
  assign sel_246131 = array_index_246086 == array_index_239382 ? add_246130 : sel_246127;
  assign add_246134 = sel_246131 + 8'h01;
  assign sel_246135 = array_index_246086 == array_index_239388 ? add_246134 : sel_246131;
  assign add_246138 = sel_246135 + 8'h01;
  assign sel_246139 = array_index_246086 == array_index_239394 ? add_246138 : sel_246135;
  assign add_246142 = sel_246139 + 8'h01;
  assign sel_246143 = array_index_246086 == array_index_239400 ? add_246142 : sel_246139;
  assign add_246146 = sel_246143 + 8'h01;
  assign sel_246147 = array_index_246086 == array_index_239406 ? add_246146 : sel_246143;
  assign add_246150 = sel_246147 + 8'h01;
  assign sel_246151 = array_index_246086 == array_index_239412 ? add_246150 : sel_246147;
  assign add_246154 = sel_246151 + 8'h01;
  assign sel_246155 = array_index_246086 == array_index_239418 ? add_246154 : sel_246151;
  assign add_246158 = sel_246155 + 8'h01;
  assign sel_246159 = array_index_246086 == array_index_239424 ? add_246158 : sel_246155;
  assign add_246162 = sel_246159 + 8'h01;
  assign sel_246163 = array_index_246086 == array_index_239430 ? add_246162 : sel_246159;
  assign add_246166 = sel_246163 + 8'h01;
  assign sel_246167 = array_index_246086 == array_index_239436 ? add_246166 : sel_246163;
  assign add_246170 = sel_246167 + 8'h01;
  assign sel_246171 = array_index_246086 == array_index_239442 ? add_246170 : sel_246167;
  assign add_246174 = sel_246171 + 8'h01;
  assign sel_246175 = array_index_246086 == array_index_239448 ? add_246174 : sel_246171;
  assign add_246178 = sel_246175 + 8'h01;
  assign sel_246179 = array_index_246086 == array_index_239454 ? add_246178 : sel_246175;
  assign add_246182 = sel_246179 + 8'h01;
  assign sel_246183 = array_index_246086 == array_index_239460 ? add_246182 : sel_246179;
  assign add_246186 = sel_246183 + 8'h01;
  assign sel_246187 = array_index_246086 == array_index_239466 ? add_246186 : sel_246183;
  assign add_246190 = sel_246187 + 8'h01;
  assign sel_246191 = array_index_246086 == array_index_239472 ? add_246190 : sel_246187;
  assign add_246194 = sel_246191 + 8'h01;
  assign sel_246195 = array_index_246086 == array_index_239478 ? add_246194 : sel_246191;
  assign add_246198 = sel_246195 + 8'h01;
  assign sel_246199 = array_index_246086 == array_index_239484 ? add_246198 : sel_246195;
  assign add_246202 = sel_246199 + 8'h01;
  assign sel_246203 = array_index_246086 == array_index_239490 ? add_246202 : sel_246199;
  assign add_246206 = sel_246203 + 8'h01;
  assign sel_246207 = array_index_246086 == array_index_239496 ? add_246206 : sel_246203;
  assign add_246210 = sel_246207 + 8'h01;
  assign sel_246211 = array_index_246086 == array_index_239502 ? add_246210 : sel_246207;
  assign add_246214 = sel_246211 + 8'h01;
  assign sel_246215 = array_index_246086 == array_index_239508 ? add_246214 : sel_246211;
  assign add_246218 = sel_246215 + 8'h01;
  assign sel_246219 = array_index_246086 == array_index_239514 ? add_246218 : sel_246215;
  assign add_246222 = sel_246219 + 8'h01;
  assign sel_246223 = array_index_246086 == array_index_239520 ? add_246222 : sel_246219;
  assign add_246226 = sel_246223 + 8'h01;
  assign sel_246227 = array_index_246086 == array_index_239526 ? add_246226 : sel_246223;
  assign add_246230 = sel_246227 + 8'h01;
  assign sel_246231 = array_index_246086 == array_index_239532 ? add_246230 : sel_246227;
  assign add_246234 = sel_246231 + 8'h01;
  assign sel_246235 = array_index_246086 == array_index_239538 ? add_246234 : sel_246231;
  assign add_246238 = sel_246235 + 8'h01;
  assign sel_246239 = array_index_246086 == array_index_239544 ? add_246238 : sel_246235;
  assign add_246242 = sel_246239 + 8'h01;
  assign sel_246243 = array_index_246086 == array_index_239550 ? add_246242 : sel_246239;
  assign add_246246 = sel_246243 + 8'h01;
  assign sel_246247 = array_index_246086 == array_index_239556 ? add_246246 : sel_246243;
  assign add_246250 = sel_246247 + 8'h01;
  assign sel_246251 = array_index_246086 == array_index_239562 ? add_246250 : sel_246247;
  assign add_246254 = sel_246251 + 8'h01;
  assign sel_246255 = array_index_246086 == array_index_239568 ? add_246254 : sel_246251;
  assign add_246258 = sel_246255 + 8'h01;
  assign sel_246259 = array_index_246086 == array_index_239574 ? add_246258 : sel_246255;
  assign add_246262 = sel_246259 + 8'h01;
  assign sel_246263 = array_index_246086 == array_index_239580 ? add_246262 : sel_246259;
  assign add_246266 = sel_246263 + 8'h01;
  assign sel_246267 = array_index_246086 == array_index_239586 ? add_246266 : sel_246263;
  assign add_246270 = sel_246267 + 8'h01;
  assign sel_246271 = array_index_246086 == array_index_239592 ? add_246270 : sel_246267;
  assign add_246274 = sel_246271 + 8'h01;
  assign sel_246275 = array_index_246086 == array_index_239598 ? add_246274 : sel_246271;
  assign add_246278 = sel_246275 + 8'h01;
  assign sel_246279 = array_index_246086 == array_index_239604 ? add_246278 : sel_246275;
  assign add_246282 = sel_246279 + 8'h01;
  assign sel_246283 = array_index_246086 == array_index_239610 ? add_246282 : sel_246279;
  assign add_246287 = sel_246283 + 8'h01;
  assign array_index_246288 = set1_unflattened[6'h22];
  assign sel_246289 = array_index_246086 == array_index_239616 ? add_246287 : sel_246283;
  assign add_246292 = sel_246289 + 8'h01;
  assign sel_246293 = array_index_246288 == array_index_239312 ? add_246292 : sel_246289;
  assign add_246296 = sel_246293 + 8'h01;
  assign sel_246297 = array_index_246288 == array_index_239316 ? add_246296 : sel_246293;
  assign add_246300 = sel_246297 + 8'h01;
  assign sel_246301 = array_index_246288 == array_index_239324 ? add_246300 : sel_246297;
  assign add_246304 = sel_246301 + 8'h01;
  assign sel_246305 = array_index_246288 == array_index_239332 ? add_246304 : sel_246301;
  assign add_246308 = sel_246305 + 8'h01;
  assign sel_246309 = array_index_246288 == array_index_239340 ? add_246308 : sel_246305;
  assign add_246312 = sel_246309 + 8'h01;
  assign sel_246313 = array_index_246288 == array_index_239348 ? add_246312 : sel_246309;
  assign add_246316 = sel_246313 + 8'h01;
  assign sel_246317 = array_index_246288 == array_index_239356 ? add_246316 : sel_246313;
  assign add_246320 = sel_246317 + 8'h01;
  assign sel_246321 = array_index_246288 == array_index_239364 ? add_246320 : sel_246317;
  assign add_246324 = sel_246321 + 8'h01;
  assign sel_246325 = array_index_246288 == array_index_239370 ? add_246324 : sel_246321;
  assign add_246328 = sel_246325 + 8'h01;
  assign sel_246329 = array_index_246288 == array_index_239376 ? add_246328 : sel_246325;
  assign add_246332 = sel_246329 + 8'h01;
  assign sel_246333 = array_index_246288 == array_index_239382 ? add_246332 : sel_246329;
  assign add_246336 = sel_246333 + 8'h01;
  assign sel_246337 = array_index_246288 == array_index_239388 ? add_246336 : sel_246333;
  assign add_246340 = sel_246337 + 8'h01;
  assign sel_246341 = array_index_246288 == array_index_239394 ? add_246340 : sel_246337;
  assign add_246344 = sel_246341 + 8'h01;
  assign sel_246345 = array_index_246288 == array_index_239400 ? add_246344 : sel_246341;
  assign add_246348 = sel_246345 + 8'h01;
  assign sel_246349 = array_index_246288 == array_index_239406 ? add_246348 : sel_246345;
  assign add_246352 = sel_246349 + 8'h01;
  assign sel_246353 = array_index_246288 == array_index_239412 ? add_246352 : sel_246349;
  assign add_246356 = sel_246353 + 8'h01;
  assign sel_246357 = array_index_246288 == array_index_239418 ? add_246356 : sel_246353;
  assign add_246360 = sel_246357 + 8'h01;
  assign sel_246361 = array_index_246288 == array_index_239424 ? add_246360 : sel_246357;
  assign add_246364 = sel_246361 + 8'h01;
  assign sel_246365 = array_index_246288 == array_index_239430 ? add_246364 : sel_246361;
  assign add_246368 = sel_246365 + 8'h01;
  assign sel_246369 = array_index_246288 == array_index_239436 ? add_246368 : sel_246365;
  assign add_246372 = sel_246369 + 8'h01;
  assign sel_246373 = array_index_246288 == array_index_239442 ? add_246372 : sel_246369;
  assign add_246376 = sel_246373 + 8'h01;
  assign sel_246377 = array_index_246288 == array_index_239448 ? add_246376 : sel_246373;
  assign add_246380 = sel_246377 + 8'h01;
  assign sel_246381 = array_index_246288 == array_index_239454 ? add_246380 : sel_246377;
  assign add_246384 = sel_246381 + 8'h01;
  assign sel_246385 = array_index_246288 == array_index_239460 ? add_246384 : sel_246381;
  assign add_246388 = sel_246385 + 8'h01;
  assign sel_246389 = array_index_246288 == array_index_239466 ? add_246388 : sel_246385;
  assign add_246392 = sel_246389 + 8'h01;
  assign sel_246393 = array_index_246288 == array_index_239472 ? add_246392 : sel_246389;
  assign add_246396 = sel_246393 + 8'h01;
  assign sel_246397 = array_index_246288 == array_index_239478 ? add_246396 : sel_246393;
  assign add_246400 = sel_246397 + 8'h01;
  assign sel_246401 = array_index_246288 == array_index_239484 ? add_246400 : sel_246397;
  assign add_246404 = sel_246401 + 8'h01;
  assign sel_246405 = array_index_246288 == array_index_239490 ? add_246404 : sel_246401;
  assign add_246408 = sel_246405 + 8'h01;
  assign sel_246409 = array_index_246288 == array_index_239496 ? add_246408 : sel_246405;
  assign add_246412 = sel_246409 + 8'h01;
  assign sel_246413 = array_index_246288 == array_index_239502 ? add_246412 : sel_246409;
  assign add_246416 = sel_246413 + 8'h01;
  assign sel_246417 = array_index_246288 == array_index_239508 ? add_246416 : sel_246413;
  assign add_246420 = sel_246417 + 8'h01;
  assign sel_246421 = array_index_246288 == array_index_239514 ? add_246420 : sel_246417;
  assign add_246424 = sel_246421 + 8'h01;
  assign sel_246425 = array_index_246288 == array_index_239520 ? add_246424 : sel_246421;
  assign add_246428 = sel_246425 + 8'h01;
  assign sel_246429 = array_index_246288 == array_index_239526 ? add_246428 : sel_246425;
  assign add_246432 = sel_246429 + 8'h01;
  assign sel_246433 = array_index_246288 == array_index_239532 ? add_246432 : sel_246429;
  assign add_246436 = sel_246433 + 8'h01;
  assign sel_246437 = array_index_246288 == array_index_239538 ? add_246436 : sel_246433;
  assign add_246440 = sel_246437 + 8'h01;
  assign sel_246441 = array_index_246288 == array_index_239544 ? add_246440 : sel_246437;
  assign add_246444 = sel_246441 + 8'h01;
  assign sel_246445 = array_index_246288 == array_index_239550 ? add_246444 : sel_246441;
  assign add_246448 = sel_246445 + 8'h01;
  assign sel_246449 = array_index_246288 == array_index_239556 ? add_246448 : sel_246445;
  assign add_246452 = sel_246449 + 8'h01;
  assign sel_246453 = array_index_246288 == array_index_239562 ? add_246452 : sel_246449;
  assign add_246456 = sel_246453 + 8'h01;
  assign sel_246457 = array_index_246288 == array_index_239568 ? add_246456 : sel_246453;
  assign add_246460 = sel_246457 + 8'h01;
  assign sel_246461 = array_index_246288 == array_index_239574 ? add_246460 : sel_246457;
  assign add_246464 = sel_246461 + 8'h01;
  assign sel_246465 = array_index_246288 == array_index_239580 ? add_246464 : sel_246461;
  assign add_246468 = sel_246465 + 8'h01;
  assign sel_246469 = array_index_246288 == array_index_239586 ? add_246468 : sel_246465;
  assign add_246472 = sel_246469 + 8'h01;
  assign sel_246473 = array_index_246288 == array_index_239592 ? add_246472 : sel_246469;
  assign add_246476 = sel_246473 + 8'h01;
  assign sel_246477 = array_index_246288 == array_index_239598 ? add_246476 : sel_246473;
  assign add_246480 = sel_246477 + 8'h01;
  assign sel_246481 = array_index_246288 == array_index_239604 ? add_246480 : sel_246477;
  assign add_246484 = sel_246481 + 8'h01;
  assign sel_246485 = array_index_246288 == array_index_239610 ? add_246484 : sel_246481;
  assign add_246489 = sel_246485 + 8'h01;
  assign array_index_246490 = set1_unflattened[6'h23];
  assign sel_246491 = array_index_246288 == array_index_239616 ? add_246489 : sel_246485;
  assign add_246494 = sel_246491 + 8'h01;
  assign sel_246495 = array_index_246490 == array_index_239312 ? add_246494 : sel_246491;
  assign add_246498 = sel_246495 + 8'h01;
  assign sel_246499 = array_index_246490 == array_index_239316 ? add_246498 : sel_246495;
  assign add_246502 = sel_246499 + 8'h01;
  assign sel_246503 = array_index_246490 == array_index_239324 ? add_246502 : sel_246499;
  assign add_246506 = sel_246503 + 8'h01;
  assign sel_246507 = array_index_246490 == array_index_239332 ? add_246506 : sel_246503;
  assign add_246510 = sel_246507 + 8'h01;
  assign sel_246511 = array_index_246490 == array_index_239340 ? add_246510 : sel_246507;
  assign add_246514 = sel_246511 + 8'h01;
  assign sel_246515 = array_index_246490 == array_index_239348 ? add_246514 : sel_246511;
  assign add_246518 = sel_246515 + 8'h01;
  assign sel_246519 = array_index_246490 == array_index_239356 ? add_246518 : sel_246515;
  assign add_246522 = sel_246519 + 8'h01;
  assign sel_246523 = array_index_246490 == array_index_239364 ? add_246522 : sel_246519;
  assign add_246526 = sel_246523 + 8'h01;
  assign sel_246527 = array_index_246490 == array_index_239370 ? add_246526 : sel_246523;
  assign add_246530 = sel_246527 + 8'h01;
  assign sel_246531 = array_index_246490 == array_index_239376 ? add_246530 : sel_246527;
  assign add_246534 = sel_246531 + 8'h01;
  assign sel_246535 = array_index_246490 == array_index_239382 ? add_246534 : sel_246531;
  assign add_246538 = sel_246535 + 8'h01;
  assign sel_246539 = array_index_246490 == array_index_239388 ? add_246538 : sel_246535;
  assign add_246542 = sel_246539 + 8'h01;
  assign sel_246543 = array_index_246490 == array_index_239394 ? add_246542 : sel_246539;
  assign add_246546 = sel_246543 + 8'h01;
  assign sel_246547 = array_index_246490 == array_index_239400 ? add_246546 : sel_246543;
  assign add_246550 = sel_246547 + 8'h01;
  assign sel_246551 = array_index_246490 == array_index_239406 ? add_246550 : sel_246547;
  assign add_246554 = sel_246551 + 8'h01;
  assign sel_246555 = array_index_246490 == array_index_239412 ? add_246554 : sel_246551;
  assign add_246558 = sel_246555 + 8'h01;
  assign sel_246559 = array_index_246490 == array_index_239418 ? add_246558 : sel_246555;
  assign add_246562 = sel_246559 + 8'h01;
  assign sel_246563 = array_index_246490 == array_index_239424 ? add_246562 : sel_246559;
  assign add_246566 = sel_246563 + 8'h01;
  assign sel_246567 = array_index_246490 == array_index_239430 ? add_246566 : sel_246563;
  assign add_246570 = sel_246567 + 8'h01;
  assign sel_246571 = array_index_246490 == array_index_239436 ? add_246570 : sel_246567;
  assign add_246574 = sel_246571 + 8'h01;
  assign sel_246575 = array_index_246490 == array_index_239442 ? add_246574 : sel_246571;
  assign add_246578 = sel_246575 + 8'h01;
  assign sel_246579 = array_index_246490 == array_index_239448 ? add_246578 : sel_246575;
  assign add_246582 = sel_246579 + 8'h01;
  assign sel_246583 = array_index_246490 == array_index_239454 ? add_246582 : sel_246579;
  assign add_246586 = sel_246583 + 8'h01;
  assign sel_246587 = array_index_246490 == array_index_239460 ? add_246586 : sel_246583;
  assign add_246590 = sel_246587 + 8'h01;
  assign sel_246591 = array_index_246490 == array_index_239466 ? add_246590 : sel_246587;
  assign add_246594 = sel_246591 + 8'h01;
  assign sel_246595 = array_index_246490 == array_index_239472 ? add_246594 : sel_246591;
  assign add_246598 = sel_246595 + 8'h01;
  assign sel_246599 = array_index_246490 == array_index_239478 ? add_246598 : sel_246595;
  assign add_246602 = sel_246599 + 8'h01;
  assign sel_246603 = array_index_246490 == array_index_239484 ? add_246602 : sel_246599;
  assign add_246606 = sel_246603 + 8'h01;
  assign sel_246607 = array_index_246490 == array_index_239490 ? add_246606 : sel_246603;
  assign add_246610 = sel_246607 + 8'h01;
  assign sel_246611 = array_index_246490 == array_index_239496 ? add_246610 : sel_246607;
  assign add_246614 = sel_246611 + 8'h01;
  assign sel_246615 = array_index_246490 == array_index_239502 ? add_246614 : sel_246611;
  assign add_246618 = sel_246615 + 8'h01;
  assign sel_246619 = array_index_246490 == array_index_239508 ? add_246618 : sel_246615;
  assign add_246622 = sel_246619 + 8'h01;
  assign sel_246623 = array_index_246490 == array_index_239514 ? add_246622 : sel_246619;
  assign add_246626 = sel_246623 + 8'h01;
  assign sel_246627 = array_index_246490 == array_index_239520 ? add_246626 : sel_246623;
  assign add_246630 = sel_246627 + 8'h01;
  assign sel_246631 = array_index_246490 == array_index_239526 ? add_246630 : sel_246627;
  assign add_246634 = sel_246631 + 8'h01;
  assign sel_246635 = array_index_246490 == array_index_239532 ? add_246634 : sel_246631;
  assign add_246638 = sel_246635 + 8'h01;
  assign sel_246639 = array_index_246490 == array_index_239538 ? add_246638 : sel_246635;
  assign add_246642 = sel_246639 + 8'h01;
  assign sel_246643 = array_index_246490 == array_index_239544 ? add_246642 : sel_246639;
  assign add_246646 = sel_246643 + 8'h01;
  assign sel_246647 = array_index_246490 == array_index_239550 ? add_246646 : sel_246643;
  assign add_246650 = sel_246647 + 8'h01;
  assign sel_246651 = array_index_246490 == array_index_239556 ? add_246650 : sel_246647;
  assign add_246654 = sel_246651 + 8'h01;
  assign sel_246655 = array_index_246490 == array_index_239562 ? add_246654 : sel_246651;
  assign add_246658 = sel_246655 + 8'h01;
  assign sel_246659 = array_index_246490 == array_index_239568 ? add_246658 : sel_246655;
  assign add_246662 = sel_246659 + 8'h01;
  assign sel_246663 = array_index_246490 == array_index_239574 ? add_246662 : sel_246659;
  assign add_246666 = sel_246663 + 8'h01;
  assign sel_246667 = array_index_246490 == array_index_239580 ? add_246666 : sel_246663;
  assign add_246670 = sel_246667 + 8'h01;
  assign sel_246671 = array_index_246490 == array_index_239586 ? add_246670 : sel_246667;
  assign add_246674 = sel_246671 + 8'h01;
  assign sel_246675 = array_index_246490 == array_index_239592 ? add_246674 : sel_246671;
  assign add_246678 = sel_246675 + 8'h01;
  assign sel_246679 = array_index_246490 == array_index_239598 ? add_246678 : sel_246675;
  assign add_246682 = sel_246679 + 8'h01;
  assign sel_246683 = array_index_246490 == array_index_239604 ? add_246682 : sel_246679;
  assign add_246686 = sel_246683 + 8'h01;
  assign sel_246687 = array_index_246490 == array_index_239610 ? add_246686 : sel_246683;
  assign add_246691 = sel_246687 + 8'h01;
  assign array_index_246692 = set1_unflattened[6'h24];
  assign sel_246693 = array_index_246490 == array_index_239616 ? add_246691 : sel_246687;
  assign add_246696 = sel_246693 + 8'h01;
  assign sel_246697 = array_index_246692 == array_index_239312 ? add_246696 : sel_246693;
  assign add_246700 = sel_246697 + 8'h01;
  assign sel_246701 = array_index_246692 == array_index_239316 ? add_246700 : sel_246697;
  assign add_246704 = sel_246701 + 8'h01;
  assign sel_246705 = array_index_246692 == array_index_239324 ? add_246704 : sel_246701;
  assign add_246708 = sel_246705 + 8'h01;
  assign sel_246709 = array_index_246692 == array_index_239332 ? add_246708 : sel_246705;
  assign add_246712 = sel_246709 + 8'h01;
  assign sel_246713 = array_index_246692 == array_index_239340 ? add_246712 : sel_246709;
  assign add_246716 = sel_246713 + 8'h01;
  assign sel_246717 = array_index_246692 == array_index_239348 ? add_246716 : sel_246713;
  assign add_246720 = sel_246717 + 8'h01;
  assign sel_246721 = array_index_246692 == array_index_239356 ? add_246720 : sel_246717;
  assign add_246724 = sel_246721 + 8'h01;
  assign sel_246725 = array_index_246692 == array_index_239364 ? add_246724 : sel_246721;
  assign add_246728 = sel_246725 + 8'h01;
  assign sel_246729 = array_index_246692 == array_index_239370 ? add_246728 : sel_246725;
  assign add_246732 = sel_246729 + 8'h01;
  assign sel_246733 = array_index_246692 == array_index_239376 ? add_246732 : sel_246729;
  assign add_246736 = sel_246733 + 8'h01;
  assign sel_246737 = array_index_246692 == array_index_239382 ? add_246736 : sel_246733;
  assign add_246740 = sel_246737 + 8'h01;
  assign sel_246741 = array_index_246692 == array_index_239388 ? add_246740 : sel_246737;
  assign add_246744 = sel_246741 + 8'h01;
  assign sel_246745 = array_index_246692 == array_index_239394 ? add_246744 : sel_246741;
  assign add_246748 = sel_246745 + 8'h01;
  assign sel_246749 = array_index_246692 == array_index_239400 ? add_246748 : sel_246745;
  assign add_246752 = sel_246749 + 8'h01;
  assign sel_246753 = array_index_246692 == array_index_239406 ? add_246752 : sel_246749;
  assign add_246756 = sel_246753 + 8'h01;
  assign sel_246757 = array_index_246692 == array_index_239412 ? add_246756 : sel_246753;
  assign add_246760 = sel_246757 + 8'h01;
  assign sel_246761 = array_index_246692 == array_index_239418 ? add_246760 : sel_246757;
  assign add_246764 = sel_246761 + 8'h01;
  assign sel_246765 = array_index_246692 == array_index_239424 ? add_246764 : sel_246761;
  assign add_246768 = sel_246765 + 8'h01;
  assign sel_246769 = array_index_246692 == array_index_239430 ? add_246768 : sel_246765;
  assign add_246772 = sel_246769 + 8'h01;
  assign sel_246773 = array_index_246692 == array_index_239436 ? add_246772 : sel_246769;
  assign add_246776 = sel_246773 + 8'h01;
  assign sel_246777 = array_index_246692 == array_index_239442 ? add_246776 : sel_246773;
  assign add_246780 = sel_246777 + 8'h01;
  assign sel_246781 = array_index_246692 == array_index_239448 ? add_246780 : sel_246777;
  assign add_246784 = sel_246781 + 8'h01;
  assign sel_246785 = array_index_246692 == array_index_239454 ? add_246784 : sel_246781;
  assign add_246788 = sel_246785 + 8'h01;
  assign sel_246789 = array_index_246692 == array_index_239460 ? add_246788 : sel_246785;
  assign add_246792 = sel_246789 + 8'h01;
  assign sel_246793 = array_index_246692 == array_index_239466 ? add_246792 : sel_246789;
  assign add_246796 = sel_246793 + 8'h01;
  assign sel_246797 = array_index_246692 == array_index_239472 ? add_246796 : sel_246793;
  assign add_246800 = sel_246797 + 8'h01;
  assign sel_246801 = array_index_246692 == array_index_239478 ? add_246800 : sel_246797;
  assign add_246804 = sel_246801 + 8'h01;
  assign sel_246805 = array_index_246692 == array_index_239484 ? add_246804 : sel_246801;
  assign add_246808 = sel_246805 + 8'h01;
  assign sel_246809 = array_index_246692 == array_index_239490 ? add_246808 : sel_246805;
  assign add_246812 = sel_246809 + 8'h01;
  assign sel_246813 = array_index_246692 == array_index_239496 ? add_246812 : sel_246809;
  assign add_246816 = sel_246813 + 8'h01;
  assign sel_246817 = array_index_246692 == array_index_239502 ? add_246816 : sel_246813;
  assign add_246820 = sel_246817 + 8'h01;
  assign sel_246821 = array_index_246692 == array_index_239508 ? add_246820 : sel_246817;
  assign add_246824 = sel_246821 + 8'h01;
  assign sel_246825 = array_index_246692 == array_index_239514 ? add_246824 : sel_246821;
  assign add_246828 = sel_246825 + 8'h01;
  assign sel_246829 = array_index_246692 == array_index_239520 ? add_246828 : sel_246825;
  assign add_246832 = sel_246829 + 8'h01;
  assign sel_246833 = array_index_246692 == array_index_239526 ? add_246832 : sel_246829;
  assign add_246836 = sel_246833 + 8'h01;
  assign sel_246837 = array_index_246692 == array_index_239532 ? add_246836 : sel_246833;
  assign add_246840 = sel_246837 + 8'h01;
  assign sel_246841 = array_index_246692 == array_index_239538 ? add_246840 : sel_246837;
  assign add_246844 = sel_246841 + 8'h01;
  assign sel_246845 = array_index_246692 == array_index_239544 ? add_246844 : sel_246841;
  assign add_246848 = sel_246845 + 8'h01;
  assign sel_246849 = array_index_246692 == array_index_239550 ? add_246848 : sel_246845;
  assign add_246852 = sel_246849 + 8'h01;
  assign sel_246853 = array_index_246692 == array_index_239556 ? add_246852 : sel_246849;
  assign add_246856 = sel_246853 + 8'h01;
  assign sel_246857 = array_index_246692 == array_index_239562 ? add_246856 : sel_246853;
  assign add_246860 = sel_246857 + 8'h01;
  assign sel_246861 = array_index_246692 == array_index_239568 ? add_246860 : sel_246857;
  assign add_246864 = sel_246861 + 8'h01;
  assign sel_246865 = array_index_246692 == array_index_239574 ? add_246864 : sel_246861;
  assign add_246868 = sel_246865 + 8'h01;
  assign sel_246869 = array_index_246692 == array_index_239580 ? add_246868 : sel_246865;
  assign add_246872 = sel_246869 + 8'h01;
  assign sel_246873 = array_index_246692 == array_index_239586 ? add_246872 : sel_246869;
  assign add_246876 = sel_246873 + 8'h01;
  assign sel_246877 = array_index_246692 == array_index_239592 ? add_246876 : sel_246873;
  assign add_246880 = sel_246877 + 8'h01;
  assign sel_246881 = array_index_246692 == array_index_239598 ? add_246880 : sel_246877;
  assign add_246884 = sel_246881 + 8'h01;
  assign sel_246885 = array_index_246692 == array_index_239604 ? add_246884 : sel_246881;
  assign add_246888 = sel_246885 + 8'h01;
  assign sel_246889 = array_index_246692 == array_index_239610 ? add_246888 : sel_246885;
  assign add_246893 = sel_246889 + 8'h01;
  assign array_index_246894 = set1_unflattened[6'h25];
  assign sel_246895 = array_index_246692 == array_index_239616 ? add_246893 : sel_246889;
  assign add_246898 = sel_246895 + 8'h01;
  assign sel_246899 = array_index_246894 == array_index_239312 ? add_246898 : sel_246895;
  assign add_246902 = sel_246899 + 8'h01;
  assign sel_246903 = array_index_246894 == array_index_239316 ? add_246902 : sel_246899;
  assign add_246906 = sel_246903 + 8'h01;
  assign sel_246907 = array_index_246894 == array_index_239324 ? add_246906 : sel_246903;
  assign add_246910 = sel_246907 + 8'h01;
  assign sel_246911 = array_index_246894 == array_index_239332 ? add_246910 : sel_246907;
  assign add_246914 = sel_246911 + 8'h01;
  assign sel_246915 = array_index_246894 == array_index_239340 ? add_246914 : sel_246911;
  assign add_246918 = sel_246915 + 8'h01;
  assign sel_246919 = array_index_246894 == array_index_239348 ? add_246918 : sel_246915;
  assign add_246922 = sel_246919 + 8'h01;
  assign sel_246923 = array_index_246894 == array_index_239356 ? add_246922 : sel_246919;
  assign add_246926 = sel_246923 + 8'h01;
  assign sel_246927 = array_index_246894 == array_index_239364 ? add_246926 : sel_246923;
  assign add_246930 = sel_246927 + 8'h01;
  assign sel_246931 = array_index_246894 == array_index_239370 ? add_246930 : sel_246927;
  assign add_246934 = sel_246931 + 8'h01;
  assign sel_246935 = array_index_246894 == array_index_239376 ? add_246934 : sel_246931;
  assign add_246938 = sel_246935 + 8'h01;
  assign sel_246939 = array_index_246894 == array_index_239382 ? add_246938 : sel_246935;
  assign add_246942 = sel_246939 + 8'h01;
  assign sel_246943 = array_index_246894 == array_index_239388 ? add_246942 : sel_246939;
  assign add_246946 = sel_246943 + 8'h01;
  assign sel_246947 = array_index_246894 == array_index_239394 ? add_246946 : sel_246943;
  assign add_246950 = sel_246947 + 8'h01;
  assign sel_246951 = array_index_246894 == array_index_239400 ? add_246950 : sel_246947;
  assign add_246954 = sel_246951 + 8'h01;
  assign sel_246955 = array_index_246894 == array_index_239406 ? add_246954 : sel_246951;
  assign add_246958 = sel_246955 + 8'h01;
  assign sel_246959 = array_index_246894 == array_index_239412 ? add_246958 : sel_246955;
  assign add_246962 = sel_246959 + 8'h01;
  assign sel_246963 = array_index_246894 == array_index_239418 ? add_246962 : sel_246959;
  assign add_246966 = sel_246963 + 8'h01;
  assign sel_246967 = array_index_246894 == array_index_239424 ? add_246966 : sel_246963;
  assign add_246970 = sel_246967 + 8'h01;
  assign sel_246971 = array_index_246894 == array_index_239430 ? add_246970 : sel_246967;
  assign add_246974 = sel_246971 + 8'h01;
  assign sel_246975 = array_index_246894 == array_index_239436 ? add_246974 : sel_246971;
  assign add_246978 = sel_246975 + 8'h01;
  assign sel_246979 = array_index_246894 == array_index_239442 ? add_246978 : sel_246975;
  assign add_246982 = sel_246979 + 8'h01;
  assign sel_246983 = array_index_246894 == array_index_239448 ? add_246982 : sel_246979;
  assign add_246986 = sel_246983 + 8'h01;
  assign sel_246987 = array_index_246894 == array_index_239454 ? add_246986 : sel_246983;
  assign add_246990 = sel_246987 + 8'h01;
  assign sel_246991 = array_index_246894 == array_index_239460 ? add_246990 : sel_246987;
  assign add_246994 = sel_246991 + 8'h01;
  assign sel_246995 = array_index_246894 == array_index_239466 ? add_246994 : sel_246991;
  assign add_246998 = sel_246995 + 8'h01;
  assign sel_246999 = array_index_246894 == array_index_239472 ? add_246998 : sel_246995;
  assign add_247002 = sel_246999 + 8'h01;
  assign sel_247003 = array_index_246894 == array_index_239478 ? add_247002 : sel_246999;
  assign add_247006 = sel_247003 + 8'h01;
  assign sel_247007 = array_index_246894 == array_index_239484 ? add_247006 : sel_247003;
  assign add_247010 = sel_247007 + 8'h01;
  assign sel_247011 = array_index_246894 == array_index_239490 ? add_247010 : sel_247007;
  assign add_247014 = sel_247011 + 8'h01;
  assign sel_247015 = array_index_246894 == array_index_239496 ? add_247014 : sel_247011;
  assign add_247018 = sel_247015 + 8'h01;
  assign sel_247019 = array_index_246894 == array_index_239502 ? add_247018 : sel_247015;
  assign add_247022 = sel_247019 + 8'h01;
  assign sel_247023 = array_index_246894 == array_index_239508 ? add_247022 : sel_247019;
  assign add_247026 = sel_247023 + 8'h01;
  assign sel_247027 = array_index_246894 == array_index_239514 ? add_247026 : sel_247023;
  assign add_247030 = sel_247027 + 8'h01;
  assign sel_247031 = array_index_246894 == array_index_239520 ? add_247030 : sel_247027;
  assign add_247034 = sel_247031 + 8'h01;
  assign sel_247035 = array_index_246894 == array_index_239526 ? add_247034 : sel_247031;
  assign add_247038 = sel_247035 + 8'h01;
  assign sel_247039 = array_index_246894 == array_index_239532 ? add_247038 : sel_247035;
  assign add_247042 = sel_247039 + 8'h01;
  assign sel_247043 = array_index_246894 == array_index_239538 ? add_247042 : sel_247039;
  assign add_247046 = sel_247043 + 8'h01;
  assign sel_247047 = array_index_246894 == array_index_239544 ? add_247046 : sel_247043;
  assign add_247050 = sel_247047 + 8'h01;
  assign sel_247051 = array_index_246894 == array_index_239550 ? add_247050 : sel_247047;
  assign add_247054 = sel_247051 + 8'h01;
  assign sel_247055 = array_index_246894 == array_index_239556 ? add_247054 : sel_247051;
  assign add_247058 = sel_247055 + 8'h01;
  assign sel_247059 = array_index_246894 == array_index_239562 ? add_247058 : sel_247055;
  assign add_247062 = sel_247059 + 8'h01;
  assign sel_247063 = array_index_246894 == array_index_239568 ? add_247062 : sel_247059;
  assign add_247066 = sel_247063 + 8'h01;
  assign sel_247067 = array_index_246894 == array_index_239574 ? add_247066 : sel_247063;
  assign add_247070 = sel_247067 + 8'h01;
  assign sel_247071 = array_index_246894 == array_index_239580 ? add_247070 : sel_247067;
  assign add_247074 = sel_247071 + 8'h01;
  assign sel_247075 = array_index_246894 == array_index_239586 ? add_247074 : sel_247071;
  assign add_247078 = sel_247075 + 8'h01;
  assign sel_247079 = array_index_246894 == array_index_239592 ? add_247078 : sel_247075;
  assign add_247082 = sel_247079 + 8'h01;
  assign sel_247083 = array_index_246894 == array_index_239598 ? add_247082 : sel_247079;
  assign add_247086 = sel_247083 + 8'h01;
  assign sel_247087 = array_index_246894 == array_index_239604 ? add_247086 : sel_247083;
  assign add_247090 = sel_247087 + 8'h01;
  assign sel_247091 = array_index_246894 == array_index_239610 ? add_247090 : sel_247087;
  assign add_247095 = sel_247091 + 8'h01;
  assign array_index_247096 = set1_unflattened[6'h26];
  assign sel_247097 = array_index_246894 == array_index_239616 ? add_247095 : sel_247091;
  assign add_247100 = sel_247097 + 8'h01;
  assign sel_247101 = array_index_247096 == array_index_239312 ? add_247100 : sel_247097;
  assign add_247104 = sel_247101 + 8'h01;
  assign sel_247105 = array_index_247096 == array_index_239316 ? add_247104 : sel_247101;
  assign add_247108 = sel_247105 + 8'h01;
  assign sel_247109 = array_index_247096 == array_index_239324 ? add_247108 : sel_247105;
  assign add_247112 = sel_247109 + 8'h01;
  assign sel_247113 = array_index_247096 == array_index_239332 ? add_247112 : sel_247109;
  assign add_247116 = sel_247113 + 8'h01;
  assign sel_247117 = array_index_247096 == array_index_239340 ? add_247116 : sel_247113;
  assign add_247120 = sel_247117 + 8'h01;
  assign sel_247121 = array_index_247096 == array_index_239348 ? add_247120 : sel_247117;
  assign add_247124 = sel_247121 + 8'h01;
  assign sel_247125 = array_index_247096 == array_index_239356 ? add_247124 : sel_247121;
  assign add_247128 = sel_247125 + 8'h01;
  assign sel_247129 = array_index_247096 == array_index_239364 ? add_247128 : sel_247125;
  assign add_247132 = sel_247129 + 8'h01;
  assign sel_247133 = array_index_247096 == array_index_239370 ? add_247132 : sel_247129;
  assign add_247136 = sel_247133 + 8'h01;
  assign sel_247137 = array_index_247096 == array_index_239376 ? add_247136 : sel_247133;
  assign add_247140 = sel_247137 + 8'h01;
  assign sel_247141 = array_index_247096 == array_index_239382 ? add_247140 : sel_247137;
  assign add_247144 = sel_247141 + 8'h01;
  assign sel_247145 = array_index_247096 == array_index_239388 ? add_247144 : sel_247141;
  assign add_247148 = sel_247145 + 8'h01;
  assign sel_247149 = array_index_247096 == array_index_239394 ? add_247148 : sel_247145;
  assign add_247152 = sel_247149 + 8'h01;
  assign sel_247153 = array_index_247096 == array_index_239400 ? add_247152 : sel_247149;
  assign add_247156 = sel_247153 + 8'h01;
  assign sel_247157 = array_index_247096 == array_index_239406 ? add_247156 : sel_247153;
  assign add_247160 = sel_247157 + 8'h01;
  assign sel_247161 = array_index_247096 == array_index_239412 ? add_247160 : sel_247157;
  assign add_247164 = sel_247161 + 8'h01;
  assign sel_247165 = array_index_247096 == array_index_239418 ? add_247164 : sel_247161;
  assign add_247168 = sel_247165 + 8'h01;
  assign sel_247169 = array_index_247096 == array_index_239424 ? add_247168 : sel_247165;
  assign add_247172 = sel_247169 + 8'h01;
  assign sel_247173 = array_index_247096 == array_index_239430 ? add_247172 : sel_247169;
  assign add_247176 = sel_247173 + 8'h01;
  assign sel_247177 = array_index_247096 == array_index_239436 ? add_247176 : sel_247173;
  assign add_247180 = sel_247177 + 8'h01;
  assign sel_247181 = array_index_247096 == array_index_239442 ? add_247180 : sel_247177;
  assign add_247184 = sel_247181 + 8'h01;
  assign sel_247185 = array_index_247096 == array_index_239448 ? add_247184 : sel_247181;
  assign add_247188 = sel_247185 + 8'h01;
  assign sel_247189 = array_index_247096 == array_index_239454 ? add_247188 : sel_247185;
  assign add_247192 = sel_247189 + 8'h01;
  assign sel_247193 = array_index_247096 == array_index_239460 ? add_247192 : sel_247189;
  assign add_247196 = sel_247193 + 8'h01;
  assign sel_247197 = array_index_247096 == array_index_239466 ? add_247196 : sel_247193;
  assign add_247200 = sel_247197 + 8'h01;
  assign sel_247201 = array_index_247096 == array_index_239472 ? add_247200 : sel_247197;
  assign add_247204 = sel_247201 + 8'h01;
  assign sel_247205 = array_index_247096 == array_index_239478 ? add_247204 : sel_247201;
  assign add_247208 = sel_247205 + 8'h01;
  assign sel_247209 = array_index_247096 == array_index_239484 ? add_247208 : sel_247205;
  assign add_247212 = sel_247209 + 8'h01;
  assign sel_247213 = array_index_247096 == array_index_239490 ? add_247212 : sel_247209;
  assign add_247216 = sel_247213 + 8'h01;
  assign sel_247217 = array_index_247096 == array_index_239496 ? add_247216 : sel_247213;
  assign add_247220 = sel_247217 + 8'h01;
  assign sel_247221 = array_index_247096 == array_index_239502 ? add_247220 : sel_247217;
  assign add_247224 = sel_247221 + 8'h01;
  assign sel_247225 = array_index_247096 == array_index_239508 ? add_247224 : sel_247221;
  assign add_247228 = sel_247225 + 8'h01;
  assign sel_247229 = array_index_247096 == array_index_239514 ? add_247228 : sel_247225;
  assign add_247232 = sel_247229 + 8'h01;
  assign sel_247233 = array_index_247096 == array_index_239520 ? add_247232 : sel_247229;
  assign add_247236 = sel_247233 + 8'h01;
  assign sel_247237 = array_index_247096 == array_index_239526 ? add_247236 : sel_247233;
  assign add_247240 = sel_247237 + 8'h01;
  assign sel_247241 = array_index_247096 == array_index_239532 ? add_247240 : sel_247237;
  assign add_247244 = sel_247241 + 8'h01;
  assign sel_247245 = array_index_247096 == array_index_239538 ? add_247244 : sel_247241;
  assign add_247248 = sel_247245 + 8'h01;
  assign sel_247249 = array_index_247096 == array_index_239544 ? add_247248 : sel_247245;
  assign add_247252 = sel_247249 + 8'h01;
  assign sel_247253 = array_index_247096 == array_index_239550 ? add_247252 : sel_247249;
  assign add_247256 = sel_247253 + 8'h01;
  assign sel_247257 = array_index_247096 == array_index_239556 ? add_247256 : sel_247253;
  assign add_247260 = sel_247257 + 8'h01;
  assign sel_247261 = array_index_247096 == array_index_239562 ? add_247260 : sel_247257;
  assign add_247264 = sel_247261 + 8'h01;
  assign sel_247265 = array_index_247096 == array_index_239568 ? add_247264 : sel_247261;
  assign add_247268 = sel_247265 + 8'h01;
  assign sel_247269 = array_index_247096 == array_index_239574 ? add_247268 : sel_247265;
  assign add_247272 = sel_247269 + 8'h01;
  assign sel_247273 = array_index_247096 == array_index_239580 ? add_247272 : sel_247269;
  assign add_247276 = sel_247273 + 8'h01;
  assign sel_247277 = array_index_247096 == array_index_239586 ? add_247276 : sel_247273;
  assign add_247280 = sel_247277 + 8'h01;
  assign sel_247281 = array_index_247096 == array_index_239592 ? add_247280 : sel_247277;
  assign add_247284 = sel_247281 + 8'h01;
  assign sel_247285 = array_index_247096 == array_index_239598 ? add_247284 : sel_247281;
  assign add_247288 = sel_247285 + 8'h01;
  assign sel_247289 = array_index_247096 == array_index_239604 ? add_247288 : sel_247285;
  assign add_247292 = sel_247289 + 8'h01;
  assign sel_247293 = array_index_247096 == array_index_239610 ? add_247292 : sel_247289;
  assign add_247297 = sel_247293 + 8'h01;
  assign array_index_247298 = set1_unflattened[6'h27];
  assign sel_247299 = array_index_247096 == array_index_239616 ? add_247297 : sel_247293;
  assign add_247302 = sel_247299 + 8'h01;
  assign sel_247303 = array_index_247298 == array_index_239312 ? add_247302 : sel_247299;
  assign add_247306 = sel_247303 + 8'h01;
  assign sel_247307 = array_index_247298 == array_index_239316 ? add_247306 : sel_247303;
  assign add_247310 = sel_247307 + 8'h01;
  assign sel_247311 = array_index_247298 == array_index_239324 ? add_247310 : sel_247307;
  assign add_247314 = sel_247311 + 8'h01;
  assign sel_247315 = array_index_247298 == array_index_239332 ? add_247314 : sel_247311;
  assign add_247318 = sel_247315 + 8'h01;
  assign sel_247319 = array_index_247298 == array_index_239340 ? add_247318 : sel_247315;
  assign add_247322 = sel_247319 + 8'h01;
  assign sel_247323 = array_index_247298 == array_index_239348 ? add_247322 : sel_247319;
  assign add_247326 = sel_247323 + 8'h01;
  assign sel_247327 = array_index_247298 == array_index_239356 ? add_247326 : sel_247323;
  assign add_247330 = sel_247327 + 8'h01;
  assign sel_247331 = array_index_247298 == array_index_239364 ? add_247330 : sel_247327;
  assign add_247334 = sel_247331 + 8'h01;
  assign sel_247335 = array_index_247298 == array_index_239370 ? add_247334 : sel_247331;
  assign add_247338 = sel_247335 + 8'h01;
  assign sel_247339 = array_index_247298 == array_index_239376 ? add_247338 : sel_247335;
  assign add_247342 = sel_247339 + 8'h01;
  assign sel_247343 = array_index_247298 == array_index_239382 ? add_247342 : sel_247339;
  assign add_247346 = sel_247343 + 8'h01;
  assign sel_247347 = array_index_247298 == array_index_239388 ? add_247346 : sel_247343;
  assign add_247350 = sel_247347 + 8'h01;
  assign sel_247351 = array_index_247298 == array_index_239394 ? add_247350 : sel_247347;
  assign add_247354 = sel_247351 + 8'h01;
  assign sel_247355 = array_index_247298 == array_index_239400 ? add_247354 : sel_247351;
  assign add_247358 = sel_247355 + 8'h01;
  assign sel_247359 = array_index_247298 == array_index_239406 ? add_247358 : sel_247355;
  assign add_247362 = sel_247359 + 8'h01;
  assign sel_247363 = array_index_247298 == array_index_239412 ? add_247362 : sel_247359;
  assign add_247366 = sel_247363 + 8'h01;
  assign sel_247367 = array_index_247298 == array_index_239418 ? add_247366 : sel_247363;
  assign add_247370 = sel_247367 + 8'h01;
  assign sel_247371 = array_index_247298 == array_index_239424 ? add_247370 : sel_247367;
  assign add_247374 = sel_247371 + 8'h01;
  assign sel_247375 = array_index_247298 == array_index_239430 ? add_247374 : sel_247371;
  assign add_247378 = sel_247375 + 8'h01;
  assign sel_247379 = array_index_247298 == array_index_239436 ? add_247378 : sel_247375;
  assign add_247382 = sel_247379 + 8'h01;
  assign sel_247383 = array_index_247298 == array_index_239442 ? add_247382 : sel_247379;
  assign add_247386 = sel_247383 + 8'h01;
  assign sel_247387 = array_index_247298 == array_index_239448 ? add_247386 : sel_247383;
  assign add_247390 = sel_247387 + 8'h01;
  assign sel_247391 = array_index_247298 == array_index_239454 ? add_247390 : sel_247387;
  assign add_247394 = sel_247391 + 8'h01;
  assign sel_247395 = array_index_247298 == array_index_239460 ? add_247394 : sel_247391;
  assign add_247398 = sel_247395 + 8'h01;
  assign sel_247399 = array_index_247298 == array_index_239466 ? add_247398 : sel_247395;
  assign add_247402 = sel_247399 + 8'h01;
  assign sel_247403 = array_index_247298 == array_index_239472 ? add_247402 : sel_247399;
  assign add_247406 = sel_247403 + 8'h01;
  assign sel_247407 = array_index_247298 == array_index_239478 ? add_247406 : sel_247403;
  assign add_247410 = sel_247407 + 8'h01;
  assign sel_247411 = array_index_247298 == array_index_239484 ? add_247410 : sel_247407;
  assign add_247414 = sel_247411 + 8'h01;
  assign sel_247415 = array_index_247298 == array_index_239490 ? add_247414 : sel_247411;
  assign add_247418 = sel_247415 + 8'h01;
  assign sel_247419 = array_index_247298 == array_index_239496 ? add_247418 : sel_247415;
  assign add_247422 = sel_247419 + 8'h01;
  assign sel_247423 = array_index_247298 == array_index_239502 ? add_247422 : sel_247419;
  assign add_247426 = sel_247423 + 8'h01;
  assign sel_247427 = array_index_247298 == array_index_239508 ? add_247426 : sel_247423;
  assign add_247430 = sel_247427 + 8'h01;
  assign sel_247431 = array_index_247298 == array_index_239514 ? add_247430 : sel_247427;
  assign add_247434 = sel_247431 + 8'h01;
  assign sel_247435 = array_index_247298 == array_index_239520 ? add_247434 : sel_247431;
  assign add_247438 = sel_247435 + 8'h01;
  assign sel_247439 = array_index_247298 == array_index_239526 ? add_247438 : sel_247435;
  assign add_247442 = sel_247439 + 8'h01;
  assign sel_247443 = array_index_247298 == array_index_239532 ? add_247442 : sel_247439;
  assign add_247446 = sel_247443 + 8'h01;
  assign sel_247447 = array_index_247298 == array_index_239538 ? add_247446 : sel_247443;
  assign add_247450 = sel_247447 + 8'h01;
  assign sel_247451 = array_index_247298 == array_index_239544 ? add_247450 : sel_247447;
  assign add_247454 = sel_247451 + 8'h01;
  assign sel_247455 = array_index_247298 == array_index_239550 ? add_247454 : sel_247451;
  assign add_247458 = sel_247455 + 8'h01;
  assign sel_247459 = array_index_247298 == array_index_239556 ? add_247458 : sel_247455;
  assign add_247462 = sel_247459 + 8'h01;
  assign sel_247463 = array_index_247298 == array_index_239562 ? add_247462 : sel_247459;
  assign add_247466 = sel_247463 + 8'h01;
  assign sel_247467 = array_index_247298 == array_index_239568 ? add_247466 : sel_247463;
  assign add_247470 = sel_247467 + 8'h01;
  assign sel_247471 = array_index_247298 == array_index_239574 ? add_247470 : sel_247467;
  assign add_247474 = sel_247471 + 8'h01;
  assign sel_247475 = array_index_247298 == array_index_239580 ? add_247474 : sel_247471;
  assign add_247478 = sel_247475 + 8'h01;
  assign sel_247479 = array_index_247298 == array_index_239586 ? add_247478 : sel_247475;
  assign add_247482 = sel_247479 + 8'h01;
  assign sel_247483 = array_index_247298 == array_index_239592 ? add_247482 : sel_247479;
  assign add_247486 = sel_247483 + 8'h01;
  assign sel_247487 = array_index_247298 == array_index_239598 ? add_247486 : sel_247483;
  assign add_247490 = sel_247487 + 8'h01;
  assign sel_247491 = array_index_247298 == array_index_239604 ? add_247490 : sel_247487;
  assign add_247494 = sel_247491 + 8'h01;
  assign sel_247495 = array_index_247298 == array_index_239610 ? add_247494 : sel_247491;
  assign add_247499 = sel_247495 + 8'h01;
  assign array_index_247500 = set1_unflattened[6'h28];
  assign sel_247501 = array_index_247298 == array_index_239616 ? add_247499 : sel_247495;
  assign add_247504 = sel_247501 + 8'h01;
  assign sel_247505 = array_index_247500 == array_index_239312 ? add_247504 : sel_247501;
  assign add_247508 = sel_247505 + 8'h01;
  assign sel_247509 = array_index_247500 == array_index_239316 ? add_247508 : sel_247505;
  assign add_247512 = sel_247509 + 8'h01;
  assign sel_247513 = array_index_247500 == array_index_239324 ? add_247512 : sel_247509;
  assign add_247516 = sel_247513 + 8'h01;
  assign sel_247517 = array_index_247500 == array_index_239332 ? add_247516 : sel_247513;
  assign add_247520 = sel_247517 + 8'h01;
  assign sel_247521 = array_index_247500 == array_index_239340 ? add_247520 : sel_247517;
  assign add_247524 = sel_247521 + 8'h01;
  assign sel_247525 = array_index_247500 == array_index_239348 ? add_247524 : sel_247521;
  assign add_247528 = sel_247525 + 8'h01;
  assign sel_247529 = array_index_247500 == array_index_239356 ? add_247528 : sel_247525;
  assign add_247532 = sel_247529 + 8'h01;
  assign sel_247533 = array_index_247500 == array_index_239364 ? add_247532 : sel_247529;
  assign add_247536 = sel_247533 + 8'h01;
  assign sel_247537 = array_index_247500 == array_index_239370 ? add_247536 : sel_247533;
  assign add_247540 = sel_247537 + 8'h01;
  assign sel_247541 = array_index_247500 == array_index_239376 ? add_247540 : sel_247537;
  assign add_247544 = sel_247541 + 8'h01;
  assign sel_247545 = array_index_247500 == array_index_239382 ? add_247544 : sel_247541;
  assign add_247548 = sel_247545 + 8'h01;
  assign sel_247549 = array_index_247500 == array_index_239388 ? add_247548 : sel_247545;
  assign add_247552 = sel_247549 + 8'h01;
  assign sel_247553 = array_index_247500 == array_index_239394 ? add_247552 : sel_247549;
  assign add_247556 = sel_247553 + 8'h01;
  assign sel_247557 = array_index_247500 == array_index_239400 ? add_247556 : sel_247553;
  assign add_247560 = sel_247557 + 8'h01;
  assign sel_247561 = array_index_247500 == array_index_239406 ? add_247560 : sel_247557;
  assign add_247564 = sel_247561 + 8'h01;
  assign sel_247565 = array_index_247500 == array_index_239412 ? add_247564 : sel_247561;
  assign add_247568 = sel_247565 + 8'h01;
  assign sel_247569 = array_index_247500 == array_index_239418 ? add_247568 : sel_247565;
  assign add_247572 = sel_247569 + 8'h01;
  assign sel_247573 = array_index_247500 == array_index_239424 ? add_247572 : sel_247569;
  assign add_247576 = sel_247573 + 8'h01;
  assign sel_247577 = array_index_247500 == array_index_239430 ? add_247576 : sel_247573;
  assign add_247580 = sel_247577 + 8'h01;
  assign sel_247581 = array_index_247500 == array_index_239436 ? add_247580 : sel_247577;
  assign add_247584 = sel_247581 + 8'h01;
  assign sel_247585 = array_index_247500 == array_index_239442 ? add_247584 : sel_247581;
  assign add_247588 = sel_247585 + 8'h01;
  assign sel_247589 = array_index_247500 == array_index_239448 ? add_247588 : sel_247585;
  assign add_247592 = sel_247589 + 8'h01;
  assign sel_247593 = array_index_247500 == array_index_239454 ? add_247592 : sel_247589;
  assign add_247596 = sel_247593 + 8'h01;
  assign sel_247597 = array_index_247500 == array_index_239460 ? add_247596 : sel_247593;
  assign add_247600 = sel_247597 + 8'h01;
  assign sel_247601 = array_index_247500 == array_index_239466 ? add_247600 : sel_247597;
  assign add_247604 = sel_247601 + 8'h01;
  assign sel_247605 = array_index_247500 == array_index_239472 ? add_247604 : sel_247601;
  assign add_247608 = sel_247605 + 8'h01;
  assign sel_247609 = array_index_247500 == array_index_239478 ? add_247608 : sel_247605;
  assign add_247612 = sel_247609 + 8'h01;
  assign sel_247613 = array_index_247500 == array_index_239484 ? add_247612 : sel_247609;
  assign add_247616 = sel_247613 + 8'h01;
  assign sel_247617 = array_index_247500 == array_index_239490 ? add_247616 : sel_247613;
  assign add_247620 = sel_247617 + 8'h01;
  assign sel_247621 = array_index_247500 == array_index_239496 ? add_247620 : sel_247617;
  assign add_247624 = sel_247621 + 8'h01;
  assign sel_247625 = array_index_247500 == array_index_239502 ? add_247624 : sel_247621;
  assign add_247628 = sel_247625 + 8'h01;
  assign sel_247629 = array_index_247500 == array_index_239508 ? add_247628 : sel_247625;
  assign add_247632 = sel_247629 + 8'h01;
  assign sel_247633 = array_index_247500 == array_index_239514 ? add_247632 : sel_247629;
  assign add_247636 = sel_247633 + 8'h01;
  assign sel_247637 = array_index_247500 == array_index_239520 ? add_247636 : sel_247633;
  assign add_247640 = sel_247637 + 8'h01;
  assign sel_247641 = array_index_247500 == array_index_239526 ? add_247640 : sel_247637;
  assign add_247644 = sel_247641 + 8'h01;
  assign sel_247645 = array_index_247500 == array_index_239532 ? add_247644 : sel_247641;
  assign add_247648 = sel_247645 + 8'h01;
  assign sel_247649 = array_index_247500 == array_index_239538 ? add_247648 : sel_247645;
  assign add_247652 = sel_247649 + 8'h01;
  assign sel_247653 = array_index_247500 == array_index_239544 ? add_247652 : sel_247649;
  assign add_247656 = sel_247653 + 8'h01;
  assign sel_247657 = array_index_247500 == array_index_239550 ? add_247656 : sel_247653;
  assign add_247660 = sel_247657 + 8'h01;
  assign sel_247661 = array_index_247500 == array_index_239556 ? add_247660 : sel_247657;
  assign add_247664 = sel_247661 + 8'h01;
  assign sel_247665 = array_index_247500 == array_index_239562 ? add_247664 : sel_247661;
  assign add_247668 = sel_247665 + 8'h01;
  assign sel_247669 = array_index_247500 == array_index_239568 ? add_247668 : sel_247665;
  assign add_247672 = sel_247669 + 8'h01;
  assign sel_247673 = array_index_247500 == array_index_239574 ? add_247672 : sel_247669;
  assign add_247676 = sel_247673 + 8'h01;
  assign sel_247677 = array_index_247500 == array_index_239580 ? add_247676 : sel_247673;
  assign add_247680 = sel_247677 + 8'h01;
  assign sel_247681 = array_index_247500 == array_index_239586 ? add_247680 : sel_247677;
  assign add_247684 = sel_247681 + 8'h01;
  assign sel_247685 = array_index_247500 == array_index_239592 ? add_247684 : sel_247681;
  assign add_247688 = sel_247685 + 8'h01;
  assign sel_247689 = array_index_247500 == array_index_239598 ? add_247688 : sel_247685;
  assign add_247692 = sel_247689 + 8'h01;
  assign sel_247693 = array_index_247500 == array_index_239604 ? add_247692 : sel_247689;
  assign add_247696 = sel_247693 + 8'h01;
  assign sel_247697 = array_index_247500 == array_index_239610 ? add_247696 : sel_247693;
  assign add_247701 = sel_247697 + 8'h01;
  assign array_index_247702 = set1_unflattened[6'h29];
  assign sel_247703 = array_index_247500 == array_index_239616 ? add_247701 : sel_247697;
  assign add_247706 = sel_247703 + 8'h01;
  assign sel_247707 = array_index_247702 == array_index_239312 ? add_247706 : sel_247703;
  assign add_247710 = sel_247707 + 8'h01;
  assign sel_247711 = array_index_247702 == array_index_239316 ? add_247710 : sel_247707;
  assign add_247714 = sel_247711 + 8'h01;
  assign sel_247715 = array_index_247702 == array_index_239324 ? add_247714 : sel_247711;
  assign add_247718 = sel_247715 + 8'h01;
  assign sel_247719 = array_index_247702 == array_index_239332 ? add_247718 : sel_247715;
  assign add_247722 = sel_247719 + 8'h01;
  assign sel_247723 = array_index_247702 == array_index_239340 ? add_247722 : sel_247719;
  assign add_247726 = sel_247723 + 8'h01;
  assign sel_247727 = array_index_247702 == array_index_239348 ? add_247726 : sel_247723;
  assign add_247730 = sel_247727 + 8'h01;
  assign sel_247731 = array_index_247702 == array_index_239356 ? add_247730 : sel_247727;
  assign add_247734 = sel_247731 + 8'h01;
  assign sel_247735 = array_index_247702 == array_index_239364 ? add_247734 : sel_247731;
  assign add_247738 = sel_247735 + 8'h01;
  assign sel_247739 = array_index_247702 == array_index_239370 ? add_247738 : sel_247735;
  assign add_247742 = sel_247739 + 8'h01;
  assign sel_247743 = array_index_247702 == array_index_239376 ? add_247742 : sel_247739;
  assign add_247746 = sel_247743 + 8'h01;
  assign sel_247747 = array_index_247702 == array_index_239382 ? add_247746 : sel_247743;
  assign add_247750 = sel_247747 + 8'h01;
  assign sel_247751 = array_index_247702 == array_index_239388 ? add_247750 : sel_247747;
  assign add_247754 = sel_247751 + 8'h01;
  assign sel_247755 = array_index_247702 == array_index_239394 ? add_247754 : sel_247751;
  assign add_247758 = sel_247755 + 8'h01;
  assign sel_247759 = array_index_247702 == array_index_239400 ? add_247758 : sel_247755;
  assign add_247762 = sel_247759 + 8'h01;
  assign sel_247763 = array_index_247702 == array_index_239406 ? add_247762 : sel_247759;
  assign add_247766 = sel_247763 + 8'h01;
  assign sel_247767 = array_index_247702 == array_index_239412 ? add_247766 : sel_247763;
  assign add_247770 = sel_247767 + 8'h01;
  assign sel_247771 = array_index_247702 == array_index_239418 ? add_247770 : sel_247767;
  assign add_247774 = sel_247771 + 8'h01;
  assign sel_247775 = array_index_247702 == array_index_239424 ? add_247774 : sel_247771;
  assign add_247778 = sel_247775 + 8'h01;
  assign sel_247779 = array_index_247702 == array_index_239430 ? add_247778 : sel_247775;
  assign add_247782 = sel_247779 + 8'h01;
  assign sel_247783 = array_index_247702 == array_index_239436 ? add_247782 : sel_247779;
  assign add_247786 = sel_247783 + 8'h01;
  assign sel_247787 = array_index_247702 == array_index_239442 ? add_247786 : sel_247783;
  assign add_247790 = sel_247787 + 8'h01;
  assign sel_247791 = array_index_247702 == array_index_239448 ? add_247790 : sel_247787;
  assign add_247794 = sel_247791 + 8'h01;
  assign sel_247795 = array_index_247702 == array_index_239454 ? add_247794 : sel_247791;
  assign add_247798 = sel_247795 + 8'h01;
  assign sel_247799 = array_index_247702 == array_index_239460 ? add_247798 : sel_247795;
  assign add_247802 = sel_247799 + 8'h01;
  assign sel_247803 = array_index_247702 == array_index_239466 ? add_247802 : sel_247799;
  assign add_247806 = sel_247803 + 8'h01;
  assign sel_247807 = array_index_247702 == array_index_239472 ? add_247806 : sel_247803;
  assign add_247810 = sel_247807 + 8'h01;
  assign sel_247811 = array_index_247702 == array_index_239478 ? add_247810 : sel_247807;
  assign add_247814 = sel_247811 + 8'h01;
  assign sel_247815 = array_index_247702 == array_index_239484 ? add_247814 : sel_247811;
  assign add_247818 = sel_247815 + 8'h01;
  assign sel_247819 = array_index_247702 == array_index_239490 ? add_247818 : sel_247815;
  assign add_247822 = sel_247819 + 8'h01;
  assign sel_247823 = array_index_247702 == array_index_239496 ? add_247822 : sel_247819;
  assign add_247826 = sel_247823 + 8'h01;
  assign sel_247827 = array_index_247702 == array_index_239502 ? add_247826 : sel_247823;
  assign add_247830 = sel_247827 + 8'h01;
  assign sel_247831 = array_index_247702 == array_index_239508 ? add_247830 : sel_247827;
  assign add_247834 = sel_247831 + 8'h01;
  assign sel_247835 = array_index_247702 == array_index_239514 ? add_247834 : sel_247831;
  assign add_247838 = sel_247835 + 8'h01;
  assign sel_247839 = array_index_247702 == array_index_239520 ? add_247838 : sel_247835;
  assign add_247842 = sel_247839 + 8'h01;
  assign sel_247843 = array_index_247702 == array_index_239526 ? add_247842 : sel_247839;
  assign add_247846 = sel_247843 + 8'h01;
  assign sel_247847 = array_index_247702 == array_index_239532 ? add_247846 : sel_247843;
  assign add_247850 = sel_247847 + 8'h01;
  assign sel_247851 = array_index_247702 == array_index_239538 ? add_247850 : sel_247847;
  assign add_247854 = sel_247851 + 8'h01;
  assign sel_247855 = array_index_247702 == array_index_239544 ? add_247854 : sel_247851;
  assign add_247858 = sel_247855 + 8'h01;
  assign sel_247859 = array_index_247702 == array_index_239550 ? add_247858 : sel_247855;
  assign add_247862 = sel_247859 + 8'h01;
  assign sel_247863 = array_index_247702 == array_index_239556 ? add_247862 : sel_247859;
  assign add_247866 = sel_247863 + 8'h01;
  assign sel_247867 = array_index_247702 == array_index_239562 ? add_247866 : sel_247863;
  assign add_247870 = sel_247867 + 8'h01;
  assign sel_247871 = array_index_247702 == array_index_239568 ? add_247870 : sel_247867;
  assign add_247874 = sel_247871 + 8'h01;
  assign sel_247875 = array_index_247702 == array_index_239574 ? add_247874 : sel_247871;
  assign add_247878 = sel_247875 + 8'h01;
  assign sel_247879 = array_index_247702 == array_index_239580 ? add_247878 : sel_247875;
  assign add_247882 = sel_247879 + 8'h01;
  assign sel_247883 = array_index_247702 == array_index_239586 ? add_247882 : sel_247879;
  assign add_247886 = sel_247883 + 8'h01;
  assign sel_247887 = array_index_247702 == array_index_239592 ? add_247886 : sel_247883;
  assign add_247890 = sel_247887 + 8'h01;
  assign sel_247891 = array_index_247702 == array_index_239598 ? add_247890 : sel_247887;
  assign add_247894 = sel_247891 + 8'h01;
  assign sel_247895 = array_index_247702 == array_index_239604 ? add_247894 : sel_247891;
  assign add_247898 = sel_247895 + 8'h01;
  assign sel_247899 = array_index_247702 == array_index_239610 ? add_247898 : sel_247895;
  assign add_247903 = sel_247899 + 8'h01;
  assign array_index_247904 = set1_unflattened[6'h2a];
  assign sel_247905 = array_index_247702 == array_index_239616 ? add_247903 : sel_247899;
  assign add_247908 = sel_247905 + 8'h01;
  assign sel_247909 = array_index_247904 == array_index_239312 ? add_247908 : sel_247905;
  assign add_247912 = sel_247909 + 8'h01;
  assign sel_247913 = array_index_247904 == array_index_239316 ? add_247912 : sel_247909;
  assign add_247916 = sel_247913 + 8'h01;
  assign sel_247917 = array_index_247904 == array_index_239324 ? add_247916 : sel_247913;
  assign add_247920 = sel_247917 + 8'h01;
  assign sel_247921 = array_index_247904 == array_index_239332 ? add_247920 : sel_247917;
  assign add_247924 = sel_247921 + 8'h01;
  assign sel_247925 = array_index_247904 == array_index_239340 ? add_247924 : sel_247921;
  assign add_247928 = sel_247925 + 8'h01;
  assign sel_247929 = array_index_247904 == array_index_239348 ? add_247928 : sel_247925;
  assign add_247932 = sel_247929 + 8'h01;
  assign sel_247933 = array_index_247904 == array_index_239356 ? add_247932 : sel_247929;
  assign add_247936 = sel_247933 + 8'h01;
  assign sel_247937 = array_index_247904 == array_index_239364 ? add_247936 : sel_247933;
  assign add_247940 = sel_247937 + 8'h01;
  assign sel_247941 = array_index_247904 == array_index_239370 ? add_247940 : sel_247937;
  assign add_247944 = sel_247941 + 8'h01;
  assign sel_247945 = array_index_247904 == array_index_239376 ? add_247944 : sel_247941;
  assign add_247948 = sel_247945 + 8'h01;
  assign sel_247949 = array_index_247904 == array_index_239382 ? add_247948 : sel_247945;
  assign add_247952 = sel_247949 + 8'h01;
  assign sel_247953 = array_index_247904 == array_index_239388 ? add_247952 : sel_247949;
  assign add_247956 = sel_247953 + 8'h01;
  assign sel_247957 = array_index_247904 == array_index_239394 ? add_247956 : sel_247953;
  assign add_247960 = sel_247957 + 8'h01;
  assign sel_247961 = array_index_247904 == array_index_239400 ? add_247960 : sel_247957;
  assign add_247964 = sel_247961 + 8'h01;
  assign sel_247965 = array_index_247904 == array_index_239406 ? add_247964 : sel_247961;
  assign add_247968 = sel_247965 + 8'h01;
  assign sel_247969 = array_index_247904 == array_index_239412 ? add_247968 : sel_247965;
  assign add_247972 = sel_247969 + 8'h01;
  assign sel_247973 = array_index_247904 == array_index_239418 ? add_247972 : sel_247969;
  assign add_247976 = sel_247973 + 8'h01;
  assign sel_247977 = array_index_247904 == array_index_239424 ? add_247976 : sel_247973;
  assign add_247980 = sel_247977 + 8'h01;
  assign sel_247981 = array_index_247904 == array_index_239430 ? add_247980 : sel_247977;
  assign add_247984 = sel_247981 + 8'h01;
  assign sel_247985 = array_index_247904 == array_index_239436 ? add_247984 : sel_247981;
  assign add_247988 = sel_247985 + 8'h01;
  assign sel_247989 = array_index_247904 == array_index_239442 ? add_247988 : sel_247985;
  assign add_247992 = sel_247989 + 8'h01;
  assign sel_247993 = array_index_247904 == array_index_239448 ? add_247992 : sel_247989;
  assign add_247996 = sel_247993 + 8'h01;
  assign sel_247997 = array_index_247904 == array_index_239454 ? add_247996 : sel_247993;
  assign add_248000 = sel_247997 + 8'h01;
  assign sel_248001 = array_index_247904 == array_index_239460 ? add_248000 : sel_247997;
  assign add_248004 = sel_248001 + 8'h01;
  assign sel_248005 = array_index_247904 == array_index_239466 ? add_248004 : sel_248001;
  assign add_248008 = sel_248005 + 8'h01;
  assign sel_248009 = array_index_247904 == array_index_239472 ? add_248008 : sel_248005;
  assign add_248012 = sel_248009 + 8'h01;
  assign sel_248013 = array_index_247904 == array_index_239478 ? add_248012 : sel_248009;
  assign add_248016 = sel_248013 + 8'h01;
  assign sel_248017 = array_index_247904 == array_index_239484 ? add_248016 : sel_248013;
  assign add_248020 = sel_248017 + 8'h01;
  assign sel_248021 = array_index_247904 == array_index_239490 ? add_248020 : sel_248017;
  assign add_248024 = sel_248021 + 8'h01;
  assign sel_248025 = array_index_247904 == array_index_239496 ? add_248024 : sel_248021;
  assign add_248028 = sel_248025 + 8'h01;
  assign sel_248029 = array_index_247904 == array_index_239502 ? add_248028 : sel_248025;
  assign add_248032 = sel_248029 + 8'h01;
  assign sel_248033 = array_index_247904 == array_index_239508 ? add_248032 : sel_248029;
  assign add_248036 = sel_248033 + 8'h01;
  assign sel_248037 = array_index_247904 == array_index_239514 ? add_248036 : sel_248033;
  assign add_248040 = sel_248037 + 8'h01;
  assign sel_248041 = array_index_247904 == array_index_239520 ? add_248040 : sel_248037;
  assign add_248044 = sel_248041 + 8'h01;
  assign sel_248045 = array_index_247904 == array_index_239526 ? add_248044 : sel_248041;
  assign add_248048 = sel_248045 + 8'h01;
  assign sel_248049 = array_index_247904 == array_index_239532 ? add_248048 : sel_248045;
  assign add_248052 = sel_248049 + 8'h01;
  assign sel_248053 = array_index_247904 == array_index_239538 ? add_248052 : sel_248049;
  assign add_248056 = sel_248053 + 8'h01;
  assign sel_248057 = array_index_247904 == array_index_239544 ? add_248056 : sel_248053;
  assign add_248060 = sel_248057 + 8'h01;
  assign sel_248061 = array_index_247904 == array_index_239550 ? add_248060 : sel_248057;
  assign add_248064 = sel_248061 + 8'h01;
  assign sel_248065 = array_index_247904 == array_index_239556 ? add_248064 : sel_248061;
  assign add_248068 = sel_248065 + 8'h01;
  assign sel_248069 = array_index_247904 == array_index_239562 ? add_248068 : sel_248065;
  assign add_248072 = sel_248069 + 8'h01;
  assign sel_248073 = array_index_247904 == array_index_239568 ? add_248072 : sel_248069;
  assign add_248076 = sel_248073 + 8'h01;
  assign sel_248077 = array_index_247904 == array_index_239574 ? add_248076 : sel_248073;
  assign add_248080 = sel_248077 + 8'h01;
  assign sel_248081 = array_index_247904 == array_index_239580 ? add_248080 : sel_248077;
  assign add_248084 = sel_248081 + 8'h01;
  assign sel_248085 = array_index_247904 == array_index_239586 ? add_248084 : sel_248081;
  assign add_248088 = sel_248085 + 8'h01;
  assign sel_248089 = array_index_247904 == array_index_239592 ? add_248088 : sel_248085;
  assign add_248092 = sel_248089 + 8'h01;
  assign sel_248093 = array_index_247904 == array_index_239598 ? add_248092 : sel_248089;
  assign add_248096 = sel_248093 + 8'h01;
  assign sel_248097 = array_index_247904 == array_index_239604 ? add_248096 : sel_248093;
  assign add_248100 = sel_248097 + 8'h01;
  assign sel_248101 = array_index_247904 == array_index_239610 ? add_248100 : sel_248097;
  assign add_248105 = sel_248101 + 8'h01;
  assign array_index_248106 = set1_unflattened[6'h2b];
  assign sel_248107 = array_index_247904 == array_index_239616 ? add_248105 : sel_248101;
  assign add_248110 = sel_248107 + 8'h01;
  assign sel_248111 = array_index_248106 == array_index_239312 ? add_248110 : sel_248107;
  assign add_248114 = sel_248111 + 8'h01;
  assign sel_248115 = array_index_248106 == array_index_239316 ? add_248114 : sel_248111;
  assign add_248118 = sel_248115 + 8'h01;
  assign sel_248119 = array_index_248106 == array_index_239324 ? add_248118 : sel_248115;
  assign add_248122 = sel_248119 + 8'h01;
  assign sel_248123 = array_index_248106 == array_index_239332 ? add_248122 : sel_248119;
  assign add_248126 = sel_248123 + 8'h01;
  assign sel_248127 = array_index_248106 == array_index_239340 ? add_248126 : sel_248123;
  assign add_248130 = sel_248127 + 8'h01;
  assign sel_248131 = array_index_248106 == array_index_239348 ? add_248130 : sel_248127;
  assign add_248134 = sel_248131 + 8'h01;
  assign sel_248135 = array_index_248106 == array_index_239356 ? add_248134 : sel_248131;
  assign add_248138 = sel_248135 + 8'h01;
  assign sel_248139 = array_index_248106 == array_index_239364 ? add_248138 : sel_248135;
  assign add_248142 = sel_248139 + 8'h01;
  assign sel_248143 = array_index_248106 == array_index_239370 ? add_248142 : sel_248139;
  assign add_248146 = sel_248143 + 8'h01;
  assign sel_248147 = array_index_248106 == array_index_239376 ? add_248146 : sel_248143;
  assign add_248150 = sel_248147 + 8'h01;
  assign sel_248151 = array_index_248106 == array_index_239382 ? add_248150 : sel_248147;
  assign add_248154 = sel_248151 + 8'h01;
  assign sel_248155 = array_index_248106 == array_index_239388 ? add_248154 : sel_248151;
  assign add_248158 = sel_248155 + 8'h01;
  assign sel_248159 = array_index_248106 == array_index_239394 ? add_248158 : sel_248155;
  assign add_248162 = sel_248159 + 8'h01;
  assign sel_248163 = array_index_248106 == array_index_239400 ? add_248162 : sel_248159;
  assign add_248166 = sel_248163 + 8'h01;
  assign sel_248167 = array_index_248106 == array_index_239406 ? add_248166 : sel_248163;
  assign add_248170 = sel_248167 + 8'h01;
  assign sel_248171 = array_index_248106 == array_index_239412 ? add_248170 : sel_248167;
  assign add_248174 = sel_248171 + 8'h01;
  assign sel_248175 = array_index_248106 == array_index_239418 ? add_248174 : sel_248171;
  assign add_248178 = sel_248175 + 8'h01;
  assign sel_248179 = array_index_248106 == array_index_239424 ? add_248178 : sel_248175;
  assign add_248182 = sel_248179 + 8'h01;
  assign sel_248183 = array_index_248106 == array_index_239430 ? add_248182 : sel_248179;
  assign add_248186 = sel_248183 + 8'h01;
  assign sel_248187 = array_index_248106 == array_index_239436 ? add_248186 : sel_248183;
  assign add_248190 = sel_248187 + 8'h01;
  assign sel_248191 = array_index_248106 == array_index_239442 ? add_248190 : sel_248187;
  assign add_248194 = sel_248191 + 8'h01;
  assign sel_248195 = array_index_248106 == array_index_239448 ? add_248194 : sel_248191;
  assign add_248198 = sel_248195 + 8'h01;
  assign sel_248199 = array_index_248106 == array_index_239454 ? add_248198 : sel_248195;
  assign add_248202 = sel_248199 + 8'h01;
  assign sel_248203 = array_index_248106 == array_index_239460 ? add_248202 : sel_248199;
  assign add_248206 = sel_248203 + 8'h01;
  assign sel_248207 = array_index_248106 == array_index_239466 ? add_248206 : sel_248203;
  assign add_248210 = sel_248207 + 8'h01;
  assign sel_248211 = array_index_248106 == array_index_239472 ? add_248210 : sel_248207;
  assign add_248214 = sel_248211 + 8'h01;
  assign sel_248215 = array_index_248106 == array_index_239478 ? add_248214 : sel_248211;
  assign add_248218 = sel_248215 + 8'h01;
  assign sel_248219 = array_index_248106 == array_index_239484 ? add_248218 : sel_248215;
  assign add_248222 = sel_248219 + 8'h01;
  assign sel_248223 = array_index_248106 == array_index_239490 ? add_248222 : sel_248219;
  assign add_248226 = sel_248223 + 8'h01;
  assign sel_248227 = array_index_248106 == array_index_239496 ? add_248226 : sel_248223;
  assign add_248230 = sel_248227 + 8'h01;
  assign sel_248231 = array_index_248106 == array_index_239502 ? add_248230 : sel_248227;
  assign add_248234 = sel_248231 + 8'h01;
  assign sel_248235 = array_index_248106 == array_index_239508 ? add_248234 : sel_248231;
  assign add_248238 = sel_248235 + 8'h01;
  assign sel_248239 = array_index_248106 == array_index_239514 ? add_248238 : sel_248235;
  assign add_248242 = sel_248239 + 8'h01;
  assign sel_248243 = array_index_248106 == array_index_239520 ? add_248242 : sel_248239;
  assign add_248246 = sel_248243 + 8'h01;
  assign sel_248247 = array_index_248106 == array_index_239526 ? add_248246 : sel_248243;
  assign add_248250 = sel_248247 + 8'h01;
  assign sel_248251 = array_index_248106 == array_index_239532 ? add_248250 : sel_248247;
  assign add_248254 = sel_248251 + 8'h01;
  assign sel_248255 = array_index_248106 == array_index_239538 ? add_248254 : sel_248251;
  assign add_248258 = sel_248255 + 8'h01;
  assign sel_248259 = array_index_248106 == array_index_239544 ? add_248258 : sel_248255;
  assign add_248262 = sel_248259 + 8'h01;
  assign sel_248263 = array_index_248106 == array_index_239550 ? add_248262 : sel_248259;
  assign add_248266 = sel_248263 + 8'h01;
  assign sel_248267 = array_index_248106 == array_index_239556 ? add_248266 : sel_248263;
  assign add_248270 = sel_248267 + 8'h01;
  assign sel_248271 = array_index_248106 == array_index_239562 ? add_248270 : sel_248267;
  assign add_248274 = sel_248271 + 8'h01;
  assign sel_248275 = array_index_248106 == array_index_239568 ? add_248274 : sel_248271;
  assign add_248278 = sel_248275 + 8'h01;
  assign sel_248279 = array_index_248106 == array_index_239574 ? add_248278 : sel_248275;
  assign add_248282 = sel_248279 + 8'h01;
  assign sel_248283 = array_index_248106 == array_index_239580 ? add_248282 : sel_248279;
  assign add_248286 = sel_248283 + 8'h01;
  assign sel_248287 = array_index_248106 == array_index_239586 ? add_248286 : sel_248283;
  assign add_248290 = sel_248287 + 8'h01;
  assign sel_248291 = array_index_248106 == array_index_239592 ? add_248290 : sel_248287;
  assign add_248294 = sel_248291 + 8'h01;
  assign sel_248295 = array_index_248106 == array_index_239598 ? add_248294 : sel_248291;
  assign add_248298 = sel_248295 + 8'h01;
  assign sel_248299 = array_index_248106 == array_index_239604 ? add_248298 : sel_248295;
  assign add_248302 = sel_248299 + 8'h01;
  assign sel_248303 = array_index_248106 == array_index_239610 ? add_248302 : sel_248299;
  assign add_248307 = sel_248303 + 8'h01;
  assign array_index_248308 = set1_unflattened[6'h2c];
  assign sel_248309 = array_index_248106 == array_index_239616 ? add_248307 : sel_248303;
  assign add_248312 = sel_248309 + 8'h01;
  assign sel_248313 = array_index_248308 == array_index_239312 ? add_248312 : sel_248309;
  assign add_248316 = sel_248313 + 8'h01;
  assign sel_248317 = array_index_248308 == array_index_239316 ? add_248316 : sel_248313;
  assign add_248320 = sel_248317 + 8'h01;
  assign sel_248321 = array_index_248308 == array_index_239324 ? add_248320 : sel_248317;
  assign add_248324 = sel_248321 + 8'h01;
  assign sel_248325 = array_index_248308 == array_index_239332 ? add_248324 : sel_248321;
  assign add_248328 = sel_248325 + 8'h01;
  assign sel_248329 = array_index_248308 == array_index_239340 ? add_248328 : sel_248325;
  assign add_248332 = sel_248329 + 8'h01;
  assign sel_248333 = array_index_248308 == array_index_239348 ? add_248332 : sel_248329;
  assign add_248336 = sel_248333 + 8'h01;
  assign sel_248337 = array_index_248308 == array_index_239356 ? add_248336 : sel_248333;
  assign add_248340 = sel_248337 + 8'h01;
  assign sel_248341 = array_index_248308 == array_index_239364 ? add_248340 : sel_248337;
  assign add_248344 = sel_248341 + 8'h01;
  assign sel_248345 = array_index_248308 == array_index_239370 ? add_248344 : sel_248341;
  assign add_248348 = sel_248345 + 8'h01;
  assign sel_248349 = array_index_248308 == array_index_239376 ? add_248348 : sel_248345;
  assign add_248352 = sel_248349 + 8'h01;
  assign sel_248353 = array_index_248308 == array_index_239382 ? add_248352 : sel_248349;
  assign add_248356 = sel_248353 + 8'h01;
  assign sel_248357 = array_index_248308 == array_index_239388 ? add_248356 : sel_248353;
  assign add_248360 = sel_248357 + 8'h01;
  assign sel_248361 = array_index_248308 == array_index_239394 ? add_248360 : sel_248357;
  assign add_248364 = sel_248361 + 8'h01;
  assign sel_248365 = array_index_248308 == array_index_239400 ? add_248364 : sel_248361;
  assign add_248368 = sel_248365 + 8'h01;
  assign sel_248369 = array_index_248308 == array_index_239406 ? add_248368 : sel_248365;
  assign add_248372 = sel_248369 + 8'h01;
  assign sel_248373 = array_index_248308 == array_index_239412 ? add_248372 : sel_248369;
  assign add_248376 = sel_248373 + 8'h01;
  assign sel_248377 = array_index_248308 == array_index_239418 ? add_248376 : sel_248373;
  assign add_248380 = sel_248377 + 8'h01;
  assign sel_248381 = array_index_248308 == array_index_239424 ? add_248380 : sel_248377;
  assign add_248384 = sel_248381 + 8'h01;
  assign sel_248385 = array_index_248308 == array_index_239430 ? add_248384 : sel_248381;
  assign add_248388 = sel_248385 + 8'h01;
  assign sel_248389 = array_index_248308 == array_index_239436 ? add_248388 : sel_248385;
  assign add_248392 = sel_248389 + 8'h01;
  assign sel_248393 = array_index_248308 == array_index_239442 ? add_248392 : sel_248389;
  assign add_248396 = sel_248393 + 8'h01;
  assign sel_248397 = array_index_248308 == array_index_239448 ? add_248396 : sel_248393;
  assign add_248400 = sel_248397 + 8'h01;
  assign sel_248401 = array_index_248308 == array_index_239454 ? add_248400 : sel_248397;
  assign add_248404 = sel_248401 + 8'h01;
  assign sel_248405 = array_index_248308 == array_index_239460 ? add_248404 : sel_248401;
  assign add_248408 = sel_248405 + 8'h01;
  assign sel_248409 = array_index_248308 == array_index_239466 ? add_248408 : sel_248405;
  assign add_248412 = sel_248409 + 8'h01;
  assign sel_248413 = array_index_248308 == array_index_239472 ? add_248412 : sel_248409;
  assign add_248416 = sel_248413 + 8'h01;
  assign sel_248417 = array_index_248308 == array_index_239478 ? add_248416 : sel_248413;
  assign add_248420 = sel_248417 + 8'h01;
  assign sel_248421 = array_index_248308 == array_index_239484 ? add_248420 : sel_248417;
  assign add_248424 = sel_248421 + 8'h01;
  assign sel_248425 = array_index_248308 == array_index_239490 ? add_248424 : sel_248421;
  assign add_248428 = sel_248425 + 8'h01;
  assign sel_248429 = array_index_248308 == array_index_239496 ? add_248428 : sel_248425;
  assign add_248432 = sel_248429 + 8'h01;
  assign sel_248433 = array_index_248308 == array_index_239502 ? add_248432 : sel_248429;
  assign add_248436 = sel_248433 + 8'h01;
  assign sel_248437 = array_index_248308 == array_index_239508 ? add_248436 : sel_248433;
  assign add_248440 = sel_248437 + 8'h01;
  assign sel_248441 = array_index_248308 == array_index_239514 ? add_248440 : sel_248437;
  assign add_248444 = sel_248441 + 8'h01;
  assign sel_248445 = array_index_248308 == array_index_239520 ? add_248444 : sel_248441;
  assign add_248448 = sel_248445 + 8'h01;
  assign sel_248449 = array_index_248308 == array_index_239526 ? add_248448 : sel_248445;
  assign add_248452 = sel_248449 + 8'h01;
  assign sel_248453 = array_index_248308 == array_index_239532 ? add_248452 : sel_248449;
  assign add_248456 = sel_248453 + 8'h01;
  assign sel_248457 = array_index_248308 == array_index_239538 ? add_248456 : sel_248453;
  assign add_248460 = sel_248457 + 8'h01;
  assign sel_248461 = array_index_248308 == array_index_239544 ? add_248460 : sel_248457;
  assign add_248464 = sel_248461 + 8'h01;
  assign sel_248465 = array_index_248308 == array_index_239550 ? add_248464 : sel_248461;
  assign add_248468 = sel_248465 + 8'h01;
  assign sel_248469 = array_index_248308 == array_index_239556 ? add_248468 : sel_248465;
  assign add_248472 = sel_248469 + 8'h01;
  assign sel_248473 = array_index_248308 == array_index_239562 ? add_248472 : sel_248469;
  assign add_248476 = sel_248473 + 8'h01;
  assign sel_248477 = array_index_248308 == array_index_239568 ? add_248476 : sel_248473;
  assign add_248480 = sel_248477 + 8'h01;
  assign sel_248481 = array_index_248308 == array_index_239574 ? add_248480 : sel_248477;
  assign add_248484 = sel_248481 + 8'h01;
  assign sel_248485 = array_index_248308 == array_index_239580 ? add_248484 : sel_248481;
  assign add_248488 = sel_248485 + 8'h01;
  assign sel_248489 = array_index_248308 == array_index_239586 ? add_248488 : sel_248485;
  assign add_248492 = sel_248489 + 8'h01;
  assign sel_248493 = array_index_248308 == array_index_239592 ? add_248492 : sel_248489;
  assign add_248496 = sel_248493 + 8'h01;
  assign sel_248497 = array_index_248308 == array_index_239598 ? add_248496 : sel_248493;
  assign add_248500 = sel_248497 + 8'h01;
  assign sel_248501 = array_index_248308 == array_index_239604 ? add_248500 : sel_248497;
  assign add_248504 = sel_248501 + 8'h01;
  assign sel_248505 = array_index_248308 == array_index_239610 ? add_248504 : sel_248501;
  assign add_248509 = sel_248505 + 8'h01;
  assign array_index_248510 = set1_unflattened[6'h2d];
  assign sel_248511 = array_index_248308 == array_index_239616 ? add_248509 : sel_248505;
  assign add_248514 = sel_248511 + 8'h01;
  assign sel_248515 = array_index_248510 == array_index_239312 ? add_248514 : sel_248511;
  assign add_248518 = sel_248515 + 8'h01;
  assign sel_248519 = array_index_248510 == array_index_239316 ? add_248518 : sel_248515;
  assign add_248522 = sel_248519 + 8'h01;
  assign sel_248523 = array_index_248510 == array_index_239324 ? add_248522 : sel_248519;
  assign add_248526 = sel_248523 + 8'h01;
  assign sel_248527 = array_index_248510 == array_index_239332 ? add_248526 : sel_248523;
  assign add_248530 = sel_248527 + 8'h01;
  assign sel_248531 = array_index_248510 == array_index_239340 ? add_248530 : sel_248527;
  assign add_248534 = sel_248531 + 8'h01;
  assign sel_248535 = array_index_248510 == array_index_239348 ? add_248534 : sel_248531;
  assign add_248538 = sel_248535 + 8'h01;
  assign sel_248539 = array_index_248510 == array_index_239356 ? add_248538 : sel_248535;
  assign add_248542 = sel_248539 + 8'h01;
  assign sel_248543 = array_index_248510 == array_index_239364 ? add_248542 : sel_248539;
  assign add_248546 = sel_248543 + 8'h01;
  assign sel_248547 = array_index_248510 == array_index_239370 ? add_248546 : sel_248543;
  assign add_248550 = sel_248547 + 8'h01;
  assign sel_248551 = array_index_248510 == array_index_239376 ? add_248550 : sel_248547;
  assign add_248554 = sel_248551 + 8'h01;
  assign sel_248555 = array_index_248510 == array_index_239382 ? add_248554 : sel_248551;
  assign add_248558 = sel_248555 + 8'h01;
  assign sel_248559 = array_index_248510 == array_index_239388 ? add_248558 : sel_248555;
  assign add_248562 = sel_248559 + 8'h01;
  assign sel_248563 = array_index_248510 == array_index_239394 ? add_248562 : sel_248559;
  assign add_248566 = sel_248563 + 8'h01;
  assign sel_248567 = array_index_248510 == array_index_239400 ? add_248566 : sel_248563;
  assign add_248570 = sel_248567 + 8'h01;
  assign sel_248571 = array_index_248510 == array_index_239406 ? add_248570 : sel_248567;
  assign add_248574 = sel_248571 + 8'h01;
  assign sel_248575 = array_index_248510 == array_index_239412 ? add_248574 : sel_248571;
  assign add_248578 = sel_248575 + 8'h01;
  assign sel_248579 = array_index_248510 == array_index_239418 ? add_248578 : sel_248575;
  assign add_248582 = sel_248579 + 8'h01;
  assign sel_248583 = array_index_248510 == array_index_239424 ? add_248582 : sel_248579;
  assign add_248586 = sel_248583 + 8'h01;
  assign sel_248587 = array_index_248510 == array_index_239430 ? add_248586 : sel_248583;
  assign add_248590 = sel_248587 + 8'h01;
  assign sel_248591 = array_index_248510 == array_index_239436 ? add_248590 : sel_248587;
  assign add_248594 = sel_248591 + 8'h01;
  assign sel_248595 = array_index_248510 == array_index_239442 ? add_248594 : sel_248591;
  assign add_248598 = sel_248595 + 8'h01;
  assign sel_248599 = array_index_248510 == array_index_239448 ? add_248598 : sel_248595;
  assign add_248602 = sel_248599 + 8'h01;
  assign sel_248603 = array_index_248510 == array_index_239454 ? add_248602 : sel_248599;
  assign add_248606 = sel_248603 + 8'h01;
  assign sel_248607 = array_index_248510 == array_index_239460 ? add_248606 : sel_248603;
  assign add_248610 = sel_248607 + 8'h01;
  assign sel_248611 = array_index_248510 == array_index_239466 ? add_248610 : sel_248607;
  assign add_248614 = sel_248611 + 8'h01;
  assign sel_248615 = array_index_248510 == array_index_239472 ? add_248614 : sel_248611;
  assign add_248618 = sel_248615 + 8'h01;
  assign sel_248619 = array_index_248510 == array_index_239478 ? add_248618 : sel_248615;
  assign add_248622 = sel_248619 + 8'h01;
  assign sel_248623 = array_index_248510 == array_index_239484 ? add_248622 : sel_248619;
  assign add_248626 = sel_248623 + 8'h01;
  assign sel_248627 = array_index_248510 == array_index_239490 ? add_248626 : sel_248623;
  assign add_248630 = sel_248627 + 8'h01;
  assign sel_248631 = array_index_248510 == array_index_239496 ? add_248630 : sel_248627;
  assign add_248634 = sel_248631 + 8'h01;
  assign sel_248635 = array_index_248510 == array_index_239502 ? add_248634 : sel_248631;
  assign add_248638 = sel_248635 + 8'h01;
  assign sel_248639 = array_index_248510 == array_index_239508 ? add_248638 : sel_248635;
  assign add_248642 = sel_248639 + 8'h01;
  assign sel_248643 = array_index_248510 == array_index_239514 ? add_248642 : sel_248639;
  assign add_248646 = sel_248643 + 8'h01;
  assign sel_248647 = array_index_248510 == array_index_239520 ? add_248646 : sel_248643;
  assign add_248650 = sel_248647 + 8'h01;
  assign sel_248651 = array_index_248510 == array_index_239526 ? add_248650 : sel_248647;
  assign add_248654 = sel_248651 + 8'h01;
  assign sel_248655 = array_index_248510 == array_index_239532 ? add_248654 : sel_248651;
  assign add_248658 = sel_248655 + 8'h01;
  assign sel_248659 = array_index_248510 == array_index_239538 ? add_248658 : sel_248655;
  assign add_248662 = sel_248659 + 8'h01;
  assign sel_248663 = array_index_248510 == array_index_239544 ? add_248662 : sel_248659;
  assign add_248666 = sel_248663 + 8'h01;
  assign sel_248667 = array_index_248510 == array_index_239550 ? add_248666 : sel_248663;
  assign add_248670 = sel_248667 + 8'h01;
  assign sel_248671 = array_index_248510 == array_index_239556 ? add_248670 : sel_248667;
  assign add_248674 = sel_248671 + 8'h01;
  assign sel_248675 = array_index_248510 == array_index_239562 ? add_248674 : sel_248671;
  assign add_248678 = sel_248675 + 8'h01;
  assign sel_248679 = array_index_248510 == array_index_239568 ? add_248678 : sel_248675;
  assign add_248682 = sel_248679 + 8'h01;
  assign sel_248683 = array_index_248510 == array_index_239574 ? add_248682 : sel_248679;
  assign add_248686 = sel_248683 + 8'h01;
  assign sel_248687 = array_index_248510 == array_index_239580 ? add_248686 : sel_248683;
  assign add_248690 = sel_248687 + 8'h01;
  assign sel_248691 = array_index_248510 == array_index_239586 ? add_248690 : sel_248687;
  assign add_248694 = sel_248691 + 8'h01;
  assign sel_248695 = array_index_248510 == array_index_239592 ? add_248694 : sel_248691;
  assign add_248698 = sel_248695 + 8'h01;
  assign sel_248699 = array_index_248510 == array_index_239598 ? add_248698 : sel_248695;
  assign add_248702 = sel_248699 + 8'h01;
  assign sel_248703 = array_index_248510 == array_index_239604 ? add_248702 : sel_248699;
  assign add_248706 = sel_248703 + 8'h01;
  assign sel_248707 = array_index_248510 == array_index_239610 ? add_248706 : sel_248703;
  assign add_248711 = sel_248707 + 8'h01;
  assign array_index_248712 = set1_unflattened[6'h2e];
  assign sel_248713 = array_index_248510 == array_index_239616 ? add_248711 : sel_248707;
  assign add_248716 = sel_248713 + 8'h01;
  assign sel_248717 = array_index_248712 == array_index_239312 ? add_248716 : sel_248713;
  assign add_248720 = sel_248717 + 8'h01;
  assign sel_248721 = array_index_248712 == array_index_239316 ? add_248720 : sel_248717;
  assign add_248724 = sel_248721 + 8'h01;
  assign sel_248725 = array_index_248712 == array_index_239324 ? add_248724 : sel_248721;
  assign add_248728 = sel_248725 + 8'h01;
  assign sel_248729 = array_index_248712 == array_index_239332 ? add_248728 : sel_248725;
  assign add_248732 = sel_248729 + 8'h01;
  assign sel_248733 = array_index_248712 == array_index_239340 ? add_248732 : sel_248729;
  assign add_248736 = sel_248733 + 8'h01;
  assign sel_248737 = array_index_248712 == array_index_239348 ? add_248736 : sel_248733;
  assign add_248740 = sel_248737 + 8'h01;
  assign sel_248741 = array_index_248712 == array_index_239356 ? add_248740 : sel_248737;
  assign add_248744 = sel_248741 + 8'h01;
  assign sel_248745 = array_index_248712 == array_index_239364 ? add_248744 : sel_248741;
  assign add_248748 = sel_248745 + 8'h01;
  assign sel_248749 = array_index_248712 == array_index_239370 ? add_248748 : sel_248745;
  assign add_248752 = sel_248749 + 8'h01;
  assign sel_248753 = array_index_248712 == array_index_239376 ? add_248752 : sel_248749;
  assign add_248756 = sel_248753 + 8'h01;
  assign sel_248757 = array_index_248712 == array_index_239382 ? add_248756 : sel_248753;
  assign add_248760 = sel_248757 + 8'h01;
  assign sel_248761 = array_index_248712 == array_index_239388 ? add_248760 : sel_248757;
  assign add_248764 = sel_248761 + 8'h01;
  assign sel_248765 = array_index_248712 == array_index_239394 ? add_248764 : sel_248761;
  assign add_248768 = sel_248765 + 8'h01;
  assign sel_248769 = array_index_248712 == array_index_239400 ? add_248768 : sel_248765;
  assign add_248772 = sel_248769 + 8'h01;
  assign sel_248773 = array_index_248712 == array_index_239406 ? add_248772 : sel_248769;
  assign add_248776 = sel_248773 + 8'h01;
  assign sel_248777 = array_index_248712 == array_index_239412 ? add_248776 : sel_248773;
  assign add_248780 = sel_248777 + 8'h01;
  assign sel_248781 = array_index_248712 == array_index_239418 ? add_248780 : sel_248777;
  assign add_248784 = sel_248781 + 8'h01;
  assign sel_248785 = array_index_248712 == array_index_239424 ? add_248784 : sel_248781;
  assign add_248788 = sel_248785 + 8'h01;
  assign sel_248789 = array_index_248712 == array_index_239430 ? add_248788 : sel_248785;
  assign add_248792 = sel_248789 + 8'h01;
  assign sel_248793 = array_index_248712 == array_index_239436 ? add_248792 : sel_248789;
  assign add_248796 = sel_248793 + 8'h01;
  assign sel_248797 = array_index_248712 == array_index_239442 ? add_248796 : sel_248793;
  assign add_248800 = sel_248797 + 8'h01;
  assign sel_248801 = array_index_248712 == array_index_239448 ? add_248800 : sel_248797;
  assign add_248804 = sel_248801 + 8'h01;
  assign sel_248805 = array_index_248712 == array_index_239454 ? add_248804 : sel_248801;
  assign add_248808 = sel_248805 + 8'h01;
  assign sel_248809 = array_index_248712 == array_index_239460 ? add_248808 : sel_248805;
  assign add_248812 = sel_248809 + 8'h01;
  assign sel_248813 = array_index_248712 == array_index_239466 ? add_248812 : sel_248809;
  assign add_248816 = sel_248813 + 8'h01;
  assign sel_248817 = array_index_248712 == array_index_239472 ? add_248816 : sel_248813;
  assign add_248820 = sel_248817 + 8'h01;
  assign sel_248821 = array_index_248712 == array_index_239478 ? add_248820 : sel_248817;
  assign add_248824 = sel_248821 + 8'h01;
  assign sel_248825 = array_index_248712 == array_index_239484 ? add_248824 : sel_248821;
  assign add_248828 = sel_248825 + 8'h01;
  assign sel_248829 = array_index_248712 == array_index_239490 ? add_248828 : sel_248825;
  assign add_248832 = sel_248829 + 8'h01;
  assign sel_248833 = array_index_248712 == array_index_239496 ? add_248832 : sel_248829;
  assign add_248836 = sel_248833 + 8'h01;
  assign sel_248837 = array_index_248712 == array_index_239502 ? add_248836 : sel_248833;
  assign add_248840 = sel_248837 + 8'h01;
  assign sel_248841 = array_index_248712 == array_index_239508 ? add_248840 : sel_248837;
  assign add_248844 = sel_248841 + 8'h01;
  assign sel_248845 = array_index_248712 == array_index_239514 ? add_248844 : sel_248841;
  assign add_248848 = sel_248845 + 8'h01;
  assign sel_248849 = array_index_248712 == array_index_239520 ? add_248848 : sel_248845;
  assign add_248852 = sel_248849 + 8'h01;
  assign sel_248853 = array_index_248712 == array_index_239526 ? add_248852 : sel_248849;
  assign add_248856 = sel_248853 + 8'h01;
  assign sel_248857 = array_index_248712 == array_index_239532 ? add_248856 : sel_248853;
  assign add_248860 = sel_248857 + 8'h01;
  assign sel_248861 = array_index_248712 == array_index_239538 ? add_248860 : sel_248857;
  assign add_248864 = sel_248861 + 8'h01;
  assign sel_248865 = array_index_248712 == array_index_239544 ? add_248864 : sel_248861;
  assign add_248868 = sel_248865 + 8'h01;
  assign sel_248869 = array_index_248712 == array_index_239550 ? add_248868 : sel_248865;
  assign add_248872 = sel_248869 + 8'h01;
  assign sel_248873 = array_index_248712 == array_index_239556 ? add_248872 : sel_248869;
  assign add_248876 = sel_248873 + 8'h01;
  assign sel_248877 = array_index_248712 == array_index_239562 ? add_248876 : sel_248873;
  assign add_248880 = sel_248877 + 8'h01;
  assign sel_248881 = array_index_248712 == array_index_239568 ? add_248880 : sel_248877;
  assign add_248884 = sel_248881 + 8'h01;
  assign sel_248885 = array_index_248712 == array_index_239574 ? add_248884 : sel_248881;
  assign add_248888 = sel_248885 + 8'h01;
  assign sel_248889 = array_index_248712 == array_index_239580 ? add_248888 : sel_248885;
  assign add_248892 = sel_248889 + 8'h01;
  assign sel_248893 = array_index_248712 == array_index_239586 ? add_248892 : sel_248889;
  assign add_248896 = sel_248893 + 8'h01;
  assign sel_248897 = array_index_248712 == array_index_239592 ? add_248896 : sel_248893;
  assign add_248900 = sel_248897 + 8'h01;
  assign sel_248901 = array_index_248712 == array_index_239598 ? add_248900 : sel_248897;
  assign add_248904 = sel_248901 + 8'h01;
  assign sel_248905 = array_index_248712 == array_index_239604 ? add_248904 : sel_248901;
  assign add_248908 = sel_248905 + 8'h01;
  assign sel_248909 = array_index_248712 == array_index_239610 ? add_248908 : sel_248905;
  assign add_248913 = sel_248909 + 8'h01;
  assign array_index_248914 = set1_unflattened[6'h2f];
  assign sel_248915 = array_index_248712 == array_index_239616 ? add_248913 : sel_248909;
  assign add_248918 = sel_248915 + 8'h01;
  assign sel_248919 = array_index_248914 == array_index_239312 ? add_248918 : sel_248915;
  assign add_248922 = sel_248919 + 8'h01;
  assign sel_248923 = array_index_248914 == array_index_239316 ? add_248922 : sel_248919;
  assign add_248926 = sel_248923 + 8'h01;
  assign sel_248927 = array_index_248914 == array_index_239324 ? add_248926 : sel_248923;
  assign add_248930 = sel_248927 + 8'h01;
  assign sel_248931 = array_index_248914 == array_index_239332 ? add_248930 : sel_248927;
  assign add_248934 = sel_248931 + 8'h01;
  assign sel_248935 = array_index_248914 == array_index_239340 ? add_248934 : sel_248931;
  assign add_248938 = sel_248935 + 8'h01;
  assign sel_248939 = array_index_248914 == array_index_239348 ? add_248938 : sel_248935;
  assign add_248942 = sel_248939 + 8'h01;
  assign sel_248943 = array_index_248914 == array_index_239356 ? add_248942 : sel_248939;
  assign add_248946 = sel_248943 + 8'h01;
  assign sel_248947 = array_index_248914 == array_index_239364 ? add_248946 : sel_248943;
  assign add_248950 = sel_248947 + 8'h01;
  assign sel_248951 = array_index_248914 == array_index_239370 ? add_248950 : sel_248947;
  assign add_248954 = sel_248951 + 8'h01;
  assign sel_248955 = array_index_248914 == array_index_239376 ? add_248954 : sel_248951;
  assign add_248958 = sel_248955 + 8'h01;
  assign sel_248959 = array_index_248914 == array_index_239382 ? add_248958 : sel_248955;
  assign add_248962 = sel_248959 + 8'h01;
  assign sel_248963 = array_index_248914 == array_index_239388 ? add_248962 : sel_248959;
  assign add_248966 = sel_248963 + 8'h01;
  assign sel_248967 = array_index_248914 == array_index_239394 ? add_248966 : sel_248963;
  assign add_248970 = sel_248967 + 8'h01;
  assign sel_248971 = array_index_248914 == array_index_239400 ? add_248970 : sel_248967;
  assign add_248974 = sel_248971 + 8'h01;
  assign sel_248975 = array_index_248914 == array_index_239406 ? add_248974 : sel_248971;
  assign add_248978 = sel_248975 + 8'h01;
  assign sel_248979 = array_index_248914 == array_index_239412 ? add_248978 : sel_248975;
  assign add_248982 = sel_248979 + 8'h01;
  assign sel_248983 = array_index_248914 == array_index_239418 ? add_248982 : sel_248979;
  assign add_248986 = sel_248983 + 8'h01;
  assign sel_248987 = array_index_248914 == array_index_239424 ? add_248986 : sel_248983;
  assign add_248990 = sel_248987 + 8'h01;
  assign sel_248991 = array_index_248914 == array_index_239430 ? add_248990 : sel_248987;
  assign add_248994 = sel_248991 + 8'h01;
  assign sel_248995 = array_index_248914 == array_index_239436 ? add_248994 : sel_248991;
  assign add_248998 = sel_248995 + 8'h01;
  assign sel_248999 = array_index_248914 == array_index_239442 ? add_248998 : sel_248995;
  assign add_249002 = sel_248999 + 8'h01;
  assign sel_249003 = array_index_248914 == array_index_239448 ? add_249002 : sel_248999;
  assign add_249006 = sel_249003 + 8'h01;
  assign sel_249007 = array_index_248914 == array_index_239454 ? add_249006 : sel_249003;
  assign add_249010 = sel_249007 + 8'h01;
  assign sel_249011 = array_index_248914 == array_index_239460 ? add_249010 : sel_249007;
  assign add_249014 = sel_249011 + 8'h01;
  assign sel_249015 = array_index_248914 == array_index_239466 ? add_249014 : sel_249011;
  assign add_249018 = sel_249015 + 8'h01;
  assign sel_249019 = array_index_248914 == array_index_239472 ? add_249018 : sel_249015;
  assign add_249022 = sel_249019 + 8'h01;
  assign sel_249023 = array_index_248914 == array_index_239478 ? add_249022 : sel_249019;
  assign add_249026 = sel_249023 + 8'h01;
  assign sel_249027 = array_index_248914 == array_index_239484 ? add_249026 : sel_249023;
  assign add_249030 = sel_249027 + 8'h01;
  assign sel_249031 = array_index_248914 == array_index_239490 ? add_249030 : sel_249027;
  assign add_249034 = sel_249031 + 8'h01;
  assign sel_249035 = array_index_248914 == array_index_239496 ? add_249034 : sel_249031;
  assign add_249038 = sel_249035 + 8'h01;
  assign sel_249039 = array_index_248914 == array_index_239502 ? add_249038 : sel_249035;
  assign add_249042 = sel_249039 + 8'h01;
  assign sel_249043 = array_index_248914 == array_index_239508 ? add_249042 : sel_249039;
  assign add_249046 = sel_249043 + 8'h01;
  assign sel_249047 = array_index_248914 == array_index_239514 ? add_249046 : sel_249043;
  assign add_249050 = sel_249047 + 8'h01;
  assign sel_249051 = array_index_248914 == array_index_239520 ? add_249050 : sel_249047;
  assign add_249054 = sel_249051 + 8'h01;
  assign sel_249055 = array_index_248914 == array_index_239526 ? add_249054 : sel_249051;
  assign add_249058 = sel_249055 + 8'h01;
  assign sel_249059 = array_index_248914 == array_index_239532 ? add_249058 : sel_249055;
  assign add_249062 = sel_249059 + 8'h01;
  assign sel_249063 = array_index_248914 == array_index_239538 ? add_249062 : sel_249059;
  assign add_249066 = sel_249063 + 8'h01;
  assign sel_249067 = array_index_248914 == array_index_239544 ? add_249066 : sel_249063;
  assign add_249070 = sel_249067 + 8'h01;
  assign sel_249071 = array_index_248914 == array_index_239550 ? add_249070 : sel_249067;
  assign add_249074 = sel_249071 + 8'h01;
  assign sel_249075 = array_index_248914 == array_index_239556 ? add_249074 : sel_249071;
  assign add_249078 = sel_249075 + 8'h01;
  assign sel_249079 = array_index_248914 == array_index_239562 ? add_249078 : sel_249075;
  assign add_249082 = sel_249079 + 8'h01;
  assign sel_249083 = array_index_248914 == array_index_239568 ? add_249082 : sel_249079;
  assign add_249086 = sel_249083 + 8'h01;
  assign sel_249087 = array_index_248914 == array_index_239574 ? add_249086 : sel_249083;
  assign add_249090 = sel_249087 + 8'h01;
  assign sel_249091 = array_index_248914 == array_index_239580 ? add_249090 : sel_249087;
  assign add_249094 = sel_249091 + 8'h01;
  assign sel_249095 = array_index_248914 == array_index_239586 ? add_249094 : sel_249091;
  assign add_249098 = sel_249095 + 8'h01;
  assign sel_249099 = array_index_248914 == array_index_239592 ? add_249098 : sel_249095;
  assign add_249102 = sel_249099 + 8'h01;
  assign sel_249103 = array_index_248914 == array_index_239598 ? add_249102 : sel_249099;
  assign add_249106 = sel_249103 + 8'h01;
  assign sel_249107 = array_index_248914 == array_index_239604 ? add_249106 : sel_249103;
  assign add_249110 = sel_249107 + 8'h01;
  assign sel_249111 = array_index_248914 == array_index_239610 ? add_249110 : sel_249107;
  assign add_249115 = sel_249111 + 8'h01;
  assign array_index_249116 = set1_unflattened[6'h30];
  assign sel_249117 = array_index_248914 == array_index_239616 ? add_249115 : sel_249111;
  assign add_249120 = sel_249117 + 8'h01;
  assign sel_249121 = array_index_249116 == array_index_239312 ? add_249120 : sel_249117;
  assign add_249124 = sel_249121 + 8'h01;
  assign sel_249125 = array_index_249116 == array_index_239316 ? add_249124 : sel_249121;
  assign add_249128 = sel_249125 + 8'h01;
  assign sel_249129 = array_index_249116 == array_index_239324 ? add_249128 : sel_249125;
  assign add_249132 = sel_249129 + 8'h01;
  assign sel_249133 = array_index_249116 == array_index_239332 ? add_249132 : sel_249129;
  assign add_249136 = sel_249133 + 8'h01;
  assign sel_249137 = array_index_249116 == array_index_239340 ? add_249136 : sel_249133;
  assign add_249140 = sel_249137 + 8'h01;
  assign sel_249141 = array_index_249116 == array_index_239348 ? add_249140 : sel_249137;
  assign add_249144 = sel_249141 + 8'h01;
  assign sel_249145 = array_index_249116 == array_index_239356 ? add_249144 : sel_249141;
  assign add_249148 = sel_249145 + 8'h01;
  assign sel_249149 = array_index_249116 == array_index_239364 ? add_249148 : sel_249145;
  assign add_249152 = sel_249149 + 8'h01;
  assign sel_249153 = array_index_249116 == array_index_239370 ? add_249152 : sel_249149;
  assign add_249156 = sel_249153 + 8'h01;
  assign sel_249157 = array_index_249116 == array_index_239376 ? add_249156 : sel_249153;
  assign add_249160 = sel_249157 + 8'h01;
  assign sel_249161 = array_index_249116 == array_index_239382 ? add_249160 : sel_249157;
  assign add_249164 = sel_249161 + 8'h01;
  assign sel_249165 = array_index_249116 == array_index_239388 ? add_249164 : sel_249161;
  assign add_249168 = sel_249165 + 8'h01;
  assign sel_249169 = array_index_249116 == array_index_239394 ? add_249168 : sel_249165;
  assign add_249172 = sel_249169 + 8'h01;
  assign sel_249173 = array_index_249116 == array_index_239400 ? add_249172 : sel_249169;
  assign add_249176 = sel_249173 + 8'h01;
  assign sel_249177 = array_index_249116 == array_index_239406 ? add_249176 : sel_249173;
  assign add_249180 = sel_249177 + 8'h01;
  assign sel_249181 = array_index_249116 == array_index_239412 ? add_249180 : sel_249177;
  assign add_249184 = sel_249181 + 8'h01;
  assign sel_249185 = array_index_249116 == array_index_239418 ? add_249184 : sel_249181;
  assign add_249188 = sel_249185 + 8'h01;
  assign sel_249189 = array_index_249116 == array_index_239424 ? add_249188 : sel_249185;
  assign add_249192 = sel_249189 + 8'h01;
  assign sel_249193 = array_index_249116 == array_index_239430 ? add_249192 : sel_249189;
  assign add_249196 = sel_249193 + 8'h01;
  assign sel_249197 = array_index_249116 == array_index_239436 ? add_249196 : sel_249193;
  assign add_249200 = sel_249197 + 8'h01;
  assign sel_249201 = array_index_249116 == array_index_239442 ? add_249200 : sel_249197;
  assign add_249204 = sel_249201 + 8'h01;
  assign sel_249205 = array_index_249116 == array_index_239448 ? add_249204 : sel_249201;
  assign add_249208 = sel_249205 + 8'h01;
  assign sel_249209 = array_index_249116 == array_index_239454 ? add_249208 : sel_249205;
  assign add_249212 = sel_249209 + 8'h01;
  assign sel_249213 = array_index_249116 == array_index_239460 ? add_249212 : sel_249209;
  assign add_249216 = sel_249213 + 8'h01;
  assign sel_249217 = array_index_249116 == array_index_239466 ? add_249216 : sel_249213;
  assign add_249220 = sel_249217 + 8'h01;
  assign sel_249221 = array_index_249116 == array_index_239472 ? add_249220 : sel_249217;
  assign add_249224 = sel_249221 + 8'h01;
  assign sel_249225 = array_index_249116 == array_index_239478 ? add_249224 : sel_249221;
  assign add_249228 = sel_249225 + 8'h01;
  assign sel_249229 = array_index_249116 == array_index_239484 ? add_249228 : sel_249225;
  assign add_249232 = sel_249229 + 8'h01;
  assign sel_249233 = array_index_249116 == array_index_239490 ? add_249232 : sel_249229;
  assign add_249236 = sel_249233 + 8'h01;
  assign sel_249237 = array_index_249116 == array_index_239496 ? add_249236 : sel_249233;
  assign add_249240 = sel_249237 + 8'h01;
  assign sel_249241 = array_index_249116 == array_index_239502 ? add_249240 : sel_249237;
  assign add_249244 = sel_249241 + 8'h01;
  assign sel_249245 = array_index_249116 == array_index_239508 ? add_249244 : sel_249241;
  assign add_249248 = sel_249245 + 8'h01;
  assign sel_249249 = array_index_249116 == array_index_239514 ? add_249248 : sel_249245;
  assign add_249252 = sel_249249 + 8'h01;
  assign sel_249253 = array_index_249116 == array_index_239520 ? add_249252 : sel_249249;
  assign add_249256 = sel_249253 + 8'h01;
  assign sel_249257 = array_index_249116 == array_index_239526 ? add_249256 : sel_249253;
  assign add_249260 = sel_249257 + 8'h01;
  assign sel_249261 = array_index_249116 == array_index_239532 ? add_249260 : sel_249257;
  assign add_249264 = sel_249261 + 8'h01;
  assign sel_249265 = array_index_249116 == array_index_239538 ? add_249264 : sel_249261;
  assign add_249268 = sel_249265 + 8'h01;
  assign sel_249269 = array_index_249116 == array_index_239544 ? add_249268 : sel_249265;
  assign add_249272 = sel_249269 + 8'h01;
  assign sel_249273 = array_index_249116 == array_index_239550 ? add_249272 : sel_249269;
  assign add_249276 = sel_249273 + 8'h01;
  assign sel_249277 = array_index_249116 == array_index_239556 ? add_249276 : sel_249273;
  assign add_249280 = sel_249277 + 8'h01;
  assign sel_249281 = array_index_249116 == array_index_239562 ? add_249280 : sel_249277;
  assign add_249284 = sel_249281 + 8'h01;
  assign sel_249285 = array_index_249116 == array_index_239568 ? add_249284 : sel_249281;
  assign add_249288 = sel_249285 + 8'h01;
  assign sel_249289 = array_index_249116 == array_index_239574 ? add_249288 : sel_249285;
  assign add_249292 = sel_249289 + 8'h01;
  assign sel_249293 = array_index_249116 == array_index_239580 ? add_249292 : sel_249289;
  assign add_249296 = sel_249293 + 8'h01;
  assign sel_249297 = array_index_249116 == array_index_239586 ? add_249296 : sel_249293;
  assign add_249300 = sel_249297 + 8'h01;
  assign sel_249301 = array_index_249116 == array_index_239592 ? add_249300 : sel_249297;
  assign add_249304 = sel_249301 + 8'h01;
  assign sel_249305 = array_index_249116 == array_index_239598 ? add_249304 : sel_249301;
  assign add_249308 = sel_249305 + 8'h01;
  assign sel_249309 = array_index_249116 == array_index_239604 ? add_249308 : sel_249305;
  assign add_249312 = sel_249309 + 8'h01;
  assign sel_249313 = array_index_249116 == array_index_239610 ? add_249312 : sel_249309;
  assign add_249317 = sel_249313 + 8'h01;
  assign array_index_249318 = set1_unflattened[6'h31];
  assign sel_249319 = array_index_249116 == array_index_239616 ? add_249317 : sel_249313;
  assign add_249322 = sel_249319 + 8'h01;
  assign sel_249323 = array_index_249318 == array_index_239312 ? add_249322 : sel_249319;
  assign add_249326 = sel_249323 + 8'h01;
  assign sel_249327 = array_index_249318 == array_index_239316 ? add_249326 : sel_249323;
  assign add_249330 = sel_249327 + 8'h01;
  assign sel_249331 = array_index_249318 == array_index_239324 ? add_249330 : sel_249327;
  assign add_249334 = sel_249331 + 8'h01;
  assign sel_249335 = array_index_249318 == array_index_239332 ? add_249334 : sel_249331;
  assign add_249338 = sel_249335 + 8'h01;
  assign sel_249339 = array_index_249318 == array_index_239340 ? add_249338 : sel_249335;
  assign add_249342 = sel_249339 + 8'h01;
  assign sel_249343 = array_index_249318 == array_index_239348 ? add_249342 : sel_249339;
  assign add_249346 = sel_249343 + 8'h01;
  assign sel_249347 = array_index_249318 == array_index_239356 ? add_249346 : sel_249343;
  assign add_249350 = sel_249347 + 8'h01;
  assign sel_249351 = array_index_249318 == array_index_239364 ? add_249350 : sel_249347;
  assign add_249354 = sel_249351 + 8'h01;
  assign sel_249355 = array_index_249318 == array_index_239370 ? add_249354 : sel_249351;
  assign add_249358 = sel_249355 + 8'h01;
  assign sel_249359 = array_index_249318 == array_index_239376 ? add_249358 : sel_249355;
  assign add_249362 = sel_249359 + 8'h01;
  assign sel_249363 = array_index_249318 == array_index_239382 ? add_249362 : sel_249359;
  assign add_249366 = sel_249363 + 8'h01;
  assign sel_249367 = array_index_249318 == array_index_239388 ? add_249366 : sel_249363;
  assign add_249370 = sel_249367 + 8'h01;
  assign sel_249371 = array_index_249318 == array_index_239394 ? add_249370 : sel_249367;
  assign add_249374 = sel_249371 + 8'h01;
  assign sel_249375 = array_index_249318 == array_index_239400 ? add_249374 : sel_249371;
  assign add_249378 = sel_249375 + 8'h01;
  assign sel_249379 = array_index_249318 == array_index_239406 ? add_249378 : sel_249375;
  assign add_249382 = sel_249379 + 8'h01;
  assign sel_249383 = array_index_249318 == array_index_239412 ? add_249382 : sel_249379;
  assign add_249386 = sel_249383 + 8'h01;
  assign sel_249387 = array_index_249318 == array_index_239418 ? add_249386 : sel_249383;
  assign add_249390 = sel_249387 + 8'h01;
  assign sel_249391 = array_index_249318 == array_index_239424 ? add_249390 : sel_249387;
  assign add_249394 = sel_249391 + 8'h01;
  assign sel_249395 = array_index_249318 == array_index_239430 ? add_249394 : sel_249391;
  assign add_249398 = sel_249395 + 8'h01;
  assign sel_249399 = array_index_249318 == array_index_239436 ? add_249398 : sel_249395;
  assign add_249402 = sel_249399 + 8'h01;
  assign sel_249403 = array_index_249318 == array_index_239442 ? add_249402 : sel_249399;
  assign add_249406 = sel_249403 + 8'h01;
  assign sel_249407 = array_index_249318 == array_index_239448 ? add_249406 : sel_249403;
  assign add_249410 = sel_249407 + 8'h01;
  assign sel_249411 = array_index_249318 == array_index_239454 ? add_249410 : sel_249407;
  assign add_249414 = sel_249411 + 8'h01;
  assign sel_249415 = array_index_249318 == array_index_239460 ? add_249414 : sel_249411;
  assign add_249418 = sel_249415 + 8'h01;
  assign sel_249419 = array_index_249318 == array_index_239466 ? add_249418 : sel_249415;
  assign add_249422 = sel_249419 + 8'h01;
  assign sel_249423 = array_index_249318 == array_index_239472 ? add_249422 : sel_249419;
  assign add_249426 = sel_249423 + 8'h01;
  assign sel_249427 = array_index_249318 == array_index_239478 ? add_249426 : sel_249423;
  assign add_249430 = sel_249427 + 8'h01;
  assign sel_249431 = array_index_249318 == array_index_239484 ? add_249430 : sel_249427;
  assign add_249434 = sel_249431 + 8'h01;
  assign sel_249435 = array_index_249318 == array_index_239490 ? add_249434 : sel_249431;
  assign add_249438 = sel_249435 + 8'h01;
  assign sel_249439 = array_index_249318 == array_index_239496 ? add_249438 : sel_249435;
  assign add_249442 = sel_249439 + 8'h01;
  assign sel_249443 = array_index_249318 == array_index_239502 ? add_249442 : sel_249439;
  assign add_249446 = sel_249443 + 8'h01;
  assign sel_249447 = array_index_249318 == array_index_239508 ? add_249446 : sel_249443;
  assign add_249450 = sel_249447 + 8'h01;
  assign sel_249451 = array_index_249318 == array_index_239514 ? add_249450 : sel_249447;
  assign add_249454 = sel_249451 + 8'h01;
  assign sel_249455 = array_index_249318 == array_index_239520 ? add_249454 : sel_249451;
  assign add_249458 = sel_249455 + 8'h01;
  assign sel_249459 = array_index_249318 == array_index_239526 ? add_249458 : sel_249455;
  assign add_249462 = sel_249459 + 8'h01;
  assign sel_249463 = array_index_249318 == array_index_239532 ? add_249462 : sel_249459;
  assign add_249466 = sel_249463 + 8'h01;
  assign sel_249467 = array_index_249318 == array_index_239538 ? add_249466 : sel_249463;
  assign add_249470 = sel_249467 + 8'h01;
  assign sel_249471 = array_index_249318 == array_index_239544 ? add_249470 : sel_249467;
  assign add_249474 = sel_249471 + 8'h01;
  assign sel_249475 = array_index_249318 == array_index_239550 ? add_249474 : sel_249471;
  assign add_249478 = sel_249475 + 8'h01;
  assign sel_249479 = array_index_249318 == array_index_239556 ? add_249478 : sel_249475;
  assign add_249482 = sel_249479 + 8'h01;
  assign sel_249483 = array_index_249318 == array_index_239562 ? add_249482 : sel_249479;
  assign add_249486 = sel_249483 + 8'h01;
  assign sel_249487 = array_index_249318 == array_index_239568 ? add_249486 : sel_249483;
  assign add_249490 = sel_249487 + 8'h01;
  assign sel_249491 = array_index_249318 == array_index_239574 ? add_249490 : sel_249487;
  assign add_249494 = sel_249491 + 8'h01;
  assign sel_249495 = array_index_249318 == array_index_239580 ? add_249494 : sel_249491;
  assign add_249498 = sel_249495 + 8'h01;
  assign sel_249499 = array_index_249318 == array_index_239586 ? add_249498 : sel_249495;
  assign add_249502 = sel_249499 + 8'h01;
  assign sel_249503 = array_index_249318 == array_index_239592 ? add_249502 : sel_249499;
  assign add_249506 = sel_249503 + 8'h01;
  assign sel_249507 = array_index_249318 == array_index_239598 ? add_249506 : sel_249503;
  assign add_249510 = sel_249507 + 8'h01;
  assign sel_249511 = array_index_249318 == array_index_239604 ? add_249510 : sel_249507;
  assign add_249514 = sel_249511 + 8'h01;
  assign sel_249515 = array_index_249318 == array_index_239610 ? add_249514 : sel_249511;
  assign add_249518 = sel_249515 + 8'h01;
  assign out = {array_index_249318 == array_index_239616 ? add_249518 : sel_249515, {set1_unflattened[49], set1_unflattened[48], set1_unflattened[47], set1_unflattened[46], set1_unflattened[45], set1_unflattened[44], set1_unflattened[43], set1_unflattened[42], set1_unflattened[41], set1_unflattened[40], set1_unflattened[39], set1_unflattened[38], set1_unflattened[37], set1_unflattened[36], set1_unflattened[35], set1_unflattened[34], set1_unflattened[33], set1_unflattened[32], set1_unflattened[31], set1_unflattened[30], set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[49], set2_unflattened[48], set2_unflattened[47], set2_unflattened[46], set2_unflattened[45], set2_unflattened[44], set2_unflattened[43], set2_unflattened[42], set2_unflattened[41], set2_unflattened[40], set2_unflattened[39], set2_unflattened[38], set2_unflattened[37], set2_unflattened[36], set2_unflattened[35], set2_unflattened[34], set2_unflattened[33], set2_unflattened[32], set2_unflattened[31], set2_unflattened[30], set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
