module min_hash(
  input wire [319:0] set1,
  input wire [319:0] set2,
  output wire [647:0] out
);
  wire [15:0] set1_unflattened[20];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  wire [15:0] set2_unflattened[20];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  wire [15:0] array_index_38821;
  wire [15:0] array_index_38822;
  wire [15:0] array_index_38826;
  wire [1:0] concat_38827;
  wire [1:0] add_38830;
  wire [15:0] array_index_38834;
  wire [2:0] concat_38835;
  wire [2:0] add_38838;
  wire [15:0] array_index_38842;
  wire [3:0] concat_38843;
  wire [3:0] add_38846;
  wire [15:0] array_index_38850;
  wire [4:0] concat_38851;
  wire [4:0] add_38854;
  wire [15:0] array_index_38858;
  wire [5:0] concat_38859;
  wire [5:0] add_38862;
  wire [15:0] array_index_38866;
  wire [6:0] concat_38867;
  wire [6:0] add_38870;
  wire [15:0] array_index_38874;
  wire [7:0] concat_38875;
  wire [7:0] add_38879;
  wire [15:0] array_index_38880;
  wire [7:0] sel_38881;
  wire [7:0] add_38885;
  wire [15:0] array_index_38886;
  wire [7:0] sel_38887;
  wire [7:0] add_38891;
  wire [15:0] array_index_38892;
  wire [7:0] sel_38893;
  wire [7:0] add_38897;
  wire [15:0] array_index_38898;
  wire [7:0] sel_38899;
  wire [7:0] add_38903;
  wire [15:0] array_index_38904;
  wire [7:0] sel_38905;
  wire [7:0] add_38909;
  wire [15:0] array_index_38910;
  wire [7:0] sel_38911;
  wire [7:0] add_38915;
  wire [15:0] array_index_38916;
  wire [7:0] sel_38917;
  wire [7:0] add_38921;
  wire [15:0] array_index_38922;
  wire [7:0] sel_38923;
  wire [7:0] add_38927;
  wire [15:0] array_index_38928;
  wire [7:0] sel_38929;
  wire [7:0] add_38933;
  wire [15:0] array_index_38934;
  wire [7:0] sel_38935;
  wire [7:0] add_38939;
  wire [15:0] array_index_38940;
  wire [7:0] sel_38941;
  wire [7:0] add_38945;
  wire [15:0] array_index_38946;
  wire [7:0] sel_38947;
  wire [7:0] add_38951;
  wire [15:0] array_index_38952;
  wire [7:0] sel_38953;
  wire [7:0] add_38956;
  wire [7:0] sel_38957;
  wire [7:0] add_38960;
  wire [7:0] sel_38961;
  wire [7:0] add_38964;
  wire [7:0] sel_38965;
  wire [7:0] add_38968;
  wire [7:0] sel_38969;
  wire [7:0] add_38972;
  wire [7:0] sel_38973;
  wire [7:0] add_38976;
  wire [7:0] sel_38977;
  wire [7:0] add_38980;
  wire [7:0] sel_38981;
  wire [7:0] add_38984;
  wire [7:0] sel_38985;
  wire [7:0] add_38988;
  wire [7:0] sel_38989;
  wire [7:0] add_38992;
  wire [7:0] sel_38993;
  wire [7:0] add_38996;
  wire [7:0] sel_38997;
  wire [7:0] add_39000;
  wire [7:0] sel_39001;
  wire [7:0] add_39004;
  wire [7:0] sel_39005;
  wire [7:0] add_39008;
  wire [7:0] sel_39009;
  wire [7:0] add_39012;
  wire [7:0] sel_39013;
  wire [7:0] add_39016;
  wire [7:0] sel_39017;
  wire [7:0] add_39020;
  wire [7:0] sel_39021;
  wire [7:0] add_39024;
  wire [7:0] sel_39025;
  wire [7:0] add_39028;
  wire [7:0] sel_39029;
  wire [7:0] add_39033;
  wire [15:0] array_index_39034;
  wire [7:0] sel_39035;
  wire [7:0] add_39038;
  wire [7:0] sel_39039;
  wire [7:0] add_39042;
  wire [7:0] sel_39043;
  wire [7:0] add_39046;
  wire [7:0] sel_39047;
  wire [7:0] add_39050;
  wire [7:0] sel_39051;
  wire [7:0] add_39054;
  wire [7:0] sel_39055;
  wire [7:0] add_39058;
  wire [7:0] sel_39059;
  wire [7:0] add_39062;
  wire [7:0] sel_39063;
  wire [7:0] add_39066;
  wire [7:0] sel_39067;
  wire [7:0] add_39070;
  wire [7:0] sel_39071;
  wire [7:0] add_39074;
  wire [7:0] sel_39075;
  wire [7:0] add_39078;
  wire [7:0] sel_39079;
  wire [7:0] add_39082;
  wire [7:0] sel_39083;
  wire [7:0] add_39086;
  wire [7:0] sel_39087;
  wire [7:0] add_39090;
  wire [7:0] sel_39091;
  wire [7:0] add_39094;
  wire [7:0] sel_39095;
  wire [7:0] add_39098;
  wire [7:0] sel_39099;
  wire [7:0] add_39102;
  wire [7:0] sel_39103;
  wire [7:0] add_39106;
  wire [7:0] sel_39107;
  wire [7:0] add_39110;
  wire [7:0] sel_39111;
  wire [7:0] add_39115;
  wire [15:0] array_index_39116;
  wire [7:0] sel_39117;
  wire [7:0] add_39120;
  wire [7:0] sel_39121;
  wire [7:0] add_39124;
  wire [7:0] sel_39125;
  wire [7:0] add_39128;
  wire [7:0] sel_39129;
  wire [7:0] add_39132;
  wire [7:0] sel_39133;
  wire [7:0] add_39136;
  wire [7:0] sel_39137;
  wire [7:0] add_39140;
  wire [7:0] sel_39141;
  wire [7:0] add_39144;
  wire [7:0] sel_39145;
  wire [7:0] add_39148;
  wire [7:0] sel_39149;
  wire [7:0] add_39152;
  wire [7:0] sel_39153;
  wire [7:0] add_39156;
  wire [7:0] sel_39157;
  wire [7:0] add_39160;
  wire [7:0] sel_39161;
  wire [7:0] add_39164;
  wire [7:0] sel_39165;
  wire [7:0] add_39168;
  wire [7:0] sel_39169;
  wire [7:0] add_39172;
  wire [7:0] sel_39173;
  wire [7:0] add_39176;
  wire [7:0] sel_39177;
  wire [7:0] add_39180;
  wire [7:0] sel_39181;
  wire [7:0] add_39184;
  wire [7:0] sel_39185;
  wire [7:0] add_39188;
  wire [7:0] sel_39189;
  wire [7:0] add_39192;
  wire [7:0] sel_39193;
  wire [7:0] add_39197;
  wire [15:0] array_index_39198;
  wire [7:0] sel_39199;
  wire [7:0] add_39202;
  wire [7:0] sel_39203;
  wire [7:0] add_39206;
  wire [7:0] sel_39207;
  wire [7:0] add_39210;
  wire [7:0] sel_39211;
  wire [7:0] add_39214;
  wire [7:0] sel_39215;
  wire [7:0] add_39218;
  wire [7:0] sel_39219;
  wire [7:0] add_39222;
  wire [7:0] sel_39223;
  wire [7:0] add_39226;
  wire [7:0] sel_39227;
  wire [7:0] add_39230;
  wire [7:0] sel_39231;
  wire [7:0] add_39234;
  wire [7:0] sel_39235;
  wire [7:0] add_39238;
  wire [7:0] sel_39239;
  wire [7:0] add_39242;
  wire [7:0] sel_39243;
  wire [7:0] add_39246;
  wire [7:0] sel_39247;
  wire [7:0] add_39250;
  wire [7:0] sel_39251;
  wire [7:0] add_39254;
  wire [7:0] sel_39255;
  wire [7:0] add_39258;
  wire [7:0] sel_39259;
  wire [7:0] add_39262;
  wire [7:0] sel_39263;
  wire [7:0] add_39266;
  wire [7:0] sel_39267;
  wire [7:0] add_39270;
  wire [7:0] sel_39271;
  wire [7:0] add_39274;
  wire [7:0] sel_39275;
  wire [7:0] add_39279;
  wire [15:0] array_index_39280;
  wire [7:0] sel_39281;
  wire [7:0] add_39284;
  wire [7:0] sel_39285;
  wire [7:0] add_39288;
  wire [7:0] sel_39289;
  wire [7:0] add_39292;
  wire [7:0] sel_39293;
  wire [7:0] add_39296;
  wire [7:0] sel_39297;
  wire [7:0] add_39300;
  wire [7:0] sel_39301;
  wire [7:0] add_39304;
  wire [7:0] sel_39305;
  wire [7:0] add_39308;
  wire [7:0] sel_39309;
  wire [7:0] add_39312;
  wire [7:0] sel_39313;
  wire [7:0] add_39316;
  wire [7:0] sel_39317;
  wire [7:0] add_39320;
  wire [7:0] sel_39321;
  wire [7:0] add_39324;
  wire [7:0] sel_39325;
  wire [7:0] add_39328;
  wire [7:0] sel_39329;
  wire [7:0] add_39332;
  wire [7:0] sel_39333;
  wire [7:0] add_39336;
  wire [7:0] sel_39337;
  wire [7:0] add_39340;
  wire [7:0] sel_39341;
  wire [7:0] add_39344;
  wire [7:0] sel_39345;
  wire [7:0] add_39348;
  wire [7:0] sel_39349;
  wire [7:0] add_39352;
  wire [7:0] sel_39353;
  wire [7:0] add_39356;
  wire [7:0] sel_39357;
  wire [7:0] add_39361;
  wire [15:0] array_index_39362;
  wire [7:0] sel_39363;
  wire [7:0] add_39366;
  wire [7:0] sel_39367;
  wire [7:0] add_39370;
  wire [7:0] sel_39371;
  wire [7:0] add_39374;
  wire [7:0] sel_39375;
  wire [7:0] add_39378;
  wire [7:0] sel_39379;
  wire [7:0] add_39382;
  wire [7:0] sel_39383;
  wire [7:0] add_39386;
  wire [7:0] sel_39387;
  wire [7:0] add_39390;
  wire [7:0] sel_39391;
  wire [7:0] add_39394;
  wire [7:0] sel_39395;
  wire [7:0] add_39398;
  wire [7:0] sel_39399;
  wire [7:0] add_39402;
  wire [7:0] sel_39403;
  wire [7:0] add_39406;
  wire [7:0] sel_39407;
  wire [7:0] add_39410;
  wire [7:0] sel_39411;
  wire [7:0] add_39414;
  wire [7:0] sel_39415;
  wire [7:0] add_39418;
  wire [7:0] sel_39419;
  wire [7:0] add_39422;
  wire [7:0] sel_39423;
  wire [7:0] add_39426;
  wire [7:0] sel_39427;
  wire [7:0] add_39430;
  wire [7:0] sel_39431;
  wire [7:0] add_39434;
  wire [7:0] sel_39435;
  wire [7:0] add_39438;
  wire [7:0] sel_39439;
  wire [7:0] add_39443;
  wire [15:0] array_index_39444;
  wire [7:0] sel_39445;
  wire [7:0] add_39448;
  wire [7:0] sel_39449;
  wire [7:0] add_39452;
  wire [7:0] sel_39453;
  wire [7:0] add_39456;
  wire [7:0] sel_39457;
  wire [7:0] add_39460;
  wire [7:0] sel_39461;
  wire [7:0] add_39464;
  wire [7:0] sel_39465;
  wire [7:0] add_39468;
  wire [7:0] sel_39469;
  wire [7:0] add_39472;
  wire [7:0] sel_39473;
  wire [7:0] add_39476;
  wire [7:0] sel_39477;
  wire [7:0] add_39480;
  wire [7:0] sel_39481;
  wire [7:0] add_39484;
  wire [7:0] sel_39485;
  wire [7:0] add_39488;
  wire [7:0] sel_39489;
  wire [7:0] add_39492;
  wire [7:0] sel_39493;
  wire [7:0] add_39496;
  wire [7:0] sel_39497;
  wire [7:0] add_39500;
  wire [7:0] sel_39501;
  wire [7:0] add_39504;
  wire [7:0] sel_39505;
  wire [7:0] add_39508;
  wire [7:0] sel_39509;
  wire [7:0] add_39512;
  wire [7:0] sel_39513;
  wire [7:0] add_39516;
  wire [7:0] sel_39517;
  wire [7:0] add_39520;
  wire [7:0] sel_39521;
  wire [7:0] add_39525;
  wire [15:0] array_index_39526;
  wire [7:0] sel_39527;
  wire [7:0] add_39530;
  wire [7:0] sel_39531;
  wire [7:0] add_39534;
  wire [7:0] sel_39535;
  wire [7:0] add_39538;
  wire [7:0] sel_39539;
  wire [7:0] add_39542;
  wire [7:0] sel_39543;
  wire [7:0] add_39546;
  wire [7:0] sel_39547;
  wire [7:0] add_39550;
  wire [7:0] sel_39551;
  wire [7:0] add_39554;
  wire [7:0] sel_39555;
  wire [7:0] add_39558;
  wire [7:0] sel_39559;
  wire [7:0] add_39562;
  wire [7:0] sel_39563;
  wire [7:0] add_39566;
  wire [7:0] sel_39567;
  wire [7:0] add_39570;
  wire [7:0] sel_39571;
  wire [7:0] add_39574;
  wire [7:0] sel_39575;
  wire [7:0] add_39578;
  wire [7:0] sel_39579;
  wire [7:0] add_39582;
  wire [7:0] sel_39583;
  wire [7:0] add_39586;
  wire [7:0] sel_39587;
  wire [7:0] add_39590;
  wire [7:0] sel_39591;
  wire [7:0] add_39594;
  wire [7:0] sel_39595;
  wire [7:0] add_39598;
  wire [7:0] sel_39599;
  wire [7:0] add_39602;
  wire [7:0] sel_39603;
  wire [7:0] add_39607;
  wire [15:0] array_index_39608;
  wire [7:0] sel_39609;
  wire [7:0] add_39612;
  wire [7:0] sel_39613;
  wire [7:0] add_39616;
  wire [7:0] sel_39617;
  wire [7:0] add_39620;
  wire [7:0] sel_39621;
  wire [7:0] add_39624;
  wire [7:0] sel_39625;
  wire [7:0] add_39628;
  wire [7:0] sel_39629;
  wire [7:0] add_39632;
  wire [7:0] sel_39633;
  wire [7:0] add_39636;
  wire [7:0] sel_39637;
  wire [7:0] add_39640;
  wire [7:0] sel_39641;
  wire [7:0] add_39644;
  wire [7:0] sel_39645;
  wire [7:0] add_39648;
  wire [7:0] sel_39649;
  wire [7:0] add_39652;
  wire [7:0] sel_39653;
  wire [7:0] add_39656;
  wire [7:0] sel_39657;
  wire [7:0] add_39660;
  wire [7:0] sel_39661;
  wire [7:0] add_39664;
  wire [7:0] sel_39665;
  wire [7:0] add_39668;
  wire [7:0] sel_39669;
  wire [7:0] add_39672;
  wire [7:0] sel_39673;
  wire [7:0] add_39676;
  wire [7:0] sel_39677;
  wire [7:0] add_39680;
  wire [7:0] sel_39681;
  wire [7:0] add_39684;
  wire [7:0] sel_39685;
  wire [7:0] add_39689;
  wire [15:0] array_index_39690;
  wire [7:0] sel_39691;
  wire [7:0] add_39694;
  wire [7:0] sel_39695;
  wire [7:0] add_39698;
  wire [7:0] sel_39699;
  wire [7:0] add_39702;
  wire [7:0] sel_39703;
  wire [7:0] add_39706;
  wire [7:0] sel_39707;
  wire [7:0] add_39710;
  wire [7:0] sel_39711;
  wire [7:0] add_39714;
  wire [7:0] sel_39715;
  wire [7:0] add_39718;
  wire [7:0] sel_39719;
  wire [7:0] add_39722;
  wire [7:0] sel_39723;
  wire [7:0] add_39726;
  wire [7:0] sel_39727;
  wire [7:0] add_39730;
  wire [7:0] sel_39731;
  wire [7:0] add_39734;
  wire [7:0] sel_39735;
  wire [7:0] add_39738;
  wire [7:0] sel_39739;
  wire [7:0] add_39742;
  wire [7:0] sel_39743;
  wire [7:0] add_39746;
  wire [7:0] sel_39747;
  wire [7:0] add_39750;
  wire [7:0] sel_39751;
  wire [7:0] add_39754;
  wire [7:0] sel_39755;
  wire [7:0] add_39758;
  wire [7:0] sel_39759;
  wire [7:0] add_39762;
  wire [7:0] sel_39763;
  wire [7:0] add_39766;
  wire [7:0] sel_39767;
  wire [7:0] add_39771;
  wire [15:0] array_index_39772;
  wire [7:0] sel_39773;
  wire [7:0] add_39776;
  wire [7:0] sel_39777;
  wire [7:0] add_39780;
  wire [7:0] sel_39781;
  wire [7:0] add_39784;
  wire [7:0] sel_39785;
  wire [7:0] add_39788;
  wire [7:0] sel_39789;
  wire [7:0] add_39792;
  wire [7:0] sel_39793;
  wire [7:0] add_39796;
  wire [7:0] sel_39797;
  wire [7:0] add_39800;
  wire [7:0] sel_39801;
  wire [7:0] add_39804;
  wire [7:0] sel_39805;
  wire [7:0] add_39808;
  wire [7:0] sel_39809;
  wire [7:0] add_39812;
  wire [7:0] sel_39813;
  wire [7:0] add_39816;
  wire [7:0] sel_39817;
  wire [7:0] add_39820;
  wire [7:0] sel_39821;
  wire [7:0] add_39824;
  wire [7:0] sel_39825;
  wire [7:0] add_39828;
  wire [7:0] sel_39829;
  wire [7:0] add_39832;
  wire [7:0] sel_39833;
  wire [7:0] add_39836;
  wire [7:0] sel_39837;
  wire [7:0] add_39840;
  wire [7:0] sel_39841;
  wire [7:0] add_39844;
  wire [7:0] sel_39845;
  wire [7:0] add_39848;
  wire [7:0] sel_39849;
  wire [7:0] add_39853;
  wire [15:0] array_index_39854;
  wire [7:0] sel_39855;
  wire [7:0] add_39858;
  wire [7:0] sel_39859;
  wire [7:0] add_39862;
  wire [7:0] sel_39863;
  wire [7:0] add_39866;
  wire [7:0] sel_39867;
  wire [7:0] add_39870;
  wire [7:0] sel_39871;
  wire [7:0] add_39874;
  wire [7:0] sel_39875;
  wire [7:0] add_39878;
  wire [7:0] sel_39879;
  wire [7:0] add_39882;
  wire [7:0] sel_39883;
  wire [7:0] add_39886;
  wire [7:0] sel_39887;
  wire [7:0] add_39890;
  wire [7:0] sel_39891;
  wire [7:0] add_39894;
  wire [7:0] sel_39895;
  wire [7:0] add_39898;
  wire [7:0] sel_39899;
  wire [7:0] add_39902;
  wire [7:0] sel_39903;
  wire [7:0] add_39906;
  wire [7:0] sel_39907;
  wire [7:0] add_39910;
  wire [7:0] sel_39911;
  wire [7:0] add_39914;
  wire [7:0] sel_39915;
  wire [7:0] add_39918;
  wire [7:0] sel_39919;
  wire [7:0] add_39922;
  wire [7:0] sel_39923;
  wire [7:0] add_39926;
  wire [7:0] sel_39927;
  wire [7:0] add_39930;
  wire [7:0] sel_39931;
  wire [7:0] add_39935;
  wire [15:0] array_index_39936;
  wire [7:0] sel_39937;
  wire [7:0] add_39940;
  wire [7:0] sel_39941;
  wire [7:0] add_39944;
  wire [7:0] sel_39945;
  wire [7:0] add_39948;
  wire [7:0] sel_39949;
  wire [7:0] add_39952;
  wire [7:0] sel_39953;
  wire [7:0] add_39956;
  wire [7:0] sel_39957;
  wire [7:0] add_39960;
  wire [7:0] sel_39961;
  wire [7:0] add_39964;
  wire [7:0] sel_39965;
  wire [7:0] add_39968;
  wire [7:0] sel_39969;
  wire [7:0] add_39972;
  wire [7:0] sel_39973;
  wire [7:0] add_39976;
  wire [7:0] sel_39977;
  wire [7:0] add_39980;
  wire [7:0] sel_39981;
  wire [7:0] add_39984;
  wire [7:0] sel_39985;
  wire [7:0] add_39988;
  wire [7:0] sel_39989;
  wire [7:0] add_39992;
  wire [7:0] sel_39993;
  wire [7:0] add_39996;
  wire [7:0] sel_39997;
  wire [7:0] add_40000;
  wire [7:0] sel_40001;
  wire [7:0] add_40004;
  wire [7:0] sel_40005;
  wire [7:0] add_40008;
  wire [7:0] sel_40009;
  wire [7:0] add_40012;
  wire [7:0] sel_40013;
  wire [7:0] add_40017;
  wire [15:0] array_index_40018;
  wire [7:0] sel_40019;
  wire [7:0] add_40022;
  wire [7:0] sel_40023;
  wire [7:0] add_40026;
  wire [7:0] sel_40027;
  wire [7:0] add_40030;
  wire [7:0] sel_40031;
  wire [7:0] add_40034;
  wire [7:0] sel_40035;
  wire [7:0] add_40038;
  wire [7:0] sel_40039;
  wire [7:0] add_40042;
  wire [7:0] sel_40043;
  wire [7:0] add_40046;
  wire [7:0] sel_40047;
  wire [7:0] add_40050;
  wire [7:0] sel_40051;
  wire [7:0] add_40054;
  wire [7:0] sel_40055;
  wire [7:0] add_40058;
  wire [7:0] sel_40059;
  wire [7:0] add_40062;
  wire [7:0] sel_40063;
  wire [7:0] add_40066;
  wire [7:0] sel_40067;
  wire [7:0] add_40070;
  wire [7:0] sel_40071;
  wire [7:0] add_40074;
  wire [7:0] sel_40075;
  wire [7:0] add_40078;
  wire [7:0] sel_40079;
  wire [7:0] add_40082;
  wire [7:0] sel_40083;
  wire [7:0] add_40086;
  wire [7:0] sel_40087;
  wire [7:0] add_40090;
  wire [7:0] sel_40091;
  wire [7:0] add_40094;
  wire [7:0] sel_40095;
  wire [7:0] add_40099;
  wire [15:0] array_index_40100;
  wire [7:0] sel_40101;
  wire [7:0] add_40104;
  wire [7:0] sel_40105;
  wire [7:0] add_40108;
  wire [7:0] sel_40109;
  wire [7:0] add_40112;
  wire [7:0] sel_40113;
  wire [7:0] add_40116;
  wire [7:0] sel_40117;
  wire [7:0] add_40120;
  wire [7:0] sel_40121;
  wire [7:0] add_40124;
  wire [7:0] sel_40125;
  wire [7:0] add_40128;
  wire [7:0] sel_40129;
  wire [7:0] add_40132;
  wire [7:0] sel_40133;
  wire [7:0] add_40136;
  wire [7:0] sel_40137;
  wire [7:0] add_40140;
  wire [7:0] sel_40141;
  wire [7:0] add_40144;
  wire [7:0] sel_40145;
  wire [7:0] add_40148;
  wire [7:0] sel_40149;
  wire [7:0] add_40152;
  wire [7:0] sel_40153;
  wire [7:0] add_40156;
  wire [7:0] sel_40157;
  wire [7:0] add_40160;
  wire [7:0] sel_40161;
  wire [7:0] add_40164;
  wire [7:0] sel_40165;
  wire [7:0] add_40168;
  wire [7:0] sel_40169;
  wire [7:0] add_40172;
  wire [7:0] sel_40173;
  wire [7:0] add_40176;
  wire [7:0] sel_40177;
  wire [7:0] add_40181;
  wire [15:0] array_index_40182;
  wire [7:0] sel_40183;
  wire [7:0] add_40186;
  wire [7:0] sel_40187;
  wire [7:0] add_40190;
  wire [7:0] sel_40191;
  wire [7:0] add_40194;
  wire [7:0] sel_40195;
  wire [7:0] add_40198;
  wire [7:0] sel_40199;
  wire [7:0] add_40202;
  wire [7:0] sel_40203;
  wire [7:0] add_40206;
  wire [7:0] sel_40207;
  wire [7:0] add_40210;
  wire [7:0] sel_40211;
  wire [7:0] add_40214;
  wire [7:0] sel_40215;
  wire [7:0] add_40218;
  wire [7:0] sel_40219;
  wire [7:0] add_40222;
  wire [7:0] sel_40223;
  wire [7:0] add_40226;
  wire [7:0] sel_40227;
  wire [7:0] add_40230;
  wire [7:0] sel_40231;
  wire [7:0] add_40234;
  wire [7:0] sel_40235;
  wire [7:0] add_40238;
  wire [7:0] sel_40239;
  wire [7:0] add_40242;
  wire [7:0] sel_40243;
  wire [7:0] add_40246;
  wire [7:0] sel_40247;
  wire [7:0] add_40250;
  wire [7:0] sel_40251;
  wire [7:0] add_40254;
  wire [7:0] sel_40255;
  wire [7:0] add_40258;
  wire [7:0] sel_40259;
  wire [7:0] add_40263;
  wire [15:0] array_index_40264;
  wire [7:0] sel_40265;
  wire [7:0] add_40268;
  wire [7:0] sel_40269;
  wire [7:0] add_40272;
  wire [7:0] sel_40273;
  wire [7:0] add_40276;
  wire [7:0] sel_40277;
  wire [7:0] add_40280;
  wire [7:0] sel_40281;
  wire [7:0] add_40284;
  wire [7:0] sel_40285;
  wire [7:0] add_40288;
  wire [7:0] sel_40289;
  wire [7:0] add_40292;
  wire [7:0] sel_40293;
  wire [7:0] add_40296;
  wire [7:0] sel_40297;
  wire [7:0] add_40300;
  wire [7:0] sel_40301;
  wire [7:0] add_40304;
  wire [7:0] sel_40305;
  wire [7:0] add_40308;
  wire [7:0] sel_40309;
  wire [7:0] add_40312;
  wire [7:0] sel_40313;
  wire [7:0] add_40316;
  wire [7:0] sel_40317;
  wire [7:0] add_40320;
  wire [7:0] sel_40321;
  wire [7:0] add_40324;
  wire [7:0] sel_40325;
  wire [7:0] add_40328;
  wire [7:0] sel_40329;
  wire [7:0] add_40332;
  wire [7:0] sel_40333;
  wire [7:0] add_40336;
  wire [7:0] sel_40337;
  wire [7:0] add_40340;
  wire [7:0] sel_40341;
  wire [7:0] add_40345;
  wire [15:0] array_index_40346;
  wire [7:0] sel_40347;
  wire [7:0] add_40350;
  wire [7:0] sel_40351;
  wire [7:0] add_40354;
  wire [7:0] sel_40355;
  wire [7:0] add_40358;
  wire [7:0] sel_40359;
  wire [7:0] add_40362;
  wire [7:0] sel_40363;
  wire [7:0] add_40366;
  wire [7:0] sel_40367;
  wire [7:0] add_40370;
  wire [7:0] sel_40371;
  wire [7:0] add_40374;
  wire [7:0] sel_40375;
  wire [7:0] add_40378;
  wire [7:0] sel_40379;
  wire [7:0] add_40382;
  wire [7:0] sel_40383;
  wire [7:0] add_40386;
  wire [7:0] sel_40387;
  wire [7:0] add_40390;
  wire [7:0] sel_40391;
  wire [7:0] add_40394;
  wire [7:0] sel_40395;
  wire [7:0] add_40398;
  wire [7:0] sel_40399;
  wire [7:0] add_40402;
  wire [7:0] sel_40403;
  wire [7:0] add_40406;
  wire [7:0] sel_40407;
  wire [7:0] add_40410;
  wire [7:0] sel_40411;
  wire [7:0] add_40414;
  wire [7:0] sel_40415;
  wire [7:0] add_40418;
  wire [7:0] sel_40419;
  wire [7:0] add_40422;
  wire [7:0] sel_40423;
  wire [7:0] add_40427;
  wire [15:0] array_index_40428;
  wire [7:0] sel_40429;
  wire [7:0] add_40432;
  wire [7:0] sel_40433;
  wire [7:0] add_40436;
  wire [7:0] sel_40437;
  wire [7:0] add_40440;
  wire [7:0] sel_40441;
  wire [7:0] add_40444;
  wire [7:0] sel_40445;
  wire [7:0] add_40448;
  wire [7:0] sel_40449;
  wire [7:0] add_40452;
  wire [7:0] sel_40453;
  wire [7:0] add_40456;
  wire [7:0] sel_40457;
  wire [7:0] add_40460;
  wire [7:0] sel_40461;
  wire [7:0] add_40464;
  wire [7:0] sel_40465;
  wire [7:0] add_40468;
  wire [7:0] sel_40469;
  wire [7:0] add_40472;
  wire [7:0] sel_40473;
  wire [7:0] add_40476;
  wire [7:0] sel_40477;
  wire [7:0] add_40480;
  wire [7:0] sel_40481;
  wire [7:0] add_40484;
  wire [7:0] sel_40485;
  wire [7:0] add_40488;
  wire [7:0] sel_40489;
  wire [7:0] add_40492;
  wire [7:0] sel_40493;
  wire [7:0] add_40496;
  wire [7:0] sel_40497;
  wire [7:0] add_40500;
  wire [7:0] sel_40501;
  wire [7:0] add_40504;
  wire [7:0] sel_40505;
  wire [7:0] add_40508;
  assign array_index_38821 = set1_unflattened[5'h00];
  assign array_index_38822 = set2_unflattened[5'h00];
  assign array_index_38826 = set2_unflattened[5'h01];
  assign concat_38827 = {1'h0, array_index_38821 == array_index_38822};
  assign add_38830 = concat_38827 + 2'h1;
  assign array_index_38834 = set2_unflattened[5'h02];
  assign concat_38835 = {1'h0, array_index_38821 == array_index_38826 ? add_38830 : concat_38827};
  assign add_38838 = concat_38835 + 3'h1;
  assign array_index_38842 = set2_unflattened[5'h03];
  assign concat_38843 = {1'h0, array_index_38821 == array_index_38834 ? add_38838 : concat_38835};
  assign add_38846 = concat_38843 + 4'h1;
  assign array_index_38850 = set2_unflattened[5'h04];
  assign concat_38851 = {1'h0, array_index_38821 == array_index_38842 ? add_38846 : concat_38843};
  assign add_38854 = concat_38851 + 5'h01;
  assign array_index_38858 = set2_unflattened[5'h05];
  assign concat_38859 = {1'h0, array_index_38821 == array_index_38850 ? add_38854 : concat_38851};
  assign add_38862 = concat_38859 + 6'h01;
  assign array_index_38866 = set2_unflattened[5'h06];
  assign concat_38867 = {1'h0, array_index_38821 == array_index_38858 ? add_38862 : concat_38859};
  assign add_38870 = concat_38867 + 7'h01;
  assign array_index_38874 = set2_unflattened[5'h07];
  assign concat_38875 = {1'h0, array_index_38821 == array_index_38866 ? add_38870 : concat_38867};
  assign add_38879 = concat_38875 + 8'h01;
  assign array_index_38880 = set2_unflattened[5'h08];
  assign sel_38881 = array_index_38821 == array_index_38874 ? add_38879 : concat_38875;
  assign add_38885 = sel_38881 + 8'h01;
  assign array_index_38886 = set2_unflattened[5'h09];
  assign sel_38887 = array_index_38821 == array_index_38880 ? add_38885 : sel_38881;
  assign add_38891 = sel_38887 + 8'h01;
  assign array_index_38892 = set2_unflattened[5'h0a];
  assign sel_38893 = array_index_38821 == array_index_38886 ? add_38891 : sel_38887;
  assign add_38897 = sel_38893 + 8'h01;
  assign array_index_38898 = set2_unflattened[5'h0b];
  assign sel_38899 = array_index_38821 == array_index_38892 ? add_38897 : sel_38893;
  assign add_38903 = sel_38899 + 8'h01;
  assign array_index_38904 = set2_unflattened[5'h0c];
  assign sel_38905 = array_index_38821 == array_index_38898 ? add_38903 : sel_38899;
  assign add_38909 = sel_38905 + 8'h01;
  assign array_index_38910 = set2_unflattened[5'h0d];
  assign sel_38911 = array_index_38821 == array_index_38904 ? add_38909 : sel_38905;
  assign add_38915 = sel_38911 + 8'h01;
  assign array_index_38916 = set2_unflattened[5'h0e];
  assign sel_38917 = array_index_38821 == array_index_38910 ? add_38915 : sel_38911;
  assign add_38921 = sel_38917 + 8'h01;
  assign array_index_38922 = set2_unflattened[5'h0f];
  assign sel_38923 = array_index_38821 == array_index_38916 ? add_38921 : sel_38917;
  assign add_38927 = sel_38923 + 8'h01;
  assign array_index_38928 = set2_unflattened[5'h10];
  assign sel_38929 = array_index_38821 == array_index_38922 ? add_38927 : sel_38923;
  assign add_38933 = sel_38929 + 8'h01;
  assign array_index_38934 = set2_unflattened[5'h11];
  assign sel_38935 = array_index_38821 == array_index_38928 ? add_38933 : sel_38929;
  assign add_38939 = sel_38935 + 8'h01;
  assign array_index_38940 = set2_unflattened[5'h12];
  assign sel_38941 = array_index_38821 == array_index_38934 ? add_38939 : sel_38935;
  assign add_38945 = sel_38941 + 8'h01;
  assign array_index_38946 = set2_unflattened[5'h13];
  assign sel_38947 = array_index_38821 == array_index_38940 ? add_38945 : sel_38941;
  assign add_38951 = sel_38947 + 8'h01;
  assign array_index_38952 = set1_unflattened[5'h01];
  assign sel_38953 = array_index_38821 == array_index_38946 ? add_38951 : sel_38947;
  assign add_38956 = sel_38953 + 8'h01;
  assign sel_38957 = array_index_38952 == array_index_38822 ? add_38956 : sel_38953;
  assign add_38960 = sel_38957 + 8'h01;
  assign sel_38961 = array_index_38952 == array_index_38826 ? add_38960 : sel_38957;
  assign add_38964 = sel_38961 + 8'h01;
  assign sel_38965 = array_index_38952 == array_index_38834 ? add_38964 : sel_38961;
  assign add_38968 = sel_38965 + 8'h01;
  assign sel_38969 = array_index_38952 == array_index_38842 ? add_38968 : sel_38965;
  assign add_38972 = sel_38969 + 8'h01;
  assign sel_38973 = array_index_38952 == array_index_38850 ? add_38972 : sel_38969;
  assign add_38976 = sel_38973 + 8'h01;
  assign sel_38977 = array_index_38952 == array_index_38858 ? add_38976 : sel_38973;
  assign add_38980 = sel_38977 + 8'h01;
  assign sel_38981 = array_index_38952 == array_index_38866 ? add_38980 : sel_38977;
  assign add_38984 = sel_38981 + 8'h01;
  assign sel_38985 = array_index_38952 == array_index_38874 ? add_38984 : sel_38981;
  assign add_38988 = sel_38985 + 8'h01;
  assign sel_38989 = array_index_38952 == array_index_38880 ? add_38988 : sel_38985;
  assign add_38992 = sel_38989 + 8'h01;
  assign sel_38993 = array_index_38952 == array_index_38886 ? add_38992 : sel_38989;
  assign add_38996 = sel_38993 + 8'h01;
  assign sel_38997 = array_index_38952 == array_index_38892 ? add_38996 : sel_38993;
  assign add_39000 = sel_38997 + 8'h01;
  assign sel_39001 = array_index_38952 == array_index_38898 ? add_39000 : sel_38997;
  assign add_39004 = sel_39001 + 8'h01;
  assign sel_39005 = array_index_38952 == array_index_38904 ? add_39004 : sel_39001;
  assign add_39008 = sel_39005 + 8'h01;
  assign sel_39009 = array_index_38952 == array_index_38910 ? add_39008 : sel_39005;
  assign add_39012 = sel_39009 + 8'h01;
  assign sel_39013 = array_index_38952 == array_index_38916 ? add_39012 : sel_39009;
  assign add_39016 = sel_39013 + 8'h01;
  assign sel_39017 = array_index_38952 == array_index_38922 ? add_39016 : sel_39013;
  assign add_39020 = sel_39017 + 8'h01;
  assign sel_39021 = array_index_38952 == array_index_38928 ? add_39020 : sel_39017;
  assign add_39024 = sel_39021 + 8'h01;
  assign sel_39025 = array_index_38952 == array_index_38934 ? add_39024 : sel_39021;
  assign add_39028 = sel_39025 + 8'h01;
  assign sel_39029 = array_index_38952 == array_index_38940 ? add_39028 : sel_39025;
  assign add_39033 = sel_39029 + 8'h01;
  assign array_index_39034 = set1_unflattened[5'h02];
  assign sel_39035 = array_index_38952 == array_index_38946 ? add_39033 : sel_39029;
  assign add_39038 = sel_39035 + 8'h01;
  assign sel_39039 = array_index_39034 == array_index_38822 ? add_39038 : sel_39035;
  assign add_39042 = sel_39039 + 8'h01;
  assign sel_39043 = array_index_39034 == array_index_38826 ? add_39042 : sel_39039;
  assign add_39046 = sel_39043 + 8'h01;
  assign sel_39047 = array_index_39034 == array_index_38834 ? add_39046 : sel_39043;
  assign add_39050 = sel_39047 + 8'h01;
  assign sel_39051 = array_index_39034 == array_index_38842 ? add_39050 : sel_39047;
  assign add_39054 = sel_39051 + 8'h01;
  assign sel_39055 = array_index_39034 == array_index_38850 ? add_39054 : sel_39051;
  assign add_39058 = sel_39055 + 8'h01;
  assign sel_39059 = array_index_39034 == array_index_38858 ? add_39058 : sel_39055;
  assign add_39062 = sel_39059 + 8'h01;
  assign sel_39063 = array_index_39034 == array_index_38866 ? add_39062 : sel_39059;
  assign add_39066 = sel_39063 + 8'h01;
  assign sel_39067 = array_index_39034 == array_index_38874 ? add_39066 : sel_39063;
  assign add_39070 = sel_39067 + 8'h01;
  assign sel_39071 = array_index_39034 == array_index_38880 ? add_39070 : sel_39067;
  assign add_39074 = sel_39071 + 8'h01;
  assign sel_39075 = array_index_39034 == array_index_38886 ? add_39074 : sel_39071;
  assign add_39078 = sel_39075 + 8'h01;
  assign sel_39079 = array_index_39034 == array_index_38892 ? add_39078 : sel_39075;
  assign add_39082 = sel_39079 + 8'h01;
  assign sel_39083 = array_index_39034 == array_index_38898 ? add_39082 : sel_39079;
  assign add_39086 = sel_39083 + 8'h01;
  assign sel_39087 = array_index_39034 == array_index_38904 ? add_39086 : sel_39083;
  assign add_39090 = sel_39087 + 8'h01;
  assign sel_39091 = array_index_39034 == array_index_38910 ? add_39090 : sel_39087;
  assign add_39094 = sel_39091 + 8'h01;
  assign sel_39095 = array_index_39034 == array_index_38916 ? add_39094 : sel_39091;
  assign add_39098 = sel_39095 + 8'h01;
  assign sel_39099 = array_index_39034 == array_index_38922 ? add_39098 : sel_39095;
  assign add_39102 = sel_39099 + 8'h01;
  assign sel_39103 = array_index_39034 == array_index_38928 ? add_39102 : sel_39099;
  assign add_39106 = sel_39103 + 8'h01;
  assign sel_39107 = array_index_39034 == array_index_38934 ? add_39106 : sel_39103;
  assign add_39110 = sel_39107 + 8'h01;
  assign sel_39111 = array_index_39034 == array_index_38940 ? add_39110 : sel_39107;
  assign add_39115 = sel_39111 + 8'h01;
  assign array_index_39116 = set1_unflattened[5'h03];
  assign sel_39117 = array_index_39034 == array_index_38946 ? add_39115 : sel_39111;
  assign add_39120 = sel_39117 + 8'h01;
  assign sel_39121 = array_index_39116 == array_index_38822 ? add_39120 : sel_39117;
  assign add_39124 = sel_39121 + 8'h01;
  assign sel_39125 = array_index_39116 == array_index_38826 ? add_39124 : sel_39121;
  assign add_39128 = sel_39125 + 8'h01;
  assign sel_39129 = array_index_39116 == array_index_38834 ? add_39128 : sel_39125;
  assign add_39132 = sel_39129 + 8'h01;
  assign sel_39133 = array_index_39116 == array_index_38842 ? add_39132 : sel_39129;
  assign add_39136 = sel_39133 + 8'h01;
  assign sel_39137 = array_index_39116 == array_index_38850 ? add_39136 : sel_39133;
  assign add_39140 = sel_39137 + 8'h01;
  assign sel_39141 = array_index_39116 == array_index_38858 ? add_39140 : sel_39137;
  assign add_39144 = sel_39141 + 8'h01;
  assign sel_39145 = array_index_39116 == array_index_38866 ? add_39144 : sel_39141;
  assign add_39148 = sel_39145 + 8'h01;
  assign sel_39149 = array_index_39116 == array_index_38874 ? add_39148 : sel_39145;
  assign add_39152 = sel_39149 + 8'h01;
  assign sel_39153 = array_index_39116 == array_index_38880 ? add_39152 : sel_39149;
  assign add_39156 = sel_39153 + 8'h01;
  assign sel_39157 = array_index_39116 == array_index_38886 ? add_39156 : sel_39153;
  assign add_39160 = sel_39157 + 8'h01;
  assign sel_39161 = array_index_39116 == array_index_38892 ? add_39160 : sel_39157;
  assign add_39164 = sel_39161 + 8'h01;
  assign sel_39165 = array_index_39116 == array_index_38898 ? add_39164 : sel_39161;
  assign add_39168 = sel_39165 + 8'h01;
  assign sel_39169 = array_index_39116 == array_index_38904 ? add_39168 : sel_39165;
  assign add_39172 = sel_39169 + 8'h01;
  assign sel_39173 = array_index_39116 == array_index_38910 ? add_39172 : sel_39169;
  assign add_39176 = sel_39173 + 8'h01;
  assign sel_39177 = array_index_39116 == array_index_38916 ? add_39176 : sel_39173;
  assign add_39180 = sel_39177 + 8'h01;
  assign sel_39181 = array_index_39116 == array_index_38922 ? add_39180 : sel_39177;
  assign add_39184 = sel_39181 + 8'h01;
  assign sel_39185 = array_index_39116 == array_index_38928 ? add_39184 : sel_39181;
  assign add_39188 = sel_39185 + 8'h01;
  assign sel_39189 = array_index_39116 == array_index_38934 ? add_39188 : sel_39185;
  assign add_39192 = sel_39189 + 8'h01;
  assign sel_39193 = array_index_39116 == array_index_38940 ? add_39192 : sel_39189;
  assign add_39197 = sel_39193 + 8'h01;
  assign array_index_39198 = set1_unflattened[5'h04];
  assign sel_39199 = array_index_39116 == array_index_38946 ? add_39197 : sel_39193;
  assign add_39202 = sel_39199 + 8'h01;
  assign sel_39203 = array_index_39198 == array_index_38822 ? add_39202 : sel_39199;
  assign add_39206 = sel_39203 + 8'h01;
  assign sel_39207 = array_index_39198 == array_index_38826 ? add_39206 : sel_39203;
  assign add_39210 = sel_39207 + 8'h01;
  assign sel_39211 = array_index_39198 == array_index_38834 ? add_39210 : sel_39207;
  assign add_39214 = sel_39211 + 8'h01;
  assign sel_39215 = array_index_39198 == array_index_38842 ? add_39214 : sel_39211;
  assign add_39218 = sel_39215 + 8'h01;
  assign sel_39219 = array_index_39198 == array_index_38850 ? add_39218 : sel_39215;
  assign add_39222 = sel_39219 + 8'h01;
  assign sel_39223 = array_index_39198 == array_index_38858 ? add_39222 : sel_39219;
  assign add_39226 = sel_39223 + 8'h01;
  assign sel_39227 = array_index_39198 == array_index_38866 ? add_39226 : sel_39223;
  assign add_39230 = sel_39227 + 8'h01;
  assign sel_39231 = array_index_39198 == array_index_38874 ? add_39230 : sel_39227;
  assign add_39234 = sel_39231 + 8'h01;
  assign sel_39235 = array_index_39198 == array_index_38880 ? add_39234 : sel_39231;
  assign add_39238 = sel_39235 + 8'h01;
  assign sel_39239 = array_index_39198 == array_index_38886 ? add_39238 : sel_39235;
  assign add_39242 = sel_39239 + 8'h01;
  assign sel_39243 = array_index_39198 == array_index_38892 ? add_39242 : sel_39239;
  assign add_39246 = sel_39243 + 8'h01;
  assign sel_39247 = array_index_39198 == array_index_38898 ? add_39246 : sel_39243;
  assign add_39250 = sel_39247 + 8'h01;
  assign sel_39251 = array_index_39198 == array_index_38904 ? add_39250 : sel_39247;
  assign add_39254 = sel_39251 + 8'h01;
  assign sel_39255 = array_index_39198 == array_index_38910 ? add_39254 : sel_39251;
  assign add_39258 = sel_39255 + 8'h01;
  assign sel_39259 = array_index_39198 == array_index_38916 ? add_39258 : sel_39255;
  assign add_39262 = sel_39259 + 8'h01;
  assign sel_39263 = array_index_39198 == array_index_38922 ? add_39262 : sel_39259;
  assign add_39266 = sel_39263 + 8'h01;
  assign sel_39267 = array_index_39198 == array_index_38928 ? add_39266 : sel_39263;
  assign add_39270 = sel_39267 + 8'h01;
  assign sel_39271 = array_index_39198 == array_index_38934 ? add_39270 : sel_39267;
  assign add_39274 = sel_39271 + 8'h01;
  assign sel_39275 = array_index_39198 == array_index_38940 ? add_39274 : sel_39271;
  assign add_39279 = sel_39275 + 8'h01;
  assign array_index_39280 = set1_unflattened[5'h05];
  assign sel_39281 = array_index_39198 == array_index_38946 ? add_39279 : sel_39275;
  assign add_39284 = sel_39281 + 8'h01;
  assign sel_39285 = array_index_39280 == array_index_38822 ? add_39284 : sel_39281;
  assign add_39288 = sel_39285 + 8'h01;
  assign sel_39289 = array_index_39280 == array_index_38826 ? add_39288 : sel_39285;
  assign add_39292 = sel_39289 + 8'h01;
  assign sel_39293 = array_index_39280 == array_index_38834 ? add_39292 : sel_39289;
  assign add_39296 = sel_39293 + 8'h01;
  assign sel_39297 = array_index_39280 == array_index_38842 ? add_39296 : sel_39293;
  assign add_39300 = sel_39297 + 8'h01;
  assign sel_39301 = array_index_39280 == array_index_38850 ? add_39300 : sel_39297;
  assign add_39304 = sel_39301 + 8'h01;
  assign sel_39305 = array_index_39280 == array_index_38858 ? add_39304 : sel_39301;
  assign add_39308 = sel_39305 + 8'h01;
  assign sel_39309 = array_index_39280 == array_index_38866 ? add_39308 : sel_39305;
  assign add_39312 = sel_39309 + 8'h01;
  assign sel_39313 = array_index_39280 == array_index_38874 ? add_39312 : sel_39309;
  assign add_39316 = sel_39313 + 8'h01;
  assign sel_39317 = array_index_39280 == array_index_38880 ? add_39316 : sel_39313;
  assign add_39320 = sel_39317 + 8'h01;
  assign sel_39321 = array_index_39280 == array_index_38886 ? add_39320 : sel_39317;
  assign add_39324 = sel_39321 + 8'h01;
  assign sel_39325 = array_index_39280 == array_index_38892 ? add_39324 : sel_39321;
  assign add_39328 = sel_39325 + 8'h01;
  assign sel_39329 = array_index_39280 == array_index_38898 ? add_39328 : sel_39325;
  assign add_39332 = sel_39329 + 8'h01;
  assign sel_39333 = array_index_39280 == array_index_38904 ? add_39332 : sel_39329;
  assign add_39336 = sel_39333 + 8'h01;
  assign sel_39337 = array_index_39280 == array_index_38910 ? add_39336 : sel_39333;
  assign add_39340 = sel_39337 + 8'h01;
  assign sel_39341 = array_index_39280 == array_index_38916 ? add_39340 : sel_39337;
  assign add_39344 = sel_39341 + 8'h01;
  assign sel_39345 = array_index_39280 == array_index_38922 ? add_39344 : sel_39341;
  assign add_39348 = sel_39345 + 8'h01;
  assign sel_39349 = array_index_39280 == array_index_38928 ? add_39348 : sel_39345;
  assign add_39352 = sel_39349 + 8'h01;
  assign sel_39353 = array_index_39280 == array_index_38934 ? add_39352 : sel_39349;
  assign add_39356 = sel_39353 + 8'h01;
  assign sel_39357 = array_index_39280 == array_index_38940 ? add_39356 : sel_39353;
  assign add_39361 = sel_39357 + 8'h01;
  assign array_index_39362 = set1_unflattened[5'h06];
  assign sel_39363 = array_index_39280 == array_index_38946 ? add_39361 : sel_39357;
  assign add_39366 = sel_39363 + 8'h01;
  assign sel_39367 = array_index_39362 == array_index_38822 ? add_39366 : sel_39363;
  assign add_39370 = sel_39367 + 8'h01;
  assign sel_39371 = array_index_39362 == array_index_38826 ? add_39370 : sel_39367;
  assign add_39374 = sel_39371 + 8'h01;
  assign sel_39375 = array_index_39362 == array_index_38834 ? add_39374 : sel_39371;
  assign add_39378 = sel_39375 + 8'h01;
  assign sel_39379 = array_index_39362 == array_index_38842 ? add_39378 : sel_39375;
  assign add_39382 = sel_39379 + 8'h01;
  assign sel_39383 = array_index_39362 == array_index_38850 ? add_39382 : sel_39379;
  assign add_39386 = sel_39383 + 8'h01;
  assign sel_39387 = array_index_39362 == array_index_38858 ? add_39386 : sel_39383;
  assign add_39390 = sel_39387 + 8'h01;
  assign sel_39391 = array_index_39362 == array_index_38866 ? add_39390 : sel_39387;
  assign add_39394 = sel_39391 + 8'h01;
  assign sel_39395 = array_index_39362 == array_index_38874 ? add_39394 : sel_39391;
  assign add_39398 = sel_39395 + 8'h01;
  assign sel_39399 = array_index_39362 == array_index_38880 ? add_39398 : sel_39395;
  assign add_39402 = sel_39399 + 8'h01;
  assign sel_39403 = array_index_39362 == array_index_38886 ? add_39402 : sel_39399;
  assign add_39406 = sel_39403 + 8'h01;
  assign sel_39407 = array_index_39362 == array_index_38892 ? add_39406 : sel_39403;
  assign add_39410 = sel_39407 + 8'h01;
  assign sel_39411 = array_index_39362 == array_index_38898 ? add_39410 : sel_39407;
  assign add_39414 = sel_39411 + 8'h01;
  assign sel_39415 = array_index_39362 == array_index_38904 ? add_39414 : sel_39411;
  assign add_39418 = sel_39415 + 8'h01;
  assign sel_39419 = array_index_39362 == array_index_38910 ? add_39418 : sel_39415;
  assign add_39422 = sel_39419 + 8'h01;
  assign sel_39423 = array_index_39362 == array_index_38916 ? add_39422 : sel_39419;
  assign add_39426 = sel_39423 + 8'h01;
  assign sel_39427 = array_index_39362 == array_index_38922 ? add_39426 : sel_39423;
  assign add_39430 = sel_39427 + 8'h01;
  assign sel_39431 = array_index_39362 == array_index_38928 ? add_39430 : sel_39427;
  assign add_39434 = sel_39431 + 8'h01;
  assign sel_39435 = array_index_39362 == array_index_38934 ? add_39434 : sel_39431;
  assign add_39438 = sel_39435 + 8'h01;
  assign sel_39439 = array_index_39362 == array_index_38940 ? add_39438 : sel_39435;
  assign add_39443 = sel_39439 + 8'h01;
  assign array_index_39444 = set1_unflattened[5'h07];
  assign sel_39445 = array_index_39362 == array_index_38946 ? add_39443 : sel_39439;
  assign add_39448 = sel_39445 + 8'h01;
  assign sel_39449 = array_index_39444 == array_index_38822 ? add_39448 : sel_39445;
  assign add_39452 = sel_39449 + 8'h01;
  assign sel_39453 = array_index_39444 == array_index_38826 ? add_39452 : sel_39449;
  assign add_39456 = sel_39453 + 8'h01;
  assign sel_39457 = array_index_39444 == array_index_38834 ? add_39456 : sel_39453;
  assign add_39460 = sel_39457 + 8'h01;
  assign sel_39461 = array_index_39444 == array_index_38842 ? add_39460 : sel_39457;
  assign add_39464 = sel_39461 + 8'h01;
  assign sel_39465 = array_index_39444 == array_index_38850 ? add_39464 : sel_39461;
  assign add_39468 = sel_39465 + 8'h01;
  assign sel_39469 = array_index_39444 == array_index_38858 ? add_39468 : sel_39465;
  assign add_39472 = sel_39469 + 8'h01;
  assign sel_39473 = array_index_39444 == array_index_38866 ? add_39472 : sel_39469;
  assign add_39476 = sel_39473 + 8'h01;
  assign sel_39477 = array_index_39444 == array_index_38874 ? add_39476 : sel_39473;
  assign add_39480 = sel_39477 + 8'h01;
  assign sel_39481 = array_index_39444 == array_index_38880 ? add_39480 : sel_39477;
  assign add_39484 = sel_39481 + 8'h01;
  assign sel_39485 = array_index_39444 == array_index_38886 ? add_39484 : sel_39481;
  assign add_39488 = sel_39485 + 8'h01;
  assign sel_39489 = array_index_39444 == array_index_38892 ? add_39488 : sel_39485;
  assign add_39492 = sel_39489 + 8'h01;
  assign sel_39493 = array_index_39444 == array_index_38898 ? add_39492 : sel_39489;
  assign add_39496 = sel_39493 + 8'h01;
  assign sel_39497 = array_index_39444 == array_index_38904 ? add_39496 : sel_39493;
  assign add_39500 = sel_39497 + 8'h01;
  assign sel_39501 = array_index_39444 == array_index_38910 ? add_39500 : sel_39497;
  assign add_39504 = sel_39501 + 8'h01;
  assign sel_39505 = array_index_39444 == array_index_38916 ? add_39504 : sel_39501;
  assign add_39508 = sel_39505 + 8'h01;
  assign sel_39509 = array_index_39444 == array_index_38922 ? add_39508 : sel_39505;
  assign add_39512 = sel_39509 + 8'h01;
  assign sel_39513 = array_index_39444 == array_index_38928 ? add_39512 : sel_39509;
  assign add_39516 = sel_39513 + 8'h01;
  assign sel_39517 = array_index_39444 == array_index_38934 ? add_39516 : sel_39513;
  assign add_39520 = sel_39517 + 8'h01;
  assign sel_39521 = array_index_39444 == array_index_38940 ? add_39520 : sel_39517;
  assign add_39525 = sel_39521 + 8'h01;
  assign array_index_39526 = set1_unflattened[5'h08];
  assign sel_39527 = array_index_39444 == array_index_38946 ? add_39525 : sel_39521;
  assign add_39530 = sel_39527 + 8'h01;
  assign sel_39531 = array_index_39526 == array_index_38822 ? add_39530 : sel_39527;
  assign add_39534 = sel_39531 + 8'h01;
  assign sel_39535 = array_index_39526 == array_index_38826 ? add_39534 : sel_39531;
  assign add_39538 = sel_39535 + 8'h01;
  assign sel_39539 = array_index_39526 == array_index_38834 ? add_39538 : sel_39535;
  assign add_39542 = sel_39539 + 8'h01;
  assign sel_39543 = array_index_39526 == array_index_38842 ? add_39542 : sel_39539;
  assign add_39546 = sel_39543 + 8'h01;
  assign sel_39547 = array_index_39526 == array_index_38850 ? add_39546 : sel_39543;
  assign add_39550 = sel_39547 + 8'h01;
  assign sel_39551 = array_index_39526 == array_index_38858 ? add_39550 : sel_39547;
  assign add_39554 = sel_39551 + 8'h01;
  assign sel_39555 = array_index_39526 == array_index_38866 ? add_39554 : sel_39551;
  assign add_39558 = sel_39555 + 8'h01;
  assign sel_39559 = array_index_39526 == array_index_38874 ? add_39558 : sel_39555;
  assign add_39562 = sel_39559 + 8'h01;
  assign sel_39563 = array_index_39526 == array_index_38880 ? add_39562 : sel_39559;
  assign add_39566 = sel_39563 + 8'h01;
  assign sel_39567 = array_index_39526 == array_index_38886 ? add_39566 : sel_39563;
  assign add_39570 = sel_39567 + 8'h01;
  assign sel_39571 = array_index_39526 == array_index_38892 ? add_39570 : sel_39567;
  assign add_39574 = sel_39571 + 8'h01;
  assign sel_39575 = array_index_39526 == array_index_38898 ? add_39574 : sel_39571;
  assign add_39578 = sel_39575 + 8'h01;
  assign sel_39579 = array_index_39526 == array_index_38904 ? add_39578 : sel_39575;
  assign add_39582 = sel_39579 + 8'h01;
  assign sel_39583 = array_index_39526 == array_index_38910 ? add_39582 : sel_39579;
  assign add_39586 = sel_39583 + 8'h01;
  assign sel_39587 = array_index_39526 == array_index_38916 ? add_39586 : sel_39583;
  assign add_39590 = sel_39587 + 8'h01;
  assign sel_39591 = array_index_39526 == array_index_38922 ? add_39590 : sel_39587;
  assign add_39594 = sel_39591 + 8'h01;
  assign sel_39595 = array_index_39526 == array_index_38928 ? add_39594 : sel_39591;
  assign add_39598 = sel_39595 + 8'h01;
  assign sel_39599 = array_index_39526 == array_index_38934 ? add_39598 : sel_39595;
  assign add_39602 = sel_39599 + 8'h01;
  assign sel_39603 = array_index_39526 == array_index_38940 ? add_39602 : sel_39599;
  assign add_39607 = sel_39603 + 8'h01;
  assign array_index_39608 = set1_unflattened[5'h09];
  assign sel_39609 = array_index_39526 == array_index_38946 ? add_39607 : sel_39603;
  assign add_39612 = sel_39609 + 8'h01;
  assign sel_39613 = array_index_39608 == array_index_38822 ? add_39612 : sel_39609;
  assign add_39616 = sel_39613 + 8'h01;
  assign sel_39617 = array_index_39608 == array_index_38826 ? add_39616 : sel_39613;
  assign add_39620 = sel_39617 + 8'h01;
  assign sel_39621 = array_index_39608 == array_index_38834 ? add_39620 : sel_39617;
  assign add_39624 = sel_39621 + 8'h01;
  assign sel_39625 = array_index_39608 == array_index_38842 ? add_39624 : sel_39621;
  assign add_39628 = sel_39625 + 8'h01;
  assign sel_39629 = array_index_39608 == array_index_38850 ? add_39628 : sel_39625;
  assign add_39632 = sel_39629 + 8'h01;
  assign sel_39633 = array_index_39608 == array_index_38858 ? add_39632 : sel_39629;
  assign add_39636 = sel_39633 + 8'h01;
  assign sel_39637 = array_index_39608 == array_index_38866 ? add_39636 : sel_39633;
  assign add_39640 = sel_39637 + 8'h01;
  assign sel_39641 = array_index_39608 == array_index_38874 ? add_39640 : sel_39637;
  assign add_39644 = sel_39641 + 8'h01;
  assign sel_39645 = array_index_39608 == array_index_38880 ? add_39644 : sel_39641;
  assign add_39648 = sel_39645 + 8'h01;
  assign sel_39649 = array_index_39608 == array_index_38886 ? add_39648 : sel_39645;
  assign add_39652 = sel_39649 + 8'h01;
  assign sel_39653 = array_index_39608 == array_index_38892 ? add_39652 : sel_39649;
  assign add_39656 = sel_39653 + 8'h01;
  assign sel_39657 = array_index_39608 == array_index_38898 ? add_39656 : sel_39653;
  assign add_39660 = sel_39657 + 8'h01;
  assign sel_39661 = array_index_39608 == array_index_38904 ? add_39660 : sel_39657;
  assign add_39664 = sel_39661 + 8'h01;
  assign sel_39665 = array_index_39608 == array_index_38910 ? add_39664 : sel_39661;
  assign add_39668 = sel_39665 + 8'h01;
  assign sel_39669 = array_index_39608 == array_index_38916 ? add_39668 : sel_39665;
  assign add_39672 = sel_39669 + 8'h01;
  assign sel_39673 = array_index_39608 == array_index_38922 ? add_39672 : sel_39669;
  assign add_39676 = sel_39673 + 8'h01;
  assign sel_39677 = array_index_39608 == array_index_38928 ? add_39676 : sel_39673;
  assign add_39680 = sel_39677 + 8'h01;
  assign sel_39681 = array_index_39608 == array_index_38934 ? add_39680 : sel_39677;
  assign add_39684 = sel_39681 + 8'h01;
  assign sel_39685 = array_index_39608 == array_index_38940 ? add_39684 : sel_39681;
  assign add_39689 = sel_39685 + 8'h01;
  assign array_index_39690 = set1_unflattened[5'h0a];
  assign sel_39691 = array_index_39608 == array_index_38946 ? add_39689 : sel_39685;
  assign add_39694 = sel_39691 + 8'h01;
  assign sel_39695 = array_index_39690 == array_index_38822 ? add_39694 : sel_39691;
  assign add_39698 = sel_39695 + 8'h01;
  assign sel_39699 = array_index_39690 == array_index_38826 ? add_39698 : sel_39695;
  assign add_39702 = sel_39699 + 8'h01;
  assign sel_39703 = array_index_39690 == array_index_38834 ? add_39702 : sel_39699;
  assign add_39706 = sel_39703 + 8'h01;
  assign sel_39707 = array_index_39690 == array_index_38842 ? add_39706 : sel_39703;
  assign add_39710 = sel_39707 + 8'h01;
  assign sel_39711 = array_index_39690 == array_index_38850 ? add_39710 : sel_39707;
  assign add_39714 = sel_39711 + 8'h01;
  assign sel_39715 = array_index_39690 == array_index_38858 ? add_39714 : sel_39711;
  assign add_39718 = sel_39715 + 8'h01;
  assign sel_39719 = array_index_39690 == array_index_38866 ? add_39718 : sel_39715;
  assign add_39722 = sel_39719 + 8'h01;
  assign sel_39723 = array_index_39690 == array_index_38874 ? add_39722 : sel_39719;
  assign add_39726 = sel_39723 + 8'h01;
  assign sel_39727 = array_index_39690 == array_index_38880 ? add_39726 : sel_39723;
  assign add_39730 = sel_39727 + 8'h01;
  assign sel_39731 = array_index_39690 == array_index_38886 ? add_39730 : sel_39727;
  assign add_39734 = sel_39731 + 8'h01;
  assign sel_39735 = array_index_39690 == array_index_38892 ? add_39734 : sel_39731;
  assign add_39738 = sel_39735 + 8'h01;
  assign sel_39739 = array_index_39690 == array_index_38898 ? add_39738 : sel_39735;
  assign add_39742 = sel_39739 + 8'h01;
  assign sel_39743 = array_index_39690 == array_index_38904 ? add_39742 : sel_39739;
  assign add_39746 = sel_39743 + 8'h01;
  assign sel_39747 = array_index_39690 == array_index_38910 ? add_39746 : sel_39743;
  assign add_39750 = sel_39747 + 8'h01;
  assign sel_39751 = array_index_39690 == array_index_38916 ? add_39750 : sel_39747;
  assign add_39754 = sel_39751 + 8'h01;
  assign sel_39755 = array_index_39690 == array_index_38922 ? add_39754 : sel_39751;
  assign add_39758 = sel_39755 + 8'h01;
  assign sel_39759 = array_index_39690 == array_index_38928 ? add_39758 : sel_39755;
  assign add_39762 = sel_39759 + 8'h01;
  assign sel_39763 = array_index_39690 == array_index_38934 ? add_39762 : sel_39759;
  assign add_39766 = sel_39763 + 8'h01;
  assign sel_39767 = array_index_39690 == array_index_38940 ? add_39766 : sel_39763;
  assign add_39771 = sel_39767 + 8'h01;
  assign array_index_39772 = set1_unflattened[5'h0b];
  assign sel_39773 = array_index_39690 == array_index_38946 ? add_39771 : sel_39767;
  assign add_39776 = sel_39773 + 8'h01;
  assign sel_39777 = array_index_39772 == array_index_38822 ? add_39776 : sel_39773;
  assign add_39780 = sel_39777 + 8'h01;
  assign sel_39781 = array_index_39772 == array_index_38826 ? add_39780 : sel_39777;
  assign add_39784 = sel_39781 + 8'h01;
  assign sel_39785 = array_index_39772 == array_index_38834 ? add_39784 : sel_39781;
  assign add_39788 = sel_39785 + 8'h01;
  assign sel_39789 = array_index_39772 == array_index_38842 ? add_39788 : sel_39785;
  assign add_39792 = sel_39789 + 8'h01;
  assign sel_39793 = array_index_39772 == array_index_38850 ? add_39792 : sel_39789;
  assign add_39796 = sel_39793 + 8'h01;
  assign sel_39797 = array_index_39772 == array_index_38858 ? add_39796 : sel_39793;
  assign add_39800 = sel_39797 + 8'h01;
  assign sel_39801 = array_index_39772 == array_index_38866 ? add_39800 : sel_39797;
  assign add_39804 = sel_39801 + 8'h01;
  assign sel_39805 = array_index_39772 == array_index_38874 ? add_39804 : sel_39801;
  assign add_39808 = sel_39805 + 8'h01;
  assign sel_39809 = array_index_39772 == array_index_38880 ? add_39808 : sel_39805;
  assign add_39812 = sel_39809 + 8'h01;
  assign sel_39813 = array_index_39772 == array_index_38886 ? add_39812 : sel_39809;
  assign add_39816 = sel_39813 + 8'h01;
  assign sel_39817 = array_index_39772 == array_index_38892 ? add_39816 : sel_39813;
  assign add_39820 = sel_39817 + 8'h01;
  assign sel_39821 = array_index_39772 == array_index_38898 ? add_39820 : sel_39817;
  assign add_39824 = sel_39821 + 8'h01;
  assign sel_39825 = array_index_39772 == array_index_38904 ? add_39824 : sel_39821;
  assign add_39828 = sel_39825 + 8'h01;
  assign sel_39829 = array_index_39772 == array_index_38910 ? add_39828 : sel_39825;
  assign add_39832 = sel_39829 + 8'h01;
  assign sel_39833 = array_index_39772 == array_index_38916 ? add_39832 : sel_39829;
  assign add_39836 = sel_39833 + 8'h01;
  assign sel_39837 = array_index_39772 == array_index_38922 ? add_39836 : sel_39833;
  assign add_39840 = sel_39837 + 8'h01;
  assign sel_39841 = array_index_39772 == array_index_38928 ? add_39840 : sel_39837;
  assign add_39844 = sel_39841 + 8'h01;
  assign sel_39845 = array_index_39772 == array_index_38934 ? add_39844 : sel_39841;
  assign add_39848 = sel_39845 + 8'h01;
  assign sel_39849 = array_index_39772 == array_index_38940 ? add_39848 : sel_39845;
  assign add_39853 = sel_39849 + 8'h01;
  assign array_index_39854 = set1_unflattened[5'h0c];
  assign sel_39855 = array_index_39772 == array_index_38946 ? add_39853 : sel_39849;
  assign add_39858 = sel_39855 + 8'h01;
  assign sel_39859 = array_index_39854 == array_index_38822 ? add_39858 : sel_39855;
  assign add_39862 = sel_39859 + 8'h01;
  assign sel_39863 = array_index_39854 == array_index_38826 ? add_39862 : sel_39859;
  assign add_39866 = sel_39863 + 8'h01;
  assign sel_39867 = array_index_39854 == array_index_38834 ? add_39866 : sel_39863;
  assign add_39870 = sel_39867 + 8'h01;
  assign sel_39871 = array_index_39854 == array_index_38842 ? add_39870 : sel_39867;
  assign add_39874 = sel_39871 + 8'h01;
  assign sel_39875 = array_index_39854 == array_index_38850 ? add_39874 : sel_39871;
  assign add_39878 = sel_39875 + 8'h01;
  assign sel_39879 = array_index_39854 == array_index_38858 ? add_39878 : sel_39875;
  assign add_39882 = sel_39879 + 8'h01;
  assign sel_39883 = array_index_39854 == array_index_38866 ? add_39882 : sel_39879;
  assign add_39886 = sel_39883 + 8'h01;
  assign sel_39887 = array_index_39854 == array_index_38874 ? add_39886 : sel_39883;
  assign add_39890 = sel_39887 + 8'h01;
  assign sel_39891 = array_index_39854 == array_index_38880 ? add_39890 : sel_39887;
  assign add_39894 = sel_39891 + 8'h01;
  assign sel_39895 = array_index_39854 == array_index_38886 ? add_39894 : sel_39891;
  assign add_39898 = sel_39895 + 8'h01;
  assign sel_39899 = array_index_39854 == array_index_38892 ? add_39898 : sel_39895;
  assign add_39902 = sel_39899 + 8'h01;
  assign sel_39903 = array_index_39854 == array_index_38898 ? add_39902 : sel_39899;
  assign add_39906 = sel_39903 + 8'h01;
  assign sel_39907 = array_index_39854 == array_index_38904 ? add_39906 : sel_39903;
  assign add_39910 = sel_39907 + 8'h01;
  assign sel_39911 = array_index_39854 == array_index_38910 ? add_39910 : sel_39907;
  assign add_39914 = sel_39911 + 8'h01;
  assign sel_39915 = array_index_39854 == array_index_38916 ? add_39914 : sel_39911;
  assign add_39918 = sel_39915 + 8'h01;
  assign sel_39919 = array_index_39854 == array_index_38922 ? add_39918 : sel_39915;
  assign add_39922 = sel_39919 + 8'h01;
  assign sel_39923 = array_index_39854 == array_index_38928 ? add_39922 : sel_39919;
  assign add_39926 = sel_39923 + 8'h01;
  assign sel_39927 = array_index_39854 == array_index_38934 ? add_39926 : sel_39923;
  assign add_39930 = sel_39927 + 8'h01;
  assign sel_39931 = array_index_39854 == array_index_38940 ? add_39930 : sel_39927;
  assign add_39935 = sel_39931 + 8'h01;
  assign array_index_39936 = set1_unflattened[5'h0d];
  assign sel_39937 = array_index_39854 == array_index_38946 ? add_39935 : sel_39931;
  assign add_39940 = sel_39937 + 8'h01;
  assign sel_39941 = array_index_39936 == array_index_38822 ? add_39940 : sel_39937;
  assign add_39944 = sel_39941 + 8'h01;
  assign sel_39945 = array_index_39936 == array_index_38826 ? add_39944 : sel_39941;
  assign add_39948 = sel_39945 + 8'h01;
  assign sel_39949 = array_index_39936 == array_index_38834 ? add_39948 : sel_39945;
  assign add_39952 = sel_39949 + 8'h01;
  assign sel_39953 = array_index_39936 == array_index_38842 ? add_39952 : sel_39949;
  assign add_39956 = sel_39953 + 8'h01;
  assign sel_39957 = array_index_39936 == array_index_38850 ? add_39956 : sel_39953;
  assign add_39960 = sel_39957 + 8'h01;
  assign sel_39961 = array_index_39936 == array_index_38858 ? add_39960 : sel_39957;
  assign add_39964 = sel_39961 + 8'h01;
  assign sel_39965 = array_index_39936 == array_index_38866 ? add_39964 : sel_39961;
  assign add_39968 = sel_39965 + 8'h01;
  assign sel_39969 = array_index_39936 == array_index_38874 ? add_39968 : sel_39965;
  assign add_39972 = sel_39969 + 8'h01;
  assign sel_39973 = array_index_39936 == array_index_38880 ? add_39972 : sel_39969;
  assign add_39976 = sel_39973 + 8'h01;
  assign sel_39977 = array_index_39936 == array_index_38886 ? add_39976 : sel_39973;
  assign add_39980 = sel_39977 + 8'h01;
  assign sel_39981 = array_index_39936 == array_index_38892 ? add_39980 : sel_39977;
  assign add_39984 = sel_39981 + 8'h01;
  assign sel_39985 = array_index_39936 == array_index_38898 ? add_39984 : sel_39981;
  assign add_39988 = sel_39985 + 8'h01;
  assign sel_39989 = array_index_39936 == array_index_38904 ? add_39988 : sel_39985;
  assign add_39992 = sel_39989 + 8'h01;
  assign sel_39993 = array_index_39936 == array_index_38910 ? add_39992 : sel_39989;
  assign add_39996 = sel_39993 + 8'h01;
  assign sel_39997 = array_index_39936 == array_index_38916 ? add_39996 : sel_39993;
  assign add_40000 = sel_39997 + 8'h01;
  assign sel_40001 = array_index_39936 == array_index_38922 ? add_40000 : sel_39997;
  assign add_40004 = sel_40001 + 8'h01;
  assign sel_40005 = array_index_39936 == array_index_38928 ? add_40004 : sel_40001;
  assign add_40008 = sel_40005 + 8'h01;
  assign sel_40009 = array_index_39936 == array_index_38934 ? add_40008 : sel_40005;
  assign add_40012 = sel_40009 + 8'h01;
  assign sel_40013 = array_index_39936 == array_index_38940 ? add_40012 : sel_40009;
  assign add_40017 = sel_40013 + 8'h01;
  assign array_index_40018 = set1_unflattened[5'h0e];
  assign sel_40019 = array_index_39936 == array_index_38946 ? add_40017 : sel_40013;
  assign add_40022 = sel_40019 + 8'h01;
  assign sel_40023 = array_index_40018 == array_index_38822 ? add_40022 : sel_40019;
  assign add_40026 = sel_40023 + 8'h01;
  assign sel_40027 = array_index_40018 == array_index_38826 ? add_40026 : sel_40023;
  assign add_40030 = sel_40027 + 8'h01;
  assign sel_40031 = array_index_40018 == array_index_38834 ? add_40030 : sel_40027;
  assign add_40034 = sel_40031 + 8'h01;
  assign sel_40035 = array_index_40018 == array_index_38842 ? add_40034 : sel_40031;
  assign add_40038 = sel_40035 + 8'h01;
  assign sel_40039 = array_index_40018 == array_index_38850 ? add_40038 : sel_40035;
  assign add_40042 = sel_40039 + 8'h01;
  assign sel_40043 = array_index_40018 == array_index_38858 ? add_40042 : sel_40039;
  assign add_40046 = sel_40043 + 8'h01;
  assign sel_40047 = array_index_40018 == array_index_38866 ? add_40046 : sel_40043;
  assign add_40050 = sel_40047 + 8'h01;
  assign sel_40051 = array_index_40018 == array_index_38874 ? add_40050 : sel_40047;
  assign add_40054 = sel_40051 + 8'h01;
  assign sel_40055 = array_index_40018 == array_index_38880 ? add_40054 : sel_40051;
  assign add_40058 = sel_40055 + 8'h01;
  assign sel_40059 = array_index_40018 == array_index_38886 ? add_40058 : sel_40055;
  assign add_40062 = sel_40059 + 8'h01;
  assign sel_40063 = array_index_40018 == array_index_38892 ? add_40062 : sel_40059;
  assign add_40066 = sel_40063 + 8'h01;
  assign sel_40067 = array_index_40018 == array_index_38898 ? add_40066 : sel_40063;
  assign add_40070 = sel_40067 + 8'h01;
  assign sel_40071 = array_index_40018 == array_index_38904 ? add_40070 : sel_40067;
  assign add_40074 = sel_40071 + 8'h01;
  assign sel_40075 = array_index_40018 == array_index_38910 ? add_40074 : sel_40071;
  assign add_40078 = sel_40075 + 8'h01;
  assign sel_40079 = array_index_40018 == array_index_38916 ? add_40078 : sel_40075;
  assign add_40082 = sel_40079 + 8'h01;
  assign sel_40083 = array_index_40018 == array_index_38922 ? add_40082 : sel_40079;
  assign add_40086 = sel_40083 + 8'h01;
  assign sel_40087 = array_index_40018 == array_index_38928 ? add_40086 : sel_40083;
  assign add_40090 = sel_40087 + 8'h01;
  assign sel_40091 = array_index_40018 == array_index_38934 ? add_40090 : sel_40087;
  assign add_40094 = sel_40091 + 8'h01;
  assign sel_40095 = array_index_40018 == array_index_38940 ? add_40094 : sel_40091;
  assign add_40099 = sel_40095 + 8'h01;
  assign array_index_40100 = set1_unflattened[5'h0f];
  assign sel_40101 = array_index_40018 == array_index_38946 ? add_40099 : sel_40095;
  assign add_40104 = sel_40101 + 8'h01;
  assign sel_40105 = array_index_40100 == array_index_38822 ? add_40104 : sel_40101;
  assign add_40108 = sel_40105 + 8'h01;
  assign sel_40109 = array_index_40100 == array_index_38826 ? add_40108 : sel_40105;
  assign add_40112 = sel_40109 + 8'h01;
  assign sel_40113 = array_index_40100 == array_index_38834 ? add_40112 : sel_40109;
  assign add_40116 = sel_40113 + 8'h01;
  assign sel_40117 = array_index_40100 == array_index_38842 ? add_40116 : sel_40113;
  assign add_40120 = sel_40117 + 8'h01;
  assign sel_40121 = array_index_40100 == array_index_38850 ? add_40120 : sel_40117;
  assign add_40124 = sel_40121 + 8'h01;
  assign sel_40125 = array_index_40100 == array_index_38858 ? add_40124 : sel_40121;
  assign add_40128 = sel_40125 + 8'h01;
  assign sel_40129 = array_index_40100 == array_index_38866 ? add_40128 : sel_40125;
  assign add_40132 = sel_40129 + 8'h01;
  assign sel_40133 = array_index_40100 == array_index_38874 ? add_40132 : sel_40129;
  assign add_40136 = sel_40133 + 8'h01;
  assign sel_40137 = array_index_40100 == array_index_38880 ? add_40136 : sel_40133;
  assign add_40140 = sel_40137 + 8'h01;
  assign sel_40141 = array_index_40100 == array_index_38886 ? add_40140 : sel_40137;
  assign add_40144 = sel_40141 + 8'h01;
  assign sel_40145 = array_index_40100 == array_index_38892 ? add_40144 : sel_40141;
  assign add_40148 = sel_40145 + 8'h01;
  assign sel_40149 = array_index_40100 == array_index_38898 ? add_40148 : sel_40145;
  assign add_40152 = sel_40149 + 8'h01;
  assign sel_40153 = array_index_40100 == array_index_38904 ? add_40152 : sel_40149;
  assign add_40156 = sel_40153 + 8'h01;
  assign sel_40157 = array_index_40100 == array_index_38910 ? add_40156 : sel_40153;
  assign add_40160 = sel_40157 + 8'h01;
  assign sel_40161 = array_index_40100 == array_index_38916 ? add_40160 : sel_40157;
  assign add_40164 = sel_40161 + 8'h01;
  assign sel_40165 = array_index_40100 == array_index_38922 ? add_40164 : sel_40161;
  assign add_40168 = sel_40165 + 8'h01;
  assign sel_40169 = array_index_40100 == array_index_38928 ? add_40168 : sel_40165;
  assign add_40172 = sel_40169 + 8'h01;
  assign sel_40173 = array_index_40100 == array_index_38934 ? add_40172 : sel_40169;
  assign add_40176 = sel_40173 + 8'h01;
  assign sel_40177 = array_index_40100 == array_index_38940 ? add_40176 : sel_40173;
  assign add_40181 = sel_40177 + 8'h01;
  assign array_index_40182 = set1_unflattened[5'h10];
  assign sel_40183 = array_index_40100 == array_index_38946 ? add_40181 : sel_40177;
  assign add_40186 = sel_40183 + 8'h01;
  assign sel_40187 = array_index_40182 == array_index_38822 ? add_40186 : sel_40183;
  assign add_40190 = sel_40187 + 8'h01;
  assign sel_40191 = array_index_40182 == array_index_38826 ? add_40190 : sel_40187;
  assign add_40194 = sel_40191 + 8'h01;
  assign sel_40195 = array_index_40182 == array_index_38834 ? add_40194 : sel_40191;
  assign add_40198 = sel_40195 + 8'h01;
  assign sel_40199 = array_index_40182 == array_index_38842 ? add_40198 : sel_40195;
  assign add_40202 = sel_40199 + 8'h01;
  assign sel_40203 = array_index_40182 == array_index_38850 ? add_40202 : sel_40199;
  assign add_40206 = sel_40203 + 8'h01;
  assign sel_40207 = array_index_40182 == array_index_38858 ? add_40206 : sel_40203;
  assign add_40210 = sel_40207 + 8'h01;
  assign sel_40211 = array_index_40182 == array_index_38866 ? add_40210 : sel_40207;
  assign add_40214 = sel_40211 + 8'h01;
  assign sel_40215 = array_index_40182 == array_index_38874 ? add_40214 : sel_40211;
  assign add_40218 = sel_40215 + 8'h01;
  assign sel_40219 = array_index_40182 == array_index_38880 ? add_40218 : sel_40215;
  assign add_40222 = sel_40219 + 8'h01;
  assign sel_40223 = array_index_40182 == array_index_38886 ? add_40222 : sel_40219;
  assign add_40226 = sel_40223 + 8'h01;
  assign sel_40227 = array_index_40182 == array_index_38892 ? add_40226 : sel_40223;
  assign add_40230 = sel_40227 + 8'h01;
  assign sel_40231 = array_index_40182 == array_index_38898 ? add_40230 : sel_40227;
  assign add_40234 = sel_40231 + 8'h01;
  assign sel_40235 = array_index_40182 == array_index_38904 ? add_40234 : sel_40231;
  assign add_40238 = sel_40235 + 8'h01;
  assign sel_40239 = array_index_40182 == array_index_38910 ? add_40238 : sel_40235;
  assign add_40242 = sel_40239 + 8'h01;
  assign sel_40243 = array_index_40182 == array_index_38916 ? add_40242 : sel_40239;
  assign add_40246 = sel_40243 + 8'h01;
  assign sel_40247 = array_index_40182 == array_index_38922 ? add_40246 : sel_40243;
  assign add_40250 = sel_40247 + 8'h01;
  assign sel_40251 = array_index_40182 == array_index_38928 ? add_40250 : sel_40247;
  assign add_40254 = sel_40251 + 8'h01;
  assign sel_40255 = array_index_40182 == array_index_38934 ? add_40254 : sel_40251;
  assign add_40258 = sel_40255 + 8'h01;
  assign sel_40259 = array_index_40182 == array_index_38940 ? add_40258 : sel_40255;
  assign add_40263 = sel_40259 + 8'h01;
  assign array_index_40264 = set1_unflattened[5'h11];
  assign sel_40265 = array_index_40182 == array_index_38946 ? add_40263 : sel_40259;
  assign add_40268 = sel_40265 + 8'h01;
  assign sel_40269 = array_index_40264 == array_index_38822 ? add_40268 : sel_40265;
  assign add_40272 = sel_40269 + 8'h01;
  assign sel_40273 = array_index_40264 == array_index_38826 ? add_40272 : sel_40269;
  assign add_40276 = sel_40273 + 8'h01;
  assign sel_40277 = array_index_40264 == array_index_38834 ? add_40276 : sel_40273;
  assign add_40280 = sel_40277 + 8'h01;
  assign sel_40281 = array_index_40264 == array_index_38842 ? add_40280 : sel_40277;
  assign add_40284 = sel_40281 + 8'h01;
  assign sel_40285 = array_index_40264 == array_index_38850 ? add_40284 : sel_40281;
  assign add_40288 = sel_40285 + 8'h01;
  assign sel_40289 = array_index_40264 == array_index_38858 ? add_40288 : sel_40285;
  assign add_40292 = sel_40289 + 8'h01;
  assign sel_40293 = array_index_40264 == array_index_38866 ? add_40292 : sel_40289;
  assign add_40296 = sel_40293 + 8'h01;
  assign sel_40297 = array_index_40264 == array_index_38874 ? add_40296 : sel_40293;
  assign add_40300 = sel_40297 + 8'h01;
  assign sel_40301 = array_index_40264 == array_index_38880 ? add_40300 : sel_40297;
  assign add_40304 = sel_40301 + 8'h01;
  assign sel_40305 = array_index_40264 == array_index_38886 ? add_40304 : sel_40301;
  assign add_40308 = sel_40305 + 8'h01;
  assign sel_40309 = array_index_40264 == array_index_38892 ? add_40308 : sel_40305;
  assign add_40312 = sel_40309 + 8'h01;
  assign sel_40313 = array_index_40264 == array_index_38898 ? add_40312 : sel_40309;
  assign add_40316 = sel_40313 + 8'h01;
  assign sel_40317 = array_index_40264 == array_index_38904 ? add_40316 : sel_40313;
  assign add_40320 = sel_40317 + 8'h01;
  assign sel_40321 = array_index_40264 == array_index_38910 ? add_40320 : sel_40317;
  assign add_40324 = sel_40321 + 8'h01;
  assign sel_40325 = array_index_40264 == array_index_38916 ? add_40324 : sel_40321;
  assign add_40328 = sel_40325 + 8'h01;
  assign sel_40329 = array_index_40264 == array_index_38922 ? add_40328 : sel_40325;
  assign add_40332 = sel_40329 + 8'h01;
  assign sel_40333 = array_index_40264 == array_index_38928 ? add_40332 : sel_40329;
  assign add_40336 = sel_40333 + 8'h01;
  assign sel_40337 = array_index_40264 == array_index_38934 ? add_40336 : sel_40333;
  assign add_40340 = sel_40337 + 8'h01;
  assign sel_40341 = array_index_40264 == array_index_38940 ? add_40340 : sel_40337;
  assign add_40345 = sel_40341 + 8'h01;
  assign array_index_40346 = set1_unflattened[5'h12];
  assign sel_40347 = array_index_40264 == array_index_38946 ? add_40345 : sel_40341;
  assign add_40350 = sel_40347 + 8'h01;
  assign sel_40351 = array_index_40346 == array_index_38822 ? add_40350 : sel_40347;
  assign add_40354 = sel_40351 + 8'h01;
  assign sel_40355 = array_index_40346 == array_index_38826 ? add_40354 : sel_40351;
  assign add_40358 = sel_40355 + 8'h01;
  assign sel_40359 = array_index_40346 == array_index_38834 ? add_40358 : sel_40355;
  assign add_40362 = sel_40359 + 8'h01;
  assign sel_40363 = array_index_40346 == array_index_38842 ? add_40362 : sel_40359;
  assign add_40366 = sel_40363 + 8'h01;
  assign sel_40367 = array_index_40346 == array_index_38850 ? add_40366 : sel_40363;
  assign add_40370 = sel_40367 + 8'h01;
  assign sel_40371 = array_index_40346 == array_index_38858 ? add_40370 : sel_40367;
  assign add_40374 = sel_40371 + 8'h01;
  assign sel_40375 = array_index_40346 == array_index_38866 ? add_40374 : sel_40371;
  assign add_40378 = sel_40375 + 8'h01;
  assign sel_40379 = array_index_40346 == array_index_38874 ? add_40378 : sel_40375;
  assign add_40382 = sel_40379 + 8'h01;
  assign sel_40383 = array_index_40346 == array_index_38880 ? add_40382 : sel_40379;
  assign add_40386 = sel_40383 + 8'h01;
  assign sel_40387 = array_index_40346 == array_index_38886 ? add_40386 : sel_40383;
  assign add_40390 = sel_40387 + 8'h01;
  assign sel_40391 = array_index_40346 == array_index_38892 ? add_40390 : sel_40387;
  assign add_40394 = sel_40391 + 8'h01;
  assign sel_40395 = array_index_40346 == array_index_38898 ? add_40394 : sel_40391;
  assign add_40398 = sel_40395 + 8'h01;
  assign sel_40399 = array_index_40346 == array_index_38904 ? add_40398 : sel_40395;
  assign add_40402 = sel_40399 + 8'h01;
  assign sel_40403 = array_index_40346 == array_index_38910 ? add_40402 : sel_40399;
  assign add_40406 = sel_40403 + 8'h01;
  assign sel_40407 = array_index_40346 == array_index_38916 ? add_40406 : sel_40403;
  assign add_40410 = sel_40407 + 8'h01;
  assign sel_40411 = array_index_40346 == array_index_38922 ? add_40410 : sel_40407;
  assign add_40414 = sel_40411 + 8'h01;
  assign sel_40415 = array_index_40346 == array_index_38928 ? add_40414 : sel_40411;
  assign add_40418 = sel_40415 + 8'h01;
  assign sel_40419 = array_index_40346 == array_index_38934 ? add_40418 : sel_40415;
  assign add_40422 = sel_40419 + 8'h01;
  assign sel_40423 = array_index_40346 == array_index_38940 ? add_40422 : sel_40419;
  assign add_40427 = sel_40423 + 8'h01;
  assign array_index_40428 = set1_unflattened[5'h13];
  assign sel_40429 = array_index_40346 == array_index_38946 ? add_40427 : sel_40423;
  assign add_40432 = sel_40429 + 8'h01;
  assign sel_40433 = array_index_40428 == array_index_38822 ? add_40432 : sel_40429;
  assign add_40436 = sel_40433 + 8'h01;
  assign sel_40437 = array_index_40428 == array_index_38826 ? add_40436 : sel_40433;
  assign add_40440 = sel_40437 + 8'h01;
  assign sel_40441 = array_index_40428 == array_index_38834 ? add_40440 : sel_40437;
  assign add_40444 = sel_40441 + 8'h01;
  assign sel_40445 = array_index_40428 == array_index_38842 ? add_40444 : sel_40441;
  assign add_40448 = sel_40445 + 8'h01;
  assign sel_40449 = array_index_40428 == array_index_38850 ? add_40448 : sel_40445;
  assign add_40452 = sel_40449 + 8'h01;
  assign sel_40453 = array_index_40428 == array_index_38858 ? add_40452 : sel_40449;
  assign add_40456 = sel_40453 + 8'h01;
  assign sel_40457 = array_index_40428 == array_index_38866 ? add_40456 : sel_40453;
  assign add_40460 = sel_40457 + 8'h01;
  assign sel_40461 = array_index_40428 == array_index_38874 ? add_40460 : sel_40457;
  assign add_40464 = sel_40461 + 8'h01;
  assign sel_40465 = array_index_40428 == array_index_38880 ? add_40464 : sel_40461;
  assign add_40468 = sel_40465 + 8'h01;
  assign sel_40469 = array_index_40428 == array_index_38886 ? add_40468 : sel_40465;
  assign add_40472 = sel_40469 + 8'h01;
  assign sel_40473 = array_index_40428 == array_index_38892 ? add_40472 : sel_40469;
  assign add_40476 = sel_40473 + 8'h01;
  assign sel_40477 = array_index_40428 == array_index_38898 ? add_40476 : sel_40473;
  assign add_40480 = sel_40477 + 8'h01;
  assign sel_40481 = array_index_40428 == array_index_38904 ? add_40480 : sel_40477;
  assign add_40484 = sel_40481 + 8'h01;
  assign sel_40485 = array_index_40428 == array_index_38910 ? add_40484 : sel_40481;
  assign add_40488 = sel_40485 + 8'h01;
  assign sel_40489 = array_index_40428 == array_index_38916 ? add_40488 : sel_40485;
  assign add_40492 = sel_40489 + 8'h01;
  assign sel_40493 = array_index_40428 == array_index_38922 ? add_40492 : sel_40489;
  assign add_40496 = sel_40493 + 8'h01;
  assign sel_40497 = array_index_40428 == array_index_38928 ? add_40496 : sel_40493;
  assign add_40500 = sel_40497 + 8'h01;
  assign sel_40501 = array_index_40428 == array_index_38934 ? add_40500 : sel_40497;
  assign add_40504 = sel_40501 + 8'h01;
  assign sel_40505 = array_index_40428 == array_index_38940 ? add_40504 : sel_40501;
  assign add_40508 = sel_40505 + 8'h01;
  assign out = {array_index_40428 == array_index_38946 ? add_40508 : sel_40505, {set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
