module min_hash(set1, set2, out);
  wire _000000_, _000001_, _000002_, _000003_, _000004_, _000005_, _000006_, _000007_, _000008_, _000009_, _000010_, _000011_, _000012_, _000013_, _000014_, _000015_, _000016_, _000017_, _000018_, _000019_, _000020_, _000021_, _000022_, _000023_, _000024_, _000025_, _000026_, _000027_, _000028_, _000029_, _000030_, _000031_, _000032_, _000033_, _000034_, _000035_, _000036_, _000037_, _000038_, _000039_, _000040_, _000041_, _000042_, _000043_, _000044_, _000045_, _000046_, _000047_, _000048_, _000049_, _000050_, _000051_, _000052_, _000053_, _000054_, _000055_, _000056_, _000057_, _000058_, _000059_, _000060_, _000061_, _000062_, _000063_, _000064_, _000065_, _000066_, _000067_, _000068_, _000069_, _000070_, _000071_, _000072_, _000073_, _000074_, _000075_, _000076_, _000077_, _000078_, _000079_, _000080_, _000081_, _000082_, _000083_, _000084_, _000085_, _000086_, _000087_, _000088_, _000089_, _000090_, _000091_, _000092_, _000093_, _000094_, _000095_, _000096_, _000097_, _000098_, _000099_, _000100_, _000101_, _000102_, _000103_, _000104_, _000105_, _000106_, _000107_, _000108_, _000109_, _000110_, _000111_, _000112_, _000113_, _000114_, _000115_, _000116_, _000117_, _000118_, _000119_, _000120_, _000121_, _000122_, _000123_, _000124_, _000125_, _000126_, _000127_, _000128_, _000129_, _000130_, _000131_, _000132_, _000133_, _000134_, _000135_, _000136_, _000137_, _000138_, _000139_, _000140_, _000141_, _000142_, _000143_, _000144_, _000145_, _000146_, _000147_, _000148_, _000149_, _000150_, _000151_, _000152_, _000153_, _000154_, _000155_, _000156_, _000157_, _000158_, _000159_, _000160_, _000161_, _000162_, _000163_, _000164_, _000165_, _000166_, _000167_, _000168_, _000169_, _000170_, _000171_, _000172_, _000173_, _000174_, _000175_, _000176_, _000177_, _000178_, _000179_, _000180_, _000181_, _000182_, _000183_, _000184_, _000185_, _000186_, _000187_, _000188_, _000189_, _000190_, _000191_, _000192_, _000193_, _000194_, _000195_, _000196_, _000197_, _000198_, _000199_, _000200_, _000201_, _000202_, _000203_, _000204_, _000205_, _000206_, _000207_, _000208_, _000209_, _000210_, _000211_, _000212_, _000213_, _000214_, _000215_, _000216_, _000217_, _000218_, _000219_, _000220_, _000221_, _000222_, _000223_, _000224_, _000225_, _000226_, _000227_, _000228_, _000229_, _000230_, _000231_, _000232_, _000233_, _000234_, _000235_, _000236_, _000237_, _000238_, _000239_, _000240_, _000241_, _000242_, _000243_, _000244_, _000245_, _000246_, _000247_, _000248_, _000249_, _000250_, _000251_, _000252_, _000253_, _000254_, _000255_, _000256_, _000257_, _000258_, _000259_, _000260_, _000261_, _000262_, _000263_, _000264_, _000265_, _000266_, _000267_, _000268_, _000269_, _000270_, _000271_, _000272_, _000273_, _000274_, _000275_, _000276_, _000277_, _000278_, _000279_, _000280_, _000281_, _000282_, _000283_, _000284_, _000285_, _000286_, _000287_, _000288_, _000289_, _000290_, _000291_, _000292_, _000293_, _000294_, _000295_, _000296_, _000297_, _000298_, _000299_, _000300_, _000301_, _000302_, _000303_, _000304_, _000305_, _000306_, _000307_, _000308_, _000309_, _000310_, _000311_, _000312_, _000313_, _000314_, _000315_, _000316_, _000317_, _000318_, _000319_, _000320_, _000321_, _000322_, _000323_, _000324_, _000325_, _000326_, _000327_, _000328_, _000329_, _000330_, _000331_, _000332_, _000333_, _000334_, _000335_, _000336_, _000337_, _000338_, _000339_, _000340_, _000341_, _000342_, _000343_, _000344_, _000345_, _000346_, _000347_, _000348_, _000349_, _000350_, _000351_, _000352_, _000353_, _000354_, _000355_, _000356_, _000357_, _000358_, _000359_, _000360_, _000361_, _000362_, _000363_, _000364_, _000365_, _000366_, _000367_, _000368_, _000369_, _000370_, _000371_, _000372_, _000373_, _000374_, _000375_, _000376_, _000377_, _000378_, _000379_, _000380_, _000381_, _000382_, _000383_, _000384_, _000385_, _000386_, _000387_, _000388_, _000389_, _000390_, _000391_, _000392_, _000393_, _000394_, _000395_, _000396_, _000397_, _000398_, _000399_, _000400_, _000401_, _000402_, _000403_, _000404_, _000405_, _000406_, _000407_, _000408_, _000409_, _000410_, _000411_, _000412_, _000413_, _000414_, _000415_, _000416_, _000417_, _000418_, _000419_, _000420_, _000421_, _000422_, _000423_, _000424_, _000425_, _000426_, _000427_, _000428_, _000429_, _000430_, _000431_, _000432_, _000433_, _000434_, _000435_, _000436_, _000437_, _000438_, _000439_, _000440_, _000441_, _000442_, _000443_, _000444_, _000445_, _000446_, _000447_, _000448_, _000449_, _000450_, _000451_, _000452_, _000453_, _000454_, _000455_, _000456_, _000457_, _000458_, _000459_, _000460_, _000461_, _000462_, _000463_, _000464_, _000465_, _000466_, _000467_, _000468_, _000469_, _000470_, _000471_, _000472_, _000473_, _000474_, _000475_, _000476_, _000477_, _000478_, _000479_, _000480_, _000481_, _000482_, _000483_, _000484_, _000485_, _000486_, _000487_, _000488_, _000489_, _000490_, _000491_, _000492_, _000493_, _000494_, _000495_, _000496_, _000497_, _000498_, _000499_, _000500_, _000501_, _000502_, _000503_, _000504_, _000505_, _000506_, _000507_, _000508_, _000509_, _000510_, _000511_, _000512_, _000513_, _000514_, _000515_, _000516_, _000517_, _000518_, _000519_, _000520_, _000521_, _000522_, _000523_, _000524_, _000525_, _000526_, _000527_, _000528_, _000529_, _000530_, _000531_, _000532_, _000533_, _000534_, _000535_, _000536_, _000537_, _000538_, _000539_, _000540_, _000541_, _000542_, _000543_, _000544_, _000545_, _000546_, _000547_, _000548_, _000549_, _000550_, _000551_, _000552_, _000553_, _000554_, _000555_, _000556_, _000557_, _000558_, _000559_, _000560_, _000561_, _000562_, _000563_, _000564_, _000565_, _000566_, _000567_, _000568_, _000569_, _000570_, _000571_, _000572_, _000573_, _000574_, _000575_, _000576_, _000577_, _000578_, _000579_, _000580_, _000581_, _000582_, _000583_, _000584_, _000585_, _000586_, _000587_, _000588_, _000589_, _000590_, _000591_, _000592_, _000593_, _000594_, _000595_, _000596_, _000597_, _000598_, _000599_, _000600_, _000601_, _000602_, _000603_, _000604_, _000605_, _000606_, _000607_, _000608_, _000609_, _000610_, _000611_, _000612_, _000613_, _000614_, _000615_, _000616_, _000617_, _000618_, _000619_, _000620_, _000621_, _000622_, _000623_, _000624_, _000625_, _000626_, _000627_, _000628_, _000629_, _000630_, _000631_, _000632_, _000633_, _000634_, _000635_, _000636_, _000637_, _000638_, _000639_, _000640_, _000641_, _000642_, _000643_, _000644_, _000645_, _000646_, _000647_, _000648_, _000649_, _000650_, _000651_, _000652_, _000653_, _000654_, _000655_, _000656_, _000657_, _000658_, _000659_, _000660_, _000661_, _000662_, _000663_, _000664_, _000665_, _000666_, _000667_, _000668_, _000669_, _000670_, _000671_, _000672_, _000673_, _000674_, _000675_, _000676_, _000677_, _000678_, _000679_, _000680_, _000681_, _000682_, _000683_, _000684_, _000685_, _000686_, _000687_, _000688_, _000689_, _000690_, _000691_, _000692_, _000693_, _000694_, _000695_, _000696_, _000697_, _000698_, _000699_, _000700_, _000701_, _000702_, _000703_, _000704_, _000705_, _000706_, _000707_, _000708_, _000709_, _000710_, _000711_, _000712_, _000713_, _000714_, _000715_, _000716_, _000717_, _000718_, _000719_, _000720_, _000721_, _000722_, _000723_, _000724_, _000725_, _000726_, _000727_, _000728_, _000729_, _000730_, _000731_, _000732_, _000733_, _000734_, _000735_, _000736_, _000737_, _000738_, _000739_, _000740_, _000741_, _000742_, _000743_, _000744_, _000745_, _000746_, _000747_, _000748_, _000749_, _000750_, _000751_, _000752_, _000753_, _000754_, _000755_, _000756_, _000757_, _000758_, _000759_, _000760_, _000761_, _000762_, _000763_, _000764_, _000765_, _000766_, _000767_, _000768_, _000769_, _000770_, _000771_, _000772_, _000773_, _000774_, _000775_, _000776_, _000777_, _000778_, _000779_, _000780_, _000781_, _000782_, _000783_, _000784_, _000785_, _000786_, _000787_, _000788_, _000789_, _000790_, _000791_, _000792_, _000793_, _000794_, _000795_, _000796_, _000797_, _000798_, _000799_, _000800_, _000801_, _000802_, _000803_, _000804_, _000805_, _000806_, _000807_, _000808_, _000809_, _000810_, _000811_, _000812_, _000813_, _000814_, _000815_, _000816_, _000817_, _000818_, _000819_, _000820_, _000821_, _000822_, _000823_, _000824_, _000825_, _000826_, _000827_, _000828_, _000829_, _000830_, _000831_, _000832_, _000833_, _000834_, _000835_, _000836_, _000837_, _000838_, _000839_, _000840_, _000841_, _000842_, _000843_, _000844_, _000845_, _000846_, _000847_, _000848_, _000849_, _000850_, _000851_, _000852_, _000853_, _000854_, _000855_, _000856_, _000857_, _000858_, _000859_, _000860_, _000861_, _000862_, _000863_, _000864_, _000865_, _000866_, _000867_, _000868_, _000869_, _000870_, _000871_, _000872_, _000873_, _000874_, _000875_, _000876_, _000877_, _000878_, _000879_, _000880_, _000881_, _000882_, _000883_, _000884_, _000885_, _000886_, _000887_, _000888_, _000889_, _000890_, _000891_, _000892_, _000893_, _000894_, _000895_, _000896_, _000897_, _000898_, _000899_, _000900_, _000901_, _000902_, _000903_, _000904_, _000905_, _000906_, _000907_, _000908_, _000909_, _000910_, _000911_, _000912_, _000913_, _000914_, _000915_, _000916_, _000917_, _000918_, _000919_, _000920_, _000921_, _000922_, _000923_, _000924_, _000925_, _000926_, _000927_, _000928_, _000929_, _000930_, _000931_, _000932_, _000933_, _000934_, _000935_, _000936_, _000937_, _000938_, _000939_, _000940_, _000941_, _000942_, _000943_, _000944_, _000945_, _000946_, _000947_, _000948_, _000949_, _000950_, _000951_, _000952_, _000953_, _000954_, _000955_, _000956_, _000957_, _000958_, _000959_, _000960_, _000961_, _000962_, _000963_, _000964_, _000965_, _000966_, _000967_, _000968_, _000969_, _000970_, _000971_, _000972_, _000973_, _000974_, _000975_, _000976_, _000977_, _000978_, _000979_, _000980_, _000981_, _000982_, _000983_, _000984_, _000985_, _000986_, _000987_, _000988_, _000989_, _000990_, _000991_, _000992_, _000993_, _000994_, _000995_, _000996_, _000997_, _000998_, _000999_, _001000_, _001001_, _001002_, _001003_, _001004_, _001005_, _001006_, _001007_, _001008_, _001009_, _001010_, _001011_, _001012_, _001013_, _001014_, _001015_, _001016_, _001017_, _001018_, _001019_, _001020_, _001021_, _001022_, _001023_, _001024_, _001025_, _001026_, _001027_, _001028_, _001029_, _001030_, _001031_, _001032_, _001033_, _001034_, _001035_, _001036_, _001037_, _001038_, _001039_, _001040_, _001041_, _001042_, _001043_, _001044_, _001045_, _001046_, _001047_, _001048_, _001049_, _001050_, _001051_, _001052_, _001053_, _001054_, _001055_, _001056_, _001057_, _001058_, _001059_, _001060_, _001061_, _001062_, _001063_, _001064_, _001065_, _001066_, _001067_, _001068_, _001069_, _001070_, _001071_, _001072_, _001073_, _001074_, _001075_, _001076_, _001077_, _001078_, _001079_, _001080_, _001081_, _001082_, _001083_, _001084_, _001085_, _001086_, _001087_, _001088_, _001089_, _001090_, _001091_, _001092_, _001093_, _001094_, _001095_, _001096_, _001097_, _001098_, _001099_, _001100_, _001101_, _001102_, _001103_, _001104_, _001105_, _001106_, _001107_, _001108_, _001109_, _001110_, _001111_, _001112_, _001113_, _001114_, _001115_, _001116_, _001117_, _001118_, _001119_, _001120_, _001121_, _001122_, _001123_, _001124_, _001125_, _001126_, _001127_, _001128_, _001129_, _001130_, _001131_, _001132_, _001133_, _001134_, _001135_, _001136_, _001137_, _001138_, _001139_, _001140_, _001141_, _001142_, _001143_, _001144_, _001145_, _001146_, _001147_, _001148_, _001149_, _001150_, _001151_, _001152_, _001153_, _001154_, _001155_, _001156_, _001157_, _001158_, _001159_, _001160_, _001161_, _001162_, _001163_, _001164_, _001165_, _001166_, _001167_, _001168_, _001169_, _001170_, _001171_, _001172_, _001173_, _001174_, _001175_, _001176_, _001177_, _001178_, _001179_, _001180_, _001181_, _001182_, _001183_, _001184_, _001185_, _001186_, _001187_, _001188_, _001189_, _001190_, _001191_, _001192_, _001193_, _001194_, _001195_, _001196_, _001197_, _001198_, _001199_, _001200_, _001201_, _001202_, _001203_, _001204_, _001205_, _001206_, _001207_, _001208_, _001209_, _001210_, _001211_, _001212_, _001213_, _001214_, _001215_, _001216_, _001217_, _001218_, _001219_, _001220_, _001221_, _001222_, _001223_, _001224_, _001225_, _001226_, _001227_, _001228_, _001229_, _001230_, _001231_, _001232_, _001233_, _001234_, _001235_, _001236_, _001237_, _001238_, _001239_, _001240_, _001241_, _001242_, _001243_, _001244_, _001245_, _001246_, _001247_, _001248_, _001249_, _001250_, _001251_, _001252_, _001253_, _001254_, _001255_, _001256_, _001257_, _001258_, _001259_, _001260_, _001261_, _001262_, _001263_, _001264_, _001265_, _001266_, _001267_, _001268_, _001269_, _001270_, _001271_, _001272_, _001273_, _001274_, _001275_, _001276_, _001277_, _001278_, _001279_, _001280_, _001281_, _001282_, _001283_, _001284_, _001285_, _001286_, _001287_, _001288_, _001289_, _001290_, _001291_, _001292_, _001293_, _001294_, _001295_, _001296_, _001297_, _001298_, _001299_, _001300_, _001301_, _001302_, _001303_, _001304_, _001305_, _001306_, _001307_, _001308_, _001309_, _001310_, _001311_, _001312_, _001313_, _001314_, _001315_, _001316_, _001317_, _001318_, _001319_, _001320_, _001321_, _001322_, _001323_, _001324_, _001325_, _001326_, _001327_, _001328_, _001329_, _001330_, _001331_, _001332_, _001333_, _001334_, _001335_, _001336_, _001337_, _001338_, _001339_, _001340_, _001341_, _001342_, _001343_, _001344_, _001345_, _001346_, _001347_, _001348_, _001349_, _001350_, _001351_, _001352_, _001353_, _001354_, _001355_, _001356_, _001357_, _001358_, _001359_, _001360_, _001361_, _001362_, _001363_, _001364_, _001365_, _001366_, _001367_, _001368_, _001369_, _001370_, _001371_, _001372_, _001373_, _001374_, _001375_, _001376_, _001377_, _001378_, _001379_, _001380_, _001381_, _001382_, _001383_, _001384_, _001385_, _001386_, _001387_, _001388_, _001389_, _001390_, _001391_, _001392_, _001393_, _001394_, _001395_, _001396_, _001397_, _001398_, _001399_, _001400_, _001401_, _001402_, _001403_, _001404_, _001405_, _001406_, _001407_, _001408_, _001409_, _001410_, _001411_, _001412_, _001413_, _001414_, _001415_, _001416_, _001417_, _001418_, _001419_, _001420_, _001421_, _001422_, _001423_, _001424_, _001425_, _001426_, _001427_, _001428_, _001429_, _001430_, _001431_, _001432_, _001433_, _001434_, _001435_, _001436_, _001437_, _001438_, _001439_, _001440_, _001441_, _001442_, _001443_, _001444_, _001445_, _001446_, _001447_, _001448_, _001449_, _001450_, _001451_, _001452_, _001453_, _001454_, _001455_, _001456_, _001457_, _001458_, _001459_, _001460_, _001461_, _001462_, _001463_, _001464_, _001465_, _001466_, _001467_, _001468_, _001469_, _001470_, _001471_, _001472_, _001473_, _001474_, _001475_, _001476_, _001477_, _001478_, _001479_, _001480_, _001481_, _001482_, _001483_, _001484_, _001485_, _001486_, _001487_, _001488_, _001489_, _001490_, _001491_, _001492_, _001493_, _001494_, _001495_, _001496_, _001497_, _001498_, _001499_, _001500_, _001501_, _001502_, _001503_, _001504_, _001505_, _001506_, _001507_, _001508_, _001509_, _001510_, _001511_, _001512_, _001513_, _001514_, _001515_, _001516_, _001517_, _001518_, _001519_, _001520_, _001521_, _001522_, _001523_, _001524_, _001525_, _001526_, _001527_, _001528_, _001529_, _001530_, _001531_, _001532_, _001533_, _001534_, _001535_, _001536_, _001537_, _001538_, _001539_, _001540_, _001541_, _001542_, _001543_, _001544_, _001545_, _001546_, _001547_, _001548_, _001549_, _001550_, _001551_, _001552_, _001553_, _001554_, _001555_, _001556_, _001557_, _001558_, _001559_, _001560_, _001561_, _001562_, _001563_, _001564_, _001565_, _001566_, _001567_, _001568_, _001569_, _001570_, _001571_, _001572_, _001573_, _001574_, _001575_, _001576_, _001577_, _001578_, _001579_, _001580_, _001581_, _001582_, _001583_, _001584_, _001585_, _001586_, _001587_, _001588_, _001589_, _001590_, _001591_, _001592_, _001593_, _001594_, _001595_, _001596_, _001597_, _001598_, _001599_, _001600_, _001601_, _001602_, _001603_, _001604_, _001605_, _001606_, _001607_, _001608_, _001609_, _001610_, _001611_, _001612_, _001613_, _001614_, _001615_, _001616_, _001617_, _001618_, _001619_, _001620_, _001621_, _001622_, _001623_, _001624_, _001625_, _001626_, _001627_, _001628_, _001629_, _001630_, _001631_, _001632_, _001633_, _001634_, _001635_, _001636_, _001637_, _001638_, _001639_, _001640_, _001641_, _001642_, _001643_, _001644_, _001645_, _001646_, _001647_, _001648_, _001649_, _001650_, _001651_, _001652_, _001653_, _001654_, _001655_, _001656_, _001657_, _001658_, _001659_, _001660_, _001661_, _001662_, _001663_, _001664_, _001665_, _001666_, _001667_, _001668_, _001669_, _001670_, _001671_, _001672_, _001673_, _001674_, _001675_, _001676_, _001677_, _001678_, _001679_, _001680_, _001681_, _001682_, _001683_, _001684_, _001685_, _001686_, _001687_, _001688_, _001689_, _001690_, _001691_, _001692_, _001693_, _001694_, _001695_, _001696_, _001697_, _001698_, _001699_, _001700_, _001701_, _001702_, _001703_, _001704_, _001705_, _001706_, _001707_, _001708_, _001709_, _001710_, _001711_, _001712_, _001713_, _001714_, _001715_, _001716_, _001717_, _001718_, _001719_, _001720_, _001721_, _001722_, _001723_, _001724_, _001725_, _001726_, _001727_, _001728_, _001729_, _001730_, _001731_, _001732_, _001733_, _001734_, _001735_, _001736_, _001737_, _001738_, _001739_, _001740_, _001741_, _001742_, _001743_, _001744_, _001745_, _001746_, _001747_, _001748_, _001749_, _001750_, _001751_, _001752_, _001753_, _001754_, _001755_, _001756_, _001757_, _001758_, _001759_, _001760_, _001761_, _001762_, _001763_, _001764_, _001765_, _001766_, _001767_, _001768_, _001769_, _001770_, _001771_, _001772_, _001773_, _001774_, _001775_, _001776_, _001777_, _001778_, _001779_, _001780_, _001781_, _001782_, _001783_, _001784_, _001785_, _001786_, _001787_, _001788_, _001789_, _001790_, _001791_, _001792_, _001793_, _001794_, _001795_, _001796_, _001797_, _001798_, _001799_, _001800_, _001801_, _001802_, _001803_, _001804_, _001805_, _001806_, _001807_, _001808_, _001809_, _001810_, _001811_, _001812_, _001813_, _001814_, _001815_, _001816_, _001817_, _001818_, _001819_, _001820_, _001821_, _001822_, _001823_, _001824_, _001825_, _001826_, _001827_, _001828_, _001829_, _001830_, _001831_, _001832_, _001833_, _001834_, _001835_, _001836_, _001837_, _001838_, _001839_, _001840_, _001841_, _001842_, _001843_, _001844_, _001845_, _001846_, _001847_, _001848_, _001849_, _001850_, _001851_, _001852_, _001853_, _001854_, _001855_, _001856_, _001857_, _001858_, _001859_, _001860_, _001861_, _001862_, _001863_, _001864_, _001865_, _001866_, _001867_, _001868_, _001869_, _001870_, _001871_, _001872_, _001873_, _001874_, _001875_, _001876_, _001877_, _001878_, _001879_, _001880_, _001881_, _001882_, _001883_, _001884_, _001885_, _001886_, _001887_, _001888_, _001889_, _001890_, _001891_, _001892_, _001893_, _001894_, _001895_, _001896_, _001897_, _001898_, _001899_, _001900_, _001901_, _001902_, _001903_, _001904_, _001905_, _001906_, _001907_, _001908_, _001909_, _001910_, _001911_, _001912_, _001913_, _001914_, _001915_, _001916_, _001917_, _001918_, _001919_, _001920_, _001921_, _001922_, _001923_, _001924_, _001925_, _001926_, _001927_, _001928_, _001929_, _001930_, _001931_, _001932_, _001933_, _001934_, _001935_, _001936_, _001937_, _001938_, _001939_, _001940_, _001941_, _001942_, _001943_, _001944_, _001945_, _001946_, _001947_, _001948_, _001949_, _001950_, _001951_, _001952_, _001953_, _001954_, _001955_, _001956_, _001957_, _001958_, _001959_, _001960_, _001961_, _001962_, _001963_, _001964_, _001965_, _001966_, _001967_, _001968_, _001969_, _001970_, _001971_, _001972_, _001973_, _001974_, _001975_, _001976_, _001977_, _001978_, _001979_, _001980_, _001981_, _001982_, _001983_, _001984_, _001985_, _001986_, _001987_, _001988_, _001989_, _001990_, _001991_, _001992_, _001993_, _001994_, _001995_, _001996_, _001997_, _001998_, _001999_, _002000_, _002001_, _002002_, _002003_, _002004_, _002005_, _002006_, _002007_, _002008_, _002009_, _002010_, _002011_, _002012_, _002013_, _002014_, _002015_, _002016_, _002017_, _002018_, _002019_, _002020_, _002021_, _002022_, _002023_, _002024_, _002025_, _002026_, _002027_, _002028_, _002029_, _002030_, _002031_, _002032_, _002033_, _002034_, _002035_, _002036_, _002037_, _002038_, _002039_, _002040_, _002041_, _002042_, _002043_, _002044_, _002045_, _002046_, _002047_, _002048_, _002049_, _002050_, _002051_, _002052_, _002053_, _002054_, _002055_, _002056_, _002057_, _002058_, _002059_, _002060_, _002061_, _002062_, _002063_, _002064_, _002065_, _002066_, _002067_, _002068_, _002069_, _002070_, _002071_, _002072_, _002073_, _002074_, _002075_, _002076_, _002077_, _002078_, _002079_, _002080_, _002081_, _002082_, _002083_, _002084_, _002085_, _002086_, _002087_, _002088_, _002089_, _002090_, _002091_, _002092_, _002093_, _002094_, _002095_, _002096_, _002097_, _002098_, _002099_, _002100_, _002101_, _002102_, _002103_, _002104_, _002105_, _002106_, _002107_, _002108_, _002109_, _002110_, _002111_, _002112_, _002113_, _002114_, _002115_, _002116_, _002117_, _002118_, _002119_, _002120_, _002121_, _002122_, _002123_, _002124_, _002125_, _002126_, _002127_, _002128_, _002129_, _002130_, _002131_, _002132_, _002133_, _002134_, _002135_, _002136_, _002137_, _002138_, _002139_, _002140_, _002141_, _002142_, _002143_, _002144_, _002145_, _002146_, _002147_, _002148_, _002149_, _002150_, _002151_, _002152_, _002153_, _002154_, _002155_, _002156_, _002157_, _002158_, _002159_, _002160_, _002161_, _002162_, _002163_, _002164_, _002165_, _002166_, _002167_, _002168_, _002169_, _002170_, _002171_, _002172_, _002173_, _002174_, _002175_, _002176_, _002177_, _002178_, _002179_, _002180_, _002181_, _002182_, _002183_, _002184_, _002185_, _002186_, _002187_, _002188_, _002189_, _002190_, _002191_, _002192_, _002193_, _002194_, _002195_, _002196_, _002197_, _002198_, _002199_, _002200_, _002201_, _002202_, _002203_, _002204_, _002205_, _002206_, _002207_, _002208_, _002209_, _002210_, _002211_, _002212_, _002213_, _002214_, _002215_, _002216_, _002217_, _002218_, _002219_, _002220_, _002221_, _002222_, _002223_, _002224_, _002225_, _002226_, _002227_, _002228_, _002229_, _002230_, _002231_, _002232_, _002233_, _002234_, _002235_, _002236_, _002237_, _002238_, _002239_, _002240_, _002241_, _002242_, _002243_, _002244_, _002245_, _002246_, _002247_, _002248_, _002249_, _002250_, _002251_, _002252_, _002253_, _002254_, _002255_, _002256_, _002257_, _002258_, _002259_, _002260_, _002261_, _002262_, _002263_, _002264_, _002265_, _002266_, _002267_, _002268_, _002269_, _002270_, _002271_, _002272_, _002273_, _002274_, _002275_, _002276_, _002277_, _002278_, _002279_, _002280_, _002281_, _002282_, _002283_, _002284_, _002285_, _002286_, _002287_, _002288_, _002289_, _002290_, _002291_, _002292_, _002293_, _002294_, _002295_, _002296_, _002297_, _002298_, _002299_, _002300_, _002301_, _002302_, _002303_, _002304_, _002305_, _002306_, _002307_, _002308_, _002309_, _002310_, _002311_, _002312_, _002313_, _002314_, _002315_, _002316_, _002317_, _002318_, _002319_, _002320_, _002321_, _002322_, _002323_, _002324_, _002325_, _002326_, _002327_, _002328_, _002329_, _002330_, _002331_, _002332_, _002333_, _002334_, _002335_, _002336_, _002337_, _002338_, _002339_, _002340_, _002341_, _002342_, _002343_, _002344_, _002345_, _002346_, _002347_, _002348_, _002349_, _002350_, _002351_, _002352_, _002353_, _002354_, _002355_, _002356_, _002357_, _002358_, _002359_, _002360_, _002361_, _002362_, _002363_, _002364_, _002365_, _002366_, _002367_, _002368_, _002369_, _002370_, _002371_, _002372_, _002373_, _002374_, _002375_, _002376_, _002377_, _002378_, _002379_, _002380_, _002381_, _002382_, _002383_, _002384_, _002385_, _002386_, _002387_, _002388_, _002389_, _002390_, _002391_, _002392_, _002393_, _002394_, _002395_, _002396_, _002397_, _002398_, _002399_, _002400_, _002401_, _002402_, _002403_, _002404_, _002405_, _002406_, _002407_, _002408_, _002409_, _002410_, _002411_, _002412_, _002413_, _002414_, _002415_, _002416_, _002417_, _002418_, _002419_, _002420_, _002421_, _002422_, _002423_, _002424_, _002425_, _002426_, _002427_, _002428_, _002429_, _002430_, _002431_, _002432_, _002433_, _002434_, _002435_, _002436_, _002437_, _002438_, _002439_, _002440_, _002441_, _002442_, _002443_, _002444_, _002445_, _002446_, _002447_, _002448_, _002449_, _002450_, _002451_, _002452_, _002453_, _002454_, _002455_, _002456_, _002457_, _002458_, _002459_, _002460_, _002461_, _002462_, _002463_, _002464_, _002465_, _002466_, _002467_, _002468_, _002469_, _002470_, _002471_, _002472_, _002473_, _002474_, _002475_, _002476_, _002477_, _002478_, _002479_, _002480_, _002481_, _002482_, _002483_, _002484_, _002485_, _002486_, _002487_, _002488_, _002489_, _002490_, _002491_, _002492_, _002493_, _002494_, _002495_, _002496_, _002497_, _002498_, _002499_, _002500_, _002501_, _002502_, _002503_, _002504_, _002505_, _002506_, _002507_, _002508_, _002509_, _002510_, _002511_, _002512_, _002513_, _002514_, _002515_, _002516_, _002517_, _002518_, _002519_, _002520_, _002521_, _002522_, _002523_, _002524_, _002525_, _002526_, _002527_, _002528_, _002529_, _002530_, _002531_, _002532_, _002533_, _002534_, _002535_, _002536_, _002537_, _002538_, _002539_, _002540_, _002541_, _002542_, _002543_, _002544_, _002545_, _002546_, _002547_, _002548_, _002549_, _002550_, _002551_, _002552_, _002553_, _002554_, _002555_, _002556_, _002557_, _002558_, _002559_, _002560_, _002561_, _002562_, _002563_, _002564_, _002565_, _002566_, _002567_, _002568_, _002569_, _002570_, _002571_, _002572_, _002573_, _002574_, _002575_, _002576_, _002577_, _002578_, _002579_, _002580_, _002581_, _002582_, _002583_, _002584_, _002585_, _002586_, _002587_, _002588_, _002589_, _002590_, _002591_, _002592_, _002593_, _002594_, _002595_, _002596_, _002597_, _002598_, _002599_, _002600_, _002601_, _002602_, _002603_, _002604_, _002605_, _002606_, _002607_, _002608_, _002609_, _002610_, _002611_, _002612_, _002613_, _002614_, _002615_, _002616_, _002617_, _002618_, _002619_, _002620_, _002621_, _002622_, _002623_, _002624_, _002625_, _002626_, _002627_, _002628_, _002629_, _002630_, _002631_, _002632_, _002633_, _002634_, _002635_, _002636_, _002637_, _002638_, _002639_, _002640_, _002641_, _002642_, _002643_, _002644_, _002645_, _002646_, _002647_, _002648_, _002649_, _002650_, _002651_, _002652_, _002653_, _002654_, _002655_, _002656_, _002657_, _002658_, _002659_, _002660_, _002661_, _002662_, _002663_, _002664_, _002665_, _002666_, _002667_, _002668_, _002669_, _002670_, _002671_, _002672_, _002673_, _002674_, _002675_, _002676_, _002677_, _002678_, _002679_, _002680_, _002681_, _002682_, _002683_, _002684_, _002685_, _002686_, _002687_, _002688_, _002689_, _002690_, _002691_, _002692_, _002693_, _002694_, _002695_, _002696_, _002697_, _002698_, _002699_, _002700_, _002701_, _002702_, _002703_, _002704_, _002705_, _002706_, _002707_, _002708_, _002709_, _002710_, _002711_, _002712_, _002713_, _002714_, _002715_, _002716_, _002717_, _002718_, _002719_, _002720_, _002721_, _002722_, _002723_, _002724_, _002725_, _002726_, _002727_, _002728_, _002729_, _002730_, _002731_, _002732_, _002733_, _002734_, _002735_, _002736_, _002737_, _002738_, _002739_, _002740_, _002741_, _002742_, _002743_, _002744_, _002745_, _002746_, _002747_, _002748_, _002749_, _002750_, _002751_, _002752_, _002753_, _002754_, _002755_, _002756_, _002757_, _002758_, _002759_, _002760_, _002761_, _002762_, _002763_, _002764_, _002765_, _002766_, _002767_, _002768_, _002769_, _002770_, _002771_, _002772_, _002773_, _002774_, _002775_, _002776_, _002777_, _002778_, _002779_, _002780_, _002781_, _002782_, _002783_, _002784_, _002785_, _002786_, _002787_, _002788_, _002789_, _002790_, _002791_, _002792_, _002793_, _002794_, _002795_, _002796_, _002797_, _002798_, _002799_, _002800_, _002801_, _002802_, _002803_, _002804_, _002805_, _002806_, _002807_, _002808_, _002809_, _002810_, _002811_, _002812_, _002813_, _002814_, _002815_, _002816_, _002817_, _002818_, _002819_, _002820_, _002821_, _002822_, _002823_, _002824_, _002825_, _002826_, _002827_, _002828_, _002829_, _002830_, _002831_, _002832_, _002833_, _002834_, _002835_, _002836_, _002837_, _002838_, _002839_, _002840_, _002841_, _002842_, _002843_, _002844_, _002845_, _002846_, _002847_, _002848_, _002849_, _002850_, _002851_, _002852_, _002853_, _002854_, _002855_, _002856_, _002857_, _002858_, _002859_, _002860_, _002861_, _002862_, _002863_, _002864_, _002865_, _002866_, _002867_, _002868_, _002869_, _002870_, _002871_, _002872_, _002873_, _002874_, _002875_, _002876_, _002877_, _002878_, _002879_, _002880_, _002881_, _002882_, _002883_, _002884_, _002885_, _002886_, _002887_, _002888_, _002889_, _002890_, _002891_, _002892_, _002893_, _002894_, _002895_, _002896_, _002897_, _002898_, _002899_, _002900_, _002901_, _002902_, _002903_, _002904_, _002905_, _002906_, _002907_, _002908_, _002909_, _002910_, _002911_, _002912_, _002913_, _002914_, _002915_, _002916_, _002917_, _002918_, _002919_, _002920_, _002921_, _002922_, _002923_, _002924_, _002925_, _002926_, _002927_, _002928_, _002929_, _002930_, _002931_, _002932_, _002933_, _002934_, _002935_, _002936_, _002937_, _002938_, _002939_, _002940_, _002941_, _002942_, _002943_, _002944_, _002945_, _002946_, _002947_, _002948_, _002949_, _002950_, _002951_, _002952_, _002953_, _002954_, _002955_, _002956_, _002957_, _002958_, _002959_, _002960_, _002961_, _002962_, _002963_, _002964_, _002965_, _002966_, _002967_, _002968_, _002969_, _002970_, _002971_, _002972_, _002973_, _002974_, _002975_, _002976_, _002977_, _002978_, _002979_, _002980_, _002981_, _002982_, _002983_, _002984_, _002985_, _002986_, _002987_, _002988_, _002989_, _002990_, _002991_, _002992_, _002993_, _002994_, _002995_, _002996_, _002997_, _002998_, _002999_, _003000_, _003001_, _003002_, _003003_, _003004_, _003005_, _003006_, _003007_, _003008_, _003009_, _003010_, _003011_, _003012_, _003013_, _003014_, _003015_, _003016_, _003017_, _003018_, _003019_, _003020_, _003021_, _003022_, _003023_, _003024_, _003025_, _003026_, _003027_, _003028_, _003029_, _003030_, _003031_, _003032_, _003033_, _003034_, _003035_, _003036_, _003037_, _003038_, _003039_, _003040_, _003041_, _003042_, _003043_, _003044_, _003045_, _003046_, _003047_, _003048_, _003049_, _003050_, _003051_, _003052_, _003053_, _003054_, _003055_, _003056_, _003057_, _003058_, _003059_, _003060_, _003061_, _003062_, _003063_, _003064_, _003065_, _003066_, _003067_, _003068_, _003069_, _003070_, _003071_, _003072_, _003073_, _003074_, _003075_, _003076_, _003077_, _003078_, _003079_, _003080_, _003081_, _003082_, _003083_, _003084_, _003085_, _003086_, _003087_, _003088_, _003089_, _003090_, _003091_, _003092_, _003093_, _003094_, _003095_, _003096_, _003097_, _003098_, _003099_, _003100_, _003101_, _003102_, _003103_, _003104_, _003105_, _003106_, _003107_, _003108_, _003109_, _003110_, _003111_, _003112_, _003113_, _003114_, _003115_, _003116_, _003117_, _003118_, _003119_, _003120_, _003121_, _003122_, _003123_, _003124_, _003125_, _003126_, _003127_, _003128_, _003129_, _003130_, _003131_, _003132_, _003133_, _003134_, _003135_, _003136_, _003137_, _003138_, _003139_, _003140_, _003141_, _003142_, _003143_, _003144_, _003145_, _003146_, _003147_, _003148_, _003149_, _003150_, _003151_, _003152_, _003153_, _003154_, _003155_, _003156_, _003157_, _003158_, _003159_, _003160_, _003161_, _003162_, _003163_, _003164_, _003165_, _003166_, _003167_, _003168_, _003169_, _003170_, _003171_, _003172_, _003173_, _003174_, _003175_, _003176_, _003177_, _003178_, _003179_, _003180_, _003181_, _003182_, _003183_, _003184_, _003185_, _003186_, _003187_, _003188_, _003189_, _003190_, _003191_, _003192_, _003193_, _003194_, _003195_, _003196_, _003197_, _003198_, _003199_, _003200_, _003201_, _003202_, _003203_, _003204_, _003205_, _003206_, _003207_, _003208_, _003209_, _003210_, _003211_, _003212_, _003213_, _003214_, _003215_, _003216_, _003217_, _003218_, _003219_, _003220_, _003221_, _003222_, _003223_, _003224_, _003225_, _003226_, _003227_, _003228_, _003229_, _003230_, _003231_, _003232_, _003233_, _003234_, _003235_, _003236_, _003237_, _003238_, _003239_, _003240_, _003241_, _003242_, _003243_, _003244_, _003245_, _003246_, _003247_, _003248_, _003249_, _003250_, _003251_, _003252_, _003253_, _003254_, _003255_, _003256_, _003257_, _003258_, _003259_, _003260_, _003261_, _003262_, _003263_, _003264_, _003265_, _003266_, _003267_, _003268_, _003269_, _003270_, _003271_, _003272_, _003273_, _003274_, _003275_, _003276_, _003277_, _003278_, _003279_, _003280_, _003281_, _003282_, _003283_, _003284_, _003285_, _003286_, _003287_, _003288_, _003289_, _003290_, _003291_, _003292_, _003293_, _003294_, _003295_, _003296_, _003297_, _003298_, _003299_, _003300_, _003301_, _003302_, _003303_, _003304_, _003305_, _003306_, _003307_, _003308_, _003309_, _003310_, _003311_, _003312_, _003313_, _003314_, _003315_, _003316_, _003317_, _003318_, _003319_, _003320_, _003321_, _003322_, _003323_, _003324_, _003325_, _003326_, _003327_, _003328_, _003329_, _003330_, _003331_, _003332_, _003333_, _003334_, _003335_, _003336_, _003337_, _003338_, _003339_, _003340_, _003341_, _003342_, _003343_, _003344_, _003345_, _003346_, _003347_, _003348_, _003349_, _003350_, _003351_, _003352_, _003353_, _003354_, _003355_, _003356_, _003357_, _003358_, _003359_, _003360_, _003361_, _003362_, _003363_, _003364_, _003365_, _003366_, _003367_, _003368_, _003369_, _003370_, _003371_, _003372_, _003373_, _003374_, _003375_, _003376_, _003377_, _003378_, _003379_, _003380_, _003381_, _003382_, _003383_, _003384_, _003385_, _003386_, _003387_, _003388_, _003389_, _003390_, _003391_, _003392_, _003393_, _003394_, _003395_, _003396_, _003397_, _003398_, _003399_, _003400_, _003401_, _003402_, _003403_, _003404_, _003405_, _003406_, _003407_, _003408_, _003409_, _003410_, _003411_, _003412_, _003413_, _003414_, _003415_, _003416_, _003417_, _003418_, _003419_, _003420_, _003421_, _003422_, _003423_, _003424_, _003425_, _003426_, _003427_, _003428_, _003429_, _003430_, _003431_, _003432_, _003433_, _003434_, _003435_, _003436_, _003437_, _003438_, _003439_, _003440_, _003441_, _003442_, _003443_, _003444_, _003445_, _003446_, _003447_, _003448_, _003449_, _003450_, _003451_, _003452_, _003453_, _003454_, _003455_, _003456_, _003457_, _003458_, _003459_, _003460_, _003461_, _003462_, _003463_, _003464_, _003465_, _003466_, _003467_, _003468_, _003469_, _003470_, _003471_, _003472_, _003473_, _003474_, _003475_, _003476_, _003477_, _003478_, _003479_, _003480_, _003481_, _003482_, _003483_, _003484_, _003485_, _003486_, _003487_, _003488_, _003489_, _003490_, _003491_, _003492_, _003493_, _003494_, _003495_, _003496_, _003497_, _003498_, _003499_, _003500_, _003501_, _003502_, _003503_, _003504_, _003505_, _003506_, _003507_, _003508_, _003509_, _003510_, _003511_, _003512_, _003513_, _003514_, _003515_, _003516_, _003517_, _003518_, _003519_, _003520_, _003521_, _003522_, _003523_, _003524_, _003525_, _003526_, _003527_, _003528_, _003529_, _003530_, _003531_, _003532_, _003533_, _003534_, _003535_, _003536_, _003537_, _003538_, _003539_, _003540_, _003541_, _003542_, _003543_, _003544_, _003545_, _003546_, _003547_, _003548_, _003549_, _003550_, _003551_, _003552_, _003553_, _003554_, _003555_, _003556_, _003557_, _003558_, _003559_, _003560_, _003561_, _003562_, _003563_, _003564_, _003565_, _003566_, _003567_, _003568_, _003569_, _003570_, _003571_, _003572_, _003573_, _003574_, _003575_, _003576_, _003577_, _003578_, _003579_, _003580_, _003581_, _003582_, _003583_, _003584_, _003585_, _003586_, _003587_, _003588_, _003589_, _003590_, _003591_, _003592_, _003593_, _003594_, _003595_, _003596_, _003597_, _003598_, _003599_, _003600_, _003601_, _003602_, _003603_, _003604_, _003605_, _003606_, _003607_, _003608_, _003609_, _003610_, _003611_, _003612_, _003613_, _003614_, _003615_, _003616_, _003617_, _003618_, _003619_, _003620_, _003621_, _003622_, _003623_, _003624_, _003625_, _003626_, _003627_, _003628_, _003629_, _003630_, _003631_, _003632_, _003633_, _003634_, _003635_, _003636_, _003637_, _003638_, _003639_, _003640_, _003641_, _003642_, _003643_, _003644_, _003645_, _003646_, _003647_, _003648_, _003649_, _003650_, _003651_, _003652_, _003653_, _003654_, _003655_, _003656_, _003657_, _003658_, _003659_, _003660_, _003661_, _003662_, _003663_, _003664_, _003665_, _003666_, _003667_, _003668_, _003669_, _003670_, _003671_, _003672_, _003673_, _003674_, _003675_, _003676_, _003677_, _003678_, _003679_, _003680_, _003681_, _003682_, _003683_, _003684_, _003685_, _003686_, _003687_, _003688_, _003689_, _003690_, _003691_, _003692_, _003693_, _003694_, _003695_, _003696_, _003697_, _003698_, _003699_, _003700_, _003701_, _003702_, _003703_, _003704_, _003705_, _003706_, _003707_, _003708_, _003709_, _003710_, _003711_, _003712_, _003713_, _003714_, _003715_, _003716_, _003717_, _003718_, _003719_, _003720_, _003721_, _003722_, _003723_, _003724_, _003725_, _003726_, _003727_, _003728_, _003729_, _003730_, _003731_, _003732_, _003733_, _003734_, _003735_, _003736_, _003737_, _003738_, _003739_, _003740_, _003741_, _003742_, _003743_, _003744_, _003745_, _003746_, _003747_, _003748_, _003749_, _003750_, _003751_, _003752_, _003753_, _003754_, _003755_, _003756_, _003757_, _003758_, _003759_, _003760_, _003761_, _003762_, _003763_, _003764_, _003765_, _003766_, _003767_, _003768_, _003769_, _003770_, _003771_, _003772_, _003773_, _003774_, _003775_, _003776_, _003777_, _003778_, _003779_, _003780_, _003781_, _003782_, _003783_, _003784_, _003785_, _003786_, _003787_, _003788_, _003789_, _003790_, _003791_, _003792_, _003793_, _003794_, _003795_, _003796_, _003797_, _003798_, _003799_, _003800_, _003801_, _003802_, _003803_, _003804_, _003805_, _003806_, _003807_, _003808_, _003809_, _003810_, _003811_, _003812_, _003813_, _003814_, _003815_, _003816_, _003817_, _003818_, _003819_, _003820_, _003821_, _003822_, _003823_, _003824_, _003825_, _003826_, _003827_, _003828_, _003829_, _003830_, _003831_, _003832_, _003833_, _003834_, _003835_, _003836_, _003837_, _003838_, _003839_, _003840_, _003841_, _003842_, _003843_, _003844_, _003845_, _003846_, _003847_, _003848_, _003849_, _003850_, _003851_, _003852_, _003853_, _003854_, _003855_, _003856_, _003857_, _003858_, _003859_, _003860_, _003861_, _003862_, _003863_, _003864_, _003865_, _003866_, _003867_, _003868_, _003869_, _003870_, _003871_, _003872_, _003873_, _003874_, _003875_, _003876_, _003877_, _003878_, _003879_, _003880_, _003881_, _003882_, _003883_, _003884_, _003885_, _003886_, _003887_, _003888_, _003889_, _003890_, _003891_, _003892_, _003893_, _003894_, _003895_, _003896_, _003897_, _003898_, _003899_, _003900_, _003901_, _003902_, _003903_, _003904_, _003905_, _003906_, _003907_, _003908_, _003909_, _003910_, _003911_, _003912_, _003913_, _003914_, _003915_, _003916_, _003917_, _003918_, _003919_, _003920_, _003921_, _003922_, _003923_, _003924_, _003925_, _003926_, _003927_, _003928_, _003929_, _003930_, _003931_, _003932_, _003933_, _003934_, _003935_, _003936_, _003937_, _003938_, _003939_, _003940_, _003941_, _003942_, _003943_, _003944_, _003945_, _003946_, _003947_, _003948_, _003949_, _003950_, _003951_, _003952_, _003953_, _003954_, _003955_, _003956_, _003957_, _003958_, _003959_, _003960_, _003961_, _003962_, _003963_, _003964_, _003965_, _003966_, _003967_, _003968_, _003969_, _003970_, _003971_, _003972_, _003973_, _003974_, _003975_, _003976_, _003977_, _003978_, _003979_, _003980_, _003981_, _003982_, _003983_, _003984_, _003985_, _003986_, _003987_, _003988_, _003989_, _003990_, _003991_, _003992_, _003993_, _003994_, _003995_, _003996_, _003997_, _003998_, _003999_, _004000_, _004001_, _004002_, _004003_, _004004_, _004005_, _004006_, _004007_, _004008_, _004009_, _004010_, _004011_, _004012_, _004013_, _004014_, _004015_, _004016_, _004017_, _004018_, _004019_, _004020_, _004021_, _004022_, _004023_, _004024_, _004025_, _004026_, _004027_, _004028_, _004029_, _004030_, _004031_, _004032_, _004033_, _004034_, _004035_, _004036_, _004037_, _004038_, _004039_, _004040_, _004041_, _004042_, _004043_, _004044_, _004045_, _004046_, _004047_, _004048_, _004049_, _004050_, _004051_, _004052_, _004053_, _004054_, _004055_, _004056_, _004057_, _004058_, _004059_, _004060_, _004061_, _004062_, _004063_, _004064_, _004065_, _004066_, _004067_, _004068_, _004069_, _004070_, _004071_, _004072_, _004073_, _004074_, _004075_, _004076_, _004077_, _004078_, _004079_, _004080_, _004081_, _004082_, _004083_, _004084_, _004085_, _004086_, _004087_, _004088_, _004089_, _004090_, _004091_, _004092_, _004093_, _004094_, _004095_, _004096_, _004097_, _004098_, _004099_, _004100_, _004101_, _004102_, _004103_, _004104_, _004105_, _004106_, _004107_, _004108_, _004109_, _004110_, _004111_, _004112_, _004113_, _004114_, _004115_, _004116_, _004117_, _004118_, _004119_, _004120_, _004121_, _004122_, _004123_, _004124_, _004125_, _004126_, _004127_, _004128_, _004129_, _004130_, _004131_, _004132_, _004133_, _004134_, _004135_, _004136_, _004137_, _004138_, _004139_, _004140_, _004141_, _004142_, _004143_, _004144_, _004145_, _004146_, _004147_, _004148_, _004149_, _004150_, _004151_, _004152_, _004153_, _004154_, _004155_, _004156_, _004157_, _004158_, _004159_, _004160_, _004161_, _004162_, _004163_, _004164_, _004165_, _004166_, _004167_, _004168_, _004169_, _004170_, _004171_, _004172_, _004173_, _004174_, _004175_, _004176_, _004177_, _004178_, _004179_, _004180_, _004181_, _004182_, _004183_, _004184_, _004185_, _004186_, _004187_, _004188_, _004189_, _004190_, _004191_, _004192_, _004193_, _004194_, _004195_, _004196_, _004197_, _004198_, _004199_, _004200_, _004201_, _004202_, _004203_, _004204_, _004205_, _004206_, _004207_, _004208_, _004209_, _004210_, _004211_, _004212_, _004213_, _004214_, _004215_, _004216_, _004217_, _004218_, _004219_, _004220_, _004221_, _004222_, _004223_, _004224_, _004225_, _004226_, _004227_, _004228_, _004229_, _004230_, _004231_, _004232_, _004233_, _004234_, _004235_, _004236_, _004237_, _004238_, _004239_, _004240_, _004241_, _004242_, _004243_, _004244_, _004245_, _004246_, _004247_, _004248_, _004249_, _004250_, _004251_, _004252_, _004253_, _004254_, _004255_, _004256_, _004257_, _004258_, _004259_, _004260_, _004261_, _004262_, _004263_, _004264_, _004265_, _004266_, _004267_, _004268_, _004269_, _004270_, _004271_, _004272_, _004273_, _004274_, _004275_, _004276_, _004277_, _004278_, _004279_, _004280_, _004281_, _004282_, _004283_, _004284_, _004285_, _004286_, _004287_, _004288_, _004289_, _004290_, _004291_, _004292_, _004293_, _004294_, _004295_, _004296_, _004297_, _004298_, _004299_, _004300_, _004301_, _004302_, _004303_, _004304_, _004305_, _004306_, _004307_, _004308_, _004309_, _004310_, _004311_, _004312_, _004313_, _004314_, _004315_, _004316_, _004317_, _004318_, _004319_, _004320_, _004321_, _004322_, _004323_, _004324_, _004325_, _004326_, _004327_, _004328_, _004329_, _004330_, _004331_, _004332_, _004333_, _004334_, _004335_, _004336_, _004337_, _004338_, _004339_, _004340_, _004341_, _004342_, _004343_, _004344_, _004345_, _004346_, _004347_, _004348_, _004349_, _004350_, _004351_, _004352_, _004353_, _004354_, _004355_, _004356_, _004357_, _004358_, _004359_, _004360_, _004361_, _004362_, _004363_, _004364_, _004365_, _004366_, _004367_, _004368_, _004369_, _004370_, _004371_, _004372_, _004373_, _004374_, _004375_, _004376_, _004377_, _004378_, _004379_, _004380_, _004381_, _004382_, _004383_, _004384_, _004385_, _004386_, _004387_, _004388_, _004389_, _004390_, _004391_, _004392_, _004393_, _004394_, _004395_, _004396_, _004397_, _004398_, _004399_, _004400_, _004401_, _004402_, _004403_, _004404_, _004405_, _004406_, _004407_, _004408_, _004409_, _004410_, _004411_, _004412_, _004413_, _004414_, _004415_, _004416_, _004417_, _004418_, _004419_, _004420_, _004421_, _004422_, _004423_, _004424_, _004425_, _004426_, _004427_, _004428_, _004429_, _004430_, _004431_, _004432_, _004433_, _004434_, _004435_, _004436_, _004437_, _004438_, _004439_, _004440_, _004441_, _004442_, _004443_, _004444_, _004445_, _004446_, _004447_, _004448_, _004449_, _004450_, _004451_, _004452_, _004453_, _004454_, _004455_, _004456_, _004457_, _004458_, _004459_, _004460_, _004461_, _004462_, _004463_, _004464_, _004465_, _004466_, _004467_, _004468_, _004469_, _004470_, _004471_, _004472_, _004473_, _004474_, _004475_, _004476_, _004477_, _004478_, _004479_, _004480_, _004481_, _004482_, _004483_, _004484_, _004485_, _004486_, _004487_, _004488_, _004489_, _004490_, _004491_, _004492_, _004493_, _004494_, _004495_, _004496_, _004497_, _004498_, _004499_, _004500_, _004501_, _004502_, _004503_, _004504_, _004505_, _004506_, _004507_, _004508_, _004509_, _004510_, _004511_, _004512_, _004513_, _004514_, _004515_, _004516_, _004517_, _004518_, _004519_, _004520_, _004521_, _004522_, _004523_, _004524_, _004525_, _004526_, _004527_, _004528_, _004529_, _004530_, _004531_, _004532_, _004533_, _004534_, _004535_, _004536_, _004537_, _004538_, _004539_, _004540_, _004541_, _004542_, _004543_, _004544_, _004545_, _004546_, _004547_, _004548_, _004549_, _004550_, _004551_, _004552_, _004553_, _004554_, _004555_, _004556_, _004557_, _004558_, _004559_, _004560_, _004561_, _004562_, _004563_, _004564_, _004565_, _004566_, _004567_, _004568_, _004569_, _004570_, _004571_, _004572_, _004573_, _004574_, _004575_, _004576_, _004577_, _004578_, _004579_, _004580_, _004581_, _004582_, _004583_, _004584_, _004585_, _004586_, _004587_, _004588_, _004589_, _004590_, _004591_, _004592_, _004593_, _004594_, _004595_, _004596_, _004597_, _004598_, _004599_, _004600_, _004601_, _004602_, _004603_, _004604_, _004605_, _004606_, _004607_, _004608_, _004609_, _004610_, _004611_, _004612_, _004613_, _004614_, _004615_, _004616_, _004617_, _004618_, _004619_, _004620_, _004621_, _004622_, _004623_, _004624_, _004625_, _004626_, _004627_, _004628_, _004629_, _004630_, _004631_, _004632_, _004633_, _004634_, _004635_, _004636_, _004637_, _004638_, _004639_, _004640_, _004641_, _004642_, _004643_, _004644_, _004645_, _004646_, _004647_, _004648_, _004649_, _004650_, _004651_, _004652_, _004653_, _004654_, _004655_, _004656_, _004657_, _004658_, _004659_, _004660_, _004661_, _004662_, _004663_, _004664_, _004665_, _004666_, _004667_, _004668_, _004669_, _004670_, _004671_, _004672_, _004673_, _004674_, _004675_, _004676_, _004677_, _004678_, _004679_, _004680_, _004681_, _004682_, _004683_, _004684_, _004685_, _004686_, _004687_, _004688_, _004689_, _004690_, _004691_, _004692_, _004693_, _004694_, _004695_, _004696_, _004697_, _004698_, _004699_, _004700_, _004701_, _004702_, _004703_, _004704_, _004705_, _004706_, _004707_, _004708_, _004709_, _004710_, _004711_, _004712_, _004713_, _004714_, _004715_, _004716_, _004717_, _004718_, _004719_, _004720_, _004721_, _004722_, _004723_, _004724_, _004725_, _004726_, _004727_, _004728_, _004729_, _004730_, _004731_, _004732_, _004733_, _004734_, _004735_, _004736_, _004737_, _004738_, _004739_, _004740_, _004741_, _004742_, _004743_, _004744_, _004745_, _004746_, _004747_, _004748_, _004749_, _004750_, _004751_, _004752_, _004753_, _004754_, _004755_, _004756_, _004757_, _004758_, _004759_, _004760_, _004761_, _004762_, _004763_, _004764_, _004765_, _004766_, _004767_, _004768_, _004769_, _004770_, _004771_, _004772_, _004773_, _004774_, _004775_, _004776_, _004777_, _004778_, _004779_, _004780_, _004781_, _004782_, _004783_, _004784_, _004785_, _004786_, _004787_, _004788_, _004789_, _004790_, _004791_, _004792_, _004793_, _004794_, _004795_, _004796_, _004797_, _004798_, _004799_, _004800_, _004801_, _004802_, _004803_, _004804_, _004805_, _004806_, _004807_, _004808_, _004809_, _004810_, _004811_, _004812_, _004813_, _004814_, _004815_, _004816_, _004817_, _004818_, _004819_, _004820_, _004821_, _004822_, _004823_, _004824_, _004825_, _004826_, _004827_, _004828_, _004829_, _004830_, _004831_, _004832_, _004833_, _004834_, _004835_, _004836_, _004837_, _004838_, _004839_, _004840_, _004841_, _004842_, _004843_, _004844_, _004845_, _004846_, _004847_, _004848_, _004849_, _004850_, _004851_, _004852_, _004853_, _004854_, _004855_, _004856_, _004857_, _004858_, _004859_, _004860_, _004861_, _004862_, _004863_, _004864_, _004865_, _004866_, _004867_, _004868_, _004869_, _004870_, _004871_, _004872_, _004873_, _004874_, _004875_, _004876_, _004877_, _004878_, _004879_, _004880_, _004881_, _004882_, _004883_, _004884_, _004885_, _004886_, _004887_, _004888_, _004889_, _004890_, _004891_, _004892_, _004893_, _004894_, _004895_, _004896_, _004897_, _004898_, _004899_, _004900_, _004901_, _004902_, _004903_, _004904_, _004905_, _004906_, _004907_, _004908_, _004909_, _004910_, _004911_, _004912_, _004913_, _004914_, _004915_, _004916_, _004917_, _004918_, _004919_, _004920_, _004921_, _004922_, _004923_, _004924_, _004925_, _004926_, _004927_, _004928_, _004929_, _004930_, _004931_, _004932_, _004933_, _004934_, _004935_, _004936_, _004937_, _004938_, _004939_, _004940_, _004941_, _004942_, _004943_, _004944_, _004945_, _004946_, _004947_, _004948_, _004949_, _004950_, _004951_, _004952_, _004953_, _004954_, _004955_, _004956_, _004957_, _004958_, _004959_, _004960_, _004961_, _004962_, _004963_, _004964_, _004965_, _004966_, _004967_, _004968_, _004969_, _004970_, _004971_, _004972_, _004973_, _004974_, _004975_, _004976_, _004977_, _004978_, _004979_, _004980_, _004981_, _004982_, _004983_, _004984_, _004985_, _004986_, _004987_, _004988_, _004989_, _004990_, _004991_, _004992_, _004993_, _004994_, _004995_, _004996_, _004997_, _004998_, _004999_, _005000_, _005001_, _005002_, _005003_, _005004_, _005005_, _005006_, _005007_, _005008_, _005009_, _005010_, _005011_, _005012_, _005013_, _005014_, _005015_, _005016_, _005017_, _005018_, _005019_, _005020_, _005021_, _005022_, _005023_, _005024_, _005025_, _005026_, _005027_, _005028_, _005029_, _005030_, _005031_, _005032_, _005033_, _005034_, _005035_, _005036_, _005037_, _005038_, _005039_, _005040_, _005041_, _005042_, _005043_, _005044_, _005045_, _005046_, _005047_, _005048_, _005049_, _005050_, _005051_, _005052_, _005053_, _005054_, _005055_, _005056_, _005057_, _005058_, _005059_, _005060_, _005061_, _005062_, _005063_, _005064_, _005065_, _005066_, _005067_, _005068_, _005069_, _005070_, _005071_, _005072_, _005073_, _005074_, _005075_, _005076_, _005077_, _005078_, _005079_, _005080_, _005081_, _005082_, _005083_, _005084_, _005085_, _005086_, _005087_, _005088_, _005089_, _005090_, _005091_, _005092_, _005093_, _005094_, _005095_, _005096_, _005097_, _005098_, _005099_, _005100_, _005101_, _005102_, _005103_, _005104_, _005105_, _005106_, _005107_, _005108_, _005109_, _005110_, _005111_, _005112_, _005113_, _005114_, _005115_, _005116_, _005117_, _005118_, _005119_, _005120_, _005121_, _005122_, _005123_, _005124_, _005125_, _005126_, _005127_, _005128_, _005129_, _005130_, _005131_, _005132_, _005133_, _005134_, _005135_, _005136_, _005137_, _005138_, _005139_, _005140_, _005141_, _005142_, _005143_, _005144_, _005145_, _005146_, _005147_, _005148_, _005149_, _005150_, _005151_, _005152_, _005153_, _005154_, _005155_, _005156_, _005157_, _005158_, _005159_, _005160_, _005161_, _005162_, _005163_, _005164_, _005165_, _005166_, _005167_, _005168_, _005169_, _005170_, _005171_, _005172_, _005173_, _005174_, _005175_, _005176_, _005177_, _005178_, _005179_, _005180_, _005181_, _005182_, _005183_, _005184_, _005185_, _005186_, _005187_, _005188_, _005189_, _005190_, _005191_, _005192_, _005193_, _005194_, _005195_, _005196_, _005197_, _005198_, _005199_, _005200_, _005201_, _005202_, _005203_, _005204_, _005205_, _005206_, _005207_, _005208_, _005209_, _005210_, _005211_, _005212_, _005213_, _005214_, _005215_, _005216_, _005217_, _005218_, _005219_, _005220_, _005221_, _005222_, _005223_, _005224_, _005225_, _005226_, _005227_, _005228_, _005229_, _005230_, _005231_, _005232_, _005233_, _005234_, _005235_, _005236_, _005237_, _005238_, _005239_, _005240_, _005241_, _005242_, _005243_, _005244_, _005245_, _005246_, _005247_, _005248_, _005249_, _005250_, _005251_, _005252_, _005253_, _005254_, _005255_, _005256_, _005257_, _005258_, _005259_, _005260_, _005261_, _005262_, _005263_, _005264_, _005265_, _005266_, _005267_, _005268_, _005269_, _005270_, _005271_, _005272_, _005273_, _005274_, _005275_, _005276_, _005277_, _005278_, _005279_, _005280_, _005281_, _005282_, _005283_, _005284_, _005285_, _005286_, _005287_, _005288_, _005289_, _005290_, _005291_, _005292_, _005293_, _005294_, _005295_, _005296_, _005297_, _005298_, _005299_, _005300_, _005301_, _005302_, _005303_, _005304_, _005305_, _005306_, _005307_, _005308_, _005309_, _005310_, _005311_, _005312_, _005313_, _005314_, _005315_, _005316_, _005317_, _005318_, _005319_, _005320_, _005321_, _005322_, _005323_, _005324_, _005325_, _005326_, _005327_, _005328_, _005329_, _005330_, _005331_, _005332_, _005333_, _005334_, _005335_, _005336_, _005337_, _005338_, _005339_, _005340_, _005341_, _005342_, _005343_, _005344_, _005345_, _005346_, _005347_, _005348_, _005349_, _005350_, _005351_, _005352_, _005353_, _005354_, _005355_, _005356_, _005357_, _005358_, _005359_, _005360_, _005361_, _005362_, _005363_, _005364_, _005365_, _005366_, _005367_, _005368_, _005369_, _005370_, _005371_, _005372_, _005373_, _005374_, _005375_, _005376_, _005377_, _005378_, _005379_, _005380_, _005381_, _005382_, _005383_, _005384_, _005385_, _005386_, _005387_, _005388_, _005389_, _005390_, _005391_, _005392_, _005393_, _005394_, _005395_, _005396_, _005397_, _005398_, _005399_, _005400_, _005401_, _005402_, _005403_, _005404_, _005405_, _005406_, _005407_, _005408_, _005409_, _005410_, _005411_, _005412_, _005413_, _005414_, _005415_, _005416_, _005417_, _005418_, _005419_, _005420_, _005421_, _005422_, _005423_, _005424_, _005425_, _005426_, _005427_, _005428_, _005429_, _005430_, _005431_, _005432_, _005433_, _005434_, _005435_, _005436_, _005437_, _005438_, _005439_, _005440_, _005441_, _005442_, _005443_, _005444_, _005445_, _005446_, _005447_, _005448_, _005449_, _005450_, _005451_, _005452_, _005453_, _005454_, _005455_, _005456_, _005457_, _005458_, _005459_, _005460_, _005461_, _005462_, _005463_, _005464_, _005465_, _005466_, _005467_, _005468_, _005469_, _005470_, _005471_, _005472_, _005473_, _005474_, _005475_, _005476_, _005477_, _005478_, _005479_, _005480_, _005481_, _005482_, _005483_, _005484_, _005485_, _005486_, _005487_, _005488_, _005489_, _005490_, _005491_, _005492_, _005493_, _005494_, _005495_, _005496_, _005497_, _005498_, _005499_, _005500_, _005501_, _005502_, _005503_, _005504_, _005505_, _005506_, _005507_, _005508_, _005509_, _005510_, _005511_, _005512_, _005513_, _005514_, _005515_, _005516_, _005517_, _005518_, _005519_, _005520_, _005521_, _005522_, _005523_, _005524_, _005525_, _005526_, _005527_, _005528_, _005529_, _005530_, _005531_, _005532_, _005533_, _005534_, _005535_, _005536_, _005537_, _005538_, _005539_, _005540_, _005541_, _005542_, _005543_, _005544_, _005545_, _005546_, _005547_, _005548_, _005549_, _005550_, _005551_, _005552_, _005553_, _005554_, _005555_, _005556_, _005557_, _005558_, _005559_, _005560_, _005561_, _005562_, _005563_, _005564_, _005565_, _005566_, _005567_, _005568_, _005569_, _005570_, _005571_, _005572_, _005573_, _005574_, _005575_, _005576_, _005577_, _005578_, _005579_, _005580_, _005581_, _005582_, _005583_, _005584_, _005585_, _005586_, _005587_, _005588_, _005589_, _005590_, _005591_, _005592_, _005593_, _005594_, _005595_, _005596_, _005597_, _005598_, _005599_, _005600_, _005601_, _005602_, _005603_, _005604_, _005605_, _005606_, _005607_, _005608_, _005609_, _005610_, _005611_, _005612_, _005613_, _005614_, _005615_, _005616_, _005617_, _005618_, _005619_, _005620_, _005621_, _005622_, _005623_, _005624_, _005625_, _005626_, _005627_, _005628_, _005629_, _005630_, _005631_, _005632_, _005633_, _005634_, _005635_, _005636_, _005637_, _005638_, _005639_, _005640_, _005641_, _005642_, _005643_, _005644_, _005645_, _005646_, _005647_, _005648_, _005649_, _005650_, _005651_, _005652_, _005653_, _005654_, _005655_, _005656_, _005657_, _005658_, _005659_, _005660_, _005661_, _005662_, _005663_, _005664_, _005665_, _005666_, _005667_, _005668_, _005669_, _005670_, _005671_, _005672_, _005673_, _005674_, _005675_, _005676_, _005677_, _005678_, _005679_, _005680_, _005681_, _005682_, _005683_, _005684_, _005685_, _005686_, _005687_, _005688_, _005689_, _005690_, _005691_, _005692_, _005693_, _005694_, _005695_, _005696_, _005697_, _005698_, _005699_, _005700_, _005701_, _005702_, _005703_, _005704_, _005705_, _005706_, _005707_, _005708_, _005709_, _005710_, _005711_, _005712_, _005713_, _005714_, _005715_, _005716_, _005717_, _005718_, _005719_, _005720_, _005721_, _005722_, _005723_, _005724_, _005725_, _005726_, _005727_, _005728_, _005729_, _005730_, _005731_, _005732_, _005733_, _005734_, _005735_, _005736_, _005737_, _005738_, _005739_, _005740_, _005741_, _005742_, _005743_, _005744_, _005745_, _005746_, _005747_, _005748_, _005749_, _005750_, _005751_, _005752_, _005753_, _005754_, _005755_, _005756_, _005757_, _005758_, _005759_, _005760_, _005761_, _005762_, _005763_, _005764_, _005765_, _005766_, _005767_, _005768_, _005769_, _005770_, _005771_, _005772_, _005773_, _005774_, _005775_, _005776_, _005777_, _005778_, _005779_, _005780_, _005781_, _005782_, _005783_, _005784_, _005785_, _005786_, _005787_, _005788_, _005789_, _005790_, _005791_, _005792_, _005793_, _005794_, _005795_, _005796_, _005797_, _005798_, _005799_, _005800_, _005801_, _005802_, _005803_, _005804_, _005805_, _005806_, _005807_, _005808_, _005809_, _005810_, _005811_, _005812_, _005813_, _005814_, _005815_, _005816_, _005817_, _005818_, _005819_, _005820_, _005821_, _005822_, _005823_, _005824_, _005825_, _005826_, _005827_, _005828_, _005829_, _005830_, _005831_, _005832_, _005833_, _005834_, _005835_, _005836_, _005837_, _005838_, _005839_, _005840_, _005841_, _005842_, _005843_, _005844_, _005845_, _005846_, _005847_, _005848_, _005849_, _005850_, _005851_, _005852_, _005853_, _005854_, _005855_, _005856_, _005857_, _005858_, _005859_, _005860_, _005861_, _005862_, _005863_, _005864_, _005865_, _005866_, _005867_, _005868_, _005869_, _005870_, _005871_, _005872_, _005873_, _005874_, _005875_, _005876_, _005877_, _005878_, _005879_, _005880_, _005881_, _005882_, _005883_, _005884_, _005885_, _005886_, _005887_, _005888_, _005889_, _005890_, _005891_, _005892_, _005893_, _005894_, _005895_, _005896_, _005897_, _005898_, _005899_, _005900_, _005901_, _005902_, _005903_, _005904_, _005905_, _005906_, _005907_, _005908_, _005909_, _005910_, _005911_, _005912_, _005913_, _005914_, _005915_, _005916_, _005917_, _005918_, _005919_, _005920_, _005921_, _005922_, _005923_, _005924_, _005925_, _005926_, _005927_, _005928_, _005929_, _005930_, _005931_, _005932_, _005933_, _005934_, _005935_, _005936_, _005937_, _005938_, _005939_, _005940_, _005941_, _005942_, _005943_, _005944_, _005945_, _005946_, _005947_, _005948_, _005949_, _005950_, _005951_, _005952_, _005953_, _005954_, _005955_, _005956_, _005957_, _005958_, _005959_, _005960_, _005961_, _005962_, _005963_, _005964_, _005965_, _005966_, _005967_, _005968_, _005969_, _005970_, _005971_, _005972_, _005973_, _005974_, _005975_, _005976_, _005977_, _005978_, _005979_, _005980_, _005981_, _005982_, _005983_, _005984_, _005985_, _005986_, _005987_, _005988_, _005989_, _005990_, _005991_, _005992_, _005993_, _005994_, _005995_, _005996_, _005997_, _005998_, _005999_, _006000_, _006001_, _006002_, _006003_, _006004_, _006005_, _006006_, _006007_, _006008_, _006009_, _006010_, _006011_, _006012_, _006013_, _006014_, _006015_, _006016_, _006017_, _006018_, _006019_, _006020_, _006021_, _006022_, _006023_, _006024_, _006025_, _006026_, _006027_, _006028_, _006029_, _006030_, _006031_, _006032_, _006033_, _006034_, _006035_, _006036_, _006037_, _006038_, _006039_, _006040_, _006041_, _006042_, _006043_, _006044_, _006045_, _006046_, _006047_, _006048_, _006049_, _006050_, _006051_, _006052_, _006053_, _006054_, _006055_, _006056_, _006057_, _006058_, _006059_, _006060_, _006061_, _006062_, _006063_, _006064_, _006065_, _006066_, _006067_, _006068_, _006069_, _006070_, _006071_, _006072_, _006073_, _006074_, _006075_, _006076_, _006077_, _006078_, _006079_, _006080_, _006081_, _006082_, _006083_, _006084_, _006085_, _006086_, _006087_, _006088_, _006089_, _006090_, _006091_, _006092_, _006093_, _006094_, _006095_, _006096_, _006097_, _006098_, _006099_, _006100_, _006101_, _006102_, _006103_, _006104_, _006105_, _006106_, _006107_, _006108_, _006109_, _006110_, _006111_, _006112_, _006113_, _006114_, _006115_, _006116_, _006117_, _006118_, _006119_, _006120_, _006121_, _006122_, _006123_, _006124_, _006125_, _006126_, _006127_, _006128_, _006129_, _006130_, _006131_, _006132_, _006133_, _006134_, _006135_, _006136_, _006137_, _006138_, _006139_, _006140_, _006141_, _006142_, _006143_, _006144_, _006145_, _006146_, _006147_, _006148_, _006149_, _006150_, _006151_, _006152_, _006153_, _006154_, _006155_, _006156_, _006157_, _006158_, _006159_, _006160_, _006161_, _006162_, _006163_, _006164_, _006165_, _006166_, _006167_, _006168_, _006169_, _006170_, _006171_, _006172_, _006173_, _006174_, _006175_, _006176_, _006177_, _006178_, _006179_, _006180_, _006181_, _006182_, _006183_, _006184_, _006185_, _006186_, _006187_, _006188_, _006189_, _006190_, _006191_, _006192_, _006193_, _006194_, _006195_, _006196_, _006197_, _006198_, _006199_, _006200_, _006201_, _006202_, _006203_, _006204_, _006205_, _006206_, _006207_, _006208_, _006209_, _006210_, _006211_, _006212_, _006213_, _006214_, _006215_, _006216_, _006217_, _006218_, _006219_, _006220_, _006221_, _006222_, _006223_, _006224_, _006225_, _006226_, _006227_, _006228_, _006229_, _006230_, _006231_, _006232_, _006233_, _006234_, _006235_, _006236_, _006237_, _006238_, _006239_, _006240_, _006241_, _006242_, _006243_, _006244_, _006245_, _006246_, _006247_, _006248_, _006249_, _006250_, _006251_, _006252_, _006253_, _006254_, _006255_, _006256_, _006257_, _006258_, _006259_, _006260_, _006261_, _006262_, _006263_, _006264_, _006265_, _006266_, _006267_, _006268_, _006269_, _006270_, _006271_, _006272_, _006273_, _006274_, _006275_, _006276_, _006277_, _006278_, _006279_, _006280_, _006281_, _006282_, _006283_, _006284_, _006285_, _006286_, _006287_, _006288_, _006289_, _006290_, _006291_, _006292_, _006293_, _006294_, _006295_, _006296_, _006297_, _006298_, _006299_, _006300_, _006301_, _006302_, _006303_, _006304_, _006305_, _006306_, _006307_, _006308_, _006309_, _006310_, _006311_, _006312_, _006313_, _006314_, _006315_, _006316_, _006317_, _006318_, _006319_, _006320_, _006321_, _006322_, _006323_, _006324_, _006325_, _006326_, _006327_, _006328_, _006329_, _006330_, _006331_, _006332_, _006333_, _006334_, _006335_, _006336_, _006337_, _006338_, _006339_, _006340_, _006341_, _006342_, _006343_, _006344_, _006345_, _006346_, _006347_, _006348_, _006349_, _006350_, _006351_, _006352_, _006353_, _006354_, _006355_, _006356_, _006357_, _006358_, _006359_, _006360_, _006361_, _006362_, _006363_, _006364_, _006365_, _006366_, _006367_, _006368_, _006369_, _006370_, _006371_, _006372_, _006373_, _006374_, _006375_, _006376_, _006377_, _006378_, _006379_, _006380_, _006381_, _006382_, _006383_, _006384_, _006385_, _006386_, _006387_, _006388_, _006389_, _006390_, _006391_, _006392_, _006393_, _006394_, _006395_, _006396_, _006397_, _006398_, _006399_, _006400_, _006401_, _006402_, _006403_, _006404_, _006405_, _006406_, _006407_, _006408_, _006409_, _006410_, _006411_, _006412_, _006413_, _006414_, _006415_, _006416_, _006417_, _006418_, _006419_, _006420_, _006421_, _006422_, _006423_, _006424_, _006425_, _006426_, _006427_, _006428_, _006429_, _006430_, _006431_, _006432_, _006433_, _006434_, _006435_, _006436_, _006437_, _006438_, _006439_, _006440_, _006441_, _006442_, _006443_, _006444_, _006445_, _006446_, _006447_, _006448_, _006449_, _006450_, _006451_, _006452_, _006453_, _006454_, _006455_, _006456_, _006457_, _006458_, _006459_, _006460_, _006461_, _006462_, _006463_, _006464_, _006465_, _006466_, _006467_, _006468_, _006469_, _006470_, _006471_, _006472_, _006473_, _006474_, _006475_, _006476_, _006477_, _006478_, _006479_, _006480_, _006481_, _006482_, _006483_, _006484_, _006485_, _006486_, _006487_, _006488_, _006489_, _006490_, _006491_, _006492_, _006493_, _006494_, _006495_, _006496_, _006497_, _006498_, _006499_, _006500_, _006501_, _006502_, _006503_, _006504_, _006505_, _006506_, _006507_, _006508_, _006509_, _006510_, _006511_, _006512_, _006513_, _006514_, _006515_, _006516_, _006517_, _006518_, _006519_, _006520_, _006521_, _006522_, _006523_, _006524_, _006525_, _006526_, _006527_, _006528_, _006529_, _006530_, _006531_, _006532_, _006533_, _006534_, _006535_, _006536_, _006537_, _006538_, _006539_, _006540_, _006541_, _006542_, _006543_, _006544_, _006545_, _006546_, _006547_, _006548_, _006549_, _006550_, _006551_, _006552_, _006553_, _006554_, _006555_, _006556_, _006557_, _006558_, _006559_, _006560_, _006561_, _006562_, _006563_, _006564_, _006565_, _006566_, _006567_, _006568_, _006569_, _006570_, _006571_, _006572_, _006573_, _006574_, _006575_, _006576_, _006577_, _006578_, _006579_, _006580_, _006581_, _006582_, _006583_, _006584_, _006585_, _006586_, _006587_, _006588_, _006589_, _006590_, _006591_, _006592_, _006593_, _006594_, _006595_, _006596_, _006597_, _006598_, _006599_, _006600_, _006601_, _006602_, _006603_, _006604_, _006605_, _006606_, _006607_, _006608_, _006609_, _006610_, _006611_, _006612_, _006613_, _006614_, _006615_, _006616_, _006617_, _006618_, _006619_, _006620_, _006621_, _006622_, _006623_, _006624_, _006625_, _006626_, _006627_, _006628_, _006629_, _006630_, _006631_, _006632_, _006633_, _006634_, _006635_, _006636_, _006637_, _006638_, _006639_, _006640_, _006641_, _006642_, _006643_, _006644_, _006645_, _006646_, _006647_, _006648_, _006649_, _006650_, _006651_, _006652_, _006653_, _006654_, _006655_, _006656_, _006657_, _006658_, _006659_, _006660_, _006661_, _006662_, _006663_, _006664_, _006665_, _006666_, _006667_, _006668_, _006669_, _006670_, _006671_, _006672_, _006673_, _006674_, _006675_, _006676_, _006677_, _006678_, _006679_, _006680_, _006681_, _006682_, _006683_, _006684_, _006685_, _006686_, _006687_, _006688_, _006689_, _006690_, _006691_, _006692_, _006693_, _006694_, _006695_, _006696_, _006697_, _006698_, _006699_, _006700_, _006701_, _006702_, _006703_, _006704_, _006705_, _006706_, _006707_, _006708_, _006709_, _006710_, _006711_, _006712_, _006713_, _006714_, _006715_, _006716_, _006717_, _006718_, _006719_, _006720_, _006721_, _006722_, _006723_, _006724_, _006725_, _006726_, _006727_, _006728_, _006729_, _006730_, _006731_, _006732_, _006733_, _006734_, _006735_, _006736_, _006737_, _006738_, _006739_, _006740_, _006741_, _006742_, _006743_, _006744_, _006745_, _006746_, _006747_, _006748_, _006749_, _006750_, _006751_, _006752_, _006753_, _006754_, _006755_, _006756_, _006757_, _006758_, _006759_, _006760_, _006761_, _006762_, _006763_, _006764_, _006765_, _006766_, _006767_, _006768_, _006769_, _006770_, _006771_, _006772_, _006773_, _006774_, _006775_, _006776_, _006777_, _006778_, _006779_, _006780_, _006781_, _006782_, _006783_, _006784_, _006785_, _006786_, _006787_, _006788_, _006789_, _006790_, _006791_, _006792_, _006793_, _006794_, _006795_, _006796_, _006797_, _006798_, _006799_, _006800_, _006801_, _006802_, _006803_, _006804_, _006805_, _006806_, _006807_, _006808_, _006809_, _006810_, _006811_, _006812_, _006813_, _006814_, _006815_, _006816_, _006817_, _006818_, _006819_, _006820_, _006821_, _006822_, _006823_, _006824_, _006825_, _006826_, _006827_, _006828_, _006829_, _006830_, _006831_, _006832_, _006833_, _006834_, _006835_, _006836_, _006837_, _006838_, _006839_, _006840_, _006841_, _006842_, _006843_, _006844_, _006845_, _006846_, _006847_, _006848_, _006849_, _006850_, _006851_, _006852_, _006853_, _006854_, _006855_, _006856_, _006857_, _006858_, _006859_, _006860_, _006861_, _006862_, _006863_, _006864_, _006865_, _006866_, _006867_, _006868_, _006869_, _006870_, _006871_, _006872_, _006873_, _006874_, _006875_, _006876_, _006877_, _006878_, _006879_, _006880_, _006881_, _006882_, _006883_, _006884_, _006885_, _006886_, _006887_, _006888_, _006889_, _006890_, _006891_, _006892_, _006893_, _006894_, _006895_, _006896_, _006897_, _006898_, _006899_, _006900_, _006901_, _006902_, _006903_, _006904_, _006905_, _006906_, _006907_, _006908_, _006909_, _006910_, _006911_, _006912_, _006913_, _006914_, _006915_, _006916_, _006917_, _006918_, _006919_, _006920_, _006921_, _006922_, _006923_, _006924_, _006925_, _006926_, _006927_, _006928_, _006929_, _006930_, _006931_, _006932_, _006933_, _006934_, _006935_, _006936_, _006937_, _006938_, _006939_, _006940_, _006941_, _006942_, _006943_, _006944_, _006945_, _006946_, _006947_, _006948_, _006949_, _006950_, _006951_, _006952_, _006953_, _006954_, _006955_, _006956_, _006957_, _006958_, _006959_, _006960_, _006961_, _006962_, _006963_, _006964_, _006965_, _006966_, _006967_, _006968_, _006969_, _006970_, _006971_, _006972_, _006973_, _006974_, _006975_, _006976_, _006977_, _006978_, _006979_, _006980_, _006981_, _006982_, _006983_, _006984_, _006985_, _006986_, _006987_, _006988_, _006989_, _006990_, _006991_, _006992_, _006993_, _006994_, _006995_, _006996_, _006997_, _006998_, _006999_, _007000_, _007001_, _007002_, _007003_, _007004_, _007005_, _007006_, _007007_, _007008_, _007009_, _007010_, _007011_, _007012_, _007013_, _007014_, _007015_, _007016_, _007017_, _007018_, _007019_, _007020_, _007021_, _007022_, _007023_, _007024_, _007025_, _007026_, _007027_, _007028_, _007029_, _007030_, _007031_, _007032_, _007033_, _007034_, _007035_, _007036_, _007037_, _007038_, _007039_, _007040_, _007041_, _007042_, _007043_, _007044_, _007045_, _007046_, _007047_, _007048_, _007049_, _007050_, _007051_, _007052_, _007053_, _007054_, _007055_, _007056_, _007057_, _007058_, _007059_, _007060_, _007061_, _007062_, _007063_, _007064_, _007065_, _007066_, _007067_, _007068_, _007069_, _007070_, _007071_, _007072_, _007073_, _007074_, _007075_, _007076_, _007077_, _007078_, _007079_, _007080_, _007081_, _007082_, _007083_, _007084_, _007085_, _007086_, _007087_, _007088_, _007089_, _007090_, _007091_, _007092_, _007093_, _007094_, _007095_, _007096_, _007097_, _007098_, _007099_, _007100_, _007101_, _007102_, _007103_, _007104_, _007105_, _007106_, _007107_, _007108_, _007109_, _007110_, _007111_, _007112_, _007113_, _007114_, _007115_, _007116_, _007117_, _007118_, _007119_, _007120_, _007121_, _007122_, _007123_, _007124_, _007125_, _007126_, _007127_, _007128_, _007129_, _007130_, _007131_, _007132_, _007133_, _007134_, _007135_, _007136_, _007137_, _007138_, _007139_, _007140_, _007141_, _007142_, _007143_, _007144_, _007145_, _007146_, _007147_, _007148_, _007149_, _007150_, _007151_, _007152_, _007153_, _007154_, _007155_, _007156_, _007157_, _007158_, _007159_, _007160_, _007161_, _007162_, _007163_, _007164_, _007165_, _007166_, _007167_, _007168_, _007169_, _007170_, _007171_, _007172_, _007173_, _007174_, _007175_, _007176_, _007177_, _007178_, _007179_, _007180_, _007181_, _007182_, _007183_, _007184_, _007185_, _007186_, _007187_, _007188_, _007189_, _007190_, _007191_, _007192_, _007193_, _007194_, _007195_, _007196_, _007197_, _007198_, _007199_, _007200_, _007201_, _007202_, _007203_, _007204_, _007205_, _007206_, _007207_, _007208_, _007209_, _007210_, _007211_, _007212_, _007213_, _007214_, _007215_, _007216_, _007217_, _007218_, _007219_, _007220_, _007221_, _007222_, _007223_, _007224_, _007225_, _007226_, _007227_, _007228_, _007229_, _007230_, _007231_, _007232_, _007233_, _007234_, _007235_, _007236_, _007237_, _007238_, _007239_, _007240_, _007241_, _007242_, _007243_, _007244_, _007245_, _007246_, _007247_, _007248_, _007249_, _007250_, _007251_, _007252_, _007253_, _007254_, _007255_, _007256_, _007257_, _007258_, _007259_, _007260_, _007261_, _007262_, _007263_, _007264_, _007265_, _007266_, _007267_, _007268_, _007269_, _007270_, _007271_, _007272_, _007273_, _007274_, _007275_, _007276_, _007277_, _007278_, _007279_, _007280_, _007281_, _007282_, _007283_, _007284_, _007285_, _007286_, _007287_, _007288_, _007289_, _007290_, _007291_, _007292_, _007293_, _007294_, _007295_, _007296_, _007297_, _007298_, _007299_, _007300_, _007301_, _007302_, _007303_, _007304_, _007305_, _007306_, _007307_, _007308_, _007309_, _007310_, _007311_, _007312_, _007313_, _007314_, _007315_, _007316_, _007317_, _007318_, _007319_, _007320_, _007321_, _007322_, _007323_, _007324_, _007325_, _007326_, _007327_, _007328_, _007329_, _007330_, _007331_, _007332_, _007333_, _007334_, _007335_, _007336_, _007337_, _007338_, _007339_, _007340_, _007341_, _007342_, _007343_, _007344_, _007345_, _007346_, _007347_, _007348_, _007349_, _007350_, _007351_, _007352_, _007353_, _007354_, _007355_, _007356_, _007357_, _007358_, _007359_, _007360_, _007361_, _007362_, _007363_, _007364_, _007365_, _007366_, _007367_, _007368_, _007369_, _007370_, _007371_, _007372_, _007373_, _007374_, _007375_, _007376_, _007377_, _007378_, _007379_, _007380_, _007381_, _007382_, _007383_, _007384_, _007385_, _007386_, _007387_, _007388_, _007389_, _007390_, _007391_, _007392_, _007393_, _007394_, _007395_, _007396_, _007397_, _007398_, _007399_, _007400_, _007401_, _007402_, _007403_, _007404_, _007405_, _007406_, _007407_, _007408_, _007409_, _007410_, _007411_, _007412_, _007413_, _007414_, _007415_, _007416_, _007417_, _007418_, _007419_, _007420_, _007421_, _007422_, _007423_, _007424_, _007425_, _007426_, _007427_, _007428_, _007429_, _007430_, _007431_, _007432_, _007433_, _007434_, _007435_, _007436_, _007437_, _007438_, _007439_, _007440_, _007441_, _007442_, _007443_, _007444_, _007445_, _007446_, _007447_, _007448_, _007449_, _007450_, _007451_, _007452_, _007453_, _007454_, _007455_, _007456_, _007457_, _007458_, _007459_, _007460_, _007461_, _007462_, _007463_, _007464_, _007465_, _007466_, _007467_, _007468_, _007469_, _007470_, _007471_, _007472_, _007473_, _007474_, _007475_, _007476_, _007477_, _007478_, _007479_, _007480_, _007481_, _007482_, _007483_, _007484_, _007485_, _007486_, _007487_, _007488_, _007489_, _007490_, _007491_, _007492_, _007493_, _007494_, _007495_, _007496_, _007497_, _007498_, _007499_, _007500_, _007501_, _007502_, _007503_, _007504_, _007505_, _007506_, _007507_, _007508_, _007509_, _007510_, _007511_, _007512_, _007513_, _007514_, _007515_, _007516_, _007517_, _007518_, _007519_, _007520_, _007521_, _007522_, _007523_, _007524_, _007525_, _007526_, _007527_, _007528_, _007529_, _007530_, _007531_, _007532_, _007533_, _007534_, _007535_, _007536_, _007537_, _007538_, _007539_, _007540_, _007541_, _007542_, _007543_, _007544_, _007545_, _007546_, _007547_, _007548_, _007549_, _007550_, _007551_, _007552_, _007553_, _007554_, _007555_, _007556_, _007557_, _007558_, _007559_, _007560_, _007561_, _007562_, _007563_, _007564_, _007565_, _007566_, _007567_, _007568_, _007569_, _007570_, _007571_, _007572_, _007573_, _007574_, _007575_, _007576_, _007577_, _007578_, _007579_, _007580_, _007581_, _007582_, _007583_, _007584_, _007585_, _007586_, _007587_, _007588_, _007589_, _007590_, _007591_, _007592_, _007593_, _007594_, _007595_, _007596_, _007597_, _007598_, _007599_, _007600_, _007601_, _007602_, _007603_, _007604_, _007605_, _007606_, _007607_, _007608_, _007609_, _007610_, _007611_, _007612_, _007613_, _007614_, _007615_, _007616_, _007617_, _007618_, _007619_, _007620_, _007621_, _007622_, _007623_, _007624_, _007625_, _007626_, _007627_, _007628_, _007629_, _007630_, _007631_, _007632_, _007633_, _007634_, _007635_, _007636_, _007637_, _007638_, _007639_, _007640_, _007641_, _007642_, _007643_, _007644_, _007645_, _007646_, _007647_, _007648_, _007649_, _007650_, _007651_, _007652_, _007653_, _007654_, _007655_, _007656_, _007657_, _007658_, _007659_, _007660_, _007661_, _007662_, _007663_, _007664_, _007665_, _007666_, _007667_, _007668_, _007669_, _007670_, _007671_, _007672_, _007673_, _007674_, _007675_, _007676_, _007677_, _007678_, _007679_, _007680_, _007681_, _007682_, _007683_, _007684_, _007685_, _007686_, _007687_, _007688_, _007689_, _007690_, _007691_, _007692_, _007693_, _007694_, _007695_, _007696_, _007697_, _007698_, _007699_, _007700_, _007701_, _007702_, _007703_, _007704_, _007705_, _007706_, _007707_, _007708_, _007709_, _007710_, _007711_, _007712_, _007713_, _007714_, _007715_, _007716_, _007717_, _007718_, _007719_, _007720_, _007721_, _007722_, _007723_, _007724_, _007725_, _007726_, _007727_, _007728_, _007729_, _007730_, _007731_, _007732_, _007733_, _007734_, _007735_, _007736_, _007737_, _007738_, _007739_, _007740_, _007741_, _007742_, _007743_, _007744_, _007745_, _007746_, _007747_, _007748_, _007749_, _007750_, _007751_, _007752_, _007753_, _007754_, _007755_, _007756_, _007757_, _007758_, _007759_, _007760_, _007761_, _007762_, _007763_, _007764_, _007765_, _007766_, _007767_, _007768_, _007769_, _007770_, _007771_, _007772_, _007773_, _007774_, _007775_, _007776_, _007777_, _007778_, _007779_, _007780_, _007781_, _007782_, _007783_, _007784_, _007785_, _007786_, _007787_, _007788_, _007789_, _007790_, _007791_, _007792_, _007793_, _007794_, _007795_, _007796_, _007797_, _007798_, _007799_, _007800_, _007801_, _007802_, _007803_, _007804_, _007805_, _007806_, _007807_, _007808_, _007809_, _007810_, _007811_, _007812_, _007813_, _007814_, _007815_, _007816_, _007817_, _007818_, _007819_, _007820_, _007821_, _007822_, _007823_, _007824_, _007825_, _007826_, _007827_, _007828_, _007829_, _007830_, _007831_, _007832_, _007833_, _007834_, _007835_, _007836_, _007837_, _007838_, _007839_, _007840_, _007841_, _007842_, _007843_, _007844_, _007845_, _007846_, _007847_, _007848_, _007849_, _007850_, _007851_, _007852_, _007853_, _007854_, _007855_, _007856_, _007857_, _007858_, _007859_, _007860_, _007861_, _007862_, _007863_, _007864_, _007865_, _007866_, _007867_, _007868_, _007869_, _007870_, _007871_, _007872_, _007873_, _007874_, _007875_, _007876_, _007877_, _007878_, _007879_, _007880_, _007881_, _007882_, _007883_, _007884_, _007885_, _007886_, _007887_, _007888_, _007889_, _007890_, _007891_, _007892_, _007893_, _007894_, _007895_, _007896_, _007897_, _007898_, _007899_, _007900_, _007901_, _007902_, _007903_, _007904_, _007905_, _007906_, _007907_, _007908_, _007909_, _007910_, _007911_, _007912_, _007913_, _007914_, _007915_, _007916_, _007917_, _007918_, _007919_, _007920_, _007921_, _007922_, _007923_, _007924_, _007925_, _007926_, _007927_, _007928_, _007929_, _007930_, _007931_, _007932_, _007933_, _007934_, _007935_, _007936_, _007937_, _007938_, _007939_, _007940_, _007941_, _007942_, _007943_, _007944_, _007945_, _007946_, _007947_, _007948_, _007949_, _007950_, _007951_, _007952_, _007953_, _007954_, _007955_, _007956_, _007957_, _007958_, _007959_, _007960_, _007961_, _007962_, _007963_, _007964_, _007965_, _007966_, _007967_, _007968_, _007969_, _007970_, _007971_, _007972_, _007973_, _007974_, _007975_, _007976_, _007977_, _007978_, _007979_, _007980_, _007981_, _007982_, _007983_, _007984_, _007985_, _007986_, _007987_, _007988_, _007989_, _007990_, _007991_, _007992_, _007993_, _007994_, _007995_, _007996_, _007997_, _007998_, _007999_, _008000_, _008001_, _008002_, _008003_, _008004_, _008005_, _008006_, _008007_, _008008_, _008009_, _008010_, _008011_, _008012_, _008013_, _008014_, _008015_, _008016_, _008017_, _008018_, _008019_, _008020_, _008021_, _008022_, _008023_, _008024_, _008025_, _008026_, _008027_, _008028_, _008029_, _008030_, _008031_, _008032_, _008033_, _008034_, _008035_, _008036_, _008037_, _008038_, _008039_, _008040_, _008041_, _008042_, _008043_, _008044_, _008045_, _008046_, _008047_, _008048_, _008049_, _008050_, _008051_, _008052_, _008053_, _008054_, _008055_, _008056_, _008057_, _008058_, _008059_, _008060_, _008061_, _008062_, _008063_, _008064_, _008065_, _008066_, _008067_, _008068_, _008069_, _008070_, _008071_, _008072_, _008073_, _008074_, _008075_, _008076_, _008077_, _008078_, _008079_, _008080_, _008081_, _008082_, _008083_, _008084_, _008085_, _008086_, _008087_, _008088_, _008089_, _008090_, _008091_, _008092_, _008093_, _008094_, _008095_, _008096_, _008097_, _008098_, _008099_, _008100_, _008101_, _008102_, _008103_, _008104_, _008105_, _008106_, _008107_, _008108_, _008109_, _008110_, _008111_, _008112_, _008113_, _008114_, _008115_, _008116_, _008117_, _008118_, _008119_, _008120_, _008121_, _008122_, _008123_, _008124_, _008125_, _008126_, _008127_, _008128_, _008129_, _008130_, _008131_, _008132_, _008133_, _008134_, _008135_, _008136_, _008137_, _008138_, _008139_, _008140_, _008141_, _008142_, _008143_, _008144_, _008145_, _008146_, _008147_, _008148_, _008149_, _008150_, _008151_, _008152_, _008153_, _008154_, _008155_, _008156_, _008157_, _008158_, _008159_, _008160_, _008161_, _008162_, _008163_, _008164_, _008165_, _008166_, _008167_, _008168_, _008169_, _008170_, _008171_, _008172_, _008173_, _008174_, _008175_, _008176_, _008177_, _008178_, _008179_, _008180_, _008181_, _008182_, _008183_, _008184_, _008185_, _008186_, _008187_, _008188_, _008189_, _008190_, _008191_, _008192_, _008193_, _008194_, _008195_, _008196_, _008197_, _008198_, _008199_, _008200_, _008201_, _008202_, _008203_, _008204_, _008205_, _008206_, _008207_, _008208_, _008209_, _008210_, _008211_, _008212_, _008213_, _008214_, _008215_, _008216_, _008217_, _008218_, _008219_, _008220_, _008221_, _008222_, _008223_, _008224_, _008225_, _008226_, _008227_, _008228_, _008229_, _008230_, _008231_, _008232_, _008233_, _008234_, _008235_, _008236_, _008237_, _008238_, _008239_, _008240_, _008241_, _008242_, _008243_, _008244_, _008245_, _008246_, _008247_, _008248_, _008249_, _008250_, _008251_, _008252_, _008253_, _008254_, _008255_, _008256_, _008257_, _008258_, _008259_, _008260_, _008261_, _008262_, _008263_, _008264_, _008265_, _008266_, _008267_, _008268_, _008269_, _008270_, _008271_, _008272_, _008273_, _008274_, _008275_, _008276_, _008277_, _008278_, _008279_, _008280_, _008281_, _008282_, _008283_, _008284_, _008285_, _008286_, _008287_, _008288_, _008289_, _008290_, _008291_, _008292_, _008293_, _008294_, _008295_, _008296_, _008297_, _008298_, _008299_, _008300_, _008301_, _008302_, _008303_, _008304_, _008305_, _008306_, _008307_, _008308_, _008309_, _008310_, _008311_, _008312_, _008313_, _008314_, _008315_, _008316_, _008317_, _008318_, _008319_, _008320_, _008321_, _008322_, _008323_, _008324_, _008325_, _008326_, _008327_, _008328_, _008329_, _008330_, _008331_, _008332_, _008333_, _008334_, _008335_, _008336_, _008337_, _008338_, _008339_, _008340_, _008341_, _008342_, _008343_, _008344_, _008345_, _008346_, _008347_, _008348_, _008349_, _008350_, _008351_, _008352_, _008353_, _008354_, _008355_, _008356_, _008357_, _008358_, _008359_, _008360_, _008361_, _008362_, _008363_, _008364_, _008365_, _008366_, _008367_, _008368_, _008369_, _008370_, _008371_, _008372_, _008373_, _008374_, _008375_, _008376_, _008377_, _008378_, _008379_, _008380_, _008381_, _008382_, _008383_, _008384_, _008385_, _008386_, _008387_, _008388_, _008389_, _008390_, _008391_, _008392_, _008393_, _008394_, _008395_, _008396_, _008397_, _008398_, _008399_, _008400_, _008401_, _008402_, _008403_, _008404_, _008405_, _008406_, _008407_, _008408_, _008409_, _008410_, _008411_, _008412_, _008413_, _008414_, _008415_, _008416_, _008417_, _008418_, _008419_, _008420_, _008421_, _008422_, _008423_, _008424_, _008425_, _008426_, _008427_, _008428_, _008429_, _008430_, _008431_, _008432_, _008433_, _008434_, _008435_, _008436_, _008437_, _008438_, _008439_, _008440_, _008441_, _008442_, _008443_, _008444_, _008445_, _008446_, _008447_, _008448_, _008449_, _008450_, _008451_, _008452_, _008453_, _008454_, _008455_, _008456_, _008457_, _008458_, _008459_, _008460_, _008461_, _008462_, _008463_, _008464_, _008465_, _008466_, _008467_, _008468_, _008469_, _008470_, _008471_, _008472_, _008473_, _008474_, _008475_, _008476_, _008477_, _008478_, _008479_, _008480_, _008481_, _008482_, _008483_, _008484_, _008485_, _008486_, _008487_, _008488_, _008489_, _008490_, _008491_, _008492_, _008493_, _008494_, _008495_, _008496_, _008497_, _008498_, _008499_, _008500_, _008501_, _008502_, _008503_, _008504_, _008505_, _008506_, _008507_, _008508_, _008509_, _008510_, _008511_, _008512_, _008513_, _008514_, _008515_, _008516_, _008517_, _008518_, _008519_, _008520_, _008521_, _008522_, _008523_, _008524_, _008525_, _008526_, _008527_, _008528_, _008529_, _008530_, _008531_, _008532_, _008533_, _008534_, _008535_, _008536_, _008537_, _008538_, _008539_, _008540_, _008541_, _008542_, _008543_, _008544_, _008545_, _008546_, _008547_, _008548_, _008549_, _008550_, _008551_, _008552_, _008553_, _008554_, _008555_, _008556_, _008557_, _008558_, _008559_, _008560_, _008561_, _008562_, _008563_, _008564_, _008565_, _008566_, _008567_, _008568_, _008569_, _008570_, _008571_, _008572_, _008573_, _008574_, _008575_, _008576_, _008577_, _008578_, _008579_, _008580_, _008581_, _008582_, _008583_, _008584_, _008585_, _008586_, _008587_, _008588_, _008589_, _008590_, _008591_, _008592_, _008593_, _008594_, _008595_, _008596_, _008597_, _008598_, _008599_, _008600_, _008601_, _008602_, _008603_, _008604_, _008605_, _008606_, _008607_, _008608_, _008609_, _008610_, _008611_, _008612_, _008613_, _008614_, _008615_, _008616_, _008617_, _008618_, _008619_, _008620_, _008621_, _008622_, _008623_, _008624_, _008625_, _008626_, _008627_, _008628_, _008629_, _008630_, _008631_, _008632_, _008633_, _008634_, _008635_, _008636_, _008637_, _008638_, _008639_, _008640_, _008641_, _008642_, _008643_, _008644_, _008645_, _008646_, _008647_, _008648_, _008649_, _008650_, _008651_, _008652_, _008653_, _008654_, _008655_, _008656_, _008657_, _008658_, _008659_, _008660_, _008661_, _008662_, _008663_, _008664_, _008665_, _008666_, _008667_, _008668_, _008669_, _008670_, _008671_, _008672_, _008673_, _008674_, _008675_, _008676_, _008677_, _008678_, _008679_, _008680_, _008681_, _008682_, _008683_, _008684_, _008685_, _008686_, _008687_, _008688_, _008689_, _008690_, _008691_, _008692_, _008693_, _008694_, _008695_, _008696_, _008697_, _008698_, _008699_, _008700_, _008701_, _008702_, _008703_, _008704_, _008705_, _008706_, _008707_, _008708_, _008709_, _008710_, _008711_, _008712_, _008713_, _008714_, _008715_, _008716_, _008717_, _008718_, _008719_, _008720_, _008721_, _008722_, _008723_, _008724_, _008725_, _008726_, _008727_, _008728_, _008729_, _008730_, _008731_, _008732_, _008733_, _008734_, _008735_, _008736_, _008737_, _008738_, _008739_, _008740_, _008741_, _008742_, _008743_, _008744_, _008745_, _008746_, _008747_, _008748_, _008749_, _008750_, _008751_, _008752_, _008753_, _008754_, _008755_, _008756_, _008757_, _008758_, _008759_, _008760_, _008761_, _008762_, _008763_, _008764_, _008765_, _008766_, _008767_, _008768_, _008769_, _008770_, _008771_, _008772_, _008773_, _008774_, _008775_, _008776_, _008777_, _008778_, _008779_, _008780_, _008781_, _008782_, _008783_, _008784_, _008785_, _008786_, _008787_, _008788_, _008789_, _008790_, _008791_, _008792_, _008793_, _008794_, _008795_, _008796_, _008797_, _008798_, _008799_, _008800_, _008801_, _008802_, _008803_, _008804_, _008805_, _008806_, _008807_, _008808_, _008809_, _008810_, _008811_, _008812_, _008813_, _008814_, _008815_, _008816_, _008817_, _008818_, _008819_, _008820_, _008821_, _008822_, _008823_, _008824_, _008825_, _008826_, _008827_, _008828_, _008829_, _008830_, _008831_, _008832_, _008833_, _008834_, _008835_, _008836_, _008837_, _008838_, _008839_, _008840_, _008841_, _008842_, _008843_, _008844_, _008845_, _008846_, _008847_, _008848_, _008849_, _008850_, _008851_, _008852_, _008853_, _008854_, _008855_, _008856_, _008857_, _008858_, _008859_, _008860_, _008861_, _008862_, _008863_, _008864_, _008865_, _008866_, _008867_, _008868_, _008869_, _008870_, _008871_, _008872_, _008873_, _008874_, _008875_, _008876_, _008877_, _008878_, _008879_, _008880_, _008881_, _008882_, _008883_, _008884_, _008885_, _008886_, _008887_, _008888_, _008889_, _008890_, _008891_, _008892_, _008893_, _008894_, _008895_, _008896_, _008897_, _008898_, _008899_, _008900_, _008901_, _008902_, _008903_, _008904_, _008905_, _008906_, _008907_, _008908_, _008909_, _008910_, _008911_, _008912_, _008913_, _008914_, _008915_, _008916_, _008917_, _008918_, _008919_, _008920_, _008921_, _008922_, _008923_, _008924_, _008925_, _008926_, _008927_, _008928_, _008929_, _008930_, _008931_, _008932_, _008933_, _008934_, _008935_, _008936_, _008937_, _008938_, _008939_, _008940_, _008941_, _008942_, _008943_, _008944_, _008945_, _008946_, _008947_, _008948_, _008949_, _008950_, _008951_, _008952_, _008953_, _008954_, _008955_, _008956_, _008957_, _008958_, _008959_, _008960_, _008961_, _008962_, _008963_, _008964_, _008965_, _008966_, _008967_, _008968_, _008969_, _008970_, _008971_, _008972_, _008973_, _008974_, _008975_, _008976_, _008977_, _008978_, _008979_, _008980_, _008981_, _008982_, _008983_, _008984_, _008985_, _008986_, _008987_, _008988_, _008989_, _008990_, _008991_, _008992_, _008993_, _008994_, _008995_, _008996_, _008997_, _008998_, _008999_, _009000_, _009001_, _009002_, _009003_, _009004_, _009005_, _009006_, _009007_, _009008_, _009009_, _009010_, _009011_, _009012_, _009013_, _009014_, _009015_, _009016_, _009017_, _009018_, _009019_, _009020_, _009021_, _009022_, _009023_, _009024_, _009025_, _009026_, _009027_, _009028_, _009029_, _009030_, _009031_, _009032_, _009033_, _009034_, _009035_, _009036_, _009037_, _009038_, _009039_, _009040_, _009041_, _009042_, _009043_, _009044_, _009045_, _009046_, _009047_, _009048_, _009049_, _009050_, _009051_, _009052_, _009053_, _009054_, _009055_, _009056_, _009057_, _009058_, _009059_, _009060_, _009061_, _009062_, _009063_, _009064_, _009065_, _009066_, _009067_, _009068_, _009069_, _009070_, _009071_, _009072_, _009073_, _009074_, _009075_, _009076_, _009077_, _009078_, _009079_, _009080_, _009081_, _009082_, _009083_, _009084_, _009085_, _009086_, _009087_, _009088_, _009089_, _009090_, _009091_, _009092_, _009093_, _009094_, _009095_, _009096_, _009097_, _009098_, _009099_, _009100_, _009101_, _009102_, _009103_, _009104_, _009105_, _009106_, _009107_, _009108_, _009109_, _009110_, _009111_, _009112_, _009113_, _009114_, _009115_, _009116_, _009117_, _009118_, _009119_, _009120_, _009121_, _009122_, _009123_, _009124_, _009125_, _009126_, _009127_, _009128_, _009129_, _009130_, _009131_, _009132_, _009133_, _009134_, _009135_, _009136_, _009137_, _009138_, _009139_, _009140_, _009141_, _009142_, _009143_, _009144_, _009145_, _009146_, _009147_, _009148_, _009149_, _009150_, _009151_, _009152_, _009153_, _009154_, _009155_, _009156_, _009157_, _009158_, _009159_, _009160_, _009161_, _009162_, _009163_, _009164_, _009165_, _009166_, _009167_, _009168_, _009169_, _009170_, _009171_, _009172_, _009173_, _009174_, _009175_, _009176_, _009177_, _009178_, _009179_, _009180_, _009181_, _009182_, _009183_, _009184_, _009185_, _009186_, _009187_, _009188_, _009189_, _009190_, _009191_, _009192_, _009193_, _009194_, _009195_, _009196_, _009197_, _009198_, _009199_, _009200_, _009201_, _009202_, _009203_, _009204_, _009205_, _009206_, _009207_, _009208_, _009209_, _009210_, _009211_, _009212_, _009213_, _009214_, _009215_, _009216_, _009217_, _009218_, _009219_, _009220_, _009221_, _009222_, _009223_, _009224_, _009225_, _009226_, _009227_, _009228_, _009229_, _009230_, _009231_, _009232_, _009233_, _009234_, _009235_, _009236_, _009237_, _009238_, _009239_, _009240_, _009241_, _009242_, _009243_, _009244_, _009245_, _009246_, _009247_, _009248_, _009249_, _009250_, _009251_, _009252_, _009253_, _009254_, _009255_, _009256_, _009257_, _009258_, _009259_, _009260_, _009261_, _009262_, _009263_, _009264_, _009265_, _009266_, _009267_, _009268_, _009269_, _009270_, _009271_, _009272_, _009273_, _009274_, _009275_, _009276_, _009277_, _009278_, _009279_, _009280_, _009281_, _009282_, _009283_, _009284_, _009285_, _009286_, _009287_, _009288_, _009289_, _009290_, _009291_, _009292_, _009293_, _009294_, _009295_, _009296_, _009297_, _009298_, _009299_, _009300_, _009301_, _009302_, _009303_, _009304_, _009305_, _009306_, _009307_, _009308_, _009309_, _009310_, _009311_, _009312_, _009313_, _009314_, _009315_, _009316_, _009317_, _009318_, _009319_, _009320_, _009321_, _009322_, _009323_, _009324_, _009325_, _009326_, _009327_, _009328_, _009329_, _009330_, _009331_, _009332_, _009333_, _009334_, _009335_, _009336_, _009337_, _009338_, _009339_, _009340_, _009341_, _009342_, _009343_, _009344_, _009345_, _009346_, _009347_, _009348_, _009349_, _009350_, _009351_, _009352_, _009353_, _009354_, _009355_, _009356_, _009357_, _009358_, _009359_, _009360_, _009361_, _009362_, _009363_, _009364_, _009365_, _009366_, _009367_, _009368_, _009369_, _009370_, _009371_, _009372_, _009373_, _009374_, _009375_, _009376_, _009377_, _009378_, _009379_, _009380_, _009381_, _009382_, _009383_, _009384_, _009385_, _009386_, _009387_, _009388_, _009389_, _009390_, _009391_, _009392_, _009393_, _009394_, _009395_, _009396_, _009397_, _009398_, _009399_, _009400_, _009401_, _009402_, _009403_, _009404_, _009405_, _009406_, _009407_, _009408_, _009409_, _009410_, _009411_, _009412_, _009413_, _009414_, _009415_, _009416_, _009417_, _009418_, _009419_, _009420_, _009421_, _009422_, _009423_, _009424_, _009425_, _009426_, _009427_, _009428_, _009429_, _009430_, _009431_, _009432_, _009433_, _009434_, _009435_, _009436_, _009437_, _009438_, _009439_, _009440_, _009441_, _009442_, _009443_, _009444_, _009445_, _009446_, _009447_, _009448_, _009449_, _009450_, _009451_, _009452_, _009453_, _009454_, _009455_, _009456_, _009457_, _009458_, _009459_, _009460_, _009461_, _009462_, _009463_, _009464_, _009465_, _009466_, _009467_, _009468_, _009469_, _009470_, _009471_, _009472_, _009473_, _009474_, _009475_, _009476_, _009477_, _009478_, _009479_, _009480_, _009481_, _009482_, _009483_, _009484_, _009485_, _009486_, _009487_, _009488_, _009489_, _009490_, _009491_, _009492_, _009493_, _009494_, _009495_, _009496_, _009497_, _009498_, _009499_, _009500_, _009501_, _009502_, _009503_, _009504_, _009505_, _009506_, _009507_, _009508_, _009509_, _009510_, _009511_, _009512_, _009513_, _009514_, _009515_, _009516_, _009517_, _009518_, _009519_, _009520_, _009521_, _009522_, _009523_, _009524_, _009525_, _009526_, _009527_, _009528_, _009529_, _009530_, _009531_, _009532_, _009533_, _009534_, _009535_, _009536_, _009537_, _009538_, _009539_, _009540_, _009541_, _009542_, _009543_, _009544_, _009545_, _009546_, _009547_, _009548_, _009549_, _009550_, _009551_, _009552_, _009553_, _009554_, _009555_, _009556_, _009557_, _009558_, _009559_, _009560_, _009561_, _009562_, _009563_, _009564_, _009565_, _009566_, _009567_, _009568_, _009569_, _009570_, _009571_, _009572_, _009573_, _009574_, _009575_, _009576_, _009577_, _009578_, _009579_, _009580_, _009581_, _009582_, _009583_, _009584_, _009585_, _009586_, _009587_, _009588_, _009589_, _009590_, _009591_, _009592_, _009593_, _009594_, _009595_, _009596_, _009597_, _009598_, _009599_, _009600_, _009601_, _009602_, _009603_, _009604_, _009605_, _009606_, _009607_, _009608_, _009609_, _009610_, _009611_, _009612_, _009613_, _009614_, _009615_, _009616_, _009617_, _009618_, _009619_, _009620_, _009621_, _009622_, _009623_, _009624_, _009625_, _009626_, _009627_, _009628_, _009629_, _009630_, _009631_, _009632_, _009633_, _009634_, _009635_, _009636_, _009637_, _009638_, _009639_, _009640_, _009641_, _009642_, _009643_, _009644_, _009645_, _009646_, _009647_, _009648_, _009649_, _009650_, _009651_, _009652_, _009653_, _009654_, _009655_, _009656_, _009657_, _009658_, _009659_, _009660_, _009661_, _009662_, _009663_, _009664_, _009665_, _009666_, _009667_, _009668_, _009669_, _009670_, _009671_, _009672_, _009673_, _009674_, _009675_, _009676_, _009677_, _009678_, _009679_, _009680_, _009681_, _009682_, _009683_, _009684_, _009685_, _009686_, _009687_, _009688_, _009689_, _009690_, _009691_, _009692_, _009693_, _009694_, _009695_, _009696_, _009697_, _009698_, _009699_, _009700_, _009701_, _009702_, _009703_, _009704_, _009705_, _009706_, _009707_, _009708_, _009709_, _009710_, _009711_, _009712_, _009713_, _009714_, _009715_, _009716_, _009717_, _009718_, _009719_, _009720_, _009721_, _009722_, _009723_, _009724_, _009725_, _009726_, _009727_, _009728_, _009729_, _009730_, _009731_, _009732_, _009733_, _009734_, _009735_, _009736_, _009737_, _009738_, _009739_, _009740_, _009741_, _009742_, _009743_, _009744_, _009745_, _009746_, _009747_, _009748_, _009749_, _009750_, _009751_, _009752_, _009753_, _009754_, _009755_, _009756_, _009757_, _009758_, _009759_, _009760_, _009761_, _009762_, _009763_, _009764_, _009765_, _009766_, _009767_, _009768_, _009769_, _009770_, _009771_, _009772_, _009773_, _009774_, _009775_, _009776_, _009777_, _009778_, _009779_, _009780_, _009781_, _009782_, _009783_, _009784_, _009785_, _009786_, _009787_, _009788_, _009789_, _009790_, _009791_, _009792_, _009793_, _009794_, _009795_, _009796_, _009797_, _009798_, _009799_, _009800_, _009801_, _009802_, _009803_, _009804_, _009805_, _009806_, _009807_, _009808_, _009809_, _009810_, _009811_, _009812_, _009813_, _009814_, _009815_, _009816_, _009817_, _009818_, _009819_, _009820_, _009821_, _009822_, _009823_, _009824_, _009825_, _009826_, _009827_, _009828_, _009829_, _009830_, _009831_, _009832_, _009833_, _009834_, _009835_, _009836_, _009837_, _009838_, _009839_, _009840_, _009841_, _009842_, _009843_, _009844_, _009845_, _009846_, _009847_, _009848_, _009849_, _009850_, _009851_, _009852_, _009853_, _009854_, _009855_, _009856_, _009857_, _009858_, _009859_, _009860_, _009861_, _009862_, _009863_, _009864_, _009865_, _009866_, _009867_, _009868_, _009869_, _009870_, _009871_, _009872_, _009873_, _009874_, _009875_, _009876_, _009877_, _009878_, _009879_, _009880_, _009881_, _009882_, _009883_, _009884_, _009885_, _009886_, _009887_, _009888_, _009889_, _009890_, _009891_, _009892_, _009893_, _009894_, _009895_, _009896_, _009897_, _009898_, _009899_, _009900_, _009901_, _009902_, _009903_, _009904_, _009905_, _009906_, _009907_, _009908_, _009909_, _009910_, _009911_, _009912_, _009913_, _009914_, _009915_, _009916_, _009917_, _009918_, _009919_, _009920_, _009921_, _009922_, _009923_, _009924_, _009925_, _009926_, _009927_, _009928_, _009929_, _009930_, _009931_, _009932_, _009933_, _009934_, _009935_, _009936_, _009937_, _009938_, _009939_, _009940_, _009941_, _009942_, _009943_, _009944_, _009945_, _009946_, _009947_, _009948_, _009949_, _009950_, _009951_, _009952_, _009953_, _009954_, _009955_, _009956_, _009957_, _009958_, _009959_, _009960_, _009961_, _009962_, _009963_, _009964_, _009965_, _009966_, _009967_, _009968_, _009969_, _009970_, _009971_, _009972_, _009973_, _009974_, _009975_, _009976_, _009977_, _009978_, _009979_, _009980_, _009981_, _009982_, _009983_, _009984_, _009985_, _009986_, _009987_, _009988_, _009989_, _009990_, _009991_, _009992_, _009993_, _009994_, _009995_, _009996_, _009997_, _009998_, _009999_, _010000_, _010001_, _010002_, _010003_, _010004_, _010005_, _010006_, _010007_, _010008_, _010009_, _010010_, _010011_, _010012_, _010013_, _010014_, _010015_, _010016_, _010017_, _010018_, _010019_, _010020_, _010021_, _010022_, _010023_, _010024_, _010025_, _010026_, _010027_, _010028_, _010029_, _010030_, _010031_, _010032_, _010033_, _010034_, _010035_, _010036_, _010037_, _010038_, _010039_, _010040_, _010041_, _010042_, _010043_, _010044_, _010045_, _010046_, _010047_, _010048_, _010049_, _010050_, _010051_, _010052_, _010053_, _010054_, _010055_, _010056_, _010057_, _010058_, _010059_, _010060_, _010061_, _010062_, _010063_, _010064_, _010065_, _010066_, _010067_, _010068_, _010069_, _010070_, _010071_, _010072_, _010073_, _010074_, _010075_, _010076_, _010077_, _010078_, _010079_, _010080_, _010081_, _010082_, _010083_, _010084_, _010085_, _010086_, _010087_, _010088_, _010089_, _010090_, _010091_, _010092_, _010093_, _010094_, _010095_, _010096_, _010097_, _010098_, _010099_, _010100_, _010101_, _010102_, _010103_, _010104_, _010105_, _010106_, _010107_, _010108_, _010109_, _010110_, _010111_, _010112_, _010113_, _010114_, _010115_, _010116_, _010117_, _010118_, _010119_, _010120_, _010121_, _010122_, _010123_, _010124_, _010125_, _010126_, _010127_, _010128_, _010129_, _010130_, _010131_, _010132_, _010133_, _010134_, _010135_, _010136_, _010137_, _010138_, _010139_, _010140_, _010141_, _010142_, _010143_, _010144_, _010145_, _010146_, _010147_, _010148_, _010149_, _010150_, _010151_, _010152_, _010153_, _010154_, _010155_, _010156_, _010157_, _010158_, _010159_, _010160_, _010161_, _010162_, _010163_, _010164_, _010165_, _010166_, _010167_, _010168_, _010169_, _010170_, _010171_, _010172_, _010173_, _010174_, _010175_, _010176_, _010177_, _010178_, _010179_, _010180_, _010181_, _010182_, _010183_, _010184_, _010185_, _010186_, _010187_, _010188_, _010189_, _010190_, _010191_, _010192_, _010193_, _010194_, _010195_, _010196_, _010197_, _010198_, _010199_, _010200_, _010201_, _010202_, _010203_, _010204_, _010205_, _010206_, _010207_, _010208_, _010209_, _010210_, _010211_, _010212_, _010213_, _010214_, _010215_, _010216_, _010217_, _010218_, _010219_, _010220_, _010221_, _010222_, _010223_, _010224_, _010225_, _010226_, _010227_, _010228_, _010229_, _010230_, _010231_, _010232_, _010233_, _010234_, _010235_, _010236_, _010237_, _010238_, _010239_, _010240_, _010241_, _010242_, _010243_, _010244_, _010245_, _010246_, _010247_, _010248_, _010249_, _010250_, _010251_, _010252_, _010253_, _010254_, _010255_, _010256_, _010257_, _010258_, _010259_, _010260_, _010261_, _010262_, _010263_, _010264_, _010265_, _010266_, _010267_, _010268_, _010269_, _010270_, _010271_, _010272_, _010273_, _010274_, _010275_, _010276_, _010277_, _010278_, _010279_, _010280_, _010281_, _010282_, _010283_, _010284_, _010285_, _010286_, _010287_, _010288_, _010289_, _010290_, _010291_, _010292_, _010293_, _010294_, _010295_, _010296_, _010297_, _010298_, _010299_, _010300_, _010301_, _010302_, _010303_, _010304_, _010305_, _010306_, _010307_, _010308_, _010309_, _010310_, _010311_, _010312_, _010313_, _010314_, _010315_, _010316_, _010317_, _010318_, _010319_, _010320_, _010321_, _010322_, _010323_, _010324_, _010325_, _010326_, _010327_, _010328_, _010329_, _010330_, _010331_, _010332_, _010333_, _010334_, _010335_, _010336_, _010337_, _010338_, _010339_, _010340_, _010341_, _010342_, _010343_, _010344_, _010345_, _010346_, _010347_, _010348_, _010349_, _010350_, _010351_, _010352_, _010353_, _010354_, _010355_, _010356_, _010357_, _010358_, _010359_, _010360_, _010361_, _010362_, _010363_, _010364_, _010365_, _010366_, _010367_, _010368_, _010369_, _010370_, _010371_, _010372_, _010373_, _010374_, _010375_, _010376_, _010377_, _010378_, _010379_, _010380_, _010381_, _010382_, _010383_, _010384_, _010385_, _010386_, _010387_, _010388_, _010389_, _010390_, _010391_, _010392_, _010393_, _010394_, _010395_, _010396_, _010397_, _010398_, _010399_, _010400_, _010401_, _010402_, _010403_, _010404_, _010405_, _010406_, _010407_, _010408_, _010409_, _010410_, _010411_, _010412_, _010413_, _010414_, _010415_, _010416_, _010417_, _010418_, _010419_, _010420_, _010421_, _010422_, _010423_, _010424_, _010425_, _010426_, _010427_, _010428_, _010429_, _010430_, _010431_, _010432_, _010433_, _010434_, _010435_, _010436_, _010437_, _010438_, _010439_, _010440_, _010441_, _010442_, _010443_, _010444_, _010445_, _010446_, _010447_, _010448_, _010449_, _010450_, _010451_, _010452_, _010453_, _010454_, _010455_, _010456_, _010457_, _010458_, _010459_, _010460_, _010461_, _010462_, _010463_, _010464_, _010465_, _010466_, _010467_, _010468_, _010469_, _010470_, _010471_, _010472_, _010473_, _010474_, _010475_, _010476_, _010477_, _010478_, _010479_, _010480_, _010481_, _010482_, _010483_, _010484_, _010485_, _010486_, _010487_, _010488_, _010489_, _010490_, _010491_, _010492_, _010493_, _010494_, _010495_, _010496_, _010497_, _010498_, _010499_, _010500_, _010501_, _010502_, _010503_, _010504_, _010505_, _010506_, _010507_, _010508_, _010509_, _010510_, _010511_, _010512_, _010513_, _010514_, _010515_, _010516_, _010517_, _010518_, _010519_, _010520_, _010521_, _010522_, _010523_, _010524_, _010525_, _010526_, _010527_, _010528_, _010529_, _010530_, _010531_, _010532_, _010533_, _010534_, _010535_, _010536_, _010537_, _010538_, _010539_, _010540_, _010541_, _010542_, _010543_, _010544_, _010545_, _010546_, _010547_, _010548_, _010549_, _010550_, _010551_, _010552_, _010553_, _010554_, _010555_, _010556_, _010557_, _010558_, _010559_, _010560_, _010561_, _010562_, _010563_, _010564_, _010565_, _010566_, _010567_, _010568_, _010569_, _010570_, _010571_, _010572_, _010573_, _010574_, _010575_, _010576_, _010577_, _010578_, _010579_, _010580_, _010581_, _010582_, _010583_, _010584_, _010585_, _010586_, _010587_, _010588_, _010589_, _010590_, _010591_, _010592_, _010593_, _010594_, _010595_, _010596_, _010597_, _010598_, _010599_, _010600_, _010601_, _010602_, _010603_, _010604_, _010605_, _010606_, _010607_, _010608_, _010609_, _010610_, _010611_, _010612_, _010613_, _010614_, _010615_, _010616_, _010617_, _010618_, _010619_, _010620_, _010621_, _010622_, _010623_, _010624_, _010625_, _010626_, _010627_, _010628_, _010629_, _010630_, _010631_, _010632_, _010633_, _010634_, _010635_, _010636_, _010637_, _010638_, _010639_, _010640_, _010641_, _010642_, _010643_, _010644_, _010645_, _010646_, _010647_, _010648_, _010649_, _010650_, _010651_, _010652_, _010653_, _010654_, _010655_, _010656_, _010657_, _010658_, _010659_, _010660_, _010661_, _010662_, _010663_, _010664_, _010665_, _010666_, _010667_, _010668_, _010669_, _010670_, _010671_, _010672_, _010673_, _010674_, _010675_, _010676_, _010677_, _010678_, _010679_, _010680_, _010681_, _010682_, _010683_, _010684_, _010685_, _010686_, _010687_, _010688_, _010689_, _010690_, _010691_, _010692_, _010693_, _010694_, _010695_, _010696_, _010697_, _010698_, _010699_, _010700_, _010701_, _010702_, _010703_, _010704_, _010705_, _010706_, _010707_, _010708_, _010709_, _010710_, _010711_, _010712_, _010713_, _010714_, _010715_, _010716_, _010717_, _010718_, _010719_, _010720_, _010721_, _010722_, _010723_, _010724_, _010725_, _010726_, _010727_, _010728_, _010729_, _010730_, _010731_, _010732_, _010733_, _010734_, _010735_, _010736_, _010737_, _010738_, _010739_, _010740_, _010741_, _010742_, _010743_, _010744_, _010745_, _010746_, _010747_, _010748_, _010749_, _010750_, _010751_, _010752_, _010753_, _010754_, _010755_, _010756_, _010757_, _010758_, _010759_, _010760_, _010761_, _010762_, _010763_, _010764_, _010765_, _010766_, _010767_, _010768_, _010769_, _010770_, _010771_, _010772_, _010773_, _010774_, _010775_, _010776_, _010777_, _010778_, _010779_, _010780_, _010781_, _010782_, _010783_, _010784_, _010785_, _010786_, _010787_, _010788_, _010789_, _010790_, _010791_, _010792_, _010793_, _010794_, _010795_, _010796_, _010797_, _010798_, _010799_, _010800_, _010801_, _010802_, _010803_, _010804_, _010805_, _010806_, _010807_, _010808_, _010809_, _010810_, _010811_, _010812_, _010813_, _010814_, _010815_, _010816_, _010817_, _010818_, _010819_, _010820_, _010821_, _010822_, _010823_, _010824_, _010825_, _010826_, _010827_, _010828_, _010829_, _010830_, _010831_, _010832_, _010833_, _010834_, _010835_, _010836_, _010837_, _010838_, _010839_, _010840_, _010841_, _010842_, _010843_, _010844_, _010845_, _010846_, _010847_, _010848_, _010849_, _010850_, _010851_, _010852_, _010853_, _010854_, _010855_, _010856_, _010857_, _010858_, _010859_, _010860_, _010861_, _010862_, _010863_, _010864_, _010865_, _010866_, _010867_, _010868_, _010869_, _010870_, _010871_, _010872_, _010873_, _010874_, _010875_, _010876_, _010877_, _010878_, _010879_, _010880_, _010881_, _010882_, _010883_, _010884_, _010885_, _010886_, _010887_, _010888_, _010889_, _010890_, _010891_, _010892_, _010893_, _010894_, _010895_, _010896_, _010897_, _010898_, _010899_, _010900_, _010901_, _010902_, _010903_, _010904_, _010905_, _010906_, _010907_, _010908_, _010909_, _010910_, _010911_, _010912_, _010913_, _010914_, _010915_, _010916_, _010917_, _010918_, _010919_, _010920_, _010921_, _010922_, _010923_, _010924_, _010925_, _010926_, _010927_, _010928_, _010929_, _010930_, _010931_, _010932_, _010933_, _010934_, _010935_, _010936_, _010937_, _010938_, _010939_, _010940_, _010941_, _010942_, _010943_, _010944_, _010945_, _010946_, _010947_, _010948_, _010949_, _010950_, _010951_, _010952_, _010953_, _010954_, _010955_, _010956_, _010957_, _010958_, _010959_, _010960_, _010961_, _010962_, _010963_, _010964_, _010965_, _010966_, _010967_, _010968_, _010969_, _010970_, _010971_, _010972_, _010973_, _010974_, _010975_, _010976_, _010977_, _010978_, _010979_, _010980_, _010981_, _010982_, _010983_, _010984_, _010985_, _010986_, _010987_, _010988_, _010989_, _010990_, _010991_, _010992_, _010993_, _010994_, _010995_, _010996_, _010997_, _010998_, _010999_, _011000_, _011001_, _011002_, _011003_, _011004_, _011005_, _011006_, _011007_, _011008_, _011009_, _011010_, _011011_, _011012_, _011013_, _011014_, _011015_, _011016_, _011017_, _011018_, _011019_, _011020_, _011021_, _011022_, _011023_, _011024_, _011025_, _011026_, _011027_, _011028_, _011029_, _011030_, _011031_, _011032_, _011033_, _011034_, _011035_, _011036_, _011037_, _011038_, _011039_, _011040_, _011041_, _011042_, _011043_, _011044_, _011045_, _011046_, _011047_, _011048_, _011049_, _011050_, _011051_, _011052_, _011053_, _011054_, _011055_, _011056_, _011057_, _011058_, _011059_, _011060_, _011061_, _011062_, _011063_, _011064_, _011065_, _011066_, _011067_, _011068_, _011069_, _011070_, _011071_, _011072_, _011073_, _011074_, _011075_, _011076_, _011077_, _011078_, _011079_, _011080_, _011081_, _011082_, _011083_, _011084_, _011085_, _011086_, _011087_, _011088_, _011089_, _011090_, _011091_, _011092_, _011093_, _011094_, _011095_, _011096_, _011097_, _011098_, _011099_, _011100_, _011101_, _011102_, _011103_, _011104_, _011105_, _011106_, _011107_, _011108_, _011109_, _011110_, _011111_, _011112_, _011113_, _011114_, _011115_, _011116_, _011117_, _011118_, _011119_, _011120_, _011121_, _011122_, _011123_, _011124_, _011125_, _011126_, _011127_, _011128_, _011129_, _011130_, _011131_, _011132_, _011133_, _011134_, _011135_, _011136_, _011137_, _011138_, _011139_, _011140_, _011141_, _011142_, _011143_, _011144_, _011145_, _011146_, _011147_, _011148_, _011149_, _011150_, _011151_, _011152_, _011153_, _011154_, _011155_, _011156_, _011157_, _011158_, _011159_, _011160_, _011161_, _011162_, _011163_, _011164_, _011165_, _011166_, _011167_, _011168_, _011169_, _011170_, _011171_, _011172_, _011173_, _011174_, _011175_, _011176_, _011177_, _011178_, _011179_, _011180_, _011181_, _011182_, _011183_, _011184_, _011185_, _011186_, _011187_, _011188_, _011189_, _011190_, _011191_, _011192_, _011193_, _011194_, _011195_, _011196_, _011197_, _011198_, _011199_, _011200_, _011201_, _011202_, _011203_, _011204_, _011205_, _011206_, _011207_, _011208_, _011209_, _011210_, _011211_, _011212_, _011213_, _011214_, _011215_, _011216_, _011217_, _011218_, _011219_, _011220_, _011221_, _011222_, _011223_, _011224_, _011225_, _011226_, _011227_, _011228_, _011229_, _011230_, _011231_, _011232_, _011233_, _011234_, _011235_, _011236_, _011237_, _011238_, _011239_, _011240_, _011241_, _011242_, _011243_, _011244_, _011245_, _011246_, _011247_, _011248_, _011249_, _011250_, _011251_, _011252_, _011253_, _011254_, _011255_, _011256_, _011257_, _011258_, _011259_, _011260_, _011261_, _011262_, _011263_, _011264_, _011265_, _011266_, _011267_, _011268_, _011269_, _011270_, _011271_, _011272_, _011273_, _011274_, _011275_, _011276_, _011277_, _011278_, _011279_, _011280_, _011281_, _011282_, _011283_, _011284_, _011285_, _011286_, _011287_, _011288_, _011289_, _011290_, _011291_, _011292_, _011293_, _011294_, _011295_, _011296_, _011297_, _011298_, _011299_, _011300_, _011301_, _011302_, _011303_, _011304_, _011305_, _011306_, _011307_, _011308_, _011309_, _011310_, _011311_, _011312_, _011313_, _011314_, _011315_, _011316_, _011317_, _011318_, _011319_, _011320_, _011321_, _011322_, _011323_, _011324_, _011325_, _011326_, _011327_, _011328_, _011329_, _011330_, _011331_, _011332_, _011333_, _011334_, _011335_, _011336_, _011337_, _011338_, _011339_, _011340_, _011341_, _011342_, _011343_, _011344_, _011345_, _011346_, _011347_, _011348_, _011349_, _011350_, _011351_, _011352_, _011353_, _011354_, _011355_, _011356_, _011357_, _011358_, _011359_, _011360_, _011361_, _011362_, _011363_, _011364_, _011365_, _011366_, _011367_, _011368_, _011369_, _011370_, _011371_, _011372_, _011373_, _011374_, _011375_, _011376_, _011377_, _011378_, _011379_, _011380_, _011381_, _011382_, _011383_, _011384_, _011385_, _011386_, _011387_, _011388_, _011389_, _011390_, _011391_, _011392_, _011393_, _011394_, _011395_, _011396_, _011397_, _011398_, _011399_, _011400_, _011401_, _011402_, _011403_, _011404_, _011405_, _011406_, _011407_, _011408_, _011409_, _011410_, _011411_, _011412_, _011413_, _011414_, _011415_, _011416_, _011417_, _011418_, _011419_, _011420_, _011421_, _011422_, _011423_, _011424_, _011425_, _011426_, _011427_, _011428_, _011429_, _011430_, _011431_, _011432_, _011433_, _011434_, _011435_, _011436_, _011437_, _011438_, _011439_, _011440_, _011441_, _011442_, _011443_, _011444_, _011445_, _011446_, _011447_, _011448_, _011449_, _011450_, _011451_, _011452_, _011453_, _011454_, _011455_, _011456_, _011457_, _011458_, _011459_, _011460_, _011461_, _011462_, _011463_, _011464_, _011465_, _011466_, _011467_, _011468_, _011469_, _011470_, _011471_, _011472_, _011473_, _011474_, _011475_, _011476_, _011477_, _011478_, _011479_, _011480_, _011481_, _011482_, _011483_, _011484_, _011485_, _011486_, _011487_, _011488_, _011489_, _011490_, _011491_, _011492_, _011493_, _011494_, _011495_, _011496_, _011497_, _011498_, _011499_, _011500_, _011501_, _011502_, _011503_, _011504_, _011505_, _011506_, _011507_, _011508_, _011509_, _011510_, _011511_, _011512_, _011513_, _011514_, _011515_, _011516_, _011517_, _011518_, _011519_, _011520_, _011521_, _011522_, _011523_, _011524_, _011525_, _011526_, _011527_, _011528_, _011529_, _011530_, _011531_, _011532_, _011533_, _011534_, _011535_, _011536_, _011537_, _011538_, _011539_, _011540_, _011541_, _011542_, _011543_, _011544_, _011545_, _011546_, _011547_, _011548_, _011549_, _011550_, _011551_, _011552_, _011553_, _011554_, _011555_, _011556_, _011557_, _011558_, _011559_, _011560_, _011561_, _011562_, _011563_, _011564_, _011565_, _011566_, _011567_, _011568_, _011569_, _011570_, _011571_, _011572_, _011573_, _011574_, _011575_, _011576_, _011577_, _011578_, _011579_, _011580_, _011581_, _011582_, _011583_, _011584_, _011585_, _011586_, _011587_, _011588_, _011589_, _011590_, _011591_, _011592_, _011593_, _011594_, _011595_, _011596_, _011597_, _011598_, _011599_, _011600_, _011601_, _011602_, _011603_, _011604_, _011605_, _011606_, _011607_, _011608_, _011609_, _011610_, _011611_, _011612_, _011613_, _011614_, _011615_, _011616_, _011617_, _011618_, _011619_, _011620_, _011621_, _011622_, _011623_, _011624_, _011625_, _011626_, _011627_, _011628_, _011629_, _011630_, _011631_, _011632_, _011633_, _011634_, _011635_, _011636_, _011637_, _011638_, _011639_, _011640_, _011641_, _011642_, _011643_, _011644_, _011645_, _011646_, _011647_, _011648_, _011649_, _011650_, _011651_, _011652_, _011653_, _011654_, _011655_, _011656_, _011657_, _011658_, _011659_, _011660_, _011661_, _011662_, _011663_, _011664_, _011665_, _011666_, _011667_, _011668_, _011669_, _011670_, _011671_, _011672_, _011673_, _011674_, _011675_, _011676_, _011677_, _011678_, _011679_, _011680_, _011681_, _011682_, _011683_, _011684_, _011685_, _011686_, _011687_, _011688_, _011689_, _011690_, _011691_, _011692_, _011693_, _011694_, _011695_, _011696_, _011697_, _011698_, _011699_, _011700_, _011701_, _011702_, _011703_, _011704_, _011705_, _011706_, _011707_, _011708_, _011709_, _011710_, _011711_, _011712_, _011713_, _011714_, _011715_, _011716_, _011717_, _011718_, _011719_, _011720_, _011721_, _011722_, _011723_, _011724_, _011725_, _011726_, _011727_, _011728_, _011729_, _011730_, _011731_, _011732_, _011733_, _011734_, _011735_, _011736_, _011737_, _011738_, _011739_, _011740_, _011741_, _011742_, _011743_, _011744_, _011745_, _011746_, _011747_, _011748_, _011749_, _011750_, _011751_, _011752_, _011753_, _011754_, _011755_, _011756_, _011757_, _011758_, _011759_, _011760_, _011761_, _011762_, _011763_, _011764_, _011765_, _011766_, _011767_, _011768_, _011769_, _011770_, _011771_, _011772_, _011773_, _011774_, _011775_, _011776_, _011777_, _011778_, _011779_, _011780_, _011781_, _011782_, _011783_, _011784_, _011785_, _011786_, _011787_, _011788_, _011789_, _011790_, _011791_, _011792_, _011793_, _011794_, _011795_, _011796_, _011797_, _011798_, _011799_, _011800_, _011801_, _011802_, _011803_, _011804_, _011805_, _011806_, _011807_, _011808_, _011809_, _011810_, _011811_, _011812_, _011813_, _011814_, _011815_, _011816_, _011817_, _011818_, _011819_, _011820_, _011821_, _011822_, _011823_, _011824_, _011825_, _011826_, _011827_, _011828_, _011829_, _011830_, _011831_, _011832_, _011833_, _011834_, _011835_, _011836_, _011837_, _011838_, _011839_, _011840_, _011841_, _011842_, _011843_, _011844_, _011845_, _011846_, _011847_, _011848_, _011849_, _011850_, _011851_, _011852_, _011853_, _011854_, _011855_, _011856_, _011857_, _011858_, _011859_, _011860_, _011861_, _011862_, _011863_, _011864_, _011865_, _011866_, _011867_, _011868_, _011869_, _011870_, _011871_, _011872_, _011873_, _011874_, _011875_, _011876_, _011877_, _011878_, _011879_, _011880_, _011881_, _011882_, _011883_, _011884_, _011885_, _011886_, _011887_, _011888_, _011889_, _011890_, _011891_, _011892_, _011893_, _011894_, _011895_, _011896_, _011897_, _011898_, _011899_, _011900_, _011901_, _011902_, _011903_, _011904_, _011905_, _011906_, _011907_, _011908_, _011909_, _011910_, _011911_, _011912_, _011913_, _011914_, _011915_, _011916_, _011917_, _011918_, _011919_, _011920_, _011921_, _011922_, _011923_, _011924_, _011925_, _011926_, _011927_, _011928_, _011929_, _011930_, _011931_, _011932_, _011933_, _011934_, _011935_, _011936_, _011937_, _011938_, _011939_, _011940_, _011941_, _011942_, _011943_, _011944_, _011945_, _011946_, _011947_, _011948_, _011949_, _011950_, _011951_, _011952_, _011953_, _011954_, _011955_, _011956_, _011957_, _011958_, _011959_, _011960_, _011961_, _011962_, _011963_, _011964_, _011965_, _011966_, _011967_, _011968_, _011969_, _011970_, _011971_, _011972_, _011973_, _011974_, _011975_, _011976_, _011977_, _011978_, _011979_, _011980_, _011981_, _011982_, _011983_, _011984_, _011985_, _011986_, _011987_, _011988_, _011989_, _011990_, _011991_, _011992_, _011993_, _011994_, _011995_, _011996_, _011997_, _011998_, _011999_, _012000_, _012001_, _012002_, _012003_, _012004_, _012005_, _012006_, _012007_, _012008_, _012009_, _012010_, _012011_, _012012_, _012013_, _012014_, _012015_, _012016_, _012017_, _012018_, _012019_, _012020_, _012021_, _012022_, _012023_, _012024_, _012025_, _012026_, _012027_, _012028_, _012029_, _012030_, _012031_, _012032_, _012033_, _012034_, _012035_, _012036_, _012037_, _012038_, _012039_, _012040_, _012041_, _012042_, _012043_, _012044_, _012045_, _012046_, _012047_, _012048_, _012049_, _012050_, _012051_, _012052_, _012053_, _012054_, _012055_, _012056_, _012057_, _012058_, _012059_, _012060_, _012061_, _012062_, _012063_, _012064_, _012065_, _012066_, _012067_, _012068_, _012069_, _012070_, _012071_, _012072_, _012073_, _012074_, _012075_, _012076_, _012077_, _012078_, _012079_, _012080_, _012081_, _012082_, _012083_, _012084_, _012085_, _012086_, _012087_, _012088_, _012089_, _012090_, _012091_, _012092_, _012093_, _012094_, _012095_, _012096_, _012097_, _012098_, _012099_, _012100_, _012101_, _012102_, _012103_, _012104_, _012105_, _012106_, _012107_, _012108_, _012109_, _012110_, _012111_, _012112_, _012113_, _012114_, _012115_, _012116_, _012117_, _012118_, _012119_, _012120_, _012121_, _012122_, _012123_, _012124_, _012125_, _012126_, _012127_, _012128_, _012129_, _012130_, _012131_, _012132_, _012133_, _012134_, _012135_, _012136_, _012137_, _012138_, _012139_, _012140_, _012141_, _012142_, _012143_, _012144_, _012145_, _012146_, _012147_, _012148_, _012149_, _012150_, _012151_, _012152_, _012153_, _012154_, _012155_, _012156_, _012157_, _012158_, _012159_, _012160_, _012161_, _012162_, _012163_, _012164_, _012165_, _012166_, _012167_, _012168_, _012169_, _012170_, _012171_, _012172_, _012173_, _012174_, _012175_, _012176_, _012177_, _012178_, _012179_, _012180_, _012181_, _012182_, _012183_, _012184_, _012185_, _012186_, _012187_, _012188_, _012189_, _012190_, _012191_, _012192_, _012193_, _012194_, _012195_, _012196_, _012197_, _012198_, _012199_, _012200_, _012201_, _012202_, _012203_, _012204_, _012205_, _012206_, _012207_, _012208_, _012209_, _012210_, _012211_, _012212_, _012213_, _012214_, _012215_, _012216_, _012217_, _012218_, _012219_, _012220_, _012221_, _012222_, _012223_, _012224_, _012225_, _012226_, _012227_, _012228_, _012229_, _012230_, _012231_, _012232_, _012233_, _012234_, _012235_, _012236_, _012237_, _012238_, _012239_, _012240_, _012241_, _012242_, _012243_, _012244_, _012245_, _012246_, _012247_, _012248_, _012249_, _012250_, _012251_, _012252_, _012253_, _012254_, _012255_, _012256_, _012257_, _012258_, _012259_, _012260_, _012261_, _012262_, _012263_, _012264_, _012265_, _012266_, _012267_, _012268_, _012269_, _012270_, _012271_, _012272_, _012273_, _012274_, _012275_, _012276_, _012277_, _012278_, _012279_, _012280_, _012281_, _012282_, _012283_, _012284_, _012285_, _012286_, _012287_, _012288_, _012289_, _012290_, _012291_, _012292_, _012293_, _012294_, _012295_, _012296_, _012297_, _012298_, _012299_, _012300_, _012301_, _012302_, _012303_, _012304_, _012305_, _012306_, _012307_, _012308_, _012309_, _012310_, _012311_, _012312_, _012313_, _012314_, _012315_, _012316_, _012317_, _012318_, _012319_, _012320_, _012321_, _012322_, _012323_, _012324_, _012325_, _012326_, _012327_, _012328_, _012329_, _012330_, _012331_, _012332_, _012333_, _012334_, _012335_, _012336_, _012337_, _012338_, _012339_, _012340_, _012341_, _012342_, _012343_, _012344_, _012345_, _012346_, _012347_, _012348_, _012349_, _012350_, _012351_, _012352_, _012353_, _012354_, _012355_, _012356_, _012357_, _012358_, _012359_, _012360_, _012361_, _012362_, _012363_, _012364_, _012365_, _012366_, _012367_, _012368_, _012369_, _012370_, _012371_, _012372_, _012373_, _012374_, _012375_, _012376_, _012377_, _012378_, _012379_, _012380_, _012381_, _012382_, _012383_, _012384_, _012385_, _012386_, _012387_, _012388_, _012389_, _012390_, _012391_, _012392_, _012393_, _012394_, _012395_, _012396_, _012397_, _012398_, _012399_, _012400_, _012401_, _012402_, _012403_, _012404_, _012405_, _012406_, _012407_, _012408_, _012409_, _012410_, _012411_, _012412_, _012413_, _012414_, _012415_, _012416_, _012417_, _012418_, _012419_, _012420_, _012421_, _012422_, _012423_, _012424_, _012425_, _012426_, _012427_, _012428_, _012429_, _012430_, _012431_, _012432_, _012433_, _012434_, _012435_, _012436_, _012437_, _012438_, _012439_, _012440_, _012441_, _012442_, _012443_, _012444_, _012445_, _012446_, _012447_, _012448_, _012449_, _012450_, _012451_, _012452_, _012453_, _012454_, _012455_, _012456_, _012457_, _012458_, _012459_, _012460_, _012461_, _012462_, _012463_, _012464_, _012465_, _012466_, _012467_, _012468_, _012469_, _012470_, _012471_, _012472_, _012473_, _012474_, _012475_, _012476_, _012477_, _012478_, _012479_, _012480_, _012481_, _012482_, _012483_, _012484_, _012485_, _012486_, _012487_, _012488_, _012489_, _012490_, _012491_, _012492_, _012493_, _012494_, _012495_, _012496_, _012497_, _012498_, _012499_, _012500_, _012501_, _012502_, _012503_, _012504_, _012505_, _012506_, _012507_, _012508_, _012509_, _012510_, _012511_, _012512_, _012513_, _012514_, _012515_, _012516_, _012517_, _012518_, _012519_, _012520_, _012521_, _012522_, _012523_, _012524_, _012525_, _012526_, _012527_, _012528_, _012529_, _012530_, _012531_, _012532_, _012533_, _012534_, _012535_, _012536_, _012537_, _012538_, _012539_, _012540_, _012541_, _012542_, _012543_, _012544_, _012545_, _012546_, _012547_, _012548_, _012549_, _012550_, _012551_, _012552_, _012553_, _012554_, _012555_, _012556_, _012557_, _012558_, _012559_, _012560_, _012561_, _012562_, _012563_, _012564_, _012565_, _012566_, _012567_, _012568_, _012569_, _012570_, _012571_, _012572_, _012573_, _012574_, _012575_, _012576_, _012577_, _012578_, _012579_, _012580_, _012581_, _012582_, _012583_, _012584_, _012585_, _012586_, _012587_, _012588_, _012589_, _012590_, _012591_, _012592_, _012593_, _012594_, _012595_, _012596_, _012597_, _012598_, _012599_, _012600_, _012601_, _012602_, _012603_, _012604_, _012605_, _012606_, _012607_, _012608_, _012609_, _012610_, _012611_, _012612_, _012613_, _012614_, _012615_, _012616_, _012617_, _012618_, _012619_, _012620_, _012621_, _012622_, _012623_, _012624_, _012625_, _012626_, _012627_, _012628_, _012629_, _012630_, _012631_, _012632_, _012633_, _012634_, _012635_, _012636_, _012637_, _012638_, _012639_, _012640_, _012641_, _012642_, _012643_, _012644_, _012645_, _012646_, _012647_, _012648_, _012649_, _012650_, _012651_, _012652_, _012653_, _012654_, _012655_, _012656_, _012657_, _012658_, _012659_, _012660_, _012661_, _012662_, _012663_, _012664_, _012665_, _012666_, _012667_, _012668_, _012669_, _012670_, _012671_, _012672_, _012673_, _012674_, _012675_, _012676_, _012677_, _012678_, _012679_, _012680_, _012681_, _012682_, _012683_, _012684_, _012685_, _012686_, _012687_, _012688_, _012689_, _012690_, _012691_, _012692_, _012693_, _012694_, _012695_, _012696_, _012697_, _012698_, _012699_, _012700_, _012701_, _012702_, _012703_, _012704_, _012705_, _012706_, _012707_, _012708_, _012709_, _012710_, _012711_, _012712_, _012713_, _012714_, _012715_, _012716_, _012717_, _012718_, _012719_, _012720_, _012721_, _012722_, _012723_, _012724_, _012725_, _012726_, _012727_, _012728_, _012729_, _012730_, _012731_, _012732_, _012733_, _012734_, _012735_, _012736_, _012737_, _012738_, _012739_, _012740_, _012741_, _012742_, _012743_, _012744_, _012745_, _012746_, _012747_, _012748_, _012749_, _012750_, _012751_, _012752_, _012753_, _012754_, _012755_, _012756_, _012757_, _012758_, _012759_, _012760_, _012761_, _012762_, _012763_, _012764_, _012765_, _012766_, _012767_, _012768_, _012769_, _012770_, _012771_, _012772_, _012773_, _012774_, _012775_, _012776_, _012777_, _012778_, _012779_, _012780_, _012781_, _012782_, _012783_, _012784_, _012785_, _012786_, _012787_, _012788_, _012789_, _012790_, _012791_, _012792_, _012793_, _012794_, _012795_, _012796_, _012797_, _012798_, _012799_, _012800_, _012801_, _012802_, _012803_, _012804_, _012805_, _012806_, _012807_, _012808_, _012809_, _012810_, _012811_, _012812_, _012813_, _012814_, _012815_, _012816_, _012817_, _012818_, _012819_, _012820_, _012821_, _012822_, _012823_, _012824_, _012825_, _012826_, _012827_, _012828_, _012829_, _012830_, _012831_, _012832_, _012833_, _012834_, _012835_, _012836_, _012837_, _012838_, _012839_, _012840_, _012841_, _012842_, _012843_, _012844_, _012845_, _012846_, _012847_, _012848_, _012849_, _012850_, _012851_, _012852_, _012853_, _012854_, _012855_, _012856_, _012857_, _012858_, _012859_, _012860_, _012861_, _012862_, _012863_, _012864_, _012865_, _012866_, _012867_, _012868_, _012869_, _012870_, _012871_, _012872_, _012873_, _012874_, _012875_, _012876_, _012877_, _012878_, _012879_, _012880_, _012881_, _012882_, _012883_, _012884_, _012885_, _012886_, _012887_, _012888_, _012889_, _012890_, _012891_, _012892_, _012893_, _012894_, _012895_, _012896_, _012897_, _012898_, _012899_, _012900_, _012901_, _012902_, _012903_, _012904_, _012905_, _012906_, _012907_, _012908_, _012909_, _012910_, _012911_, _012912_, _012913_, _012914_, _012915_, _012916_, _012917_, _012918_, _012919_, _012920_, _012921_, _012922_, _012923_, _012924_, _012925_, _012926_, _012927_, _012928_, _012929_, _012930_, _012931_, _012932_, _012933_, _012934_, _012935_, _012936_, _012937_, _012938_, _012939_, _012940_, _012941_, _012942_, _012943_, _012944_, _012945_, _012946_, _012947_, _012948_, _012949_, _012950_, _012951_, _012952_, _012953_, _012954_, _012955_, _012956_, _012957_, _012958_, _012959_, _012960_, _012961_, _012962_, _012963_, _012964_, _012965_, _012966_, _012967_, _012968_, _012969_, _012970_, _012971_, _012972_, _012973_, _012974_, _012975_, _012976_, _012977_, _012978_, _012979_, _012980_, _012981_, _012982_, _012983_, _012984_, _012985_, _012986_, _012987_, _012988_, _012989_, _012990_, _012991_, _012992_, _012993_, _012994_, _012995_, _012996_, _012997_, _012998_, _012999_, _013000_, _013001_, _013002_, _013003_, _013004_, _013005_, _013006_, _013007_, _013008_, _013009_, _013010_, _013011_, _013012_, _013013_, _013014_, _013015_, _013016_, _013017_, _013018_, _013019_, _013020_, _013021_, _013022_, _013023_, _013024_, _013025_, _013026_, _013027_, _013028_, _013029_, _013030_, _013031_, _013032_, _013033_, _013034_, _013035_, _013036_, _013037_, _013038_, _013039_, _013040_, _013041_, _013042_, _013043_, _013044_, _013045_, _013046_, _013047_, _013048_, _013049_, _013050_, _013051_, _013052_, _013053_, _013054_, _013055_, _013056_, _013057_, _013058_, _013059_, _013060_, _013061_, _013062_, _013063_, _013064_, _013065_, _013066_, _013067_, _013068_, _013069_, _013070_, _013071_, _013072_, _013073_, _013074_, _013075_, _013076_, _013077_, _013078_, _013079_, _013080_, _013081_, _013082_, _013083_, _013084_, _013085_, _013086_, _013087_, _013088_, _013089_, _013090_, _013091_, _013092_, _013093_, _013094_, _013095_, _013096_, _013097_, _013098_, _013099_, _013100_, _013101_, _013102_, _013103_, _013104_, _013105_, _013106_, _013107_, _013108_, _013109_, _013110_, _013111_, _013112_, _013113_, _013114_, _013115_, _013116_, _013117_, _013118_, _013119_, _013120_, _013121_, _013122_, _013123_, _013124_, _013125_, _013126_, _013127_, _013128_, _013129_, _013130_, _013131_, _013132_, _013133_, _013134_, _013135_, _013136_, _013137_, _013138_, _013139_, _013140_, _013141_, _013142_, _013143_, _013144_, _013145_, _013146_, _013147_, _013148_, _013149_, _013150_, _013151_, _013152_, _013153_, _013154_, _013155_, _013156_, _013157_, _013158_, _013159_, _013160_, _013161_, _013162_, _013163_, _013164_, _013165_, _013166_, _013167_, _013168_, _013169_, _013170_, _013171_, _013172_, _013173_, _013174_, _013175_, _013176_, _013177_, _013178_, _013179_, _013180_, _013181_, _013182_, _013183_, _013184_, _013185_, _013186_, _013187_, _013188_, _013189_, _013190_, _013191_, _013192_, _013193_, _013194_, _013195_, _013196_, _013197_, _013198_, _013199_, _013200_, _013201_, _013202_, _013203_, _013204_, _013205_, _013206_, _013207_, _013208_, _013209_, _013210_, _013211_, _013212_, _013213_, _013214_, _013215_, _013216_, _013217_, _013218_, _013219_, _013220_, _013221_, _013222_, _013223_, _013224_, _013225_, _013226_, _013227_, _013228_, _013229_, _013230_, _013231_, _013232_, _013233_, _013234_, _013235_, _013236_, _013237_, _013238_, _013239_, _013240_, _013241_, _013242_, _013243_, _013244_, _013245_, _013246_, _013247_, _013248_, _013249_, _013250_, _013251_, _013252_, _013253_, _013254_, _013255_, _013256_, _013257_, _013258_, _013259_, _013260_, _013261_, _013262_, _013263_, _013264_, _013265_, _013266_, _013267_, _013268_, _013269_, _013270_, _013271_, _013272_, _013273_, _013274_, _013275_, _013276_, _013277_, _013278_, _013279_, _013280_, _013281_, _013282_, _013283_, _013284_, _013285_, _013286_, _013287_, _013288_, _013289_, _013290_, _013291_, _013292_, _013293_, _013294_, _013295_, _013296_, _013297_, _013298_, _013299_, _013300_, _013301_, _013302_, _013303_, _013304_, _013305_, _013306_, _013307_, _013308_, _013309_, _013310_, _013311_, _013312_, _013313_, _013314_, _013315_, _013316_, _013317_, _013318_, _013319_, _013320_, _013321_, _013322_, _013323_, _013324_, _013325_, _013326_, _013327_, _013328_, _013329_, _013330_, _013331_, _013332_, _013333_, _013334_, _013335_, _013336_, _013337_, _013338_, _013339_, _013340_, _013341_, _013342_, _013343_, _013344_, _013345_, _013346_, _013347_, _013348_, _013349_, _013350_, _013351_, _013352_, _013353_, _013354_, _013355_, _013356_, _013357_, _013358_, _013359_, _013360_, _013361_, _013362_, _013363_, _013364_, _013365_, _013366_, _013367_, _013368_, _013369_, _013370_, _013371_, _013372_, _013373_, _013374_, _013375_, _013376_, _013377_, _013378_, _013379_, _013380_, _013381_, _013382_, _013383_, _013384_, _013385_, _013386_, _013387_, _013388_, _013389_, _013390_, _013391_, _013392_, _013393_, _013394_, _013395_, _013396_, _013397_, _013398_, _013399_, _013400_, _013401_, _013402_, _013403_, _013404_, _013405_, _013406_, _013407_, _013408_, _013409_, _013410_, _013411_, _013412_, _013413_, _013414_, _013415_, _013416_, _013417_, _013418_, _013419_, _013420_, _013421_, _013422_, _013423_, _013424_, _013425_, _013426_, _013427_, _013428_, _013429_, _013430_, _013431_, _013432_, _013433_, _013434_, _013435_, _013436_, _013437_, _013438_, _013439_, _013440_, _013441_, _013442_, _013443_, _013444_, _013445_, _013446_, _013447_, _013448_, _013449_, _013450_, _013451_, _013452_, _013453_, _013454_, _013455_, _013456_, _013457_, _013458_, _013459_, _013460_, _013461_, _013462_, _013463_, _013464_, _013465_, _013466_, _013467_, _013468_, _013469_, _013470_, _013471_, _013472_, _013473_, _013474_, _013475_, _013476_, _013477_, _013478_, _013479_, _013480_, _013481_, _013482_, _013483_, _013484_, _013485_, _013486_, _013487_, _013488_, _013489_, _013490_, _013491_, _013492_, _013493_, _013494_, _013495_, _013496_, _013497_, _013498_, _013499_, _013500_, _013501_, _013502_, _013503_, _013504_, _013505_, _013506_, _013507_, _013508_, _013509_, _013510_, _013511_, _013512_, _013513_, _013514_, _013515_, _013516_, _013517_, _013518_, _013519_, _013520_, _013521_, _013522_, _013523_, _013524_, _013525_, _013526_, _013527_, _013528_, _013529_, _013530_, _013531_, _013532_, _013533_, _013534_, _013535_, _013536_, _013537_, _013538_, _013539_, _013540_, _013541_, _013542_, _013543_, _013544_, _013545_, _013546_, _013547_, _013548_, _013549_, _013550_, _013551_, _013552_, _013553_, _013554_, _013555_, _013556_, _013557_, _013558_, _013559_, _013560_, _013561_, _013562_, _013563_, _013564_, _013565_, _013566_, _013567_, _013568_, _013569_, _013570_, _013571_, _013572_, _013573_, _013574_, _013575_, _013576_, _013577_, _013578_, _013579_, _013580_, _013581_, _013582_, _013583_, _013584_, _013585_, _013586_, _013587_, _013588_, _013589_, _013590_, _013591_, _013592_, _013593_, _013594_, _013595_, _013596_, _013597_, _013598_, _013599_, _013600_, _013601_, _013602_, _013603_, _013604_, _013605_, _013606_, _013607_, _013608_, _013609_, _013610_, _013611_, _013612_, _013613_, _013614_, _013615_, _013616_, _013617_, _013618_, _013619_, _013620_, _013621_, _013622_, _013623_, _013624_, _013625_, _013626_, _013627_, _013628_, _013629_, _013630_, _013631_, _013632_, _013633_, _013634_, _013635_, _013636_, _013637_, _013638_, _013639_, _013640_, _013641_, _013642_, _013643_, _013644_, _013645_, _013646_, _013647_, _013648_, _013649_, _013650_, _013651_, _013652_, _013653_, _013654_, _013655_, _013656_, _013657_, _013658_, _013659_, _013660_, _013661_, _013662_, _013663_, _013664_, _013665_, _013666_, _013667_, _013668_, _013669_, _013670_, _013671_, _013672_, _013673_, _013674_, _013675_, _013676_, _013677_, _013678_, _013679_, _013680_, _013681_, _013682_, _013683_, _013684_, _013685_, _013686_, _013687_, _013688_, _013689_, _013690_, _013691_, _013692_, _013693_, _013694_, _013695_, _013696_, _013697_, _013698_, _013699_, _013700_, _013701_, _013702_, _013703_, _013704_, _013705_, _013706_, _013707_, _013708_, _013709_, _013710_, _013711_, _013712_, _013713_, _013714_, _013715_, _013716_, _013717_, _013718_, _013719_, _013720_, _013721_, _013722_, _013723_, _013724_, _013725_, _013726_, _013727_, _013728_, _013729_, _013730_, _013731_, _013732_, _013733_, _013734_, _013735_, _013736_, _013737_, _013738_, _013739_, _013740_, _013741_, _013742_, _013743_, _013744_, _013745_, _013746_, _013747_, _013748_, _013749_, _013750_, _013751_, _013752_, _013753_, _013754_, _013755_, _013756_, _013757_, _013758_, _013759_, _013760_, _013761_, _013762_, _013763_, _013764_, _013765_, _013766_, _013767_, _013768_, _013769_, _013770_, _013771_, _013772_, _013773_, _013774_, _013775_, _013776_, _013777_, _013778_, _013779_, _013780_, _013781_, _013782_, _013783_, _013784_, _013785_, _013786_, _013787_, _013788_, _013789_, _013790_, _013791_, _013792_, _013793_, _013794_, _013795_, _013796_, _013797_, _013798_, _013799_, _013800_, _013801_, _013802_, _013803_, _013804_, _013805_, _013806_, _013807_, _013808_, _013809_, _013810_, _013811_, _013812_, _013813_, _013814_, _013815_, _013816_, _013817_, _013818_, _013819_, _013820_, _013821_, _013822_, _013823_, _013824_, _013825_, _013826_, _013827_, _013828_, _013829_, _013830_, _013831_, _013832_, _013833_, _013834_, _013835_, _013836_, _013837_, _013838_, _013839_, _013840_, _013841_, _013842_, _013843_, _013844_, _013845_, _013846_, _013847_, _013848_, _013849_, _013850_, _013851_, _013852_, _013853_, _013854_, _013855_, _013856_, _013857_, _013858_, _013859_, _013860_, _013861_, _013862_, _013863_, _013864_, _013865_, _013866_, _013867_, _013868_, _013869_, _013870_, _013871_, _013872_, _013873_, _013874_, _013875_, _013876_, _013877_, _013878_, _013879_, _013880_, _013881_, _013882_, _013883_, _013884_, _013885_, _013886_, _013887_, _013888_, _013889_, _013890_, _013891_, _013892_, _013893_, _013894_, _013895_, _013896_, _013897_, _013898_, _013899_, _013900_, _013901_, _013902_, _013903_, _013904_, _013905_, _013906_, _013907_, _013908_, _013909_, _013910_, _013911_, _013912_, _013913_, _013914_, _013915_, _013916_, _013917_, _013918_, _013919_, _013920_, _013921_, _013922_, _013923_, _013924_, _013925_, _013926_, _013927_, _013928_, _013929_, _013930_, _013931_, _013932_, _013933_, _013934_, _013935_, _013936_, _013937_, _013938_, _013939_, _013940_, _013941_, _013942_, _013943_, _013944_, _013945_, _013946_, _013947_, _013948_, _013949_, _013950_, _013951_, _013952_, _013953_, _013954_, _013955_, _013956_, _013957_, _013958_, _013959_, _013960_, _013961_, _013962_, _013963_, _013964_, _013965_, _013966_, _013967_, _013968_, _013969_, _013970_, _013971_, _013972_, _013973_, _013974_, _013975_, _013976_, _013977_, _013978_, _013979_, _013980_, _013981_, _013982_, _013983_, _013984_, _013985_, _013986_, _013987_, _013988_, _013989_, _013990_, _013991_, _013992_, _013993_, _013994_, _013995_, _013996_, _013997_, _013998_, _013999_, _014000_, _014001_, _014002_, _014003_, _014004_, _014005_, _014006_, _014007_, _014008_, _014009_, _014010_, _014011_, _014012_, _014013_, _014014_, _014015_, _014016_, _014017_, _014018_, _014019_, _014020_, _014021_, _014022_, _014023_, _014024_, _014025_, _014026_, _014027_, _014028_, _014029_, _014030_, _014031_, _014032_, _014033_, _014034_, _014035_, _014036_, _014037_, _014038_, _014039_, _014040_, _014041_, _014042_, _014043_, _014044_, _014045_, _014046_, _014047_, _014048_, _014049_, _014050_, _014051_, _014052_, _014053_, _014054_, _014055_, _014056_, _014057_, _014058_, _014059_, _014060_, _014061_, _014062_, _014063_, _014064_, _014065_, _014066_, _014067_, _014068_, _014069_, _014070_, _014071_, _014072_, _014073_, _014074_, _014075_, _014076_, _014077_, _014078_, _014079_, _014080_, _014081_, _014082_, _014083_, _014084_, _014085_, _014086_, _014087_, _014088_, _014089_, _014090_, _014091_, _014092_, _014093_, _014094_, _014095_, _014096_, _014097_, _014098_, _014099_, _014100_, _014101_, _014102_, _014103_, _014104_, _014105_, _014106_, _014107_, _014108_, _014109_, _014110_, _014111_, _014112_, _014113_, _014114_, _014115_, _014116_, _014117_, _014118_, _014119_, _014120_, _014121_, _014122_, _014123_, _014124_, _014125_, _014126_, _014127_, _014128_, _014129_, _014130_, _014131_, _014132_, _014133_, _014134_, _014135_, _014136_, _014137_, _014138_, _014139_, _014140_, _014141_, _014142_, _014143_, _014144_, _014145_, _014146_, _014147_, _014148_, _014149_, _014150_, _014151_, _014152_, _014153_, _014154_, _014155_, _014156_, _014157_, _014158_, _014159_, _014160_, _014161_, _014162_, _014163_, _014164_, _014165_, _014166_, _014167_, _014168_, _014169_, _014170_, _014171_, _014172_, _014173_, _014174_, _014175_, _014176_, _014177_, _014178_, _014179_, _014180_, _014181_, _014182_, _014183_, _014184_, _014185_, _014186_, _014187_, _014188_, _014189_, _014190_, _014191_, _014192_, _014193_, _014194_, _014195_, _014196_, _014197_, _014198_, _014199_, _014200_, _014201_, _014202_, _014203_, _014204_, _014205_, _014206_, _014207_, _014208_, _014209_, _014210_, _014211_, _014212_, _014213_, _014214_, _014215_, _014216_, _014217_, _014218_, _014219_, _014220_, _014221_, _014222_, _014223_, _014224_, _014225_, _014226_, _014227_, _014228_, _014229_, _014230_, _014231_, _014232_, _014233_, _014234_, _014235_, _014236_, _014237_, _014238_, _014239_, _014240_, _014241_, _014242_, _014243_, _014244_, _014245_, _014246_, _014247_, _014248_, _014249_, _014250_, _014251_, _014252_, _014253_, _014254_, _014255_, _014256_, _014257_, _014258_, _014259_, _014260_, _014261_, _014262_, _014263_, _014264_, _014265_, _014266_, _014267_, _014268_, _014269_, _014270_, _014271_, _014272_, _014273_, _014274_, _014275_, _014276_, _014277_, _014278_, _014279_, _014280_, _014281_, _014282_, _014283_, _014284_, _014285_, _014286_, _014287_, _014288_, _014289_, _014290_, _014291_, _014292_, _014293_, _014294_, _014295_, _014296_, _014297_, _014298_, _014299_, _014300_, _014301_, _014302_, _014303_, _014304_, _014305_, _014306_, _014307_, _014308_, _014309_, _014310_, _014311_, _014312_, _014313_, _014314_, _014315_, _014316_, _014317_, _014318_, _014319_, _014320_, _014321_, _014322_, _014323_, _014324_, _014325_, _014326_, _014327_, _014328_, _014329_, _014330_, _014331_, _014332_, _014333_, _014334_, _014335_, _014336_, _014337_, _014338_, _014339_, _014340_, _014341_, _014342_, _014343_, _014344_, _014345_, _014346_, _014347_, _014348_, _014349_, _014350_, _014351_, _014352_, _014353_, _014354_, _014355_, _014356_, _014357_, _014358_, _014359_, _014360_, _014361_, _014362_, _014363_, _014364_, _014365_, _014366_, _014367_, _014368_, _014369_, _014370_, _014371_, _014372_, _014373_, _014374_, _014375_, _014376_, _014377_, _014378_, _014379_, _014380_, _014381_, _014382_, _014383_, _014384_, _014385_, _014386_, _014387_, _014388_, _014389_, _014390_, _014391_, _014392_, _014393_, _014394_, _014395_, _014396_, _014397_, _014398_, _014399_, _014400_, _014401_, _014402_, _014403_, _014404_, _014405_, _014406_, _014407_, _014408_, _014409_, _014410_, _014411_, _014412_, _014413_, _014414_, _014415_, _014416_, _014417_, _014418_, _014419_, _014420_, _014421_, _014422_, _014423_, _014424_, _014425_, _014426_, _014427_, _014428_, _014429_, _014430_, _014431_, _014432_, _014433_, _014434_, _014435_, _014436_, _014437_, _014438_, _014439_, _014440_, _014441_, _014442_, _014443_, _014444_, _014445_, _014446_, _014447_, _014448_, _014449_, _014450_, _014451_, _014452_, _014453_, _014454_, _014455_, _014456_, _014457_, _014458_, _014459_, _014460_, _014461_, _014462_, _014463_, _014464_, _014465_, _014466_, _014467_, _014468_, _014469_, _014470_, _014471_, _014472_, _014473_, _014474_, _014475_, _014476_, _014477_, _014478_, _014479_, _014480_, _014481_, _014482_, _014483_, _014484_, _014485_, _014486_, _014487_, _014488_, _014489_, _014490_, _014491_, _014492_, _014493_, _014494_, _014495_, _014496_, _014497_, _014498_, _014499_, _014500_, _014501_, _014502_, _014503_, _014504_, _014505_, _014506_, _014507_, _014508_, _014509_, _014510_, _014511_, _014512_, _014513_, _014514_, _014515_, _014516_, _014517_, _014518_, _014519_, _014520_, _014521_, _014522_, _014523_, _014524_, _014525_, _014526_, _014527_, _014528_, _014529_, _014530_, _014531_, _014532_, _014533_, _014534_, _014535_, _014536_, _014537_, _014538_, _014539_, _014540_, _014541_, _014542_, _014543_, _014544_, _014545_, _014546_, _014547_, _014548_, _014549_, _014550_, _014551_, _014552_, _014553_, _014554_, _014555_, _014556_, _014557_, _014558_, _014559_, _014560_, _014561_, _014562_, _014563_, _014564_, _014565_, _014566_, _014567_, _014568_, _014569_, _014570_, _014571_, _014572_, _014573_, _014574_, _014575_, _014576_, _014577_, _014578_, _014579_, _014580_, _014581_, _014582_, _014583_, _014584_, _014585_, _014586_, _014587_, _014588_, _014589_, _014590_, _014591_, _014592_, _014593_, _014594_, _014595_, _014596_, _014597_, _014598_, _014599_, _014600_, _014601_, _014602_, _014603_, _014604_, _014605_, _014606_, _014607_, _014608_, _014609_, _014610_, _014611_, _014612_, _014613_, _014614_, _014615_, _014616_, _014617_, _014618_, _014619_, _014620_, _014621_, _014622_, _014623_, _014624_, _014625_, _014626_, _014627_, _014628_, _014629_, _014630_, _014631_, _014632_, _014633_, _014634_, _014635_, _014636_, _014637_, _014638_, _014639_, _014640_, _014641_, _014642_, _014643_, _014644_, _014645_, _014646_, _014647_, _014648_, _014649_, _014650_, _014651_, _014652_, _014653_, _014654_, _014655_, _014656_, _014657_, _014658_, _014659_, _014660_, _014661_, _014662_, _014663_, _014664_, _014665_, _014666_, _014667_, _014668_, _014669_, _014670_, _014671_, _014672_, _014673_, _014674_, _014675_, _014676_, _014677_, _014678_, _014679_, _014680_, _014681_, _014682_, _014683_, _014684_, _014685_, _014686_, _014687_, _014688_, _014689_, _014690_, _014691_, _014692_, _014693_, _014694_, _014695_, _014696_, _014697_, _014698_, _014699_, _014700_, _014701_, _014702_, _014703_, _014704_, _014705_, _014706_, _014707_, _014708_, _014709_, _014710_, _014711_, _014712_, _014713_, _014714_, _014715_, _014716_, _014717_, _014718_, _014719_, _014720_, _014721_, _014722_, _014723_, _014724_, _014725_, _014726_, _014727_, _014728_, _014729_, _014730_, _014731_, _014732_, _014733_, _014734_, _014735_, _014736_, _014737_, _014738_, _014739_, _014740_, _014741_, _014742_, _014743_, _014744_, _014745_, _014746_, _014747_, _014748_, _014749_, _014750_, _014751_, _014752_, _014753_, _014754_, _014755_, _014756_, _014757_, _014758_, _014759_, _014760_, _014761_, _014762_, _014763_, _014764_, _014765_, _014766_, _014767_, _014768_, _014769_, _014770_, _014771_, _014772_, _014773_, _014774_, _014775_, _014776_, _014777_, _014778_, _014779_, _014780_, _014781_, _014782_, _014783_, _014784_, _014785_, _014786_, _014787_, _014788_, _014789_, _014790_, _014791_, _014792_, _014793_, _014794_, _014795_, _014796_, _014797_, _014798_, _014799_, _014800_, _014801_, _014802_, _014803_, _014804_, _014805_, _014806_, _014807_, _014808_, _014809_, _014810_, _014811_, _014812_, _014813_, _014814_, _014815_, _014816_, _014817_, _014818_, _014819_, _014820_, _014821_, _014822_, _014823_, _014824_, _014825_, _014826_, _014827_, _014828_, _014829_, _014830_, _014831_, _014832_, _014833_, _014834_, _014835_, _014836_, _014837_, _014838_, _014839_, _014840_, _014841_, _014842_, _014843_, _014844_, _014845_, _014846_, _014847_, _014848_, _014849_, _014850_, _014851_, _014852_, _014853_, _014854_, _014855_, _014856_, _014857_, _014858_, _014859_, _014860_, _014861_, _014862_, _014863_, _014864_, _014865_, _014866_, _014867_, _014868_, _014869_, _014870_, _014871_, _014872_, _014873_, _014874_, _014875_, _014876_, _014877_, _014878_, _014879_, _014880_, _014881_, _014882_, _014883_, _014884_, _014885_, _014886_, _014887_, _014888_, _014889_, _014890_, _014891_, _014892_, _014893_, _014894_, _014895_, _014896_, _014897_, _014898_, _014899_, _014900_, _014901_, _014902_, _014903_, _014904_, _014905_, _014906_, _014907_, _014908_, _014909_, _014910_, _014911_, _014912_, _014913_, _014914_, _014915_, _014916_, _014917_, _014918_, _014919_, _014920_, _014921_, _014922_, _014923_, _014924_, _014925_, _014926_, _014927_, _014928_, _014929_, _014930_, _014931_, _014932_, _014933_, _014934_, _014935_, _014936_, _014937_, _014938_, _014939_, _014940_, _014941_, _014942_, _014943_, _014944_, _014945_, _014946_, _014947_, _014948_, _014949_, _014950_, _014951_, _014952_, _014953_, _014954_, _014955_, _014956_, _014957_, _014958_, _014959_, _014960_, _014961_, _014962_, _014963_, _014964_, _014965_, _014966_, _014967_, _014968_, _014969_, _014970_, _014971_, _014972_, _014973_, _014974_, _014975_, _014976_, _014977_, _014978_, _014979_, _014980_, _014981_, _014982_, _014983_, _014984_, _014985_, _014986_, _014987_, _014988_, _014989_, _014990_, _014991_, _014992_, _014993_, _014994_, _014995_, _014996_, _014997_, _014998_, _014999_, _015000_, _015001_, _015002_, _015003_, _015004_, _015005_, _015006_, _015007_, _015008_, _015009_, _015010_, _015011_, _015012_, _015013_, _015014_, _015015_, _015016_, _015017_, _015018_, _015019_, _015020_, _015021_, _015022_, _015023_, _015024_, _015025_, _015026_, _015027_, _015028_, _015029_, _015030_, _015031_, _015032_, _015033_, _015034_, _015035_, _015036_, _015037_, _015038_, _015039_, _015040_, _015041_, _015042_, _015043_, _015044_, _015045_, _015046_, _015047_, _015048_, _015049_, _015050_, _015051_, _015052_, _015053_, _015054_, _015055_, _015056_, _015057_, _015058_, _015059_, _015060_, _015061_, _015062_, _015063_, _015064_, _015065_, _015066_, _015067_, _015068_, _015069_, _015070_, _015071_, _015072_, _015073_, _015074_, _015075_, _015076_, _015077_, _015078_, _015079_, _015080_, _015081_, _015082_, _015083_, _015084_, _015085_, _015086_, _015087_, _015088_, _015089_, _015090_, _015091_, _015092_, _015093_, _015094_, _015095_, _015096_, _015097_, _015098_, _015099_, _015100_, _015101_, _015102_, _015103_, _015104_, _015105_, _015106_, _015107_, _015108_, _015109_, _015110_, _015111_, _015112_, _015113_, _015114_, _015115_, _015116_, _015117_, _015118_, _015119_, _015120_, _015121_, _015122_, _015123_, _015124_, _015125_, _015126_, _015127_, _015128_, _015129_, _015130_, _015131_, _015132_, _015133_, _015134_, _015135_, _015136_, _015137_, _015138_, _015139_, _015140_, _015141_, _015142_, _015143_, _015144_, _015145_, _015146_, _015147_, _015148_, _015149_, _015150_, _015151_, _015152_, _015153_, _015154_, _015155_, _015156_, _015157_, _015158_, _015159_, _015160_, _015161_, _015162_, _015163_, _015164_, _015165_, _015166_, _015167_, _015168_, _015169_, _015170_, _015171_, _015172_, _015173_, _015174_, _015175_, _015176_, _015177_, _015178_, _015179_, _015180_, _015181_, _015182_, _015183_, _015184_, _015185_, _015186_, _015187_, _015188_, _015189_, _015190_, _015191_, _015192_, _015193_, _015194_, _015195_, _015196_, _015197_, _015198_, _015199_, _015200_, _015201_, _015202_, _015203_, _015204_, _015205_, _015206_, _015207_, _015208_, _015209_, _015210_, _015211_, _015212_, _015213_, _015214_, _015215_, _015216_, _015217_, _015218_, _015219_, _015220_, _015221_, _015222_, _015223_, _015224_, _015225_, _015226_, _015227_, _015228_, _015229_, _015230_, _015231_, _015232_, _015233_, _015234_, _015235_, _015236_, _015237_, _015238_, _015239_, _015240_, _015241_, _015242_, _015243_, _015244_, _015245_, _015246_, _015247_, _015248_, _015249_, _015250_, _015251_, _015252_, _015253_, _015254_, _015255_, _015256_, _015257_, _015258_, _015259_, _015260_, _015261_, _015262_, _015263_, _015264_, _015265_, _015266_, _015267_, _015268_, _015269_, _015270_, _015271_, _015272_, _015273_, _015274_, _015275_, _015276_, _015277_, _015278_, _015279_, _015280_, _015281_, _015282_, _015283_, _015284_, _015285_, _015286_, _015287_, _015288_, _015289_, _015290_, _015291_, _015292_, _015293_, _015294_, _015295_, _015296_, _015297_, _015298_, _015299_, _015300_, _015301_, _015302_, _015303_, _015304_, _015305_, _015306_, _015307_, _015308_, _015309_, _015310_, _015311_, _015312_, _015313_, _015314_, _015315_, _015316_, _015317_, _015318_, _015319_, _015320_, _015321_, _015322_, _015323_, _015324_, _015325_, _015326_, _015327_, _015328_, _015329_, _015330_, _015331_, _015332_, _015333_, _015334_, _015335_, _015336_, _015337_, _015338_, _015339_, _015340_, _015341_, _015342_, _015343_, _015344_, _015345_, _015346_, _015347_, _015348_, _015349_, _015350_, _015351_, _015352_, _015353_, _015354_, _015355_, _015356_, _015357_, _015358_, _015359_, _015360_, _015361_, _015362_, _015363_, _015364_, _015365_, _015366_, _015367_, _015368_, _015369_, _015370_, _015371_, _015372_, _015373_, _015374_, _015375_, _015376_, _015377_, _015378_, _015379_, _015380_, _015381_, _015382_, _015383_, _015384_, _015385_, _015386_, _015387_, _015388_, _015389_, _015390_, _015391_, _015392_, _015393_, _015394_, _015395_, _015396_, _015397_, _015398_, _015399_, _015400_, _015401_, _015402_, _015403_, _015404_, _015405_, _015406_, _015407_, _015408_, _015409_, _015410_, _015411_, _015412_, _015413_, _015414_, _015415_, _015416_, _015417_, _015418_, _015419_, _015420_, _015421_, _015422_, _015423_, _015424_, _015425_, _015426_, _015427_, _015428_, _015429_, _015430_, _015431_, _015432_, _015433_, _015434_, _015435_, _015436_, _015437_, _015438_, _015439_, _015440_, _015441_, _015442_, _015443_, _015444_, _015445_, _015446_, _015447_, _015448_, _015449_, _015450_, _015451_, _015452_, _015453_, _015454_, _015455_, _015456_, _015457_, _015458_, _015459_, _015460_, _015461_, _015462_, _015463_, _015464_, _015465_, _015466_, _015467_, _015468_, _015469_, _015470_, _015471_, _015472_, _015473_, _015474_, _015475_, _015476_, _015477_, _015478_, _015479_, _015480_, _015481_, _015482_, _015483_, _015484_, _015485_, _015486_, _015487_, _015488_, _015489_, _015490_, _015491_, _015492_, _015493_, _015494_, _015495_, _015496_, _015497_, _015498_, _015499_, _015500_, _015501_, _015502_, _015503_, _015504_, _015505_, _015506_, _015507_, _015508_, _015509_, _015510_, _015511_, _015512_, _015513_, _015514_, _015515_, _015516_, _015517_, _015518_, _015519_, _015520_, _015521_, _015522_, _015523_, _015524_, _015525_, _015526_, _015527_, _015528_, _015529_, _015530_, _015531_, _015532_, _015533_, _015534_, _015535_, _015536_, _015537_, _015538_, _015539_, _015540_, _015541_, _015542_, _015543_, _015544_, _015545_, _015546_, _015547_, _015548_, _015549_, _015550_, _015551_, _015552_, _015553_, _015554_, _015555_, _015556_, _015557_, _015558_, _015559_, _015560_, _015561_, _015562_, _015563_, _015564_, _015565_, _015566_, _015567_, _015568_, _015569_, _015570_, _015571_, _015572_, _015573_, _015574_, _015575_, _015576_, _015577_, _015578_, _015579_, _015580_, _015581_, _015582_, _015583_, _015584_, _015585_, _015586_, _015587_, _015588_, _015589_, _015590_, _015591_, _015592_, _015593_, _015594_, _015595_, _015596_, _015597_, _015598_, _015599_, _015600_, _015601_, _015602_, _015603_, _015604_, _015605_, _015606_, _015607_, _015608_, _015609_, _015610_, _015611_, _015612_, _015613_, _015614_, _015615_, _015616_, _015617_, _015618_, _015619_, _015620_, _015621_, _015622_, _015623_, _015624_, _015625_, _015626_, _015627_, _015628_, _015629_, _015630_, _015631_, _015632_, _015633_, _015634_, _015635_, _015636_, _015637_, _015638_, _015639_, _015640_, _015641_, _015642_, _015643_, _015644_, _015645_, _015646_, _015647_, _015648_, _015649_, _015650_, _015651_, _015652_, _015653_, _015654_, _015655_, _015656_, _015657_, _015658_, _015659_, _015660_, _015661_, _015662_, _015663_, _015664_, _015665_, _015666_, _015667_, _015668_, _015669_, _015670_, _015671_, _015672_, _015673_, _015674_, _015675_, _015676_, _015677_, _015678_, _015679_, _015680_, _015681_, _015682_, _015683_, _015684_, _015685_, _015686_, _015687_, _015688_, _015689_, _015690_, _015691_, _015692_, _015693_, _015694_, _015695_, _015696_, _015697_, _015698_, _015699_, _015700_, _015701_, _015702_, _015703_, _015704_, _015705_, _015706_, _015707_, _015708_, _015709_, _015710_, _015711_, _015712_, _015713_, _015714_, _015715_, _015716_, _015717_, _015718_, _015719_, _015720_, _015721_, _015722_, _015723_, _015724_, _015725_, _015726_, _015727_, _015728_, _015729_, _015730_, _015731_, _015732_, _015733_, _015734_, _015735_, _015736_, _015737_, _015738_, _015739_, _015740_, _015741_, _015742_, _015743_, _015744_, _015745_, _015746_, _015747_, _015748_, _015749_, _015750_, _015751_, _015752_, _015753_, _015754_, _015755_, _015756_, _015757_, _015758_, _015759_, _015760_, _015761_, _015762_, _015763_, _015764_, _015765_, _015766_, _015767_, _015768_, _015769_, _015770_, _015771_, _015772_, _015773_, _015774_, _015775_, _015776_, _015777_, _015778_, _015779_, _015780_, _015781_, _015782_, _015783_, _015784_, _015785_, _015786_, _015787_, _015788_, _015789_, _015790_, _015791_, _015792_, _015793_, _015794_, _015795_, _015796_, _015797_, _015798_, _015799_, _015800_, _015801_, _015802_, _015803_, _015804_, _015805_, _015806_, _015807_, _015808_, _015809_, _015810_, _015811_, _015812_, _015813_, _015814_, _015815_, _015816_, _015817_, _015818_, _015819_, _015820_, _015821_, _015822_, _015823_, _015824_, _015825_, _015826_, _015827_, _015828_, _015829_, _015830_, _015831_, _015832_, _015833_, _015834_, _015835_, _015836_, _015837_, _015838_, _015839_, _015840_, _015841_, _015842_, _015843_, _015844_, _015845_, _015846_, _015847_, _015848_, _015849_, _015850_, _015851_, _015852_, _015853_, _015854_, _015855_, _015856_, _015857_, _015858_, _015859_, _015860_, _015861_, _015862_, _015863_, _015864_, _015865_, _015866_, _015867_, _015868_, _015869_, _015870_, _015871_, _015872_, _015873_, _015874_, _015875_, _015876_, _015877_, _015878_, _015879_, _015880_, _015881_, _015882_, _015883_, _015884_, _015885_, _015886_, _015887_, _015888_, _015889_, _015890_, _015891_, _015892_, _015893_, _015894_, _015895_, _015896_, _015897_, _015898_, _015899_, _015900_, _015901_, _015902_, _015903_, _015904_, _015905_, _015906_, _015907_, _015908_, _015909_, _015910_, _015911_, _015912_, _015913_, _015914_, _015915_, _015916_, _015917_, _015918_, _015919_, _015920_, _015921_, _015922_, _015923_, _015924_, _015925_, _015926_, _015927_, _015928_, _015929_, _015930_, _015931_, _015932_, _015933_, _015934_, _015935_, _015936_, _015937_, _015938_, _015939_, _015940_, _015941_, _015942_, _015943_, _015944_, _015945_, _015946_, _015947_, _015948_, _015949_, _015950_, _015951_, _015952_, _015953_, _015954_, _015955_, _015956_, _015957_, _015958_, _015959_, _015960_, _015961_, _015962_, _015963_, _015964_, _015965_, _015966_, _015967_, _015968_, _015969_, _015970_, _015971_, _015972_, _015973_, _015974_, _015975_, _015976_, _015977_, _015978_, _015979_, _015980_, _015981_, _015982_, _015983_, _015984_, _015985_, _015986_, _015987_, _015988_, _015989_, _015990_, _015991_, _015992_, _015993_, _015994_, _015995_, _015996_, _015997_, _015998_, _015999_, _016000_, _016001_, _016002_, _016003_, _016004_, _016005_, _016006_, _016007_, _016008_, _016009_, _016010_, _016011_, _016012_, _016013_, _016014_, _016015_, _016016_, _016017_, _016018_, _016019_, _016020_, _016021_, _016022_, _016023_, _016024_, _016025_, _016026_, _016027_, _016028_, _016029_, _016030_, _016031_, _016032_, _016033_, _016034_, _016035_, _016036_, _016037_, _016038_, _016039_, _016040_, _016041_, _016042_, _016043_, _016044_, _016045_, _016046_, _016047_, _016048_, _016049_, _016050_, _016051_, _016052_, _016053_, _016054_, _016055_, _016056_, _016057_, _016058_, _016059_, _016060_, _016061_, _016062_, _016063_, _016064_, _016065_, _016066_, _016067_, _016068_, _016069_, _016070_, _016071_, _016072_, _016073_, _016074_, _016075_, _016076_, _016077_, _016078_, _016079_, _016080_, _016081_, _016082_, _016083_, _016084_, _016085_, _016086_, _016087_, _016088_, _016089_, _016090_, _016091_, _016092_, _016093_, _016094_, _016095_, _016096_, _016097_, _016098_, _016099_, _016100_, _016101_, _016102_, _016103_, _016104_, _016105_, _016106_, _016107_, _016108_, _016109_, _016110_, _016111_, _016112_, _016113_, _016114_, _016115_, _016116_, _016117_, _016118_, _016119_, _016120_, _016121_, _016122_, _016123_, _016124_, _016125_, _016126_, _016127_, _016128_, _016129_, _016130_, _016131_, _016132_, _016133_, _016134_, _016135_, _016136_, _016137_, _016138_, _016139_, _016140_, _016141_, _016142_, _016143_, _016144_, _016145_, _016146_, _016147_, _016148_, _016149_, _016150_, _016151_, _016152_, _016153_, _016154_, _016155_, _016156_, _016157_, _016158_, _016159_, _016160_, _016161_, _016162_, _016163_, _016164_, _016165_, _016166_, _016167_, _016168_, _016169_, _016170_, _016171_, _016172_, _016173_, _016174_, _016175_, _016176_, _016177_, _016178_, _016179_, _016180_, _016181_, _016182_, _016183_, _016184_, _016185_, _016186_, _016187_, _016188_, _016189_, _016190_, _016191_, _016192_, _016193_, _016194_, _016195_, _016196_, _016197_, _016198_, _016199_, _016200_, _016201_, _016202_, _016203_, _016204_, _016205_, _016206_, _016207_, _016208_, _016209_, _016210_, _016211_, _016212_, _016213_, _016214_, _016215_, _016216_, _016217_, _016218_, _016219_, _016220_, _016221_, _016222_, _016223_, _016224_, _016225_, _016226_, _016227_, _016228_, _016229_, _016230_, _016231_, _016232_, _016233_, _016234_, _016235_, _016236_, _016237_, _016238_, _016239_, _016240_, _016241_, _016242_, _016243_, _016244_, _016245_, _016246_, _016247_, _016248_, _016249_, _016250_, _016251_, _016252_, _016253_, _016254_, _016255_, _016256_, _016257_, _016258_, _016259_, _016260_, _016261_, _016262_, _016263_, _016264_, _016265_, _016266_, _016267_, _016268_, _016269_, _016270_, _016271_, _016272_, _016273_, _016274_, _016275_, _016276_, _016277_, _016278_, _016279_, _016280_, _016281_, _016282_, _016283_, _016284_, _016285_, _016286_, _016287_, _016288_, _016289_, _016290_, _016291_, _016292_, _016293_, _016294_, _016295_, _016296_, _016297_, _016298_, _016299_, _016300_, _016301_, _016302_, _016303_, _016304_, _016305_, _016306_, _016307_, _016308_, _016309_, _016310_, _016311_, _016312_, _016313_, _016314_, _016315_, _016316_, _016317_, _016318_, _016319_, _016320_, _016321_, _016322_, _016323_, _016324_, _016325_, _016326_, _016327_, _016328_, _016329_, _016330_, _016331_, _016332_, _016333_, _016334_, _016335_, _016336_, _016337_, _016338_, _016339_, _016340_, _016341_, _016342_, _016343_, _016344_, _016345_, _016346_, _016347_, _016348_, _016349_, _016350_, _016351_, _016352_, _016353_, _016354_, _016355_, _016356_, _016357_, _016358_, _016359_, _016360_, _016361_, _016362_, _016363_, _016364_, _016365_, _016366_, _016367_, _016368_, _016369_, _016370_, _016371_, _016372_, _016373_, _016374_, _016375_, _016376_, _016377_, _016378_, _016379_, _016380_, _016381_, _016382_, _016383_, _016384_, _016385_, _016386_, _016387_, _016388_, _016389_, _016390_, _016391_, _016392_, _016393_, _016394_, _016395_, _016396_, _016397_, _016398_, _016399_, _016400_, _016401_, _016402_, _016403_, _016404_, _016405_, _016406_, _016407_, _016408_, _016409_, _016410_, _016411_, _016412_, _016413_, _016414_, _016415_, _016416_, _016417_, _016418_, _016419_, _016420_, _016421_, _016422_, _016423_, _016424_, _016425_, _016426_, _016427_, _016428_, _016429_, _016430_, _016431_, _016432_, _016433_, _016434_, _016435_, _016436_, _016437_, _016438_, _016439_, _016440_, _016441_, _016442_, _016443_, _016444_, _016445_, _016446_, _016447_, _016448_, _016449_, _016450_, _016451_, _016452_, _016453_, _016454_, _016455_, _016456_, _016457_, _016458_, _016459_, _016460_, _016461_, _016462_, _016463_, _016464_, _016465_, _016466_, _016467_, _016468_, _016469_, _016470_, _016471_, _016472_, _016473_, _016474_, _016475_, _016476_, _016477_, _016478_, _016479_, _016480_, _016481_, _016482_, _016483_, _016484_, _016485_, _016486_, _016487_, _016488_, _016489_, _016490_, _016491_, _016492_, _016493_, _016494_, _016495_, _016496_, _016497_, _016498_, _016499_, _016500_, _016501_, _016502_, _016503_, _016504_, _016505_, _016506_, _016507_, _016508_, _016509_, _016510_, _016511_, _016512_, _016513_, _016514_, _016515_, _016516_, _016517_, _016518_, _016519_, _016520_, _016521_, _016522_, _016523_, _016524_, _016525_, _016526_, _016527_, _016528_, _016529_, _016530_, _016531_, _016532_, _016533_, _016534_, _016535_, _016536_, _016537_, _016538_, _016539_, _016540_, _016541_, _016542_, _016543_, _016544_, _016545_, _016546_, _016547_, _016548_, _016549_, _016550_, _016551_, _016552_, _016553_, _016554_, _016555_, _016556_, _016557_, _016558_, _016559_, _016560_, _016561_, _016562_, _016563_, _016564_, _016565_, _016566_, _016567_, _016568_, _016569_, _016570_, _016571_, _016572_, _016573_, _016574_, _016575_, _016576_, _016577_, _016578_, _016579_, _016580_, _016581_, _016582_, _016583_, _016584_, _016585_, _016586_, _016587_, _016588_, _016589_, _016590_, _016591_, _016592_, _016593_, _016594_, _016595_, _016596_, _016597_, _016598_, _016599_, _016600_, _016601_, _016602_, _016603_, _016604_, _016605_, _016606_, _016607_, _016608_, _016609_, _016610_, _016611_, _016612_, _016613_, _016614_, _016615_, _016616_, _016617_, _016618_, _016619_, _016620_, _016621_, _016622_, _016623_, _016624_, _016625_, _016626_, _016627_, _016628_, _016629_, _016630_, _016631_, _016632_, _016633_, _016634_, _016635_, _016636_, _016637_, _016638_, _016639_, _016640_, _016641_, _016642_, _016643_, _016644_, _016645_, _016646_, _016647_, _016648_, _016649_, _016650_, _016651_, _016652_, _016653_, _016654_, _016655_, _016656_, _016657_, _016658_, _016659_, _016660_, _016661_, _016662_, _016663_, _016664_, _016665_, _016666_, _016667_, _016668_, _016669_, _016670_, _016671_, _016672_, _016673_, _016674_, _016675_, _016676_, _016677_, _016678_, _016679_, _016680_, _016681_, _016682_, _016683_, _016684_, _016685_, _016686_, _016687_, _016688_, _016689_, _016690_, _016691_, _016692_, _016693_, _016694_, _016695_, _016696_, _016697_, _016698_, _016699_, _016700_, _016701_, _016702_, _016703_, _016704_, _016705_, _016706_, _016707_, _016708_, _016709_, _016710_, _016711_, _016712_, _016713_, _016714_, _016715_, _016716_, _016717_, _016718_, _016719_, _016720_, _016721_, _016722_, _016723_, _016724_, _016725_, _016726_, _016727_, _016728_, _016729_, _016730_, _016731_, _016732_, _016733_, _016734_, _016735_, _016736_, _016737_, _016738_, _016739_, _016740_, _016741_, _016742_, _016743_, _016744_, _016745_, _016746_, _016747_, _016748_, _016749_, _016750_, _016751_, _016752_, _016753_, _016754_, _016755_, _016756_, _016757_, _016758_, _016759_, _016760_, _016761_, _016762_, _016763_, _016764_, _016765_, _016766_, _016767_, _016768_, _016769_, _016770_, _016771_, _016772_, _016773_, _016774_, _016775_, _016776_, _016777_, _016778_, _016779_, _016780_, _016781_, _016782_, _016783_, _016784_, _016785_, _016786_, _016787_, _016788_, _016789_, _016790_, _016791_, _016792_, _016793_, _016794_, _016795_, _016796_, _016797_, _016798_, _016799_, _016800_, _016801_, _016802_, _016803_, _016804_, _016805_, _016806_, _016807_, _016808_, _016809_, _016810_, _016811_, _016812_, _016813_, _016814_, _016815_, _016816_, _016817_, _016818_, _016819_, _016820_, _016821_, _016822_, _016823_, _016824_, _016825_, _016826_, _016827_, _016828_, _016829_, _016830_, _016831_, _016832_, _016833_, _016834_, _016835_, _016836_, _016837_, _016838_, _016839_, _016840_, _016841_, _016842_, _016843_, _016844_, _016845_, _016846_, _016847_, _016848_, _016849_, _016850_, _016851_, _016852_, _016853_, _016854_, _016855_, _016856_, _016857_, _016858_, _016859_, _016860_, _016861_, _016862_, _016863_, _016864_, _016865_, _016866_, _016867_, _016868_, _016869_, _016870_, _016871_, _016872_, _016873_, _016874_, _016875_, _016876_, _016877_, _016878_, _016879_, _016880_, _016881_, _016882_, _016883_, _016884_, _016885_, _016886_, _016887_, _016888_, _016889_, _016890_, _016891_, _016892_, _016893_, _016894_, _016895_, _016896_, _016897_, _016898_, _016899_, _016900_, _016901_, _016902_, _016903_, _016904_, _016905_, _016906_, _016907_, _016908_, _016909_, _016910_, _016911_, _016912_, _016913_, _016914_, _016915_, _016916_, _016917_, _016918_, _016919_, _016920_, _016921_, _016922_, _016923_, _016924_, _016925_, _016926_, _016927_, _016928_, _016929_, _016930_, _016931_, _016932_, _016933_, _016934_, _016935_, _016936_, _016937_, _016938_, _016939_, _016940_, _016941_, _016942_, _016943_, _016944_, _016945_, _016946_, _016947_, _016948_, _016949_, _016950_, _016951_, _016952_, _016953_, _016954_, _016955_, _016956_, _016957_, _016958_, _016959_, _016960_, _016961_, _016962_, _016963_, _016964_, _016965_, _016966_, _016967_, _016968_, _016969_, _016970_, _016971_, _016972_, _016973_, _016974_, _016975_, _016976_, _016977_, _016978_, _016979_, _016980_, _016981_, _016982_, _016983_, _016984_, _016985_, _016986_, _016987_, _016988_, _016989_, _016990_, _016991_, _016992_, _016993_, _016994_, _016995_, _016996_, _016997_, _016998_, _016999_, _017000_, _017001_, _017002_, _017003_, _017004_, _017005_, _017006_, _017007_, _017008_, _017009_, _017010_, _017011_, _017012_, _017013_, _017014_, _017015_, _017016_, _017017_, _017018_, _017019_, _017020_, _017021_, _017022_, _017023_, _017024_, _017025_, _017026_, _017027_, _017028_, _017029_, _017030_, _017031_, _017032_, _017033_, _017034_, _017035_, _017036_, _017037_, _017038_, _017039_, _017040_, _017041_, _017042_, _017043_, _017044_, _017045_, _017046_, _017047_, _017048_, _017049_, _017050_, _017051_, _017052_, _017053_, _017054_, _017055_, _017056_, _017057_, _017058_, _017059_, _017060_, _017061_, _017062_, _017063_, _017064_, _017065_, _017066_, _017067_, _017068_, _017069_, _017070_, _017071_, _017072_, _017073_, _017074_, _017075_, _017076_, _017077_, _017078_, _017079_, _017080_, _017081_, _017082_, _017083_, _017084_, _017085_, _017086_, _017087_, _017088_, _017089_, _017090_, _017091_, _017092_, _017093_, _017094_, _017095_, _017096_, _017097_, _017098_, _017099_, _017100_, _017101_, _017102_, _017103_, _017104_, _017105_, _017106_, _017107_, _017108_, _017109_, _017110_, _017111_, _017112_, _017113_, _017114_, _017115_, _017116_, _017117_, _017118_, _017119_, _017120_, _017121_, _017122_, _017123_, _017124_, _017125_, _017126_, _017127_, _017128_, _017129_, _017130_, _017131_, _017132_, _017133_, _017134_, _017135_, _017136_, _017137_, _017138_, _017139_, _017140_, _017141_, _017142_, _017143_, _017144_, _017145_, _017146_, _017147_, _017148_, _017149_, _017150_, _017151_, _017152_, _017153_, _017154_, _017155_, _017156_, _017157_, _017158_, _017159_, _017160_, _017161_, _017162_, _017163_, _017164_, _017165_, _017166_, _017167_, _017168_, _017169_, _017170_, _017171_, _017172_, _017173_, _017174_, _017175_, _017176_, _017177_, _017178_, _017179_, _017180_, _017181_, _017182_, _017183_, _017184_, _017185_, _017186_, _017187_, _017188_, _017189_, _017190_, _017191_, _017192_, _017193_, _017194_, _017195_, _017196_, _017197_, _017198_, _017199_, _017200_, _017201_, _017202_, _017203_, _017204_, _017205_, _017206_, _017207_, _017208_, _017209_, _017210_, _017211_, _017212_, _017213_, _017214_, _017215_, _017216_, _017217_, _017218_, _017219_, _017220_, _017221_, _017222_, _017223_, _017224_, _017225_, _017226_, _017227_, _017228_, _017229_, _017230_, _017231_, _017232_, _017233_, _017234_, _017235_, _017236_, _017237_, _017238_, _017239_, _017240_, _017241_, _017242_, _017243_, _017244_, _017245_, _017246_, _017247_, _017248_, _017249_, _017250_, _017251_, _017252_, _017253_, _017254_, _017255_, _017256_, _017257_, _017258_, _017259_, _017260_, _017261_, _017262_, _017263_, _017264_, _017265_, _017266_, _017267_, _017268_, _017269_, _017270_, _017271_, _017272_, _017273_, _017274_, _017275_, _017276_, _017277_, _017278_, _017279_, _017280_, _017281_, _017282_, _017283_, _017284_, _017285_, _017286_, _017287_, _017288_, _017289_, _017290_, _017291_, _017292_, _017293_, _017294_, _017295_, _017296_, _017297_, _017298_, _017299_, _017300_, _017301_, _017302_, _017303_, _017304_, _017305_, _017306_, _017307_, _017308_, _017309_, _017310_, _017311_, _017312_, _017313_, _017314_, _017315_, _017316_, _017317_, _017318_, _017319_, _017320_, _017321_, _017322_, _017323_, _017324_, _017325_, _017326_, _017327_, _017328_, _017329_, _017330_, _017331_, _017332_, _017333_, _017334_, _017335_, _017336_, _017337_, _017338_, _017339_, _017340_, _017341_, _017342_, _017343_, _017344_, _017345_, _017346_, _017347_, _017348_, _017349_, _017350_, _017351_, _017352_, _017353_, _017354_, _017355_, _017356_, _017357_, _017358_, _017359_, _017360_, _017361_, _017362_, _017363_, _017364_, _017365_, _017366_, _017367_, _017368_, _017369_, _017370_, _017371_, _017372_, _017373_, _017374_, _017375_, _017376_, _017377_, _017378_, _017379_, _017380_, _017381_, _017382_, _017383_, _017384_, _017385_, _017386_, _017387_, _017388_, _017389_, _017390_, _017391_, _017392_, _017393_, _017394_, _017395_, _017396_, _017397_, _017398_, _017399_, _017400_, _017401_, _017402_, _017403_, _017404_, _017405_, _017406_, _017407_, _017408_, _017409_, _017410_, _017411_, _017412_, _017413_, _017414_, _017415_, _017416_, _017417_, _017418_, _017419_, _017420_, _017421_, _017422_, _017423_, _017424_, _017425_, _017426_, _017427_, _017428_, _017429_, _017430_, _017431_, _017432_, _017433_, _017434_, _017435_, _017436_, _017437_, _017438_, _017439_, _017440_, _017441_, _017442_, _017443_, _017444_, _017445_, _017446_, _017447_, _017448_, _017449_, _017450_, _017451_, _017452_, _017453_, _017454_, _017455_, _017456_, _017457_, _017458_, _017459_, _017460_, _017461_, _017462_, _017463_, _017464_, _017465_, _017466_, _017467_, _017468_, _017469_, _017470_, _017471_, _017472_, _017473_, _017474_, _017475_, _017476_, _017477_, _017478_, _017479_, _017480_, _017481_, _017482_, _017483_, _017484_, _017485_, _017486_, _017487_, _017488_, _017489_, _017490_, _017491_, _017492_, _017493_, _017494_, _017495_, _017496_, _017497_, _017498_, _017499_, _017500_, _017501_, _017502_, _017503_, _017504_, _017505_, _017506_, _017507_, _017508_, _017509_, _017510_, _017511_, _017512_, _017513_, _017514_, _017515_, _017516_, _017517_, _017518_, _017519_, _017520_, _017521_, _017522_, _017523_, _017524_, _017525_, _017526_, _017527_, _017528_, _017529_, _017530_, _017531_, _017532_, _017533_, _017534_, _017535_, _017536_, _017537_, _017538_, _017539_, _017540_, _017541_, _017542_, _017543_, _017544_, _017545_, _017546_, _017547_, _017548_, _017549_, _017550_, _017551_, _017552_, _017553_, _017554_, _017555_, _017556_, _017557_, _017558_, _017559_, _017560_, _017561_, _017562_, _017563_, _017564_, _017565_, _017566_, _017567_, _017568_, _017569_, _017570_, _017571_, _017572_, _017573_, _017574_, _017575_, _017576_, _017577_, _017578_, _017579_, _017580_, _017581_, _017582_, _017583_, _017584_, _017585_, _017586_, _017587_, _017588_, _017589_, _017590_, _017591_, _017592_, _017593_, _017594_, _017595_, _017596_, _017597_, _017598_, _017599_, _017600_, _017601_, _017602_, _017603_, _017604_, _017605_, _017606_, _017607_, _017608_, _017609_, _017610_, _017611_, _017612_, _017613_, _017614_, _017615_, _017616_, _017617_, _017618_, _017619_, _017620_, _017621_, _017622_, _017623_, _017624_, _017625_, _017626_, _017627_, _017628_, _017629_, _017630_, _017631_, _017632_, _017633_, _017634_, _017635_, _017636_, _017637_, _017638_, _017639_, _017640_, _017641_, _017642_, _017643_, _017644_, _017645_, _017646_, _017647_, _017648_, _017649_, _017650_, _017651_, _017652_, _017653_, _017654_, _017655_, _017656_, _017657_, _017658_, _017659_, _017660_, _017661_, _017662_, _017663_, _017664_, _017665_, _017666_, _017667_, _017668_, _017669_, _017670_, _017671_, _017672_, _017673_, _017674_, _017675_, _017676_, _017677_, _017678_, _017679_, _017680_, _017681_, _017682_, _017683_, _017684_, _017685_, _017686_, _017687_, _017688_, _017689_, _017690_, _017691_, _017692_, _017693_, _017694_, _017695_, _017696_, _017697_, _017698_, _017699_, _017700_, _017701_, _017702_, _017703_, _017704_, _017705_, _017706_, _017707_, _017708_, _017709_, _017710_, _017711_, _017712_, _017713_, _017714_, _017715_, _017716_, _017717_, _017718_, _017719_, _017720_, _017721_, _017722_, _017723_, _017724_, _017725_, _017726_, _017727_, _017728_, _017729_, _017730_, _017731_, _017732_, _017733_, _017734_, _017735_, _017736_, _017737_, _017738_, _017739_, _017740_, _017741_, _017742_, _017743_, _017744_, _017745_, _017746_, _017747_, _017748_, _017749_, _017750_, _017751_, _017752_, _017753_, _017754_, _017755_, _017756_, _017757_, _017758_, _017759_, _017760_, _017761_, _017762_, _017763_, _017764_, _017765_, _017766_, _017767_, _017768_, _017769_, _017770_, _017771_, _017772_, _017773_, _017774_, _017775_, _017776_, _017777_, _017778_, _017779_, _017780_, _017781_, _017782_, _017783_, _017784_, _017785_, _017786_, _017787_, _017788_, _017789_, _017790_, _017791_, _017792_, _017793_, _017794_, _017795_, _017796_, _017797_, _017798_, _017799_, _017800_, _017801_, _017802_, _017803_, _017804_, _017805_, _017806_, _017807_, _017808_, _017809_, _017810_, _017811_, _017812_, _017813_, _017814_, _017815_, _017816_, _017817_, _017818_, _017819_, _017820_, _017821_, _017822_, _017823_, _017824_, _017825_, _017826_, _017827_, _017828_, _017829_, _017830_, _017831_, _017832_, _017833_, _017834_, _017835_, _017836_, _017837_, _017838_, _017839_, _017840_, _017841_, _017842_, _017843_, _017844_, _017845_, _017846_, _017847_, _017848_, _017849_, _017850_, _017851_, _017852_, _017853_, _017854_, _017855_, _017856_, _017857_, _017858_, _017859_, _017860_, _017861_, _017862_, _017863_, _017864_, _017865_, _017866_, _017867_, _017868_, _017869_, _017870_, _017871_, _017872_, _017873_, _017874_, _017875_, _017876_, _017877_, _017878_, _017879_, _017880_, _017881_, _017882_, _017883_, _017884_, _017885_, _017886_, _017887_, _017888_, _017889_, _017890_, _017891_, _017892_, _017893_, _017894_, _017895_, _017896_, _017897_, _017898_, _017899_, _017900_, _017901_, _017902_, _017903_, _017904_, _017905_, _017906_, _017907_, _017908_, _017909_, _017910_, _017911_, _017912_, _017913_, _017914_, _017915_, _017916_, _017917_, _017918_, _017919_, _017920_, _017921_, _017922_, _017923_, _017924_, _017925_, _017926_, _017927_, _017928_, _017929_, _017930_, _017931_, _017932_, _017933_, _017934_, _017935_, _017936_, _017937_, _017938_, _017939_, _017940_, _017941_, _017942_, _017943_, _017944_, _017945_, _017946_, _017947_, _017948_, _017949_, _017950_, _017951_, _017952_, _017953_, _017954_, _017955_, _017956_, _017957_, _017958_, _017959_, _017960_, _017961_, _017962_, _017963_, _017964_, _017965_, _017966_, _017967_, _017968_, _017969_, _017970_, _017971_, _017972_, _017973_, _017974_, _017975_, _017976_, _017977_, _017978_, _017979_, _017980_, _017981_, _017982_, _017983_, _017984_, _017985_, _017986_, _017987_, _017988_, _017989_, _017990_, _017991_, _017992_, _017993_, _017994_, _017995_, _017996_, _017997_, _017998_, _017999_, _018000_, _018001_, _018002_, _018003_, _018004_, _018005_, _018006_, _018007_, _018008_, _018009_, _018010_, _018011_, _018012_, _018013_, _018014_, _018015_, _018016_, _018017_, _018018_, _018019_, _018020_, _018021_, _018022_, _018023_, _018024_, _018025_, _018026_, _018027_, _018028_, _018029_, _018030_, _018031_, _018032_, _018033_, _018034_, _018035_, _018036_, _018037_, _018038_, _018039_, _018040_, _018041_, _018042_, _018043_, _018044_, _018045_, _018046_, _018047_, _018048_, _018049_, _018050_, _018051_, _018052_, _018053_, _018054_, _018055_, _018056_, _018057_, _018058_, _018059_, _018060_, _018061_, _018062_, _018063_, _018064_, _018065_, _018066_, _018067_, _018068_, _018069_, _018070_, _018071_, _018072_, _018073_, _018074_, _018075_, _018076_, _018077_, _018078_, _018079_, _018080_, _018081_, _018082_, _018083_, _018084_, _018085_, _018086_, _018087_, _018088_, _018089_, _018090_, _018091_, _018092_, _018093_, _018094_, _018095_, _018096_, _018097_, _018098_, _018099_, _018100_, _018101_, _018102_, _018103_, _018104_, _018105_, _018106_, _018107_, _018108_, _018109_, _018110_, _018111_, _018112_, _018113_, _018114_, _018115_, _018116_, _018117_, _018118_, _018119_, _018120_, _018121_, _018122_, _018123_, _018124_, _018125_, _018126_, _018127_, _018128_, _018129_, _018130_, _018131_, _018132_, _018133_, _018134_, _018135_, _018136_, _018137_, _018138_, _018139_, _018140_, _018141_, _018142_, _018143_, _018144_, _018145_, _018146_, _018147_, _018148_, _018149_, _018150_, _018151_, _018152_, _018153_, _018154_, _018155_, _018156_, _018157_, _018158_, _018159_, _018160_, _018161_, _018162_, _018163_, _018164_, _018165_, _018166_, _018167_, _018168_, _018169_, _018170_, _018171_, _018172_, _018173_, _018174_, _018175_, _018176_, _018177_, _018178_, _018179_, _018180_, _018181_, _018182_, _018183_, _018184_, _018185_, _018186_, _018187_, _018188_, _018189_, _018190_, _018191_, _018192_, _018193_, _018194_, _018195_, _018196_, _018197_, _018198_, _018199_, _018200_, _018201_, _018202_, _018203_, _018204_, _018205_, _018206_, _018207_, _018208_, _018209_, _018210_, _018211_, _018212_, _018213_, _018214_, _018215_, _018216_, _018217_, _018218_, _018219_, _018220_, _018221_, _018222_, _018223_, _018224_, _018225_, _018226_, _018227_, _018228_, _018229_, _018230_, _018231_, _018232_, _018233_, _018234_, _018235_, _018236_, _018237_, _018238_, _018239_, _018240_, _018241_, _018242_, _018243_, _018244_, _018245_, _018246_, _018247_, _018248_, _018249_, _018250_, _018251_, _018252_, _018253_, _018254_, _018255_, _018256_, _018257_, _018258_, _018259_, _018260_, _018261_, _018262_, _018263_, _018264_, _018265_, _018266_, _018267_, _018268_, _018269_, _018270_, _018271_, _018272_, _018273_, _018274_, _018275_, _018276_, _018277_, _018278_, _018279_, _018280_, _018281_, _018282_, _018283_, _018284_, _018285_, _018286_, _018287_, _018288_, _018289_, _018290_, _018291_, _018292_, _018293_, _018294_, _018295_, _018296_, _018297_, _018298_, _018299_, _018300_, _018301_, _018302_, _018303_, _018304_, _018305_, _018306_, _018307_, _018308_, _018309_, _018310_, _018311_, _018312_, _018313_, _018314_, _018315_, _018316_, _018317_, _018318_, _018319_, _018320_, _018321_, _018322_, _018323_, _018324_, _018325_, _018326_, _018327_, _018328_, _018329_, _018330_, _018331_, _018332_, _018333_, _018334_, _018335_, _018336_, _018337_, _018338_, _018339_, _018340_, _018341_, _018342_, _018343_, _018344_, _018345_, _018346_, _018347_, _018348_, _018349_, _018350_, _018351_, _018352_, _018353_, _018354_, _018355_, _018356_, _018357_, _018358_, _018359_, _018360_, _018361_, _018362_, _018363_, _018364_, _018365_, _018366_, _018367_, _018368_, _018369_, _018370_, _018371_, _018372_, _018373_, _018374_, _018375_, _018376_, _018377_, _018378_, _018379_, _018380_, _018381_, _018382_, _018383_, _018384_, _018385_, _018386_, _018387_, _018388_, _018389_, _018390_, _018391_, _018392_, _018393_, _018394_, _018395_, _018396_, _018397_, _018398_, _018399_, _018400_, _018401_, _018402_, _018403_, _018404_, _018405_, _018406_, _018407_, _018408_, _018409_, _018410_, _018411_, _018412_, _018413_, _018414_, _018415_, _018416_, _018417_, _018418_, _018419_, _018420_, _018421_, _018422_, _018423_, _018424_, _018425_, _018426_, _018427_, _018428_, _018429_, _018430_, _018431_, _018432_, _018433_, _018434_, _018435_, _018436_, _018437_, _018438_, _018439_, _018440_, _018441_, _018442_, _018443_, _018444_, _018445_, _018446_, _018447_, _018448_, _018449_, _018450_, _018451_, _018452_, _018453_, _018454_, _018455_, _018456_, _018457_, _018458_, _018459_, _018460_, _018461_, _018462_, _018463_, _018464_, _018465_, _018466_, _018467_, _018468_, _018469_, _018470_, _018471_, _018472_, _018473_, _018474_, _018475_, _018476_, _018477_, _018478_, _018479_, _018480_, _018481_, _018482_, _018483_, _018484_, _018485_, _018486_, _018487_, _018488_, _018489_, _018490_, _018491_, _018492_, _018493_, _018494_, _018495_, _018496_, _018497_, _018498_, _018499_, _018500_, _018501_, _018502_, _018503_, _018504_, _018505_, _018506_, _018507_, _018508_, _018509_, _018510_, _018511_, _018512_, _018513_, _018514_, _018515_, _018516_, _018517_, _018518_, _018519_, _018520_, _018521_, _018522_, _018523_, _018524_, _018525_, _018526_, _018527_, _018528_, _018529_, _018530_, _018531_, _018532_, _018533_, _018534_, _018535_, _018536_, _018537_, _018538_, _018539_, _018540_, _018541_, _018542_, _018543_, _018544_, _018545_, _018546_, _018547_, _018548_, _018549_, _018550_, _018551_, _018552_, _018553_, _018554_, _018555_, _018556_, _018557_, _018558_, _018559_, _018560_, _018561_, _018562_, _018563_, _018564_, _018565_, _018566_, _018567_, _018568_, _018569_, _018570_, _018571_, _018572_, _018573_, _018574_, _018575_, _018576_, _018577_, _018578_, _018579_, _018580_, _018581_, _018582_, _018583_, _018584_, _018585_, _018586_, _018587_, _018588_, _018589_, _018590_, _018591_, _018592_, _018593_, _018594_, _018595_, _018596_, _018597_, _018598_, _018599_, _018600_, _018601_, _018602_, _018603_, _018604_, _018605_, _018606_, _018607_, _018608_, _018609_, _018610_, _018611_, _018612_, _018613_, _018614_, _018615_, _018616_, _018617_, _018618_, _018619_, _018620_, _018621_, _018622_, _018623_, _018624_, _018625_, _018626_, _018627_, _018628_, _018629_, _018630_, _018631_, _018632_, _018633_, _018634_, _018635_, _018636_, _018637_, _018638_, _018639_, _018640_, _018641_, _018642_, _018643_, _018644_, _018645_, _018646_, _018647_, _018648_, _018649_, _018650_, _018651_, _018652_, _018653_, _018654_, _018655_, _018656_, _018657_, _018658_, _018659_, _018660_, _018661_, _018662_, _018663_, _018664_, _018665_, _018666_, _018667_, _018668_, _018669_, _018670_, _018671_, _018672_, _018673_, _018674_, _018675_, _018676_, _018677_, _018678_, _018679_, _018680_, _018681_, _018682_, _018683_, _018684_, _018685_, _018686_, _018687_, _018688_, _018689_, _018690_, _018691_, _018692_, _018693_, _018694_, _018695_, _018696_, _018697_, _018698_, _018699_, _018700_, _018701_, _018702_, _018703_, _018704_, _018705_, _018706_, _018707_, _018708_, _018709_, _018710_, _018711_, _018712_, _018713_, _018714_, _018715_, _018716_, _018717_, _018718_, _018719_, _018720_, _018721_, _018722_, _018723_, _018724_, _018725_, _018726_, _018727_, _018728_, _018729_, _018730_, _018731_, _018732_, _018733_, _018734_, _018735_, _018736_, _018737_, _018738_, _018739_, _018740_, _018741_, _018742_, _018743_, _018744_, _018745_, _018746_, _018747_, _018748_, _018749_, _018750_, _018751_, _018752_, _018753_, _018754_, _018755_, _018756_, _018757_, _018758_, _018759_, _018760_, _018761_, _018762_, _018763_, _018764_, _018765_, _018766_, _018767_, _018768_, _018769_, _018770_, _018771_, _018772_, _018773_, _018774_, _018775_, _018776_, _018777_, _018778_, _018779_, _018780_, _018781_, _018782_, _018783_, _018784_, _018785_, _018786_, _018787_, _018788_, _018789_, _018790_, _018791_, _018792_, _018793_, _018794_, _018795_, _018796_, _018797_, _018798_, _018799_, _018800_, _018801_, _018802_, _018803_, _018804_, _018805_, _018806_, _018807_, _018808_, _018809_, _018810_, _018811_, _018812_, _018813_, _018814_, _018815_, _018816_, _018817_, _018818_, _018819_, _018820_, _018821_, _018822_, _018823_, _018824_, _018825_, _018826_, _018827_, _018828_, _018829_, _018830_, _018831_, _018832_, _018833_, _018834_, _018835_, _018836_, _018837_, _018838_, _018839_, _018840_, _018841_, _018842_, _018843_, _018844_, _018845_, _018846_, _018847_, _018848_, _018849_, _018850_, _018851_, _018852_, _018853_, _018854_, _018855_, _018856_, _018857_, _018858_, _018859_, _018860_, _018861_, _018862_, _018863_, _018864_, _018865_, _018866_, _018867_, _018868_, _018869_, _018870_, _018871_, _018872_, _018873_, _018874_, _018875_, _018876_, _018877_, _018878_, _018879_, _018880_, _018881_, _018882_, _018883_, _018884_, _018885_, _018886_, _018887_, _018888_, _018889_, _018890_, _018891_, _018892_, _018893_, _018894_, _018895_, _018896_, _018897_, _018898_, _018899_, _018900_, _018901_, _018902_, _018903_, _018904_, _018905_, _018906_, _018907_, _018908_, _018909_, _018910_, _018911_, _018912_, _018913_, _018914_, _018915_, _018916_, _018917_, _018918_, _018919_, _018920_, _018921_, _018922_, _018923_, _018924_, _018925_, _018926_, _018927_, _018928_, _018929_, _018930_, _018931_, _018932_, _018933_, _018934_, _018935_, _018936_, _018937_, _018938_, _018939_, _018940_, _018941_, _018942_, _018943_, _018944_, _018945_, _018946_, _018947_, _018948_, _018949_, _018950_, _018951_, _018952_, _018953_, _018954_, _018955_, _018956_, _018957_, _018958_, _018959_, _018960_, _018961_, _018962_, _018963_, _018964_, _018965_, _018966_, _018967_, _018968_, _018969_, _018970_, _018971_, _018972_, _018973_, _018974_, _018975_, _018976_, _018977_, _018978_, _018979_, _018980_, _018981_, _018982_, _018983_, _018984_, _018985_, _018986_, _018987_, _018988_, _018989_, _018990_, _018991_, _018992_, _018993_, _018994_, _018995_, _018996_, _018997_, _018998_, _018999_, _019000_, _019001_, _019002_, _019003_, _019004_, _019005_, _019006_, _019007_, _019008_, _019009_, _019010_, _019011_, _019012_, _019013_, _019014_, _019015_, _019016_, _019017_, _019018_, _019019_, _019020_, _019021_, _019022_, _019023_, _019024_, _019025_, _019026_, _019027_, _019028_, _019029_, _019030_, _019031_, _019032_, _019033_, _019034_, _019035_, _019036_, _019037_, _019038_, _019039_, _019040_, _019041_, _019042_, _019043_, _019044_, _019045_, _019046_, _019047_, _019048_, _019049_, _019050_, _019051_, _019052_, _019053_, _019054_, _019055_, _019056_, _019057_, _019058_, _019059_, _019060_, _019061_, _019062_, _019063_, _019064_, _019065_, _019066_, _019067_, _019068_, _019069_, _019070_, _019071_, _019072_, _019073_, _019074_, _019075_, _019076_, _019077_, _019078_, _019079_, _019080_, _019081_, _019082_, _019083_, _019084_, _019085_, _019086_, _019087_, _019088_, _019089_, _019090_, _019091_, _019092_, _019093_, _019094_, _019095_, _019096_, _019097_, _019098_, _019099_, _019100_, _019101_, _019102_, _019103_, _019104_, _019105_, _019106_, _019107_, _019108_, _019109_, _019110_, _019111_, _019112_, _019113_, _019114_, _019115_, _019116_, _019117_, _019118_, _019119_, _019120_, _019121_, _019122_, _019123_, _019124_, _019125_, _019126_, _019127_, _019128_, _019129_, _019130_, _019131_, _019132_, _019133_, _019134_, _019135_, _019136_, _019137_, _019138_, _019139_, _019140_, _019141_, _019142_, _019143_, _019144_, _019145_, _019146_, _019147_, _019148_, _019149_, _019150_, _019151_, _019152_, _019153_, _019154_, _019155_, _019156_, _019157_, _019158_, _019159_, _019160_, _019161_, _019162_, _019163_, _019164_, _019165_, _019166_, _019167_, _019168_, _019169_, _019170_, _019171_, _019172_, _019173_, _019174_, _019175_, _019176_, _019177_, _019178_, _019179_, _019180_, _019181_, _019182_, _019183_, _019184_, _019185_, _019186_, _019187_, _019188_, _019189_, _019190_, _019191_, _019192_, _019193_, _019194_, _019195_, _019196_, _019197_, _019198_, _019199_, _019200_, _019201_, _019202_, _019203_, _019204_, _019205_, _019206_, _019207_, _019208_, _019209_, _019210_, _019211_, _019212_, _019213_, _019214_, _019215_, _019216_, _019217_, _019218_, _019219_, _019220_, _019221_, _019222_, _019223_, _019224_, _019225_, _019226_, _019227_, _019228_, _019229_, _019230_, _019231_, _019232_, _019233_, _019234_, _019235_, _019236_, _019237_, _019238_, _019239_, _019240_, _019241_, _019242_, _019243_, _019244_, _019245_, _019246_, _019247_, _019248_, _019249_, _019250_, _019251_, _019252_, _019253_, _019254_, _019255_, _019256_, _019257_, _019258_, _019259_, _019260_, _019261_, _019262_, _019263_, _019264_, _019265_, _019266_, _019267_, _019268_, _019269_, _019270_, _019271_, _019272_, _019273_, _019274_, _019275_, _019276_, _019277_, _019278_, _019279_, _019280_, _019281_, _019282_, _019283_, _019284_, _019285_, _019286_, _019287_, _019288_, _019289_, _019290_, _019291_, _019292_, _019293_, _019294_, _019295_, _019296_, _019297_, _019298_, _019299_, _019300_, _019301_, _019302_, _019303_, _019304_, _019305_, _019306_, _019307_, _019308_, _019309_, _019310_, _019311_, _019312_, _019313_, _019314_, _019315_, _019316_, _019317_, _019318_, _019319_, _019320_, _019321_, _019322_, _019323_, _019324_, _019325_, _019326_, _019327_, _019328_, _019329_, _019330_, _019331_, _019332_, _019333_, _019334_, _019335_, _019336_, _019337_, _019338_, _019339_, _019340_, _019341_, _019342_, _019343_, _019344_, _019345_, _019346_, _019347_, _019348_, _019349_, _019350_, _019351_, _019352_, _019353_, _019354_, _019355_, _019356_, _019357_, _019358_, _019359_, _019360_, _019361_, _019362_, _019363_, _019364_, _019365_, _019366_, _019367_, _019368_, _019369_, _019370_, _019371_, _019372_, _019373_, _019374_, _019375_, _019376_, _019377_, _019378_, _019379_, _019380_, _019381_, _019382_, _019383_, _019384_, _019385_, _019386_, _019387_, _019388_, _019389_, _019390_, _019391_, _019392_, _019393_, _019394_, _019395_, _019396_, _019397_, _019398_, _019399_, _019400_, _019401_, _019402_, _019403_, _019404_, _019405_, _019406_, _019407_, _019408_, _019409_, _019410_, _019411_, _019412_, _019413_, _019414_, _019415_, _019416_, _019417_, _019418_, _019419_, _019420_, _019421_, _019422_, _019423_, _019424_, _019425_, _019426_, _019427_, _019428_, _019429_, _019430_, _019431_, _019432_, _019433_, _019434_, _019435_, _019436_, _019437_, _019438_, _019439_, _019440_, _019441_, _019442_, _019443_, _019444_, _019445_, _019446_, _019447_, _019448_, _019449_, _019450_, _019451_, _019452_, _019453_, _019454_, _019455_, _019456_, _019457_, _019458_, _019459_, _019460_, _019461_, _019462_, _019463_, _019464_, _019465_, _019466_, _019467_, _019468_, _019469_, _019470_, _019471_, _019472_, _019473_, _019474_, _019475_, _019476_, _019477_, _019478_, _019479_, _019480_, _019481_, _019482_, _019483_, _019484_, _019485_, _019486_, _019487_, _019488_, _019489_, _019490_, _019491_, _019492_, _019493_, _019494_, _019495_, _019496_, _019497_, _019498_, _019499_, _019500_, _019501_, _019502_, _019503_, _019504_, _019505_, _019506_, _019507_, _019508_, _019509_, _019510_, _019511_, _019512_, _019513_, _019514_, _019515_, _019516_, _019517_, _019518_, _019519_, _019520_, _019521_, _019522_, _019523_, _019524_, _019525_, _019526_, _019527_, _019528_, _019529_, _019530_, _019531_, _019532_, _019533_, _019534_, _019535_, _019536_, _019537_, _019538_, _019539_, _019540_, _019541_, _019542_, _019543_, _019544_, _019545_, _019546_, _019547_, _019548_, _019549_, _019550_, _019551_, _019552_, _019553_, _019554_, _019555_, _019556_, _019557_, _019558_, _019559_, _019560_, _019561_, _019562_, _019563_, _019564_, _019565_, _019566_, _019567_, _019568_, _019569_, _019570_, _019571_, _019572_, _019573_, _019574_, _019575_, _019576_, _019577_, _019578_, _019579_, _019580_, _019581_, _019582_, _019583_, _019584_, _019585_, _019586_, _019587_, _019588_, _019589_, _019590_, _019591_, _019592_, _019593_, _019594_, _019595_, _019596_, _019597_, _019598_, _019599_, _019600_, _019601_, _019602_, _019603_, _019604_, _019605_, _019606_, _019607_, _019608_, _019609_, _019610_, _019611_, _019612_, _019613_, _019614_, _019615_, _019616_, _019617_, _019618_, _019619_, _019620_, _019621_, _019622_, _019623_, _019624_, _019625_, _019626_, _019627_, _019628_, _019629_, _019630_, _019631_, _019632_, _019633_, _019634_, _019635_, _019636_, _019637_, _019638_, _019639_, _019640_, _019641_, _019642_, _019643_, _019644_, _019645_, _019646_, _019647_, _019648_, _019649_, _019650_, _019651_, _019652_, _019653_, _019654_, _019655_, _019656_, _019657_, _019658_, _019659_, _019660_, _019661_, _019662_, _019663_, _019664_, _019665_, _019666_, _019667_, _019668_, _019669_, _019670_, _019671_, _019672_, _019673_, _019674_, _019675_, _019676_, _019677_, _019678_, _019679_, _019680_, _019681_, _019682_, _019683_, _019684_, _019685_, _019686_, _019687_, _019688_, _019689_, _019690_, _019691_, _019692_, _019693_, _019694_, _019695_, _019696_, _019697_, _019698_, _019699_, _019700_, _019701_, _019702_, _019703_, _019704_, _019705_, _019706_, _019707_, _019708_, _019709_, _019710_, _019711_, _019712_, _019713_, _019714_, _019715_, _019716_, _019717_, _019718_, _019719_, _019720_, _019721_, _019722_, _019723_, _019724_, _019725_, _019726_, _019727_, _019728_, _019729_, _019730_, _019731_, _019732_, _019733_, _019734_, _019735_, _019736_, _019737_, _019738_, _019739_, _019740_, _019741_, _019742_, _019743_, _019744_, _019745_, _019746_, _019747_, _019748_, _019749_, _019750_, _019751_, _019752_, _019753_, _019754_, _019755_, _019756_, _019757_, _019758_, _019759_, _019760_, _019761_, _019762_, _019763_, _019764_, _019765_, _019766_, _019767_, _019768_, _019769_, _019770_, _019771_, _019772_, _019773_, _019774_, _019775_, _019776_, _019777_, _019778_, _019779_, _019780_, _019781_, _019782_, _019783_, _019784_, _019785_, _019786_, _019787_, _019788_, _019789_, _019790_, _019791_, _019792_, _019793_, _019794_, _019795_, _019796_, _019797_, _019798_, _019799_, _019800_, _019801_, _019802_, _019803_, _019804_, _019805_, _019806_, _019807_, _019808_, _019809_, _019810_, _019811_, _019812_, _019813_, _019814_, _019815_, _019816_, _019817_, _019818_, _019819_, _019820_, _019821_, _019822_, _019823_, _019824_, _019825_, _019826_, _019827_, _019828_, _019829_, _019830_, _019831_, _019832_, _019833_, _019834_, _019835_, _019836_, _019837_, _019838_, _019839_, _019840_, _019841_, _019842_, _019843_, _019844_, _019845_, _019846_, _019847_, _019848_, _019849_, _019850_, _019851_, _019852_, _019853_, _019854_, _019855_, _019856_, _019857_, _019858_, _019859_, _019860_, _019861_, _019862_, _019863_, _019864_, _019865_, _019866_, _019867_, _019868_, _019869_, _019870_, _019871_, _019872_, _019873_, _019874_, _019875_, _019876_, _019877_, _019878_, _019879_, _019880_, _019881_, _019882_, _019883_, _019884_, _019885_, _019886_, _019887_, _019888_, _019889_, _019890_, _019891_, _019892_, _019893_, _019894_, _019895_, _019896_, _019897_, _019898_, _019899_, _019900_, _019901_, _019902_, _019903_, _019904_, _019905_, _019906_, _019907_, _019908_, _019909_, _019910_, _019911_, _019912_, _019913_, _019914_, _019915_, _019916_, _019917_, _019918_, _019919_, _019920_, _019921_, _019922_, _019923_, _019924_, _019925_, _019926_, _019927_, _019928_, _019929_, _019930_, _019931_, _019932_, _019933_, _019934_, _019935_, _019936_, _019937_, _019938_, _019939_, _019940_, _019941_, _019942_, _019943_, _019944_, _019945_, _019946_, _019947_, _019948_, _019949_, _019950_, _019951_, _019952_, _019953_, _019954_, _019955_, _019956_, _019957_, _019958_, _019959_, _019960_, _019961_, _019962_, _019963_, _019964_, _019965_, _019966_, _019967_, _019968_, _019969_, _019970_, _019971_, _019972_, _019973_, _019974_, _019975_, _019976_, _019977_, _019978_, _019979_, _019980_, _019981_, _019982_, _019983_, _019984_, _019985_, _019986_, _019987_, _019988_, _019989_, _019990_, _019991_, _019992_, _019993_, _019994_, _019995_, _019996_, _019997_, _019998_, _019999_, _020000_, _020001_, _020002_, _020003_, _020004_, _020005_, _020006_, _020007_, _020008_, _020009_, _020010_, _020011_, _020012_, _020013_, _020014_, _020015_, _020016_, _020017_, _020018_, _020019_, _020020_, _020021_, _020022_, _020023_, _020024_, _020025_, _020026_, _020027_, _020028_, _020029_, _020030_, _020031_, _020032_, _020033_, _020034_, _020035_, _020036_, _020037_, _020038_, _020039_, _020040_, _020041_, _020042_, _020043_, _020044_, _020045_, _020046_, _020047_, _020048_, _020049_, _020050_, _020051_, _020052_, _020053_, _020054_, _020055_, _020056_, _020057_, _020058_, _020059_, _020060_, _020061_, _020062_, _020063_, _020064_, _020065_, _020066_, _020067_, _020068_, _020069_, _020070_, _020071_, _020072_, _020073_, _020074_, _020075_, _020076_, _020077_, _020078_, _020079_, _020080_, _020081_, _020082_, _020083_, _020084_, _020085_, _020086_, _020087_, _020088_, _020089_, _020090_, _020091_, _020092_, _020093_, _020094_, _020095_, _020096_, _020097_, _020098_, _020099_, _020100_, _020101_, _020102_, _020103_, _020104_, _020105_, _020106_, _020107_, _020108_, _020109_, _020110_, _020111_, _020112_, _020113_, _020114_, _020115_, _020116_, _020117_, _020118_, _020119_, _020120_, _020121_, _020122_, _020123_, _020124_, _020125_, _020126_, _020127_, _020128_, _020129_, _020130_, _020131_, _020132_, _020133_, _020134_, _020135_, _020136_, _020137_, _020138_, _020139_, _020140_, _020141_, _020142_, _020143_, _020144_, _020145_, _020146_, _020147_, _020148_, _020149_, _020150_, _020151_, _020152_, _020153_, _020154_, _020155_, _020156_, _020157_, _020158_, _020159_, _020160_, _020161_, _020162_, _020163_, _020164_, _020165_, _020166_, _020167_, _020168_, _020169_, _020170_, _020171_, _020172_, _020173_, _020174_, _020175_, _020176_, _020177_, _020178_, _020179_, _020180_, _020181_, _020182_, _020183_, _020184_, _020185_, _020186_, _020187_, _020188_, _020189_, _020190_, _020191_, _020192_, _020193_, _020194_, _020195_, _020196_, _020197_, _020198_, _020199_, _020200_, _020201_, _020202_, _020203_, _020204_, _020205_, _020206_, _020207_, _020208_, _020209_, _020210_, _020211_, _020212_, _020213_, _020214_, _020215_, _020216_, _020217_, _020218_, _020219_, _020220_, _020221_, _020222_, _020223_, _020224_, _020225_, _020226_, _020227_, _020228_, _020229_, _020230_, _020231_, _020232_, _020233_, _020234_, _020235_, _020236_, _020237_, _020238_, _020239_, _020240_, _020241_, _020242_, _020243_, _020244_, _020245_, _020246_, _020247_, _020248_, _020249_, _020250_, _020251_, _020252_, _020253_, _020254_, _020255_, _020256_, _020257_, _020258_, _020259_, _020260_, _020261_, _020262_, _020263_, _020264_, _020265_, _020266_, _020267_, _020268_, _020269_, _020270_, _020271_, _020272_, _020273_, _020274_, _020275_, _020276_, _020277_, _020278_, _020279_, _020280_, _020281_, _020282_, _020283_, _020284_, _020285_, _020286_, _020287_, _020288_, _020289_, _020290_, _020291_, _020292_, _020293_, _020294_, _020295_, _020296_, _020297_, _020298_, _020299_, _020300_, _020301_, _020302_, _020303_, _020304_, _020305_, _020306_, _020307_, _020308_, _020309_, _020310_, _020311_, _020312_, _020313_, _020314_, _020315_, _020316_, _020317_, _020318_, _020319_, _020320_, _020321_, _020322_, _020323_, _020324_, _020325_, _020326_, _020327_, _020328_, _020329_, _020330_, _020331_, _020332_, _020333_, _020334_, _020335_, _020336_, _020337_, _020338_, _020339_, _020340_, _020341_, _020342_, _020343_, _020344_, _020345_, _020346_, _020347_, _020348_, _020349_, _020350_, _020351_, _020352_, _020353_, _020354_, _020355_, _020356_, _020357_, _020358_, _020359_, _020360_, _020361_, _020362_, _020363_, _020364_, _020365_, _020366_, _020367_, _020368_, _020369_, _020370_, _020371_, _020372_, _020373_, _020374_, _020375_, _020376_, _020377_, _020378_, _020379_, _020380_, _020381_, _020382_, _020383_, _020384_, _020385_, _020386_, _020387_, _020388_, _020389_, _020390_, _020391_, _020392_, _020393_, _020394_, _020395_, _020396_, _020397_, _020398_, _020399_, _020400_, _020401_, _020402_, _020403_, _020404_, _020405_, _020406_, _020407_, _020408_, _020409_, _020410_, _020411_, _020412_, _020413_, _020414_, _020415_, _020416_, _020417_, _020418_, _020419_, _020420_, _020421_, _020422_, _020423_, _020424_, _020425_, _020426_, _020427_, _020428_, _020429_, _020430_, _020431_, _020432_, _020433_, _020434_, _020435_, _020436_, _020437_, _020438_, _020439_, _020440_, _020441_, _020442_, _020443_, _020444_, _020445_, _020446_, _020447_, _020448_, _020449_, _020450_, _020451_, _020452_, _020453_, _020454_, _020455_, _020456_, _020457_, _020458_, _020459_, _020460_, _020461_, _020462_, _020463_, _020464_, _020465_, _020466_, _020467_, _020468_, _020469_, _020470_, _020471_, _020472_, _020473_, _020474_, _020475_, _020476_, _020477_, _020478_, _020479_, _020480_, _020481_, _020482_, _020483_, _020484_, _020485_, _020486_, _020487_, _020488_, _020489_, _020490_, _020491_, _020492_, _020493_, _020494_, _020495_, _020496_, _020497_, _020498_, _020499_, _020500_, _020501_, _020502_, _020503_, _020504_, _020505_, _020506_, _020507_, _020508_, _020509_, _020510_, _020511_, _020512_, _020513_, _020514_, _020515_, _020516_, _020517_, _020518_, _020519_, _020520_, _020521_, _020522_, _020523_, _020524_, _020525_, _020526_, _020527_, _020528_, _020529_, _020530_, _020531_, _020532_, _020533_, _020534_, _020535_, _020536_, _020537_, _020538_, _020539_, _020540_, _020541_, _020542_, _020543_, _020544_, _020545_, _020546_, _020547_, _020548_, _020549_, _020550_, _020551_, _020552_, _020553_, _020554_, _020555_, _020556_, _020557_, _020558_, _020559_, _020560_, _020561_, _020562_, _020563_, _020564_, _020565_, _020566_, _020567_, _020568_, _020569_, _020570_, _020571_, _020572_, _020573_, _020574_, _020575_, _020576_, _020577_, _020578_, _020579_, _020580_, _020581_, _020582_, _020583_, _020584_, _020585_, _020586_, _020587_, _020588_, _020589_, _020590_, _020591_, _020592_, _020593_, _020594_, _020595_, _020596_, _020597_, _020598_, _020599_, _020600_, _020601_, _020602_, _020603_, _020604_, _020605_, _020606_, _020607_, _020608_, _020609_, _020610_, _020611_, _020612_, _020613_, _020614_, _020615_, _020616_, _020617_, _020618_, _020619_, _020620_, _020621_, _020622_, _020623_, _020624_, _020625_, _020626_, _020627_, _020628_, _020629_, _020630_, _020631_, _020632_, _020633_, _020634_, _020635_, _020636_, _020637_, _020638_, _020639_, _020640_, _020641_, _020642_, _020643_, _020644_, _020645_, _020646_, _020647_, _020648_, _020649_, _020650_, _020651_, _020652_, _020653_, _020654_, _020655_, _020656_, _020657_, _020658_, _020659_, _020660_, _020661_, _020662_, _020663_, _020664_, _020665_, _020666_, _020667_, _020668_, _020669_, _020670_, _020671_, _020672_, _020673_, _020674_, _020675_, _020676_, _020677_, _020678_, _020679_, _020680_, _020681_, _020682_, _020683_, _020684_, _020685_, _020686_, _020687_, _020688_, _020689_, _020690_, _020691_, _020692_, _020693_, _020694_, _020695_, _020696_, _020697_, _020698_, _020699_, _020700_, _020701_, _020702_, _020703_, _020704_, _020705_, _020706_, _020707_, _020708_, _020709_, _020710_, _020711_, _020712_, _020713_, _020714_, _020715_, _020716_, _020717_, _020718_, _020719_, _020720_, _020721_, _020722_, _020723_, _020724_, _020725_, _020726_, _020727_, _020728_, _020729_, _020730_, _020731_, _020732_, _020733_, _020734_, _020735_, _020736_, _020737_, _020738_, _020739_, _020740_, _020741_, _020742_, _020743_, _020744_, _020745_, _020746_, _020747_, _020748_, _020749_, _020750_, _020751_, _020752_, _020753_, _020754_, _020755_, _020756_, _020757_, _020758_, _020759_, _020760_, _020761_, _020762_, _020763_, _020764_, _020765_, _020766_, _020767_, _020768_, _020769_, _020770_, _020771_, _020772_, _020773_, _020774_, _020775_, _020776_, _020777_, _020778_, _020779_, _020780_, _020781_, _020782_, _020783_, _020784_, _020785_, _020786_, _020787_, _020788_, _020789_, _020790_, _020791_, _020792_, _020793_, _020794_, _020795_, _020796_, _020797_, _020798_, _020799_, _020800_, _020801_, _020802_, _020803_, _020804_, _020805_, _020806_, _020807_, _020808_, _020809_, _020810_, _020811_, _020812_, _020813_, _020814_, _020815_, _020816_, _020817_, _020818_, _020819_, _020820_, _020821_, _020822_, _020823_, _020824_, _020825_, _020826_, _020827_, _020828_, _020829_, _020830_, _020831_, _020832_, _020833_, _020834_, _020835_, _020836_, _020837_, _020838_, _020839_, _020840_, _020841_, _020842_, _020843_, _020844_, _020845_, _020846_, _020847_, _020848_, _020849_, _020850_, _020851_, _020852_, _020853_, _020854_, _020855_, _020856_, _020857_, _020858_, _020859_, _020860_, _020861_, _020862_, _020863_, _020864_, _020865_, _020866_, _020867_, _020868_, _020869_, _020870_, _020871_, _020872_, _020873_, _020874_, _020875_, _020876_, _020877_, _020878_, _020879_, _020880_, _020881_, _020882_, _020883_, _020884_, _020885_, _020886_, _020887_, _020888_, _020889_, _020890_, _020891_, _020892_, _020893_, _020894_, _020895_, _020896_, _020897_, _020898_, _020899_, _020900_, _020901_, _020902_, _020903_, _020904_, _020905_, _020906_, _020907_, _020908_, _020909_, _020910_, _020911_, _020912_, _020913_, _020914_, _020915_, _020916_, _020917_, _020918_, _020919_, _020920_, _020921_, _020922_, _020923_, _020924_, _020925_, _020926_, _020927_, _020928_, _020929_, _020930_, _020931_, _020932_, _020933_, _020934_, _020935_, _020936_, _020937_, _020938_, _020939_, _020940_, _020941_, _020942_, _020943_, _020944_, _020945_, _020946_, _020947_, _020948_, _020949_, _020950_, _020951_, _020952_, _020953_, _020954_, _020955_, _020956_, _020957_, _020958_, _020959_, _020960_, _020961_, _020962_, _020963_, _020964_, _020965_, _020966_, _020967_, _020968_, _020969_, _020970_, _020971_, _020972_, _020973_, _020974_, _020975_, _020976_, _020977_, _020978_, _020979_, _020980_, _020981_, _020982_, _020983_, _020984_, _020985_, _020986_, _020987_, _020988_, _020989_, _020990_, _020991_, _020992_, _020993_, _020994_, _020995_, _020996_, _020997_, _020998_, _020999_, _021000_, _021001_, _021002_, _021003_, _021004_, _021005_, _021006_, _021007_, _021008_, _021009_, _021010_, _021011_, _021012_, _021013_, _021014_, _021015_, _021016_, _021017_, _021018_, _021019_, _021020_, _021021_, _021022_, _021023_, _021024_, _021025_, _021026_, _021027_, _021028_, _021029_, _021030_, _021031_, _021032_, _021033_, _021034_, _021035_, _021036_, _021037_, _021038_, _021039_, _021040_, _021041_, _021042_, _021043_, _021044_, _021045_, _021046_, _021047_, _021048_, _021049_, _021050_, _021051_, _021052_, _021053_, _021054_, _021055_, _021056_, _021057_, _021058_, _021059_, _021060_, _021061_, _021062_, _021063_, _021064_, _021065_, _021066_, _021067_, _021068_, _021069_, _021070_, _021071_, _021072_, _021073_, _021074_, _021075_, _021076_, _021077_, _021078_, _021079_, _021080_, _021081_, _021082_, _021083_, _021084_, _021085_, _021086_, _021087_, _021088_, _021089_, _021090_, _021091_, _021092_, _021093_, _021094_, _021095_, _021096_, _021097_, _021098_, _021099_, _021100_, _021101_, _021102_, _021103_, _021104_, _021105_, _021106_, _021107_, _021108_, _021109_, _021110_, _021111_, _021112_, _021113_, _021114_, _021115_, _021116_, _021117_, _021118_, _021119_, _021120_, _021121_, _021122_, _021123_, _021124_, _021125_, _021126_, _021127_, _021128_, _021129_, _021130_, _021131_, _021132_, _021133_, _021134_, _021135_, _021136_, _021137_, _021138_, _021139_, _021140_, _021141_, _021142_, _021143_, _021144_, _021145_, _021146_, _021147_, _021148_, _021149_, _021150_, _021151_, _021152_, _021153_, _021154_, _021155_, _021156_, _021157_, _021158_, _021159_, _021160_, _021161_, _021162_, _021163_, _021164_, _021165_, _021166_, _021167_, _021168_, _021169_, _021170_, _021171_, _021172_, _021173_, _021174_, _021175_, _021176_, _021177_, _021178_, _021179_, _021180_, _021181_, _021182_, _021183_, _021184_, _021185_, _021186_, _021187_, _021188_, _021189_, _021190_, _021191_, _021192_, _021193_, _021194_, _021195_, _021196_, _021197_, _021198_, _021199_, _021200_, _021201_, _021202_, _021203_, _021204_, _021205_, _021206_, _021207_, _021208_, _021209_, _021210_, _021211_, _021212_, _021213_, _021214_, _021215_, _021216_, _021217_, _021218_, _021219_, _021220_, _021221_, _021222_, _021223_, _021224_, _021225_, _021226_, _021227_, _021228_, _021229_, _021230_, _021231_, _021232_, _021233_, _021234_, _021235_, _021236_, _021237_, _021238_, _021239_, _021240_, _021241_, _021242_, _021243_, _021244_, _021245_, _021246_, _021247_, _021248_, _021249_, _021250_, _021251_, _021252_, _021253_, _021254_, _021255_, _021256_, _021257_, _021258_, _021259_, _021260_, _021261_, _021262_, _021263_, _021264_, _021265_, _021266_, _021267_, _021268_, _021269_, _021270_, _021271_, _021272_, _021273_, _021274_, _021275_, _021276_, _021277_, _021278_, _021279_, _021280_, _021281_, _021282_, _021283_, _021284_, _021285_, _021286_, _021287_, _021288_, _021289_, _021290_, _021291_, _021292_, _021293_, _021294_, _021295_, _021296_, _021297_, _021298_, _021299_, _021300_, _021301_, _021302_, _021303_, _021304_, _021305_, _021306_, _021307_, _021308_, _021309_, _021310_, _021311_, _021312_, _021313_, _021314_, _021315_, _021316_, _021317_, _021318_, _021319_, _021320_, _021321_, _021322_, _021323_, _021324_, _021325_, _021326_, _021327_, _021328_, _021329_, _021330_, _021331_, _021332_, _021333_, _021334_, _021335_, _021336_, _021337_, _021338_, _021339_, _021340_, _021341_, _021342_, _021343_, _021344_, _021345_, _021346_, _021347_, _021348_, _021349_, _021350_, _021351_, _021352_, _021353_, _021354_, _021355_, _021356_, _021357_, _021358_, _021359_, _021360_, _021361_, _021362_, _021363_, _021364_, _021365_, _021366_, _021367_, _021368_, _021369_, _021370_, _021371_, _021372_, _021373_, _021374_, _021375_, _021376_, _021377_, _021378_, _021379_, _021380_, _021381_, _021382_, _021383_, _021384_, _021385_, _021386_, _021387_, _021388_, _021389_, _021390_, _021391_, _021392_, _021393_, _021394_, _021395_, _021396_, _021397_, _021398_, _021399_, _021400_, _021401_, _021402_, _021403_, _021404_, _021405_, _021406_, _021407_, _021408_, _021409_, _021410_, _021411_, _021412_, _021413_, _021414_, _021415_, _021416_, _021417_, _021418_, _021419_, _021420_, _021421_, _021422_, _021423_, _021424_, _021425_, _021426_, _021427_, _021428_, _021429_, _021430_, _021431_, _021432_, _021433_, _021434_, _021435_, _021436_, _021437_, _021438_, _021439_, _021440_, _021441_, _021442_, _021443_, _021444_, _021445_, _021446_, _021447_, _021448_, _021449_, _021450_, _021451_, _021452_, _021453_, _021454_, _021455_, _021456_, _021457_, _021458_, _021459_, _021460_, _021461_, _021462_, _021463_, _021464_, _021465_, _021466_, _021467_, _021468_, _021469_, _021470_, _021471_, _021472_, _021473_, _021474_, _021475_, _021476_, _021477_, _021478_, _021479_, _021480_, _021481_, _021482_, _021483_, _021484_, _021485_, _021486_, _021487_, _021488_, _021489_, _021490_, _021491_, _021492_, _021493_, _021494_, _021495_, _021496_, _021497_, _021498_, _021499_, _021500_, _021501_, _021502_, _021503_, _021504_, _021505_, _021506_, _021507_, _021508_, _021509_, _021510_, _021511_, _021512_, _021513_, _021514_, _021515_, _021516_, _021517_, _021518_, _021519_, _021520_, _021521_, _021522_, _021523_, _021524_, _021525_, _021526_, _021527_, _021528_, _021529_, _021530_, _021531_, _021532_, _021533_, _021534_, _021535_, _021536_, _021537_, _021538_, _021539_, _021540_, _021541_, _021542_, _021543_, _021544_, _021545_, _021546_, _021547_, _021548_, _021549_, _021550_, _021551_, _021552_, _021553_, _021554_, _021555_, _021556_, _021557_, _021558_, _021559_, _021560_, _021561_, _021562_, _021563_, _021564_, _021565_, _021566_, _021567_, _021568_, _021569_, _021570_, _021571_, _021572_, _021573_, _021574_, _021575_, _021576_, _021577_, _021578_, _021579_, _021580_, _021581_, _021582_, _021583_, _021584_, _021585_, _021586_, _021587_, _021588_, _021589_, _021590_, _021591_, _021592_, _021593_, _021594_, _021595_, _021596_, _021597_, _021598_, _021599_, _021600_, _021601_, _021602_, _021603_, _021604_, _021605_, _021606_, _021607_, _021608_, _021609_, _021610_, _021611_, _021612_, _021613_, _021614_, _021615_, _021616_, _021617_, _021618_, _021619_, _021620_, _021621_, _021622_, _021623_, _021624_, _021625_, _021626_, _021627_, _021628_, _021629_, _021630_, _021631_, _021632_, _021633_, _021634_, _021635_, _021636_, _021637_, _021638_, _021639_, _021640_, _021641_, _021642_, _021643_, _021644_, _021645_, _021646_, _021647_, _021648_, _021649_, _021650_, _021651_, _021652_, _021653_, _021654_, _021655_, _021656_, _021657_, _021658_, _021659_, _021660_, _021661_, _021662_, _021663_, _021664_, _021665_, _021666_, _021667_, _021668_, _021669_, _021670_, _021671_, _021672_, _021673_, _021674_, _021675_, _021676_, _021677_, _021678_, _021679_, _021680_, _021681_, _021682_, _021683_, _021684_, _021685_, _021686_, _021687_, _021688_, _021689_, _021690_, _021691_, _021692_, _021693_, _021694_, _021695_, _021696_, _021697_, _021698_, _021699_, _021700_, _021701_, _021702_, _021703_, _021704_, _021705_, _021706_, _021707_, _021708_, _021709_, _021710_, _021711_, _021712_, _021713_, _021714_, _021715_, _021716_, _021717_, _021718_, _021719_, _021720_, _021721_, _021722_, _021723_, _021724_, _021725_, _021726_, _021727_, _021728_, _021729_, _021730_, _021731_, _021732_, _021733_, _021734_, _021735_, _021736_, _021737_, _021738_, _021739_, _021740_, _021741_, _021742_, _021743_, _021744_, _021745_, _021746_, _021747_, _021748_, _021749_, _021750_, _021751_, _021752_, _021753_, _021754_, _021755_, _021756_, _021757_, _021758_, _021759_, _021760_, _021761_, _021762_, _021763_, _021764_, _021765_, _021766_, _021767_, _021768_, _021769_, _021770_, _021771_, _021772_, _021773_, _021774_, _021775_, _021776_, _021777_, _021778_, _021779_, _021780_, _021781_, _021782_, _021783_, _021784_, _021785_, _021786_, _021787_, _021788_, _021789_, _021790_, _021791_, _021792_, _021793_, _021794_, _021795_, _021796_, _021797_, _021798_, _021799_, _021800_, _021801_, _021802_, _021803_, _021804_, _021805_, _021806_, _021807_, _021808_, _021809_, _021810_, _021811_, _021812_, _021813_, _021814_, _021815_, _021816_, _021817_, _021818_, _021819_, _021820_, _021821_, _021822_, _021823_, _021824_, _021825_, _021826_, _021827_, _021828_, _021829_, _021830_, _021831_, _021832_, _021833_, _021834_, _021835_, _021836_, _021837_, _021838_, _021839_, _021840_, _021841_, _021842_, _021843_, _021844_, _021845_, _021846_, _021847_, _021848_, _021849_, _021850_, _021851_, _021852_, _021853_, _021854_, _021855_, _021856_, _021857_, _021858_, _021859_, _021860_, _021861_, _021862_, _021863_, _021864_, _021865_, _021866_, _021867_, _021868_, _021869_, _021870_, _021871_, _021872_, _021873_, _021874_, _021875_, _021876_, _021877_, _021878_, _021879_, _021880_, _021881_, _021882_, _021883_, _021884_, _021885_, _021886_, _021887_, _021888_, _021889_, _021890_, _021891_, _021892_, _021893_, _021894_, _021895_, _021896_, _021897_, _021898_, _021899_, _021900_, _021901_, _021902_, _021903_, _021904_, _021905_, _021906_, _021907_, _021908_, _021909_, _021910_, _021911_, _021912_, _021913_, _021914_, _021915_, _021916_, _021917_, _021918_, _021919_, _021920_, _021921_, _021922_, _021923_, _021924_, _021925_, _021926_, _021927_, _021928_, _021929_, _021930_, _021931_, _021932_, _021933_, _021934_, _021935_, _021936_, _021937_, _021938_, _021939_, _021940_, _021941_, _021942_, _021943_, _021944_, _021945_, _021946_, _021947_, _021948_, _021949_, _021950_, _021951_, _021952_, _021953_, _021954_, _021955_, _021956_, _021957_, _021958_, _021959_, _021960_, _021961_, _021962_, _021963_, _021964_, _021965_, _021966_, _021967_, _021968_, _021969_, _021970_, _021971_, _021972_, _021973_, _021974_, _021975_, _021976_, _021977_, _021978_, _021979_, _021980_, _021981_, _021982_, _021983_, _021984_, _021985_, _021986_, _021987_, _021988_, _021989_, _021990_, _021991_, _021992_, _021993_, _021994_, _021995_, _021996_, _021997_, _021998_, _021999_, _022000_, _022001_, _022002_, _022003_, _022004_, _022005_, _022006_, _022007_, _022008_, _022009_, _022010_, _022011_, _022012_, _022013_, _022014_, _022015_, _022016_, _022017_, _022018_, _022019_, _022020_, _022021_, _022022_, _022023_, _022024_, _022025_, _022026_, _022027_, _022028_, _022029_, _022030_, _022031_, _022032_, _022033_, _022034_, _022035_, _022036_, _022037_, _022038_, _022039_, _022040_, _022041_, _022042_, _022043_, _022044_, _022045_, _022046_, _022047_, _022048_, _022049_, _022050_, _022051_, _022052_, _022053_, _022054_, _022055_, _022056_, _022057_, _022058_, _022059_, _022060_, _022061_, _022062_, _022063_, _022064_, _022065_, _022066_, _022067_, _022068_, _022069_, _022070_, _022071_, _022072_, _022073_, _022074_, _022075_, _022076_, _022077_, _022078_, _022079_, _022080_, _022081_, _022082_, _022083_, _022084_, _022085_, _022086_, _022087_, _022088_, _022089_, _022090_, _022091_, _022092_, _022093_, _022094_, _022095_, _022096_, _022097_, _022098_, _022099_, _022100_, _022101_, _022102_, _022103_, _022104_, _022105_, _022106_, _022107_, _022108_, _022109_, _022110_, _022111_, _022112_, _022113_, _022114_, _022115_, _022116_, _022117_, _022118_, _022119_, _022120_, _022121_, _022122_, _022123_, _022124_, _022125_, _022126_, _022127_, _022128_, _022129_, _022130_, _022131_, _022132_, _022133_, _022134_, _022135_, _022136_, _022137_, _022138_, _022139_, _022140_, _022141_, _022142_, _022143_, _022144_, _022145_, _022146_, _022147_, _022148_, _022149_, _022150_, _022151_, _022152_, _022153_, _022154_, _022155_, _022156_, _022157_, _022158_, _022159_, _022160_, _022161_, _022162_, _022163_, _022164_, _022165_, _022166_, _022167_, _022168_, _022169_, _022170_, _022171_, _022172_, _022173_, _022174_, _022175_, _022176_, _022177_, _022178_, _022179_, _022180_, _022181_, _022182_, _022183_, _022184_, _022185_, _022186_, _022187_, _022188_, _022189_, _022190_, _022191_, _022192_, _022193_, _022194_, _022195_, _022196_, _022197_, _022198_, _022199_, _022200_, _022201_, _022202_, _022203_, _022204_, _022205_, _022206_, _022207_, _022208_, _022209_, _022210_, _022211_, _022212_, _022213_, _022214_, _022215_, _022216_, _022217_, _022218_, _022219_, _022220_, _022221_, _022222_, _022223_, _022224_, _022225_, _022226_, _022227_, _022228_, _022229_, _022230_, _022231_, _022232_, _022233_, _022234_, _022235_, _022236_, _022237_, _022238_, _022239_, _022240_, _022241_, _022242_, _022243_, _022244_, _022245_, _022246_, _022247_, _022248_, _022249_, _022250_, _022251_, _022252_, _022253_, _022254_, _022255_, _022256_, _022257_, _022258_, _022259_, _022260_, _022261_, _022262_, _022263_, _022264_, _022265_, _022266_, _022267_, _022268_, _022269_, _022270_, _022271_, _022272_, _022273_, _022274_, _022275_, _022276_, _022277_, _022278_, _022279_, _022280_, _022281_, _022282_, _022283_, _022284_, _022285_, _022286_, _022287_, _022288_, _022289_, _022290_, _022291_, _022292_, _022293_, _022294_, _022295_, _022296_, _022297_, _022298_, _022299_, _022300_, _022301_, _022302_, _022303_, _022304_, _022305_, _022306_, _022307_, _022308_, _022309_, _022310_, _022311_, _022312_, _022313_, _022314_, _022315_, _022316_, _022317_, _022318_, _022319_, _022320_, _022321_, _022322_, _022323_, _022324_, _022325_, _022326_, _022327_, _022328_, _022329_, _022330_, _022331_, _022332_, _022333_, _022334_, _022335_, _022336_, _022337_, _022338_, _022339_, _022340_, _022341_, _022342_, _022343_, _022344_, _022345_, _022346_, _022347_, _022348_, _022349_, _022350_, _022351_, _022352_, _022353_, _022354_, _022355_, _022356_, _022357_, _022358_, _022359_, _022360_, _022361_, _022362_, _022363_, _022364_, _022365_, _022366_, _022367_, _022368_, _022369_, _022370_, _022371_, _022372_, _022373_, _022374_, _022375_, _022376_, _022377_, _022378_, _022379_, _022380_, _022381_, _022382_, _022383_, _022384_, _022385_, _022386_, _022387_, _022388_, _022389_, _022390_, _022391_, _022392_, _022393_, _022394_, _022395_, _022396_, _022397_, _022398_, _022399_, _022400_, _022401_, _022402_, _022403_, _022404_, _022405_, _022406_, _022407_, _022408_, _022409_, _022410_, _022411_, _022412_, _022413_, _022414_, _022415_, _022416_, _022417_, _022418_, _022419_, _022420_, _022421_, _022422_, _022423_, _022424_, _022425_, _022426_, _022427_, _022428_, _022429_, _022430_, _022431_, _022432_, _022433_, _022434_, _022435_, _022436_, _022437_, _022438_, _022439_, _022440_, _022441_, _022442_, _022443_, _022444_, _022445_, _022446_, _022447_, _022448_, _022449_, _022450_, _022451_, _022452_, _022453_, _022454_, _022455_, _022456_, _022457_, _022458_, _022459_, _022460_, _022461_, _022462_, _022463_, _022464_, _022465_, _022466_, _022467_, _022468_, _022469_, _022470_, _022471_, _022472_, _022473_, _022474_, _022475_, _022476_, _022477_, _022478_, _022479_, _022480_, _022481_, _022482_, _022483_, _022484_, _022485_, _022486_, _022487_, _022488_, _022489_, _022490_, _022491_, _022492_, _022493_, _022494_, _022495_, _022496_, _022497_, _022498_, _022499_, _022500_, _022501_, _022502_, _022503_, _022504_, _022505_, _022506_, _022507_, _022508_, _022509_, _022510_, _022511_, _022512_, _022513_, _022514_, _022515_, _022516_, _022517_, _022518_, _022519_, _022520_, _022521_, _022522_, _022523_, _022524_, _022525_, _022526_, _022527_, _022528_, _022529_, _022530_, _022531_, _022532_, _022533_, _022534_, _022535_, _022536_, _022537_, _022538_, _022539_, _022540_, _022541_, _022542_, _022543_, _022544_, _022545_, _022546_, _022547_, _022548_, _022549_, _022550_, _022551_, _022552_, _022553_, _022554_, _022555_, _022556_, _022557_, _022558_, _022559_, _022560_, _022561_, _022562_, _022563_, _022564_, _022565_, _022566_, _022567_, _022568_, _022569_, _022570_, _022571_, _022572_, _022573_, _022574_, _022575_, _022576_, _022577_, _022578_, _022579_, _022580_, _022581_, _022582_, _022583_, _022584_, _022585_, _022586_, _022587_, _022588_, _022589_, _022590_, _022591_, _022592_, _022593_, _022594_, _022595_, _022596_, _022597_, _022598_, _022599_, _022600_, _022601_, _022602_, _022603_, _022604_, _022605_, _022606_, _022607_, _022608_, _022609_, _022610_, _022611_, _022612_, _022613_, _022614_, _022615_, _022616_, _022617_, _022618_, _022619_, _022620_, _022621_, _022622_, _022623_, _022624_, _022625_, _022626_, _022627_, _022628_, _022629_, _022630_, _022631_, _022632_, _022633_, _022634_, _022635_, _022636_, _022637_, _022638_, _022639_, _022640_, _022641_, _022642_, _022643_, _022644_, _022645_, _022646_, _022647_, _022648_, _022649_, _022650_, _022651_, _022652_, _022653_, _022654_, _022655_, _022656_, _022657_, _022658_, _022659_, _022660_, _022661_, _022662_, _022663_, _022664_, _022665_, _022666_, _022667_, _022668_, _022669_, _022670_, _022671_, _022672_, _022673_, _022674_, _022675_, _022676_, _022677_, _022678_, _022679_, _022680_, _022681_, _022682_, _022683_, _022684_, _022685_, _022686_, _022687_, _022688_, _022689_, _022690_, _022691_, _022692_, _022693_, _022694_, _022695_, _022696_, _022697_, _022698_, _022699_, _022700_, _022701_, _022702_, _022703_, _022704_, _022705_, _022706_, _022707_, _022708_, _022709_, _022710_, _022711_, _022712_, _022713_, _022714_, _022715_, _022716_, _022717_, _022718_, _022719_, _022720_, _022721_, _022722_, _022723_, _022724_, _022725_, _022726_, _022727_, _022728_, _022729_, _022730_, _022731_, _022732_, _022733_, _022734_, _022735_, _022736_, _022737_, _022738_, _022739_, _022740_, _022741_, _022742_, _022743_, _022744_, _022745_, _022746_, _022747_, _022748_, _022749_, _022750_, _022751_, _022752_, _022753_, _022754_, _022755_, _022756_, _022757_, _022758_, _022759_, _022760_, _022761_, _022762_, _022763_, _022764_, _022765_, _022766_, _022767_, _022768_, _022769_, _022770_, _022771_, _022772_, _022773_, _022774_, _022775_, _022776_, _022777_, _022778_, _022779_, _022780_, _022781_, _022782_, _022783_, _022784_, _022785_, _022786_, _022787_, _022788_, _022789_, _022790_, _022791_, _022792_, _022793_, _022794_, _022795_, _022796_, _022797_, _022798_, _022799_, _022800_, _022801_, _022802_, _022803_, _022804_, _022805_, _022806_, _022807_, _022808_, _022809_, _022810_, _022811_, _022812_, _022813_, _022814_, _022815_, _022816_, _022817_, _022818_, _022819_, _022820_, _022821_, _022822_, _022823_, _022824_, _022825_, _022826_, _022827_, _022828_, _022829_, _022830_, _022831_, _022832_, _022833_, _022834_, _022835_, _022836_, _022837_, _022838_, _022839_, _022840_, _022841_, _022842_, _022843_, _022844_, _022845_, _022846_, _022847_, _022848_, _022849_, _022850_, _022851_, _022852_, _022853_, _022854_, _022855_, _022856_, _022857_, _022858_, _022859_, _022860_, _022861_, _022862_, _022863_, _022864_, _022865_, _022866_, _022867_, _022868_, _022869_, _022870_, _022871_, _022872_, _022873_, _022874_, _022875_, _022876_, _022877_, _022878_, _022879_, _022880_, _022881_, _022882_, _022883_, _022884_, _022885_, _022886_, _022887_, _022888_, _022889_, _022890_, _022891_, _022892_, _022893_, _022894_, _022895_, _022896_, _022897_, _022898_, _022899_, _022900_, _022901_, _022902_, _022903_, _022904_, _022905_, _022906_, _022907_, _022908_, _022909_, _022910_, _022911_, _022912_, _022913_, _022914_, _022915_, _022916_, _022917_, _022918_, _022919_, _022920_, _022921_, _022922_, _022923_, _022924_, _022925_, _022926_, _022927_, _022928_, _022929_, _022930_, _022931_, _022932_, _022933_, _022934_, _022935_, _022936_, _022937_, _022938_, _022939_, _022940_, _022941_, _022942_, _022943_, _022944_, _022945_, _022946_, _022947_, _022948_, _022949_, _022950_, _022951_, _022952_, _022953_, _022954_, _022955_, _022956_, _022957_, _022958_, _022959_, _022960_, _022961_, _022962_, _022963_, _022964_, _022965_, _022966_, _022967_, _022968_, _022969_, _022970_, _022971_, _022972_, _022973_, _022974_, _022975_, _022976_, _022977_, _022978_, _022979_, _022980_, _022981_, _022982_, _022983_, _022984_, _022985_, _022986_, _022987_, _022988_, _022989_, _022990_, _022991_, _022992_, _022993_, _022994_, _022995_, _022996_, _022997_, _022998_, _022999_, _023000_, _023001_, _023002_, _023003_, _023004_, _023005_, _023006_, _023007_, _023008_, _023009_, _023010_, _023011_, _023012_, _023013_, _023014_, _023015_, _023016_, _023017_, _023018_, _023019_, _023020_, _023021_, _023022_, _023023_, _023024_, _023025_, _023026_, _023027_, _023028_, _023029_, _023030_, _023031_, _023032_, _023033_, _023034_, _023035_, _023036_, _023037_, _023038_, _023039_, _023040_, _023041_, _023042_, _023043_, _023044_, _023045_, _023046_, _023047_, _023048_, _023049_, _023050_, _023051_, _023052_, _023053_, _023054_, _023055_, _023056_, _023057_, _023058_, _023059_, _023060_, _023061_, _023062_, _023063_, _023064_, _023065_, _023066_, _023067_, _023068_, _023069_, _023070_, _023071_, _023072_, _023073_, _023074_, _023075_, _023076_, _023077_, _023078_, _023079_, _023080_, _023081_, _023082_, _023083_, _023084_, _023085_, _023086_, _023087_, _023088_, _023089_, _023090_, _023091_, _023092_, _023093_, _023094_, _023095_, _023096_, _023097_, _023098_, _023099_, _023100_, _023101_, _023102_, _023103_, _023104_, _023105_, _023106_, _023107_, _023108_, _023109_, _023110_, _023111_, _023112_, _023113_, _023114_, _023115_, _023116_, _023117_, _023118_, _023119_, _023120_, _023121_, _023122_, _023123_, _023124_, _023125_, _023126_, _023127_, _023128_, _023129_, _023130_, _023131_, _023132_, _023133_, _023134_, _023135_, _023136_, _023137_, _023138_, _023139_, _023140_, _023141_, _023142_, _023143_, _023144_, _023145_, _023146_, _023147_, _023148_, _023149_, _023150_, _023151_, _023152_, _023153_, _023154_, _023155_, _023156_, _023157_, _023158_, _023159_, _023160_, _023161_, _023162_, _023163_, _023164_, _023165_, _023166_, _023167_, _023168_, _023169_, _023170_, _023171_, _023172_, _023173_, _023174_, _023175_, _023176_, _023177_, _023178_, _023179_, _023180_, _023181_, _023182_, _023183_, _023184_, _023185_, _023186_, _023187_, _023188_, _023189_, _023190_, _023191_, _023192_, _023193_, _023194_, _023195_, _023196_, _023197_, _023198_, _023199_, _023200_, _023201_, _023202_, _023203_, _023204_, _023205_, _023206_, _023207_, _023208_, _023209_, _023210_, _023211_, _023212_, _023213_, _023214_, _023215_, _023216_, _023217_, _023218_, _023219_, _023220_, _023221_, _023222_, _023223_, _023224_, _023225_, _023226_, _023227_, _023228_, _023229_, _023230_, _023231_, _023232_, _023233_, _023234_, _023235_, _023236_, _023237_, _023238_, _023239_, _023240_, _023241_, _023242_, _023243_, _023244_, _023245_, _023246_, _023247_, _023248_, _023249_, _023250_, _023251_, _023252_, _023253_, _023254_, _023255_, _023256_, _023257_, _023258_, _023259_, _023260_, _023261_, _023262_, _023263_, _023264_, _023265_, _023266_, _023267_, _023268_, _023269_, _023270_, _023271_, _023272_, _023273_, _023274_, _023275_, _023276_, _023277_, _023278_, _023279_, _023280_, _023281_, _023282_, _023283_, _023284_, _023285_, _023286_, _023287_, _023288_, _023289_, _023290_, _023291_, _023292_, _023293_, _023294_, _023295_, _023296_, _023297_, _023298_, _023299_, _023300_, _023301_, _023302_, _023303_, _023304_, _023305_, _023306_, _023307_, _023308_, _023309_, _023310_, _023311_, _023312_, _023313_, _023314_, _023315_, _023316_, _023317_, _023318_, _023319_, _023320_, _023321_, _023322_, _023323_, _023324_, _023325_, _023326_, _023327_, _023328_, _023329_, _023330_, _023331_, _023332_, _023333_, _023334_, _023335_, _023336_, _023337_, _023338_, _023339_, _023340_, _023341_, _023342_, _023343_, _023344_, _023345_, _023346_, _023347_, _023348_, _023349_, _023350_, _023351_, _023352_, _023353_, _023354_, _023355_, _023356_, _023357_, _023358_, _023359_, _023360_, _023361_, _023362_, _023363_, _023364_, _023365_, _023366_, _023367_, _023368_, _023369_, _023370_, _023371_, _023372_, _023373_, _023374_, _023375_, _023376_, _023377_, _023378_, _023379_, _023380_, _023381_, _023382_, _023383_, _023384_, _023385_, _023386_, _023387_, _023388_, _023389_, _023390_, _023391_, _023392_, _023393_, _023394_, _023395_, _023396_, _023397_, _023398_, _023399_, _023400_, _023401_, _023402_, _023403_, _023404_, _023405_, _023406_, _023407_, _023408_, _023409_, _023410_, _023411_, _023412_, _023413_, _023414_, _023415_, _023416_, _023417_, _023418_, _023419_, _023420_, _023421_, _023422_, _023423_, _023424_, _023425_, _023426_, _023427_, _023428_, _023429_, _023430_, _023431_, _023432_, _023433_, _023434_, _023435_, _023436_, _023437_, _023438_, _023439_, _023440_, _023441_, _023442_, _023443_, _023444_, _023445_, _023446_, _023447_, _023448_, _023449_, _023450_, _023451_, _023452_, _023453_, _023454_, _023455_, _023456_, _023457_, _023458_, _023459_, _023460_, _023461_, _023462_, _023463_, _023464_, _023465_, _023466_, _023467_, _023468_, _023469_, _023470_, _023471_, _023472_, _023473_, _023474_, _023475_, _023476_, _023477_, _023478_, _023479_, _023480_, _023481_, _023482_, _023483_, _023484_, _023485_, _023486_, _023487_, _023488_, _023489_, _023490_, _023491_, _023492_, _023493_, _023494_, _023495_, _023496_, _023497_, _023498_, _023499_, _023500_, _023501_, _023502_, _023503_, _023504_, _023505_, _023506_, _023507_, _023508_, _023509_, _023510_, _023511_, _023512_, _023513_, _023514_, _023515_, _023516_, _023517_, _023518_, _023519_, _023520_, _023521_, _023522_, _023523_, _023524_, _023525_, _023526_, _023527_, _023528_, _023529_, _023530_, _023531_, _023532_, _023533_, _023534_, _023535_, _023536_, _023537_, _023538_, _023539_, _023540_, _023541_, _023542_, _023543_, _023544_, _023545_, _023546_, _023547_, _023548_, _023549_, _023550_, _023551_, _023552_, _023553_, _023554_, _023555_, _023556_, _023557_, _023558_, _023559_, _023560_, _023561_, _023562_, _023563_, _023564_, _023565_, _023566_, _023567_, _023568_, _023569_, _023570_, _023571_, _023572_, _023573_, _023574_, _023575_, _023576_, _023577_, _023578_, _023579_, _023580_, _023581_, _023582_, _023583_, _023584_, _023585_, _023586_, _023587_, _023588_, _023589_, _023590_, _023591_, _023592_, _023593_, _023594_, _023595_, _023596_, _023597_, _023598_, _023599_, _023600_, _023601_, _023602_, _023603_, _023604_, _023605_, _023606_, _023607_, _023608_, _023609_, _023610_, _023611_, _023612_, _023613_, _023614_, _023615_, _023616_, _023617_, _023618_, _023619_, _023620_, _023621_, _023622_, _023623_, _023624_, _023625_, _023626_, _023627_, _023628_, _023629_, _023630_, _023631_, _023632_, _023633_, _023634_, _023635_, _023636_, _023637_, _023638_, _023639_, _023640_, _023641_, _023642_, _023643_, _023644_, _023645_, _023646_, _023647_, _023648_, _023649_, _023650_, _023651_, _023652_, _023653_, _023654_, _023655_, _023656_, _023657_, _023658_, _023659_, _023660_, _023661_, _023662_, _023663_, _023664_, _023665_, _023666_, _023667_, _023668_, _023669_, _023670_, _023671_, _023672_, _023673_, _023674_, _023675_, _023676_, _023677_, _023678_, _023679_, _023680_, _023681_, _023682_, _023683_, _023684_, _023685_, _023686_, _023687_, _023688_, _023689_, _023690_, _023691_, _023692_, _023693_, _023694_, _023695_, _023696_, _023697_, _023698_, _023699_, _023700_, _023701_, _023702_, _023703_, _023704_, _023705_, _023706_, _023707_, _023708_, _023709_, _023710_, _023711_, _023712_, _023713_, _023714_, _023715_, _023716_, _023717_, _023718_, _023719_, _023720_, _023721_, _023722_, _023723_, _023724_, _023725_, _023726_, _023727_, _023728_, _023729_, _023730_, _023731_, _023732_, _023733_, _023734_, _023735_, _023736_, _023737_, _023738_, _023739_, _023740_, _023741_, _023742_, _023743_, _023744_, _023745_, _023746_, _023747_, _023748_, _023749_, _023750_, _023751_, _023752_, _023753_, _023754_, _023755_, _023756_, _023757_, _023758_, _023759_, _023760_, _023761_, _023762_, _023763_, _023764_, _023765_, _023766_, _023767_, _023768_, _023769_, _023770_, _023771_, _023772_, _023773_, _023774_, _023775_, _023776_, _023777_, _023778_, _023779_, _023780_, _023781_, _023782_, _023783_, _023784_, _023785_, _023786_, _023787_, _023788_, _023789_, _023790_, _023791_, _023792_, _023793_, _023794_, _023795_, _023796_, _023797_, _023798_, _023799_, _023800_, _023801_, _023802_, _023803_, _023804_, _023805_, _023806_, _023807_, _023808_, _023809_, _023810_, _023811_, _023812_, _023813_, _023814_, _023815_, _023816_, _023817_, _023818_, _023819_, _023820_, _023821_, _023822_, _023823_, _023824_, _023825_, _023826_, _023827_, _023828_, _023829_, _023830_, _023831_, _023832_, _023833_, _023834_, _023835_, _023836_, _023837_, _023838_, _023839_, _023840_, _023841_, _023842_, _023843_, _023844_, _023845_, _023846_, _023847_, _023848_, _023849_, _023850_, _023851_, _023852_, _023853_, _023854_, _023855_, _023856_, _023857_, _023858_, _023859_, _023860_, _023861_, _023862_, _023863_, _023864_, _023865_, _023866_, _023867_, _023868_, _023869_, _023870_, _023871_, _023872_, _023873_, _023874_, _023875_, _023876_, _023877_, _023878_, _023879_, _023880_, _023881_, _023882_, _023883_, _023884_, _023885_, _023886_, _023887_, _023888_, _023889_, _023890_, _023891_, _023892_, _023893_, _023894_, _023895_, _023896_, _023897_, _023898_, _023899_, _023900_, _023901_, _023902_, _023903_, _023904_, _023905_, _023906_, _023907_, _023908_, _023909_, _023910_, _023911_, _023912_, _023913_, _023914_, _023915_, _023916_, _023917_, _023918_, _023919_, _023920_, _023921_, _023922_, _023923_, _023924_, _023925_, _023926_, _023927_, _023928_, _023929_, _023930_, _023931_, _023932_, _023933_, _023934_, _023935_, _023936_, _023937_, _023938_, _023939_, _023940_, _023941_, _023942_, _023943_, _023944_, _023945_, _023946_, _023947_, _023948_, _023949_, _023950_, _023951_, _023952_, _023953_, _023954_, _023955_, _023956_, _023957_, _023958_, _023959_, _023960_, _023961_, _023962_, _023963_, _023964_, _023965_, _023966_, _023967_, _023968_, _023969_, _023970_, _023971_, _023972_, _023973_, _023974_, _023975_, _023976_, _023977_, _023978_, _023979_, _023980_, _023981_, _023982_, _023983_, _023984_, _023985_, _023986_, _023987_, _023988_, _023989_, _023990_, _023991_, _023992_, _023993_, _023994_, _023995_, _023996_, _023997_, _023998_, _023999_, _024000_, _024001_, _024002_, _024003_, _024004_, _024005_, _024006_, _024007_, _024008_, _024009_, _024010_, _024011_, _024012_, _024013_, _024014_, _024015_, _024016_, _024017_, _024018_, _024019_, _024020_, _024021_, _024022_, _024023_, _024024_, _024025_, _024026_, _024027_, _024028_, _024029_, _024030_, _024031_, _024032_, _024033_, _024034_, _024035_, _024036_, _024037_, _024038_, _024039_, _024040_, _024041_, _024042_, _024043_, _024044_, _024045_, _024046_, _024047_, _024048_, _024049_, _024050_, _024051_, _024052_, _024053_, _024054_, _024055_, _024056_, _024057_, _024058_, _024059_, _024060_, _024061_, _024062_, _024063_, _024064_, _024065_, _024066_, _024067_, _024068_, _024069_, _024070_, _024071_, _024072_, _024073_, _024074_, _024075_, _024076_, _024077_, _024078_, _024079_, _024080_, _024081_, _024082_, _024083_, _024084_, _024085_, _024086_, _024087_, _024088_, _024089_, _024090_, _024091_, _024092_, _024093_, _024094_, _024095_, _024096_, _024097_, _024098_, _024099_, _024100_, _024101_, _024102_, _024103_, _024104_, _024105_, _024106_, _024107_, _024108_, _024109_, _024110_, _024111_, _024112_, _024113_, _024114_, _024115_, _024116_, _024117_, _024118_, _024119_, _024120_, _024121_, _024122_, _024123_, _024124_, _024125_, _024126_, _024127_, _024128_, _024129_, _024130_, _024131_, _024132_, _024133_, _024134_, _024135_, _024136_, _024137_, _024138_, _024139_, _024140_, _024141_, _024142_, _024143_, _024144_, _024145_, _024146_, _024147_, _024148_, _024149_, _024150_, _024151_, _024152_, _024153_, _024154_, _024155_, _024156_, _024157_, _024158_, _024159_, _024160_, _024161_, _024162_, _024163_, _024164_, _024165_, _024166_, _024167_, _024168_, _024169_, _024170_, _024171_, _024172_, _024173_, _024174_, _024175_, _024176_, _024177_, _024178_, _024179_, _024180_, _024181_, _024182_, _024183_, _024184_, _024185_, _024186_, _024187_, _024188_, _024189_, _024190_, _024191_, _024192_, _024193_, _024194_, _024195_, _024196_, _024197_, _024198_, _024199_, _024200_, _024201_, _024202_, _024203_, _024204_, _024205_, _024206_, _024207_, _024208_, _024209_, _024210_, _024211_, _024212_, _024213_, _024214_, _024215_, _024216_, _024217_, _024218_, _024219_, _024220_, _024221_, _024222_, _024223_, _024224_, _024225_, _024226_, _024227_, _024228_, _024229_, _024230_, _024231_, _024232_, _024233_, _024234_, _024235_, _024236_, _024237_, _024238_, _024239_, _024240_, _024241_, _024242_, _024243_, _024244_, _024245_, _024246_, _024247_, _024248_, _024249_, _024250_, _024251_, _024252_, _024253_, _024254_, _024255_, _024256_, _024257_, _024258_, _024259_, _024260_, _024261_, _024262_, _024263_, _024264_, _024265_, _024266_, _024267_, _024268_, _024269_, _024270_, _024271_, _024272_, _024273_, _024274_, _024275_, _024276_, _024277_, _024278_, _024279_, _024280_, _024281_, _024282_, _024283_, _024284_, _024285_, _024286_, _024287_, _024288_, _024289_, _024290_, _024291_, _024292_, _024293_, _024294_, _024295_, _024296_, _024297_, _024298_, _024299_, _024300_, _024301_, _024302_, _024303_, _024304_, _024305_, _024306_, _024307_, _024308_, _024309_, _024310_, _024311_, _024312_, _024313_, _024314_, _024315_, _024316_, _024317_, _024318_, _024319_, _024320_, _024321_, _024322_, _024323_, _024324_, _024325_, _024326_, _024327_, _024328_, _024329_, _024330_, _024331_, _024332_, _024333_, _024334_, _024335_, _024336_, _024337_, _024338_, _024339_, _024340_, _024341_, _024342_, _024343_, _024344_, _024345_, _024346_, _024347_, _024348_, _024349_, _024350_, _024351_, _024352_, _024353_, _024354_, _024355_, _024356_, _024357_, _024358_, _024359_, _024360_, _024361_, _024362_, _024363_, _024364_, _024365_, _024366_, _024367_, _024368_, _024369_, _024370_, _024371_, _024372_, _024373_, _024374_, _024375_, _024376_, _024377_, _024378_, _024379_, _024380_, _024381_, _024382_, _024383_, _024384_, _024385_, _024386_, _024387_, _024388_, _024389_, _024390_, _024391_, _024392_, _024393_, _024394_, _024395_, _024396_, _024397_, _024398_, _024399_, _024400_, _024401_, _024402_, _024403_, _024404_, _024405_, _024406_, _024407_, _024408_, _024409_, _024410_, _024411_, _024412_, _024413_, _024414_, _024415_, _024416_, _024417_, _024418_, _024419_, _024420_, _024421_, _024422_, _024423_, _024424_, _024425_, _024426_, _024427_, _024428_, _024429_, _024430_, _024431_, _024432_, _024433_, _024434_, _024435_, _024436_, _024437_, _024438_, _024439_, _024440_, _024441_, _024442_, _024443_, _024444_, _024445_, _024446_, _024447_, _024448_, _024449_, _024450_, _024451_, _024452_, _024453_, _024454_, _024455_, _024456_, _024457_, _024458_, _024459_, _024460_, _024461_, _024462_, _024463_, _024464_, _024465_, _024466_, _024467_, _024468_, _024469_, _024470_, _024471_, _024472_, _024473_, _024474_, _024475_, _024476_, _024477_, _024478_, _024479_, _024480_, _024481_, _024482_, _024483_, _024484_, _024485_, _024486_, _024487_, _024488_, _024489_, _024490_, _024491_, _024492_, _024493_, _024494_, _024495_, _024496_, _024497_, _024498_, _024499_, _024500_, _024501_, _024502_, _024503_, _024504_, _024505_, _024506_, _024507_, _024508_, _024509_, _024510_, _024511_, _024512_, _024513_, _024514_, _024515_, _024516_, _024517_, _024518_, _024519_, _024520_, _024521_, _024522_, _024523_, _024524_, _024525_, _024526_, _024527_, _024528_, _024529_, _024530_, _024531_, _024532_, _024533_, _024534_, _024535_, _024536_, _024537_, _024538_, _024539_, _024540_, _024541_, _024542_, _024543_, _024544_, _024545_, _024546_, _024547_, _024548_, _024549_, _024550_, _024551_, _024552_, _024553_, _024554_, _024555_, _024556_, _024557_, _024558_, _024559_, _024560_, _024561_, _024562_, _024563_, _024564_, _024565_, _024566_, _024567_, _024568_, _024569_, _024570_, _024571_, _024572_, _024573_, _024574_, _024575_, _024576_, _024577_, _024578_, _024579_, _024580_, _024581_, _024582_, _024583_, _024584_, _024585_, _024586_, _024587_, _024588_, _024589_, _024590_, _024591_, _024592_, _024593_, _024594_, _024595_, _024596_, _024597_, _024598_, _024599_, _024600_, _024601_, _024602_, _024603_, _024604_, _024605_, _024606_, _024607_, _024608_, _024609_, _024610_, _024611_, _024612_, _024613_, _024614_, _024615_, _024616_, _024617_, _024618_, _024619_, _024620_, _024621_, _024622_, _024623_, _024624_, _024625_, _024626_, _024627_, _024628_, _024629_, _024630_, _024631_, _024632_, _024633_, _024634_, _024635_, _024636_, _024637_, _024638_, _024639_, _024640_, _024641_, _024642_, _024643_, _024644_, _024645_, _024646_, _024647_, _024648_, _024649_, _024650_, _024651_, _024652_, _024653_, _024654_, _024655_, _024656_, _024657_, _024658_, _024659_, _024660_, _024661_, _024662_, _024663_, _024664_, _024665_, _024666_, _024667_, _024668_, _024669_, _024670_, _024671_, _024672_, _024673_, _024674_, _024675_, _024676_, _024677_, _024678_, _024679_, _024680_, _024681_, _024682_, _024683_, _024684_, _024685_, _024686_, _024687_, _024688_, _024689_, _024690_, _024691_, _024692_, _024693_, _024694_, _024695_, _024696_, _024697_, _024698_, _024699_, _024700_, _024701_, _024702_, _024703_, _024704_, _024705_, _024706_, _024707_, _024708_, _024709_, _024710_, _024711_, _024712_, _024713_, _024714_, _024715_, _024716_, _024717_, _024718_, _024719_, _024720_, _024721_, _024722_, _024723_, _024724_, _024725_, _024726_, _024727_, _024728_, _024729_, _024730_, _024731_, _024732_, _024733_, _024734_, _024735_, _024736_, _024737_, _024738_, _024739_, _024740_, _024741_, _024742_, _024743_, _024744_, _024745_, _024746_, _024747_, _024748_, _024749_, _024750_, _024751_, _024752_, _024753_, _024754_, _024755_, _024756_, _024757_, _024758_, _024759_, _024760_, _024761_, _024762_, _024763_, _024764_, _024765_, _024766_, _024767_, _024768_, _024769_, _024770_, _024771_, _024772_, _024773_, _024774_, _024775_, _024776_, _024777_, _024778_, _024779_, _024780_, _024781_, _024782_, _024783_, _024784_, _024785_, _024786_, _024787_, _024788_, _024789_, _024790_, _024791_, _024792_, _024793_, _024794_, _024795_, _024796_, _024797_, _024798_, _024799_, _024800_, _024801_, _024802_, _024803_, _024804_, _024805_, _024806_, _024807_, _024808_, _024809_, _024810_, _024811_, _024812_, _024813_, _024814_, _024815_, _024816_, _024817_, _024818_, _024819_, _024820_, _024821_, _024822_, _024823_, _024824_, _024825_, _024826_, _024827_, _024828_, _024829_, _024830_, _024831_, _024832_, _024833_, _024834_, _024835_, _024836_, _024837_, _024838_, _024839_, _024840_, _024841_, _024842_, _024843_, _024844_, _024845_, _024846_, _024847_, _024848_, _024849_, _024850_, _024851_, _024852_, _024853_, _024854_, _024855_, _024856_, _024857_, _024858_, _024859_, _024860_, _024861_, _024862_, _024863_, _024864_, _024865_, _024866_, _024867_, _024868_, _024869_, _024870_, _024871_, _024872_, _024873_, _024874_, _024875_, _024876_, _024877_, _024878_, _024879_, _024880_, _024881_, _024882_, _024883_, _024884_, _024885_, _024886_, _024887_, _024888_, _024889_, _024890_, _024891_, _024892_, _024893_, _024894_, _024895_, _024896_, _024897_, _024898_, _024899_, _024900_, _024901_, _024902_, _024903_, _024904_, _024905_, _024906_, _024907_, _024908_, _024909_, _024910_, _024911_, _024912_, _024913_, _024914_, _024915_, _024916_, _024917_, _024918_, _024919_, _024920_, _024921_, _024922_, _024923_, _024924_, _024925_, _024926_, _024927_, _024928_, _024929_, _024930_, _024931_, _024932_, _024933_, _024934_, _024935_, _024936_, _024937_, _024938_, _024939_, _024940_, _024941_, _024942_, _024943_, _024944_, _024945_, _024946_, _024947_, _024948_, _024949_, _024950_, _024951_, _024952_, _024953_, _024954_, _024955_, _024956_, _024957_, _024958_, _024959_, _024960_, _024961_, _024962_, _024963_, _024964_, _024965_, _024966_, _024967_, _024968_, _024969_, _024970_, _024971_, _024972_, _024973_, _024974_, _024975_, _024976_, _024977_, _024978_, _024979_, _024980_, _024981_, _024982_, _024983_, _024984_, _024985_, _024986_, _024987_, _024988_, _024989_, _024990_, _024991_, _024992_, _024993_, _024994_, _024995_, _024996_, _024997_, _024998_, _024999_, _025000_, _025001_, _025002_, _025003_, _025004_, _025005_, _025006_, _025007_, _025008_, _025009_, _025010_, _025011_, _025012_, _025013_, _025014_, _025015_, _025016_, _025017_, _025018_, _025019_, _025020_, _025021_, _025022_, _025023_, _025024_, _025025_, _025026_, _025027_, _025028_, _025029_, _025030_, _025031_, _025032_, _025033_, _025034_, _025035_, _025036_, _025037_, _025038_, _025039_, _025040_, _025041_, _025042_, _025043_, _025044_, _025045_, _025046_, _025047_, _025048_, _025049_, _025050_, _025051_, _025052_, _025053_, _025054_, _025055_, _025056_, _025057_, _025058_, _025059_, _025060_, _025061_, _025062_, _025063_, _025064_, _025065_, _025066_, _025067_, _025068_, _025069_, _025070_, _025071_, _025072_, _025073_, _025074_, _025075_, _025076_, _025077_, _025078_, _025079_, _025080_, _025081_, _025082_, _025083_, _025084_, _025085_, _025086_, _025087_, _025088_, _025089_, _025090_, _025091_, _025092_, _025093_, _025094_, _025095_, _025096_, _025097_, _025098_, _025099_, _025100_, _025101_, _025102_, _025103_, _025104_, _025105_, _025106_, _025107_, _025108_, _025109_, _025110_, _025111_, _025112_, _025113_, _025114_, _025115_, _025116_, _025117_, _025118_, _025119_, _025120_, _025121_, _025122_, _025123_, _025124_, _025125_, _025126_, _025127_, _025128_, _025129_, _025130_, _025131_, _025132_, _025133_, _025134_, _025135_, _025136_, _025137_, _025138_, _025139_, _025140_, _025141_, _025142_, _025143_, _025144_, _025145_, _025146_, _025147_, _025148_, _025149_, _025150_, _025151_, _025152_, _025153_, _025154_, _025155_, _025156_, _025157_, _025158_, _025159_, _025160_, _025161_, _025162_, _025163_, _025164_, _025165_, _025166_, _025167_, _025168_, _025169_, _025170_, _025171_, _025172_, _025173_, _025174_, _025175_, _025176_, _025177_, _025178_, _025179_, _025180_, _025181_, _025182_, _025183_, _025184_, _025185_, _025186_, _025187_, _025188_, _025189_, _025190_, _025191_, _025192_, _025193_, _025194_, _025195_, _025196_, _025197_, _025198_, _025199_, _025200_, _025201_, _025202_, _025203_, _025204_, _025205_, _025206_, _025207_, _025208_, _025209_, _025210_, _025211_, _025212_, _025213_, _025214_, _025215_, _025216_, _025217_, _025218_, _025219_, _025220_, _025221_, _025222_, _025223_, _025224_, _025225_, _025226_, _025227_, _025228_, _025229_, _025230_, _025231_, _025232_, _025233_, _025234_, _025235_, _025236_, _025237_, _025238_, _025239_, _025240_, _025241_, _025242_, _025243_, _025244_, _025245_, _025246_, _025247_, _025248_, _025249_, _025250_, _025251_, _025252_, _025253_, _025254_, _025255_, _025256_, _025257_, _025258_, _025259_, _025260_, _025261_, _025262_, _025263_, _025264_, _025265_, _025266_, _025267_, _025268_, _025269_, _025270_, _025271_, _025272_, _025273_, _025274_, _025275_, _025276_, _025277_, _025278_, _025279_, _025280_, _025281_, _025282_, _025283_, _025284_, _025285_, _025286_, _025287_, _025288_, _025289_, _025290_, _025291_, _025292_, _025293_, _025294_, _025295_, _025296_, _025297_, _025298_, _025299_, _025300_, _025301_, _025302_, _025303_, _025304_, _025305_, _025306_, _025307_, _025308_, _025309_, _025310_, _025311_, _025312_, _025313_, _025314_, _025315_, _025316_, _025317_, _025318_, _025319_, _025320_, _025321_, _025322_, _025323_, _025324_, _025325_, _025326_, _025327_, _025328_, _025329_, _025330_, _025331_, _025332_, _025333_, _025334_, _025335_, _025336_, _025337_, _025338_, _025339_, _025340_, _025341_, _025342_, _025343_, _025344_, _025345_, _025346_, _025347_, _025348_, _025349_, _025350_, _025351_, _025352_, _025353_, _025354_, _025355_, _025356_, _025357_, _025358_, _025359_, _025360_, _025361_, _025362_, _025363_, _025364_, _025365_, _025366_, _025367_, _025368_, _025369_, _025370_, _025371_, _025372_, _025373_, _025374_, _025375_, _025376_, _025377_, _025378_, _025379_, _025380_, _025381_, _025382_, _025383_, _025384_, _025385_, _025386_, _025387_, _025388_, _025389_, _025390_, _025391_, _025392_, _025393_, _025394_, _025395_, _025396_, _025397_, _025398_, _025399_, _025400_, _025401_, _025402_, _025403_, _025404_, _025405_, _025406_, _025407_, _025408_, _025409_, _025410_, _025411_, _025412_, _025413_, _025414_, _025415_, _025416_, _025417_, _025418_, _025419_, _025420_, _025421_, _025422_, _025423_, _025424_, _025425_, _025426_, _025427_, _025428_, _025429_, _025430_, _025431_, _025432_, _025433_, _025434_, _025435_, _025436_, _025437_, _025438_, _025439_, _025440_, _025441_, _025442_, _025443_, _025444_, _025445_, _025446_, _025447_, _025448_, _025449_, _025450_, _025451_, _025452_, _025453_, _025454_, _025455_, _025456_, _025457_, _025458_, _025459_, _025460_, _025461_, _025462_, _025463_, _025464_, _025465_, _025466_, _025467_, _025468_, _025469_, _025470_, _025471_, _025472_, _025473_, _025474_, _025475_, _025476_, _025477_, _025478_, _025479_, _025480_, _025481_, _025482_, _025483_, _025484_, _025485_, _025486_, _025487_, _025488_, _025489_, _025490_, _025491_, _025492_, _025493_, _025494_, _025495_, _025496_, _025497_, _025498_, _025499_, _025500_, _025501_, _025502_, _025503_, _025504_, _025505_, _025506_, _025507_, _025508_, _025509_, _025510_, _025511_, _025512_, _025513_, _025514_, _025515_, _025516_, _025517_, _025518_, _025519_, _025520_, _025521_, _025522_, _025523_, _025524_, _025525_, _025526_, _025527_, _025528_, _025529_, _025530_, _025531_, _025532_, _025533_, _025534_, _025535_, _025536_, _025537_, _025538_, _025539_, _025540_, _025541_, _025542_, _025543_, _025544_, _025545_, _025546_, _025547_, _025548_, _025549_, _025550_, _025551_, _025552_, _025553_, _025554_, _025555_, _025556_, _025557_, _025558_, _025559_, _025560_, _025561_, _025562_, _025563_, _025564_, _025565_, _025566_, _025567_, _025568_, _025569_, _025570_, _025571_, _025572_, _025573_, _025574_, _025575_, _025576_, _025577_, _025578_, _025579_, _025580_, _025581_, _025582_, _025583_, _025584_, _025585_, _025586_, _025587_, _025588_, _025589_, _025590_, _025591_, _025592_, _025593_, _025594_, _025595_, _025596_, _025597_, _025598_, _025599_, _025600_, _025601_, _025602_, _025603_, _025604_, _025605_, _025606_, _025607_, _025608_, _025609_, _025610_, _025611_, _025612_, _025613_, _025614_, _025615_, _025616_, _025617_, _025618_, _025619_, _025620_, _025621_, _025622_, _025623_, _025624_, _025625_, _025626_, _025627_, _025628_, _025629_, _025630_, _025631_, _025632_, _025633_, _025634_, _025635_, _025636_, _025637_, _025638_, _025639_, _025640_, _025641_, _025642_, _025643_, _025644_, _025645_, _025646_, _025647_, _025648_, _025649_, _025650_, _025651_, _025652_, _025653_, _025654_, _025655_, _025656_, _025657_, _025658_, _025659_, _025660_, _025661_, _025662_, _025663_, _025664_, _025665_, _025666_, _025667_, _025668_, _025669_, _025670_, _025671_, _025672_, _025673_, _025674_, _025675_, _025676_, _025677_, _025678_, _025679_, _025680_, _025681_, _025682_, _025683_, _025684_, _025685_, _025686_, _025687_, _025688_, _025689_, _025690_, _025691_, _025692_, _025693_, _025694_, _025695_, _025696_, _025697_, _025698_, _025699_, _025700_, _025701_, _025702_, _025703_, _025704_, _025705_, _025706_, _025707_, _025708_, _025709_, _025710_, _025711_, _025712_, _025713_, _025714_, _025715_, _025716_, _025717_, _025718_, _025719_, _025720_, _025721_, _025722_, _025723_, _025724_, _025725_, _025726_, _025727_, _025728_, _025729_, _025730_, _025731_, _025732_, _025733_, _025734_, _025735_, _025736_, _025737_, _025738_, _025739_, _025740_, _025741_, _025742_, _025743_, _025744_, _025745_, _025746_, _025747_, _025748_, _025749_, _025750_, _025751_, _025752_, _025753_, _025754_, _025755_, _025756_, _025757_, _025758_, _025759_, _025760_, _025761_, _025762_, _025763_, _025764_, _025765_, _025766_, _025767_, _025768_, _025769_, _025770_, _025771_, _025772_, _025773_, _025774_, _025775_, _025776_, _025777_, _025778_, _025779_, _025780_, _025781_, _025782_, _025783_, _025784_, _025785_, _025786_, _025787_, _025788_, _025789_, _025790_, _025791_, _025792_, _025793_, _025794_, _025795_, _025796_, _025797_, _025798_, _025799_, _025800_, _025801_, _025802_, _025803_, _025804_, _025805_, _025806_, _025807_, _025808_, _025809_, _025810_, _025811_, _025812_, _025813_, _025814_, _025815_, _025816_, _025817_, _025818_, _025819_, _025820_, _025821_, _025822_, _025823_, _025824_, _025825_, _025826_, _025827_, _025828_, _025829_, _025830_, _025831_, _025832_, _025833_, _025834_, _025835_, _025836_, _025837_, _025838_, _025839_, _025840_, _025841_, _025842_, _025843_, _025844_, _025845_, _025846_, _025847_, _025848_, _025849_, _025850_, _025851_, _025852_, _025853_, _025854_, _025855_, _025856_, _025857_, _025858_, _025859_, _025860_, _025861_, _025862_, _025863_, _025864_, _025865_, _025866_, _025867_, _025868_, _025869_, _025870_, _025871_, _025872_, _025873_, _025874_, _025875_, _025876_, _025877_, _025878_, _025879_, _025880_, _025881_, _025882_, _025883_, _025884_, _025885_, _025886_, _025887_, _025888_, _025889_, _025890_, _025891_, _025892_, _025893_, _025894_, _025895_, _025896_, _025897_, _025898_, _025899_, _025900_, _025901_, _025902_, _025903_, _025904_, _025905_, _025906_, _025907_, _025908_, _025909_, _025910_, _025911_, _025912_, _025913_, _025914_, _025915_, _025916_, _025917_, _025918_, _025919_, _025920_, _025921_, _025922_, _025923_, _025924_, _025925_, _025926_, _025927_, _025928_, _025929_, _025930_, _025931_, _025932_, _025933_, _025934_, _025935_, _025936_, _025937_, _025938_, _025939_, _025940_, _025941_, _025942_, _025943_, _025944_, _025945_, _025946_, _025947_, _025948_, _025949_, _025950_, _025951_, _025952_, _025953_, _025954_, _025955_, _025956_, _025957_, _025958_, _025959_, _025960_, _025961_, _025962_, _025963_, _025964_, _025965_, _025966_, _025967_, _025968_, _025969_, _025970_, _025971_, _025972_, _025973_, _025974_, _025975_, _025976_, _025977_, _025978_, _025979_, _025980_, _025981_, _025982_, _025983_, _025984_, _025985_, _025986_, _025987_, _025988_, _025989_, _025990_, _025991_, _025992_, _025993_, _025994_, _025995_, _025996_, _025997_, _025998_, _025999_, _026000_, _026001_, _026002_, _026003_, _026004_, _026005_, _026006_, _026007_, _026008_, _026009_, _026010_, _026011_, _026012_, _026013_, _026014_, _026015_, _026016_, _026017_, _026018_, _026019_, _026020_, _026021_, _026022_, _026023_, _026024_, _026025_, _026026_, _026027_, _026028_, _026029_, _026030_, _026031_, _026032_, _026033_, _026034_, _026035_, _026036_, _026037_, _026038_, _026039_, _026040_, _026041_, _026042_, _026043_, _026044_, _026045_, _026046_, _026047_, _026048_, _026049_, _026050_, _026051_, _026052_, _026053_, _026054_, _026055_, _026056_, _026057_, _026058_, _026059_, _026060_, _026061_, _026062_, _026063_, _026064_, _026065_, _026066_, _026067_, _026068_, _026069_, _026070_, _026071_, _026072_, _026073_, _026074_, _026075_, _026076_, _026077_, _026078_, _026079_, _026080_, _026081_, _026082_, _026083_, _026084_, _026085_, _026086_, _026087_, _026088_, _026089_, _026090_, _026091_, _026092_, _026093_, _026094_, _026095_, _026096_, _026097_, _026098_, _026099_, _026100_, _026101_, _026102_, _026103_, _026104_, _026105_, _026106_, _026107_, _026108_, _026109_, _026110_, _026111_, _026112_, _026113_, _026114_, _026115_, _026116_, _026117_, _026118_, _026119_, _026120_, _026121_, _026122_, _026123_, _026124_, _026125_, _026126_, _026127_, _026128_, _026129_, _026130_, _026131_, _026132_, _026133_, _026134_, _026135_, _026136_, _026137_, _026138_, _026139_, _026140_, _026141_, _026142_, _026143_, _026144_, _026145_, _026146_, _026147_, _026148_, _026149_, _026150_, _026151_, _026152_, _026153_, _026154_, _026155_, _026156_, _026157_, _026158_, _026159_, _026160_, _026161_, _026162_, _026163_, _026164_, _026165_, _026166_, _026167_, _026168_, _026169_, _026170_, _026171_, _026172_, _026173_, _026174_, _026175_, _026176_, _026177_, _026178_, _026179_, _026180_, _026181_, _026182_, _026183_, _026184_, _026185_, _026186_, _026187_, _026188_, _026189_, _026190_, _026191_, _026192_, _026193_, _026194_, _026195_, _026196_, _026197_, _026198_, _026199_, _026200_, _026201_, _026202_, _026203_, _026204_, _026205_, _026206_, _026207_, _026208_, _026209_, _026210_, _026211_, _026212_, _026213_, _026214_, _026215_, _026216_, _026217_, _026218_, _026219_, _026220_, _026221_, _026222_, _026223_, _026224_, _026225_, _026226_, _026227_, _026228_, _026229_, _026230_, _026231_, _026232_, _026233_, _026234_, _026235_, _026236_, _026237_, _026238_, _026239_, _026240_, _026241_, _026242_, _026243_, _026244_, _026245_, _026246_, _026247_, _026248_, _026249_, _026250_, _026251_, _026252_, _026253_, _026254_, _026255_, _026256_, _026257_, _026258_, _026259_, _026260_, _026261_, _026262_, _026263_, _026264_, _026265_, _026266_, _026267_, _026268_, _026269_, _026270_, _026271_, _026272_, _026273_, _026274_, _026275_, _026276_, _026277_, _026278_, _026279_, _026280_, _026281_, _026282_, _026283_, _026284_, _026285_, _026286_, _026287_, _026288_, _026289_, _026290_, _026291_, _026292_, _026293_, _026294_, _026295_, _026296_, _026297_, _026298_, _026299_, _026300_, _026301_, _026302_, _026303_, _026304_, _026305_, _026306_, _026307_, _026308_, _026309_, _026310_, _026311_, _026312_, _026313_, _026314_, _026315_, _026316_, _026317_, _026318_, _026319_, _026320_, _026321_, _026322_, _026323_, _026324_, _026325_, _026326_, _026327_, _026328_, _026329_, _026330_, _026331_, _026332_, _026333_, _026334_, _026335_, _026336_, _026337_, _026338_, _026339_, _026340_, _026341_, _026342_, _026343_, _026344_, _026345_, _026346_, _026347_, _026348_, _026349_, _026350_, _026351_, _026352_, _026353_, _026354_, _026355_, _026356_, _026357_, _026358_, _026359_, _026360_, _026361_, _026362_, _026363_, _026364_, _026365_, _026366_, _026367_, _026368_, _026369_, _026370_, _026371_, _026372_, _026373_, _026374_, _026375_, _026376_, _026377_, _026378_, _026379_, _026380_, _026381_, _026382_, _026383_, _026384_, _026385_, _026386_, _026387_, _026388_, _026389_, _026390_, _026391_, _026392_, _026393_, _026394_, _026395_, _026396_, _026397_, _026398_, _026399_, _026400_, _026401_, _026402_, _026403_, _026404_, _026405_, _026406_, _026407_, _026408_, _026409_, _026410_, _026411_, _026412_, _026413_, _026414_, _026415_, _026416_, _026417_, _026418_, _026419_, _026420_, _026421_, _026422_, _026423_, _026424_, _026425_, _026426_, _026427_, _026428_, _026429_, _026430_, _026431_, _026432_, _026433_, _026434_, _026435_, _026436_, _026437_, _026438_, _026439_, _026440_, _026441_, _026442_, _026443_, _026444_, _026445_, _026446_, _026447_, _026448_, _026449_, _026450_, _026451_, _026452_, _026453_, _026454_, _026455_, _026456_, _026457_, _026458_, _026459_, _026460_, _026461_, _026462_, _026463_, _026464_, _026465_, _026466_, _026467_, _026468_, _026469_, _026470_, _026471_, _026472_, _026473_, _026474_, _026475_, _026476_, _026477_, _026478_, _026479_, _026480_, _026481_, _026482_, _026483_, _026484_, _026485_, _026486_, _026487_, _026488_, _026489_, _026490_, _026491_, _026492_, _026493_, _026494_, _026495_, _026496_, _026497_, _026498_, _026499_, _026500_, _026501_, _026502_, _026503_, _026504_, _026505_, _026506_, _026507_, _026508_, _026509_, _026510_, _026511_, _026512_, _026513_, _026514_, _026515_, _026516_, _026517_, _026518_, _026519_, _026520_, _026521_, _026522_, _026523_, _026524_, _026525_, _026526_, _026527_, _026528_, _026529_, _026530_, _026531_, _026532_, _026533_, _026534_, _026535_, _026536_, _026537_, _026538_, _026539_, _026540_, _026541_, _026542_, _026543_, _026544_, _026545_, _026546_, _026547_, _026548_, _026549_, _026550_, _026551_, _026552_, _026553_, _026554_, _026555_, _026556_, _026557_, _026558_, _026559_, _026560_, _026561_, _026562_, _026563_, _026564_, _026565_, _026566_, _026567_, _026568_, _026569_, _026570_, _026571_, _026572_, _026573_, _026574_, _026575_, _026576_, _026577_, _026578_, _026579_, _026580_, _026581_, _026582_, _026583_, _026584_, _026585_, _026586_, _026587_, _026588_, _026589_, _026590_, _026591_, _026592_, _026593_, _026594_, _026595_, _026596_, _026597_, _026598_, _026599_, _026600_, _026601_, _026602_, _026603_, _026604_, _026605_, _026606_, _026607_, _026608_, _026609_, _026610_, _026611_, _026612_, _026613_, _026614_, _026615_, _026616_, _026617_, _026618_, _026619_, _026620_, _026621_, _026622_, _026623_, _026624_, _026625_, _026626_, _026627_, _026628_, _026629_, _026630_, _026631_, _026632_, _026633_, _026634_, _026635_, _026636_, _026637_, _026638_, _026639_, _026640_, _026641_, _026642_, _026643_, _026644_, _026645_, _026646_, _026647_, _026648_, _026649_, _026650_, _026651_, _026652_, _026653_, _026654_, _026655_, _026656_, _026657_, _026658_, _026659_, _026660_, _026661_, _026662_, _026663_, _026664_, _026665_, _026666_, _026667_, _026668_, _026669_, _026670_, _026671_, _026672_, _026673_, _026674_, _026675_, _026676_, _026677_, _026678_, _026679_, _026680_, _026681_, _026682_, _026683_, _026684_, _026685_, _026686_, _026687_, _026688_, _026689_, _026690_, _026691_, _026692_, _026693_, _026694_, _026695_, _026696_, _026697_, _026698_, _026699_, _026700_, _026701_, _026702_, _026703_, _026704_, _026705_, _026706_, _026707_, _026708_, _026709_, _026710_, _026711_, _026712_, _026713_, _026714_, _026715_, _026716_, _026717_, _026718_, _026719_, _026720_, _026721_, _026722_, _026723_, _026724_, _026725_, _026726_, _026727_, _026728_, _026729_, _026730_, _026731_, _026732_, _026733_, _026734_, _026735_, _026736_, _026737_, _026738_, _026739_, _026740_, _026741_, _026742_, _026743_, _026744_, _026745_, _026746_, _026747_, _026748_, _026749_, _026750_, _026751_, _026752_, _026753_, _026754_, _026755_, _026756_, _026757_, _026758_, _026759_, _026760_, _026761_, _026762_, _026763_, _026764_, _026765_, _026766_, _026767_, _026768_, _026769_, _026770_, _026771_, _026772_, _026773_, _026774_, _026775_, _026776_, _026777_, _026778_, _026779_, _026780_, _026781_, _026782_, _026783_, _026784_, _026785_, _026786_, _026787_, _026788_, _026789_, _026790_, _026791_, _026792_, _026793_, _026794_, _026795_, _026796_, _026797_, _026798_, _026799_, _026800_, _026801_, _026802_, _026803_, _026804_, _026805_, _026806_, _026807_, _026808_, _026809_, _026810_, _026811_, _026812_, _026813_, _026814_, _026815_, _026816_, _026817_, _026818_, _026819_, _026820_, _026821_, _026822_, _026823_, _026824_, _026825_, _026826_, _026827_, _026828_, _026829_, _026830_, _026831_, _026832_, _026833_, _026834_, _026835_, _026836_, _026837_, _026838_, _026839_, _026840_, _026841_, _026842_, _026843_, _026844_, _026845_, _026846_, _026847_, _026848_, _026849_, _026850_, _026851_, _026852_, _026853_, _026854_, _026855_, _026856_, _026857_, _026858_, _026859_, _026860_, _026861_, _026862_, _026863_, _026864_, _026865_, _026866_, _026867_, _026868_, _026869_, _026870_, _026871_, _026872_, _026873_, _026874_, _026875_, _026876_, _026877_, _026878_, _026879_, _026880_, _026881_, _026882_, _026883_, _026884_, _026885_, _026886_, _026887_, _026888_, _026889_, _026890_, _026891_, _026892_, _026893_, _026894_, _026895_, _026896_, _026897_, _026898_, _026899_, _026900_, _026901_, _026902_, _026903_, _026904_, _026905_, _026906_, _026907_, _026908_, _026909_, _026910_, _026911_, _026912_, _026913_, _026914_, _026915_, _026916_, _026917_, _026918_, _026919_, _026920_, _026921_, _026922_, _026923_, _026924_, _026925_, _026926_, _026927_, _026928_, _026929_, _026930_, _026931_, _026932_, _026933_, _026934_, _026935_, _026936_, _026937_, _026938_, _026939_, _026940_, _026941_, _026942_, _026943_, _026944_, _026945_, _026946_, _026947_, _026948_, _026949_, _026950_, _026951_, _026952_, _026953_, _026954_, _026955_, _026956_, _026957_, _026958_, _026959_, _026960_, _026961_, _026962_, _026963_, _026964_, _026965_, _026966_, _026967_, _026968_, _026969_, _026970_, _026971_, _026972_, _026973_, _026974_, _026975_, _026976_, _026977_, _026978_, _026979_, _026980_, _026981_, _026982_, _026983_, _026984_, _026985_, _026986_, _026987_, _026988_, _026989_, _026990_, _026991_, _026992_, _026993_, _026994_, _026995_, _026996_, _026997_, _026998_, _026999_, _027000_, _027001_, _027002_, _027003_, _027004_, _027005_, _027006_, _027007_, _027008_, _027009_, _027010_, _027011_, _027012_, _027013_, _027014_, _027015_, _027016_, _027017_, _027018_, _027019_, _027020_, _027021_, _027022_, _027023_, _027024_, _027025_, _027026_, _027027_, _027028_, _027029_, _027030_, _027031_, _027032_, _027033_, _027034_, _027035_, _027036_, _027037_, _027038_, _027039_, _027040_, _027041_, _027042_, _027043_, _027044_, _027045_, _027046_, _027047_, _027048_, _027049_, _027050_, _027051_, _027052_, _027053_, _027054_, _027055_, _027056_, _027057_, _027058_, _027059_, _027060_, _027061_, _027062_, _027063_, _027064_, _027065_, _027066_, _027067_, _027068_, _027069_, _027070_, _027071_, _027072_, _027073_, _027074_, _027075_, _027076_, _027077_, _027078_, _027079_, _027080_, _027081_, _027082_, _027083_, _027084_, _027085_, _027086_, _027087_, _027088_, _027089_, _027090_, _027091_, _027092_, _027093_, _027094_, _027095_, _027096_, _027097_, _027098_, _027099_, _027100_, _027101_, _027102_, _027103_, _027104_, _027105_, _027106_, _027107_, _027108_, _027109_, _027110_, _027111_, _027112_, _027113_, _027114_, _027115_, _027116_, _027117_, _027118_, _027119_, _027120_, _027121_, _027122_, _027123_, _027124_, _027125_, _027126_, _027127_, _027128_, _027129_, _027130_, _027131_, _027132_, _027133_, _027134_, _027135_, _027136_, _027137_, _027138_, _027139_, _027140_, _027141_, _027142_, _027143_, _027144_, _027145_, _027146_, _027147_, _027148_, _027149_, _027150_, _027151_, _027152_, _027153_, _027154_, _027155_, _027156_, _027157_, _027158_, _027159_, _027160_, _027161_, _027162_, _027163_, _027164_, _027165_, _027166_, _027167_, _027168_, _027169_, _027170_, _027171_, _027172_, _027173_, _027174_, _027175_, _027176_, _027177_, _027178_, _027179_, _027180_, _027181_, _027182_, _027183_, _027184_, _027185_, _027186_, _027187_, _027188_, _027189_, _027190_, _027191_, _027192_, _027193_, _027194_, _027195_, _027196_, _027197_, _027198_, _027199_, _027200_, _027201_, _027202_, _027203_, _027204_, _027205_, _027206_, _027207_, _027208_, _027209_, _027210_, _027211_, _027212_, _027213_, _027214_, _027215_, _027216_, _027217_, _027218_, _027219_, _027220_, _027221_, _027222_, _027223_, _027224_, _027225_, _027226_, _027227_, _027228_, _027229_, _027230_, _027231_, _027232_, _027233_, _027234_, _027235_, _027236_, _027237_, _027238_, _027239_, _027240_, _027241_, _027242_, _027243_, _027244_, _027245_, _027246_, _027247_, _027248_, _027249_, _027250_, _027251_, _027252_, _027253_, _027254_, _027255_, _027256_, _027257_, _027258_, _027259_, _027260_, _027261_, _027262_, _027263_, _027264_, _027265_, _027266_, _027267_, _027268_, _027269_, _027270_, _027271_, _027272_, _027273_, _027274_, _027275_, _027276_, _027277_, _027278_, _027279_, _027280_, _027281_, _027282_, _027283_, _027284_, _027285_, _027286_, _027287_, _027288_, _027289_, _027290_, _027291_, _027292_, _027293_, _027294_, _027295_, _027296_, _027297_, _027298_, _027299_, _027300_, _027301_, _027302_, _027303_, _027304_, _027305_, _027306_, _027307_, _027308_, _027309_, _027310_, _027311_, _027312_, _027313_, _027314_, _027315_, _027316_, _027317_, _027318_, _027319_, _027320_, _027321_, _027322_, _027323_, _027324_, _027325_, _027326_, _027327_, _027328_, _027329_, _027330_, _027331_, _027332_, _027333_, _027334_, _027335_, _027336_, _027337_, _027338_, _027339_, _027340_, _027341_, _027342_, _027343_, _027344_, _027345_, _027346_, _027347_, _027348_, _027349_, _027350_, _027351_, _027352_, _027353_, _027354_, _027355_, _027356_, _027357_, _027358_, _027359_, _027360_, _027361_, _027362_, _027363_, _027364_, _027365_, _027366_, _027367_, _027368_, _027369_, _027370_, _027371_, _027372_, _027373_, _027374_, _027375_, _027376_, _027377_, _027378_, _027379_, _027380_, _027381_, _027382_, _027383_, _027384_, _027385_, _027386_, _027387_, _027388_, _027389_, _027390_, _027391_, _027392_, _027393_, _027394_, _027395_, _027396_, _027397_, _027398_, _027399_, _027400_, _027401_, _027402_, _027403_, _027404_, _027405_, _027406_, _027407_, _027408_, _027409_, _027410_, _027411_, _027412_, _027413_, _027414_, _027415_, _027416_, _027417_, _027418_, _027419_, _027420_, _027421_, _027422_, _027423_, _027424_, _027425_, _027426_, _027427_, _027428_, _027429_, _027430_, _027431_, _027432_, _027433_, _027434_, _027435_, _027436_, _027437_, _027438_, _027439_, _027440_, _027441_, _027442_, _027443_, _027444_, _027445_, _027446_, _027447_, _027448_, _027449_, _027450_, _027451_, _027452_, _027453_, _027454_, _027455_, _027456_, _027457_, _027458_, _027459_, _027460_, _027461_, _027462_, _027463_, _027464_, _027465_, _027466_, _027467_, _027468_, _027469_, _027470_, _027471_, _027472_, _027473_, _027474_, _027475_, _027476_, _027477_, _027478_, _027479_, _027480_, _027481_, _027482_, _027483_, _027484_, _027485_, _027486_, _027487_, _027488_, _027489_, _027490_, _027491_, _027492_, _027493_, _027494_, _027495_, _027496_, _027497_, _027498_, _027499_, _027500_, _027501_, _027502_, _027503_, _027504_, _027505_, _027506_, _027507_, _027508_, _027509_, _027510_, _027511_, _027512_, _027513_, _027514_, _027515_, _027516_, _027517_, _027518_, _027519_, _027520_, _027521_, _027522_, _027523_, _027524_, _027525_, _027526_, _027527_, _027528_, _027529_, _027530_, _027531_, _027532_, _027533_, _027534_, _027535_, _027536_, _027537_, _027538_, _027539_, _027540_, _027541_, _027542_, _027543_, _027544_, _027545_, _027546_, _027547_, _027548_, _027549_, _027550_, _027551_, _027552_, _027553_, _027554_, _027555_, _027556_, _027557_, _027558_, _027559_, _027560_, _027561_, _027562_, _027563_, _027564_, _027565_, _027566_, _027567_, _027568_, _027569_, _027570_, _027571_, _027572_, _027573_, _027574_, _027575_, _027576_, _027577_, _027578_, _027579_, _027580_, _027581_, _027582_, _027583_, _027584_, _027585_, _027586_, _027587_, _027588_, _027589_, _027590_, _027591_, _027592_, _027593_, _027594_, _027595_, _027596_, _027597_, _027598_, _027599_, _027600_, _027601_, _027602_, _027603_, _027604_, _027605_, _027606_, _027607_, _027608_, _027609_, _027610_, _027611_, _027612_, _027613_, _027614_, _027615_, _027616_, _027617_, _027618_, _027619_, _027620_, _027621_, _027622_, _027623_, _027624_, _027625_, _027626_, _027627_, _027628_, _027629_, _027630_, _027631_, _027632_, _027633_, _027634_, _027635_, _027636_, _027637_, _027638_, _027639_, _027640_, _027641_, _027642_, _027643_, _027644_, _027645_, _027646_, _027647_, _027648_, _027649_, _027650_, _027651_, _027652_, _027653_, _027654_, _027655_, _027656_, _027657_, _027658_, _027659_, _027660_, _027661_, _027662_, _027663_, _027664_, _027665_, _027666_, _027667_, _027668_, _027669_, _027670_, _027671_, _027672_, _027673_, _027674_, _027675_, _027676_, _027677_, _027678_, _027679_, _027680_, _027681_, _027682_, _027683_, _027684_, _027685_, _027686_, _027687_, _027688_, _027689_, _027690_, _027691_, _027692_, _027693_, _027694_, _027695_, _027696_, _027697_, _027698_, _027699_, _027700_, _027701_, _027702_, _027703_, _027704_, _027705_, _027706_, _027707_, _027708_, _027709_, _027710_, _027711_, _027712_, _027713_, _027714_, _027715_, _027716_, _027717_, _027718_, _027719_, _027720_, _027721_, _027722_, _027723_, _027724_, _027725_, _027726_, _027727_, _027728_, _027729_, _027730_, _027731_, _027732_, _027733_, _027734_, _027735_, _027736_, _027737_, _027738_, _027739_, _027740_, _027741_, _027742_, _027743_, _027744_, _027745_, _027746_, _027747_, _027748_, _027749_, _027750_, _027751_, _027752_, _027753_, _027754_, _027755_, _027756_, _027757_, _027758_, _027759_, _027760_, _027761_, _027762_, _027763_, _027764_, _027765_, _027766_, _027767_, _027768_, _027769_, _027770_, _027771_, _027772_, _027773_, _027774_, _027775_, _027776_, _027777_, _027778_, _027779_, _027780_, _027781_, _027782_, _027783_, _027784_, _027785_, _027786_, _027787_, _027788_, _027789_, _027790_, _027791_, _027792_, _027793_, _027794_, _027795_, _027796_, _027797_, _027798_, _027799_, _027800_, _027801_, _027802_, _027803_, _027804_, _027805_, _027806_, _027807_, _027808_, _027809_, _027810_, _027811_, _027812_, _027813_, _027814_, _027815_, _027816_, _027817_, _027818_, _027819_, _027820_, _027821_, _027822_, _027823_, _027824_, _027825_, _027826_, _027827_, _027828_, _027829_, _027830_, _027831_, _027832_, _027833_, _027834_, _027835_, _027836_, _027837_, _027838_, _027839_, _027840_, _027841_, _027842_, _027843_, _027844_, _027845_, _027846_, _027847_, _027848_, _027849_, _027850_, _027851_, _027852_, _027853_, _027854_, _027855_, _027856_, _027857_, _027858_, _027859_, _027860_, _027861_, _027862_, _027863_, _027864_, _027865_, _027866_, _027867_, _027868_, _027869_, _027870_, _027871_, _027872_, _027873_, _027874_, _027875_, _027876_, _027877_, _027878_, _027879_, _027880_, _027881_, _027882_, _027883_, _027884_, _027885_, _027886_, _027887_, _027888_, _027889_, _027890_, _027891_, _027892_, _027893_, _027894_, _027895_, _027896_, _027897_, _027898_, _027899_, _027900_, _027901_, _027902_, _027903_, _027904_, _027905_, _027906_, _027907_, _027908_, _027909_, _027910_, _027911_, _027912_, _027913_, _027914_, _027915_, _027916_, _027917_, _027918_, _027919_, _027920_, _027921_, _027922_, _027923_, _027924_, _027925_, _027926_, _027927_, _027928_, _027929_, _027930_, _027931_, _027932_, _027933_, _027934_, _027935_, _027936_, _027937_, _027938_, _027939_, _027940_, _027941_, _027942_, _027943_, _027944_, _027945_, _027946_, _027947_, _027948_, _027949_, _027950_, _027951_, _027952_, _027953_, _027954_, _027955_, _027956_, _027957_, _027958_, _027959_, _027960_, _027961_, _027962_, _027963_, _027964_, _027965_, _027966_, _027967_, _027968_, _027969_, _027970_, _027971_, _027972_, _027973_, _027974_, _027975_, _027976_, _027977_, _027978_, _027979_, _027980_, _027981_, _027982_, _027983_, _027984_, _027985_, _027986_, _027987_, _027988_, _027989_, _027990_, _027991_, _027992_, _027993_, _027994_, _027995_, _027996_, _027997_, _027998_, _027999_, _028000_, _028001_, _028002_, _028003_, _028004_, _028005_, _028006_, _028007_, _028008_, _028009_, _028010_, _028011_, _028012_, _028013_, _028014_, _028015_, _028016_, _028017_, _028018_, _028019_, _028020_, _028021_, _028022_, _028023_, _028024_, _028025_, _028026_, _028027_, _028028_, _028029_, _028030_, _028031_, _028032_, _028033_, _028034_, _028035_, _028036_, _028037_, _028038_, _028039_, _028040_, _028041_, _028042_, _028043_, _028044_, _028045_, _028046_, _028047_, _028048_, _028049_, _028050_, _028051_, _028052_, _028053_, _028054_, _028055_, _028056_, _028057_, _028058_, _028059_, _028060_, _028061_, _028062_, _028063_, _028064_, _028065_, _028066_, _028067_, _028068_, _028069_, _028070_, _028071_, _028072_, _028073_, _028074_, _028075_, _028076_, _028077_, _028078_, _028079_, _028080_, _028081_, _028082_, _028083_, _028084_, _028085_, _028086_, _028087_, _028088_, _028089_, _028090_, _028091_, _028092_, _028093_, _028094_, _028095_, _028096_, _028097_, _028098_, _028099_, _028100_, _028101_, _028102_, _028103_, _028104_, _028105_, _028106_, _028107_, _028108_, _028109_, _028110_, _028111_, _028112_, _028113_, _028114_, _028115_, _028116_, _028117_, _028118_, _028119_, _028120_, _028121_, _028122_, _028123_, _028124_, _028125_, _028126_, _028127_, _028128_, _028129_, _028130_, _028131_, _028132_, _028133_, _028134_, _028135_, _028136_, _028137_, _028138_, _028139_, _028140_, _028141_, _028142_, _028143_, _028144_, _028145_, _028146_, _028147_, _028148_, _028149_, _028150_, _028151_, _028152_, _028153_, _028154_, _028155_, _028156_, _028157_, _028158_, _028159_, _028160_, _028161_, _028162_, _028163_, _028164_, _028165_, _028166_, _028167_, _028168_, _028169_, _028170_, _028171_, _028172_, _028173_, _028174_, _028175_, _028176_, _028177_, _028178_, _028179_, _028180_, _028181_, _028182_, _028183_, _028184_, _028185_, _028186_, _028187_, _028188_, _028189_, _028190_, _028191_, _028192_, _028193_, _028194_, _028195_, _028196_, _028197_, _028198_, _028199_, _028200_, _028201_, _028202_, _028203_, _028204_, _028205_, _028206_, _028207_, _028208_, _028209_, _028210_, _028211_, _028212_, _028213_, _028214_, _028215_, _028216_, _028217_, _028218_, _028219_, _028220_, _028221_, _028222_, _028223_, _028224_, _028225_, _028226_, _028227_, _028228_, _028229_, _028230_, _028231_, _028232_, _028233_, _028234_, _028235_, _028236_, _028237_, _028238_, _028239_, _028240_, _028241_, _028242_, _028243_, _028244_, _028245_, _028246_, _028247_, _028248_, _028249_, _028250_, _028251_, _028252_, _028253_, _028254_, _028255_, _028256_, _028257_, _028258_, _028259_, _028260_, _028261_, _028262_, _028263_, _028264_, _028265_, _028266_, _028267_, _028268_, _028269_, _028270_, _028271_, _028272_, _028273_, _028274_, _028275_, _028276_, _028277_, _028278_, _028279_, _028280_, _028281_, _028282_, _028283_, _028284_, _028285_, _028286_, _028287_, _028288_, _028289_, _028290_, _028291_, _028292_, _028293_, _028294_, _028295_, _028296_, _028297_, _028298_, _028299_, _028300_, _028301_, _028302_, _028303_, _028304_, _028305_, _028306_, _028307_, _028308_, _028309_, _028310_, _028311_, _028312_, _028313_, _028314_, _028315_, _028316_, _028317_, _028318_, _028319_, _028320_, _028321_, _028322_, _028323_, _028324_, _028325_, _028326_, _028327_, _028328_, _028329_, _028330_, _028331_, _028332_, _028333_, _028334_, _028335_, _028336_, _028337_, _028338_, _028339_, _028340_, _028341_, _028342_, _028343_, _028344_, _028345_, _028346_, _028347_, _028348_, _028349_, _028350_, _028351_, _028352_, _028353_, _028354_, _028355_, _028356_, _028357_, _028358_, _028359_, _028360_, _028361_, _028362_, _028363_, _028364_, _028365_, _028366_, _028367_, _028368_, _028369_, _028370_, _028371_, _028372_, _028373_, _028374_, _028375_, _028376_, _028377_, _028378_, _028379_, _028380_, _028381_, _028382_, _028383_, _028384_, _028385_, _028386_, _028387_, _028388_, _028389_, _028390_, _028391_, _028392_, _028393_, _028394_, _028395_, _028396_, _028397_, _028398_, _028399_, _028400_, _028401_, _028402_, _028403_, _028404_, _028405_, _028406_, _028407_, _028408_, _028409_, _028410_, _028411_, _028412_, _028413_, _028414_, _028415_, _028416_, _028417_, _028418_, _028419_, _028420_, _028421_, _028422_, _028423_, _028424_, _028425_, _028426_, _028427_, _028428_, _028429_, _028430_, _028431_, _028432_, _028433_, _028434_, _028435_, _028436_, _028437_, _028438_, _028439_, _028440_, _028441_, _028442_, _028443_, _028444_, _028445_, _028446_, _028447_, _028448_, _028449_, _028450_, _028451_, _028452_, _028453_, _028454_, _028455_, _028456_, _028457_, _028458_, _028459_, _028460_, _028461_, _028462_, _028463_, _028464_, _028465_, _028466_, _028467_, _028468_, _028469_, _028470_, _028471_, _028472_, _028473_, _028474_, _028475_, _028476_, _028477_, _028478_, _028479_, _028480_, _028481_, _028482_, _028483_, _028484_, _028485_, _028486_, _028487_, _028488_, _028489_, _028490_, _028491_, _028492_, _028493_, _028494_, _028495_, _028496_, _028497_, _028498_, _028499_, _028500_, _028501_, _028502_, _028503_, _028504_, _028505_, _028506_, _028507_, _028508_, _028509_, _028510_, _028511_, _028512_, _028513_, _028514_, _028515_, _028516_, _028517_, _028518_, _028519_, _028520_, _028521_, _028522_, _028523_, _028524_, _028525_, _028526_, _028527_, _028528_, _028529_, _028530_, _028531_, _028532_, _028533_, _028534_, _028535_, _028536_, _028537_, _028538_, _028539_, _028540_, _028541_, _028542_, _028543_, _028544_, _028545_, _028546_, _028547_, _028548_, _028549_, _028550_, _028551_, _028552_, _028553_, _028554_, _028555_, _028556_, _028557_, _028558_, _028559_, _028560_, _028561_, _028562_, _028563_, _028564_, _028565_, _028566_, _028567_, _028568_, _028569_, _028570_, _028571_, _028572_, _028573_, _028574_, _028575_, _028576_, _028577_, _028578_, _028579_, _028580_, _028581_, _028582_, _028583_, _028584_, _028585_, _028586_, _028587_, _028588_, _028589_, _028590_, _028591_, _028592_, _028593_, _028594_, _028595_, _028596_, _028597_, _028598_, _028599_, _028600_, _028601_, _028602_, _028603_, _028604_, _028605_, _028606_, _028607_, _028608_, _028609_, _028610_, _028611_, _028612_, _028613_, _028614_, _028615_, _028616_, _028617_, _028618_, _028619_, _028620_, _028621_, _028622_, _028623_, _028624_, _028625_, _028626_, _028627_, _028628_, _028629_, _028630_, _028631_, _028632_, _028633_, _028634_, _028635_, _028636_, _028637_, _028638_, _028639_, _028640_, _028641_, _028642_, _028643_, _028644_, _028645_, _028646_, _028647_, _028648_, _028649_, _028650_, _028651_, _028652_, _028653_, _028654_, _028655_, _028656_, _028657_, _028658_, _028659_, _028660_, _028661_, _028662_, _028663_, _028664_, _028665_, _028666_, _028667_, _028668_, _028669_, _028670_, _028671_, _028672_, _028673_, _028674_, _028675_, _028676_, _028677_, _028678_, _028679_, _028680_, _028681_, _028682_, _028683_, _028684_, _028685_, _028686_, _028687_, _028688_, _028689_, _028690_, _028691_, _028692_, _028693_, _028694_, _028695_, _028696_, _028697_, _028698_, _028699_, _028700_, _028701_, _028702_, _028703_, _028704_, _028705_, _028706_, _028707_, _028708_, _028709_, _028710_, _028711_, _028712_, _028713_, _028714_, _028715_, _028716_, _028717_, _028718_, _028719_, _028720_, _028721_, _028722_, _028723_, _028724_, _028725_, _028726_, _028727_, _028728_, _028729_, _028730_, _028731_, _028732_, _028733_, _028734_, _028735_, _028736_, _028737_, _028738_, _028739_, _028740_, _028741_, _028742_, _028743_, _028744_, _028745_, _028746_, _028747_, _028748_, _028749_, _028750_, _028751_, _028752_, _028753_, _028754_, _028755_, _028756_, _028757_, _028758_, _028759_, _028760_, _028761_, _028762_, _028763_, _028764_, _028765_, _028766_, _028767_, _028768_, _028769_, _028770_, _028771_, _028772_, _028773_, _028774_, _028775_, _028776_, _028777_, _028778_, _028779_, _028780_, _028781_, _028782_, _028783_, _028784_, _028785_, _028786_, _028787_, _028788_, _028789_, _028790_, _028791_, _028792_, _028793_, _028794_, _028795_, _028796_, _028797_, _028798_, _028799_, _028800_, _028801_, _028802_, _028803_, _028804_, _028805_, _028806_, _028807_, _028808_, _028809_, _028810_, _028811_, _028812_, _028813_, _028814_, _028815_, _028816_, _028817_, _028818_, _028819_, _028820_, _028821_, _028822_, _028823_, _028824_, _028825_, _028826_, _028827_, _028828_, _028829_, _028830_, _028831_, _028832_, _028833_, _028834_, _028835_, _028836_, _028837_, _028838_, _028839_, _028840_, _028841_, _028842_, _028843_, _028844_, _028845_, _028846_, _028847_, _028848_, _028849_, _028850_, _028851_, _028852_, _028853_, _028854_, _028855_, _028856_, _028857_, _028858_, _028859_, _028860_, _028861_, _028862_, _028863_, _028864_, _028865_, _028866_, _028867_, _028868_, _028869_, _028870_, _028871_, _028872_, _028873_, _028874_, _028875_, _028876_, _028877_, _028878_, _028879_, _028880_, _028881_, _028882_, _028883_, _028884_, _028885_, _028886_, _028887_, _028888_, _028889_, _028890_, _028891_, _028892_, _028893_, _028894_, _028895_, _028896_, _028897_, _028898_, _028899_, _028900_, _028901_, _028902_, _028903_, _028904_, _028905_, _028906_, _028907_, _028908_, _028909_, _028910_, _028911_, _028912_, _028913_, _028914_, _028915_, _028916_, _028917_, _028918_, _028919_, _028920_, _028921_, _028922_, _028923_, _028924_, _028925_, _028926_, _028927_, _028928_, _028929_, _028930_, _028931_, _028932_, _028933_, _028934_, _028935_, _028936_, _028937_, _028938_, _028939_, _028940_, _028941_, _028942_, _028943_, _028944_, _028945_, _028946_, _028947_, _028948_, _028949_, _028950_, _028951_, _028952_, _028953_, _028954_, _028955_, _028956_, _028957_, _028958_, _028959_, _028960_, _028961_, _028962_, _028963_, _028964_, _028965_, _028966_, _028967_, _028968_, _028969_, _028970_, _028971_, _028972_, _028973_, _028974_, _028975_, _028976_, _028977_, _028978_, _028979_, _028980_, _028981_, _028982_, _028983_, _028984_, _028985_, _028986_, _028987_, _028988_, _028989_, _028990_, _028991_, _028992_, _028993_, _028994_, _028995_, _028996_, _028997_, _028998_, _028999_, _029000_, _029001_, _029002_, _029003_, _029004_, _029005_, _029006_, _029007_, _029008_, _029009_, _029010_, _029011_, _029012_, _029013_, _029014_, _029015_, _029016_, _029017_, _029018_, _029019_, _029020_, _029021_, _029022_, _029023_, _029024_, _029025_, _029026_, _029027_, _029028_, _029029_, _029030_, _029031_, _029032_, _029033_, _029034_, _029035_, _029036_, _029037_, _029038_, _029039_, _029040_, _029041_, _029042_, _029043_, _029044_, _029045_, _029046_, _029047_, _029048_, _029049_, _029050_, _029051_, _029052_, _029053_, _029054_, _029055_, _029056_, _029057_, _029058_, _029059_, _029060_, _029061_, _029062_, _029063_, _029064_, _029065_, _029066_, _029067_, _029068_, _029069_, _029070_, _029071_, _029072_, _029073_, _029074_, _029075_, _029076_, _029077_, _029078_, _029079_, _029080_, _029081_, _029082_, _029083_, _029084_, _029085_, _029086_, _029087_, _029088_, _029089_, _029090_, _029091_, _029092_, _029093_, _029094_, _029095_, _029096_, _029097_, _029098_, _029099_, _029100_, _029101_, _029102_, _029103_, _029104_, _029105_, _029106_, _029107_, _029108_, _029109_, _029110_, _029111_, _029112_, _029113_, _029114_, _029115_, _029116_, _029117_, _029118_, _029119_, _029120_, _029121_, _029122_, _029123_, _029124_, _029125_, _029126_, _029127_, _029128_, _029129_, _029130_, _029131_, _029132_, _029133_, _029134_, _029135_, _029136_, _029137_, _029138_, _029139_, _029140_, _029141_, _029142_, _029143_, _029144_, _029145_, _029146_, _029147_, _029148_, _029149_, _029150_, _029151_, _029152_, _029153_, _029154_, _029155_, _029156_, _029157_, _029158_, _029159_, _029160_, _029161_, _029162_, _029163_, _029164_, _029165_, _029166_, _029167_, _029168_, _029169_, _029170_, _029171_, _029172_, _029173_, _029174_, _029175_, _029176_, _029177_, _029178_, _029179_, _029180_, _029181_, _029182_, _029183_, _029184_, _029185_, _029186_, _029187_, _029188_, _029189_, _029190_, _029191_, _029192_, _029193_, _029194_, _029195_, _029196_, _029197_, _029198_, _029199_, _029200_, _029201_, _029202_, _029203_, _029204_, _029205_, _029206_, _029207_, _029208_, _029209_, _029210_, _029211_, _029212_, _029213_, _029214_, _029215_, _029216_, _029217_, _029218_, _029219_, _029220_, _029221_, _029222_, _029223_, _029224_, _029225_, _029226_, _029227_, _029228_, _029229_, _029230_, _029231_, _029232_, _029233_, _029234_, _029235_, _029236_, _029237_, _029238_, _029239_, _029240_, _029241_, _029242_, _029243_, _029244_, _029245_, _029246_, _029247_, _029248_, _029249_, _029250_, _029251_, _029252_, _029253_, _029254_, _029255_, _029256_, _029257_, _029258_, _029259_, _029260_, _029261_, _029262_, _029263_, _029264_, _029265_, _029266_, _029267_, _029268_, _029269_, _029270_, _029271_, _029272_, _029273_, _029274_, _029275_, _029276_, _029277_, _029278_, _029279_, _029280_, _029281_, _029282_, _029283_, _029284_, _029285_, _029286_, _029287_, _029288_, _029289_, _029290_, _029291_, _029292_, _029293_, _029294_, _029295_, _029296_, _029297_, _029298_, _029299_, _029300_, _029301_, _029302_, _029303_, _029304_, _029305_, _029306_, _029307_, _029308_, _029309_, _029310_, _029311_, _029312_, _029313_, _029314_, _029315_, _029316_, _029317_, _029318_, _029319_, _029320_, _029321_, _029322_, _029323_, _029324_, _029325_, _029326_, _029327_, _029328_, _029329_, _029330_, _029331_, _029332_, _029333_, _029334_, _029335_, _029336_, _029337_, _029338_, _029339_, _029340_, _029341_, _029342_, _029343_, _029344_, _029345_, _029346_, _029347_, _029348_, _029349_, _029350_, _029351_, _029352_, _029353_, _029354_, _029355_, _029356_, _029357_, _029358_, _029359_, _029360_, _029361_, _029362_, _029363_, _029364_, _029365_, _029366_, _029367_, _029368_, _029369_, _029370_, _029371_, _029372_, _029373_, _029374_, _029375_, _029376_, _029377_, _029378_, _029379_, _029380_, _029381_, _029382_, _029383_, _029384_, _029385_, _029386_, _029387_, _029388_, _029389_, _029390_, _029391_, _029392_, _029393_, _029394_, _029395_, _029396_, _029397_, _029398_, _029399_, _029400_, _029401_, _029402_, _029403_, _029404_, _029405_, _029406_, _029407_, _029408_, _029409_, _029410_, _029411_, _029412_, _029413_, _029414_, _029415_, _029416_, _029417_, _029418_, _029419_, _029420_, _029421_, _029422_, _029423_, _029424_, _029425_, _029426_, _029427_, _029428_, _029429_, _029430_, _029431_, _029432_, _029433_, _029434_, _029435_, _029436_, _029437_, _029438_, _029439_, _029440_, _029441_, _029442_, _029443_, _029444_, _029445_, _029446_, _029447_, _029448_, _029449_, _029450_, _029451_, _029452_, _029453_, _029454_, _029455_, _029456_, _029457_, _029458_, _029459_, _029460_, _029461_, _029462_, _029463_, _029464_, _029465_, _029466_, _029467_, _029468_, _029469_, _029470_, _029471_, _029472_, _029473_, _029474_, _029475_, _029476_, _029477_, _029478_, _029479_, _029480_, _029481_, _029482_, _029483_, _029484_, _029485_, _029486_, _029487_, _029488_, _029489_, _029490_, _029491_, _029492_, _029493_, _029494_, _029495_, _029496_, _029497_, _029498_, _029499_, _029500_, _029501_, _029502_, _029503_, _029504_, _029505_, _029506_, _029507_, _029508_, _029509_, _029510_, _029511_, _029512_, _029513_, _029514_, _029515_, _029516_, _029517_, _029518_, _029519_, _029520_, _029521_, _029522_, _029523_, _029524_, _029525_, _029526_, _029527_, _029528_, _029529_, _029530_, _029531_, _029532_, _029533_, _029534_, _029535_, _029536_, _029537_, _029538_, _029539_, _029540_, _029541_, _029542_, _029543_, _029544_, _029545_, _029546_, _029547_, _029548_, _029549_, _029550_, _029551_, _029552_, _029553_, _029554_, _029555_, _029556_, _029557_, _029558_, _029559_, _029560_, _029561_, _029562_, _029563_, _029564_, _029565_, _029566_, _029567_, _029568_, _029569_, _029570_, _029571_, _029572_, _029573_, _029574_, _029575_, _029576_, _029577_, _029578_, _029579_, _029580_, _029581_, _029582_, _029583_, _029584_, _029585_, _029586_, _029587_, _029588_, _029589_, _029590_, _029591_, _029592_, _029593_, _029594_, _029595_, _029596_, _029597_, _029598_, _029599_, _029600_, _029601_, _029602_, _029603_, _029604_, _029605_, _029606_, _029607_, _029608_, _029609_, _029610_, _029611_, _029612_, _029613_, _029614_, _029615_, _029616_, _029617_, _029618_, _029619_, _029620_, _029621_, _029622_, _029623_, _029624_, _029625_, _029626_, _029627_, _029628_, _029629_, _029630_, _029631_, _029632_, _029633_, _029634_, _029635_, _029636_, _029637_, _029638_, _029639_, _029640_, _029641_, _029642_, _029643_, _029644_, _029645_, _029646_, _029647_, _029648_, _029649_, _029650_, _029651_, _029652_, _029653_, _029654_, _029655_, _029656_, _029657_, _029658_, _029659_, _029660_, _029661_, _029662_, _029663_, _029664_, _029665_, _029666_, _029667_, _029668_, _029669_, _029670_, _029671_, _029672_, _029673_, _029674_, _029675_, _029676_, _029677_, _029678_, _029679_, _029680_, _029681_, _029682_, _029683_, _029684_, _029685_, _029686_, _029687_, _029688_, _029689_, _029690_, _029691_, _029692_, _029693_, _029694_, _029695_, _029696_, _029697_, _029698_, _029699_, _029700_, _029701_, _029702_, _029703_, _029704_, _029705_, _029706_, _029707_, _029708_, _029709_, _029710_, _029711_, _029712_, _029713_, _029714_, _029715_, _029716_, _029717_, _029718_, _029719_, _029720_, _029721_, _029722_, _029723_, _029724_, _029725_, _029726_, _029727_, _029728_, _029729_, _029730_, _029731_, _029732_, _029733_, _029734_, _029735_, _029736_, _029737_, _029738_, _029739_, _029740_, _029741_, _029742_, _029743_, _029744_, _029745_, _029746_, _029747_, _029748_, _029749_, _029750_, _029751_, _029752_, _029753_, _029754_, _029755_, _029756_, _029757_, _029758_, _029759_, _029760_, _029761_, _029762_, _029763_, _029764_, _029765_, _029766_, _029767_, _029768_, _029769_, _029770_, _029771_, _029772_, _029773_, _029774_, _029775_, _029776_, _029777_, _029778_, _029779_, _029780_, _029781_, _029782_, _029783_, _029784_, _029785_, _029786_, _029787_, _029788_, _029789_, _029790_, _029791_, _029792_, _029793_, _029794_, _029795_, _029796_, _029797_, _029798_, _029799_, _029800_, _029801_, _029802_, _029803_, _029804_, _029805_, _029806_, _029807_, _029808_, _029809_, _029810_, _029811_, _029812_, _029813_, _029814_, _029815_, _029816_, _029817_, _029818_, _029819_, _029820_, _029821_, _029822_, _029823_, _029824_, _029825_, _029826_, _029827_, _029828_, _029829_, _029830_, _029831_, _029832_, _029833_, _029834_, _029835_, _029836_, _029837_, _029838_, _029839_, _029840_, _029841_, _029842_, _029843_, _029844_, _029845_, _029846_, _029847_, _029848_, _029849_, _029850_, _029851_, _029852_, _029853_, _029854_, _029855_, _029856_, _029857_, _029858_, _029859_, _029860_, _029861_, _029862_, _029863_, _029864_, _029865_, _029866_, _029867_, _029868_, _029869_, _029870_, _029871_, _029872_, _029873_, _029874_, _029875_, _029876_, _029877_, _029878_, _029879_, _029880_, _029881_, _029882_, _029883_, _029884_, _029885_, _029886_, _029887_, _029888_, _029889_, _029890_, _029891_, _029892_, _029893_, _029894_, _029895_, _029896_, _029897_, _029898_, _029899_, _029900_, _029901_, _029902_, _029903_, _029904_, _029905_, _029906_, _029907_, _029908_, _029909_, _029910_, _029911_, _029912_, _029913_, _029914_, _029915_, _029916_, _029917_, _029918_, _029919_, _029920_, _029921_, _029922_, _029923_, _029924_, _029925_, _029926_, _029927_, _029928_, _029929_, _029930_, _029931_, _029932_, _029933_, _029934_, _029935_, _029936_, _029937_, _029938_, _029939_, _029940_, _029941_, _029942_, _029943_, _029944_, _029945_, _029946_, _029947_, _029948_, _029949_, _029950_, _029951_, _029952_, _029953_, _029954_, _029955_, _029956_, _029957_, _029958_, _029959_, _029960_, _029961_, _029962_, _029963_, _029964_, _029965_, _029966_, _029967_, _029968_, _029969_, _029970_, _029971_, _029972_, _029973_, _029974_, _029975_, _029976_, _029977_, _029978_, _029979_, _029980_, _029981_, _029982_, _029983_, _029984_, _029985_, _029986_, _029987_, _029988_, _029989_, _029990_, _029991_, _029992_, _029993_, _029994_, _029995_, _029996_, _029997_, _029998_, _029999_, _030000_, _030001_, _030002_, _030003_, _030004_, _030005_, _030006_, _030007_, _030008_, _030009_, _030010_, _030011_, _030012_, _030013_, _030014_, _030015_, _030016_, _030017_, _030018_, _030019_, _030020_, _030021_, _030022_, _030023_, _030024_, _030025_, _030026_, _030027_, _030028_, _030029_, _030030_, _030031_, _030032_, _030033_, _030034_, _030035_, _030036_, _030037_, _030038_, _030039_, _030040_, _030041_, _030042_, _030043_, _030044_, _030045_, _030046_, _030047_, _030048_, _030049_, _030050_, _030051_, _030052_, _030053_, _030054_, _030055_, _030056_, _030057_, _030058_, _030059_, _030060_, _030061_, _030062_, _030063_, _030064_, _030065_, _030066_, _030067_, _030068_, _030069_, _030070_, _030071_, _030072_, _030073_, _030074_, _030075_, _030076_, _030077_, _030078_, _030079_, _030080_, _030081_, _030082_, _030083_, _030084_, _030085_, _030086_, _030087_, _030088_, _030089_, _030090_, _030091_, _030092_, _030093_, _030094_, _030095_, _030096_, _030097_, _030098_, _030099_, _030100_, _030101_, _030102_, _030103_, _030104_, _030105_, _030106_, _030107_, _030108_, _030109_, _030110_, _030111_, _030112_, _030113_, _030114_, _030115_, _030116_, _030117_, _030118_, _030119_, _030120_, _030121_, _030122_, _030123_, _030124_, _030125_, _030126_, _030127_, _030128_, _030129_, _030130_, _030131_, _030132_, _030133_, _030134_, _030135_, _030136_, _030137_, _030138_, _030139_, _030140_, _030141_, _030142_, _030143_, _030144_, _030145_, _030146_, _030147_, _030148_, _030149_, _030150_, _030151_, _030152_, _030153_, _030154_, _030155_, _030156_, _030157_, _030158_, _030159_, _030160_, _030161_, _030162_, _030163_, _030164_, _030165_, _030166_, _030167_, _030168_, _030169_, _030170_, _030171_, _030172_, _030173_, _030174_, _030175_, _030176_, _030177_, _030178_, _030179_, _030180_, _030181_, _030182_, _030183_, _030184_, _030185_, _030186_, _030187_, _030188_, _030189_, _030190_, _030191_, _030192_, _030193_, _030194_, _030195_, _030196_, _030197_, _030198_, _030199_, _030200_, _030201_, _030202_, _030203_, _030204_, _030205_, _030206_, _030207_, _030208_, _030209_, _030210_, _030211_, _030212_, _030213_, _030214_, _030215_, _030216_, _030217_, _030218_, _030219_, _030220_, _030221_, _030222_, _030223_, _030224_, _030225_, _030226_, _030227_, _030228_, _030229_, _030230_, _030231_, _030232_, _030233_, _030234_, _030235_, _030236_, _030237_, _030238_, _030239_, _030240_, _030241_, _030242_, _030243_, _030244_, _030245_, _030246_, _030247_, _030248_, _030249_, _030250_, _030251_, _030252_, _030253_, _030254_, _030255_, _030256_, _030257_, _030258_, _030259_, _030260_, _030261_, _030262_, _030263_, _030264_, _030265_, _030266_, _030267_, _030268_, _030269_, _030270_, _030271_, _030272_, _030273_, _030274_, _030275_, _030276_, _030277_, _030278_, _030279_, _030280_, _030281_, _030282_, _030283_, _030284_, _030285_, _030286_, _030287_, _030288_, _030289_, _030290_, _030291_, _030292_, _030293_, _030294_, _030295_, _030296_, _030297_, _030298_, _030299_, _030300_, _030301_, _030302_, _030303_, _030304_, _030305_, _030306_, _030307_, _030308_, _030309_, _030310_, _030311_, _030312_, _030313_, _030314_, _030315_, _030316_, _030317_, _030318_, _030319_, _030320_, _030321_, _030322_, _030323_, _030324_, _030325_, _030326_, _030327_, _030328_, _030329_, _030330_, _030331_, _030332_, _030333_, _030334_, _030335_, _030336_, _030337_, _030338_, _030339_, _030340_, _030341_, _030342_, _030343_, _030344_, _030345_, _030346_, _030347_, _030348_, _030349_, _030350_, _030351_, _030352_, _030353_, _030354_, _030355_, _030356_, _030357_, _030358_, _030359_, _030360_, _030361_, _030362_, _030363_, _030364_, _030365_, _030366_, _030367_, _030368_, _030369_, _030370_, _030371_, _030372_, _030373_, _030374_, _030375_, _030376_, _030377_, _030378_, _030379_, _030380_, _030381_, _030382_, _030383_, _030384_, _030385_, _030386_, _030387_, _030388_, _030389_, _030390_, _030391_, _030392_, _030393_, _030394_, _030395_, _030396_, _030397_, _030398_, _030399_, _030400_, _030401_, _030402_, _030403_, _030404_, _030405_, _030406_, _030407_, _030408_, _030409_, _030410_, _030411_, _030412_, _030413_, _030414_, _030415_, _030416_, _030417_, _030418_, _030419_, _030420_, _030421_, _030422_, _030423_, _030424_, _030425_, _030426_, _030427_, _030428_, _030429_, _030430_, _030431_, _030432_, _030433_, _030434_, _030435_, _030436_, _030437_, _030438_, _030439_, _030440_, _030441_, _030442_, _030443_, _030444_, _030445_, _030446_, _030447_, _030448_, _030449_, _030450_, _030451_, _030452_, _030453_, _030454_, _030455_, _030456_, _030457_, _030458_, _030459_, _030460_, _030461_, _030462_, _030463_, _030464_, _030465_, _030466_, _030467_, _030468_, _030469_, _030470_, _030471_, _030472_, _030473_, _030474_, _030475_, _030476_, _030477_, _030478_, _030479_, _030480_, _030481_, _030482_, _030483_, _030484_, _030485_, _030486_, _030487_, _030488_, _030489_, _030490_, _030491_, _030492_, _030493_, _030494_, _030495_, _030496_, _030497_, _030498_, _030499_, _030500_, _030501_, _030502_, _030503_, _030504_, _030505_, _030506_, _030507_, _030508_, _030509_, _030510_, _030511_, _030512_, _030513_, _030514_, _030515_, _030516_, _030517_, _030518_, _030519_, _030520_, _030521_, _030522_, _030523_, _030524_, _030525_, _030526_, _030527_, _030528_, _030529_, _030530_, _030531_, _030532_, _030533_, _030534_, _030535_, _030536_, _030537_, _030538_, _030539_, _030540_, _030541_, _030542_, _030543_, _030544_, _030545_, _030546_, _030547_, _030548_, _030549_, _030550_, _030551_, _030552_, _030553_, _030554_, _030555_, _030556_, _030557_, _030558_, _030559_, _030560_, _030561_, _030562_, _030563_, _030564_, _030565_, _030566_, _030567_, _030568_, _030569_, _030570_, _030571_, _030572_, _030573_, _030574_, _030575_, _030576_, _030577_, _030578_, _030579_, _030580_, _030581_, _030582_, _030583_, _030584_, _030585_, _030586_, _030587_, _030588_, _030589_, _030590_, _030591_, _030592_, _030593_, _030594_, _030595_, _030596_, _030597_, _030598_, _030599_, _030600_, _030601_, _030602_, _030603_, _030604_, _030605_, _030606_, _030607_, _030608_, _030609_, _030610_, _030611_, _030612_, _030613_, _030614_, _030615_, _030616_, _030617_, _030618_, _030619_, _030620_, _030621_, _030622_, _030623_, _030624_, _030625_, _030626_, _030627_, _030628_, _030629_, _030630_, _030631_, _030632_, _030633_, _030634_, _030635_, _030636_, _030637_, _030638_, _030639_, _030640_, _030641_, _030642_, _030643_, _030644_, _030645_, _030646_, _030647_, _030648_, _030649_, _030650_, _030651_, _030652_, _030653_, _030654_, _030655_, _030656_, _030657_, _030658_, _030659_, _030660_, _030661_, _030662_, _030663_, _030664_, _030665_, _030666_, _030667_, _030668_, _030669_, _030670_, _030671_, _030672_, _030673_, _030674_, _030675_, _030676_, _030677_, _030678_, _030679_, _030680_, _030681_, _030682_, _030683_, _030684_, _030685_, _030686_, _030687_, _030688_, _030689_, _030690_, _030691_, _030692_, _030693_, _030694_, _030695_, _030696_, _030697_, _030698_, _030699_, _030700_, _030701_, _030702_, _030703_, _030704_, _030705_, _030706_, _030707_, _030708_, _030709_, _030710_, _030711_, _030712_, _030713_, _030714_, _030715_, _030716_, _030717_, _030718_, _030719_, _030720_, _030721_, _030722_, _030723_, _030724_, _030725_, _030726_, _030727_, _030728_, _030729_, _030730_, _030731_, _030732_, _030733_, _030734_, _030735_, _030736_, _030737_, _030738_, _030739_, _030740_, _030741_, _030742_, _030743_, _030744_, _030745_, _030746_, _030747_, _030748_, _030749_, _030750_, _030751_, _030752_, _030753_, _030754_, _030755_, _030756_, _030757_, _030758_, _030759_, _030760_, _030761_, _030762_, _030763_, _030764_, _030765_, _030766_, _030767_, _030768_, _030769_, _030770_, _030771_, _030772_, _030773_, _030774_, _030775_, _030776_, _030777_, _030778_, _030779_, _030780_, _030781_, _030782_, _030783_, _030784_, _030785_, _030786_, _030787_, _030788_, _030789_, _030790_, _030791_, _030792_, _030793_, _030794_, _030795_, _030796_, _030797_, _030798_, _030799_, _030800_, _030801_, _030802_, _030803_, _030804_, _030805_, _030806_, _030807_, _030808_, _030809_, _030810_, _030811_, _030812_, _030813_, _030814_, _030815_, _030816_, _030817_, _030818_, _030819_, _030820_, _030821_, _030822_, _030823_, _030824_, _030825_, _030826_, _030827_, _030828_, _030829_, _030830_, _030831_, _030832_, _030833_, _030834_, _030835_, _030836_, _030837_, _030838_, _030839_, _030840_, _030841_, _030842_, _030843_, _030844_, _030845_, _030846_, _030847_, _030848_, _030849_, _030850_, _030851_, _030852_, _030853_, _030854_, _030855_, _030856_, _030857_, _030858_, _030859_, _030860_, _030861_, _030862_, _030863_, _030864_, _030865_, _030866_, _030867_, _030868_, _030869_, _030870_, _030871_, _030872_, _030873_, _030874_, _030875_, _030876_, _030877_, _030878_, _030879_, _030880_, _030881_, _030882_, _030883_, _030884_, _030885_, _030886_, _030887_, _030888_, _030889_, _030890_, _030891_, _030892_, _030893_, _030894_, _030895_, _030896_, _030897_, _030898_, _030899_, _030900_, _030901_, _030902_, _030903_, _030904_, _030905_, _030906_, _030907_, _030908_, _030909_, _030910_, _030911_, _030912_, _030913_, _030914_, _030915_, _030916_, _030917_, _030918_, _030919_, _030920_, _030921_, _030922_, _030923_, _030924_, _030925_, _030926_, _030927_, _030928_, _030929_, _030930_, _030931_, _030932_, _030933_, _030934_, _030935_, _030936_, _030937_, _030938_, _030939_, _030940_, _030941_, _030942_, _030943_, _030944_, _030945_, _030946_, _030947_, _030948_, _030949_, _030950_, _030951_, _030952_, _030953_, _030954_, _030955_, _030956_, _030957_, _030958_, _030959_, _030960_, _030961_, _030962_, _030963_, _030964_, _030965_, _030966_, _030967_, _030968_, _030969_, _030970_, _030971_, _030972_, _030973_, _030974_, _030975_, _030976_, _030977_, _030978_, _030979_, _030980_, _030981_, _030982_, _030983_, _030984_, _030985_, _030986_, _030987_, _030988_, _030989_, _030990_, _030991_, _030992_, _030993_, _030994_, _030995_, _030996_, _030997_, _030998_, _030999_, _031000_, _031001_, _031002_, _031003_, _031004_, _031005_, _031006_, _031007_, _031008_, _031009_, _031010_, _031011_, _031012_, _031013_, _031014_, _031015_, _031016_, _031017_, _031018_, _031019_, _031020_, _031021_, _031022_, _031023_, _031024_, _031025_, _031026_, _031027_, _031028_, _031029_, _031030_, _031031_, _031032_, _031033_, _031034_, _031035_, _031036_, _031037_, _031038_, _031039_, _031040_, _031041_, _031042_, _031043_, _031044_, _031045_, _031046_, _031047_, _031048_, _031049_, _031050_, _031051_, _031052_, _031053_, _031054_, _031055_, _031056_, _031057_, _031058_, _031059_, _031060_, _031061_, _031062_, _031063_, _031064_, _031065_, _031066_, _031067_, _031068_, _031069_, _031070_, _031071_, _031072_, _031073_, _031074_, _031075_, _031076_, _031077_, _031078_, _031079_, _031080_, _031081_, _031082_, _031083_, _031084_, _031085_, _031086_, _031087_, _031088_, _031089_, _031090_, _031091_, _031092_, _031093_, _031094_, _031095_, _031096_, _031097_, _031098_, _031099_, _031100_, _031101_, _031102_, _031103_, _031104_, _031105_, _031106_, _031107_, _031108_, _031109_, _031110_, _031111_, _031112_, _031113_, _031114_, _031115_, _031116_, _031117_, _031118_, _031119_, _031120_, _031121_, _031122_, _031123_, _031124_, _031125_, _031126_, _031127_, _031128_, _031129_, _031130_, _031131_, _031132_, _031133_, _031134_, _031135_, _031136_, _031137_, _031138_, _031139_, _031140_, _031141_, _031142_, _031143_, _031144_, _031145_, _031146_, _031147_, _031148_, _031149_, _031150_, _031151_, _031152_, _031153_, _031154_, _031155_, _031156_, _031157_, _031158_, _031159_, _031160_, _031161_, _031162_, _031163_, _031164_, _031165_, _031166_, _031167_, _031168_, _031169_, _031170_, _031171_, _031172_, _031173_, _031174_, _031175_, _031176_, _031177_, _031178_, _031179_, _031180_, _031181_, _031182_, _031183_, _031184_, _031185_, _031186_, _031187_, _031188_, _031189_, _031190_, _031191_, _031192_, _031193_, _031194_, _031195_, _031196_, _031197_, _031198_, _031199_, _031200_, _031201_, _031202_, _031203_, _031204_, _031205_, _031206_, _031207_, _031208_, _031209_, _031210_, _031211_, _031212_, _031213_, _031214_, _031215_, _031216_, _031217_, _031218_, _031219_, _031220_, _031221_, _031222_, _031223_, _031224_, _031225_, _031226_, _031227_, _031228_, _031229_, _031230_, _031231_, _031232_, _031233_, _031234_, _031235_, _031236_, _031237_, _031238_, _031239_, _031240_, _031241_, _031242_, _031243_, _031244_, _031245_, _031246_, _031247_, _031248_, _031249_, _031250_, _031251_, _031252_, _031253_, _031254_, _031255_, _031256_, _031257_, _031258_, _031259_, _031260_, _031261_, _031262_, _031263_, _031264_, _031265_, _031266_, _031267_, _031268_, _031269_, _031270_, _031271_, _031272_, _031273_, _031274_, _031275_, _031276_, _031277_, _031278_, _031279_, _031280_, _031281_, _031282_, _031283_, _031284_, _031285_, _031286_, _031287_, _031288_, _031289_, _031290_, _031291_, _031292_, _031293_, _031294_, _031295_, _031296_, _031297_, _031298_, _031299_, _031300_, _031301_, _031302_, _031303_, _031304_, _031305_, _031306_, _031307_, _031308_, _031309_, _031310_, _031311_, _031312_, _031313_, _031314_, _031315_, _031316_, _031317_, _031318_, _031319_, _031320_, _031321_, _031322_, _031323_, _031324_, _031325_, _031326_, _031327_, _031328_, _031329_, _031330_, _031331_, _031332_, _031333_, _031334_, _031335_, _031336_, _031337_, _031338_, _031339_, _031340_, _031341_, _031342_, _031343_, _031344_, _031345_, _031346_, _031347_, _031348_, _031349_, _031350_, _031351_, _031352_, _031353_, _031354_, _031355_, _031356_, _031357_, _031358_, _031359_, _031360_, _031361_, _031362_, _031363_, _031364_, _031365_, _031366_, _031367_, _031368_, _031369_, _031370_, _031371_, _031372_, _031373_, _031374_, _031375_, _031376_, _031377_, _031378_, _031379_, _031380_, _031381_, _031382_, _031383_, _031384_, _031385_, _031386_, _031387_, _031388_, _031389_, _031390_, _031391_, _031392_, _031393_, _031394_, _031395_, _031396_, _031397_, _031398_, _031399_, _031400_, _031401_, _031402_, _031403_, _031404_, _031405_, _031406_, _031407_, _031408_, _031409_, _031410_, _031411_, _031412_, _031413_, _031414_, _031415_, _031416_, _031417_, _031418_, _031419_, _031420_, _031421_, _031422_, _031423_, _031424_, _031425_, _031426_, _031427_, _031428_, _031429_, _031430_, _031431_, _031432_, _031433_, _031434_, _031435_, _031436_, _031437_, _031438_, _031439_, _031440_, _031441_, _031442_, _031443_, _031444_, _031445_, _031446_, _031447_, _031448_, _031449_, _031450_, _031451_, _031452_, _031453_, _031454_, _031455_, _031456_, _031457_, _031458_, _031459_, _031460_, _031461_, _031462_, _031463_, _031464_, _031465_, _031466_, _031467_, _031468_, _031469_, _031470_, _031471_, _031472_, _031473_, _031474_, _031475_, _031476_, _031477_, _031478_, _031479_, _031480_, _031481_, _031482_, _031483_, _031484_, _031485_, _031486_, _031487_, _031488_, _031489_, _031490_, _031491_, _031492_, _031493_, _031494_, _031495_, _031496_, _031497_, _031498_, _031499_, _031500_, _031501_, _031502_, _031503_, _031504_, _031505_, _031506_, _031507_, _031508_, _031509_, _031510_, _031511_, _031512_, _031513_, _031514_, _031515_, _031516_, _031517_, _031518_, _031519_, _031520_, _031521_, _031522_, _031523_, _031524_, _031525_, _031526_, _031527_, _031528_, _031529_, _031530_, _031531_, _031532_, _031533_, _031534_, _031535_, _031536_, _031537_, _031538_, _031539_, _031540_, _031541_, _031542_, _031543_, _031544_, _031545_, _031546_, _031547_, _031548_, _031549_, _031550_, _031551_, _031552_, _031553_, _031554_, _031555_, _031556_, _031557_, _031558_, _031559_, _031560_, _031561_, _031562_, _031563_, _031564_, _031565_, _031566_, _031567_, _031568_, _031569_, _031570_, _031571_, _031572_, _031573_, _031574_, _031575_, _031576_, _031577_, _031578_, _031579_, _031580_, _031581_, _031582_, _031583_, _031584_, _031585_, _031586_, _031587_, _031588_, _031589_, _031590_, _031591_, _031592_, _031593_, _031594_, _031595_, _031596_, _031597_, _031598_, _031599_, _031600_, _031601_, _031602_, _031603_, _031604_, _031605_, _031606_, _031607_, _031608_, _031609_, _031610_, _031611_, _031612_, _031613_, _031614_, _031615_, _031616_, _031617_, _031618_, _031619_, _031620_, _031621_, _031622_, _031623_, _031624_, _031625_, _031626_, _031627_, _031628_, _031629_, _031630_, _031631_, _031632_, _031633_, _031634_, _031635_, _031636_, _031637_, _031638_, _031639_, _031640_, _031641_, _031642_, _031643_, _031644_, _031645_, _031646_, _031647_, _031648_, _031649_, _031650_, _031651_, _031652_, _031653_, _031654_, _031655_, _031656_, _031657_, _031658_, _031659_, _031660_, _031661_, _031662_, _031663_, _031664_, _031665_, _031666_, _031667_, _031668_, _031669_, _031670_, _031671_, _031672_, _031673_, _031674_, _031675_, _031676_, _031677_, _031678_, _031679_, _031680_, _031681_, _031682_, _031683_, _031684_, _031685_, _031686_, _031687_, _031688_, _031689_, _031690_, _031691_, _031692_, _031693_, _031694_, _031695_, _031696_, _031697_, _031698_, _031699_, _031700_, _031701_, _031702_, _031703_, _031704_, _031705_, _031706_, _031707_, _031708_, _031709_, _031710_, _031711_, _031712_, _031713_, _031714_, _031715_, _031716_, _031717_, _031718_, _031719_, _031720_, _031721_, _031722_, _031723_, _031724_, _031725_, _031726_, _031727_, _031728_, _031729_, _031730_, _031731_, _031732_, _031733_, _031734_, _031735_, _031736_, _031737_, _031738_, _031739_, _031740_, _031741_, _031742_, _031743_, _031744_, _031745_, _031746_, _031747_, _031748_, _031749_, _031750_, _031751_, _031752_, _031753_, _031754_, _031755_, _031756_, _031757_, _031758_, _031759_, _031760_, _031761_, _031762_, _031763_, _031764_, _031765_, _031766_, _031767_, _031768_, _031769_, _031770_, _031771_, _031772_, _031773_, _031774_, _031775_, _031776_, _031777_, _031778_, _031779_, _031780_, _031781_, _031782_, _031783_, _031784_, _031785_, _031786_, _031787_, _031788_, _031789_, _031790_, _031791_, _031792_, _031793_, _031794_, _031795_, _031796_, _031797_, _031798_, _031799_, _031800_, _031801_, _031802_, _031803_, _031804_, _031805_, _031806_, _031807_, _031808_, _031809_, _031810_, _031811_, _031812_, _031813_, _031814_, _031815_, _031816_, _031817_, _031818_, _031819_, _031820_, _031821_, _031822_, _031823_, _031824_, _031825_, _031826_, _031827_, _031828_, _031829_, _031830_, _031831_, _031832_, _031833_, _031834_, _031835_, _031836_, _031837_, _031838_, _031839_, _031840_, _031841_, _031842_, _031843_, _031844_, _031845_, _031846_, _031847_, _031848_, _031849_, _031850_, _031851_, _031852_, _031853_, _031854_, _031855_, _031856_, _031857_, _031858_, _031859_, _031860_, _031861_, _031862_, _031863_, _031864_, _031865_, _031866_, _031867_, _031868_, _031869_, _031870_, _031871_, _031872_, _031873_, _031874_, _031875_, _031876_, _031877_, _031878_, _031879_, _031880_, _031881_, _031882_, _031883_, _031884_, _031885_, _031886_, _031887_, _031888_, _031889_, _031890_, _031891_, _031892_, _031893_, _031894_, _031895_, _031896_, _031897_, _031898_, _031899_, _031900_, _031901_, _031902_, _031903_, _031904_, _031905_, _031906_, _031907_, _031908_, _031909_, _031910_, _031911_, _031912_, _031913_, _031914_, _031915_, _031916_, _031917_, _031918_, _031919_, _031920_, _031921_, _031922_, _031923_, _031924_, _031925_, _031926_, _031927_, _031928_, _031929_, _031930_, _031931_, _031932_, _031933_, _031934_, _031935_, _031936_, _031937_, _031938_, _031939_, _031940_, _031941_, _031942_, _031943_, _031944_, _031945_, _031946_, _031947_, _031948_, _031949_, _031950_, _031951_, _031952_, _031953_, _031954_, _031955_, _031956_, _031957_, _031958_, _031959_, _031960_, _031961_, _031962_, _031963_, _031964_, _031965_, _031966_, _031967_, _031968_, _031969_, _031970_, _031971_, _031972_, _031973_, _031974_, _031975_, _031976_, _031977_, _031978_, _031979_, _031980_, _031981_, _031982_, _031983_, _031984_, _031985_, _031986_, _031987_, _031988_, _031989_, _031990_, _031991_, _031992_, _031993_, _031994_, _031995_, _031996_, _031997_, _031998_, _031999_, _032000_, _032001_, _032002_, _032003_, _032004_, _032005_, _032006_, _032007_, _032008_, _032009_, _032010_, _032011_, _032012_, _032013_, _032014_, _032015_, _032016_, _032017_, _032018_, _032019_, _032020_, _032021_, _032022_, _032023_, _032024_, _032025_, _032026_, _032027_, _032028_, _032029_, _032030_, _032031_, _032032_, _032033_, _032034_, _032035_, _032036_, _032037_, _032038_, _032039_, _032040_, _032041_, _032042_, _032043_, _032044_, _032045_, _032046_, _032047_, _032048_, _032049_, _032050_, _032051_, _032052_, _032053_, _032054_, _032055_, _032056_, _032057_, _032058_, _032059_, _032060_, _032061_, _032062_, _032063_, _032064_, _032065_, _032066_, _032067_, _032068_, _032069_, _032070_, _032071_, _032072_, _032073_, _032074_, _032075_, _032076_, _032077_, _032078_, _032079_, _032080_, _032081_, _032082_, _032083_, _032084_, _032085_, _032086_, _032087_, _032088_, _032089_, _032090_, _032091_, _032092_, _032093_, _032094_, _032095_, _032096_, _032097_, _032098_, _032099_, _032100_, _032101_, _032102_, _032103_, _032104_, _032105_, _032106_, _032107_, _032108_, _032109_, _032110_, _032111_, _032112_, _032113_, _032114_, _032115_, _032116_, _032117_, _032118_, _032119_, _032120_, _032121_, _032122_, _032123_, _032124_, _032125_, _032126_, _032127_, _032128_, _032129_, _032130_, _032131_, _032132_, _032133_, _032134_, _032135_, _032136_, _032137_, _032138_, _032139_, _032140_, _032141_, _032142_, _032143_, _032144_, _032145_, _032146_, _032147_, _032148_, _032149_, _032150_, _032151_, _032152_, _032153_, _032154_, _032155_, _032156_, _032157_, _032158_, _032159_, _032160_, _032161_, _032162_, _032163_, _032164_, _032165_, _032166_, _032167_, _032168_, _032169_, _032170_, _032171_, _032172_, _032173_, _032174_, _032175_, _032176_, _032177_, _032178_, _032179_, _032180_, _032181_, _032182_, _032183_, _032184_, _032185_, _032186_, _032187_, _032188_, _032189_, _032190_, _032191_, _032192_, _032193_, _032194_, _032195_, _032196_, _032197_, _032198_, _032199_, _032200_, _032201_, _032202_, _032203_, _032204_, _032205_, _032206_, _032207_, _032208_, _032209_, _032210_, _032211_, _032212_, _032213_, _032214_, _032215_, _032216_, _032217_, _032218_, _032219_, _032220_, _032221_, _032222_, _032223_, _032224_, _032225_, _032226_, _032227_, _032228_, _032229_, _032230_, _032231_, _032232_, _032233_, _032234_, _032235_, _032236_, _032237_, _032238_, _032239_, _032240_, _032241_, _032242_, _032243_, _032244_, _032245_, _032246_, _032247_, _032248_, _032249_, _032250_, _032251_, _032252_, _032253_, _032254_, _032255_, _032256_, _032257_, _032258_, _032259_, _032260_, _032261_, _032262_, _032263_, _032264_, _032265_, _032266_, _032267_, _032268_, _032269_, _032270_, _032271_, _032272_, _032273_, _032274_, _032275_, _032276_, _032277_, _032278_, _032279_, _032280_, _032281_, _032282_, _032283_, _032284_, _032285_, _032286_, _032287_, _032288_, _032289_, _032290_, _032291_, _032292_, _032293_, _032294_, _032295_, _032296_, _032297_, _032298_, _032299_, _032300_, _032301_, _032302_, _032303_, _032304_, _032305_, _032306_, _032307_, _032308_, _032309_, _032310_, _032311_, _032312_, _032313_, _032314_, _032315_, _032316_, _032317_, _032318_, _032319_, _032320_, _032321_, _032322_, _032323_, _032324_, _032325_, _032326_, _032327_, _032328_, _032329_, _032330_, _032331_, _032332_, _032333_, _032334_, _032335_, _032336_, _032337_, _032338_, _032339_, _032340_, _032341_, _032342_, _032343_, _032344_, _032345_, _032346_, _032347_, _032348_, _032349_, _032350_, _032351_, _032352_, _032353_, _032354_, _032355_, _032356_, _032357_, _032358_, _032359_, _032360_, _032361_, _032362_, _032363_, _032364_, _032365_, _032366_, _032367_, _032368_, _032369_, _032370_, _032371_, _032372_, _032373_, _032374_, _032375_, _032376_, _032377_, _032378_, _032379_, _032380_, _032381_, _032382_, _032383_, _032384_, _032385_, _032386_, _032387_, _032388_, _032389_, _032390_, _032391_, _032392_, _032393_, _032394_, _032395_, _032396_, _032397_, _032398_, _032399_, _032400_, _032401_, _032402_, _032403_, _032404_, _032405_, _032406_, _032407_, _032408_, _032409_, _032410_, _032411_, _032412_, _032413_, _032414_, _032415_, _032416_, _032417_, _032418_, _032419_, _032420_, _032421_, _032422_, _032423_, _032424_, _032425_, _032426_, _032427_, _032428_, _032429_, _032430_, _032431_, _032432_, _032433_, _032434_, _032435_, _032436_, _032437_, _032438_, _032439_, _032440_, _032441_, _032442_, _032443_, _032444_, _032445_, _032446_, _032447_, _032448_, _032449_, _032450_, _032451_, _032452_, _032453_, _032454_, _032455_, _032456_, _032457_, _032458_, _032459_, _032460_, _032461_, _032462_, _032463_, _032464_, _032465_, _032466_, _032467_, _032468_, _032469_, _032470_, _032471_, _032472_, _032473_, _032474_, _032475_, _032476_, _032477_, _032478_, _032479_, _032480_, _032481_, _032482_, _032483_, _032484_, _032485_, _032486_, _032487_, _032488_, _032489_, _032490_, _032491_, _032492_, _032493_, _032494_, _032495_, _032496_, _032497_, _032498_, _032499_, _032500_, _032501_, _032502_, _032503_, _032504_, _032505_, _032506_, _032507_, _032508_, _032509_, _032510_, _032511_, _032512_, _032513_, _032514_, _032515_, _032516_, _032517_, _032518_, _032519_, _032520_, _032521_, _032522_, _032523_, _032524_, _032525_, _032526_, _032527_, _032528_, _032529_, _032530_, _032531_, _032532_, _032533_, _032534_, _032535_, _032536_, _032537_, _032538_, _032539_, _032540_, _032541_, _032542_, _032543_, _032544_, _032545_, _032546_, _032547_, _032548_, _032549_, _032550_, _032551_, _032552_, _032553_, _032554_, _032555_, _032556_, _032557_, _032558_, _032559_, _032560_, _032561_, _032562_, _032563_, _032564_, _032565_, _032566_, _032567_, _032568_, _032569_, _032570_, _032571_, _032572_, _032573_, _032574_, _032575_, _032576_, _032577_, _032578_, _032579_, _032580_, _032581_, _032582_, _032583_, _032584_, _032585_, _032586_, _032587_, _032588_, _032589_, _032590_, _032591_, _032592_, _032593_, _032594_, _032595_, _032596_, _032597_, _032598_, _032599_, _032600_, _032601_, _032602_, _032603_, _032604_, _032605_, _032606_, _032607_, _032608_, _032609_, _032610_, _032611_, _032612_, _032613_, _032614_, _032615_, _032616_, _032617_, _032618_, _032619_, _032620_, _032621_, _032622_, _032623_, _032624_, _032625_, _032626_, _032627_, _032628_, _032629_, _032630_, _032631_, _032632_, _032633_, _032634_, _032635_, _032636_, _032637_, _032638_, _032639_, _032640_, _032641_, _032642_, _032643_, _032644_, _032645_, _032646_, _032647_, _032648_, _032649_, _032650_, _032651_, _032652_, _032653_, _032654_, _032655_, _032656_, _032657_, _032658_, _032659_, _032660_, _032661_, _032662_, _032663_, _032664_, _032665_, _032666_, _032667_, _032668_, _032669_, _032670_, _032671_, _032672_, _032673_, _032674_, _032675_, _032676_, _032677_, _032678_, _032679_, _032680_, _032681_, _032682_, _032683_, _032684_, _032685_, _032686_, _032687_, _032688_, _032689_, _032690_, _032691_, _032692_, _032693_, _032694_, _032695_, _032696_, _032697_, _032698_, _032699_, _032700_, _032701_, _032702_, _032703_, _032704_, _032705_, _032706_, _032707_, _032708_, _032709_, _032710_, _032711_, _032712_, _032713_, _032714_, _032715_, _032716_, _032717_, _032718_, _032719_, _032720_, _032721_, _032722_, _032723_, _032724_, _032725_, _032726_, _032727_, _032728_, _032729_, _032730_, _032731_, _032732_, _032733_, _032734_, _032735_, _032736_, _032737_, _032738_, _032739_, _032740_, _032741_, _032742_, _032743_, _032744_, _032745_, _032746_, _032747_, _032748_, _032749_, _032750_, _032751_, _032752_, _032753_, _032754_, _032755_, _032756_, _032757_, _032758_, _032759_, _032760_, _032761_, _032762_, _032763_, _032764_, _032765_, _032766_, _032767_, _032768_, _032769_, _032770_, _032771_, _032772_, _032773_, _032774_, _032775_, _032776_, _032777_, _032778_, _032779_, _032780_, _032781_, _032782_, _032783_, _032784_, _032785_, _032786_, _032787_, _032788_, _032789_, _032790_, _032791_, _032792_, _032793_, _032794_, _032795_, _032796_, _032797_, _032798_, _032799_, _032800_, _032801_, _032802_, _032803_, _032804_, _032805_, _032806_, _032807_, _032808_, _032809_, _032810_, _032811_, _032812_, _032813_, _032814_, _032815_, _032816_, _032817_, _032818_, _032819_, _032820_, _032821_, _032822_, _032823_, _032824_, _032825_, _032826_, _032827_, _032828_, _032829_, _032830_, _032831_, _032832_, _032833_, _032834_, _032835_, _032836_, _032837_, _032838_, _032839_, _032840_, _032841_, _032842_, _032843_, _032844_, _032845_, _032846_, _032847_, _032848_, _032849_, _032850_, _032851_, _032852_, _032853_, _032854_, _032855_, _032856_, _032857_, _032858_, _032859_, _032860_, _032861_, _032862_, _032863_, _032864_, _032865_, _032866_, _032867_, _032868_, _032869_, _032870_, _032871_, _032872_, _032873_, _032874_, _032875_, _032876_, _032877_, _032878_, _032879_, _032880_, _032881_, _032882_, _032883_, _032884_, _032885_, _032886_, _032887_, _032888_, _032889_, _032890_, _032891_, _032892_, _032893_, _032894_, _032895_, _032896_, _032897_, _032898_, _032899_, _032900_, _032901_, _032902_, _032903_, _032904_, _032905_, _032906_, _032907_, _032908_, _032909_, _032910_, _032911_, _032912_, _032913_, _032914_, _032915_, _032916_, _032917_, _032918_, _032919_, _032920_, _032921_, _032922_, _032923_, _032924_, _032925_, _032926_, _032927_, _032928_, _032929_, _032930_, _032931_, _032932_, _032933_, _032934_, _032935_, _032936_, _032937_, _032938_, _032939_, _032940_, _032941_, _032942_, _032943_, _032944_, _032945_, _032946_, _032947_, _032948_, _032949_, _032950_, _032951_, _032952_, _032953_, _032954_, _032955_, _032956_, _032957_, _032958_, _032959_, _032960_, _032961_, _032962_, _032963_, _032964_, _032965_, _032966_, _032967_, _032968_, _032969_, _032970_, _032971_, _032972_, _032973_, _032974_, _032975_, _032976_, _032977_, _032978_, _032979_, _032980_, _032981_, _032982_, _032983_, _032984_, _032985_, _032986_, _032987_, _032988_, _032989_, _032990_, _032991_, _032992_, _032993_, _032994_, _032995_, _032996_, _032997_, _032998_, _032999_, _033000_, _033001_, _033002_, _033003_, _033004_, _033005_, _033006_, _033007_, _033008_, _033009_, _033010_, _033011_, _033012_, _033013_, _033014_, _033015_, _033016_, _033017_, _033018_, _033019_, _033020_, _033021_, _033022_, _033023_, _033024_, _033025_, _033026_, _033027_, _033028_, _033029_, _033030_, _033031_, _033032_, _033033_, _033034_, _033035_, _033036_, _033037_, _033038_, _033039_, _033040_, _033041_, _033042_, _033043_, _033044_, _033045_, _033046_, _033047_, _033048_, _033049_, _033050_, _033051_, _033052_, _033053_, _033054_, _033055_, _033056_, _033057_, _033058_, _033059_, _033060_, _033061_, _033062_, _033063_, _033064_, _033065_, _033066_, _033067_, _033068_, _033069_, _033070_, _033071_, _033072_, _033073_, _033074_, _033075_, _033076_, _033077_, _033078_, _033079_, _033080_, _033081_, _033082_, _033083_, _033084_, _033085_, _033086_, _033087_, _033088_, _033089_, _033090_, _033091_, _033092_, _033093_, _033094_, _033095_, _033096_, _033097_, _033098_, _033099_, _033100_, _033101_, _033102_, _033103_, _033104_, _033105_, _033106_, _033107_, _033108_, _033109_, _033110_, _033111_, _033112_, _033113_, _033114_, _033115_, _033116_, _033117_, _033118_, _033119_, _033120_, _033121_, _033122_, _033123_, _033124_, _033125_, _033126_, _033127_, _033128_, _033129_, _033130_, _033131_, _033132_, _033133_, _033134_, _033135_, _033136_, _033137_, _033138_, _033139_, _033140_, _033141_, _033142_, _033143_, _033144_, _033145_, _033146_, _033147_, _033148_, _033149_, _033150_, _033151_, _033152_, _033153_, _033154_, _033155_, _033156_, _033157_, _033158_, _033159_, _033160_, _033161_, _033162_, _033163_, _033164_, _033165_, _033166_, _033167_, _033168_, _033169_, _033170_, _033171_, _033172_, _033173_, _033174_, _033175_, _033176_, _033177_, _033178_, _033179_, _033180_, _033181_, _033182_, _033183_, _033184_, _033185_, _033186_, _033187_, _033188_, _033189_, _033190_, _033191_, _033192_, _033193_, _033194_, _033195_, _033196_, _033197_, _033198_, _033199_, _033200_, _033201_, _033202_, _033203_, _033204_, _033205_, _033206_, _033207_, _033208_, _033209_, _033210_, _033211_, _033212_, _033213_, _033214_, _033215_, _033216_, _033217_, _033218_, _033219_, _033220_, _033221_, _033222_, _033223_, _033224_, _033225_, _033226_, _033227_, _033228_, _033229_, _033230_, _033231_, _033232_, _033233_, _033234_, _033235_, _033236_, _033237_, _033238_, _033239_, _033240_, _033241_, _033242_, _033243_, _033244_, _033245_, _033246_, _033247_, _033248_, _033249_, _033250_, _033251_, _033252_, _033253_, _033254_, _033255_, _033256_, _033257_, _033258_, _033259_, _033260_, _033261_, _033262_, _033263_, _033264_, _033265_, _033266_, _033267_, _033268_, _033269_, _033270_, _033271_, _033272_, _033273_, _033274_, _033275_, _033276_, _033277_, _033278_, _033279_, _033280_, _033281_, _033282_, _033283_, _033284_, _033285_, _033286_, _033287_, _033288_, _033289_, _033290_, _033291_, _033292_, _033293_, _033294_, _033295_, _033296_, _033297_, _033298_, _033299_, _033300_, _033301_, _033302_, _033303_, _033304_, _033305_, _033306_, _033307_, _033308_, _033309_, _033310_, _033311_, _033312_, _033313_, _033314_, _033315_, _033316_, _033317_, _033318_, _033319_, _033320_, _033321_, _033322_, _033323_, _033324_, _033325_, _033326_, _033327_, _033328_, _033329_, _033330_, _033331_, _033332_, _033333_, _033334_, _033335_, _033336_, _033337_, _033338_, _033339_, _033340_, _033341_, _033342_, _033343_, _033344_, _033345_, _033346_, _033347_, _033348_, _033349_, _033350_, _033351_, _033352_, _033353_, _033354_, _033355_, _033356_, _033357_, _033358_, _033359_, _033360_, _033361_, _033362_, _033363_, _033364_, _033365_, _033366_, _033367_, _033368_, _033369_, _033370_, _033371_, _033372_, _033373_, _033374_, _033375_, _033376_, _033377_, _033378_, _033379_, _033380_, _033381_, _033382_, _033383_, _033384_, _033385_, _033386_, _033387_, _033388_, _033389_, _033390_, _033391_, _033392_, _033393_, _033394_, _033395_, _033396_, _033397_, _033398_, _033399_, _033400_, _033401_, _033402_, _033403_, _033404_, _033405_, _033406_, _033407_, _033408_, _033409_, _033410_, _033411_, _033412_, _033413_, _033414_, _033415_, _033416_, _033417_, _033418_, _033419_, _033420_, _033421_, _033422_, _033423_, _033424_, _033425_, _033426_, _033427_, _033428_, _033429_, _033430_, _033431_, _033432_, _033433_, _033434_, _033435_, _033436_, _033437_, _033438_, _033439_, _033440_, _033441_, _033442_, _033443_, _033444_, _033445_, _033446_, _033447_, _033448_, _033449_, _033450_, _033451_, _033452_, _033453_, _033454_, _033455_, _033456_, _033457_, _033458_, _033459_, _033460_, _033461_, _033462_, _033463_, _033464_, _033465_, _033466_, _033467_, _033468_, _033469_, _033470_, _033471_, _033472_, _033473_, _033474_, _033475_, _033476_, _033477_, _033478_, _033479_, _033480_, _033481_, _033482_, _033483_, _033484_, _033485_, _033486_, _033487_, _033488_, _033489_, _033490_, _033491_, _033492_, _033493_, _033494_, _033495_, _033496_, _033497_, _033498_, _033499_, _033500_, _033501_, _033502_, _033503_, _033504_, _033505_, _033506_, _033507_, _033508_, _033509_, _033510_, _033511_, _033512_, _033513_, _033514_, _033515_, _033516_, _033517_, _033518_, _033519_, _033520_, _033521_, _033522_, _033523_, _033524_, _033525_, _033526_, _033527_, _033528_, _033529_, _033530_, _033531_, _033532_, _033533_, _033534_, _033535_, _033536_, _033537_, _033538_, _033539_, _033540_, _033541_, _033542_, _033543_, _033544_, _033545_, _033546_, _033547_, _033548_, _033549_, _033550_, _033551_, _033552_, _033553_, _033554_, _033555_, _033556_, _033557_, _033558_, _033559_, _033560_, _033561_, _033562_, _033563_, _033564_, _033565_, _033566_, _033567_, _033568_, _033569_, _033570_, _033571_, _033572_, _033573_, _033574_, _033575_, _033576_, _033577_, _033578_, _033579_, _033580_, _033581_, _033582_, _033583_, _033584_, _033585_, _033586_, _033587_, _033588_, _033589_, _033590_, _033591_, _033592_, _033593_, _033594_, _033595_, _033596_, _033597_, _033598_, _033599_, _033600_, _033601_, _033602_, _033603_, _033604_, _033605_, _033606_, _033607_, _033608_, _033609_, _033610_, _033611_, _033612_, _033613_, _033614_, _033615_, _033616_, _033617_, _033618_, _033619_, _033620_, _033621_, _033622_, _033623_, _033624_, _033625_, _033626_, _033627_, _033628_, _033629_, _033630_, _033631_, _033632_, _033633_, _033634_, _033635_, _033636_, _033637_, _033638_, _033639_, _033640_, _033641_, _033642_, _033643_, _033644_, _033645_, _033646_, _033647_, _033648_, _033649_, _033650_, _033651_, _033652_, _033653_, _033654_, _033655_, _033656_, _033657_, _033658_, _033659_, _033660_, _033661_, _033662_, _033663_, _033664_, _033665_, _033666_, _033667_, _033668_, _033669_, _033670_, _033671_, _033672_, _033673_, _033674_, _033675_, _033676_, _033677_, _033678_, _033679_, _033680_, _033681_, _033682_, _033683_, _033684_, _033685_, _033686_, _033687_, _033688_, _033689_, _033690_, _033691_, _033692_, _033693_, _033694_, _033695_, _033696_, _033697_, _033698_, _033699_, _033700_, _033701_, _033702_, _033703_, _033704_, _033705_, _033706_, _033707_, _033708_, _033709_, _033710_, _033711_, _033712_, _033713_, _033714_, _033715_, _033716_, _033717_, _033718_, _033719_, _033720_, _033721_, _033722_, _033723_, _033724_, _033725_, _033726_, _033727_, _033728_, _033729_, _033730_, _033731_, _033732_, _033733_, _033734_, _033735_, _033736_, _033737_, _033738_, _033739_, _033740_, _033741_, _033742_, _033743_, _033744_, _033745_, _033746_, _033747_, _033748_, _033749_, _033750_, _033751_, _033752_, _033753_, _033754_, _033755_, _033756_, _033757_, _033758_, _033759_, _033760_, _033761_, _033762_, _033763_, _033764_, _033765_, _033766_, _033767_, _033768_, _033769_, _033770_, _033771_, _033772_, _033773_, _033774_, _033775_, _033776_, _033777_, _033778_, _033779_, _033780_, _033781_, _033782_, _033783_, _033784_, _033785_, _033786_, _033787_, _033788_, _033789_, _033790_, _033791_, _033792_, _033793_, _033794_, _033795_, _033796_, _033797_, _033798_, _033799_, _033800_, _033801_, _033802_, _033803_, _033804_, _033805_, _033806_, _033807_, _033808_, _033809_, _033810_, _033811_, _033812_, _033813_, _033814_, _033815_, _033816_, _033817_, _033818_, _033819_, _033820_, _033821_, _033822_, _033823_, _033824_, _033825_, _033826_, _033827_, _033828_, _033829_, _033830_, _033831_, _033832_, _033833_, _033834_, _033835_, _033836_, _033837_, _033838_, _033839_, _033840_, _033841_, _033842_, _033843_, _033844_, _033845_, _033846_, _033847_, _033848_, _033849_, _033850_, _033851_, _033852_, _033853_, _033854_, _033855_, _033856_, _033857_, _033858_, _033859_, _033860_, _033861_, _033862_, _033863_, _033864_, _033865_, _033866_, _033867_, _033868_, _033869_, _033870_, _033871_, _033872_, _033873_, _033874_, _033875_, _033876_, _033877_, _033878_, _033879_, _033880_, _033881_, _033882_, _033883_, _033884_, _033885_, _033886_, _033887_, _033888_, _033889_, _033890_, _033891_, _033892_, _033893_, _033894_, _033895_, _033896_, _033897_, _033898_, _033899_, _033900_, _033901_, _033902_, _033903_, _033904_, _033905_, _033906_, _033907_, _033908_, _033909_, _033910_, _033911_, _033912_, _033913_, _033914_, _033915_, _033916_, _033917_, _033918_, _033919_, _033920_, _033921_, _033922_, _033923_, _033924_, _033925_, _033926_, _033927_, _033928_, _033929_, _033930_, _033931_, _033932_, _033933_, _033934_, _033935_, _033936_, _033937_, _033938_, _033939_, _033940_, _033941_, _033942_, _033943_, _033944_, _033945_, _033946_, _033947_, _033948_, _033949_, _033950_, _033951_, _033952_, _033953_, _033954_, _033955_, _033956_, _033957_, _033958_, _033959_, _033960_, _033961_, _033962_, _033963_, _033964_, _033965_, _033966_, _033967_, _033968_, _033969_, _033970_, _033971_, _033972_, _033973_, _033974_, _033975_, _033976_, _033977_, _033978_, _033979_, _033980_, _033981_, _033982_, _033983_, _033984_, _033985_, _033986_, _033987_, _033988_, _033989_, _033990_, _033991_, _033992_, _033993_, _033994_, _033995_, _033996_, _033997_, _033998_, _033999_, _034000_, _034001_, _034002_, _034003_, _034004_, _034005_, _034006_, _034007_, _034008_, _034009_, _034010_, _034011_, _034012_, _034013_, _034014_, _034015_, _034016_, _034017_, _034018_, _034019_, _034020_, _034021_, _034022_, _034023_, _034024_, _034025_, _034026_, _034027_, _034028_, _034029_, _034030_, _034031_, _034032_, _034033_, _034034_, _034035_, _034036_, _034037_, _034038_, _034039_, _034040_, _034041_, _034042_, _034043_, _034044_, _034045_, _034046_, _034047_, _034048_, _034049_, _034050_, _034051_, _034052_, _034053_, _034054_, _034055_, _034056_, _034057_, _034058_, _034059_, _034060_, _034061_, _034062_, _034063_, _034064_, _034065_, _034066_, _034067_, _034068_, _034069_, _034070_, _034071_, _034072_, _034073_, _034074_, _034075_, _034076_, _034077_, _034078_, _034079_, _034080_, _034081_, _034082_, _034083_, _034084_, _034085_, _034086_, _034087_, _034088_, _034089_, _034090_, _034091_, _034092_, _034093_, _034094_, _034095_, _034096_, _034097_, _034098_, _034099_, _034100_, _034101_, _034102_, _034103_, _034104_, _034105_, _034106_, _034107_, _034108_, _034109_, _034110_, _034111_, _034112_, _034113_, _034114_, _034115_, _034116_, _034117_, _034118_, _034119_, _034120_, _034121_, _034122_, _034123_, _034124_, _034125_, _034126_, _034127_, _034128_, _034129_, _034130_, _034131_, _034132_, _034133_, _034134_, _034135_, _034136_, _034137_, _034138_, _034139_, _034140_, _034141_, _034142_, _034143_, _034144_, _034145_, _034146_, _034147_, _034148_, _034149_, _034150_, _034151_, _034152_, _034153_, _034154_, _034155_, _034156_, _034157_, _034158_, _034159_, _034160_, _034161_, _034162_, _034163_, _034164_, _034165_, _034166_, _034167_, _034168_, _034169_, _034170_, _034171_, _034172_, _034173_, _034174_, _034175_, _034176_, _034177_, _034178_, _034179_, _034180_, _034181_, _034182_, _034183_, _034184_, _034185_, _034186_, _034187_, _034188_, _034189_, _034190_, _034191_, _034192_, _034193_, _034194_, _034195_, _034196_, _034197_, _034198_, _034199_, _034200_, _034201_, _034202_, _034203_, _034204_, _034205_, _034206_, _034207_, _034208_, _034209_, _034210_, _034211_, _034212_, _034213_, _034214_, _034215_, _034216_, _034217_, _034218_, _034219_, _034220_, _034221_, _034222_, _034223_, _034224_, _034225_, _034226_, _034227_, _034228_, _034229_, _034230_, _034231_, _034232_, _034233_, _034234_, _034235_, _034236_, _034237_, _034238_, _034239_, _034240_, _034241_, _034242_, _034243_, _034244_, _034245_, _034246_, _034247_, _034248_, _034249_, _034250_, _034251_, _034252_, _034253_, _034254_, _034255_, _034256_, _034257_, _034258_, _034259_, _034260_, _034261_, _034262_, _034263_, _034264_, _034265_, _034266_, _034267_, _034268_, _034269_, _034270_, _034271_, _034272_, _034273_, _034274_, _034275_, _034276_, _034277_, _034278_, _034279_, _034280_, _034281_, _034282_, _034283_, _034284_, _034285_, _034286_, _034287_, _034288_, _034289_, _034290_, _034291_, _034292_, _034293_, _034294_, _034295_, _034296_, _034297_, _034298_, _034299_, _034300_, _034301_, _034302_, _034303_, _034304_, _034305_, _034306_, _034307_, _034308_, _034309_, _034310_, _034311_, _034312_, _034313_, _034314_, _034315_, _034316_, _034317_, _034318_, _034319_, _034320_, _034321_, _034322_, _034323_, _034324_, _034325_, _034326_, _034327_, _034328_, _034329_, _034330_, _034331_, _034332_, _034333_, _034334_, _034335_, _034336_, _034337_, _034338_, _034339_, _034340_, _034341_, _034342_, _034343_, _034344_, _034345_, _034346_, _034347_, _034348_, _034349_, _034350_, _034351_, _034352_, _034353_, _034354_, _034355_, _034356_, _034357_, _034358_, _034359_, _034360_, _034361_, _034362_, _034363_, _034364_, _034365_, _034366_, _034367_, _034368_, _034369_, _034370_, _034371_, _034372_, _034373_, _034374_, _034375_, _034376_, _034377_, _034378_, _034379_, _034380_, _034381_, _034382_, _034383_, _034384_, _034385_, _034386_, _034387_, _034388_, _034389_, _034390_, _034391_, _034392_, _034393_, _034394_, _034395_, _034396_, _034397_, _034398_, _034399_, _034400_, _034401_, _034402_, _034403_, _034404_, _034405_, _034406_, _034407_, _034408_, _034409_, _034410_, _034411_, _034412_, _034413_, _034414_, _034415_, _034416_, _034417_, _034418_, _034419_, _034420_, _034421_, _034422_, _034423_, _034424_, _034425_, _034426_, _034427_, _034428_, _034429_, _034430_, _034431_, _034432_, _034433_, _034434_, _034435_, _034436_, _034437_, _034438_, _034439_, _034440_, _034441_, _034442_, _034443_, _034444_, _034445_, _034446_, _034447_, _034448_, _034449_, _034450_, _034451_, _034452_, _034453_, _034454_, _034455_, _034456_, _034457_, _034458_, _034459_, _034460_, _034461_, _034462_, _034463_, _034464_, _034465_, _034466_, _034467_, _034468_, _034469_, _034470_, _034471_, _034472_, _034473_, _034474_, _034475_, _034476_, _034477_, _034478_, _034479_, _034480_, _034481_, _034482_, _034483_, _034484_, _034485_, _034486_, _034487_, _034488_, _034489_, _034490_, _034491_, _034492_, _034493_, _034494_, _034495_, _034496_, _034497_, _034498_, _034499_, _034500_, _034501_, _034502_, _034503_, _034504_, _034505_, _034506_, _034507_, _034508_, _034509_, _034510_, _034511_, _034512_, _034513_, _034514_, _034515_, _034516_, _034517_, _034518_, _034519_, _034520_, _034521_, _034522_, _034523_, _034524_, _034525_, _034526_, _034527_, _034528_, _034529_, _034530_, _034531_, _034532_, _034533_, _034534_, _034535_, _034536_, _034537_, _034538_, _034539_, _034540_, _034541_, _034542_, _034543_, _034544_, _034545_, _034546_, _034547_, _034548_, _034549_, _034550_, _034551_, _034552_, _034553_, _034554_, _034555_, _034556_, _034557_, _034558_, _034559_, _034560_, _034561_, _034562_, _034563_, _034564_, _034565_, _034566_, _034567_, _034568_, _034569_, _034570_, _034571_, _034572_, _034573_, _034574_, _034575_, _034576_, _034577_, _034578_, _034579_, _034580_, _034581_, _034582_, _034583_, _034584_, _034585_, _034586_, _034587_, _034588_, _034589_, _034590_, _034591_, _034592_, _034593_, _034594_, _034595_, _034596_, _034597_, _034598_, _034599_, _034600_, _034601_, _034602_, _034603_, _034604_, _034605_, _034606_, _034607_, _034608_, _034609_, _034610_, _034611_, _034612_, _034613_, _034614_, _034615_, _034616_, _034617_, _034618_, _034619_, _034620_, _034621_, _034622_, _034623_, _034624_, _034625_, _034626_, _034627_, _034628_, _034629_, _034630_, _034631_, _034632_, _034633_, _034634_, _034635_, _034636_, _034637_, _034638_, _034639_, _034640_, _034641_, _034642_, _034643_, _034644_, _034645_, _034646_, _034647_, _034648_, _034649_, _034650_, _034651_, _034652_, _034653_, _034654_, _034655_, _034656_, _034657_, _034658_, _034659_, _034660_, _034661_, _034662_, _034663_, _034664_, _034665_, _034666_, _034667_, _034668_, _034669_, _034670_, _034671_, _034672_, _034673_, _034674_, _034675_, _034676_, _034677_, _034678_, _034679_, _034680_, _034681_, _034682_, _034683_, _034684_, _034685_, _034686_, _034687_, _034688_, _034689_, _034690_, _034691_, _034692_, _034693_, _034694_, _034695_, _034696_, _034697_, _034698_, _034699_, _034700_, _034701_, _034702_, _034703_, _034704_, _034705_, _034706_, _034707_, _034708_, _034709_, _034710_, _034711_, _034712_, _034713_, _034714_, _034715_, _034716_, _034717_, _034718_, _034719_, _034720_, _034721_, _034722_, _034723_, _034724_, _034725_, _034726_, _034727_, _034728_, _034729_, _034730_, _034731_, _034732_, _034733_, _034734_, _034735_, _034736_, _034737_, _034738_, _034739_, _034740_, _034741_, _034742_, _034743_, _034744_, _034745_, _034746_, _034747_, _034748_, _034749_, _034750_, _034751_, _034752_, _034753_, _034754_, _034755_, _034756_, _034757_, _034758_, _034759_, _034760_, _034761_, _034762_, _034763_, _034764_, _034765_, _034766_, _034767_, _034768_, _034769_, _034770_, _034771_, _034772_, _034773_, _034774_, _034775_, _034776_, _034777_, _034778_, _034779_, _034780_, _034781_, _034782_, _034783_, _034784_, _034785_, _034786_, _034787_, _034788_, _034789_, _034790_, _034791_, _034792_, _034793_, _034794_, _034795_, _034796_, _034797_, _034798_, _034799_, _034800_, _034801_, _034802_, _034803_, _034804_, _034805_, _034806_, _034807_, _034808_, _034809_, _034810_, _034811_, _034812_, _034813_, _034814_, _034815_, _034816_, _034817_, _034818_, _034819_, _034820_, _034821_, _034822_, _034823_, _034824_, _034825_, _034826_, _034827_, _034828_, _034829_, _034830_, _034831_, _034832_, _034833_, _034834_, _034835_, _034836_, _034837_, _034838_, _034839_, _034840_, _034841_, _034842_, _034843_, _034844_, _034845_, _034846_, _034847_, _034848_, _034849_, _034850_, _034851_, _034852_, _034853_, _034854_, _034855_, _034856_, _034857_, _034858_, _034859_, _034860_, _034861_, _034862_, _034863_, _034864_, _034865_, _034866_, _034867_, _034868_, _034869_, _034870_, _034871_, _034872_, _034873_, _034874_, _034875_, _034876_, _034877_, _034878_, _034879_, _034880_, _034881_, _034882_, _034883_, _034884_, _034885_, _034886_, _034887_, _034888_, _034889_, _034890_, _034891_, _034892_, _034893_, _034894_, _034895_, _034896_, _034897_, _034898_, _034899_, _034900_, _034901_, _034902_, _034903_, _034904_, _034905_, _034906_, _034907_, _034908_, _034909_, _034910_, _034911_, _034912_, _034913_, _034914_, _034915_, _034916_, _034917_, _034918_, _034919_, _034920_, _034921_, _034922_, _034923_, _034924_, _034925_, _034926_, _034927_, _034928_, _034929_, _034930_, _034931_, _034932_, _034933_, _034934_, _034935_, _034936_, _034937_, _034938_, _034939_, _034940_, _034941_, _034942_, _034943_, _034944_, _034945_, _034946_, _034947_, _034948_, _034949_, _034950_, _034951_, _034952_, _034953_, _034954_, _034955_, _034956_, _034957_, _034958_, _034959_, _034960_, _034961_, _034962_, _034963_, _034964_, _034965_, _034966_, _034967_, _034968_, _034969_, _034970_, _034971_, _034972_, _034973_, _034974_, _034975_, _034976_, _034977_, _034978_, _034979_, _034980_, _034981_, _034982_, _034983_, _034984_, _034985_, _034986_, _034987_, _034988_, _034989_, _034990_, _034991_, _034992_, _034993_, _034994_, _034995_, _034996_, _034997_, _034998_, _034999_, _035000_, _035001_, _035002_, _035003_, _035004_, _035005_, _035006_, _035007_, _035008_, _035009_, _035010_, _035011_, _035012_, _035013_, _035014_, _035015_, _035016_, _035017_, _035018_, _035019_, _035020_, _035021_, _035022_, _035023_, _035024_, _035025_, _035026_, _035027_, _035028_, _035029_, _035030_, _035031_, _035032_, _035033_, _035034_, _035035_, _035036_, _035037_, _035038_, _035039_, _035040_, _035041_, _035042_, _035043_, _035044_, _035045_, _035046_, _035047_, _035048_, _035049_, _035050_, _035051_, _035052_, _035053_, _035054_, _035055_, _035056_, _035057_, _035058_, _035059_, _035060_, _035061_, _035062_, _035063_, _035064_, _035065_, _035066_, _035067_, _035068_, _035069_, _035070_, _035071_, _035072_, _035073_, _035074_, _035075_, _035076_, _035077_, _035078_, _035079_, _035080_, _035081_, _035082_, _035083_, _035084_, _035085_, _035086_, _035087_, _035088_, _035089_, _035090_, _035091_, _035092_, _035093_, _035094_, _035095_, _035096_, _035097_, _035098_, _035099_, _035100_, _035101_, _035102_, _035103_, _035104_, _035105_, _035106_, _035107_, _035108_, _035109_, _035110_, _035111_, _035112_, _035113_, _035114_, _035115_, _035116_, _035117_, _035118_, _035119_, _035120_, _035121_, _035122_, _035123_, _035124_, _035125_, _035126_, _035127_, _035128_, _035129_, _035130_, _035131_, _035132_, _035133_, _035134_, _035135_, _035136_, _035137_, _035138_, _035139_, _035140_, _035141_, _035142_, _035143_, _035144_, _035145_, _035146_, _035147_, _035148_, _035149_, _035150_, _035151_, _035152_, _035153_, _035154_, _035155_, _035156_, _035157_, _035158_, _035159_, _035160_, _035161_, _035162_, _035163_, _035164_, _035165_, _035166_, _035167_, _035168_, _035169_, _035170_, _035171_, _035172_, _035173_, _035174_, _035175_, _035176_, _035177_, _035178_, _035179_, _035180_, _035181_, _035182_, _035183_, _035184_, _035185_, _035186_, _035187_, _035188_, _035189_, _035190_, _035191_, _035192_, _035193_, _035194_, _035195_, _035196_, _035197_, _035198_, _035199_, _035200_, _035201_, _035202_, _035203_, _035204_, _035205_, _035206_, _035207_, _035208_, _035209_, _035210_, _035211_, _035212_, _035213_, _035214_, _035215_, _035216_, _035217_, _035218_, _035219_, _035220_, _035221_, _035222_, _035223_, _035224_, _035225_, _035226_, _035227_, _035228_, _035229_, _035230_, _035231_, _035232_, _035233_, _035234_, _035235_, _035236_, _035237_, _035238_, _035239_, _035240_, _035241_, _035242_, _035243_, _035244_, _035245_, _035246_, _035247_, _035248_, _035249_, _035250_, _035251_, _035252_, _035253_, _035254_, _035255_, _035256_, _035257_, _035258_, _035259_, _035260_, _035261_, _035262_, _035263_, _035264_, _035265_, _035266_, _035267_, _035268_, _035269_, _035270_, _035271_, _035272_, _035273_, _035274_, _035275_, _035276_, _035277_, _035278_, _035279_, _035280_, _035281_, _035282_, _035283_, _035284_, _035285_, _035286_, _035287_, _035288_, _035289_, _035290_, _035291_, _035292_, _035293_, _035294_, _035295_, _035296_, _035297_, _035298_, _035299_, _035300_, _035301_, _035302_, _035303_, _035304_, _035305_, _035306_, _035307_, _035308_, _035309_, _035310_, _035311_, _035312_, _035313_, _035314_, _035315_, _035316_, _035317_, _035318_, _035319_, _035320_, _035321_, _035322_, _035323_, _035324_, _035325_, _035326_, _035327_, _035328_, _035329_, _035330_, _035331_, _035332_, _035333_, _035334_, _035335_, _035336_, _035337_, _035338_, _035339_, _035340_, _035341_, _035342_, _035343_, _035344_, _035345_, _035346_, _035347_, _035348_, _035349_, _035350_, _035351_, _035352_, _035353_, _035354_, _035355_, _035356_, _035357_, _035358_, _035359_, _035360_, _035361_, _035362_, _035363_, _035364_, _035365_, _035366_, _035367_, _035368_, _035369_, _035370_, _035371_, _035372_, _035373_, _035374_, _035375_, _035376_, _035377_, _035378_, _035379_, _035380_, _035381_, _035382_, _035383_, _035384_, _035385_, _035386_, _035387_, _035388_, _035389_, _035390_, _035391_, _035392_, _035393_, _035394_, _035395_, _035396_, _035397_, _035398_, _035399_, _035400_, _035401_, _035402_, _035403_, _035404_, _035405_, _035406_, _035407_, _035408_, _035409_, _035410_, _035411_, _035412_, _035413_, _035414_, _035415_, _035416_, _035417_, _035418_, _035419_, _035420_, _035421_, _035422_, _035423_, _035424_, _035425_, _035426_, _035427_, _035428_, _035429_, _035430_, _035431_, _035432_, _035433_, _035434_, _035435_, _035436_, _035437_, _035438_, _035439_, _035440_, _035441_, _035442_, _035443_, _035444_, _035445_, _035446_, _035447_, _035448_, _035449_, _035450_, _035451_, _035452_, _035453_, _035454_, _035455_, _035456_, _035457_, _035458_, _035459_, _035460_, _035461_, _035462_, _035463_, _035464_, _035465_, _035466_, _035467_, _035468_, _035469_, _035470_, _035471_, _035472_, _035473_, _035474_, _035475_, _035476_, _035477_, _035478_, _035479_, _035480_, _035481_, _035482_, _035483_, _035484_, _035485_, _035486_, _035487_, _035488_, _035489_, _035490_, _035491_, _035492_, _035493_, _035494_, _035495_, _035496_, _035497_, _035498_, _035499_, _035500_, _035501_, _035502_, _035503_, _035504_, _035505_, _035506_, _035507_, _035508_, _035509_, _035510_, _035511_, _035512_, _035513_, _035514_, _035515_, _035516_, _035517_, _035518_, _035519_, _035520_, _035521_, _035522_, _035523_, _035524_, _035525_, _035526_, _035527_, _035528_, _035529_, _035530_, _035531_, _035532_, _035533_, _035534_, _035535_, _035536_, _035537_, _035538_, _035539_, _035540_, _035541_, _035542_, _035543_, _035544_, _035545_, _035546_, _035547_, _035548_, _035549_, _035550_, _035551_, _035552_, _035553_, _035554_, _035555_, _035556_, _035557_, _035558_, _035559_, _035560_, _035561_, _035562_, _035563_, _035564_, _035565_, _035566_, _035567_, _035568_, _035569_, _035570_, _035571_, _035572_, _035573_, _035574_, _035575_, _035576_, _035577_, _035578_, _035579_, _035580_, _035581_, _035582_, _035583_, _035584_, _035585_, _035586_, _035587_, _035588_, _035589_, _035590_, _035591_, _035592_, _035593_, _035594_, _035595_, _035596_, _035597_, _035598_, _035599_, _035600_, _035601_, _035602_, _035603_, _035604_, _035605_, _035606_, _035607_, _035608_, _035609_, _035610_, _035611_, _035612_, _035613_, _035614_, _035615_, _035616_, _035617_, _035618_, _035619_, _035620_, _035621_, _035622_, _035623_, _035624_, _035625_, _035626_, _035627_, _035628_, _035629_, _035630_, _035631_, _035632_, _035633_, _035634_, _035635_, _035636_, _035637_, _035638_, _035639_, _035640_, _035641_, _035642_, _035643_, _035644_, _035645_, _035646_, _035647_, _035648_, _035649_, _035650_, _035651_, _035652_, _035653_, _035654_, _035655_, _035656_, _035657_, _035658_, _035659_, _035660_, _035661_, _035662_, _035663_, _035664_, _035665_, _035666_, _035667_, _035668_, _035669_, _035670_, _035671_, _035672_, _035673_, _035674_, _035675_, _035676_, _035677_, _035678_, _035679_, _035680_, _035681_, _035682_, _035683_, _035684_, _035685_, _035686_, _035687_, _035688_, _035689_, _035690_, _035691_, _035692_, _035693_, _035694_, _035695_, _035696_, _035697_, _035698_, _035699_, _035700_, _035701_, _035702_, _035703_, _035704_, _035705_, _035706_, _035707_, _035708_, _035709_, _035710_, _035711_, _035712_, _035713_, _035714_, _035715_, _035716_, _035717_, _035718_, _035719_, _035720_, _035721_, _035722_, _035723_, _035724_, _035725_, _035726_, _035727_, _035728_, _035729_, _035730_, _035731_, _035732_, _035733_, _035734_, _035735_, _035736_, _035737_, _035738_, _035739_, _035740_, _035741_, _035742_, _035743_, _035744_, _035745_, _035746_, _035747_, _035748_, _035749_, _035750_, _035751_, _035752_, _035753_, _035754_, _035755_, _035756_, _035757_, _035758_, _035759_, _035760_, _035761_, _035762_, _035763_, _035764_, _035765_, _035766_, _035767_, _035768_, _035769_, _035770_, _035771_, _035772_, _035773_, _035774_, _035775_, _035776_, _035777_, _035778_, _035779_, _035780_, _035781_, _035782_, _035783_, _035784_, _035785_, _035786_, _035787_, _035788_, _035789_, _035790_, _035791_, _035792_, _035793_, _035794_, _035795_, _035796_, _035797_, _035798_, _035799_, _035800_, _035801_, _035802_, _035803_, _035804_, _035805_, _035806_, _035807_, _035808_, _035809_, _035810_, _035811_, _035812_, _035813_, _035814_, _035815_, _035816_, _035817_, _035818_, _035819_, _035820_, _035821_, _035822_, _035823_, _035824_, _035825_, _035826_, _035827_, _035828_, _035829_, _035830_, _035831_, _035832_, _035833_, _035834_, _035835_, _035836_, _035837_, _035838_, _035839_, _035840_, _035841_, _035842_, _035843_, _035844_, _035845_, _035846_, _035847_, _035848_, _035849_, _035850_, _035851_, _035852_, _035853_, _035854_, _035855_, _035856_, _035857_, _035858_, _035859_, _035860_, _035861_, _035862_, _035863_, _035864_, _035865_, _035866_, _035867_, _035868_, _035869_, _035870_, _035871_, _035872_, _035873_, _035874_, _035875_, _035876_, _035877_, _035878_, _035879_, _035880_, _035881_, _035882_, _035883_, _035884_, _035885_, _035886_, _035887_, _035888_, _035889_, _035890_, _035891_, _035892_, _035893_, _035894_, _035895_, _035896_, _035897_, _035898_, _035899_, _035900_, _035901_, _035902_, _035903_, _035904_, _035905_, _035906_, _035907_, _035908_, _035909_, _035910_, _035911_, _035912_, _035913_, _035914_, _035915_, _035916_, _035917_, _035918_, _035919_, _035920_, _035921_, _035922_, _035923_, _035924_, _035925_, _035926_, _035927_, _035928_, _035929_, _035930_, _035931_, _035932_, _035933_, _035934_, _035935_, _035936_, _035937_, _035938_, _035939_, _035940_, _035941_, _035942_, _035943_, _035944_, _035945_, _035946_, _035947_, _035948_, _035949_, _035950_, _035951_, _035952_, _035953_, _035954_, _035955_, _035956_, _035957_, _035958_, _035959_, _035960_, _035961_, _035962_, _035963_, _035964_, _035965_, _035966_, _035967_, _035968_, _035969_, _035970_, _035971_, _035972_, _035973_, _035974_, _035975_, _035976_, _035977_, _035978_, _035979_, _035980_, _035981_, _035982_, _035983_, _035984_, _035985_, _035986_, _035987_, _035988_, _035989_, _035990_, _035991_, _035992_, _035993_, _035994_, _035995_, _035996_, _035997_, _035998_, _035999_, _036000_, _036001_, _036002_, _036003_, _036004_, _036005_, _036006_, _036007_, _036008_, _036009_, _036010_, _036011_, _036012_, _036013_, _036014_, _036015_, _036016_, _036017_, _036018_, _036019_, _036020_, _036021_, _036022_, _036023_, _036024_, _036025_, _036026_, _036027_, _036028_, _036029_, _036030_, _036031_, _036032_, _036033_, _036034_, _036035_, _036036_, _036037_, _036038_, _036039_, _036040_, _036041_, _036042_, _036043_, _036044_, _036045_, _036046_, _036047_, _036048_, _036049_, _036050_, _036051_, _036052_, _036053_, _036054_, _036055_, _036056_, _036057_, _036058_, _036059_, _036060_, _036061_, _036062_, _036063_, _036064_, _036065_, _036066_, _036067_, _036068_, _036069_, _036070_, _036071_, _036072_, _036073_, _036074_, _036075_, _036076_, _036077_, _036078_, _036079_, _036080_, _036081_, _036082_, _036083_, _036084_, _036085_, _036086_, _036087_, _036088_, _036089_, _036090_, _036091_, _036092_, _036093_, _036094_, _036095_, _036096_, _036097_, _036098_, _036099_, _036100_, _036101_, _036102_, _036103_, _036104_, _036105_, _036106_, _036107_, _036108_, _036109_, _036110_, _036111_, _036112_, _036113_, _036114_, _036115_, _036116_, _036117_, _036118_, _036119_, _036120_, _036121_, _036122_, _036123_, _036124_, _036125_, _036126_, _036127_, _036128_, _036129_, _036130_, _036131_, _036132_, _036133_, _036134_, _036135_, _036136_, _036137_, _036138_, _036139_, _036140_, _036141_, _036142_, _036143_, _036144_, _036145_, _036146_, _036147_, _036148_, _036149_, _036150_, _036151_, _036152_, _036153_, _036154_, _036155_, _036156_, _036157_, _036158_, _036159_, _036160_, _036161_, _036162_, _036163_, _036164_, _036165_, _036166_, _036167_, _036168_, _036169_, _036170_, _036171_, _036172_, _036173_, _036174_, _036175_, _036176_, _036177_, _036178_, _036179_, _036180_, _036181_, _036182_, _036183_, _036184_, _036185_, _036186_, _036187_, _036188_, _036189_, _036190_, _036191_, _036192_, _036193_, _036194_, _036195_, _036196_, _036197_, _036198_, _036199_, _036200_, _036201_, _036202_, _036203_, _036204_, _036205_, _036206_, _036207_, _036208_, _036209_, _036210_, _036211_, _036212_, _036213_, _036214_, _036215_, _036216_, _036217_, _036218_, _036219_, _036220_, _036221_, _036222_, _036223_, _036224_, _036225_, _036226_, _036227_, _036228_, _036229_, _036230_, _036231_, _036232_, _036233_, _036234_, _036235_, _036236_, _036237_, _036238_, _036239_, _036240_, _036241_, _036242_, _036243_, _036244_, _036245_, _036246_, _036247_, _036248_, _036249_, _036250_, _036251_, _036252_, _036253_, _036254_, _036255_, _036256_, _036257_, _036258_, _036259_, _036260_, _036261_, _036262_, _036263_, _036264_, _036265_, _036266_, _036267_, _036268_, _036269_, _036270_, _036271_, _036272_, _036273_, _036274_, _036275_, _036276_, _036277_, _036278_, _036279_, _036280_, _036281_, _036282_, _036283_, _036284_, _036285_, _036286_, _036287_, _036288_, _036289_, _036290_, _036291_, _036292_, _036293_, _036294_, _036295_, _036296_, _036297_, _036298_, _036299_, _036300_, _036301_, _036302_, _036303_, _036304_, _036305_, _036306_, _036307_, _036308_, _036309_, _036310_, _036311_, _036312_, _036313_, _036314_, _036315_, _036316_, _036317_, _036318_, _036319_, _036320_, _036321_, _036322_, _036323_, _036324_, _036325_, _036326_, _036327_, _036328_, _036329_, _036330_, _036331_, _036332_, _036333_, _036334_, _036335_, _036336_, _036337_, _036338_, _036339_, _036340_, _036341_, _036342_, _036343_, _036344_, _036345_, _036346_, _036347_, _036348_, _036349_, _036350_, _036351_, _036352_, _036353_, _036354_, _036355_, _036356_, _036357_, _036358_, _036359_, _036360_, _036361_, _036362_, _036363_, _036364_, _036365_, _036366_, _036367_, _036368_, _036369_, _036370_, _036371_, _036372_, _036373_, _036374_, _036375_, _036376_, _036377_, _036378_, _036379_, _036380_, _036381_, _036382_, _036383_, _036384_, _036385_, _036386_, _036387_, _036388_, _036389_, _036390_, _036391_, _036392_, _036393_, _036394_, _036395_, _036396_, _036397_, _036398_, _036399_, _036400_, _036401_, _036402_, _036403_, _036404_, _036405_, _036406_, _036407_, _036408_, _036409_, _036410_, _036411_, _036412_, _036413_, _036414_, _036415_, _036416_, _036417_, _036418_, _036419_, _036420_, _036421_, _036422_, _036423_, _036424_, _036425_, _036426_, _036427_, _036428_, _036429_, _036430_, _036431_, _036432_, _036433_, _036434_, _036435_, _036436_, _036437_, _036438_, _036439_, _036440_, _036441_, _036442_, _036443_, _036444_, _036445_, _036446_, _036447_, _036448_, _036449_, _036450_, _036451_, _036452_, _036453_, _036454_, _036455_, _036456_, _036457_, _036458_, _036459_, _036460_, _036461_, _036462_, _036463_, _036464_, _036465_, _036466_, _036467_, _036468_, _036469_, _036470_, _036471_, _036472_, _036473_, _036474_, _036475_, _036476_, _036477_, _036478_, _036479_, _036480_, _036481_, _036482_, _036483_, _036484_, _036485_, _036486_, _036487_, _036488_, _036489_, _036490_, _036491_, _036492_, _036493_, _036494_, _036495_, _036496_, _036497_, _036498_, _036499_, _036500_, _036501_, _036502_, _036503_, _036504_, _036505_, _036506_, _036507_, _036508_, _036509_, _036510_, _036511_, _036512_, _036513_, _036514_, _036515_, _036516_, _036517_, _036518_, _036519_, _036520_, _036521_, _036522_, _036523_, _036524_, _036525_, _036526_, _036527_, _036528_, _036529_, _036530_, _036531_, _036532_, _036533_, _036534_, _036535_, _036536_, _036537_, _036538_, _036539_, _036540_, _036541_, _036542_, _036543_, _036544_, _036545_, _036546_, _036547_, _036548_, _036549_, _036550_, _036551_, _036552_, _036553_, _036554_, _036555_, _036556_, _036557_, _036558_, _036559_, _036560_, _036561_, _036562_, _036563_, _036564_, _036565_, _036566_, _036567_, _036568_, _036569_, _036570_, _036571_, _036572_, _036573_, _036574_, _036575_, _036576_, _036577_, _036578_, _036579_, _036580_, _036581_, _036582_, _036583_, _036584_, _036585_, _036586_, _036587_, _036588_, _036589_, _036590_, _036591_, _036592_, _036593_, _036594_, _036595_, _036596_, _036597_, _036598_, _036599_, _036600_, _036601_, _036602_, _036603_, _036604_, _036605_, _036606_, _036607_, _036608_, _036609_, _036610_, _036611_, _036612_, _036613_, _036614_, _036615_, _036616_, _036617_, _036618_, _036619_, _036620_, _036621_, _036622_, _036623_, _036624_, _036625_, _036626_, _036627_, _036628_, _036629_, _036630_, _036631_, _036632_, _036633_, _036634_, _036635_, _036636_, _036637_, _036638_, _036639_, _036640_, _036641_, _036642_, _036643_, _036644_, _036645_, _036646_, _036647_, _036648_, _036649_, _036650_, _036651_, _036652_, _036653_, _036654_, _036655_, _036656_, _036657_, _036658_, _036659_, _036660_, _036661_, _036662_, _036663_, _036664_, _036665_, _036666_, _036667_, _036668_, _036669_, _036670_, _036671_, _036672_, _036673_, _036674_, _036675_, _036676_, _036677_, _036678_, _036679_, _036680_, _036681_, _036682_, _036683_, _036684_, _036685_, _036686_, _036687_, _036688_, _036689_, _036690_, _036691_, _036692_, _036693_, _036694_, _036695_, _036696_, _036697_, _036698_, _036699_, _036700_, _036701_, _036702_, _036703_, _036704_, _036705_, _036706_, _036707_, _036708_, _036709_, _036710_, _036711_, _036712_, _036713_, _036714_, _036715_, _036716_, _036717_, _036718_, _036719_, _036720_, _036721_, _036722_, _036723_, _036724_, _036725_, _036726_, _036727_, _036728_, _036729_, _036730_, _036731_, _036732_, _036733_, _036734_, _036735_, _036736_, _036737_, _036738_, _036739_, _036740_, _036741_, _036742_, _036743_, _036744_, _036745_, _036746_, _036747_, _036748_, _036749_, _036750_, _036751_, _036752_, _036753_, _036754_, _036755_, _036756_, _036757_, _036758_, _036759_, _036760_, _036761_, _036762_, _036763_, _036764_, _036765_, _036766_, _036767_, _036768_, _036769_, _036770_, _036771_, _036772_, _036773_, _036774_, _036775_, _036776_, _036777_, _036778_, _036779_, _036780_, _036781_, _036782_, _036783_, _036784_, _036785_, _036786_, _036787_, _036788_, _036789_, _036790_, _036791_, _036792_, _036793_, _036794_, _036795_, _036796_, _036797_, _036798_, _036799_, _036800_, _036801_, _036802_, _036803_, _036804_, _036805_, _036806_, _036807_, _036808_, _036809_, _036810_, _036811_, _036812_, _036813_, _036814_, _036815_, _036816_, _036817_, _036818_, _036819_, _036820_, _036821_, _036822_, _036823_, _036824_, _036825_, _036826_, _036827_, _036828_, _036829_, _036830_, _036831_, _036832_, _036833_, _036834_, _036835_, _036836_, _036837_, _036838_, _036839_, _036840_, _036841_, _036842_, _036843_, _036844_, _036845_, _036846_, _036847_, _036848_, _036849_, _036850_, _036851_, _036852_, _036853_, _036854_, _036855_, _036856_, _036857_, _036858_, _036859_, _036860_, _036861_, _036862_, _036863_, _036864_, _036865_, _036866_, _036867_, _036868_, _036869_, _036870_, _036871_, _036872_, _036873_, _036874_, _036875_, _036876_, _036877_, _036878_, _036879_, _036880_, _036881_, _036882_, _036883_, _036884_, _036885_, _036886_, _036887_, _036888_, _036889_, _036890_, _036891_, _036892_, _036893_, _036894_, _036895_, _036896_, _036897_, _036898_, _036899_, _036900_, _036901_, _036902_, _036903_, _036904_, _036905_, _036906_, _036907_, _036908_, _036909_, _036910_, _036911_, _036912_, _036913_, _036914_, _036915_, _036916_, _036917_, _036918_, _036919_, _036920_, _036921_, _036922_, _036923_, _036924_, _036925_, _036926_, _036927_, _036928_, _036929_, _036930_, _036931_, _036932_, _036933_, _036934_, _036935_, _036936_, _036937_, _036938_, _036939_, _036940_, _036941_, _036942_, _036943_, _036944_, _036945_, _036946_, _036947_, _036948_, _036949_, _036950_, _036951_, _036952_, _036953_, _036954_, _036955_, _036956_, _036957_, _036958_, _036959_, _036960_, _036961_, _036962_, _036963_, _036964_, _036965_, _036966_, _036967_, _036968_, _036969_, _036970_, _036971_, _036972_, _036973_, _036974_, _036975_, _036976_, _036977_, _036978_, _036979_, _036980_, _036981_, _036982_, _036983_, _036984_, _036985_, _036986_, _036987_, _036988_, _036989_, _036990_, _036991_, _036992_, _036993_, _036994_, _036995_, _036996_, _036997_, _036998_, _036999_, _037000_, _037001_, _037002_, _037003_, _037004_, _037005_, _037006_, _037007_, _037008_, _037009_, _037010_, _037011_, _037012_, _037013_, _037014_, _037015_, _037016_, _037017_, _037018_, _037019_, _037020_, _037021_, _037022_, _037023_, _037024_, _037025_, _037026_, _037027_, _037028_, _037029_, _037030_, _037031_, _037032_, _037033_, _037034_, _037035_, _037036_, _037037_, _037038_, _037039_, _037040_, _037041_, _037042_, _037043_, _037044_, _037045_, _037046_, _037047_, _037048_, _037049_, _037050_, _037051_, _037052_, _037053_, _037054_, _037055_, _037056_, _037057_, _037058_, _037059_, _037060_, _037061_, _037062_, _037063_, _037064_, _037065_, _037066_, _037067_, _037068_, _037069_, _037070_, _037071_, _037072_, _037073_, _037074_, _037075_, _037076_, _037077_, _037078_, _037079_, _037080_, _037081_, _037082_, _037083_, _037084_, _037085_, _037086_, _037087_, _037088_, _037089_, _037090_, _037091_, _037092_, _037093_, _037094_, _037095_, _037096_, _037097_, _037098_, _037099_, _037100_, _037101_, _037102_, _037103_, _037104_, _037105_, _037106_, _037107_, _037108_, _037109_, _037110_, _037111_, _037112_, _037113_, _037114_, _037115_, _037116_, _037117_, _037118_, _037119_, _037120_, _037121_, _037122_, _037123_, _037124_, _037125_, _037126_, _037127_, _037128_, _037129_, _037130_, _037131_, _037132_, _037133_, _037134_, _037135_, _037136_, _037137_, _037138_, _037139_, _037140_, _037141_, _037142_, _037143_, _037144_, _037145_, _037146_, _037147_, _037148_, _037149_, _037150_, _037151_, _037152_, _037153_, _037154_, _037155_, _037156_, _037157_, _037158_, _037159_, _037160_, _037161_, _037162_, _037163_, _037164_, _037165_, _037166_, _037167_, _037168_, _037169_, _037170_, _037171_, _037172_, _037173_, _037174_, _037175_, _037176_, _037177_, _037178_, _037179_, _037180_, _037181_, _037182_, _037183_, _037184_, _037185_, _037186_, _037187_, _037188_, _037189_, _037190_, _037191_, _037192_, _037193_, _037194_, _037195_, _037196_, _037197_, _037198_, _037199_, _037200_, _037201_, _037202_, _037203_, _037204_, _037205_, _037206_, _037207_, _037208_, _037209_, _037210_, _037211_, _037212_, _037213_, _037214_, _037215_, _037216_, _037217_, _037218_, _037219_, _037220_, _037221_, _037222_, _037223_, _037224_, _037225_, _037226_, _037227_, _037228_, _037229_, _037230_, _037231_, _037232_, _037233_, _037234_, _037235_, _037236_, _037237_, _037238_, _037239_, _037240_, _037241_, _037242_, _037243_, _037244_, _037245_, _037246_, _037247_, _037248_, _037249_, _037250_, _037251_, _037252_, _037253_, _037254_, _037255_, _037256_, _037257_, _037258_, _037259_, _037260_, _037261_, _037262_, _037263_, _037264_, _037265_, _037266_, _037267_, _037268_, _037269_, _037270_, _037271_, _037272_, _037273_, _037274_, _037275_, _037276_, _037277_, _037278_, _037279_, _037280_, _037281_, _037282_, _037283_, _037284_, _037285_, _037286_, _037287_, _037288_, _037289_, _037290_, _037291_, _037292_, _037293_, _037294_, _037295_, _037296_, _037297_, _037298_, _037299_, _037300_, _037301_, _037302_, _037303_, _037304_, _037305_, _037306_, _037307_, _037308_, _037309_, _037310_, _037311_, _037312_, _037313_, _037314_, _037315_, _037316_, _037317_, _037318_, _037319_, _037320_, _037321_, _037322_, _037323_, _037324_, _037325_, _037326_, _037327_, _037328_, _037329_, _037330_, _037331_, _037332_, _037333_, _037334_, _037335_, _037336_, _037337_, _037338_, _037339_, _037340_, _037341_, _037342_, _037343_, _037344_, _037345_, _037346_, _037347_, _037348_, _037349_, _037350_, _037351_, _037352_, _037353_, _037354_, _037355_, _037356_, _037357_, _037358_, _037359_, _037360_, _037361_, _037362_, _037363_, _037364_, _037365_, _037366_, _037367_, _037368_, _037369_, _037370_, _037371_, _037372_, _037373_, _037374_, _037375_, _037376_, _037377_, _037378_, _037379_, _037380_, _037381_, _037382_, _037383_, _037384_, _037385_, _037386_, _037387_, _037388_, _037389_, _037390_, _037391_, _037392_, _037393_, _037394_, _037395_, _037396_, _037397_, _037398_, _037399_, _037400_, _037401_, _037402_, _037403_, _037404_, _037405_, _037406_, _037407_, _037408_, _037409_, _037410_, _037411_, _037412_, _037413_, _037414_, _037415_, _037416_, _037417_, _037418_, _037419_, _037420_, _037421_, _037422_, _037423_, _037424_, _037425_, _037426_, _037427_, _037428_, _037429_, _037430_, _037431_, _037432_, _037433_, _037434_, _037435_, _037436_, _037437_, _037438_, _037439_, _037440_, _037441_, _037442_, _037443_, _037444_, _037445_, _037446_, _037447_, _037448_, _037449_, _037450_, _037451_, _037452_, _037453_, _037454_, _037455_, _037456_, _037457_, _037458_, _037459_, _037460_, _037461_, _037462_, _037463_, _037464_, _037465_, _037466_, _037467_, _037468_, _037469_, _037470_, _037471_, _037472_, _037473_, _037474_, _037475_, _037476_, _037477_, _037478_, _037479_, _037480_, _037481_, _037482_, _037483_, _037484_, _037485_, _037486_, _037487_, _037488_, _037489_, _037490_, _037491_, _037492_, _037493_, _037494_, _037495_, _037496_, _037497_, _037498_, _037499_, _037500_, _037501_, _037502_, _037503_, _037504_, _037505_, _037506_, _037507_, _037508_, _037509_, _037510_, _037511_, _037512_, _037513_, _037514_, _037515_, _037516_, _037517_, _037518_, _037519_, _037520_, _037521_, _037522_, _037523_, _037524_, _037525_, _037526_, _037527_, _037528_, _037529_, _037530_, _037531_, _037532_, _037533_, _037534_, _037535_, _037536_, _037537_, _037538_, _037539_, _037540_, _037541_, _037542_, _037543_, _037544_, _037545_, _037546_, _037547_, _037548_, _037549_, _037550_, _037551_, _037552_, _037553_, _037554_, _037555_, _037556_, _037557_, _037558_, _037559_, _037560_, _037561_, _037562_, _037563_, _037564_, _037565_, _037566_, _037567_, _037568_, _037569_, _037570_, _037571_, _037572_, _037573_, _037574_, _037575_, _037576_, _037577_, _037578_, _037579_, _037580_, _037581_, _037582_, _037583_, _037584_, _037585_, _037586_, _037587_, _037588_, _037589_, _037590_, _037591_, _037592_, _037593_, _037594_, _037595_, _037596_, _037597_, _037598_, _037599_, _037600_, _037601_, _037602_, _037603_, _037604_, _037605_, _037606_, _037607_, _037608_, _037609_, _037610_, _037611_, _037612_, _037613_, _037614_, _037615_, _037616_, _037617_, _037618_, _037619_, _037620_, _037621_, _037622_, _037623_, _037624_, _037625_, _037626_, _037627_, _037628_, _037629_, _037630_, _037631_, _037632_, _037633_, _037634_, _037635_, _037636_, _037637_, _037638_, _037639_, _037640_, _037641_, _037642_, _037643_, _037644_, _037645_, _037646_, _037647_, _037648_, _037649_, _037650_, _037651_, _037652_, _037653_, _037654_, _037655_, _037656_, _037657_, _037658_, _037659_, _037660_, _037661_, _037662_, _037663_, _037664_, _037665_, _037666_, _037667_, _037668_, _037669_, _037670_, _037671_, _037672_, _037673_, _037674_, _037675_, _037676_, _037677_, _037678_, _037679_, _037680_, _037681_, _037682_, _037683_, _037684_, _037685_, _037686_, _037687_, _037688_, _037689_, _037690_, _037691_, _037692_, _037693_, _037694_, _037695_, _037696_, _037697_, _037698_, _037699_, _037700_, _037701_, _037702_, _037703_, _037704_, _037705_, _037706_, _037707_, _037708_, _037709_, _037710_, _037711_, _037712_, _037713_, _037714_, _037715_, _037716_, _037717_, _037718_, _037719_, _037720_, _037721_, _037722_, _037723_, _037724_, _037725_, _037726_, _037727_, _037728_, _037729_, _037730_, _037731_, _037732_, _037733_, _037734_, _037735_, _037736_, _037737_, _037738_, _037739_, _037740_, _037741_, _037742_, _037743_, _037744_, _037745_, _037746_, _037747_, _037748_, _037749_, _037750_, _037751_, _037752_, _037753_, _037754_, _037755_, _037756_, _037757_, _037758_, _037759_, _037760_, _037761_, _037762_, _037763_, _037764_, _037765_, _037766_, _037767_, _037768_, _037769_, _037770_, _037771_, _037772_, _037773_, _037774_, _037775_, _037776_, _037777_, _037778_, _037779_, _037780_, _037781_, _037782_, _037783_, _037784_, _037785_, _037786_, _037787_, _037788_, _037789_, _037790_, _037791_, _037792_, _037793_, _037794_, _037795_, _037796_, _037797_, _037798_, _037799_, _037800_, _037801_, _037802_, _037803_, _037804_, _037805_, _037806_, _037807_, _037808_, _037809_, _037810_, _037811_, _037812_, _037813_, _037814_, _037815_, _037816_, _037817_, _037818_, _037819_, _037820_, _037821_, _037822_, _037823_, _037824_, _037825_, _037826_, _037827_, _037828_, _037829_, _037830_, _037831_, _037832_, _037833_, _037834_, _037835_, _037836_, _037837_, _037838_, _037839_, _037840_, _037841_, _037842_, _037843_, _037844_, _037845_, _037846_, _037847_, _037848_, _037849_, _037850_, _037851_, _037852_, _037853_, _037854_, _037855_, _037856_, _037857_, _037858_, _037859_, _037860_, _037861_, _037862_, _037863_, _037864_, _037865_, _037866_, _037867_, _037868_, _037869_, _037870_, _037871_, _037872_, _037873_, _037874_, _037875_, _037876_, _037877_, _037878_, _037879_, _037880_, _037881_, _037882_, _037883_, _037884_, _037885_, _037886_, _037887_, _037888_, _037889_, _037890_, _037891_, _037892_, _037893_, _037894_, _037895_, _037896_, _037897_, _037898_, _037899_, _037900_, _037901_, _037902_, _037903_, _037904_, _037905_, _037906_, _037907_, _037908_, _037909_, _037910_, _037911_, _037912_, _037913_, _037914_, _037915_, _037916_, _037917_, _037918_, _037919_, _037920_, _037921_, _037922_, _037923_, _037924_, _037925_, _037926_, _037927_, _037928_, _037929_, _037930_, _037931_, _037932_, _037933_, _037934_, _037935_, _037936_, _037937_, _037938_, _037939_, _037940_, _037941_, _037942_, _037943_, _037944_, _037945_, _037946_, _037947_, _037948_, _037949_, _037950_, _037951_, _037952_, _037953_, _037954_, _037955_, _037956_, _037957_, _037958_, _037959_, _037960_, _037961_, _037962_, _037963_, _037964_, _037965_, _037966_, _037967_, _037968_, _037969_, _037970_, _037971_, _037972_, _037973_, _037974_, _037975_, _037976_, _037977_, _037978_, _037979_, _037980_, _037981_, _037982_, _037983_, _037984_, _037985_, _037986_, _037987_, _037988_, _037989_, _037990_, _037991_, _037992_, _037993_, _037994_, _037995_, _037996_, _037997_, _037998_, _037999_, _038000_, _038001_, _038002_, _038003_, _038004_, _038005_, _038006_, _038007_, _038008_, _038009_, _038010_, _038011_, _038012_, _038013_, _038014_, _038015_, _038016_, _038017_, _038018_, _038019_, _038020_, _038021_, _038022_, _038023_, _038024_, _038025_, _038026_, _038027_, _038028_, _038029_, _038030_, _038031_, _038032_, _038033_, _038034_, _038035_, _038036_, _038037_, _038038_, _038039_, _038040_, _038041_, _038042_, _038043_, _038044_, _038045_, _038046_, _038047_, _038048_, _038049_, _038050_, _038051_, _038052_, _038053_, _038054_, _038055_, _038056_, _038057_, _038058_, _038059_, _038060_, _038061_, _038062_, _038063_, _038064_, _038065_, _038066_, _038067_, _038068_, _038069_, _038070_, _038071_, _038072_, _038073_, _038074_, _038075_, _038076_, _038077_, _038078_, _038079_, _038080_, _038081_, _038082_, _038083_, _038084_, _038085_, _038086_, _038087_, _038088_, _038089_, _038090_, _038091_, _038092_, _038093_, _038094_, _038095_, _038096_, _038097_, _038098_, _038099_, _038100_, _038101_, _038102_, _038103_, _038104_, _038105_, _038106_, _038107_, _038108_, _038109_, _038110_, _038111_, _038112_, _038113_, _038114_, _038115_, _038116_, _038117_, _038118_, _038119_, _038120_, _038121_, _038122_, _038123_, _038124_, _038125_, _038126_, _038127_, _038128_, _038129_, _038130_, _038131_, _038132_, _038133_, _038134_, _038135_, _038136_, _038137_, _038138_, _038139_, _038140_, _038141_, _038142_, _038143_, _038144_, _038145_, _038146_, _038147_, _038148_, _038149_, _038150_, _038151_, _038152_, _038153_, _038154_, _038155_, _038156_, _038157_, _038158_, _038159_, _038160_, _038161_, _038162_, _038163_, _038164_, _038165_, _038166_, _038167_, _038168_, _038169_, _038170_, _038171_, _038172_, _038173_, _038174_, _038175_, _038176_, _038177_, _038178_, _038179_, _038180_, _038181_, _038182_, _038183_, _038184_, _038185_, _038186_, _038187_, _038188_, _038189_, _038190_, _038191_, _038192_, _038193_, _038194_, _038195_, _038196_, _038197_, _038198_, _038199_, _038200_, _038201_, _038202_, _038203_, _038204_, _038205_, _038206_, _038207_, _038208_, _038209_, _038210_, _038211_, _038212_, _038213_, _038214_, _038215_, _038216_, _038217_, _038218_, _038219_, _038220_, _038221_, _038222_, _038223_, _038224_, _038225_, _038226_, _038227_, _038228_, _038229_, _038230_, _038231_, _038232_, _038233_, _038234_, _038235_, _038236_, _038237_, _038238_, _038239_, _038240_, _038241_, _038242_, _038243_, _038244_, _038245_, _038246_, _038247_, _038248_, _038249_, _038250_, _038251_, _038252_, _038253_, _038254_, _038255_, _038256_, _038257_, _038258_, _038259_, _038260_, _038261_, _038262_, _038263_, _038264_, _038265_, _038266_, _038267_, _038268_, _038269_, _038270_, _038271_, _038272_, _038273_, _038274_, _038275_, _038276_, _038277_, _038278_, _038279_, _038280_, _038281_, _038282_, _038283_, _038284_, _038285_, _038286_, _038287_, _038288_, _038289_, _038290_, _038291_, _038292_, _038293_, _038294_, _038295_, _038296_, _038297_, _038298_, _038299_, _038300_, _038301_, _038302_, _038303_, _038304_, _038305_, _038306_, _038307_, _038308_, _038309_, _038310_, _038311_, _038312_, _038313_, _038314_, _038315_, _038316_, _038317_, _038318_, _038319_, _038320_, _038321_, _038322_, _038323_, _038324_, _038325_, _038326_, _038327_, _038328_, _038329_, _038330_, _038331_, _038332_, _038333_, _038334_, _038335_, _038336_, _038337_, _038338_, _038339_, _038340_, _038341_, _038342_, _038343_, _038344_, _038345_, _038346_, _038347_, _038348_, _038349_, _038350_, _038351_, _038352_, _038353_, _038354_, _038355_, _038356_, _038357_, _038358_, _038359_, _038360_, _038361_, _038362_, _038363_, _038364_, _038365_, _038366_, _038367_, _038368_, _038369_, _038370_, _038371_, _038372_, _038373_, _038374_, _038375_, _038376_, _038377_, _038378_, _038379_, _038380_, _038381_, _038382_, _038383_, _038384_, _038385_, _038386_, _038387_, _038388_, _038389_, _038390_, _038391_, _038392_, _038393_, _038394_, _038395_, _038396_, _038397_, _038398_, _038399_, _038400_, _038401_, _038402_, _038403_, _038404_, _038405_, _038406_, _038407_, _038408_, _038409_, _038410_, _038411_, _038412_, _038413_, _038414_, _038415_, _038416_, _038417_, _038418_, _038419_, _038420_, _038421_, _038422_, _038423_, _038424_, _038425_, _038426_, _038427_, _038428_, _038429_, _038430_, _038431_, _038432_, _038433_, _038434_, _038435_, _038436_, _038437_, _038438_, _038439_, _038440_, _038441_, _038442_, _038443_, _038444_, _038445_, _038446_, _038447_, _038448_, _038449_, _038450_, _038451_, _038452_, _038453_, _038454_, _038455_, _038456_, _038457_, _038458_, _038459_, _038460_, _038461_, _038462_, _038463_, _038464_, _038465_, _038466_, _038467_, _038468_, _038469_, _038470_, _038471_, _038472_, _038473_, _038474_, _038475_, _038476_, _038477_, _038478_, _038479_, _038480_, _038481_, _038482_, _038483_, _038484_, _038485_, _038486_, _038487_, _038488_, _038489_, _038490_, _038491_, _038492_, _038493_, _038494_, _038495_, _038496_, _038497_, _038498_, _038499_, _038500_, _038501_, _038502_, _038503_, _038504_, _038505_, _038506_, _038507_, _038508_, _038509_, _038510_, _038511_, _038512_, _038513_, _038514_, _038515_, _038516_, _038517_, _038518_, _038519_, _038520_, _038521_, _038522_, _038523_, _038524_, _038525_, _038526_, _038527_, _038528_, _038529_, _038530_, _038531_, _038532_, _038533_, _038534_, _038535_, _038536_, _038537_, _038538_, _038539_, _038540_, _038541_, _038542_, _038543_, _038544_, _038545_, _038546_, _038547_, _038548_, _038549_, _038550_, _038551_, _038552_, _038553_, _038554_, _038555_, _038556_, _038557_, _038558_, _038559_, _038560_, _038561_, _038562_, _038563_, _038564_, _038565_, _038566_, _038567_, _038568_, _038569_, _038570_, _038571_, _038572_, _038573_, _038574_, _038575_, _038576_, _038577_, _038578_, _038579_, _038580_, _038581_, _038582_, _038583_, _038584_, _038585_, _038586_, _038587_, _038588_, _038589_, _038590_, _038591_, _038592_, _038593_, _038594_, _038595_, _038596_, _038597_, _038598_, _038599_, _038600_, _038601_, _038602_, _038603_, _038604_, _038605_, _038606_, _038607_, _038608_, _038609_, _038610_, _038611_, _038612_, _038613_, _038614_, _038615_, _038616_, _038617_, _038618_, _038619_, _038620_, _038621_, _038622_, _038623_, _038624_, _038625_, _038626_, _038627_, _038628_, _038629_, _038630_, _038631_, _038632_, _038633_, _038634_, _038635_, _038636_, _038637_, _038638_, _038639_, _038640_, _038641_, _038642_, _038643_, _038644_, _038645_, _038646_, _038647_, _038648_, _038649_, _038650_, _038651_, _038652_, _038653_, _038654_, _038655_, _038656_, _038657_, _038658_, _038659_, _038660_, _038661_, _038662_, _038663_, _038664_, _038665_, _038666_, _038667_, _038668_, _038669_, _038670_, _038671_, _038672_, _038673_, _038674_, _038675_, _038676_, _038677_, _038678_, _038679_, _038680_, _038681_, _038682_, _038683_, _038684_, _038685_, _038686_, _038687_, _038688_, _038689_, _038690_, _038691_, _038692_, _038693_, _038694_, _038695_, _038696_, _038697_, _038698_, _038699_, _038700_, _038701_, _038702_, _038703_, _038704_, _038705_, _038706_, _038707_, _038708_, _038709_, _038710_, _038711_, _038712_, _038713_, _038714_, _038715_, _038716_, _038717_, _038718_, _038719_, _038720_, _038721_, _038722_, _038723_, _038724_, _038725_, _038726_, _038727_, _038728_, _038729_, _038730_, _038731_, _038732_, _038733_, _038734_, _038735_, _038736_, _038737_, _038738_, _038739_, _038740_, _038741_, _038742_, _038743_, _038744_, _038745_, _038746_, _038747_, _038748_, _038749_, _038750_, _038751_, _038752_, _038753_, _038754_, _038755_, _038756_, _038757_, _038758_, _038759_, _038760_, _038761_, _038762_, _038763_, _038764_, _038765_, _038766_, _038767_, _038768_, _038769_, _038770_, _038771_, _038772_, _038773_, _038774_, _038775_, _038776_, _038777_, _038778_, _038779_, _038780_, _038781_, _038782_, _038783_, _038784_, _038785_, _038786_, _038787_, _038788_, _038789_, _038790_, _038791_, _038792_, _038793_, _038794_, _038795_, _038796_, _038797_, _038798_, _038799_, _038800_, _038801_, _038802_, _038803_, _038804_, _038805_, _038806_, _038807_, _038808_, _038809_, _038810_, _038811_, _038812_, _038813_, _038814_, _038815_, _038816_, _038817_, _038818_, _038819_, _038820_, _038821_, _038822_, _038823_, _038824_, _038825_, _038826_, _038827_, _038828_, _038829_, _038830_, _038831_, _038832_, _038833_, _038834_, _038835_, _038836_, _038837_, _038838_, _038839_, _038840_, _038841_, _038842_, _038843_, _038844_, _038845_, _038846_, _038847_, _038848_, _038849_, _038850_, _038851_, _038852_, _038853_, _038854_, _038855_, _038856_, _038857_, _038858_, _038859_, _038860_, _038861_, _038862_, _038863_, _038864_, _038865_, _038866_, _038867_, _038868_, _038869_, _038870_, _038871_, _038872_, _038873_, _038874_, _038875_, _038876_, _038877_, _038878_, _038879_, _038880_, _038881_, _038882_, _038883_, _038884_, _038885_, _038886_, _038887_, _038888_, _038889_, _038890_, _038891_, _038892_, _038893_, _038894_, _038895_, _038896_, _038897_, _038898_, _038899_, _038900_, _038901_, _038902_, _038903_, _038904_, _038905_, _038906_, _038907_, _038908_, _038909_, _038910_, _038911_, _038912_, _038913_, _038914_, _038915_, _038916_, _038917_, _038918_, _038919_, _038920_, _038921_, _038922_, _038923_, _038924_, _038925_, _038926_, _038927_, _038928_, _038929_, _038930_, _038931_, _038932_, _038933_, _038934_, _038935_, _038936_, _038937_, _038938_, _038939_, _038940_, _038941_, _038942_, _038943_, _038944_, _038945_, _038946_, _038947_, _038948_, _038949_, _038950_, _038951_, _038952_, _038953_, _038954_, _038955_, _038956_, _038957_, _038958_, _038959_, _038960_, _038961_, _038962_, _038963_, _038964_, _038965_, _038966_, _038967_, _038968_, _038969_, _038970_, _038971_, _038972_, _038973_, _038974_, _038975_, _038976_, _038977_, _038978_, _038979_, _038980_, _038981_, _038982_, _038983_, _038984_, _038985_, _038986_, _038987_, _038988_, _038989_, _038990_, _038991_, _038992_, _038993_, _038994_, _038995_, _038996_, _038997_, _038998_, _038999_, _039000_, _039001_, _039002_, _039003_, _039004_, _039005_, _039006_, _039007_, _039008_, _039009_, _039010_, _039011_, _039012_, _039013_, _039014_, _039015_, _039016_, _039017_, _039018_, _039019_, _039020_, _039021_, _039022_, _039023_, _039024_, _039025_, _039026_, _039027_, _039028_, _039029_, _039030_, _039031_, _039032_, _039033_, _039034_, _039035_, _039036_, _039037_, _039038_, _039039_, _039040_, _039041_, _039042_, _039043_, _039044_, _039045_, _039046_, _039047_, _039048_, _039049_, _039050_, _039051_, _039052_, _039053_, _039054_, _039055_, _039056_, _039057_, _039058_, _039059_, _039060_, _039061_, _039062_, _039063_, _039064_, _039065_, _039066_, _039067_, _039068_, _039069_, _039070_, _039071_, _039072_, _039073_, _039074_, _039075_, _039076_, _039077_, _039078_, _039079_, _039080_, _039081_, _039082_, _039083_, _039084_, _039085_, _039086_, _039087_, _039088_, _039089_, _039090_, _039091_, _039092_, _039093_, _039094_, _039095_, _039096_, _039097_, _039098_, _039099_, _039100_, _039101_, _039102_, _039103_, _039104_, _039105_, _039106_, _039107_, _039108_, _039109_, _039110_, _039111_, _039112_, _039113_, _039114_, _039115_, _039116_, _039117_, _039118_, _039119_, _039120_, _039121_, _039122_, _039123_, _039124_, _039125_, _039126_, _039127_, _039128_, _039129_, _039130_, _039131_, _039132_, _039133_, _039134_, _039135_, _039136_, _039137_, _039138_, _039139_, _039140_, _039141_, _039142_, _039143_, _039144_, _039145_, _039146_, _039147_, _039148_, _039149_, _039150_, _039151_, _039152_, _039153_, _039154_, _039155_, _039156_, _039157_, _039158_, _039159_, _039160_, _039161_, _039162_, _039163_, _039164_, _039165_, _039166_, _039167_, _039168_, _039169_, _039170_, _039171_, _039172_, _039173_, _039174_, _039175_, _039176_, _039177_, _039178_, _039179_, _039180_, _039181_, _039182_, _039183_, _039184_, _039185_, _039186_, _039187_, _039188_, _039189_, _039190_, _039191_, _039192_, _039193_, _039194_, _039195_, _039196_, _039197_, _039198_, _039199_, _039200_, _039201_, _039202_, _039203_, _039204_, _039205_, _039206_, _039207_, _039208_, _039209_, _039210_, _039211_, _039212_, _039213_, _039214_, _039215_, _039216_, _039217_, _039218_, _039219_, _039220_, _039221_, _039222_, _039223_, _039224_, _039225_, _039226_, _039227_, _039228_, _039229_, _039230_, _039231_, _039232_, _039233_, _039234_, _039235_, _039236_, _039237_, _039238_, _039239_, _039240_, _039241_, _039242_, _039243_, _039244_, _039245_, _039246_, _039247_, _039248_, _039249_, _039250_, _039251_, _039252_, _039253_, _039254_, _039255_, _039256_, _039257_, _039258_, _039259_, _039260_, _039261_, _039262_, _039263_, _039264_, _039265_, _039266_, _039267_, _039268_, _039269_, _039270_, _039271_, _039272_, _039273_, _039274_, _039275_, _039276_, _039277_, _039278_, _039279_, _039280_, _039281_, _039282_, _039283_, _039284_, _039285_, _039286_, _039287_, _039288_, _039289_, _039290_, _039291_, _039292_, _039293_, _039294_, _039295_, _039296_, _039297_, _039298_, _039299_, _039300_, _039301_, _039302_, _039303_, _039304_, _039305_, _039306_, _039307_, _039308_, _039309_, _039310_, _039311_, _039312_, _039313_, _039314_, _039315_, _039316_, _039317_, _039318_, _039319_, _039320_, _039321_, _039322_, _039323_, _039324_, _039325_, _039326_, _039327_, _039328_, _039329_, _039330_, _039331_, _039332_, _039333_, _039334_, _039335_, _039336_, _039337_, _039338_, _039339_, _039340_, _039341_, _039342_, _039343_, _039344_, _039345_, _039346_, _039347_, _039348_, _039349_, _039350_, _039351_, _039352_, _039353_, _039354_, _039355_, _039356_, _039357_, _039358_, _039359_, _039360_, _039361_, _039362_, _039363_, _039364_, _039365_, _039366_, _039367_, _039368_, _039369_, _039370_, _039371_, _039372_, _039373_, _039374_, _039375_, _039376_, _039377_, _039378_, _039379_, _039380_, _039381_, _039382_, _039383_, _039384_, _039385_, _039386_, _039387_, _039388_, _039389_, _039390_, _039391_, _039392_, _039393_, _039394_, _039395_, _039396_, _039397_, _039398_, _039399_, _039400_, _039401_, _039402_, _039403_, _039404_, _039405_, _039406_, _039407_, _039408_, _039409_, _039410_, _039411_, _039412_, _039413_, _039414_, _039415_, _039416_, _039417_, _039418_, _039419_, _039420_, _039421_, _039422_, _039423_, _039424_, _039425_, _039426_, _039427_, _039428_, _039429_, _039430_, _039431_, _039432_, _039433_, _039434_, _039435_, _039436_, _039437_, _039438_, _039439_, _039440_, _039441_, _039442_, _039443_, _039444_, _039445_, _039446_, _039447_, _039448_, _039449_, _039450_, _039451_, _039452_, _039453_, _039454_, _039455_, _039456_, _039457_, _039458_, _039459_, _039460_, _039461_, _039462_, _039463_, _039464_, _039465_, _039466_, _039467_, _039468_, _039469_, _039470_, _039471_, _039472_, _039473_, _039474_, _039475_, _039476_, _039477_, _039478_, _039479_, _039480_, _039481_, _039482_, _039483_, _039484_, _039485_, _039486_, _039487_, _039488_, _039489_, _039490_, _039491_, _039492_, _039493_, _039494_, _039495_, _039496_, _039497_, _039498_, _039499_, _039500_, _039501_, _039502_, _039503_, _039504_, _039505_, _039506_, _039507_, _039508_, _039509_, _039510_, _039511_, _039512_, _039513_, _039514_, _039515_, _039516_, _039517_, _039518_, _039519_, _039520_, _039521_, _039522_, _039523_, _039524_, _039525_, _039526_, _039527_, _039528_, _039529_, _039530_, _039531_, _039532_, _039533_, _039534_, _039535_, _039536_, _039537_, _039538_, _039539_, _039540_, _039541_, _039542_, _039543_, _039544_, _039545_, _039546_, _039547_, _039548_, _039549_, _039550_, _039551_, _039552_, _039553_, _039554_, _039555_, _039556_, _039557_, _039558_, _039559_, _039560_, _039561_, _039562_, _039563_, _039564_, _039565_, _039566_, _039567_, _039568_, _039569_, _039570_, _039571_, _039572_, _039573_, _039574_, _039575_, _039576_, _039577_, _039578_, _039579_, _039580_, _039581_, _039582_, _039583_, _039584_, _039585_, _039586_, _039587_, _039588_, _039589_, _039590_, _039591_, _039592_, _039593_, _039594_, _039595_, _039596_, _039597_, _039598_, _039599_, _039600_, _039601_, _039602_, _039603_, _039604_, _039605_, _039606_, _039607_, _039608_, _039609_, _039610_, _039611_, _039612_, _039613_, _039614_, _039615_, _039616_, _039617_, _039618_, _039619_, _039620_, _039621_, _039622_, _039623_, _039624_, _039625_, _039626_, _039627_, _039628_, _039629_, _039630_, _039631_, _039632_, _039633_, _039634_, _039635_, _039636_, _039637_, _039638_, _039639_, _039640_, _039641_, _039642_, _039643_, _039644_, _039645_, _039646_, _039647_, _039648_, _039649_, _039650_, _039651_, _039652_, _039653_, _039654_, _039655_, _039656_, _039657_, _039658_, _039659_, _039660_, _039661_, _039662_, _039663_, _039664_, _039665_, _039666_, _039667_, _039668_, _039669_, _039670_, _039671_, _039672_, _039673_, _039674_, _039675_, _039676_, _039677_, _039678_, _039679_, _039680_, _039681_, _039682_, _039683_, _039684_, _039685_, _039686_, _039687_, _039688_, _039689_, _039690_, _039691_, _039692_, _039693_, _039694_, _039695_, _039696_, _039697_, _039698_, _039699_, _039700_, _039701_, _039702_, _039703_, _039704_, _039705_, _039706_, _039707_, _039708_, _039709_, _039710_, _039711_, _039712_, _039713_, _039714_, _039715_, _039716_, _039717_, _039718_, _039719_, _039720_, _039721_, _039722_, _039723_, _039724_, _039725_, _039726_, _039727_, _039728_, _039729_, _039730_, _039731_, _039732_, _039733_, _039734_, _039735_, _039736_, _039737_, _039738_, _039739_, _039740_, _039741_, _039742_, _039743_, _039744_, _039745_, _039746_, _039747_, _039748_, _039749_, _039750_, _039751_, _039752_, _039753_, _039754_, _039755_, _039756_, _039757_, _039758_, _039759_, _039760_, _039761_, _039762_, _039763_, _039764_, _039765_, _039766_, _039767_, _039768_, _039769_, _039770_, _039771_, _039772_, _039773_, _039774_, _039775_, _039776_, _039777_, _039778_, _039779_, _039780_, _039781_, _039782_, _039783_, _039784_, _039785_, _039786_, _039787_, _039788_, _039789_, _039790_, _039791_, _039792_, _039793_, _039794_, _039795_, _039796_, _039797_, _039798_, _039799_, _039800_, _039801_, _039802_, _039803_, _039804_, _039805_, _039806_, _039807_, _039808_, _039809_, _039810_, _039811_, _039812_, _039813_, _039814_, _039815_, _039816_, _039817_, _039818_, _039819_, _039820_, _039821_, _039822_, _039823_, _039824_, _039825_, _039826_, _039827_, _039828_, _039829_, _039830_, _039831_, _039832_, _039833_, _039834_, _039835_, _039836_, _039837_, _039838_, _039839_, _039840_, _039841_, _039842_, _039843_, _039844_, _039845_, _039846_, _039847_, _039848_, _039849_, _039850_, _039851_, _039852_, _039853_, _039854_, _039855_, _039856_, _039857_, _039858_, _039859_, _039860_, _039861_, _039862_, _039863_, _039864_, _039865_, _039866_, _039867_, _039868_, _039869_, _039870_, _039871_, _039872_, _039873_, _039874_, _039875_, _039876_, _039877_, _039878_, _039879_, _039880_, _039881_, _039882_, _039883_, _039884_, _039885_, _039886_, _039887_, _039888_, _039889_, _039890_, _039891_, _039892_, _039893_, _039894_, _039895_, _039896_, _039897_, _039898_, _039899_, _039900_, _039901_, _039902_, _039903_, _039904_, _039905_, _039906_, _039907_, _039908_, _039909_, _039910_, _039911_, _039912_, _039913_, _039914_, _039915_, _039916_, _039917_, _039918_, _039919_, _039920_, _039921_, _039922_, _039923_, _039924_, _039925_, _039926_, _039927_, _039928_, _039929_, _039930_, _039931_, _039932_, _039933_, _039934_, _039935_, _039936_, _039937_, _039938_, _039939_, _039940_, _039941_, _039942_, _039943_, _039944_, _039945_, _039946_, _039947_, _039948_, _039949_, _039950_, _039951_, _039952_, _039953_, _039954_, _039955_, _039956_, _039957_, _039958_, _039959_, _039960_, _039961_, _039962_, _039963_, _039964_, _039965_, _039966_, _039967_, _039968_, _039969_, _039970_, _039971_, _039972_, _039973_, _039974_, _039975_, _039976_, _039977_, _039978_, _039979_, _039980_, _039981_, _039982_, _039983_, _039984_, _039985_, _039986_, _039987_, _039988_, _039989_, _039990_, _039991_, _039992_, _039993_, _039994_, _039995_, _039996_, _039997_, _039998_, _039999_, _040000_, _040001_, _040002_, _040003_, _040004_, _040005_, _040006_, _040007_, _040008_, _040009_, _040010_, _040011_, _040012_, _040013_, _040014_, _040015_, _040016_, _040017_, _040018_, _040019_, _040020_, _040021_, _040022_, _040023_, _040024_, _040025_, _040026_, _040027_, _040028_, _040029_, _040030_, _040031_, _040032_, _040033_, _040034_, _040035_, _040036_, _040037_, _040038_, _040039_, _040040_, _040041_, _040042_, _040043_, _040044_, _040045_, _040046_, _040047_, _040048_, _040049_, _040050_, _040051_, _040052_, _040053_, _040054_, _040055_, _040056_, _040057_, _040058_, _040059_, _040060_, _040061_, _040062_, _040063_, _040064_, _040065_, _040066_, _040067_, _040068_, _040069_, _040070_, _040071_, _040072_, _040073_, _040074_, _040075_, _040076_, _040077_, _040078_, _040079_, _040080_, _040081_, _040082_, _040083_, _040084_, _040085_, _040086_, _040087_, _040088_, _040089_, _040090_, _040091_, _040092_, _040093_, _040094_, _040095_, _040096_, _040097_, _040098_, _040099_, _040100_, _040101_, _040102_, _040103_, _040104_, _040105_, _040106_, _040107_, _040108_, _040109_, _040110_, _040111_, _040112_, _040113_, _040114_, _040115_, _040116_, _040117_, _040118_, _040119_, _040120_, _040121_, _040122_, _040123_, _040124_, _040125_, _040126_, _040127_, _040128_, _040129_, _040130_, _040131_, _040132_, _040133_, _040134_, _040135_, _040136_, _040137_, _040138_, _040139_, _040140_, _040141_, _040142_, _040143_, _040144_, _040145_, _040146_, _040147_, _040148_, _040149_, _040150_, _040151_, _040152_, _040153_, _040154_, _040155_, _040156_, _040157_, _040158_, _040159_, _040160_, _040161_, _040162_, _040163_, _040164_, _040165_, _040166_, _040167_, _040168_, _040169_, _040170_, _040171_, _040172_, _040173_, _040174_, _040175_, _040176_, _040177_, _040178_, _040179_, _040180_, _040181_, _040182_, _040183_, _040184_, _040185_, _040186_, _040187_, _040188_, _040189_, _040190_, _040191_, _040192_, _040193_, _040194_, _040195_, _040196_, _040197_, _040198_, _040199_, _040200_, _040201_, _040202_, _040203_, _040204_, _040205_, _040206_, _040207_, _040208_, _040209_, _040210_, _040211_, _040212_, _040213_, _040214_, _040215_, _040216_, _040217_, _040218_, _040219_, _040220_, _040221_, _040222_, _040223_, _040224_, _040225_, _040226_, _040227_, _040228_, _040229_, _040230_, _040231_, _040232_, _040233_, _040234_, _040235_, _040236_, _040237_, _040238_, _040239_, _040240_, _040241_, _040242_, _040243_, _040244_, _040245_, _040246_, _040247_, _040248_, _040249_, _040250_, _040251_, _040252_, _040253_, _040254_, _040255_, _040256_, _040257_, _040258_, _040259_, _040260_, _040261_, _040262_, _040263_, _040264_, _040265_, _040266_, _040267_, _040268_, _040269_, _040270_, _040271_, _040272_, _040273_, _040274_, _040275_, _040276_, _040277_, _040278_, _040279_, _040280_, _040281_, _040282_, _040283_, _040284_, _040285_, _040286_, _040287_, _040288_, _040289_, _040290_, _040291_, _040292_, _040293_, _040294_, _040295_, _040296_, _040297_, _040298_, _040299_, _040300_, _040301_, _040302_, _040303_, _040304_, _040305_, _040306_, _040307_, _040308_, _040309_, _040310_, _040311_, _040312_, _040313_, _040314_, _040315_, _040316_, _040317_, _040318_, _040319_, _040320_, _040321_, _040322_, _040323_, _040324_, _040325_, _040326_, _040327_, _040328_, _040329_, _040330_, _040331_, _040332_, _040333_, _040334_, _040335_, _040336_, _040337_, _040338_, _040339_, _040340_, _040341_, _040342_, _040343_, _040344_, _040345_, _040346_, _040347_, _040348_, _040349_, _040350_, _040351_, _040352_, _040353_, _040354_, _040355_, _040356_, _040357_, _040358_, _040359_, _040360_, _040361_, _040362_, _040363_, _040364_, _040365_, _040366_, _040367_, _040368_, _040369_, _040370_, _040371_, _040372_, _040373_, _040374_, _040375_, _040376_, _040377_, _040378_, _040379_, _040380_, _040381_, _040382_, _040383_, _040384_, _040385_, _040386_, _040387_, _040388_, _040389_, _040390_, _040391_, _040392_, _040393_, _040394_, _040395_, _040396_, _040397_, _040398_, _040399_, _040400_, _040401_, _040402_, _040403_, _040404_, _040405_, _040406_, _040407_, _040408_, _040409_, _040410_, _040411_, _040412_, _040413_, _040414_, _040415_, _040416_, _040417_, _040418_, _040419_, _040420_, _040421_, _040422_, _040423_, _040424_, _040425_, _040426_, _040427_, _040428_, _040429_, _040430_, _040431_, _040432_, _040433_, _040434_, _040435_, _040436_, _040437_, _040438_, _040439_, _040440_, _040441_, _040442_, _040443_, _040444_, _040445_, _040446_, _040447_, _040448_, _040449_, _040450_, _040451_, _040452_, _040453_, _040454_, _040455_, _040456_, _040457_, _040458_, _040459_, _040460_, _040461_, _040462_, _040463_, _040464_, _040465_, _040466_, _040467_, _040468_, _040469_, _040470_, _040471_, _040472_, _040473_, _040474_, _040475_, _040476_, _040477_, _040478_, _040479_, _040480_, _040481_, _040482_, _040483_, _040484_, _040485_, _040486_, _040487_, _040488_, _040489_, _040490_, _040491_, _040492_, _040493_, _040494_, _040495_, _040496_, _040497_, _040498_, _040499_, _040500_, _040501_, _040502_, _040503_, _040504_, _040505_, _040506_, _040507_, _040508_, _040509_, _040510_, _040511_, _040512_, _040513_, _040514_, _040515_, _040516_, _040517_, _040518_, _040519_, _040520_, _040521_, _040522_, _040523_, _040524_, _040525_, _040526_, _040527_, _040528_, _040529_, _040530_, _040531_, _040532_, _040533_, _040534_, _040535_, _040536_, _040537_, _040538_, _040539_, _040540_, _040541_, _040542_, _040543_, _040544_, _040545_, _040546_, _040547_, _040548_, _040549_, _040550_, _040551_, _040552_, _040553_, _040554_, _040555_, _040556_, _040557_, _040558_, _040559_, _040560_, _040561_, _040562_, _040563_, _040564_, _040565_, _040566_, _040567_, _040568_, _040569_, _040570_, _040571_, _040572_, _040573_, _040574_, _040575_, _040576_, _040577_, _040578_, _040579_, _040580_, _040581_, _040582_, _040583_, _040584_, _040585_, _040586_, _040587_, _040588_, _040589_, _040590_, _040591_, _040592_, _040593_, _040594_, _040595_, _040596_, _040597_, _040598_, _040599_, _040600_, _040601_, _040602_, _040603_, _040604_, _040605_, _040606_, _040607_, _040608_, _040609_, _040610_, _040611_, _040612_, _040613_, _040614_, _040615_, _040616_, _040617_, _040618_, _040619_, _040620_, _040621_, _040622_, _040623_, _040624_, _040625_, _040626_, _040627_, _040628_, _040629_, _040630_, _040631_, _040632_, _040633_, _040634_, _040635_, _040636_, _040637_, _040638_, _040639_, _040640_, _040641_, _040642_, _040643_, _040644_, _040645_, _040646_, _040647_, _040648_, _040649_, _040650_, _040651_, _040652_, _040653_, _040654_, _040655_, _040656_, _040657_, _040658_, _040659_, _040660_, _040661_, _040662_, _040663_, _040664_, _040665_, _040666_, _040667_, _040668_, _040669_, _040670_, _040671_, _040672_, _040673_, _040674_, _040675_, _040676_, _040677_, _040678_, _040679_, _040680_, _040681_, _040682_, _040683_, _040684_, _040685_, _040686_, _040687_, _040688_, _040689_, _040690_, _040691_, _040692_, _040693_, _040694_, _040695_, _040696_, _040697_, _040698_, _040699_, _040700_, _040701_, _040702_, _040703_, _040704_, _040705_, _040706_, _040707_, _040708_, _040709_, _040710_, _040711_, _040712_, _040713_, _040714_, _040715_, _040716_, _040717_, _040718_, _040719_, _040720_, _040721_, _040722_, _040723_, _040724_, _040725_, _040726_, _040727_, _040728_, _040729_, _040730_, _040731_, _040732_, _040733_, _040734_, _040735_, _040736_, _040737_, _040738_, _040739_, _040740_, _040741_, _040742_, _040743_, _040744_, _040745_, _040746_, _040747_, _040748_, _040749_, _040750_, _040751_, _040752_, _040753_, _040754_, _040755_, _040756_, _040757_, _040758_, _040759_, _040760_, _040761_, _040762_, _040763_, _040764_, _040765_, _040766_, _040767_, _040768_, _040769_, _040770_, _040771_, _040772_, _040773_, _040774_, _040775_, _040776_, _040777_, _040778_, _040779_, _040780_, _040781_, _040782_, _040783_, _040784_, _040785_, _040786_, _040787_, _040788_, _040789_, _040790_, _040791_, _040792_, _040793_, _040794_, _040795_, _040796_, _040797_, _040798_, _040799_, _040800_, _040801_, _040802_, _040803_, _040804_, _040805_, _040806_, _040807_, _040808_, _040809_, _040810_, _040811_, _040812_, _040813_, _040814_, _040815_, _040816_, _040817_, _040818_, _040819_, _040820_, _040821_, _040822_, _040823_, _040824_, _040825_, _040826_, _040827_, _040828_, _040829_, _040830_, _040831_, _040832_, _040833_, _040834_, _040835_, _040836_, _040837_, _040838_, _040839_, _040840_, _040841_, _040842_, _040843_, _040844_, _040845_, _040846_, _040847_, _040848_, _040849_, _040850_, _040851_, _040852_, _040853_, _040854_, _040855_, _040856_, _040857_, _040858_, _040859_, _040860_, _040861_, _040862_, _040863_, _040864_, _040865_, _040866_, _040867_, _040868_, _040869_, _040870_, _040871_, _040872_, _040873_, _040874_, _040875_, _040876_, _040877_, _040878_, _040879_, _040880_, _040881_, _040882_, _040883_, _040884_, _040885_, _040886_, _040887_, _040888_, _040889_, _040890_, _040891_, _040892_, _040893_, _040894_, _040895_, _040896_, _040897_, _040898_, _040899_, _040900_, _040901_, _040902_, _040903_, _040904_, _040905_, _040906_, _040907_, _040908_, _040909_, _040910_, _040911_, _040912_, _040913_, _040914_, _040915_, _040916_, _040917_, _040918_, _040919_, _040920_, _040921_, _040922_, _040923_, _040924_, _040925_, _040926_, _040927_, _040928_, _040929_, _040930_, _040931_, _040932_, _040933_, _040934_, _040935_, _040936_, _040937_, _040938_, _040939_, _040940_, _040941_, _040942_, _040943_, _040944_, _040945_, _040946_, _040947_, _040948_, _040949_, _040950_, _040951_, _040952_, _040953_, _040954_, _040955_, _040956_, _040957_, _040958_, _040959_, _040960_, _040961_, _040962_, _040963_, _040964_, _040965_, _040966_, _040967_, _040968_, _040969_, _040970_, _040971_, _040972_, _040973_, _040974_, _040975_, _040976_, _040977_, _040978_, _040979_, _040980_, _040981_, _040982_, _040983_, _040984_, _040985_, _040986_, _040987_, _040988_, _040989_, _040990_, _040991_, _040992_, _040993_, _040994_, _040995_, _040996_, _040997_, _040998_, _040999_, _041000_, _041001_, _041002_, _041003_, _041004_, _041005_, _041006_, _041007_, _041008_, _041009_, _041010_, _041011_, _041012_, _041013_, _041014_, _041015_, _041016_, _041017_, _041018_, _041019_, _041020_, _041021_, _041022_, _041023_, _041024_, _041025_, _041026_, _041027_, _041028_, _041029_, _041030_, _041031_, _041032_, _041033_, _041034_, _041035_, _041036_, _041037_, _041038_, _041039_, _041040_, _041041_, _041042_, _041043_, _041044_, _041045_, _041046_, _041047_, _041048_, _041049_, _041050_, _041051_, _041052_, _041053_, _041054_, _041055_, _041056_, _041057_, _041058_, _041059_, _041060_, _041061_, _041062_, _041063_, _041064_, _041065_, _041066_, _041067_, _041068_, _041069_, _041070_, _041071_, _041072_, _041073_, _041074_, _041075_, _041076_, _041077_, _041078_, _041079_, _041080_, _041081_, _041082_, _041083_, _041084_, _041085_, _041086_, _041087_, _041088_, _041089_, _041090_, _041091_, _041092_, _041093_, _041094_, _041095_, _041096_, _041097_, _041098_, _041099_, _041100_, _041101_, _041102_, _041103_, _041104_, _041105_, _041106_, _041107_, _041108_, _041109_, _041110_, _041111_, _041112_, _041113_, _041114_, _041115_, _041116_, _041117_, _041118_, _041119_, _041120_, _041121_, _041122_, _041123_, _041124_, _041125_, _041126_, _041127_, _041128_, _041129_, _041130_, _041131_, _041132_, _041133_, _041134_, _041135_, _041136_, _041137_, _041138_, _041139_, _041140_, _041141_, _041142_, _041143_, _041144_, _041145_, _041146_, _041147_, _041148_, _041149_, _041150_, _041151_, _041152_, _041153_, _041154_, _041155_, _041156_, _041157_, _041158_, _041159_, _041160_, _041161_, _041162_, _041163_, _041164_, _041165_, _041166_, _041167_, _041168_, _041169_, _041170_, _041171_, _041172_, _041173_, _041174_, _041175_, _041176_, _041177_, _041178_, _041179_, _041180_, _041181_, _041182_, _041183_, _041184_, _041185_, _041186_, _041187_, _041188_, _041189_, _041190_, _041191_, _041192_, _041193_, _041194_, _041195_, _041196_, _041197_, _041198_, _041199_, _041200_, _041201_, _041202_, _041203_, _041204_, _041205_, _041206_, _041207_, _041208_, _041209_, _041210_, _041211_, _041212_, _041213_, _041214_, _041215_, _041216_, _041217_, _041218_, _041219_, _041220_, _041221_, _041222_, _041223_, _041224_, _041225_, _041226_, _041227_, _041228_, _041229_, _041230_, _041231_, _041232_, _041233_, _041234_, _041235_, _041236_, _041237_, _041238_, _041239_, _041240_, _041241_, _041242_, _041243_, _041244_, _041245_, _041246_, _041247_, _041248_, _041249_, _041250_, _041251_, _041252_, _041253_, _041254_, _041255_, _041256_, _041257_, _041258_, _041259_, _041260_, _041261_, _041262_, _041263_, _041264_, _041265_, _041266_, _041267_, _041268_, _041269_, _041270_, _041271_, _041272_, _041273_, _041274_, _041275_, _041276_, _041277_, _041278_, _041279_, _041280_, _041281_, _041282_, _041283_, _041284_, _041285_, _041286_, _041287_, _041288_, _041289_, _041290_, _041291_, _041292_, _041293_, _041294_, _041295_, _041296_, _041297_, _041298_, _041299_, _041300_, _041301_, _041302_, _041303_, _041304_, _041305_, _041306_, _041307_, _041308_, _041309_, _041310_, _041311_, _041312_, _041313_, _041314_, _041315_, _041316_, _041317_, _041318_, _041319_, _041320_, _041321_, _041322_, _041323_, _041324_, _041325_, _041326_, _041327_, _041328_, _041329_, _041330_, _041331_, _041332_, _041333_, _041334_, _041335_, _041336_, _041337_, _041338_, _041339_, _041340_, _041341_, _041342_, _041343_, _041344_, _041345_, _041346_, _041347_, _041348_, _041349_, _041350_, _041351_, _041352_, _041353_, _041354_, _041355_, _041356_, _041357_, _041358_, _041359_, _041360_, _041361_, _041362_, _041363_, _041364_, _041365_, _041366_, _041367_, _041368_, _041369_, _041370_, _041371_, _041372_, _041373_, _041374_, _041375_, _041376_, _041377_, _041378_, _041379_, _041380_, _041381_, _041382_, _041383_, _041384_, _041385_, _041386_, _041387_, _041388_, _041389_, _041390_, _041391_, _041392_, _041393_, _041394_, _041395_, _041396_, _041397_, _041398_, _041399_, _041400_, _041401_, _041402_, _041403_, _041404_, _041405_, _041406_, _041407_, _041408_, _041409_, _041410_, _041411_, _041412_, _041413_, _041414_, _041415_, _041416_, _041417_, _041418_, _041419_, _041420_, _041421_, _041422_, _041423_, _041424_, _041425_, _041426_, _041427_, _041428_, _041429_, _041430_, _041431_, _041432_, _041433_, _041434_, _041435_, _041436_, _041437_, _041438_, _041439_, _041440_, _041441_, _041442_, _041443_, _041444_, _041445_, _041446_, _041447_, _041448_, _041449_, _041450_, _041451_, _041452_, _041453_, _041454_, _041455_, _041456_, _041457_, _041458_, _041459_, _041460_, _041461_, _041462_, _041463_, _041464_, _041465_, _041466_, _041467_, _041468_, _041469_, _041470_, _041471_, _041472_, _041473_, _041474_, _041475_, _041476_, _041477_, _041478_, _041479_, _041480_, _041481_, _041482_, _041483_, _041484_, _041485_, _041486_, _041487_, _041488_, _041489_, _041490_, _041491_, _041492_, _041493_, _041494_, _041495_, _041496_, _041497_, _041498_, _041499_, _041500_, _041501_, _041502_, _041503_, _041504_, _041505_, _041506_, _041507_, _041508_, _041509_, _041510_, _041511_, _041512_, _041513_, _041514_, _041515_, _041516_, _041517_, _041518_, _041519_, _041520_, _041521_, _041522_, _041523_, _041524_, _041525_, _041526_, _041527_, _041528_, _041529_, _041530_, _041531_, _041532_, _041533_, _041534_, _041535_, _041536_, _041537_, _041538_, _041539_, _041540_, _041541_, _041542_, _041543_, _041544_, _041545_, _041546_, _041547_, _041548_, _041549_, _041550_, _041551_, _041552_, _041553_, _041554_, _041555_, _041556_, _041557_, _041558_, _041559_, _041560_, _041561_, _041562_, _041563_, _041564_, _041565_, _041566_, _041567_, _041568_, _041569_, _041570_, _041571_, _041572_, _041573_, _041574_, _041575_, _041576_, _041577_, _041578_, _041579_, _041580_, _041581_, _041582_, _041583_, _041584_, _041585_, _041586_, _041587_, _041588_, _041589_, _041590_, _041591_, _041592_, _041593_, _041594_, _041595_, _041596_, _041597_, _041598_, _041599_, _041600_, _041601_, _041602_, _041603_, _041604_, _041605_, _041606_, _041607_, _041608_, _041609_, _041610_, _041611_, _041612_, _041613_, _041614_, _041615_, _041616_, _041617_, _041618_, _041619_, _041620_, _041621_, _041622_, _041623_, _041624_, _041625_, _041626_, _041627_, _041628_, _041629_, _041630_, _041631_, _041632_, _041633_, _041634_, _041635_, _041636_, _041637_, _041638_, _041639_, _041640_, _041641_, _041642_, _041643_, _041644_, _041645_, _041646_, _041647_, _041648_, _041649_, _041650_, _041651_, _041652_, _041653_, _041654_, _041655_, _041656_, _041657_, _041658_, _041659_, _041660_, _041661_, _041662_, _041663_, _041664_, _041665_, _041666_, _041667_, _041668_, _041669_, _041670_, _041671_, _041672_, _041673_, _041674_, _041675_, _041676_, _041677_, _041678_, _041679_, _041680_, _041681_, _041682_, _041683_, _041684_, _041685_, _041686_, _041687_, _041688_, _041689_, _041690_, _041691_, _041692_, _041693_, _041694_, _041695_, _041696_, _041697_, _041698_, _041699_, _041700_, _041701_, _041702_, _041703_, _041704_, _041705_, _041706_, _041707_, _041708_, _041709_, _041710_, _041711_, _041712_, _041713_, _041714_, _041715_, _041716_, _041717_, _041718_, _041719_, _041720_, _041721_, _041722_, _041723_, _041724_, _041725_, _041726_, _041727_, _041728_, _041729_, _041730_, _041731_, _041732_, _041733_, _041734_, _041735_, _041736_, _041737_, _041738_, _041739_, _041740_, _041741_, _041742_, _041743_, _041744_, _041745_, _041746_, _041747_, _041748_, _041749_, _041750_, _041751_, _041752_, _041753_, _041754_, _041755_, _041756_, _041757_, _041758_, _041759_, _041760_, _041761_, _041762_, _041763_, _041764_, _041765_, _041766_, _041767_, _041768_, _041769_, _041770_, _041771_, _041772_, _041773_, _041774_, _041775_, _041776_, _041777_, _041778_, _041779_, _041780_, _041781_, _041782_, _041783_, _041784_, _041785_, _041786_, _041787_, _041788_, _041789_, _041790_, _041791_, _041792_, _041793_, _041794_, _041795_, _041796_, _041797_, _041798_, _041799_, _041800_, _041801_, _041802_, _041803_, _041804_, _041805_, _041806_, _041807_, _041808_, _041809_, _041810_, _041811_, _041812_, _041813_, _041814_, _041815_, _041816_, _041817_, _041818_, _041819_, _041820_, _041821_, _041822_, _041823_, _041824_, _041825_, _041826_, _041827_, _041828_, _041829_, _041830_, _041831_, _041832_, _041833_, _041834_, _041835_, _041836_, _041837_, _041838_, _041839_, _041840_, _041841_, _041842_, _041843_, _041844_, _041845_, _041846_, _041847_, _041848_, _041849_, _041850_, _041851_, _041852_, _041853_, _041854_, _041855_, _041856_, _041857_, _041858_, _041859_, _041860_, _041861_, _041862_, _041863_, _041864_, _041865_, _041866_, _041867_, _041868_, _041869_, _041870_, _041871_, _041872_, _041873_, _041874_, _041875_, _041876_, _041877_, _041878_, _041879_, _041880_, _041881_, _041882_, _041883_, _041884_, _041885_, _041886_, _041887_, _041888_, _041889_, _041890_, _041891_, _041892_, _041893_, _041894_, _041895_, _041896_, _041897_, _041898_, _041899_, _041900_, _041901_, _041902_, _041903_, _041904_, _041905_, _041906_, _041907_, _041908_, _041909_, _041910_, _041911_, _041912_, _041913_, _041914_, _041915_, _041916_, _041917_, _041918_, _041919_, _041920_, _041921_, _041922_, _041923_, _041924_, _041925_, _041926_, _041927_, _041928_, _041929_, _041930_, _041931_, _041932_, _041933_, _041934_, _041935_, _041936_, _041937_, _041938_, _041939_, _041940_, _041941_, _041942_, _041943_, _041944_, _041945_, _041946_, _041947_, _041948_, _041949_, _041950_, _041951_, _041952_, _041953_, _041954_, _041955_, _041956_, _041957_, _041958_, _041959_, _041960_, _041961_, _041962_, _041963_, _041964_, _041965_, _041966_, _041967_, _041968_, _041969_, _041970_, _041971_, _041972_, _041973_, _041974_, _041975_, _041976_, _041977_, _041978_, _041979_, _041980_, _041981_, _041982_, _041983_, _041984_, _041985_, _041986_, _041987_, _041988_, _041989_, _041990_, _041991_, _041992_, _041993_, _041994_, _041995_, _041996_, _041997_, _041998_, _041999_, _042000_, _042001_, _042002_, _042003_, _042004_, _042005_, _042006_, _042007_, _042008_, _042009_, _042010_, _042011_, _042012_, _042013_, _042014_, _042015_, _042016_, _042017_, _042018_, _042019_, _042020_, _042021_, _042022_, _042023_, _042024_, _042025_, _042026_, _042027_, _042028_, _042029_, _042030_, _042031_, _042032_, _042033_, _042034_, _042035_, _042036_, _042037_, _042038_, _042039_, _042040_, _042041_, _042042_, _042043_, _042044_, _042045_, _042046_, _042047_, _042048_, _042049_, _042050_, _042051_, _042052_, _042053_, _042054_, _042055_, _042056_, _042057_, _042058_, _042059_, _042060_, _042061_, _042062_, _042063_, _042064_, _042065_, _042066_, _042067_, _042068_, _042069_, _042070_, _042071_, _042072_, _042073_, _042074_, _042075_, _042076_, _042077_, _042078_, _042079_, _042080_, _042081_, _042082_, _042083_, _042084_, _042085_, _042086_, _042087_, _042088_, _042089_, _042090_, _042091_, _042092_, _042093_, _042094_, _042095_, _042096_, _042097_, _042098_, _042099_, _042100_, _042101_, _042102_, _042103_, _042104_, _042105_, _042106_, _042107_, _042108_, _042109_, _042110_, _042111_, _042112_, _042113_, _042114_, _042115_, _042116_, _042117_, _042118_, _042119_, _042120_, _042121_, _042122_, _042123_, _042124_, _042125_, _042126_, _042127_, _042128_, _042129_, _042130_, _042131_, _042132_, _042133_, _042134_, _042135_, _042136_, _042137_, _042138_, _042139_, _042140_, _042141_, _042142_, _042143_, _042144_, _042145_, _042146_, _042147_, _042148_, _042149_, _042150_, _042151_, _042152_, _042153_, _042154_, _042155_, _042156_, _042157_, _042158_, _042159_, _042160_, _042161_, _042162_, _042163_, _042164_, _042165_, _042166_, _042167_, _042168_, _042169_, _042170_, _042171_, _042172_, _042173_, _042174_, _042175_, _042176_, _042177_, _042178_, _042179_, _042180_, _042181_, _042182_, _042183_, _042184_, _042185_, _042186_, _042187_, _042188_, _042189_, _042190_, _042191_, _042192_, _042193_, _042194_, _042195_, _042196_, _042197_, _042198_, _042199_, _042200_, _042201_, _042202_, _042203_, _042204_, _042205_, _042206_, _042207_, _042208_, _042209_, _042210_, _042211_, _042212_, _042213_, _042214_, _042215_, _042216_, _042217_, _042218_, _042219_, _042220_, _042221_, _042222_, _042223_, _042224_, _042225_, _042226_, _042227_, _042228_, _042229_, _042230_, _042231_, _042232_, _042233_, _042234_, _042235_, _042236_, _042237_, _042238_, _042239_, _042240_, _042241_, _042242_, _042243_, _042244_, _042245_, _042246_, _042247_, _042248_, _042249_, _042250_, _042251_, _042252_, _042253_, _042254_, _042255_, _042256_, _042257_, _042258_, _042259_, _042260_, _042261_, _042262_, _042263_, _042264_, _042265_, _042266_, _042267_, _042268_, _042269_, _042270_, _042271_, _042272_, _042273_, _042274_, _042275_, _042276_, _042277_, _042278_, _042279_, _042280_, _042281_, _042282_, _042283_, _042284_, _042285_, _042286_, _042287_, _042288_, _042289_, _042290_, _042291_, _042292_, _042293_, _042294_, _042295_, _042296_, _042297_, _042298_, _042299_, _042300_, _042301_, _042302_, _042303_, _042304_, _042305_, _042306_, _042307_, _042308_, _042309_, _042310_, _042311_, _042312_, _042313_, _042314_, _042315_, _042316_, _042317_, _042318_, _042319_, _042320_, _042321_, _042322_, _042323_, _042324_, _042325_, _042326_, _042327_, _042328_, _042329_, _042330_, _042331_, _042332_, _042333_, _042334_, _042335_, _042336_, _042337_, _042338_, _042339_, _042340_, _042341_, _042342_, _042343_, _042344_, _042345_, _042346_, _042347_, _042348_, _042349_, _042350_, _042351_, _042352_, _042353_, _042354_, _042355_, _042356_, _042357_, _042358_, _042359_, _042360_, _042361_, _042362_, _042363_, _042364_, _042365_, _042366_, _042367_, _042368_, _042369_, _042370_, _042371_, _042372_, _042373_, _042374_, _042375_, _042376_, _042377_, _042378_, _042379_, _042380_, _042381_, _042382_, _042383_, _042384_, _042385_, _042386_, _042387_, _042388_, _042389_, _042390_, _042391_, _042392_, _042393_, _042394_, _042395_, _042396_, _042397_, _042398_, _042399_, _042400_, _042401_, _042402_, _042403_, _042404_, _042405_, _042406_, _042407_, _042408_, _042409_, _042410_, _042411_, _042412_, _042413_, _042414_, _042415_, _042416_, _042417_, _042418_, _042419_, _042420_, _042421_, _042422_, _042423_, _042424_, _042425_, _042426_, _042427_, _042428_, _042429_, _042430_, _042431_, _042432_, _042433_, _042434_, _042435_, _042436_, _042437_, _042438_, _042439_, _042440_, _042441_, _042442_, _042443_, _042444_, _042445_, _042446_, _042447_, _042448_, _042449_, _042450_, _042451_, _042452_, _042453_, _042454_, _042455_, _042456_, _042457_, _042458_, _042459_, _042460_, _042461_, _042462_, _042463_, _042464_, _042465_, _042466_, _042467_, _042468_, _042469_, _042470_, _042471_, _042472_, _042473_, _042474_, _042475_, _042476_, _042477_, _042478_, _042479_, _042480_, _042481_, _042482_, _042483_, _042484_, _042485_, _042486_, _042487_, _042488_, _042489_, _042490_, _042491_, _042492_, _042493_, _042494_, _042495_, _042496_, _042497_, _042498_, _042499_, _042500_, _042501_, _042502_, _042503_, _042504_, _042505_, _042506_, _042507_, _042508_, _042509_, _042510_, _042511_, _042512_, _042513_, _042514_, _042515_, _042516_, _042517_, _042518_, _042519_, _042520_, _042521_, _042522_, _042523_, _042524_, _042525_, _042526_, _042527_, _042528_, _042529_, _042530_, _042531_, _042532_, _042533_, _042534_, _042535_, _042536_, _042537_, _042538_, _042539_, _042540_, _042541_, _042542_, _042543_, _042544_, _042545_, _042546_, _042547_, _042548_, _042549_, _042550_, _042551_, _042552_, _042553_, _042554_, _042555_, _042556_, _042557_, _042558_, _042559_, _042560_, _042561_, _042562_, _042563_, _042564_, _042565_, _042566_, _042567_, _042568_, _042569_, _042570_, _042571_, _042572_, _042573_, _042574_, _042575_, _042576_, _042577_, _042578_, _042579_, _042580_, _042581_, _042582_, _042583_, _042584_, _042585_, _042586_, _042587_, _042588_, _042589_, _042590_, _042591_, _042592_, _042593_, _042594_, _042595_, _042596_, _042597_, _042598_, _042599_, _042600_, _042601_, _042602_, _042603_, _042604_, _042605_, _042606_, _042607_, _042608_, _042609_, _042610_, _042611_, _042612_, _042613_, _042614_, _042615_, _042616_, _042617_, _042618_, _042619_, _042620_, _042621_, _042622_, _042623_, _042624_, _042625_, _042626_, _042627_, _042628_, _042629_, _042630_, _042631_, _042632_, _042633_, _042634_, _042635_, _042636_, _042637_, _042638_, _042639_, _042640_, _042641_, _042642_, _042643_, _042644_, _042645_, _042646_, _042647_, _042648_, _042649_, _042650_, _042651_, _042652_, _042653_, _042654_, _042655_, _042656_, _042657_, _042658_, _042659_, _042660_, _042661_, _042662_, _042663_, _042664_, _042665_, _042666_, _042667_, _042668_, _042669_, _042670_, _042671_, _042672_, _042673_, _042674_, _042675_, _042676_, _042677_, _042678_, _042679_, _042680_, _042681_, _042682_, _042683_, _042684_, _042685_, _042686_, _042687_, _042688_, _042689_, _042690_, _042691_, _042692_, _042693_, _042694_, _042695_, _042696_, _042697_, _042698_, _042699_, _042700_, _042701_, _042702_, _042703_, _042704_, _042705_, _042706_, _042707_, _042708_, _042709_, _042710_, _042711_, _042712_, _042713_, _042714_, _042715_, _042716_, _042717_, _042718_, _042719_, _042720_, _042721_, _042722_, _042723_, _042724_, _042725_, _042726_, _042727_, _042728_, _042729_, _042730_, _042731_, _042732_, _042733_, _042734_, _042735_, _042736_, _042737_, _042738_, _042739_, _042740_, _042741_, _042742_, _042743_, _042744_, _042745_, _042746_, _042747_, _042748_, _042749_, _042750_, _042751_, _042752_, _042753_, _042754_, _042755_, _042756_, _042757_, _042758_, _042759_, _042760_, _042761_, _042762_, _042763_, _042764_, _042765_, _042766_, _042767_, _042768_, _042769_, _042770_, _042771_, _042772_, _042773_, _042774_, _042775_, _042776_, _042777_, _042778_, _042779_, _042780_, _042781_, _042782_, _042783_, _042784_, _042785_, _042786_, _042787_, _042788_, _042789_, _042790_, _042791_, _042792_, _042793_, _042794_, _042795_, _042796_, _042797_, _042798_, _042799_, _042800_, _042801_, _042802_, _042803_, _042804_, _042805_, _042806_, _042807_, _042808_, _042809_, _042810_, _042811_, _042812_, _042813_, _042814_, _042815_, _042816_, _042817_, _042818_, _042819_, _042820_, _042821_, _042822_, _042823_, _042824_, _042825_, _042826_, _042827_, _042828_, _042829_, _042830_, _042831_, _042832_, _042833_, _042834_, _042835_, _042836_, _042837_, _042838_, _042839_, _042840_, _042841_, _042842_, _042843_, _042844_, _042845_, _042846_, _042847_, _042848_, _042849_, _042850_, _042851_, _042852_, _042853_, _042854_, _042855_, _042856_, _042857_, _042858_, _042859_, _042860_, _042861_, _042862_, _042863_, _042864_, _042865_, _042866_, _042867_, _042868_, _042869_, _042870_, _042871_, _042872_, _042873_, _042874_, _042875_, _042876_, _042877_, _042878_, _042879_, _042880_, _042881_, _042882_, _042883_, _042884_, _042885_, _042886_, _042887_, _042888_, _042889_, _042890_, _042891_, _042892_, _042893_, _042894_, _042895_, _042896_, _042897_, _042898_, _042899_, _042900_, _042901_, _042902_, _042903_, _042904_, _042905_, _042906_, _042907_, _042908_, _042909_, _042910_, _042911_, _042912_, _042913_, _042914_, _042915_, _042916_, _042917_, _042918_, _042919_, _042920_, _042921_, _042922_, _042923_, _042924_, _042925_, _042926_, _042927_, _042928_, _042929_, _042930_, _042931_, _042932_, _042933_, _042934_, _042935_, _042936_, _042937_, _042938_, _042939_, _042940_, _042941_, _042942_, _042943_, _042944_, _042945_, _042946_, _042947_, _042948_, _042949_, _042950_, _042951_, _042952_, _042953_, _042954_, _042955_, _042956_, _042957_, _042958_, _042959_, _042960_, _042961_, _042962_, _042963_, _042964_, _042965_, _042966_, _042967_, _042968_, _042969_, _042970_, _042971_, _042972_, _042973_, _042974_, _042975_, _042976_, _042977_, _042978_, _042979_, _042980_, _042981_, _042982_, _042983_, _042984_, _042985_, _042986_, _042987_, _042988_, _042989_, _042990_, _042991_, _042992_, _042993_, _042994_, _042995_, _042996_, _042997_, _042998_, _042999_, _043000_, _043001_, _043002_, _043003_, _043004_, _043005_, _043006_, _043007_, _043008_, _043009_, _043010_, _043011_, _043012_, _043013_, _043014_, _043015_, _043016_, _043017_, _043018_, _043019_, _043020_, _043021_, _043022_, _043023_, _043024_, _043025_, _043026_, _043027_, _043028_, _043029_, _043030_, _043031_, _043032_, _043033_, _043034_, _043035_, _043036_, _043037_, _043038_, _043039_, _043040_, _043041_, _043042_, _043043_, _043044_, _043045_, _043046_, _043047_, _043048_, _043049_, _043050_, _043051_, _043052_, _043053_, _043054_, _043055_, _043056_, _043057_, _043058_, _043059_, _043060_, _043061_, _043062_, _043063_, _043064_, _043065_, _043066_, _043067_, _043068_, _043069_, _043070_, _043071_, _043072_, _043073_, _043074_, _043075_, _043076_, _043077_, _043078_, _043079_, _043080_, _043081_, _043082_, _043083_, _043084_, _043085_, _043086_, _043087_, _043088_, _043089_, _043090_, _043091_, _043092_, _043093_, _043094_, _043095_, _043096_, _043097_, _043098_, _043099_, _043100_, _043101_, _043102_, _043103_, _043104_, _043105_, _043106_, _043107_, _043108_, _043109_, _043110_, _043111_, _043112_, _043113_, _043114_, _043115_, _043116_, _043117_, _043118_, _043119_, _043120_, _043121_, _043122_, _043123_, _043124_, _043125_, _043126_, _043127_, _043128_, _043129_, _043130_, _043131_, _043132_, _043133_, _043134_, _043135_, _043136_, _043137_, _043138_, _043139_, _043140_, _043141_, _043142_, _043143_, _043144_, _043145_, _043146_, _043147_, _043148_, _043149_, _043150_, _043151_, _043152_, _043153_, _043154_, _043155_, _043156_, _043157_, _043158_, _043159_, _043160_, _043161_, _043162_, _043163_, _043164_, _043165_, _043166_, _043167_, _043168_, _043169_, _043170_, _043171_, _043172_, _043173_, _043174_, _043175_, _043176_, _043177_, _043178_, _043179_, _043180_, _043181_, _043182_, _043183_, _043184_, _043185_, _043186_, _043187_, _043188_, _043189_, _043190_, _043191_, _043192_, _043193_, _043194_, _043195_, _043196_, _043197_, _043198_, _043199_, _043200_, _043201_, _043202_, _043203_, _043204_, _043205_, _043206_, _043207_, _043208_, _043209_, _043210_, _043211_, _043212_, _043213_, _043214_, _043215_, _043216_, _043217_, _043218_, _043219_, _043220_, _043221_, _043222_, _043223_, _043224_, _043225_, _043226_, _043227_, _043228_, _043229_, _043230_, _043231_, _043232_, _043233_, _043234_, _043235_, _043236_, _043237_, _043238_, _043239_, _043240_, _043241_, _043242_, _043243_, _043244_, _043245_, _043246_, _043247_, _043248_, _043249_, _043250_, _043251_, _043252_, _043253_, _043254_, _043255_, _043256_, _043257_, _043258_, _043259_, _043260_, _043261_, _043262_, _043263_, _043264_, _043265_, _043266_, _043267_, _043268_, _043269_, _043270_, _043271_, _043272_, _043273_, _043274_, _043275_, _043276_, _043277_, _043278_, _043279_, _043280_, _043281_, _043282_, _043283_, _043284_, _043285_, _043286_, _043287_, _043288_, _043289_, _043290_, _043291_, _043292_, _043293_, _043294_, _043295_, _043296_, _043297_, _043298_, _043299_, _043300_, _043301_, _043302_, _043303_, _043304_, _043305_, _043306_, _043307_, _043308_, _043309_, _043310_, _043311_, _043312_, _043313_, _043314_, _043315_, _043316_, _043317_, _043318_, _043319_, _043320_, _043321_, _043322_, _043323_, _043324_, _043325_, _043326_, _043327_, _043328_, _043329_, _043330_, _043331_, _043332_, _043333_, _043334_, _043335_, _043336_, _043337_, _043338_, _043339_, _043340_, _043341_, _043342_, _043343_, _043344_, _043345_, _043346_, _043347_, _043348_, _043349_, _043350_, _043351_, _043352_, _043353_, _043354_, _043355_, _043356_, _043357_, _043358_, _043359_, _043360_, _043361_, _043362_, _043363_, _043364_, _043365_, _043366_, _043367_, _043368_, _043369_, _043370_, _043371_, _043372_, _043373_, _043374_, _043375_, _043376_, _043377_, _043378_, _043379_, _043380_, _043381_, _043382_, _043383_, _043384_, _043385_, _043386_, _043387_, _043388_, _043389_, _043390_, _043391_, _043392_, _043393_, _043394_, _043395_, _043396_, _043397_, _043398_, _043399_, _043400_, _043401_, _043402_, _043403_, _043404_, _043405_, _043406_, _043407_, _043408_, _043409_, _043410_, _043411_, _043412_, _043413_, _043414_, _043415_, _043416_, _043417_, _043418_, _043419_, _043420_, _043421_, _043422_, _043423_, _043424_, _043425_, _043426_, _043427_, _043428_, _043429_, _043430_, _043431_, _043432_, _043433_, _043434_, _043435_, _043436_, _043437_, _043438_, _043439_, _043440_, _043441_, _043442_, _043443_, _043444_, _043445_, _043446_, _043447_, _043448_, _043449_, _043450_, _043451_, _043452_, _043453_, _043454_, _043455_, _043456_, _043457_, _043458_, _043459_, _043460_, _043461_, _043462_, _043463_, _043464_, _043465_, _043466_, _043467_, _043468_, _043469_, _043470_, _043471_, _043472_, _043473_, _043474_, _043475_, _043476_, _043477_, _043478_, _043479_, _043480_, _043481_, _043482_, _043483_, _043484_, _043485_, _043486_, _043487_, _043488_, _043489_, _043490_, _043491_, _043492_, _043493_, _043494_, _043495_, _043496_, _043497_, _043498_, _043499_, _043500_, _043501_, _043502_, _043503_, _043504_, _043505_, _043506_, _043507_, _043508_, _043509_, _043510_, _043511_, _043512_, _043513_, _043514_, _043515_, _043516_, _043517_, _043518_, _043519_, _043520_, _043521_, _043522_, _043523_, _043524_, _043525_, _043526_, _043527_, _043528_, _043529_, _043530_, _043531_, _043532_, _043533_, _043534_, _043535_, _043536_, _043537_, _043538_, _043539_, _043540_, _043541_, _043542_, _043543_, _043544_, _043545_, _043546_, _043547_, _043548_, _043549_, _043550_, _043551_, _043552_, _043553_, _043554_, _043555_, _043556_, _043557_, _043558_, _043559_, _043560_, _043561_, _043562_, _043563_, _043564_, _043565_, _043566_, _043567_, _043568_, _043569_, _043570_, _043571_, _043572_, _043573_, _043574_, _043575_, _043576_, _043577_, _043578_, _043579_, _043580_, _043581_, _043582_, _043583_, _043584_, _043585_, _043586_, _043587_, _043588_, _043589_, _043590_, _043591_, _043592_, _043593_, _043594_, _043595_, _043596_, _043597_, _043598_, _043599_, _043600_, _043601_, _043602_, _043603_, _043604_, _043605_, _043606_, _043607_, _043608_, _043609_, _043610_, _043611_, _043612_, _043613_, _043614_, _043615_, _043616_, _043617_, _043618_, _043619_, _043620_, _043621_, _043622_, _043623_, _043624_, _043625_, _043626_, _043627_, _043628_, _043629_, _043630_, _043631_, _043632_, _043633_, _043634_, _043635_, _043636_, _043637_, _043638_, _043639_, _043640_, _043641_, _043642_, _043643_, _043644_, _043645_, _043646_, _043647_, _043648_, _043649_, _043650_, _043651_, _043652_, _043653_, _043654_, _043655_, _043656_, _043657_, _043658_, _043659_, _043660_, _043661_, _043662_, _043663_, _043664_, _043665_, _043666_, _043667_, _043668_, _043669_, _043670_, _043671_, _043672_, _043673_, _043674_, _043675_, _043676_, _043677_, _043678_, _043679_, _043680_, _043681_, _043682_, _043683_, _043684_, _043685_, _043686_, _043687_, _043688_, _043689_, _043690_, _043691_, _043692_, _043693_, _043694_, _043695_, _043696_, _043697_, _043698_, _043699_, _043700_, _043701_, _043702_, _043703_, _043704_, _043705_, _043706_, _043707_, _043708_, _043709_, _043710_, _043711_, _043712_, _043713_, _043714_, _043715_, _043716_, _043717_, _043718_, _043719_, _043720_, _043721_, _043722_, _043723_, _043724_, _043725_, _043726_, _043727_, _043728_, _043729_, _043730_, _043731_, _043732_, _043733_, _043734_, _043735_, _043736_, _043737_, _043738_, _043739_, _043740_, _043741_, _043742_, _043743_, _043744_, _043745_, _043746_, _043747_, _043748_, _043749_, _043750_, _043751_, _043752_, _043753_, _043754_, _043755_, _043756_, _043757_, _043758_, _043759_, _043760_, _043761_, _043762_, _043763_, _043764_, _043765_, _043766_, _043767_, _043768_, _043769_, _043770_, _043771_, _043772_, _043773_, _043774_, _043775_, _043776_, _043777_, _043778_, _043779_, _043780_, _043781_, _043782_, _043783_, _043784_, _043785_, _043786_, _043787_, _043788_, _043789_, _043790_, _043791_, _043792_, _043793_, _043794_, _043795_, _043796_, _043797_, _043798_, _043799_, _043800_, _043801_, _043802_, _043803_, _043804_, _043805_, _043806_, _043807_, _043808_, _043809_, _043810_, _043811_, _043812_, _043813_, _043814_, _043815_, _043816_, _043817_, _043818_, _043819_, _043820_, _043821_, _043822_, _043823_, _043824_, _043825_, _043826_, _043827_, _043828_, _043829_, _043830_, _043831_, _043832_, _043833_, _043834_, _043835_, _043836_, _043837_, _043838_, _043839_, _043840_, _043841_, _043842_, _043843_, _043844_, _043845_, _043846_, _043847_, _043848_, _043849_, _043850_, _043851_, _043852_, _043853_, _043854_, _043855_, _043856_, _043857_, _043858_, _043859_, _043860_, _043861_, _043862_, _043863_, _043864_, _043865_, _043866_, _043867_, _043868_, _043869_, _043870_, _043871_, _043872_, _043873_, _043874_, _043875_, _043876_, _043877_, _043878_, _043879_, _043880_, _043881_, _043882_, _043883_, _043884_, _043885_, _043886_, _043887_, _043888_, _043889_, _043890_, _043891_, _043892_, _043893_, _043894_, _043895_, _043896_, _043897_, _043898_, _043899_, _043900_, _043901_, _043902_, _043903_, _043904_, _043905_, _043906_, _043907_, _043908_, _043909_, _043910_, _043911_, _043912_, _043913_, _043914_, _043915_, _043916_, _043917_, _043918_, _043919_, _043920_, _043921_, _043922_, _043923_, _043924_, _043925_, _043926_, _043927_, _043928_, _043929_, _043930_, _043931_, _043932_, _043933_, _043934_, _043935_, _043936_, _043937_, _043938_, _043939_, _043940_, _043941_, _043942_, _043943_, _043944_, _043945_, _043946_, _043947_, _043948_, _043949_, _043950_, _043951_, _043952_, _043953_, _043954_, _043955_, _043956_, _043957_, _043958_, _043959_, _043960_, _043961_, _043962_, _043963_, _043964_, _043965_, _043966_, _043967_, _043968_, _043969_, _043970_, _043971_, _043972_, _043973_, _043974_, _043975_, _043976_, _043977_, _043978_, _043979_, _043980_, _043981_, _043982_, _043983_, _043984_, _043985_, _043986_, _043987_, _043988_, _043989_, _043990_, _043991_, _043992_, _043993_, _043994_, _043995_, _043996_, _043997_, _043998_, _043999_, _044000_, _044001_, _044002_, _044003_, _044004_, _044005_, _044006_, _044007_, _044008_, _044009_, _044010_, _044011_, _044012_, _044013_, _044014_, _044015_, _044016_, _044017_, _044018_, _044019_, _044020_, _044021_, _044022_, _044023_, _044024_, _044025_, _044026_, _044027_, _044028_, _044029_, _044030_, _044031_, _044032_, _044033_, _044034_, _044035_, _044036_, _044037_, _044038_, _044039_, _044040_, _044041_, _044042_, _044043_, _044044_, _044045_, _044046_, _044047_, _044048_, _044049_, _044050_, _044051_, _044052_, _044053_, _044054_, _044055_, _044056_, _044057_, _044058_, _044059_, _044060_, _044061_, _044062_, _044063_, _044064_, _044065_, _044066_, _044067_, _044068_, _044069_, _044070_, _044071_, _044072_, _044073_, _044074_, _044075_, _044076_, _044077_, _044078_, _044079_, _044080_, _044081_, _044082_, _044083_, _044084_, _044085_, _044086_, _044087_, _044088_, _044089_, _044090_, _044091_, _044092_, _044093_, _044094_, _044095_, _044096_, _044097_, _044098_, _044099_, _044100_, _044101_, _044102_, _044103_, _044104_, _044105_, _044106_, _044107_, _044108_, _044109_, _044110_, _044111_, _044112_, _044113_, _044114_, _044115_, _044116_, _044117_, _044118_, _044119_, _044120_, _044121_, _044122_, _044123_, _044124_, _044125_, _044126_, _044127_, _044128_, _044129_, _044130_, _044131_, _044132_, _044133_, _044134_, _044135_, _044136_, _044137_, _044138_, _044139_, _044140_, _044141_, _044142_, _044143_, _044144_, _044145_, _044146_, _044147_, _044148_, _044149_, _044150_, _044151_, _044152_, _044153_, _044154_, _044155_, _044156_, _044157_, _044158_, _044159_, _044160_, _044161_, _044162_, _044163_, _044164_, _044165_, _044166_, _044167_, _044168_, _044169_, _044170_, _044171_, _044172_, _044173_, _044174_, _044175_, _044176_, _044177_, _044178_, _044179_, _044180_, _044181_, _044182_, _044183_, _044184_, _044185_, _044186_, _044187_, _044188_, _044189_, _044190_, _044191_, _044192_, _044193_, _044194_, _044195_, _044196_, _044197_, _044198_, _044199_, _044200_, _044201_, _044202_, _044203_, _044204_, _044205_, _044206_, _044207_, _044208_, _044209_, _044210_, _044211_, _044212_, _044213_, _044214_, _044215_, _044216_, _044217_, _044218_, _044219_, _044220_, _044221_, _044222_, _044223_, _044224_, _044225_, _044226_, _044227_, _044228_, _044229_, _044230_, _044231_, _044232_, _044233_, _044234_, _044235_, _044236_, _044237_, _044238_, _044239_, _044240_, _044241_, _044242_, _044243_, _044244_, _044245_, _044246_, _044247_, _044248_, _044249_, _044250_, _044251_, _044252_, _044253_, _044254_, _044255_, _044256_, _044257_, _044258_, _044259_, _044260_, _044261_, _044262_, _044263_, _044264_, _044265_, _044266_, _044267_, _044268_, _044269_, _044270_, _044271_, _044272_, _044273_, _044274_, _044275_, _044276_, _044277_, _044278_, _044279_, _044280_, _044281_, _044282_, _044283_, _044284_, _044285_, _044286_, _044287_, _044288_, _044289_, _044290_, _044291_, _044292_, _044293_, _044294_, _044295_, _044296_, _044297_, _044298_, _044299_, _044300_, _044301_, _044302_, _044303_, _044304_, _044305_, _044306_, _044307_, _044308_, _044309_, _044310_, _044311_, _044312_, _044313_, _044314_, _044315_, _044316_, _044317_, _044318_, _044319_, _044320_, _044321_, _044322_, _044323_, _044324_, _044325_, _044326_, _044327_, _044328_, _044329_, _044330_, _044331_, _044332_, _044333_, _044334_, _044335_, _044336_, _044337_, _044338_, _044339_, _044340_, _044341_, _044342_, _044343_, _044344_, _044345_, _044346_, _044347_, _044348_, _044349_, _044350_, _044351_, _044352_, _044353_, _044354_, _044355_, _044356_, _044357_, _044358_, _044359_, _044360_, _044361_, _044362_, _044363_, _044364_, _044365_, _044366_, _044367_, _044368_, _044369_, _044370_, _044371_, _044372_, _044373_, _044374_, _044375_, _044376_, _044377_, _044378_, _044379_, _044380_, _044381_, _044382_, _044383_, _044384_, _044385_, _044386_, _044387_, _044388_, _044389_, _044390_, _044391_, _044392_, _044393_, _044394_, _044395_, _044396_, _044397_, _044398_, _044399_, _044400_, _044401_, _044402_, _044403_, _044404_, _044405_, _044406_, _044407_, _044408_, _044409_, _044410_, _044411_, _044412_, _044413_, _044414_, _044415_, _044416_, _044417_, _044418_, _044419_, _044420_, _044421_, _044422_, _044423_, _044424_, _044425_, _044426_, _044427_, _044428_, _044429_, _044430_, _044431_, _044432_, _044433_, _044434_, _044435_, _044436_, _044437_, _044438_, _044439_, _044440_, _044441_, _044442_, _044443_, _044444_, _044445_, _044446_, _044447_, _044448_, _044449_, _044450_, _044451_, _044452_, _044453_, _044454_, _044455_, _044456_, _044457_, _044458_, _044459_, _044460_, _044461_, _044462_, _044463_, _044464_, _044465_, _044466_, _044467_, _044468_, _044469_, _044470_, _044471_, _044472_, _044473_, _044474_, _044475_, _044476_, _044477_, _044478_, _044479_, _044480_, _044481_, _044482_, _044483_, _044484_, _044485_, _044486_, _044487_, _044488_, _044489_, _044490_, _044491_, _044492_, _044493_, _044494_, _044495_, _044496_, _044497_, _044498_, _044499_, _044500_, _044501_, _044502_, _044503_, _044504_, _044505_, _044506_, _044507_, _044508_, _044509_, _044510_, _044511_, _044512_, _044513_, _044514_, _044515_, _044516_, _044517_, _044518_, _044519_, _044520_, _044521_, _044522_, _044523_, _044524_, _044525_, _044526_, _044527_, _044528_, _044529_, _044530_, _044531_, _044532_, _044533_, _044534_, _044535_, _044536_, _044537_, _044538_, _044539_, _044540_, _044541_, _044542_, _044543_, _044544_, _044545_, _044546_, _044547_, _044548_, _044549_, _044550_, _044551_, _044552_, _044553_, _044554_, _044555_, _044556_, _044557_, _044558_, _044559_, _044560_, _044561_, _044562_, _044563_, _044564_, _044565_, _044566_, _044567_, _044568_, _044569_, _044570_, _044571_, _044572_, _044573_, _044574_, _044575_, _044576_, _044577_, _044578_, _044579_, _044580_, _044581_, _044582_, _044583_, _044584_, _044585_, _044586_, _044587_, _044588_, _044589_, _044590_, _044591_, _044592_, _044593_, _044594_, _044595_, _044596_, _044597_, _044598_, _044599_, _044600_, _044601_, _044602_, _044603_, _044604_, _044605_, _044606_, _044607_, _044608_, _044609_, _044610_, _044611_, _044612_, _044613_, _044614_, _044615_, _044616_, _044617_, _044618_, _044619_, _044620_, _044621_, _044622_, _044623_, _044624_, _044625_, _044626_, _044627_, _044628_, _044629_, _044630_, _044631_, _044632_, _044633_, _044634_, _044635_, _044636_, _044637_, _044638_, _044639_, _044640_, _044641_, _044642_, _044643_, _044644_, _044645_, _044646_, _044647_, _044648_, _044649_, _044650_, _044651_, _044652_, _044653_, _044654_, _044655_, _044656_, _044657_, _044658_, _044659_, _044660_, _044661_, _044662_, _044663_, _044664_, _044665_, _044666_, _044667_, _044668_, _044669_, _044670_, _044671_, _044672_, _044673_, _044674_, _044675_, _044676_, _044677_, _044678_, _044679_, _044680_, _044681_, _044682_, _044683_, _044684_, _044685_, _044686_, _044687_, _044688_, _044689_, _044690_, _044691_, _044692_, _044693_, _044694_, _044695_, _044696_, _044697_, _044698_, _044699_, _044700_, _044701_, _044702_, _044703_, _044704_, _044705_, _044706_, _044707_, _044708_, _044709_, _044710_, _044711_, _044712_, _044713_, _044714_, _044715_, _044716_, _044717_, _044718_, _044719_, _044720_, _044721_, _044722_, _044723_, _044724_, _044725_, _044726_, _044727_, _044728_, _044729_, _044730_, _044731_, _044732_, _044733_, _044734_, _044735_, _044736_, _044737_, _044738_, _044739_, _044740_, _044741_, _044742_, _044743_, _044744_, _044745_, _044746_, _044747_, _044748_, _044749_, _044750_, _044751_, _044752_, _044753_, _044754_, _044755_, _044756_, _044757_, _044758_, _044759_, _044760_, _044761_, _044762_, _044763_, _044764_, _044765_, _044766_, _044767_, _044768_, _044769_, _044770_, _044771_, _044772_, _044773_, _044774_, _044775_, _044776_, _044777_, _044778_, _044779_, _044780_, _044781_, _044782_, _044783_, _044784_, _044785_, _044786_, _044787_, _044788_, _044789_, _044790_, _044791_, _044792_, _044793_, _044794_, _044795_, _044796_, _044797_, _044798_, _044799_, _044800_, _044801_, _044802_, _044803_, _044804_, _044805_, _044806_, _044807_, _044808_, _044809_, _044810_, _044811_, _044812_, _044813_, _044814_, _044815_, _044816_, _044817_, _044818_, _044819_, _044820_, _044821_, _044822_, _044823_, _044824_, _044825_, _044826_, _044827_, _044828_, _044829_, _044830_, _044831_, _044832_, _044833_, _044834_, _044835_, _044836_, _044837_, _044838_, _044839_, _044840_, _044841_, _044842_, _044843_, _044844_, _044845_, _044846_, _044847_, _044848_, _044849_, _044850_, _044851_, _044852_, _044853_, _044854_, _044855_, _044856_, _044857_, _044858_, _044859_, _044860_, _044861_, _044862_, _044863_, _044864_, _044865_, _044866_, _044867_, _044868_, _044869_, _044870_, _044871_, _044872_, _044873_, _044874_, _044875_, _044876_, _044877_, _044878_, _044879_, _044880_, _044881_, _044882_, _044883_, _044884_, _044885_, _044886_, _044887_, _044888_, _044889_, _044890_, _044891_, _044892_, _044893_, _044894_, _044895_, _044896_, _044897_, _044898_, _044899_, _044900_, _044901_, _044902_, _044903_, _044904_, _044905_, _044906_, _044907_, _044908_, _044909_, _044910_, _044911_, _044912_, _044913_, _044914_, _044915_, _044916_, _044917_, _044918_, _044919_, _044920_, _044921_, _044922_, _044923_, _044924_, _044925_, _044926_, _044927_, _044928_, _044929_, _044930_, _044931_, _044932_, _044933_, _044934_, _044935_, _044936_, _044937_, _044938_, _044939_, _044940_, _044941_, _044942_, _044943_, _044944_, _044945_, _044946_, _044947_, _044948_, _044949_, _044950_, _044951_, _044952_, _044953_, _044954_, _044955_, _044956_, _044957_, _044958_, _044959_, _044960_, _044961_, _044962_, _044963_, _044964_, _044965_, _044966_, _044967_, _044968_, _044969_, _044970_, _044971_, _044972_, _044973_, _044974_, _044975_, _044976_, _044977_, _044978_, _044979_, _044980_, _044981_, _044982_, _044983_, _044984_, _044985_, _044986_, _044987_, _044988_, _044989_, _044990_, _044991_, _044992_, _044993_, _044994_, _044995_, _044996_, _044997_, _044998_, _044999_, _045000_, _045001_, _045002_, _045003_, _045004_, _045005_, _045006_, _045007_, _045008_, _045009_, _045010_, _045011_, _045012_, _045013_, _045014_, _045015_, _045016_, _045017_, _045018_, _045019_, _045020_, _045021_, _045022_, _045023_, _045024_, _045025_, _045026_, _045027_, _045028_, _045029_, _045030_, _045031_, _045032_, _045033_, _045034_, _045035_, _045036_, _045037_, _045038_, _045039_, _045040_, _045041_, _045042_, _045043_, _045044_, _045045_, _045046_, _045047_, _045048_, _045049_, _045050_, _045051_, _045052_, _045053_, _045054_, _045055_, _045056_, _045057_, _045058_, _045059_, _045060_, _045061_, _045062_, _045063_, _045064_, _045065_, _045066_, _045067_, _045068_, _045069_, _045070_, _045071_, _045072_, _045073_, _045074_, _045075_, _045076_, _045077_, _045078_, _045079_, _045080_, _045081_, _045082_, _045083_, _045084_, _045085_, _045086_, _045087_, _045088_, _045089_, _045090_, _045091_, _045092_, _045093_, _045094_, _045095_, _045096_, _045097_, _045098_, _045099_, _045100_, _045101_, _045102_, _045103_, _045104_, _045105_, _045106_, _045107_, _045108_, _045109_, _045110_, _045111_, _045112_, _045113_, _045114_, _045115_, _045116_, _045117_, _045118_, _045119_, _045120_, _045121_, _045122_, _045123_, _045124_, _045125_, _045126_, _045127_, _045128_, _045129_, _045130_, _045131_, _045132_, _045133_, _045134_, _045135_, _045136_, _045137_, _045138_, _045139_, _045140_, _045141_, _045142_, _045143_, _045144_, _045145_, _045146_, _045147_, _045148_, _045149_, _045150_, _045151_, _045152_, _045153_, _045154_, _045155_, _045156_, _045157_, _045158_, _045159_, _045160_, _045161_, _045162_, _045163_, _045164_, _045165_, _045166_, _045167_, _045168_, _045169_, _045170_, _045171_, _045172_, _045173_, _045174_, _045175_, _045176_, _045177_, _045178_, _045179_, _045180_, _045181_, _045182_, _045183_, _045184_, _045185_, _045186_, _045187_, _045188_, _045189_, _045190_, _045191_, _045192_, _045193_, _045194_, _045195_, _045196_, _045197_, _045198_, _045199_, _045200_, _045201_, _045202_, _045203_, _045204_, _045205_, _045206_, _045207_, _045208_, _045209_, _045210_, _045211_, _045212_, _045213_, _045214_, _045215_, _045216_, _045217_, _045218_, _045219_, _045220_, _045221_, _045222_, _045223_, _045224_, _045225_, _045226_, _045227_, _045228_, _045229_, _045230_, _045231_, _045232_, _045233_, _045234_, _045235_, _045236_, _045237_, _045238_, _045239_, _045240_, _045241_, _045242_, _045243_, _045244_, _045245_, _045246_, _045247_, _045248_, _045249_, _045250_, _045251_, _045252_, _045253_, _045254_, _045255_, _045256_, _045257_, _045258_, _045259_, _045260_, _045261_, _045262_, _045263_, _045264_, _045265_, _045266_, _045267_, _045268_, _045269_, _045270_, _045271_, _045272_, _045273_, _045274_, _045275_, _045276_, _045277_, _045278_, _045279_, _045280_, _045281_, _045282_, _045283_, _045284_, _045285_, _045286_, _045287_, _045288_, _045289_, _045290_, _045291_, _045292_, _045293_, _045294_, _045295_, _045296_, _045297_, _045298_, _045299_, _045300_, _045301_, _045302_, _045303_, _045304_, _045305_, _045306_, _045307_, _045308_, _045309_, _045310_, _045311_, _045312_, _045313_, _045314_, _045315_, _045316_, _045317_, _045318_, _045319_, _045320_, _045321_, _045322_, _045323_, _045324_, _045325_, _045326_, _045327_, _045328_, _045329_, _045330_, _045331_, _045332_, _045333_, _045334_, _045335_, _045336_, _045337_, _045338_, _045339_, _045340_, _045341_, _045342_, _045343_, _045344_, _045345_, _045346_, _045347_, _045348_, _045349_, _045350_, _045351_, _045352_, _045353_, _045354_, _045355_, _045356_, _045357_, _045358_, _045359_, _045360_, _045361_, _045362_, _045363_, _045364_, _045365_, _045366_, _045367_, _045368_, _045369_, _045370_, _045371_, _045372_, _045373_, _045374_, _045375_, _045376_, _045377_, _045378_, _045379_, _045380_, _045381_, _045382_, _045383_, _045384_, _045385_, _045386_, _045387_, _045388_, _045389_, _045390_, _045391_, _045392_, _045393_, _045394_, _045395_, _045396_, _045397_, _045398_, _045399_, _045400_, _045401_, _045402_, _045403_, _045404_, _045405_, _045406_, _045407_, _045408_, _045409_, _045410_, _045411_, _045412_, _045413_, _045414_, _045415_, _045416_, _045417_, _045418_, _045419_, _045420_, _045421_, _045422_, _045423_, _045424_, _045425_, _045426_, _045427_, _045428_, _045429_, _045430_, _045431_, _045432_, _045433_, _045434_, _045435_, _045436_, _045437_, _045438_, _045439_, _045440_, _045441_, _045442_, _045443_, _045444_, _045445_, _045446_, _045447_, _045448_, _045449_, _045450_, _045451_, _045452_, _045453_, _045454_, _045455_, _045456_, _045457_, _045458_, _045459_, _045460_, _045461_, _045462_, _045463_, _045464_, _045465_, _045466_, _045467_, _045468_, _045469_, _045470_, _045471_, _045472_, _045473_, _045474_, _045475_, _045476_, _045477_, _045478_, _045479_, _045480_, _045481_, _045482_, _045483_, _045484_, _045485_, _045486_, _045487_, _045488_, _045489_, _045490_, _045491_, _045492_, _045493_, _045494_, _045495_, _045496_, _045497_, _045498_, _045499_, _045500_, _045501_, _045502_, _045503_, _045504_, _045505_, _045506_, _045507_, _045508_, _045509_, _045510_, _045511_, _045512_, _045513_, _045514_, _045515_, _045516_, _045517_, _045518_, _045519_, _045520_, _045521_, _045522_, _045523_, _045524_, _045525_, _045526_, _045527_, _045528_, _045529_, _045530_, _045531_, _045532_, _045533_, _045534_, _045535_, _045536_, _045537_, _045538_, _045539_, _045540_, _045541_, _045542_, _045543_, _045544_, _045545_, _045546_, _045547_, _045548_, _045549_, _045550_, _045551_, _045552_, _045553_, _045554_, _045555_, _045556_, _045557_, _045558_, _045559_, _045560_, _045561_, _045562_, _045563_, _045564_, _045565_, _045566_, _045567_, _045568_, _045569_, _045570_, _045571_, _045572_, _045573_, _045574_, _045575_, _045576_, _045577_, _045578_, _045579_, _045580_, _045581_, _045582_, _045583_, _045584_, _045585_, _045586_, _045587_, _045588_, _045589_, _045590_, _045591_, _045592_, _045593_, _045594_, _045595_, _045596_, _045597_, _045598_, _045599_, _045600_, _045601_, _045602_, _045603_, _045604_, _045605_, _045606_, _045607_, _045608_, _045609_, _045610_, _045611_, _045612_, _045613_, _045614_, _045615_, _045616_, _045617_, _045618_, _045619_, _045620_, _045621_, _045622_, _045623_, _045624_, _045625_, _045626_, _045627_, _045628_, _045629_, _045630_, _045631_, _045632_, _045633_, _045634_, _045635_, _045636_, _045637_, _045638_, _045639_, _045640_, _045641_, _045642_, _045643_, _045644_, _045645_, _045646_, _045647_, _045648_, _045649_, _045650_, _045651_, _045652_, _045653_, _045654_, _045655_, _045656_, _045657_, _045658_, _045659_, _045660_, _045661_, _045662_, _045663_, _045664_, _045665_, _045666_, _045667_, _045668_, _045669_, _045670_, _045671_, _045672_, _045673_, _045674_, _045675_, _045676_, _045677_, _045678_, _045679_, _045680_, _045681_, _045682_, _045683_, _045684_, _045685_, _045686_, _045687_, _045688_, _045689_, _045690_, _045691_, _045692_, _045693_, _045694_, _045695_, _045696_, _045697_, _045698_, _045699_, _045700_, _045701_, _045702_, _045703_, _045704_, _045705_, _045706_, _045707_, _045708_, _045709_, _045710_, _045711_, _045712_, _045713_, _045714_, _045715_, _045716_, _045717_, _045718_, _045719_, _045720_, _045721_, _045722_, _045723_, _045724_, _045725_, _045726_, _045727_, _045728_, _045729_, _045730_, _045731_, _045732_, _045733_, _045734_, _045735_, _045736_, _045737_, _045738_, _045739_, _045740_, _045741_, _045742_, _045743_, _045744_, _045745_, _045746_, _045747_, _045748_, _045749_, _045750_, _045751_, _045752_, _045753_, _045754_, _045755_, _045756_, _045757_, _045758_, _045759_, _045760_, _045761_, _045762_, _045763_, _045764_, _045765_, _045766_, _045767_, _045768_, _045769_, _045770_, _045771_, _045772_, _045773_, _045774_, _045775_, _045776_, _045777_, _045778_, _045779_, _045780_, _045781_, _045782_, _045783_, _045784_, _045785_, _045786_, _045787_, _045788_, _045789_, _045790_, _045791_, _045792_, _045793_, _045794_, _045795_, _045796_, _045797_, _045798_, _045799_, _045800_, _045801_, _045802_, _045803_, _045804_, _045805_, _045806_, _045807_, _045808_, _045809_, _045810_, _045811_, _045812_, _045813_, _045814_, _045815_, _045816_, _045817_, _045818_, _045819_, _045820_, _045821_, _045822_, _045823_, _045824_, _045825_, _045826_, _045827_, _045828_, _045829_, _045830_, _045831_, _045832_, _045833_, _045834_, _045835_, _045836_, _045837_, _045838_, _045839_, _045840_, _045841_, _045842_, _045843_, _045844_, _045845_, _045846_, _045847_, _045848_, _045849_, _045850_, _045851_, _045852_, _045853_, _045854_, _045855_, _045856_, _045857_, _045858_, _045859_, _045860_, _045861_, _045862_, _045863_, _045864_, _045865_, _045866_, _045867_, _045868_, _045869_, _045870_, _045871_, _045872_, _045873_, _045874_, _045875_, _045876_, _045877_, _045878_, _045879_, _045880_, _045881_, _045882_, _045883_, _045884_, _045885_, _045886_, _045887_, _045888_, _045889_, _045890_, _045891_, _045892_, _045893_, _045894_, _045895_, _045896_, _045897_, _045898_, _045899_, _045900_, _045901_, _045902_, _045903_, _045904_, _045905_, _045906_, _045907_, _045908_, _045909_, _045910_, _045911_, _045912_, _045913_, _045914_, _045915_, _045916_, _045917_, _045918_, _045919_, _045920_, _045921_, _045922_, _045923_, _045924_, _045925_, _045926_, _045927_, _045928_, _045929_, _045930_, _045931_, _045932_, _045933_, _045934_, _045935_, _045936_, _045937_, _045938_, _045939_, _045940_, _045941_, _045942_, _045943_, _045944_, _045945_, _045946_, _045947_, _045948_, _045949_, _045950_, _045951_, _045952_, _045953_, _045954_, _045955_, _045956_, _045957_, _045958_, _045959_, _045960_, _045961_, _045962_, _045963_, _045964_, _045965_, _045966_, _045967_, _045968_, _045969_, _045970_, _045971_, _045972_, _045973_, _045974_, _045975_, _045976_, _045977_, _045978_, _045979_, _045980_, _045981_, _045982_, _045983_, _045984_, _045985_, _045986_, _045987_, _045988_, _045989_, _045990_, _045991_, _045992_, _045993_, _045994_, _045995_, _045996_, _045997_, _045998_, _045999_, _046000_, _046001_, _046002_, _046003_, _046004_, _046005_, _046006_, _046007_, _046008_, _046009_, _046010_, _046011_, _046012_, _046013_, _046014_, _046015_, _046016_, _046017_, _046018_, _046019_, _046020_, _046021_, _046022_, _046023_, _046024_, _046025_, _046026_, _046027_, _046028_, _046029_, _046030_, _046031_, _046032_, _046033_, _046034_, _046035_, _046036_, _046037_, _046038_, _046039_, _046040_, _046041_, _046042_, _046043_, _046044_, _046045_, _046046_, _046047_, _046048_, _046049_, _046050_, _046051_, _046052_, _046053_, _046054_, _046055_, _046056_, _046057_, _046058_, _046059_, _046060_, _046061_, _046062_, _046063_, _046064_, _046065_, _046066_, _046067_, _046068_, _046069_, _046070_, _046071_, _046072_, _046073_, _046074_, _046075_, _046076_, _046077_, _046078_, _046079_, _046080_, _046081_, _046082_, _046083_, _046084_, _046085_, _046086_, _046087_, _046088_, _046089_, _046090_, _046091_, _046092_, _046093_, _046094_, _046095_, _046096_, _046097_, _046098_, _046099_, _046100_, _046101_, _046102_, _046103_, _046104_, _046105_, _046106_, _046107_, _046108_, _046109_, _046110_, _046111_, _046112_, _046113_, _046114_, _046115_, _046116_, _046117_, _046118_, _046119_, _046120_, _046121_, _046122_, _046123_, _046124_, _046125_, _046126_, _046127_, _046128_, _046129_, _046130_, _046131_, _046132_, _046133_, _046134_, _046135_, _046136_, _046137_, _046138_, _046139_, _046140_, _046141_, _046142_, _046143_, _046144_, _046145_, _046146_, _046147_, _046148_, _046149_, _046150_, _046151_, _046152_, _046153_, _046154_, _046155_, _046156_, _046157_, _046158_, _046159_, _046160_, _046161_, _046162_, _046163_, _046164_, _046165_, _046166_, _046167_, _046168_, _046169_, _046170_, _046171_, _046172_, _046173_, _046174_, _046175_, _046176_, _046177_, _046178_, _046179_, _046180_, _046181_, _046182_, _046183_, _046184_, _046185_, _046186_, _046187_, _046188_, _046189_, _046190_, _046191_, _046192_, _046193_, _046194_, _046195_, _046196_, _046197_, _046198_, _046199_, _046200_, _046201_, _046202_, _046203_, _046204_, _046205_, _046206_, _046207_, _046208_, _046209_, _046210_, _046211_, _046212_, _046213_, _046214_, _046215_, _046216_, _046217_, _046218_, _046219_, _046220_, _046221_, _046222_, _046223_, _046224_, _046225_, _046226_, _046227_, _046228_, _046229_, _046230_, _046231_, _046232_, _046233_, _046234_, _046235_, _046236_, _046237_, _046238_, _046239_, _046240_, _046241_, _046242_, _046243_, _046244_, _046245_, _046246_, _046247_, _046248_, _046249_, _046250_, _046251_, _046252_, _046253_, _046254_, _046255_, _046256_, _046257_, _046258_, _046259_, _046260_, _046261_, _046262_, _046263_, _046264_, _046265_, _046266_, _046267_, _046268_, _046269_, _046270_, _046271_, _046272_, _046273_, _046274_, _046275_, _046276_, _046277_, _046278_, _046279_, _046280_, _046281_, _046282_, _046283_, _046284_, _046285_, _046286_, _046287_, _046288_, _046289_, _046290_, _046291_, _046292_, _046293_, _046294_, _046295_, _046296_, _046297_, _046298_, _046299_, _046300_, _046301_, _046302_, _046303_, _046304_, _046305_, _046306_, _046307_, _046308_, _046309_, _046310_, _046311_, _046312_, _046313_, _046314_, _046315_, _046316_, _046317_, _046318_, _046319_, _046320_, _046321_, _046322_, _046323_, _046324_, _046325_, _046326_, _046327_, _046328_, _046329_, _046330_, _046331_, _046332_, _046333_, _046334_, _046335_, _046336_, _046337_, _046338_, _046339_, _046340_, _046341_, _046342_, _046343_, _046344_, _046345_, _046346_, _046347_, _046348_, _046349_, _046350_, _046351_, _046352_, _046353_, _046354_, _046355_, _046356_, _046357_, _046358_, _046359_, _046360_, _046361_, _046362_, _046363_, _046364_, _046365_, _046366_, _046367_, _046368_, _046369_, _046370_, _046371_, _046372_, _046373_, _046374_, _046375_, _046376_, _046377_, _046378_, _046379_, _046380_, _046381_, _046382_, _046383_, _046384_, _046385_, _046386_, _046387_, _046388_, _046389_, _046390_, _046391_, _046392_, _046393_, _046394_, _046395_, _046396_, _046397_, _046398_, _046399_, _046400_, _046401_, _046402_, _046403_, _046404_, _046405_, _046406_, _046407_, _046408_, _046409_, _046410_, _046411_, _046412_, _046413_, _046414_, _046415_, _046416_, _046417_, _046418_, _046419_, _046420_, _046421_, _046422_, _046423_, _046424_, _046425_, _046426_, _046427_, _046428_, _046429_, _046430_, _046431_, _046432_, _046433_, _046434_, _046435_, _046436_, _046437_, _046438_, _046439_, _046440_, _046441_, _046442_, _046443_, _046444_, _046445_, _046446_, _046447_, _046448_, _046449_, _046450_, _046451_, _046452_, _046453_, _046454_, _046455_, _046456_, _046457_, _046458_, _046459_, _046460_, _046461_, _046462_, _046463_, _046464_, _046465_, _046466_, _046467_, _046468_, _046469_, _046470_, _046471_, _046472_, _046473_, _046474_, _046475_, _046476_, _046477_, _046478_, _046479_, _046480_, _046481_, _046482_, _046483_, _046484_, _046485_, _046486_, _046487_, _046488_, _046489_, _046490_, _046491_, _046492_, _046493_, _046494_, _046495_, _046496_, _046497_, _046498_, _046499_, _046500_, _046501_, _046502_, _046503_, _046504_, _046505_, _046506_, _046507_, _046508_, _046509_, _046510_, _046511_, _046512_, _046513_, _046514_, _046515_, _046516_, _046517_, _046518_, _046519_, _046520_, _046521_, _046522_, _046523_, _046524_, _046525_, _046526_, _046527_, _046528_, _046529_, _046530_, _046531_, _046532_, _046533_, _046534_, _046535_, _046536_, _046537_, _046538_, _046539_, _046540_, _046541_, _046542_, _046543_, _046544_, _046545_, _046546_, _046547_, _046548_, _046549_, _046550_, _046551_, _046552_, _046553_, _046554_, _046555_, _046556_, _046557_, _046558_, _046559_, _046560_, _046561_, _046562_, _046563_, _046564_, _046565_, _046566_, _046567_, _046568_, _046569_, _046570_, _046571_, _046572_, _046573_, _046574_, _046575_, _046576_, _046577_, _046578_, _046579_, _046580_, _046581_, _046582_, _046583_, _046584_, _046585_, _046586_, _046587_, _046588_, _046589_, _046590_, _046591_, _046592_, _046593_, _046594_, _046595_, _046596_, _046597_, _046598_, _046599_, _046600_, _046601_, _046602_, _046603_, _046604_, _046605_, _046606_, _046607_, _046608_, _046609_, _046610_, _046611_, _046612_, _046613_, _046614_, _046615_, _046616_, _046617_, _046618_, _046619_, _046620_, _046621_, _046622_, _046623_, _046624_, _046625_, _046626_, _046627_, _046628_, _046629_, _046630_, _046631_, _046632_, _046633_, _046634_, _046635_, _046636_, _046637_, _046638_, _046639_, _046640_, _046641_, _046642_, _046643_, _046644_, _046645_, _046646_, _046647_, _046648_, _046649_, _046650_, _046651_, _046652_, _046653_, _046654_, _046655_, _046656_, _046657_, _046658_, _046659_, _046660_, _046661_, _046662_, _046663_, _046664_, _046665_, _046666_, _046667_, _046668_, _046669_, _046670_, _046671_, _046672_, _046673_, _046674_, _046675_, _046676_, _046677_, _046678_, _046679_, _046680_, _046681_, _046682_, _046683_, _046684_, _046685_, _046686_, _046687_, _046688_, _046689_, _046690_, _046691_, _046692_, _046693_, _046694_, _046695_, _046696_, _046697_, _046698_, _046699_, _046700_, _046701_, _046702_, _046703_, _046704_, _046705_, _046706_, _046707_, _046708_, _046709_, _046710_, _046711_, _046712_, _046713_, _046714_, _046715_, _046716_, _046717_, _046718_, _046719_, _046720_, _046721_, _046722_, _046723_, _046724_, _046725_, _046726_, _046727_, _046728_, _046729_, _046730_, _046731_, _046732_, _046733_, _046734_, _046735_, _046736_, _046737_, _046738_, _046739_, _046740_, _046741_, _046742_, _046743_, _046744_, _046745_, _046746_, _046747_, _046748_, _046749_, _046750_, _046751_, _046752_, _046753_, _046754_, _046755_, _046756_, _046757_, _046758_, _046759_, _046760_, _046761_, _046762_, _046763_, _046764_, _046765_, _046766_, _046767_, _046768_, _046769_, _046770_, _046771_, _046772_, _046773_, _046774_, _046775_, _046776_, _046777_, _046778_, _046779_, _046780_, _046781_, _046782_, _046783_, _046784_, _046785_, _046786_, _046787_, _046788_, _046789_, _046790_, _046791_, _046792_, _046793_, _046794_, _046795_, _046796_, _046797_, _046798_, _046799_, _046800_, _046801_, _046802_, _046803_, _046804_, _046805_, _046806_, _046807_, _046808_, _046809_, _046810_, _046811_, _046812_, _046813_, _046814_, _046815_, _046816_, _046817_, _046818_, _046819_, _046820_, _046821_, _046822_, _046823_, _046824_, _046825_, _046826_, _046827_, _046828_, _046829_, _046830_, _046831_, _046832_, _046833_, _046834_, _046835_, _046836_, _046837_, _046838_, _046839_, _046840_, _046841_, _046842_, _046843_, _046844_, _046845_, _046846_, _046847_, _046848_, _046849_, _046850_, _046851_, _046852_, _046853_, _046854_, _046855_, _046856_, _046857_, _046858_, _046859_, _046860_, _046861_, _046862_, _046863_, _046864_, _046865_, _046866_, _046867_, _046868_, _046869_, _046870_, _046871_, _046872_, _046873_, _046874_, _046875_, _046876_, _046877_, _046878_, _046879_, _046880_, _046881_, _046882_, _046883_, _046884_, _046885_, _046886_, _046887_, _046888_, _046889_, _046890_, _046891_, _046892_, _046893_, _046894_, _046895_, _046896_, _046897_, _046898_, _046899_, _046900_, _046901_, _046902_, _046903_, _046904_, _046905_, _046906_, _046907_, _046908_, _046909_, _046910_, _046911_, _046912_, _046913_, _046914_, _046915_, _046916_, _046917_, _046918_, _046919_, _046920_, _046921_, _046922_, _046923_, _046924_, _046925_, _046926_, _046927_, _046928_, _046929_, _046930_, _046931_, _046932_, _046933_, _046934_, _046935_, _046936_, _046937_, _046938_, _046939_, _046940_, _046941_, _046942_, _046943_, _046944_, _046945_, _046946_, _046947_, _046948_, _046949_, _046950_, _046951_, _046952_, _046953_, _046954_, _046955_, _046956_, _046957_, _046958_, _046959_, _046960_, _046961_, _046962_, _046963_, _046964_, _046965_, _046966_, _046967_, _046968_, _046969_, _046970_, _046971_, _046972_, _046973_, _046974_, _046975_, _046976_, _046977_, _046978_, _046979_, _046980_, _046981_, _046982_, _046983_, _046984_, _046985_, _046986_, _046987_, _046988_, _046989_, _046990_, _046991_, _046992_, _046993_, _046994_, _046995_, _046996_, _046997_, _046998_, _046999_, _047000_, _047001_, _047002_, _047003_, _047004_, _047005_, _047006_, _047007_, _047008_, _047009_, _047010_, _047011_, _047012_, _047013_, _047014_, _047015_, _047016_, _047017_, _047018_, _047019_, _047020_, _047021_, _047022_, _047023_, _047024_, _047025_, _047026_, _047027_, _047028_, _047029_, _047030_, _047031_, _047032_, _047033_, _047034_, _047035_, _047036_, _047037_, _047038_, _047039_, _047040_, _047041_, _047042_, _047043_, _047044_, _047045_, _047046_, _047047_, _047048_, _047049_, _047050_, _047051_, _047052_, _047053_, _047054_, _047055_, _047056_, _047057_, _047058_, _047059_, _047060_, _047061_, _047062_, _047063_, _047064_, _047065_, _047066_, _047067_, _047068_, _047069_, _047070_, _047071_, _047072_, _047073_, _047074_, _047075_, _047076_, _047077_, _047078_, _047079_, _047080_, _047081_, _047082_, _047083_, _047084_, _047085_, _047086_, _047087_, _047088_, _047089_, _047090_, _047091_, _047092_, _047093_, _047094_, _047095_, _047096_, _047097_, _047098_, _047099_, _047100_, _047101_, _047102_, _047103_, _047104_, _047105_, _047106_, _047107_, _047108_, _047109_, _047110_, _047111_, _047112_, _047113_, _047114_, _047115_, _047116_, _047117_, _047118_, _047119_, _047120_, _047121_, _047122_, _047123_, _047124_, _047125_, _047126_, _047127_, _047128_, _047129_, _047130_, _047131_, _047132_, _047133_, _047134_, _047135_, _047136_, _047137_, _047138_, _047139_, _047140_, _047141_, _047142_, _047143_, _047144_, _047145_, _047146_, _047147_, _047148_, _047149_, _047150_, _047151_, _047152_, _047153_, _047154_, _047155_, _047156_, _047157_, _047158_, _047159_, _047160_, _047161_, _047162_, _047163_, _047164_, _047165_, _047166_, _047167_, _047168_, _047169_, _047170_, _047171_, _047172_, _047173_, _047174_, _047175_, _047176_, _047177_, _047178_, _047179_, _047180_, _047181_, _047182_, _047183_, _047184_, _047185_, _047186_, _047187_, _047188_, _047189_, _047190_, _047191_, _047192_, _047193_, _047194_, _047195_, _047196_, _047197_, _047198_, _047199_, _047200_, _047201_, _047202_, _047203_, _047204_, _047205_, _047206_, _047207_, _047208_, _047209_, _047210_, _047211_, _047212_, _047213_, _047214_, _047215_, _047216_, _047217_, _047218_, _047219_, _047220_, _047221_, _047222_, _047223_, _047224_, _047225_, _047226_, _047227_, _047228_, _047229_, _047230_, _047231_, _047232_, _047233_, _047234_, _047235_, _047236_, _047237_, _047238_, _047239_, _047240_, _047241_, _047242_, _047243_, _047244_, _047245_, _047246_, _047247_, _047248_, _047249_, _047250_, _047251_, _047252_, _047253_, _047254_, _047255_, _047256_, _047257_, _047258_, _047259_, _047260_, _047261_, _047262_, _047263_, _047264_, _047265_, _047266_, _047267_, _047268_, _047269_, _047270_, _047271_, _047272_, _047273_, _047274_, _047275_, _047276_, _047277_, _047278_, _047279_, _047280_, _047281_, _047282_, _047283_, _047284_, _047285_, _047286_, _047287_, _047288_, _047289_, _047290_, _047291_, _047292_, _047293_, _047294_, _047295_, _047296_, _047297_, _047298_, _047299_, _047300_, _047301_, _047302_, _047303_, _047304_, _047305_, _047306_, _047307_, _047308_, _047309_, _047310_, _047311_, _047312_, _047313_, _047314_, _047315_, _047316_, _047317_, _047318_, _047319_, _047320_, _047321_, _047322_, _047323_, _047324_, _047325_, _047326_, _047327_, _047328_, _047329_, _047330_, _047331_, _047332_, _047333_, _047334_, _047335_, _047336_, _047337_, _047338_, _047339_, _047340_, _047341_, _047342_, _047343_, _047344_, _047345_, _047346_, _047347_, _047348_, _047349_, _047350_, _047351_, _047352_, _047353_, _047354_, _047355_, _047356_, _047357_, _047358_, _047359_, _047360_, _047361_, _047362_, _047363_, _047364_, _047365_, _047366_, _047367_, _047368_, _047369_, _047370_, _047371_, _047372_, _047373_, _047374_, _047375_, _047376_, _047377_, _047378_, _047379_, _047380_, _047381_, _047382_, _047383_, _047384_, _047385_, _047386_, _047387_, _047388_, _047389_, _047390_, _047391_, _047392_, _047393_, _047394_, _047395_, _047396_, _047397_, _047398_, _047399_, _047400_, _047401_, _047402_, _047403_, _047404_, _047405_, _047406_, _047407_, _047408_, _047409_, _047410_, _047411_, _047412_, _047413_, _047414_, _047415_, _047416_, _047417_, _047418_, _047419_, _047420_, _047421_, _047422_, _047423_, _047424_, _047425_, _047426_, _047427_, _047428_, _047429_, _047430_, _047431_, _047432_, _047433_, _047434_, _047435_, _047436_, _047437_, _047438_, _047439_, _047440_, _047441_, _047442_, _047443_, _047444_, _047445_, _047446_, _047447_, _047448_, _047449_, _047450_, _047451_, _047452_, _047453_, _047454_, _047455_, _047456_, _047457_, _047458_, _047459_, _047460_, _047461_, _047462_, _047463_, _047464_, _047465_, _047466_, _047467_, _047468_, _047469_, _047470_, _047471_, _047472_, _047473_, _047474_, _047475_, _047476_, _047477_, _047478_, _047479_, _047480_, _047481_, _047482_, _047483_, _047484_, _047485_, _047486_, _047487_, _047488_, _047489_, _047490_, _047491_, _047492_, _047493_, _047494_, _047495_, _047496_, _047497_, _047498_, _047499_, _047500_, _047501_, _047502_, _047503_, _047504_, _047505_, _047506_, _047507_, _047508_, _047509_, _047510_, _047511_, _047512_, _047513_, _047514_, _047515_, _047516_, _047517_, _047518_, _047519_, _047520_, _047521_, _047522_, _047523_, _047524_, _047525_, _047526_, _047527_, _047528_, _047529_, _047530_, _047531_, _047532_, _047533_, _047534_, _047535_, _047536_, _047537_, _047538_, _047539_, _047540_, _047541_, _047542_, _047543_, _047544_, _047545_, _047546_, _047547_, _047548_, _047549_, _047550_, _047551_, _047552_, _047553_, _047554_, _047555_, _047556_, _047557_, _047558_, _047559_, _047560_, _047561_, _047562_, _047563_, _047564_, _047565_, _047566_, _047567_, _047568_, _047569_, _047570_, _047571_, _047572_, _047573_, _047574_, _047575_, _047576_, _047577_, _047578_, _047579_, _047580_, _047581_, _047582_, _047583_, _047584_, _047585_, _047586_, _047587_, _047588_, _047589_, _047590_, _047591_, _047592_, _047593_, _047594_, _047595_, _047596_, _047597_, _047598_, _047599_, _047600_, _047601_, _047602_, _047603_, _047604_, _047605_, _047606_, _047607_, _047608_, _047609_, _047610_, _047611_, _047612_, _047613_, _047614_, _047615_, _047616_, _047617_, _047618_, _047619_, _047620_, _047621_, _047622_, _047623_, _047624_, _047625_, _047626_, _047627_, _047628_, _047629_, _047630_, _047631_, _047632_, _047633_, _047634_, _047635_, _047636_, _047637_, _047638_, _047639_, _047640_, _047641_, _047642_, _047643_, _047644_, _047645_, _047646_, _047647_, _047648_, _047649_, _047650_, _047651_, _047652_, _047653_, _047654_, _047655_, _047656_, _047657_, _047658_, _047659_, _047660_, _047661_, _047662_, _047663_, _047664_, _047665_, _047666_, _047667_, _047668_, _047669_, _047670_, _047671_, _047672_, _047673_, _047674_, _047675_, _047676_, _047677_, _047678_, _047679_, _047680_, _047681_, _047682_, _047683_, _047684_, _047685_, _047686_, _047687_, _047688_, _047689_, _047690_, _047691_, _047692_, _047693_, _047694_, _047695_, _047696_, _047697_, _047698_, _047699_, _047700_, _047701_, _047702_, _047703_, _047704_, _047705_, _047706_, _047707_, _047708_, _047709_, _047710_, _047711_, _047712_, _047713_, _047714_, _047715_, _047716_, _047717_, _047718_, _047719_, _047720_, _047721_, _047722_, _047723_, _047724_, _047725_, _047726_, _047727_, _047728_, _047729_, _047730_, _047731_, _047732_, _047733_, _047734_, _047735_, _047736_, _047737_, _047738_, _047739_, _047740_, _047741_, _047742_, _047743_, _047744_, _047745_, _047746_, _047747_, _047748_, _047749_, _047750_, _047751_, _047752_, _047753_, _047754_, _047755_, _047756_, _047757_, _047758_, _047759_, _047760_, _047761_, _047762_, _047763_, _047764_, _047765_, _047766_, _047767_, _047768_, _047769_, _047770_, _047771_, _047772_, _047773_, _047774_, _047775_, _047776_, _047777_, _047778_, _047779_, _047780_, _047781_, _047782_, _047783_, _047784_, _047785_, _047786_, _047787_, _047788_, _047789_, _047790_, _047791_, _047792_, _047793_, _047794_, _047795_, _047796_, _047797_, _047798_, _047799_, _047800_, _047801_, _047802_, _047803_, _047804_, _047805_, _047806_, _047807_, _047808_, _047809_, _047810_, _047811_, _047812_, _047813_, _047814_, _047815_, _047816_, _047817_, _047818_, _047819_, _047820_, _047821_, _047822_, _047823_, _047824_, _047825_, _047826_, _047827_, _047828_, _047829_, _047830_, _047831_, _047832_, _047833_, _047834_, _047835_, _047836_, _047837_, _047838_, _047839_, _047840_, _047841_, _047842_, _047843_, _047844_, _047845_, _047846_, _047847_, _047848_, _047849_, _047850_, _047851_, _047852_, _047853_, _047854_, _047855_, _047856_, _047857_, _047858_, _047859_, _047860_, _047861_, _047862_, _047863_, _047864_, _047865_, _047866_, _047867_, _047868_, _047869_, _047870_, _047871_, _047872_, _047873_, _047874_, _047875_, _047876_, _047877_, _047878_, _047879_, _047880_, _047881_, _047882_, _047883_, _047884_, _047885_, _047886_, _047887_, _047888_, _047889_, _047890_, _047891_, _047892_, _047893_, _047894_, _047895_, _047896_, _047897_, _047898_, _047899_, _047900_, _047901_, _047902_, _047903_, _047904_, _047905_, _047906_, _047907_, _047908_, _047909_, _047910_, _047911_, _047912_, _047913_, _047914_, _047915_, _047916_, _047917_, _047918_, _047919_, _047920_, _047921_, _047922_, _047923_, _047924_, _047925_, _047926_, _047927_, _047928_, _047929_, _047930_, _047931_, _047932_, _047933_, _047934_, _047935_, _047936_, _047937_, _047938_, _047939_, _047940_, _047941_, _047942_, _047943_, _047944_, _047945_, _047946_, _047947_, _047948_, _047949_, _047950_, _047951_, _047952_, _047953_, _047954_, _047955_, _047956_, _047957_, _047958_, _047959_, _047960_, _047961_, _047962_, _047963_, _047964_, _047965_, _047966_, _047967_, _047968_, _047969_, _047970_, _047971_, _047972_, _047973_, _047974_, _047975_, _047976_, _047977_, _047978_, _047979_, _047980_, _047981_, _047982_, _047983_, _047984_, _047985_, _047986_, _047987_, _047988_, _047989_, _047990_, _047991_, _047992_, _047993_, _047994_, _047995_, _047996_, _047997_, _047998_, _047999_, _048000_, _048001_, _048002_, _048003_, _048004_, _048005_, _048006_, _048007_, _048008_, _048009_, _048010_, _048011_, _048012_, _048013_, _048014_, _048015_, _048016_, _048017_, _048018_, _048019_, _048020_, _048021_, _048022_, _048023_, _048024_, _048025_, _048026_, _048027_, _048028_, _048029_, _048030_, _048031_, _048032_, _048033_, _048034_, _048035_, _048036_, _048037_, _048038_, _048039_, _048040_, _048041_, _048042_, _048043_, _048044_, _048045_, _048046_, _048047_, _048048_, _048049_, _048050_, _048051_, _048052_, _048053_, _048054_, _048055_, _048056_, _048057_, _048058_, _048059_, _048060_, _048061_, _048062_, _048063_, _048064_, _048065_, _048066_, _048067_, _048068_, _048069_, _048070_, _048071_, _048072_, _048073_, _048074_, _048075_, _048076_, _048077_, _048078_, _048079_, _048080_, _048081_, _048082_, _048083_, _048084_, _048085_, _048086_, _048087_, _048088_, _048089_, _048090_, _048091_, _048092_, _048093_, _048094_, _048095_, _048096_, _048097_, _048098_, _048099_, _048100_, _048101_, _048102_, _048103_, _048104_, _048105_, _048106_, _048107_, _048108_, _048109_, _048110_, _048111_, _048112_, _048113_, _048114_, _048115_, _048116_, _048117_, _048118_, _048119_, _048120_, _048121_, _048122_, _048123_, _048124_, _048125_, _048126_, _048127_, _048128_, _048129_, _048130_, _048131_, _048132_, _048133_, _048134_, _048135_, _048136_, _048137_, _048138_, _048139_, _048140_, _048141_, _048142_, _048143_, _048144_, _048145_, _048146_, _048147_, _048148_, _048149_, _048150_, _048151_, _048152_, _048153_, _048154_, _048155_, _048156_, _048157_, _048158_, _048159_, _048160_, _048161_, _048162_, _048163_, _048164_, _048165_, _048166_, _048167_, _048168_, _048169_, _048170_, _048171_, _048172_, _048173_, _048174_, _048175_, _048176_, _048177_, _048178_, _048179_, _048180_, _048181_, _048182_, _048183_, _048184_, _048185_, _048186_, _048187_, _048188_, _048189_, _048190_, _048191_, _048192_, _048193_, _048194_, _048195_, _048196_, _048197_, _048198_, _048199_, _048200_, _048201_, _048202_, _048203_, _048204_, _048205_, _048206_, _048207_, _048208_, _048209_, _048210_, _048211_, _048212_, _048213_, _048214_, _048215_, _048216_, _048217_, _048218_, _048219_, _048220_, _048221_, _048222_, _048223_, _048224_, _048225_, _048226_, _048227_, _048228_, _048229_, _048230_, _048231_, _048232_, _048233_, _048234_, _048235_, _048236_, _048237_, _048238_, _048239_, _048240_, _048241_, _048242_, _048243_, _048244_, _048245_, _048246_, _048247_, _048248_, _048249_, _048250_, _048251_, _048252_, _048253_, _048254_, _048255_, _048256_, _048257_, _048258_, _048259_, _048260_, _048261_, _048262_, _048263_, _048264_, _048265_, _048266_, _048267_, _048268_, _048269_, _048270_, _048271_, _048272_, _048273_, _048274_, _048275_, _048276_, _048277_, _048278_, _048279_, _048280_, _048281_, _048282_, _048283_, _048284_, _048285_, _048286_, _048287_, _048288_, _048289_, _048290_, _048291_, _048292_, _048293_, _048294_, _048295_, _048296_, _048297_, _048298_, _048299_, _048300_, _048301_, _048302_, _048303_, _048304_, _048305_, _048306_, _048307_, _048308_, _048309_, _048310_, _048311_, _048312_, _048313_, _048314_, _048315_, _048316_, _048317_, _048318_, _048319_, _048320_, _048321_, _048322_, _048323_, _048324_, _048325_, _048326_, _048327_, _048328_, _048329_, _048330_, _048331_, _048332_, _048333_, _048334_, _048335_, _048336_, _048337_, _048338_, _048339_, _048340_, _048341_, _048342_, _048343_, _048344_, _048345_, _048346_, _048347_, _048348_, _048349_, _048350_, _048351_, _048352_, _048353_, _048354_, _048355_, _048356_, _048357_, _048358_, _048359_, _048360_, _048361_, _048362_, _048363_, _048364_, _048365_, _048366_, _048367_, _048368_, _048369_, _048370_, _048371_, _048372_, _048373_, _048374_, _048375_, _048376_, _048377_, _048378_, _048379_, _048380_, _048381_, _048382_, _048383_, _048384_, _048385_, _048386_, _048387_, _048388_, _048389_, _048390_, _048391_, _048392_, _048393_, _048394_, _048395_, _048396_, _048397_, _048398_, _048399_, _048400_, _048401_, _048402_, _048403_, _048404_, _048405_, _048406_, _048407_, _048408_, _048409_, _048410_, _048411_, _048412_, _048413_, _048414_, _048415_, _048416_, _048417_, _048418_, _048419_, _048420_, _048421_, _048422_, _048423_, _048424_, _048425_, _048426_, _048427_, _048428_, _048429_, _048430_, _048431_, _048432_, _048433_, _048434_, _048435_, _048436_, _048437_, _048438_, _048439_, _048440_, _048441_, _048442_, _048443_, _048444_, _048445_, _048446_, _048447_, _048448_, _048449_, _048450_, _048451_, _048452_, _048453_, _048454_, _048455_, _048456_, _048457_, _048458_, _048459_, _048460_, _048461_, _048462_, _048463_, _048464_, _048465_, _048466_, _048467_, _048468_, _048469_, _048470_, _048471_, _048472_, _048473_, _048474_, _048475_, _048476_, _048477_, _048478_, _048479_, _048480_, _048481_, _048482_, _048483_, _048484_, _048485_, _048486_, _048487_, _048488_, _048489_, _048490_, _048491_, _048492_, _048493_, _048494_, _048495_, _048496_, _048497_, _048498_, _048499_, _048500_, _048501_, _048502_, _048503_, _048504_, _048505_, _048506_, _048507_, _048508_, _048509_, _048510_, _048511_, _048512_, _048513_, _048514_, _048515_, _048516_, _048517_, _048518_, _048519_, _048520_, _048521_, _048522_, _048523_, _048524_, _048525_, _048526_, _048527_, _048528_, _048529_, _048530_, _048531_, _048532_, _048533_, _048534_, _048535_, _048536_, _048537_, _048538_, _048539_, _048540_, _048541_, _048542_, _048543_, _048544_, _048545_, _048546_, _048547_, _048548_, _048549_, _048550_, _048551_, _048552_, _048553_, _048554_, _048555_, _048556_, _048557_, _048558_, _048559_, _048560_, _048561_, _048562_, _048563_, _048564_, _048565_, _048566_, _048567_, _048568_, _048569_, _048570_, _048571_, _048572_, _048573_, _048574_, _048575_, _048576_, _048577_, _048578_, _048579_, _048580_, _048581_, _048582_, _048583_, _048584_, _048585_, _048586_, _048587_, _048588_, _048589_, _048590_, _048591_, _048592_, _048593_, _048594_, _048595_, _048596_, _048597_, _048598_, _048599_, _048600_, _048601_, _048602_, _048603_, _048604_, _048605_, _048606_, _048607_, _048608_, _048609_, _048610_, _048611_, _048612_, _048613_, _048614_, _048615_, _048616_, _048617_, _048618_, _048619_, _048620_, _048621_, _048622_, _048623_, _048624_, _048625_, _048626_, _048627_, _048628_, _048629_, _048630_, _048631_, _048632_, _048633_, _048634_, _048635_, _048636_, _048637_, _048638_, _048639_, _048640_, _048641_, _048642_, _048643_, _048644_, _048645_, _048646_, _048647_, _048648_, _048649_, _048650_, _048651_, _048652_, _048653_, _048654_, _048655_, _048656_, _048657_, _048658_, _048659_, _048660_, _048661_, _048662_, _048663_, _048664_, _048665_, _048666_, _048667_, _048668_, _048669_, _048670_, _048671_, _048672_, _048673_, _048674_, _048675_, _048676_, _048677_, _048678_, _048679_, _048680_, _048681_, _048682_, _048683_, _048684_, _048685_, _048686_, _048687_, _048688_, _048689_, _048690_, _048691_, _048692_, _048693_, _048694_, _048695_, _048696_, _048697_, _048698_, _048699_, _048700_, _048701_, _048702_, _048703_, _048704_, _048705_, _048706_, _048707_, _048708_, _048709_, _048710_, _048711_, _048712_, _048713_, _048714_, _048715_, _048716_, _048717_, _048718_, _048719_, _048720_, _048721_, _048722_, _048723_, _048724_, _048725_, _048726_, _048727_, _048728_, _048729_, _048730_, _048731_, _048732_, _048733_, _048734_, _048735_, _048736_, _048737_, _048738_, _048739_, _048740_, _048741_, _048742_, _048743_, _048744_, _048745_, _048746_, _048747_, _048748_, _048749_, _048750_, _048751_, _048752_, _048753_, _048754_, _048755_, _048756_, _048757_, _048758_, _048759_, _048760_, _048761_, _048762_, _048763_, _048764_, _048765_, _048766_, _048767_, _048768_, _048769_, _048770_, _048771_, _048772_, _048773_, _048774_, _048775_, _048776_, _048777_, _048778_, _048779_, _048780_, _048781_, _048782_, _048783_, _048784_, _048785_, _048786_, _048787_, _048788_, _048789_, _048790_, _048791_, _048792_, _048793_, _048794_, _048795_, _048796_, _048797_, _048798_, _048799_, _048800_, _048801_, _048802_, _048803_, _048804_, _048805_, _048806_, _048807_, _048808_, _048809_, _048810_, _048811_, _048812_, _048813_, _048814_, _048815_, _048816_, _048817_, _048818_, _048819_, _048820_, _048821_, _048822_, _048823_, _048824_, _048825_, _048826_, _048827_, _048828_, _048829_, _048830_, _048831_, _048832_, _048833_, _048834_, _048835_, _048836_, _048837_, _048838_, _048839_, _048840_, _048841_, _048842_, _048843_, _048844_, _048845_, _048846_, _048847_, _048848_, _048849_, _048850_, _048851_, _048852_, _048853_, _048854_, _048855_, _048856_, _048857_, _048858_, _048859_, _048860_, _048861_, _048862_, _048863_, _048864_, _048865_, _048866_, _048867_, _048868_, _048869_, _048870_, _048871_, _048872_, _048873_, _048874_, _048875_, _048876_, _048877_, _048878_, _048879_, _048880_, _048881_, _048882_, _048883_, _048884_, _048885_, _048886_, _048887_, _048888_, _048889_, _048890_, _048891_, _048892_, _048893_, _048894_, _048895_, _048896_, _048897_, _048898_, _048899_, _048900_, _048901_, _048902_, _048903_, _048904_, _048905_, _048906_, _048907_, _048908_, _048909_, _048910_, _048911_, _048912_, _048913_, _048914_, _048915_, _048916_, _048917_, _048918_, _048919_, _048920_, _048921_, _048922_, _048923_, _048924_, _048925_, _048926_, _048927_, _048928_, _048929_, _048930_, _048931_, _048932_, _048933_, _048934_, _048935_, _048936_, _048937_, _048938_, _048939_, _048940_, _048941_, _048942_, _048943_, _048944_, _048945_, _048946_, _048947_, _048948_, _048949_, _048950_, _048951_, _048952_, _048953_, _048954_, _048955_, _048956_, _048957_, _048958_, _048959_, _048960_, _048961_, _048962_, _048963_, _048964_, _048965_, _048966_, _048967_, _048968_, _048969_, _048970_, _048971_, _048972_, _048973_, _048974_, _048975_, _048976_, _048977_, _048978_, _048979_, _048980_, _048981_, _048982_, _048983_, _048984_, _048985_, _048986_, _048987_, _048988_, _048989_, _048990_, _048991_, _048992_, _048993_, _048994_, _048995_, _048996_, _048997_, _048998_, _048999_, _049000_, _049001_, _049002_, _049003_, _049004_, _049005_, _049006_, _049007_, _049008_, _049009_, _049010_, _049011_, _049012_, _049013_, _049014_, _049015_, _049016_, _049017_, _049018_, _049019_, _049020_, _049021_, _049022_, _049023_, _049024_, _049025_, _049026_, _049027_, _049028_, _049029_, _049030_, _049031_, _049032_, _049033_, _049034_, _049035_, _049036_, _049037_, _049038_, _049039_, _049040_, _049041_, _049042_, _049043_, _049044_, _049045_, _049046_, _049047_, _049048_, _049049_, _049050_, _049051_, _049052_, _049053_, _049054_, _049055_, _049056_, _049057_, _049058_, _049059_, _049060_, _049061_, _049062_, _049063_, _049064_, _049065_, _049066_, _049067_, _049068_, _049069_, _049070_, _049071_, _049072_, _049073_, _049074_, _049075_, _049076_, _049077_, _049078_, _049079_, _049080_, _049081_, _049082_, _049083_, _049084_, _049085_, _049086_, _049087_, _049088_, _049089_, _049090_, _049091_, _049092_, _049093_, _049094_, _049095_, _049096_, _049097_, _049098_, _049099_, _049100_, _049101_, _049102_, _049103_, _049104_, _049105_, _049106_, _049107_, _049108_, _049109_, _049110_, _049111_, _049112_, _049113_, _049114_, _049115_, _049116_, _049117_, _049118_, _049119_, _049120_, _049121_, _049122_, _049123_, _049124_, _049125_, _049126_, _049127_, _049128_, _049129_, _049130_, _049131_, _049132_, _049133_, _049134_, _049135_, _049136_, _049137_, _049138_, _049139_, _049140_, _049141_, _049142_, _049143_, _049144_, _049145_, _049146_, _049147_, _049148_, _049149_, _049150_, _049151_, _049152_, _049153_, _049154_, _049155_, _049156_, _049157_, _049158_, _049159_, _049160_, _049161_, _049162_, _049163_, _049164_, _049165_, _049166_, _049167_, _049168_, _049169_, _049170_, _049171_, _049172_, _049173_, _049174_, _049175_, _049176_, _049177_, _049178_, _049179_, _049180_, _049181_, _049182_, _049183_, _049184_, _049185_, _049186_, _049187_, _049188_, _049189_, _049190_, _049191_, _049192_, _049193_, _049194_, _049195_, _049196_, _049197_, _049198_, _049199_, _049200_, _049201_, _049202_, _049203_, _049204_, _049205_, _049206_, _049207_, _049208_, _049209_, _049210_, _049211_, _049212_, _049213_, _049214_, _049215_, _049216_, _049217_, _049218_, _049219_, _049220_, _049221_, _049222_, _049223_, _049224_, _049225_, _049226_, _049227_, _049228_, _049229_, _049230_, _049231_, _049232_, _049233_, _049234_, _049235_, _049236_, _049237_, _049238_, _049239_, _049240_, _049241_, _049242_, _049243_, _049244_, _049245_, _049246_, _049247_, _049248_, _049249_, _049250_, _049251_, _049252_, _049253_, _049254_, _049255_, _049256_, _049257_, _049258_, _049259_, _049260_, _049261_, _049262_, _049263_, _049264_, _049265_, _049266_, _049267_, _049268_, _049269_, _049270_, _049271_, _049272_, _049273_, _049274_, _049275_, _049276_, _049277_, _049278_, _049279_, _049280_, _049281_, _049282_, _049283_, _049284_, _049285_, _049286_, _049287_, _049288_, _049289_, _049290_, _049291_, _049292_, _049293_, _049294_, _049295_, _049296_, _049297_, _049298_, _049299_, _049300_, _049301_, _049302_, _049303_, _049304_, _049305_, _049306_, _049307_, _049308_, _049309_, _049310_, _049311_, _049312_, _049313_, _049314_, _049315_, _049316_, _049317_, _049318_, _049319_, _049320_, _049321_, _049322_, _049323_, _049324_, _049325_, _049326_, _049327_, _049328_, _049329_, _049330_, _049331_, _049332_, _049333_, _049334_, _049335_, _049336_, _049337_, _049338_, _049339_, _049340_, _049341_, _049342_, _049343_, _049344_, _049345_, _049346_, _049347_, _049348_, _049349_, _049350_, _049351_, _049352_, _049353_, _049354_, _049355_, _049356_, _049357_, _049358_, _049359_, _049360_, _049361_, _049362_, _049363_, _049364_, _049365_, _049366_, _049367_, _049368_, _049369_, _049370_, _049371_, _049372_, _049373_, _049374_, _049375_, _049376_, _049377_, _049378_, _049379_, _049380_, _049381_, _049382_, _049383_, _049384_, _049385_, _049386_, _049387_, _049388_, _049389_, _049390_, _049391_, _049392_, _049393_, _049394_, _049395_, _049396_, _049397_, _049398_, _049399_, _049400_, _049401_, _049402_, _049403_, _049404_, _049405_, _049406_, _049407_, _049408_, _049409_, _049410_, _049411_, _049412_, _049413_, _049414_, _049415_, _049416_, _049417_, _049418_, _049419_, _049420_, _049421_, _049422_, _049423_, _049424_, _049425_, _049426_, _049427_, _049428_, _049429_, _049430_, _049431_, _049432_, _049433_, _049434_, _049435_, _049436_, _049437_, _049438_, _049439_, _049440_, _049441_, _049442_, _049443_, _049444_, _049445_, _049446_, _049447_, _049448_, _049449_, _049450_, _049451_, _049452_, _049453_, _049454_, _049455_, _049456_, _049457_, _049458_, _049459_, _049460_, _049461_, _049462_, _049463_, _049464_, _049465_, _049466_, _049467_, _049468_, _049469_, _049470_, _049471_, _049472_, _049473_, _049474_, _049475_, _049476_, _049477_, _049478_, _049479_, _049480_, _049481_, _049482_, _049483_, _049484_, _049485_, _049486_, _049487_, _049488_, _049489_, _049490_, _049491_, _049492_, _049493_, _049494_, _049495_, _049496_, _049497_, _049498_, _049499_, _049500_, _049501_, _049502_, _049503_, _049504_, _049505_, _049506_, _049507_, _049508_, _049509_, _049510_, _049511_, _049512_, _049513_, _049514_, _049515_, _049516_, _049517_, _049518_, _049519_, _049520_, _049521_, _049522_, _049523_, _049524_, _049525_, _049526_, _049527_, _049528_, _049529_, _049530_, _049531_, _049532_, _049533_, _049534_, _049535_, _049536_, _049537_, _049538_, _049539_, _049540_, _049541_, _049542_, _049543_, _049544_, _049545_, _049546_, _049547_, _049548_, _049549_, _049550_, _049551_, _049552_, _049553_, _049554_, _049555_, _049556_, _049557_, _049558_, _049559_, _049560_, _049561_, _049562_, _049563_, _049564_, _049565_, _049566_, _049567_, _049568_, _049569_, _049570_, _049571_, _049572_, _049573_, _049574_, _049575_, _049576_, _049577_, _049578_, _049579_, _049580_, _049581_, _049582_, _049583_, _049584_, _049585_, _049586_, _049587_, _049588_, _049589_, _049590_, _049591_, _049592_, _049593_, _049594_, _049595_, _049596_, _049597_, _049598_, _049599_, _049600_, _049601_, _049602_, _049603_, _049604_, _049605_, _049606_, _049607_, _049608_, _049609_, _049610_, _049611_, _049612_, _049613_, _049614_, _049615_, _049616_, _049617_, _049618_, _049619_, _049620_, _049621_, _049622_, _049623_, _049624_, _049625_, _049626_, _049627_, _049628_, _049629_, _049630_, _049631_, _049632_, _049633_, _049634_, _049635_, _049636_, _049637_, _049638_, _049639_, _049640_, _049641_, _049642_, _049643_, _049644_, _049645_, _049646_, _049647_, _049648_, _049649_, _049650_, _049651_, _049652_, _049653_, _049654_, _049655_, _049656_, _049657_, _049658_, _049659_, _049660_, _049661_, _049662_, _049663_, _049664_, _049665_, _049666_, _049667_, _049668_, _049669_, _049670_, _049671_, _049672_, _049673_, _049674_, _049675_, _049676_, _049677_, _049678_, _049679_, _049680_, _049681_, _049682_, _049683_, _049684_, _049685_, _049686_, _049687_, _049688_, _049689_, _049690_, _049691_, _049692_, _049693_, _049694_, _049695_, _049696_, _049697_, _049698_, _049699_, _049700_, _049701_, _049702_, _049703_, _049704_, _049705_, _049706_, _049707_, _049708_, _049709_, _049710_, _049711_, _049712_, _049713_, _049714_, _049715_, _049716_, _049717_, _049718_, _049719_, _049720_, _049721_, _049722_, _049723_, _049724_, _049725_, _049726_, _049727_, _049728_, _049729_, _049730_, _049731_, _049732_, _049733_, _049734_, _049735_, _049736_, _049737_, _049738_, _049739_, _049740_, _049741_, _049742_, _049743_, _049744_, _049745_, _049746_, _049747_, _049748_, _049749_, _049750_, _049751_, _049752_, _049753_, _049754_, _049755_, _049756_, _049757_, _049758_, _049759_, _049760_, _049761_, _049762_, _049763_, _049764_, _049765_, _049766_, _049767_, _049768_, _049769_, _049770_, _049771_, _049772_, _049773_, _049774_, _049775_, _049776_, _049777_, _049778_, _049779_, _049780_, _049781_, _049782_, _049783_, _049784_, _049785_, _049786_, _049787_, _049788_, _049789_, _049790_, _049791_, _049792_, _049793_, _049794_, _049795_, _049796_, _049797_, _049798_, _049799_, _049800_, _049801_, _049802_, _049803_, _049804_, _049805_, _049806_, _049807_, _049808_, _049809_, _049810_, _049811_, _049812_, _049813_, _049814_, _049815_, _049816_, _049817_, _049818_, _049819_, _049820_, _049821_, _049822_, _049823_, _049824_, _049825_, _049826_, _049827_, _049828_, _049829_, _049830_, _049831_, _049832_, _049833_, _049834_, _049835_, _049836_, _049837_, _049838_, _049839_, _049840_, _049841_, _049842_, _049843_, _049844_, _049845_, _049846_, _049847_, _049848_, _049849_, _049850_, _049851_, _049852_, _049853_, _049854_, _049855_, _049856_, _049857_, _049858_, _049859_, _049860_, _049861_, _049862_, _049863_, _049864_, _049865_, _049866_, _049867_, _049868_, _049869_, _049870_, _049871_, _049872_, _049873_, _049874_, _049875_, _049876_, _049877_, _049878_, _049879_, _049880_, _049881_, _049882_, _049883_, _049884_, _049885_, _049886_, _049887_, _049888_, _049889_, _049890_, _049891_, _049892_, _049893_, _049894_, _049895_, _049896_, _049897_, _049898_, _049899_, _049900_, _049901_, _049902_, _049903_, _049904_, _049905_, _049906_, _049907_, _049908_, _049909_, _049910_, _049911_, _049912_, _049913_, _049914_, _049915_, _049916_, _049917_, _049918_, _049919_, _049920_, _049921_, _049922_, _049923_, _049924_, _049925_, _049926_, _049927_, _049928_, _049929_, _049930_, _049931_, _049932_, _049933_, _049934_, _049935_, _049936_, _049937_, _049938_, _049939_, _049940_, _049941_, _049942_, _049943_, _049944_, _049945_, _049946_, _049947_, _049948_, _049949_, _049950_, _049951_, _049952_, _049953_, _049954_, _049955_, _049956_, _049957_, _049958_, _049959_, _049960_, _049961_, _049962_, _049963_, _049964_, _049965_, _049966_, _049967_, _049968_, _049969_, _049970_, _049971_, _049972_, _049973_, _049974_, _049975_, _049976_, _049977_, _049978_, _049979_, _049980_, _049981_, _049982_, _049983_, _049984_, _049985_, _049986_, _049987_, _049988_, _049989_, _049990_, _049991_, _049992_, _049993_, _049994_, _049995_, _049996_, _049997_, _049998_, _049999_, _050000_, _050001_, _050002_, _050003_, _050004_, _050005_, _050006_, _050007_, _050008_, _050009_, _050010_, _050011_, _050012_, _050013_, _050014_, _050015_, _050016_, _050017_, _050018_, _050019_, _050020_, _050021_, _050022_, _050023_, _050024_, _050025_, _050026_, _050027_, _050028_, _050029_, _050030_, _050031_, _050032_, _050033_, _050034_, _050035_, _050036_, _050037_, _050038_, _050039_, _050040_, _050041_, _050042_, _050043_, _050044_, _050045_, _050046_, _050047_, _050048_, _050049_, _050050_, _050051_, _050052_, _050053_, _050054_, _050055_, _050056_, _050057_, _050058_, _050059_, _050060_, _050061_, _050062_, _050063_, _050064_, _050065_, _050066_, _050067_, _050068_, _050069_, _050070_, _050071_, _050072_, _050073_, _050074_, _050075_, _050076_, _050077_, _050078_, _050079_, _050080_, _050081_, _050082_, _050083_, _050084_, _050085_, _050086_, _050087_, _050088_, _050089_, _050090_, _050091_, _050092_, _050093_, _050094_, _050095_, _050096_, _050097_, _050098_, _050099_, _050100_, _050101_, _050102_, _050103_, _050104_, _050105_, _050106_, _050107_, _050108_, _050109_, _050110_, _050111_, _050112_, _050113_, _050114_, _050115_, _050116_, _050117_, _050118_, _050119_, _050120_, _050121_, _050122_, _050123_, _050124_, _050125_, _050126_, _050127_, _050128_, _050129_, _050130_, _050131_, _050132_, _050133_, _050134_, _050135_, _050136_, _050137_, _050138_, _050139_, _050140_, _050141_, _050142_, _050143_, _050144_, _050145_, _050146_, _050147_, _050148_, _050149_, _050150_, _050151_, _050152_, _050153_, _050154_, _050155_, _050156_, _050157_, _050158_, _050159_, _050160_, _050161_, _050162_, _050163_, _050164_, _050165_, _050166_, _050167_, _050168_, _050169_, _050170_, _050171_, _050172_, _050173_, _050174_, _050175_, _050176_, _050177_, _050178_, _050179_, _050180_, _050181_, _050182_, _050183_, _050184_, _050185_, _050186_, _050187_, _050188_, _050189_, _050190_, _050191_, _050192_, _050193_, _050194_, _050195_, _050196_, _050197_, _050198_, _050199_, _050200_, _050201_, _050202_, _050203_, _050204_, _050205_, _050206_, _050207_, _050208_, _050209_, _050210_, _050211_, _050212_, _050213_, _050214_, _050215_, _050216_, _050217_, _050218_, _050219_, _050220_, _050221_, _050222_, _050223_, _050224_, _050225_, _050226_, _050227_, _050228_, _050229_, _050230_, _050231_, _050232_, _050233_, _050234_, _050235_, _050236_, _050237_, _050238_, _050239_, _050240_, _050241_, _050242_, _050243_, _050244_, _050245_, _050246_, _050247_, _050248_, _050249_, _050250_, _050251_, _050252_, _050253_, _050254_, _050255_, _050256_, _050257_, _050258_, _050259_, _050260_, _050261_, _050262_, _050263_, _050264_, _050265_, _050266_, _050267_, _050268_, _050269_, _050270_, _050271_, _050272_, _050273_, _050274_, _050275_, _050276_, _050277_, _050278_, _050279_, _050280_, _050281_, _050282_, _050283_, _050284_, _050285_, _050286_, _050287_, _050288_, _050289_, _050290_, _050291_, _050292_, _050293_, _050294_, _050295_, _050296_, _050297_, _050298_, _050299_, _050300_, _050301_, _050302_, _050303_, _050304_, _050305_, _050306_, _050307_, _050308_, _050309_, _050310_, _050311_, _050312_, _050313_, _050314_, _050315_, _050316_, _050317_, _050318_, _050319_, _050320_, _050321_, _050322_, _050323_, _050324_, _050325_, _050326_, _050327_, _050328_, _050329_, _050330_, _050331_, _050332_, _050333_, _050334_, _050335_, _050336_, _050337_, _050338_, _050339_, _050340_, _050341_, _050342_, _050343_, _050344_, _050345_, _050346_, _050347_, _050348_, _050349_, _050350_, _050351_, _050352_, _050353_, _050354_, _050355_, _050356_, _050357_, _050358_, _050359_, _050360_, _050361_, _050362_, _050363_, _050364_, _050365_, _050366_, _050367_, _050368_, _050369_, _050370_, _050371_, _050372_, _050373_, _050374_, _050375_, _050376_, _050377_, _050378_, _050379_, _050380_, _050381_, _050382_, _050383_, _050384_, _050385_, _050386_, _050387_, _050388_, _050389_, _050390_, _050391_, _050392_, _050393_, _050394_, _050395_, _050396_, _050397_, _050398_, _050399_, _050400_, _050401_, _050402_, _050403_, _050404_, _050405_, _050406_, _050407_, _050408_, _050409_, _050410_, _050411_, _050412_, _050413_, _050414_, _050415_, _050416_, _050417_, _050418_, _050419_, _050420_, _050421_, _050422_, _050423_, _050424_, _050425_, _050426_, _050427_, _050428_, _050429_, _050430_, _050431_, _050432_, _050433_, _050434_, _050435_, _050436_, _050437_, _050438_, _050439_, _050440_, _050441_, _050442_, _050443_, _050444_, _050445_, _050446_, _050447_, _050448_, _050449_, _050450_, _050451_, _050452_, _050453_, _050454_, _050455_, _050456_, _050457_, _050458_, _050459_, _050460_, _050461_, _050462_, _050463_, _050464_, _050465_, _050466_, _050467_, _050468_, _050469_, _050470_, _050471_, _050472_, _050473_, _050474_, _050475_, _050476_, _050477_, _050478_, _050479_, _050480_, _050481_, _050482_, _050483_, _050484_, _050485_, _050486_, _050487_, _050488_, _050489_, _050490_, _050491_, _050492_, _050493_, _050494_, _050495_, _050496_, _050497_, _050498_, _050499_, _050500_, _050501_, _050502_, _050503_, _050504_, _050505_, _050506_, _050507_, _050508_, _050509_, _050510_, _050511_, _050512_, _050513_, _050514_, _050515_, _050516_, _050517_, _050518_, _050519_, _050520_, _050521_, _050522_, _050523_, _050524_, _050525_, _050526_, _050527_, _050528_, _050529_, _050530_, _050531_, _050532_, _050533_, _050534_, _050535_, _050536_, _050537_, _050538_, _050539_, _050540_, _050541_, _050542_, _050543_, _050544_, _050545_, _050546_, _050547_, _050548_, _050549_, _050550_, _050551_, _050552_, _050553_, _050554_, _050555_, _050556_, _050557_, _050558_, _050559_, _050560_, _050561_, _050562_, _050563_, _050564_, _050565_, _050566_, _050567_, _050568_, _050569_, _050570_, _050571_, _050572_, _050573_, _050574_, _050575_, _050576_, _050577_, _050578_, _050579_, _050580_, _050581_, _050582_, _050583_, _050584_, _050585_, _050586_, _050587_, _050588_, _050589_, _050590_, _050591_, _050592_, _050593_, _050594_, _050595_, _050596_, _050597_, _050598_, _050599_, _050600_, _050601_, _050602_, _050603_, _050604_, _050605_, _050606_, _050607_, _050608_, _050609_, _050610_, _050611_, _050612_, _050613_, _050614_, _050615_, _050616_, _050617_, _050618_, _050619_, _050620_, _050621_, _050622_, _050623_, _050624_, _050625_, _050626_, _050627_, _050628_, _050629_, _050630_, _050631_, _050632_, _050633_, _050634_, _050635_, _050636_, _050637_, _050638_, _050639_, _050640_, _050641_, _050642_, _050643_, _050644_, _050645_, _050646_, _050647_, _050648_, _050649_, _050650_, _050651_, _050652_, _050653_, _050654_, _050655_, _050656_, _050657_, _050658_, _050659_, _050660_, _050661_, _050662_, _050663_, _050664_, _050665_, _050666_, _050667_, _050668_, _050669_, _050670_, _050671_, _050672_, _050673_, _050674_, _050675_, _050676_, _050677_, _050678_, _050679_, _050680_, _050681_, _050682_, _050683_, _050684_, _050685_, _050686_, _050687_, _050688_, _050689_, _050690_, _050691_, _050692_, _050693_, _050694_, _050695_, _050696_, _050697_, _050698_, _050699_, _050700_, _050701_, _050702_, _050703_, _050704_, _050705_, _050706_, _050707_, _050708_, _050709_, _050710_, _050711_, _050712_, _050713_, _050714_, _050715_, _050716_, _050717_, _050718_, _050719_, _050720_, _050721_, _050722_, _050723_, _050724_, _050725_, _050726_, _050727_, _050728_, _050729_, _050730_, _050731_, _050732_, _050733_, _050734_, _050735_, _050736_, _050737_, _050738_, _050739_, _050740_, _050741_, _050742_, _050743_, _050744_, _050745_, _050746_, _050747_, _050748_, _050749_, _050750_, _050751_, _050752_, _050753_, _050754_, _050755_, _050756_, _050757_, _050758_, _050759_, _050760_, _050761_, _050762_, _050763_, _050764_, _050765_, _050766_, _050767_, _050768_, _050769_, _050770_, _050771_, _050772_, _050773_, _050774_, _050775_, _050776_, _050777_, _050778_, _050779_, _050780_, _050781_, _050782_, _050783_, _050784_, _050785_, _050786_, _050787_, _050788_, _050789_, _050790_, _050791_, _050792_, _050793_, _050794_, _050795_, _050796_, _050797_, _050798_, _050799_, _050800_, _050801_, _050802_, _050803_, _050804_, _050805_, _050806_, _050807_, _050808_, _050809_, _050810_, _050811_, _050812_, _050813_, _050814_, _050815_, _050816_, _050817_, _050818_, _050819_, _050820_, _050821_, _050822_, _050823_, _050824_, _050825_, _050826_, _050827_, _050828_, _050829_, _050830_, _050831_, _050832_, _050833_, _050834_, _050835_, _050836_, _050837_, _050838_, _050839_, _050840_, _050841_, _050842_, _050843_, _050844_, _050845_, _050846_, _050847_, _050848_, _050849_, _050850_, _050851_, _050852_, _050853_, _050854_, _050855_, _050856_, _050857_, _050858_, _050859_, _050860_, _050861_, _050862_, _050863_, _050864_, _050865_, _050866_, _050867_, _050868_, _050869_, _050870_, _050871_, _050872_, _050873_, _050874_, _050875_, _050876_, _050877_, _050878_, _050879_, _050880_, _050881_, _050882_, _050883_, _050884_, _050885_, _050886_, _050887_, _050888_, _050889_, _050890_, _050891_, _050892_, _050893_, _050894_, _050895_, _050896_, _050897_, _050898_, _050899_, _050900_, _050901_, _050902_, _050903_, _050904_, _050905_, _050906_, _050907_, _050908_, _050909_, _050910_, _050911_, _050912_, _050913_, _050914_, _050915_, _050916_, _050917_, _050918_, _050919_, _050920_, _050921_, _050922_, _050923_, _050924_, _050925_, _050926_, _050927_, _050928_, _050929_, _050930_, _050931_, _050932_, _050933_, _050934_, _050935_, _050936_, _050937_, _050938_, _050939_, _050940_, _050941_, _050942_, _050943_, _050944_, _050945_, _050946_, _050947_, _050948_, _050949_, _050950_, _050951_, _050952_, _050953_, _050954_, _050955_, _050956_, _050957_, _050958_, _050959_, _050960_, _050961_, _050962_, _050963_, _050964_, _050965_, _050966_, _050967_, _050968_, _050969_, _050970_, _050971_, _050972_, _050973_, _050974_, _050975_, _050976_, _050977_, _050978_, _050979_, _050980_, _050981_, _050982_, _050983_, _050984_, _050985_, _050986_, _050987_, _050988_, _050989_, _050990_, _050991_, _050992_, _050993_, _050994_, _050995_, _050996_, _050997_, _050998_, _050999_, _051000_, _051001_, _051002_, _051003_, _051004_, _051005_, _051006_, _051007_, _051008_, _051009_, _051010_, _051011_, _051012_, _051013_, _051014_, _051015_, _051016_, _051017_, _051018_, _051019_, _051020_, _051021_, _051022_, _051023_, _051024_, _051025_, _051026_, _051027_, _051028_, _051029_, _051030_, _051031_, _051032_, _051033_, _051034_, _051035_, _051036_, _051037_, _051038_, _051039_, _051040_, _051041_, _051042_, _051043_, _051044_, _051045_, _051046_, _051047_, _051048_, _051049_, _051050_, _051051_, _051052_, _051053_, _051054_, _051055_, _051056_, _051057_, _051058_, _051059_, _051060_, _051061_, _051062_, _051063_, _051064_, _051065_, _051066_, _051067_, _051068_, _051069_, _051070_, _051071_, _051072_, _051073_, _051074_, _051075_, _051076_, _051077_, _051078_, _051079_, _051080_, _051081_, _051082_, _051083_, _051084_, _051085_, _051086_, _051087_, _051088_, _051089_, _051090_, _051091_, _051092_, _051093_, _051094_, _051095_, _051096_, _051097_, _051098_, _051099_, _051100_, _051101_, _051102_, _051103_, _051104_, _051105_, _051106_, _051107_, _051108_, _051109_, _051110_, _051111_, _051112_, _051113_, _051114_, _051115_, _051116_, _051117_, _051118_, _051119_, _051120_, _051121_, _051122_, _051123_, _051124_, _051125_, _051126_, _051127_, _051128_, _051129_, _051130_, _051131_, _051132_, _051133_, _051134_, _051135_, _051136_, _051137_, _051138_, _051139_, _051140_, _051141_, _051142_, _051143_, _051144_, _051145_, _051146_, _051147_, _051148_, _051149_, _051150_, _051151_, _051152_, _051153_, _051154_, _051155_, _051156_, _051157_, _051158_, _051159_, _051160_, _051161_, _051162_, _051163_, _051164_, _051165_, _051166_, _051167_, _051168_, _051169_, _051170_, _051171_, _051172_, _051173_, _051174_, _051175_, _051176_, _051177_, _051178_, _051179_, _051180_, _051181_, _051182_, _051183_, _051184_, _051185_, _051186_, _051187_, _051188_, _051189_, _051190_, _051191_, _051192_, _051193_, _051194_, _051195_, _051196_, _051197_, _051198_, _051199_, _051200_, _051201_, _051202_, _051203_, _051204_, _051205_, _051206_, _051207_, _051208_, _051209_, _051210_, _051211_, _051212_, _051213_, _051214_, _051215_, _051216_, _051217_, _051218_, _051219_, _051220_, _051221_, _051222_, _051223_, _051224_, _051225_, _051226_, _051227_, _051228_, _051229_, _051230_, _051231_, _051232_, _051233_, _051234_, _051235_, _051236_, _051237_, _051238_, _051239_, _051240_, _051241_, _051242_, _051243_, _051244_, _051245_, _051246_, _051247_, _051248_, _051249_, _051250_, _051251_, _051252_, _051253_, _051254_, _051255_, _051256_, _051257_, _051258_, _051259_, _051260_, _051261_, _051262_, _051263_, _051264_, _051265_, _051266_, _051267_, _051268_, _051269_, _051270_, _051271_, _051272_, _051273_, _051274_, _051275_, _051276_, _051277_, _051278_, _051279_, _051280_, _051281_, _051282_, _051283_, _051284_, _051285_, _051286_, _051287_, _051288_, _051289_, _051290_, _051291_, _051292_, _051293_, _051294_, _051295_, _051296_, _051297_, _051298_, _051299_, _051300_, _051301_, _051302_, _051303_, _051304_, _051305_, _051306_, _051307_, _051308_, _051309_, _051310_, _051311_, _051312_, _051313_, _051314_, _051315_, _051316_, _051317_, _051318_, _051319_, _051320_, _051321_, _051322_, _051323_, _051324_, _051325_, _051326_, _051327_, _051328_, _051329_, _051330_, _051331_, _051332_, _051333_, _051334_, _051335_, _051336_, _051337_, _051338_, _051339_, _051340_, _051341_, _051342_, _051343_, _051344_, _051345_, _051346_, _051347_, _051348_, _051349_, _051350_, _051351_, _051352_, _051353_, _051354_, _051355_, _051356_, _051357_, _051358_, _051359_, _051360_, _051361_, _051362_, _051363_, _051364_, _051365_, _051366_, _051367_, _051368_, _051369_, _051370_, _051371_, _051372_, _051373_, _051374_, _051375_, _051376_, _051377_, _051378_, _051379_, _051380_, _051381_, _051382_, _051383_, _051384_, _051385_, _051386_, _051387_, _051388_, _051389_, _051390_, _051391_, _051392_, _051393_, _051394_, _051395_, _051396_, _051397_, _051398_, _051399_, _051400_, _051401_, _051402_, _051403_, _051404_, _051405_, _051406_, _051407_, _051408_, _051409_, _051410_, _051411_, _051412_, _051413_, _051414_, _051415_, _051416_, _051417_, _051418_, _051419_, _051420_, _051421_, _051422_, _051423_, _051424_, _051425_, _051426_, _051427_, _051428_, _051429_, _051430_, _051431_, _051432_, _051433_, _051434_, _051435_, _051436_, _051437_, _051438_, _051439_, _051440_, _051441_, _051442_, _051443_, _051444_, _051445_, _051446_, _051447_, _051448_, _051449_, _051450_, _051451_, _051452_, _051453_, _051454_, _051455_, _051456_, _051457_, _051458_, _051459_, _051460_, _051461_, _051462_, _051463_, _051464_, _051465_, _051466_, _051467_, _051468_, _051469_, _051470_, _051471_, _051472_, _051473_, _051474_, _051475_, _051476_, _051477_, _051478_, _051479_, _051480_, _051481_, _051482_, _051483_, _051484_, _051485_, _051486_, _051487_, _051488_, _051489_, _051490_, _051491_, _051492_, _051493_, _051494_, _051495_, _051496_, _051497_, _051498_, _051499_, _051500_, _051501_, _051502_, _051503_, _051504_, _051505_, _051506_, _051507_, _051508_, _051509_, _051510_, _051511_, _051512_, _051513_, _051514_, _051515_, _051516_, _051517_, _051518_, _051519_, _051520_, _051521_, _051522_, _051523_, _051524_, _051525_, _051526_, _051527_, _051528_, _051529_, _051530_, _051531_, _051532_, _051533_, _051534_, _051535_, _051536_, _051537_, _051538_, _051539_, _051540_, _051541_, _051542_, _051543_, _051544_, _051545_, _051546_, _051547_, _051548_, _051549_, _051550_, _051551_, _051552_, _051553_, _051554_, _051555_, _051556_, _051557_, _051558_, _051559_, _051560_, _051561_, _051562_, _051563_, _051564_, _051565_, _051566_, _051567_, _051568_, _051569_, _051570_, _051571_, _051572_, _051573_, _051574_, _051575_, _051576_, _051577_, _051578_, _051579_, _051580_, _051581_, _051582_, _051583_, _051584_, _051585_, _051586_, _051587_, _051588_, _051589_, _051590_, _051591_, _051592_, _051593_, _051594_, _051595_, _051596_, _051597_, _051598_, _051599_, _051600_, _051601_, _051602_, _051603_, _051604_, _051605_, _051606_, _051607_, _051608_, _051609_, _051610_, _051611_, _051612_, _051613_, _051614_, _051615_, _051616_, _051617_, _051618_, _051619_, _051620_, _051621_, _051622_, _051623_, _051624_, _051625_, _051626_, _051627_, _051628_, _051629_, _051630_, _051631_, _051632_, _051633_, _051634_, _051635_, _051636_, _051637_, _051638_, _051639_, _051640_, _051641_, _051642_, _051643_, _051644_, _051645_, _051646_, _051647_, _051648_, _051649_, _051650_, _051651_, _051652_, _051653_, _051654_, _051655_, _051656_, _051657_, _051658_, _051659_, _051660_, _051661_, _051662_, _051663_, _051664_, _051665_, _051666_, _051667_, _051668_, _051669_, _051670_, _051671_, _051672_, _051673_, _051674_, _051675_, _051676_, _051677_, _051678_, _051679_, _051680_, _051681_, _051682_, _051683_, _051684_, _051685_, _051686_, _051687_, _051688_, _051689_, _051690_, _051691_, _051692_, _051693_, _051694_, _051695_, _051696_, _051697_, _051698_, _051699_, _051700_, _051701_, _051702_, _051703_, _051704_, _051705_, _051706_, _051707_, _051708_, _051709_, _051710_, _051711_, _051712_, _051713_, _051714_, _051715_, _051716_, _051717_, _051718_, _051719_, _051720_, _051721_, _051722_, _051723_, _051724_, _051725_, _051726_, _051727_, _051728_, _051729_, _051730_, _051731_, _051732_, _051733_, _051734_, _051735_, _051736_, _051737_, _051738_, _051739_, _051740_, _051741_, _051742_, _051743_, _051744_, _051745_, _051746_, _051747_, _051748_, _051749_, _051750_, _051751_, _051752_, _051753_, _051754_, _051755_, _051756_, _051757_, _051758_, _051759_, _051760_, _051761_, _051762_, _051763_, _051764_, _051765_, _051766_, _051767_, _051768_, _051769_, _051770_, _051771_, _051772_, _051773_, _051774_, _051775_, _051776_, _051777_, _051778_, _051779_, _051780_, _051781_, _051782_, _051783_, _051784_, _051785_, _051786_, _051787_, _051788_, _051789_, _051790_, _051791_, _051792_, _051793_, _051794_, _051795_, _051796_, _051797_, _051798_, _051799_, _051800_, _051801_, _051802_, _051803_, _051804_, _051805_, _051806_, _051807_, _051808_, _051809_, _051810_, _051811_, _051812_, _051813_, _051814_, _051815_, _051816_, _051817_, _051818_, _051819_, _051820_, _051821_, _051822_, _051823_, _051824_, _051825_, _051826_, _051827_, _051828_, _051829_, _051830_, _051831_, _051832_, _051833_, _051834_, _051835_, _051836_, _051837_, _051838_, _051839_, _051840_, _051841_, _051842_, _051843_, _051844_, _051845_, _051846_, _051847_, _051848_, _051849_, _051850_, _051851_, _051852_, _051853_, _051854_, _051855_, _051856_, _051857_, _051858_, _051859_, _051860_, _051861_, _051862_, _051863_, _051864_, _051865_, _051866_, _051867_, _051868_, _051869_, _051870_, _051871_, _051872_, _051873_, _051874_, _051875_, _051876_, _051877_, _051878_, _051879_, _051880_, _051881_, _051882_, _051883_, _051884_, _051885_, _051886_, _051887_, _051888_, _051889_, _051890_, _051891_, _051892_, _051893_, _051894_, _051895_, _051896_, _051897_, _051898_, _051899_, _051900_, _051901_, _051902_, _051903_, _051904_, _051905_, _051906_, _051907_, _051908_, _051909_, _051910_, _051911_, _051912_, _051913_, _051914_, _051915_, _051916_, _051917_, _051918_, _051919_, _051920_, _051921_, _051922_, _051923_, _051924_, _051925_, _051926_, _051927_, _051928_, _051929_, _051930_, _051931_, _051932_, _051933_, _051934_, _051935_, _051936_, _051937_, _051938_, _051939_, _051940_, _051941_, _051942_, _051943_, _051944_, _051945_, _051946_, _051947_, _051948_, _051949_, _051950_, _051951_, _051952_, _051953_, _051954_, _051955_, _051956_, _051957_, _051958_, _051959_, _051960_, _051961_, _051962_, _051963_, _051964_, _051965_, _051966_, _051967_, _051968_, _051969_, _051970_, _051971_, _051972_, _051973_, _051974_, _051975_, _051976_, _051977_, _051978_, _051979_, _051980_, _051981_, _051982_, _051983_, _051984_, _051985_, _051986_, _051987_, _051988_, _051989_, _051990_, _051991_, _051992_, _051993_, _051994_, _051995_, _051996_, _051997_, _051998_, _051999_, _052000_, _052001_, _052002_, _052003_, _052004_, _052005_, _052006_, _052007_, _052008_, _052009_, _052010_, _052011_, _052012_, _052013_, _052014_, _052015_, _052016_, _052017_, _052018_, _052019_, _052020_, _052021_, _052022_, _052023_, _052024_, _052025_, _052026_, _052027_, _052028_, _052029_, _052030_, _052031_, _052032_, _052033_, _052034_, _052035_, _052036_, _052037_, _052038_, _052039_, _052040_, _052041_, _052042_, _052043_, _052044_, _052045_, _052046_, _052047_, _052048_, _052049_, _052050_, _052051_, _052052_, _052053_, _052054_, _052055_, _052056_, _052057_, _052058_, _052059_, _052060_, _052061_, _052062_, _052063_, _052064_, _052065_, _052066_, _052067_, _052068_, _052069_, _052070_, _052071_, _052072_, _052073_, _052074_, _052075_, _052076_, _052077_, _052078_, _052079_, _052080_, _052081_, _052082_, _052083_, _052084_, _052085_, _052086_, _052087_, _052088_, _052089_, _052090_, _052091_, _052092_, _052093_, _052094_, _052095_, _052096_, _052097_, _052098_, _052099_, _052100_, _052101_, _052102_, _052103_, _052104_, _052105_, _052106_, _052107_, _052108_, _052109_, _052110_, _052111_, _052112_, _052113_, _052114_, _052115_, _052116_, _052117_, _052118_, _052119_, _052120_, _052121_, _052122_, _052123_, _052124_, _052125_, _052126_, _052127_, _052128_, _052129_, _052130_, _052131_, _052132_, _052133_, _052134_, _052135_, _052136_, _052137_, _052138_, _052139_, _052140_, _052141_, _052142_, _052143_, _052144_, _052145_, _052146_, _052147_, _052148_, _052149_, _052150_, _052151_, _052152_, _052153_, _052154_, _052155_, _052156_, _052157_, _052158_, _052159_, _052160_, _052161_, _052162_, _052163_, _052164_, _052165_, _052166_, _052167_, _052168_, _052169_, _052170_, _052171_, _052172_, _052173_, _052174_, _052175_, _052176_, _052177_, _052178_, _052179_, _052180_, _052181_, _052182_, _052183_, _052184_, _052185_, _052186_, _052187_, _052188_, _052189_, _052190_, _052191_, _052192_, _052193_, _052194_, _052195_, _052196_, _052197_, _052198_, _052199_, _052200_, _052201_, _052202_, _052203_, _052204_, _052205_, _052206_, _052207_, _052208_, _052209_, _052210_, _052211_, _052212_, _052213_, _052214_, _052215_, _052216_, _052217_, _052218_, _052219_, _052220_, _052221_, _052222_, _052223_, _052224_, _052225_, _052226_, _052227_, _052228_, _052229_, _052230_, _052231_, _052232_, _052233_, _052234_, _052235_, _052236_, _052237_, _052238_, _052239_, _052240_, _052241_, _052242_, _052243_, _052244_, _052245_, _052246_, _052247_, _052248_, _052249_, _052250_, _052251_, _052252_, _052253_, _052254_, _052255_, _052256_, _052257_, _052258_, _052259_, _052260_, _052261_, _052262_, _052263_, _052264_, _052265_, _052266_, _052267_, _052268_, _052269_, _052270_, _052271_, _052272_, _052273_, _052274_, _052275_, _052276_, _052277_, _052278_, _052279_, _052280_, _052281_, _052282_, _052283_, _052284_, _052285_, _052286_, _052287_, _052288_, _052289_, _052290_, _052291_, _052292_, _052293_, _052294_, _052295_, _052296_, _052297_, _052298_, _052299_, _052300_, _052301_, _052302_, _052303_, _052304_, _052305_, _052306_, _052307_, _052308_, _052309_, _052310_, _052311_, _052312_, _052313_, _052314_, _052315_, _052316_, _052317_, _052318_, _052319_, _052320_, _052321_, _052322_, _052323_, _052324_, _052325_, _052326_, _052327_, _052328_, _052329_, _052330_, _052331_, _052332_, _052333_, _052334_, _052335_, _052336_, _052337_, _052338_, _052339_, _052340_, _052341_, _052342_, _052343_, _052344_, _052345_, _052346_, _052347_, _052348_, _052349_, _052350_, _052351_, _052352_, _052353_, _052354_, _052355_, _052356_, _052357_, _052358_, _052359_, _052360_, _052361_, _052362_, _052363_, _052364_, _052365_, _052366_, _052367_, _052368_, _052369_, _052370_, _052371_, _052372_, _052373_, _052374_, _052375_, _052376_, _052377_, _052378_, _052379_, _052380_, _052381_, _052382_, _052383_, _052384_, _052385_, _052386_, _052387_, _052388_, _052389_, _052390_, _052391_, _052392_, _052393_, _052394_, _052395_, _052396_, _052397_, _052398_, _052399_, _052400_, _052401_, _052402_, _052403_, _052404_, _052405_, _052406_, _052407_, _052408_, _052409_, _052410_, _052411_, _052412_, _052413_, _052414_, _052415_, _052416_, _052417_, _052418_, _052419_, _052420_, _052421_, _052422_, _052423_, _052424_, _052425_, _052426_, _052427_, _052428_, _052429_, _052430_, _052431_, _052432_, _052433_, _052434_, _052435_, _052436_, _052437_, _052438_, _052439_, _052440_, _052441_, _052442_, _052443_, _052444_, _052445_, _052446_, _052447_, _052448_, _052449_, _052450_, _052451_, _052452_, _052453_, _052454_, _052455_, _052456_, _052457_, _052458_, _052459_, _052460_, _052461_, _052462_, _052463_, _052464_, _052465_, _052466_, _052467_, _052468_, _052469_, _052470_, _052471_, _052472_, _052473_, _052474_, _052475_, _052476_, _052477_, _052478_, _052479_, _052480_, _052481_, _052482_, _052483_, _052484_, _052485_, _052486_, _052487_, _052488_, _052489_, _052490_, _052491_, _052492_, _052493_, _052494_, _052495_, _052496_, _052497_, _052498_, _052499_, _052500_, _052501_, _052502_, _052503_, _052504_, _052505_, _052506_, _052507_, _052508_, _052509_, _052510_, _052511_, _052512_, _052513_, _052514_, _052515_, _052516_, _052517_, _052518_, _052519_, _052520_, _052521_, _052522_, _052523_, _052524_, _052525_, _052526_, _052527_, _052528_, _052529_, _052530_, _052531_, _052532_, _052533_, _052534_, _052535_, _052536_, _052537_, _052538_, _052539_, _052540_, _052541_, _052542_, _052543_, _052544_, _052545_, _052546_, _052547_, _052548_, _052549_, _052550_, _052551_, _052552_, _052553_, _052554_, _052555_, _052556_, _052557_, _052558_, _052559_, _052560_, _052561_, _052562_, _052563_, _052564_, _052565_, _052566_, _052567_, _052568_, _052569_, _052570_, _052571_, _052572_, _052573_, _052574_, _052575_, _052576_, _052577_, _052578_, _052579_, _052580_, _052581_, _052582_, _052583_, _052584_, _052585_, _052586_, _052587_, _052588_, _052589_, _052590_, _052591_, _052592_, _052593_, _052594_, _052595_, _052596_, _052597_, _052598_, _052599_, _052600_, _052601_, _052602_, _052603_, _052604_, _052605_, _052606_, _052607_, _052608_, _052609_, _052610_, _052611_, _052612_, _052613_, _052614_, _052615_, _052616_, _052617_, _052618_, _052619_, _052620_, _052621_, _052622_, _052623_, _052624_, _052625_, _052626_, _052627_, _052628_, _052629_, _052630_, _052631_, _052632_, _052633_, _052634_, _052635_, _052636_, _052637_, _052638_, _052639_, _052640_, _052641_, _052642_, _052643_, _052644_, _052645_, _052646_, _052647_, _052648_, _052649_, _052650_, _052651_, _052652_, _052653_, _052654_, _052655_, _052656_, _052657_, _052658_, _052659_, _052660_, _052661_, _052662_, _052663_, _052664_, _052665_, _052666_, _052667_, _052668_, _052669_, _052670_, _052671_, _052672_, _052673_, _052674_, _052675_, _052676_, _052677_, _052678_, _052679_, _052680_, _052681_, _052682_, _052683_, _052684_, _052685_, _052686_, _052687_, _052688_, _052689_, _052690_, _052691_, _052692_, _052693_, _052694_, _052695_, _052696_, _052697_, _052698_, _052699_, _052700_, _052701_, _052702_, _052703_, _052704_, _052705_, _052706_, _052707_, _052708_, _052709_, _052710_, _052711_, _052712_, _052713_, _052714_, _052715_, _052716_, _052717_, _052718_, _052719_, _052720_, _052721_, _052722_, _052723_, _052724_, _052725_, _052726_, _052727_, _052728_, _052729_, _052730_, _052731_, _052732_, _052733_, _052734_, _052735_, _052736_, _052737_, _052738_, _052739_, _052740_, _052741_, _052742_, _052743_, _052744_, _052745_, _052746_, _052747_, _052748_, _052749_, _052750_, _052751_, _052752_, _052753_, _052754_, _052755_, _052756_, _052757_, _052758_, _052759_, _052760_, _052761_, _052762_, _052763_, _052764_, _052765_, _052766_, _052767_, _052768_, _052769_, _052770_, _052771_, _052772_, _052773_, _052774_, _052775_, _052776_, _052777_, _052778_, _052779_, _052780_, _052781_, _052782_, _052783_, _052784_, _052785_, _052786_, _052787_, _052788_, _052789_, _052790_, _052791_, _052792_, _052793_, _052794_, _052795_, _052796_, _052797_, _052798_, _052799_, _052800_, _052801_, _052802_, _052803_, _052804_, _052805_, _052806_, _052807_, _052808_, _052809_, _052810_, _052811_, _052812_, _052813_, _052814_, _052815_, _052816_, _052817_, _052818_, _052819_, _052820_, _052821_, _052822_, _052823_, _052824_, _052825_, _052826_, _052827_, _052828_, _052829_, _052830_, _052831_, _052832_, _052833_, _052834_, _052835_, _052836_, _052837_, _052838_, _052839_, _052840_, _052841_, _052842_, _052843_, _052844_, _052845_, _052846_, _052847_, _052848_, _052849_, _052850_, _052851_, _052852_, _052853_, _052854_, _052855_, _052856_, _052857_, _052858_, _052859_, _052860_, _052861_, _052862_, _052863_, _052864_, _052865_, _052866_, _052867_, _052868_, _052869_, _052870_, _052871_, _052872_, _052873_, _052874_, _052875_, _052876_, _052877_, _052878_, _052879_, _052880_, _052881_, _052882_, _052883_, _052884_, _052885_, _052886_, _052887_, _052888_, _052889_, _052890_, _052891_, _052892_, _052893_, _052894_, _052895_, _052896_, _052897_, _052898_, _052899_, _052900_, _052901_, _052902_, _052903_, _052904_, _052905_, _052906_, _052907_, _052908_, _052909_, _052910_, _052911_, _052912_, _052913_, _052914_, _052915_, _052916_, _052917_, _052918_, _052919_, _052920_, _052921_, _052922_, _052923_, _052924_, _052925_, _052926_, _052927_, _052928_, _052929_, _052930_, _052931_, _052932_, _052933_, _052934_, _052935_, _052936_, _052937_, _052938_, _052939_, _052940_, _052941_, _052942_, _052943_, _052944_, _052945_, _052946_, _052947_, _052948_, _052949_, _052950_, _052951_, _052952_, _052953_, _052954_, _052955_, _052956_, _052957_, _052958_, _052959_, _052960_, _052961_, _052962_, _052963_, _052964_, _052965_, _052966_, _052967_, _052968_, _052969_, _052970_, _052971_, _052972_, _052973_, _052974_, _052975_, _052976_, _052977_, _052978_, _052979_, _052980_, _052981_, _052982_, _052983_, _052984_, _052985_, _052986_, _052987_, _052988_, _052989_, _052990_, _052991_, _052992_, _052993_, _052994_, _052995_, _052996_, _052997_, _052998_, _052999_, _053000_, _053001_, _053002_, _053003_, _053004_, _053005_, _053006_, _053007_, _053008_, _053009_, _053010_, _053011_, _053012_, _053013_, _053014_, _053015_, _053016_, _053017_, _053018_, _053019_, _053020_, _053021_, _053022_, _053023_, _053024_, _053025_, _053026_, _053027_, _053028_, _053029_, _053030_, _053031_, _053032_, _053033_, _053034_, _053035_, _053036_, _053037_, _053038_, _053039_, _053040_, _053041_, _053042_, _053043_, _053044_, _053045_, _053046_, _053047_, _053048_, _053049_, _053050_, _053051_, _053052_, _053053_, _053054_, _053055_, _053056_, _053057_, _053058_, _053059_, _053060_, _053061_, _053062_, _053063_, _053064_, _053065_, _053066_, _053067_, _053068_, _053069_, _053070_, _053071_, _053072_, _053073_, _053074_, _053075_, _053076_, _053077_, _053078_, _053079_, _053080_, _053081_, _053082_, _053083_, _053084_, _053085_, _053086_, _053087_, _053088_, _053089_, _053090_, _053091_, _053092_, _053093_, _053094_, _053095_, _053096_, _053097_, _053098_, _053099_, _053100_, _053101_, _053102_, _053103_, _053104_, _053105_, _053106_, _053107_, _053108_, _053109_, _053110_, _053111_, _053112_, _053113_, _053114_, _053115_, _053116_, _053117_, _053118_, _053119_, _053120_, _053121_, _053122_, _053123_, _053124_, _053125_, _053126_, _053127_, _053128_, _053129_, _053130_, _053131_, _053132_, _053133_, _053134_, _053135_, _053136_, _053137_, _053138_, _053139_, _053140_, _053141_, _053142_, _053143_, _053144_, _053145_, _053146_, _053147_, _053148_, _053149_, _053150_, _053151_, _053152_, _053153_, _053154_, _053155_, _053156_, _053157_, _053158_, _053159_, _053160_, _053161_, _053162_, _053163_, _053164_, _053165_, _053166_, _053167_, _053168_, _053169_, _053170_, _053171_, _053172_, _053173_, _053174_, _053175_, _053176_, _053177_, _053178_, _053179_, _053180_, _053181_, _053182_, _053183_, _053184_, _053185_, _053186_, _053187_, _053188_, _053189_, _053190_, _053191_, _053192_, _053193_, _053194_, _053195_, _053196_, _053197_, _053198_, _053199_, _053200_, _053201_, _053202_, _053203_, _053204_, _053205_, _053206_, _053207_, _053208_, _053209_, _053210_, _053211_, _053212_, _053213_, _053214_, _053215_, _053216_, _053217_, _053218_, _053219_, _053220_, _053221_, _053222_, _053223_, _053224_, _053225_, _053226_, _053227_, _053228_, _053229_, _053230_, _053231_, _053232_, _053233_, _053234_, _053235_, _053236_, _053237_, _053238_, _053239_, _053240_, _053241_, _053242_, _053243_, _053244_, _053245_, _053246_, _053247_, _053248_, _053249_, _053250_, _053251_, _053252_, _053253_, _053254_, _053255_, _053256_, _053257_, _053258_, _053259_, _053260_, _053261_, _053262_, _053263_, _053264_, _053265_, _053266_, _053267_, _053268_, _053269_, _053270_, _053271_, _053272_, _053273_, _053274_, _053275_, _053276_, _053277_, _053278_, _053279_, _053280_, _053281_, _053282_, _053283_, _053284_, _053285_, _053286_, _053287_, _053288_, _053289_, _053290_, _053291_, _053292_, _053293_, _053294_, _053295_, _053296_, _053297_, _053298_, _053299_, _053300_, _053301_, _053302_, _053303_, _053304_, _053305_, _053306_, _053307_, _053308_, _053309_, _053310_, _053311_, _053312_, _053313_, _053314_, _053315_, _053316_, _053317_, _053318_, _053319_, _053320_, _053321_, _053322_, _053323_, _053324_, _053325_, _053326_, _053327_, _053328_, _053329_, _053330_, _053331_, _053332_, _053333_, _053334_, _053335_, _053336_, _053337_, _053338_, _053339_, _053340_, _053341_, _053342_, _053343_, _053344_, _053345_, _053346_, _053347_, _053348_, _053349_, _053350_, _053351_, _053352_, _053353_, _053354_, _053355_, _053356_, _053357_, _053358_, _053359_, _053360_, _053361_, _053362_, _053363_, _053364_, _053365_, _053366_, _053367_, _053368_, _053369_, _053370_, _053371_, _053372_, _053373_, _053374_, _053375_, _053376_, _053377_, _053378_, _053379_, _053380_, _053381_, _053382_, _053383_, _053384_, _053385_, _053386_, _053387_, _053388_, _053389_, _053390_, _053391_, _053392_, _053393_, _053394_, _053395_, _053396_, _053397_, _053398_, _053399_, _053400_, _053401_, _053402_, _053403_, _053404_, _053405_, _053406_, _053407_, _053408_, _053409_, _053410_, _053411_, _053412_, _053413_, _053414_, _053415_, _053416_, _053417_, _053418_, _053419_, _053420_, _053421_, _053422_, _053423_, _053424_, _053425_, _053426_, _053427_, _053428_, _053429_, _053430_, _053431_, _053432_, _053433_, _053434_, _053435_, _053436_, _053437_, _053438_, _053439_, _053440_, _053441_, _053442_, _053443_, _053444_, _053445_, _053446_, _053447_, _053448_, _053449_, _053450_, _053451_, _053452_, _053453_, _053454_, _053455_, _053456_, _053457_, _053458_, _053459_, _053460_, _053461_, _053462_, _053463_, _053464_, _053465_, _053466_, _053467_, _053468_, _053469_, _053470_, _053471_, _053472_, _053473_, _053474_, _053475_, _053476_, _053477_, _053478_, _053479_, _053480_, _053481_, _053482_, _053483_, _053484_, _053485_, _053486_, _053487_, _053488_, _053489_, _053490_, _053491_, _053492_, _053493_, _053494_, _053495_, _053496_, _053497_, _053498_, _053499_, _053500_, _053501_, _053502_, _053503_, _053504_, _053505_, _053506_, _053507_, _053508_, _053509_, _053510_, _053511_, _053512_, _053513_, _053514_, _053515_, _053516_, _053517_, _053518_, _053519_, _053520_, _053521_, _053522_, _053523_, _053524_, _053525_, _053526_, _053527_, _053528_, _053529_, _053530_, _053531_, _053532_, _053533_, _053534_, _053535_, _053536_, _053537_, _053538_, _053539_, _053540_, _053541_, _053542_, _053543_, _053544_, _053545_, _053546_, _053547_, _053548_, _053549_, _053550_, _053551_, _053552_, _053553_, _053554_, _053555_, _053556_, _053557_, _053558_, _053559_, _053560_, _053561_, _053562_, _053563_, _053564_, _053565_, _053566_, _053567_, _053568_, _053569_, _053570_, _053571_, _053572_, _053573_, _053574_, _053575_, _053576_, _053577_, _053578_, _053579_, _053580_, _053581_, _053582_, _053583_, _053584_, _053585_, _053586_, _053587_, _053588_, _053589_, _053590_, _053591_, _053592_, _053593_, _053594_, _053595_, _053596_, _053597_, _053598_, _053599_, _053600_, _053601_, _053602_, _053603_, _053604_, _053605_, _053606_, _053607_, _053608_, _053609_, _053610_, _053611_, _053612_, _053613_, _053614_, _053615_, _053616_, _053617_, _053618_, _053619_, _053620_, _053621_, _053622_, _053623_, _053624_, _053625_, _053626_, _053627_, _053628_, _053629_, _053630_, _053631_, _053632_, _053633_, _053634_, _053635_, _053636_, _053637_, _053638_, _053639_, _053640_, _053641_, _053642_, _053643_, _053644_, _053645_, _053646_, _053647_, _053648_, _053649_, _053650_, _053651_, _053652_, _053653_, _053654_, _053655_, _053656_, _053657_, _053658_, _053659_, _053660_, _053661_, _053662_, _053663_, _053664_, _053665_, _053666_, _053667_, _053668_, _053669_, _053670_, _053671_, _053672_, _053673_, _053674_, _053675_, _053676_, _053677_, _053678_, _053679_, _053680_, _053681_, _053682_, _053683_, _053684_, _053685_, _053686_, _053687_, _053688_, _053689_, _053690_, _053691_, _053692_, _053693_, _053694_, _053695_, _053696_, _053697_, _053698_, _053699_, _053700_, _053701_, _053702_, _053703_, _053704_, _053705_, _053706_, _053707_, _053708_, _053709_, _053710_, _053711_, _053712_, _053713_, _053714_, _053715_, _053716_, _053717_, _053718_, _053719_, _053720_, _053721_, _053722_, _053723_, _053724_, _053725_, _053726_, _053727_, _053728_, _053729_, _053730_, _053731_, _053732_, _053733_, _053734_, _053735_, _053736_, _053737_, _053738_, _053739_, _053740_, _053741_, _053742_, _053743_, _053744_, _053745_, _053746_, _053747_, _053748_, _053749_, _053750_, _053751_, _053752_, _053753_, _053754_, _053755_, _053756_, _053757_, _053758_, _053759_, _053760_, _053761_, _053762_, _053763_, _053764_, _053765_, _053766_, _053767_, _053768_, _053769_, _053770_, _053771_, _053772_, _053773_, _053774_, _053775_, _053776_, _053777_, _053778_, _053779_, _053780_, _053781_, _053782_, _053783_, _053784_, _053785_, _053786_, _053787_, _053788_, _053789_, _053790_, _053791_, _053792_, _053793_, _053794_, _053795_, _053796_, _053797_, _053798_, _053799_, _053800_, _053801_, _053802_, _053803_, _053804_, _053805_, _053806_, _053807_, _053808_, _053809_, _053810_, _053811_, _053812_, _053813_, _053814_, _053815_, _053816_, _053817_, _053818_, _053819_, _053820_, _053821_, _053822_, _053823_, _053824_, _053825_, _053826_, _053827_, _053828_, _053829_, _053830_, _053831_, _053832_, _053833_, _053834_, _053835_, _053836_, _053837_, _053838_, _053839_, _053840_, _053841_, _053842_, _053843_, _053844_, _053845_, _053846_, _053847_, _053848_, _053849_, _053850_, _053851_, _053852_, _053853_, _053854_, _053855_, _053856_, _053857_, _053858_, _053859_, _053860_, _053861_, _053862_, _053863_, _053864_, _053865_, _053866_, _053867_, _053868_, _053869_, _053870_, _053871_, _053872_, _053873_, _053874_, _053875_, _053876_, _053877_, _053878_, _053879_, _053880_, _053881_, _053882_, _053883_, _053884_, _053885_, _053886_, _053887_, _053888_, _053889_, _053890_, _053891_, _053892_, _053893_, _053894_, _053895_, _053896_, _053897_, _053898_, _053899_, _053900_, _053901_, _053902_, _053903_, _053904_, _053905_, _053906_, _053907_, _053908_, _053909_, _053910_, _053911_, _053912_, _053913_, _053914_, _053915_, _053916_, _053917_, _053918_, _053919_, _053920_, _053921_, _053922_, _053923_, _053924_, _053925_, _053926_, _053927_, _053928_, _053929_, _053930_, _053931_, _053932_, _053933_, _053934_, _053935_, _053936_, _053937_, _053938_, _053939_, _053940_, _053941_, _053942_, _053943_, _053944_, _053945_, _053946_, _053947_, _053948_, _053949_, _053950_, _053951_, _053952_, _053953_, _053954_, _053955_, _053956_, _053957_, _053958_, _053959_, _053960_, _053961_, _053962_, _053963_, _053964_, _053965_, _053966_, _053967_, _053968_, _053969_, _053970_, _053971_, _053972_, _053973_, _053974_, _053975_, _053976_, _053977_, _053978_, _053979_, _053980_, _053981_, _053982_, _053983_, _053984_, _053985_, _053986_, _053987_, _053988_, _053989_, _053990_, _053991_, _053992_, _053993_, _053994_, _053995_, _053996_, _053997_, _053998_, _053999_, _054000_, _054001_, _054002_, _054003_, _054004_, _054005_, _054006_, _054007_, _054008_, _054009_, _054010_, _054011_, _054012_, _054013_, _054014_, _054015_, _054016_, _054017_, _054018_, _054019_, _054020_, _054021_, _054022_, _054023_, _054024_, _054025_, _054026_, _054027_, _054028_, _054029_, _054030_, _054031_, _054032_, _054033_, _054034_, _054035_, _054036_, _054037_, _054038_, _054039_, _054040_, _054041_, _054042_, _054043_, _054044_, _054045_, _054046_, _054047_, _054048_, _054049_, _054050_, _054051_, _054052_, _054053_, _054054_, _054055_, _054056_, _054057_, _054058_, _054059_, _054060_, _054061_, _054062_, _054063_, _054064_, _054065_, _054066_, _054067_, _054068_, _054069_, _054070_, _054071_, _054072_, _054073_, _054074_, _054075_, _054076_, _054077_, _054078_, _054079_, _054080_, _054081_, _054082_, _054083_, _054084_, _054085_, _054086_, _054087_, _054088_, _054089_, _054090_, _054091_, _054092_, _054093_, _054094_, _054095_, _054096_, _054097_, _054098_, _054099_, _054100_, _054101_, _054102_, _054103_, _054104_, _054105_, _054106_, _054107_, _054108_, _054109_, _054110_, _054111_, _054112_, _054113_, _054114_, _054115_, _054116_, _054117_, _054118_, _054119_, _054120_, _054121_, _054122_, _054123_, _054124_, _054125_, _054126_, _054127_, _054128_, _054129_, _054130_, _054131_, _054132_, _054133_, _054134_, _054135_, _054136_, _054137_, _054138_, _054139_, _054140_, _054141_, _054142_, _054143_, _054144_, _054145_, _054146_, _054147_, _054148_, _054149_, _054150_, _054151_, _054152_, _054153_, _054154_, _054155_, _054156_, _054157_, _054158_, _054159_, _054160_, _054161_, _054162_, _054163_, _054164_, _054165_, _054166_, _054167_, _054168_, _054169_, _054170_, _054171_, _054172_, _054173_, _054174_, _054175_, _054176_, _054177_, _054178_, _054179_, _054180_, _054181_, _054182_, _054183_, _054184_, _054185_, _054186_, _054187_, _054188_, _054189_, _054190_, _054191_, _054192_, _054193_, _054194_, _054195_, _054196_, _054197_, _054198_, _054199_, _054200_, _054201_, _054202_, _054203_, _054204_, _054205_, _054206_, _054207_, _054208_, _054209_, _054210_, _054211_, _054212_, _054213_, _054214_, _054215_, _054216_, _054217_, _054218_, _054219_, _054220_, _054221_, _054222_, _054223_, _054224_, _054225_, _054226_, _054227_, _054228_, _054229_, _054230_, _054231_, _054232_, _054233_, _054234_, _054235_, _054236_, _054237_, _054238_, _054239_, _054240_, _054241_, _054242_, _054243_, _054244_, _054245_, _054246_, _054247_, _054248_, _054249_, _054250_, _054251_, _054252_, _054253_, _054254_, _054255_, _054256_, _054257_, _054258_, _054259_, _054260_, _054261_, _054262_, _054263_, _054264_, _054265_, _054266_, _054267_, _054268_, _054269_, _054270_, _054271_, _054272_, _054273_, _054274_, _054275_, _054276_, _054277_, _054278_, _054279_, _054280_, _054281_, _054282_, _054283_, _054284_, _054285_, _054286_, _054287_, _054288_, _054289_, _054290_, _054291_, _054292_, _054293_, _054294_, _054295_, _054296_, _054297_, _054298_, _054299_, _054300_, _054301_, _054302_, _054303_, _054304_, _054305_, _054306_, _054307_, _054308_, _054309_, _054310_, _054311_, _054312_, _054313_, _054314_, _054315_, _054316_, _054317_, _054318_, _054319_, _054320_, _054321_, _054322_, _054323_, _054324_, _054325_, _054326_, _054327_, _054328_, _054329_, _054330_, _054331_, _054332_, _054333_, _054334_, _054335_, _054336_, _054337_, _054338_, _054339_, _054340_, _054341_, _054342_, _054343_, _054344_, _054345_, _054346_, _054347_, _054348_, _054349_, _054350_, _054351_, _054352_, _054353_, _054354_, _054355_, _054356_, _054357_, _054358_, _054359_, _054360_, _054361_, _054362_, _054363_, _054364_, _054365_, _054366_, _054367_, _054368_, _054369_, _054370_, _054371_, _054372_, _054373_, _054374_, _054375_, _054376_, _054377_, _054378_, _054379_, _054380_, _054381_, _054382_, _054383_, _054384_, _054385_, _054386_, _054387_, _054388_, _054389_, _054390_, _054391_, _054392_, _054393_, _054394_, _054395_, _054396_, _054397_, _054398_, _054399_, _054400_, _054401_, _054402_, _054403_, _054404_, _054405_, _054406_, _054407_, _054408_, _054409_, _054410_, _054411_, _054412_, _054413_, _054414_, _054415_, _054416_, _054417_, _054418_, _054419_, _054420_, _054421_, _054422_, _054423_, _054424_, _054425_, _054426_, _054427_, _054428_, _054429_, _054430_, _054431_, _054432_, _054433_, _054434_, _054435_, _054436_, _054437_, _054438_, _054439_, _054440_, _054441_, _054442_, _054443_, _054444_, _054445_, _054446_, _054447_, _054448_, _054449_, _054450_, _054451_, _054452_, _054453_, _054454_, _054455_, _054456_, _054457_, _054458_, _054459_, _054460_, _054461_, _054462_, _054463_, _054464_, _054465_, _054466_, _054467_, _054468_, _054469_, _054470_, _054471_, _054472_, _054473_, _054474_, _054475_, _054476_, _054477_, _054478_, _054479_, _054480_, _054481_, _054482_, _054483_, _054484_, _054485_, _054486_, _054487_, _054488_, _054489_, _054490_, _054491_, _054492_, _054493_, _054494_, _054495_, _054496_, _054497_, _054498_, _054499_, _054500_, _054501_, _054502_, _054503_, _054504_, _054505_, _054506_, _054507_, _054508_, _054509_, _054510_, _054511_, _054512_, _054513_, _054514_, _054515_, _054516_, _054517_, _054518_, _054519_, _054520_, _054521_, _054522_, _054523_, _054524_, _054525_, _054526_, _054527_, _054528_, _054529_, _054530_, _054531_, _054532_, _054533_, _054534_, _054535_, _054536_, _054537_, _054538_, _054539_, _054540_, _054541_, _054542_, _054543_, _054544_, _054545_, _054546_, _054547_, _054548_, _054549_, _054550_, _054551_, _054552_, _054553_, _054554_, _054555_, _054556_, _054557_, _054558_, _054559_, _054560_, _054561_, _054562_, _054563_, _054564_, _054565_, _054566_, _054567_, _054568_, _054569_, _054570_, _054571_, _054572_, _054573_, _054574_, _054575_, _054576_, _054577_, _054578_, _054579_, _054580_, _054581_, _054582_, _054583_, _054584_, _054585_, _054586_, _054587_, _054588_, _054589_, _054590_, _054591_, _054592_, _054593_, _054594_, _054595_, _054596_, _054597_, _054598_, _054599_, _054600_, _054601_, _054602_, _054603_, _054604_, _054605_, _054606_, _054607_, _054608_, _054609_, _054610_, _054611_, _054612_, _054613_, _054614_, _054615_, _054616_, _054617_, _054618_, _054619_, _054620_, _054621_, _054622_, _054623_, _054624_, _054625_, _054626_, _054627_, _054628_, _054629_, _054630_, _054631_, _054632_, _054633_, _054634_, _054635_, _054636_, _054637_, _054638_, _054639_, _054640_, _054641_, _054642_, _054643_, _054644_, _054645_, _054646_, _054647_, _054648_, _054649_, _054650_, _054651_, _054652_, _054653_, _054654_, _054655_, _054656_, _054657_, _054658_, _054659_, _054660_, _054661_, _054662_, _054663_, _054664_, _054665_, _054666_, _054667_, _054668_, _054669_, _054670_, _054671_, _054672_, _054673_, _054674_, _054675_, _054676_, _054677_, _054678_, _054679_, _054680_, _054681_, _054682_, _054683_, _054684_, _054685_, _054686_, _054687_, _054688_, _054689_, _054690_, _054691_, _054692_, _054693_, _054694_, _054695_, _054696_, _054697_, _054698_, _054699_, _054700_, _054701_, _054702_, _054703_, _054704_, _054705_, _054706_, _054707_, _054708_, _054709_, _054710_, _054711_, _054712_, _054713_, _054714_, _054715_, _054716_, _054717_, _054718_, _054719_, _054720_, _054721_, _054722_, _054723_, _054724_, _054725_, _054726_, _054727_, _054728_, _054729_, _054730_, _054731_, _054732_, _054733_, _054734_, _054735_, _054736_, _054737_, _054738_, _054739_, _054740_, _054741_, _054742_, _054743_, _054744_, _054745_, _054746_, _054747_, _054748_, _054749_, _054750_, _054751_, _054752_, _054753_, _054754_, _054755_, _054756_, _054757_, _054758_, _054759_, _054760_, _054761_, _054762_, _054763_, _054764_, _054765_, _054766_, _054767_, _054768_, _054769_, _054770_, _054771_, _054772_, _054773_, _054774_, _054775_, _054776_, _054777_, _054778_, _054779_, _054780_, _054781_, _054782_, _054783_, _054784_, _054785_, _054786_, _054787_, _054788_, _054789_, _054790_, _054791_, _054792_, _054793_, _054794_, _054795_, _054796_, _054797_, _054798_, _054799_, _054800_, _054801_, _054802_, _054803_, _054804_, _054805_, _054806_, _054807_, _054808_, _054809_, _054810_, _054811_, _054812_, _054813_, _054814_, _054815_, _054816_, _054817_, _054818_, _054819_, _054820_, _054821_, _054822_, _054823_, _054824_, _054825_, _054826_, _054827_, _054828_, _054829_, _054830_, _054831_, _054832_, _054833_, _054834_, _054835_, _054836_, _054837_, _054838_, _054839_, _054840_, _054841_, _054842_, _054843_, _054844_, _054845_, _054846_, _054847_, _054848_, _054849_, _054850_, _054851_, _054852_, _054853_, _054854_, _054855_, _054856_, _054857_, _054858_, _054859_, _054860_, _054861_, _054862_, _054863_, _054864_, _054865_, _054866_, _054867_, _054868_, _054869_, _054870_, _054871_, _054872_, _054873_, _054874_, _054875_, _054876_, _054877_, _054878_, _054879_, _054880_, _054881_, _054882_, _054883_, _054884_, _054885_, _054886_, _054887_, _054888_, _054889_, _054890_, _054891_, _054892_, _054893_, _054894_, _054895_, _054896_, _054897_, _054898_, _054899_, _054900_, _054901_, _054902_, _054903_, _054904_, _054905_, _054906_, _054907_, _054908_, _054909_, _054910_, _054911_, _054912_, _054913_, _054914_, _054915_, _054916_, _054917_, _054918_, _054919_, _054920_, _054921_, _054922_, _054923_, _054924_, _054925_, _054926_, _054927_, _054928_, _054929_, _054930_, _054931_, _054932_, _054933_, _054934_, _054935_, _054936_, _054937_, _054938_, _054939_, _054940_, _054941_, _054942_, _054943_, _054944_, _054945_, _054946_, _054947_, _054948_, _054949_, _054950_, _054951_, _054952_, _054953_, _054954_, _054955_, _054956_, _054957_, _054958_, _054959_, _054960_, _054961_, _054962_, _054963_, _054964_, _054965_, _054966_, _054967_, _054968_, _054969_, _054970_, _054971_, _054972_, _054973_, _054974_, _054975_, _054976_, _054977_, _054978_, _054979_, _054980_, _054981_, _054982_, _054983_, _054984_, _054985_, _054986_, _054987_, _054988_, _054989_, _054990_, _054991_, _054992_, _054993_, _054994_, _054995_, _054996_, _054997_, _054998_, _054999_, _055000_, _055001_, _055002_, _055003_, _055004_, _055005_, _055006_, _055007_, _055008_, _055009_, _055010_, _055011_, _055012_, _055013_, _055014_, _055015_, _055016_, _055017_, _055018_, _055019_, _055020_, _055021_, _055022_, _055023_, _055024_, _055025_, _055026_, _055027_, _055028_, _055029_, _055030_, _055031_, _055032_, _055033_, _055034_, _055035_, _055036_, _055037_, _055038_, _055039_, _055040_, _055041_, _055042_, _055043_, _055044_, _055045_, _055046_, _055047_, _055048_, _055049_, _055050_, _055051_, _055052_, _055053_, _055054_, _055055_, _055056_, _055057_, _055058_, _055059_, _055060_, _055061_, _055062_, _055063_, _055064_, _055065_, _055066_, _055067_, _055068_, _055069_, _055070_, _055071_, _055072_, _055073_, _055074_, _055075_, _055076_, _055077_, _055078_, _055079_, _055080_, _055081_, _055082_, _055083_, _055084_, _055085_, _055086_, _055087_, _055088_, _055089_, _055090_, _055091_, _055092_, _055093_, _055094_, _055095_, _055096_, _055097_, _055098_, _055099_, _055100_, _055101_, _055102_, _055103_, _055104_, _055105_, _055106_, _055107_, _055108_, _055109_, _055110_, _055111_, _055112_, _055113_, _055114_, _055115_, _055116_, _055117_, _055118_, _055119_, _055120_, _055121_, _055122_, _055123_, _055124_, _055125_, _055126_, _055127_, _055128_, _055129_, _055130_, _055131_, _055132_, _055133_, _055134_, _055135_, _055136_, _055137_, _055138_, _055139_, _055140_, _055141_, _055142_, _055143_, _055144_, _055145_, _055146_, _055147_, _055148_, _055149_, _055150_, _055151_, _055152_, _055153_, _055154_, _055155_, _055156_, _055157_, _055158_, _055159_, _055160_, _055161_, _055162_, _055163_, _055164_, _055165_, _055166_, _055167_, _055168_, _055169_, _055170_, _055171_, _055172_, _055173_, _055174_, _055175_, _055176_, _055177_, _055178_, _055179_, _055180_, _055181_, _055182_, _055183_, _055184_, _055185_, _055186_, _055187_, _055188_, _055189_, _055190_, _055191_, _055192_, _055193_, _055194_, _055195_, _055196_, _055197_, _055198_, _055199_, _055200_, _055201_, _055202_, _055203_, _055204_, _055205_, _055206_, _055207_, _055208_, _055209_, _055210_, _055211_, _055212_, _055213_, _055214_, _055215_, _055216_, _055217_, _055218_, _055219_, _055220_, _055221_, _055222_, _055223_, _055224_, _055225_, _055226_, _055227_, _055228_, _055229_, _055230_, _055231_, _055232_, _055233_, _055234_, _055235_, _055236_, _055237_, _055238_, _055239_, _055240_, _055241_, _055242_, _055243_, _055244_, _055245_, _055246_, _055247_, _055248_, _055249_, _055250_, _055251_, _055252_, _055253_, _055254_, _055255_, _055256_, _055257_, _055258_, _055259_, _055260_, _055261_, _055262_, _055263_, _055264_, _055265_, _055266_, _055267_, _055268_, _055269_, _055270_, _055271_, _055272_, _055273_, _055274_, _055275_, _055276_, _055277_, _055278_, _055279_, _055280_, _055281_, _055282_, _055283_, _055284_, _055285_, _055286_, _055287_, _055288_, _055289_, _055290_, _055291_, _055292_, _055293_, _055294_, _055295_, _055296_, _055297_, _055298_, _055299_, _055300_, _055301_, _055302_, _055303_, _055304_, _055305_, _055306_, _055307_, _055308_, _055309_, _055310_, _055311_, _055312_, _055313_, _055314_, _055315_, _055316_, _055317_, _055318_, _055319_, _055320_, _055321_, _055322_, _055323_, _055324_, _055325_, _055326_, _055327_, _055328_, _055329_, _055330_, _055331_, _055332_, _055333_, _055334_, _055335_, _055336_, _055337_, _055338_, _055339_, _055340_, _055341_, _055342_, _055343_, _055344_, _055345_, _055346_, _055347_, _055348_, _055349_, _055350_, _055351_, _055352_, _055353_, _055354_, _055355_, _055356_, _055357_, _055358_, _055359_, _055360_, _055361_, _055362_, _055363_, _055364_, _055365_, _055366_, _055367_, _055368_, _055369_, _055370_, _055371_, _055372_, _055373_, _055374_, _055375_, _055376_, _055377_, _055378_, _055379_, _055380_, _055381_, _055382_, _055383_, _055384_, _055385_, _055386_, _055387_, _055388_, _055389_, _055390_, _055391_, _055392_, _055393_, _055394_, _055395_, _055396_, _055397_, _055398_, _055399_, _055400_, _055401_, _055402_, _055403_, _055404_, _055405_, _055406_, _055407_, _055408_, _055409_, _055410_, _055411_, _055412_, _055413_, _055414_, _055415_, _055416_, _055417_, _055418_, _055419_, _055420_, _055421_, _055422_, _055423_, _055424_, _055425_, _055426_, _055427_, _055428_, _055429_, _055430_, _055431_, _055432_, _055433_, _055434_, _055435_, _055436_, _055437_, _055438_, _055439_, _055440_, _055441_, _055442_, _055443_, _055444_, _055445_, _055446_, _055447_, _055448_, _055449_, _055450_, _055451_, _055452_, _055453_, _055454_, _055455_, _055456_, _055457_, _055458_, _055459_, _055460_, _055461_, _055462_, _055463_, _055464_, _055465_, _055466_, _055467_, _055468_, _055469_, _055470_, _055471_, _055472_, _055473_, _055474_, _055475_, _055476_, _055477_, _055478_, _055479_, _055480_, _055481_, _055482_, _055483_, _055484_, _055485_, _055486_, _055487_, _055488_, _055489_, _055490_, _055491_, _055492_, _055493_, _055494_, _055495_, _055496_, _055497_, _055498_, _055499_, _055500_, _055501_, _055502_, _055503_, _055504_, _055505_, _055506_, _055507_, _055508_, _055509_, _055510_, _055511_, _055512_, _055513_, _055514_, _055515_, _055516_, _055517_, _055518_, _055519_, _055520_, _055521_, _055522_, _055523_, _055524_, _055525_, _055526_, _055527_, _055528_, _055529_, _055530_, _055531_, _055532_, _055533_, _055534_, _055535_, _055536_, _055537_, _055538_, _055539_, _055540_, _055541_, _055542_, _055543_, _055544_, _055545_, _055546_, _055547_, _055548_, _055549_, _055550_, _055551_, _055552_, _055553_, _055554_, _055555_, _055556_, _055557_, _055558_, _055559_, _055560_, _055561_, _055562_, _055563_, _055564_, _055565_, _055566_, _055567_, _055568_, _055569_, _055570_, _055571_, _055572_, _055573_, _055574_, _055575_, _055576_, _055577_, _055578_, _055579_, _055580_, _055581_, _055582_, _055583_, _055584_, _055585_, _055586_, _055587_, _055588_, _055589_, _055590_, _055591_, _055592_, _055593_, _055594_, _055595_, _055596_, _055597_, _055598_, _055599_, _055600_, _055601_, _055602_, _055603_, _055604_, _055605_, _055606_, _055607_, _055608_, _055609_, _055610_, _055611_, _055612_, _055613_, _055614_, _055615_, _055616_, _055617_, _055618_, _055619_, _055620_, _055621_, _055622_, _055623_, _055624_, _055625_, _055626_, _055627_, _055628_, _055629_, _055630_, _055631_, _055632_, _055633_, _055634_, _055635_, _055636_, _055637_, _055638_, _055639_, _055640_, _055641_, _055642_, _055643_, _055644_, _055645_, _055646_, _055647_, _055648_, _055649_, _055650_, _055651_, _055652_, _055653_, _055654_, _055655_, _055656_, _055657_, _055658_, _055659_, _055660_, _055661_, _055662_, _055663_, _055664_, _055665_, _055666_, _055667_, _055668_, _055669_, _055670_, _055671_, _055672_, _055673_, _055674_, _055675_, _055676_, _055677_, _055678_, _055679_, _055680_, _055681_, _055682_, _055683_, _055684_, _055685_, _055686_, _055687_, _055688_, _055689_, _055690_, _055691_, _055692_, _055693_, _055694_, _055695_, _055696_, _055697_, _055698_, _055699_, _055700_, _055701_, _055702_, _055703_, _055704_, _055705_, _055706_, _055707_, _055708_, _055709_, _055710_, _055711_, _055712_, _055713_, _055714_, _055715_, _055716_, _055717_, _055718_, _055719_, _055720_, _055721_, _055722_, _055723_, _055724_, _055725_, _055726_, _055727_, _055728_, _055729_, _055730_, _055731_, _055732_, _055733_, _055734_, _055735_, _055736_, _055737_, _055738_, _055739_, _055740_, _055741_, _055742_, _055743_, _055744_, _055745_, _055746_, _055747_, _055748_, _055749_, _055750_, _055751_, _055752_, _055753_, _055754_, _055755_, _055756_, _055757_, _055758_, _055759_, _055760_, _055761_, _055762_, _055763_, _055764_, _055765_, _055766_, _055767_, _055768_, _055769_, _055770_, _055771_, _055772_, _055773_, _055774_, _055775_, _055776_, _055777_, _055778_, _055779_, _055780_, _055781_, _055782_, _055783_, _055784_, _055785_, _055786_, _055787_, _055788_, _055789_, _055790_, _055791_, _055792_, _055793_, _055794_, _055795_, _055796_, _055797_, _055798_, _055799_, _055800_, _055801_, _055802_, _055803_, _055804_, _055805_, _055806_, _055807_, _055808_, _055809_, _055810_, _055811_, _055812_, _055813_, _055814_, _055815_, _055816_, _055817_, _055818_, _055819_, _055820_, _055821_, _055822_, _055823_, _055824_, _055825_, _055826_, _055827_, _055828_, _055829_, _055830_, _055831_, _055832_, _055833_, _055834_, _055835_, _055836_, _055837_, _055838_, _055839_, _055840_, _055841_, _055842_, _055843_, _055844_, _055845_, _055846_, _055847_, _055848_, _055849_, _055850_, _055851_, _055852_, _055853_, _055854_, _055855_, _055856_, _055857_, _055858_, _055859_, _055860_, _055861_, _055862_, _055863_, _055864_, _055865_, _055866_, _055867_, _055868_, _055869_, _055870_, _055871_, _055872_, _055873_, _055874_, _055875_, _055876_, _055877_, _055878_, _055879_, _055880_, _055881_, _055882_, _055883_, _055884_, _055885_, _055886_, _055887_, _055888_, _055889_, _055890_, _055891_, _055892_, _055893_, _055894_, _055895_, _055896_, _055897_, _055898_, _055899_, _055900_, _055901_, _055902_, _055903_, _055904_, _055905_, _055906_, _055907_, _055908_, _055909_, _055910_, _055911_, _055912_, _055913_, _055914_, _055915_, _055916_, _055917_, _055918_, _055919_, _055920_, _055921_, _055922_, _055923_, _055924_, _055925_, _055926_, _055927_, _055928_, _055929_, _055930_, _055931_, _055932_, _055933_, _055934_, _055935_, _055936_, _055937_, _055938_, _055939_, _055940_, _055941_, _055942_, _055943_, _055944_, _055945_, _055946_, _055947_, _055948_, _055949_, _055950_, _055951_, _055952_, _055953_, _055954_, _055955_, _055956_, _055957_, _055958_, _055959_, _055960_, _055961_, _055962_, _055963_, _055964_, _055965_, _055966_, _055967_, _055968_, _055969_, _055970_, _055971_, _055972_, _055973_, _055974_, _055975_, _055976_, _055977_, _055978_, _055979_, _055980_, _055981_, _055982_, _055983_, _055984_, _055985_, _055986_, _055987_, _055988_, _055989_, _055990_, _055991_, _055992_, _055993_, _055994_, _055995_, _055996_, _055997_, _055998_, _055999_, _056000_, _056001_, _056002_, _056003_, _056004_, _056005_, _056006_, _056007_, _056008_, _056009_, _056010_, _056011_, _056012_, _056013_, _056014_, _056015_, _056016_, _056017_, _056018_, _056019_, _056020_, _056021_, _056022_, _056023_, _056024_, _056025_, _056026_, _056027_, _056028_, _056029_, _056030_, _056031_, _056032_, _056033_, _056034_, _056035_, _056036_, _056037_, _056038_, _056039_, _056040_, _056041_, _056042_, _056043_, _056044_, _056045_, _056046_, _056047_, _056048_, _056049_, _056050_, _056051_, _056052_, _056053_, _056054_, _056055_, _056056_, _056057_, _056058_, _056059_, _056060_, _056061_, _056062_, _056063_, _056064_, _056065_, _056066_, _056067_, _056068_, _056069_, _056070_, _056071_, _056072_, _056073_, _056074_, _056075_, _056076_, _056077_, _056078_, _056079_, _056080_, _056081_, _056082_, _056083_, _056084_, _056085_, _056086_, _056087_, _056088_, _056089_, _056090_, _056091_, _056092_, _056093_, _056094_, _056095_, _056096_, _056097_, _056098_, _056099_, _056100_, _056101_, _056102_, _056103_, _056104_, _056105_, _056106_, _056107_, _056108_, _056109_, _056110_, _056111_, _056112_, _056113_, _056114_, _056115_, _056116_, _056117_, _056118_, _056119_, _056120_, _056121_, _056122_, _056123_, _056124_, _056125_, _056126_, _056127_, _056128_, _056129_, _056130_, _056131_, _056132_, _056133_, _056134_, _056135_, _056136_, _056137_, _056138_, _056139_, _056140_, _056141_, _056142_, _056143_, _056144_, _056145_, _056146_, _056147_, _056148_, _056149_, _056150_, _056151_, _056152_, _056153_, _056154_, _056155_, _056156_, _056157_, _056158_, _056159_, _056160_, _056161_, _056162_, _056163_, _056164_, _056165_, _056166_, _056167_, _056168_, _056169_, _056170_, _056171_, _056172_, _056173_, _056174_, _056175_, _056176_, _056177_, _056178_, _056179_, _056180_, _056181_, _056182_, _056183_, _056184_, _056185_, _056186_, _056187_, _056188_, _056189_, _056190_, _056191_, _056192_, _056193_, _056194_, _056195_, _056196_, _056197_, _056198_, _056199_, _056200_, _056201_, _056202_, _056203_, _056204_, _056205_, _056206_, _056207_, _056208_, _056209_, _056210_, _056211_, _056212_, _056213_, _056214_, _056215_, _056216_, _056217_, _056218_, _056219_, _056220_, _056221_, _056222_, _056223_, _056224_, _056225_, _056226_, _056227_, _056228_, _056229_, _056230_, _056231_, _056232_, _056233_, _056234_, _056235_, _056236_, _056237_, _056238_, _056239_, _056240_, _056241_, _056242_, _056243_, _056244_, _056245_, _056246_, _056247_, _056248_, _056249_, _056250_, _056251_, _056252_, _056253_, _056254_, _056255_, _056256_, _056257_, _056258_, _056259_, _056260_, _056261_, _056262_, _056263_, _056264_, _056265_, _056266_, _056267_, _056268_, _056269_, _056270_, _056271_, _056272_, _056273_, _056274_, _056275_, _056276_, _056277_, _056278_, _056279_, _056280_, _056281_, _056282_, _056283_, _056284_, _056285_, _056286_, _056287_, _056288_, _056289_, _056290_, _056291_, _056292_, _056293_, _056294_, _056295_, _056296_, _056297_, _056298_, _056299_, _056300_, _056301_, _056302_, _056303_, _056304_, _056305_, _056306_, _056307_, _056308_, _056309_, _056310_, _056311_, _056312_, _056313_, _056314_, _056315_, _056316_, _056317_, _056318_, _056319_, _056320_, _056321_, _056322_, _056323_, _056324_, _056325_, _056326_, _056327_, _056328_, _056329_, _056330_, _056331_, _056332_, _056333_, _056334_, _056335_, _056336_, _056337_, _056338_, _056339_, _056340_, _056341_, _056342_, _056343_, _056344_, _056345_, _056346_, _056347_, _056348_, _056349_, _056350_, _056351_, _056352_, _056353_, _056354_, _056355_, _056356_, _056357_, _056358_, _056359_, _056360_, _056361_, _056362_, _056363_, _056364_, _056365_, _056366_, _056367_, _056368_, _056369_, _056370_, _056371_, _056372_, _056373_, _056374_, _056375_, _056376_, _056377_, _056378_, _056379_, _056380_, _056381_, _056382_, _056383_, _056384_, _056385_, _056386_, _056387_, _056388_, _056389_, _056390_, _056391_, _056392_, _056393_, _056394_, _056395_, _056396_, _056397_, _056398_, _056399_, _056400_, _056401_, _056402_, _056403_, _056404_, _056405_, _056406_, _056407_, _056408_, _056409_, _056410_, _056411_, _056412_, _056413_, _056414_, _056415_, _056416_, _056417_, _056418_, _056419_, _056420_, _056421_, _056422_, _056423_, _056424_, _056425_, _056426_, _056427_, _056428_, _056429_, _056430_, _056431_, _056432_, _056433_, _056434_, _056435_, _056436_, _056437_, _056438_, _056439_, _056440_, _056441_, _056442_, _056443_, _056444_, _056445_, _056446_, _056447_, _056448_, _056449_, _056450_, _056451_, _056452_, _056453_, _056454_, _056455_, _056456_, _056457_, _056458_, _056459_, _056460_, _056461_, _056462_, _056463_, _056464_, _056465_, _056466_, _056467_, _056468_, _056469_, _056470_, _056471_, _056472_, _056473_, _056474_, _056475_, _056476_, _056477_, _056478_, _056479_, _056480_, _056481_, _056482_, _056483_, _056484_, _056485_, _056486_, _056487_, _056488_, _056489_, _056490_, _056491_, _056492_, _056493_, _056494_, _056495_, _056496_, _056497_, _056498_, _056499_, _056500_, _056501_, _056502_, _056503_, _056504_, _056505_, _056506_, _056507_, _056508_, _056509_, _056510_, _056511_, _056512_, _056513_, _056514_, _056515_, _056516_, _056517_, _056518_, _056519_, _056520_, _056521_, _056522_, _056523_, _056524_, _056525_, _056526_, _056527_, _056528_, _056529_, _056530_, _056531_, _056532_, _056533_, _056534_, _056535_, _056536_, _056537_, _056538_, _056539_, _056540_, _056541_, _056542_, _056543_, _056544_, _056545_, _056546_, _056547_, _056548_, _056549_, _056550_, _056551_, _056552_, _056553_, _056554_, _056555_, _056556_, _056557_, _056558_, _056559_, _056560_, _056561_, _056562_, _056563_, _056564_, _056565_, _056566_, _056567_, _056568_, _056569_, _056570_, _056571_, _056572_, _056573_, _056574_, _056575_, _056576_, _056577_, _056578_, _056579_, _056580_, _056581_, _056582_, _056583_, _056584_, _056585_, _056586_, _056587_, _056588_, _056589_, _056590_, _056591_, _056592_, _056593_, _056594_, _056595_, _056596_, _056597_, _056598_, _056599_, _056600_, _056601_, _056602_, _056603_, _056604_, _056605_, _056606_, _056607_, _056608_, _056609_, _056610_, _056611_, _056612_, _056613_, _056614_, _056615_, _056616_, _056617_, _056618_, _056619_, _056620_, _056621_, _056622_, _056623_, _056624_, _056625_, _056626_, _056627_, _056628_, _056629_, _056630_, _056631_, _056632_, _056633_, _056634_, _056635_, _056636_, _056637_, _056638_, _056639_, _056640_, _056641_, _056642_, _056643_, _056644_, _056645_, _056646_, _056647_, _056648_, _056649_, _056650_, _056651_, _056652_, _056653_, _056654_, _056655_, _056656_, _056657_, _056658_, _056659_, _056660_, _056661_, _056662_, _056663_, _056664_, _056665_, _056666_, _056667_, _056668_, _056669_, _056670_, _056671_, _056672_, _056673_, _056674_, _056675_, _056676_, _056677_, _056678_, _056679_, _056680_, _056681_, _056682_, _056683_, _056684_, _056685_, _056686_, _056687_, _056688_, _056689_, _056690_, _056691_, _056692_, _056693_, _056694_, _056695_, _056696_, _056697_, _056698_, _056699_, _056700_, _056701_, _056702_, _056703_, _056704_, _056705_, _056706_, _056707_, _056708_, _056709_, _056710_, _056711_, _056712_, _056713_, _056714_, _056715_, _056716_, _056717_, _056718_, _056719_, _056720_, _056721_, _056722_, _056723_, _056724_, _056725_, _056726_, _056727_, _056728_, _056729_, _056730_, _056731_, _056732_, _056733_, _056734_, _056735_, _056736_, _056737_, _056738_, _056739_, _056740_, _056741_, _056742_, _056743_, _056744_, _056745_, _056746_, _056747_, _056748_, _056749_, _056750_, _056751_, _056752_, _056753_, _056754_, _056755_, _056756_, _056757_, _056758_, _056759_, _056760_, _056761_, _056762_, _056763_, _056764_, _056765_, _056766_, _056767_, _056768_, _056769_, _056770_, _056771_, _056772_, _056773_, _056774_, _056775_, _056776_, _056777_, _056778_, _056779_, _056780_, _056781_, _056782_, _056783_, _056784_, _056785_, _056786_, _056787_, _056788_, _056789_, _056790_, _056791_, _056792_, _056793_, _056794_, _056795_, _056796_, _056797_, _056798_, _056799_, _056800_, _056801_, _056802_, _056803_, _056804_, _056805_, _056806_, _056807_, _056808_, _056809_, _056810_, _056811_, _056812_, _056813_, _056814_, _056815_, _056816_, _056817_, _056818_, _056819_, _056820_, _056821_, _056822_, _056823_, _056824_, _056825_, _056826_, _056827_, _056828_, _056829_, _056830_, _056831_, _056832_, _056833_, _056834_, _056835_, _056836_, _056837_, _056838_, _056839_, _056840_, _056841_, _056842_, _056843_, _056844_, _056845_, _056846_, _056847_, _056848_, _056849_, _056850_, _056851_, _056852_, _056853_, _056854_, _056855_, _056856_, _056857_, _056858_, _056859_, _056860_, _056861_, _056862_, _056863_, _056864_, _056865_, _056866_, _056867_, _056868_, _056869_, _056870_, _056871_, _056872_, _056873_, _056874_, _056875_, _056876_, _056877_, _056878_, _056879_, _056880_, _056881_, _056882_, _056883_, _056884_, _056885_, _056886_, _056887_, _056888_, _056889_, _056890_, _056891_, _056892_, _056893_, _056894_, _056895_, _056896_, _056897_, _056898_, _056899_, _056900_, _056901_, _056902_, _056903_, _056904_, _056905_, _056906_, _056907_, _056908_, _056909_, _056910_, _056911_, _056912_, _056913_, _056914_, _056915_, _056916_, _056917_, _056918_, _056919_, _056920_, _056921_, _056922_, _056923_, _056924_, _056925_, _056926_, _056927_, _056928_, _056929_, _056930_, _056931_, _056932_, _056933_, _056934_, _056935_, _056936_, _056937_, _056938_, _056939_, _056940_, _056941_, _056942_, _056943_, _056944_, _056945_, _056946_, _056947_, _056948_, _056949_, _056950_, _056951_, _056952_, _056953_, _056954_, _056955_, _056956_, _056957_, _056958_, _056959_, _056960_, _056961_, _056962_, _056963_, _056964_, _056965_, _056966_, _056967_, _056968_, _056969_, _056970_, _056971_, _056972_, _056973_, _056974_, _056975_, _056976_, _056977_, _056978_, _056979_, _056980_, _056981_, _056982_, _056983_, _056984_, _056985_, _056986_, _056987_, _056988_, _056989_, _056990_, _056991_, _056992_, _056993_, _056994_, _056995_, _056996_, _056997_, _056998_, _056999_, _057000_, _057001_, _057002_, _057003_, _057004_, _057005_, _057006_, _057007_, _057008_, _057009_, _057010_, _057011_, _057012_, _057013_, _057014_, _057015_, _057016_, _057017_, _057018_, _057019_, _057020_, _057021_, _057022_, _057023_, _057024_, _057025_, _057026_, _057027_, _057028_, _057029_, _057030_, _057031_, _057032_, _057033_, _057034_, _057035_, _057036_, _057037_, _057038_, _057039_, _057040_, _057041_, _057042_, _057043_, _057044_, _057045_, _057046_, _057047_, _057048_, _057049_, _057050_, _057051_, _057052_, _057053_, _057054_, _057055_, _057056_, _057057_, _057058_, _057059_, _057060_, _057061_, _057062_, _057063_, _057064_, _057065_, _057066_, _057067_, _057068_, _057069_, _057070_, _057071_, _057072_, _057073_, _057074_, _057075_, _057076_, _057077_, _057078_, _057079_, _057080_, _057081_, _057082_, _057083_, _057084_, _057085_, _057086_, _057087_, _057088_, _057089_, _057090_, _057091_, _057092_, _057093_, _057094_, _057095_, _057096_, _057097_, _057098_, _057099_, _057100_, _057101_, _057102_, _057103_, _057104_, _057105_, _057106_, _057107_, _057108_, _057109_, _057110_, _057111_, _057112_, _057113_, _057114_, _057115_, _057116_, _057117_, _057118_, _057119_, _057120_, _057121_, _057122_, _057123_, _057124_, _057125_, _057126_, _057127_, _057128_, _057129_, _057130_, _057131_, _057132_, _057133_, _057134_, _057135_, _057136_, _057137_, _057138_, _057139_, _057140_, _057141_, _057142_, _057143_, _057144_, _057145_, _057146_, _057147_, _057148_, _057149_, _057150_, _057151_, _057152_, _057153_, _057154_, _057155_, _057156_, _057157_, _057158_, _057159_, _057160_, _057161_, _057162_, _057163_, _057164_, _057165_, _057166_, _057167_, _057168_, _057169_, _057170_, _057171_, _057172_, _057173_, _057174_, _057175_, _057176_, _057177_, _057178_, _057179_, _057180_, _057181_, _057182_, _057183_, _057184_, _057185_, _057186_, _057187_, _057188_, _057189_, _057190_, _057191_, _057192_, _057193_, _057194_, _057195_, _057196_, _057197_, _057198_, _057199_, _057200_, _057201_, _057202_, _057203_, _057204_, _057205_, _057206_, _057207_, _057208_, _057209_, _057210_, _057211_, _057212_, _057213_, _057214_, _057215_, _057216_, _057217_, _057218_, _057219_, _057220_, _057221_, _057222_, _057223_, _057224_, _057225_, _057226_, _057227_, _057228_, _057229_, _057230_, _057231_, _057232_, _057233_, _057234_, _057235_, _057236_, _057237_, _057238_, _057239_, _057240_, _057241_, _057242_, _057243_, _057244_, _057245_, _057246_, _057247_, _057248_, _057249_, _057250_, _057251_, _057252_, _057253_, _057254_, _057255_, _057256_, _057257_, _057258_, _057259_, _057260_, _057261_, _057262_, _057263_, _057264_, _057265_, _057266_, _057267_, _057268_, _057269_, _057270_, _057271_, _057272_, _057273_, _057274_, _057275_, _057276_, _057277_, _057278_, _057279_, _057280_, _057281_, _057282_, _057283_, _057284_, _057285_, _057286_, _057287_, _057288_, _057289_, _057290_, _057291_, _057292_, _057293_, _057294_, _057295_, _057296_, _057297_, _057298_, _057299_, _057300_, _057301_, _057302_, _057303_, _057304_, _057305_, _057306_, _057307_, _057308_, _057309_, _057310_, _057311_, _057312_, _057313_, _057314_, _057315_, _057316_, _057317_, _057318_, _057319_, _057320_, _057321_, _057322_, _057323_, _057324_, _057325_, _057326_, _057327_, _057328_, _057329_, _057330_, _057331_, _057332_, _057333_, _057334_, _057335_, _057336_, _057337_, _057338_, _057339_, _057340_, _057341_, _057342_, _057343_, _057344_, _057345_, _057346_, _057347_, _057348_, _057349_, _057350_, _057351_, _057352_, _057353_, _057354_, _057355_, _057356_, _057357_, _057358_, _057359_, _057360_, _057361_, _057362_, _057363_, _057364_, _057365_, _057366_, _057367_, _057368_, _057369_, _057370_, _057371_, _057372_, _057373_, _057374_, _057375_, _057376_, _057377_, _057378_, _057379_, _057380_, _057381_, _057382_, _057383_, _057384_, _057385_, _057386_, _057387_, _057388_, _057389_, _057390_, _057391_, _057392_, _057393_, _057394_, _057395_, _057396_, _057397_, _057398_, _057399_, _057400_, _057401_, _057402_, _057403_, _057404_, _057405_, _057406_, _057407_, _057408_, _057409_, _057410_, _057411_, _057412_, _057413_, _057414_, _057415_, _057416_, _057417_, _057418_, _057419_, _057420_, _057421_, _057422_, _057423_, _057424_, _057425_, _057426_, _057427_, _057428_, _057429_, _057430_, _057431_, _057432_, _057433_, _057434_, _057435_, _057436_, _057437_, _057438_, _057439_, _057440_, _057441_, _057442_, _057443_, _057444_, _057445_, _057446_, _057447_, _057448_, _057449_, _057450_, _057451_, _057452_, _057453_, _057454_, _057455_, _057456_, _057457_, _057458_, _057459_, _057460_, _057461_, _057462_, _057463_, _057464_, _057465_, _057466_, _057467_, _057468_, _057469_, _057470_, _057471_, _057472_, _057473_, _057474_, _057475_, _057476_, _057477_, _057478_, _057479_, _057480_, _057481_, _057482_, _057483_, _057484_, _057485_, _057486_, _057487_, _057488_, _057489_, _057490_, _057491_, _057492_, _057493_, _057494_, _057495_, _057496_, _057497_, _057498_, _057499_, _057500_, _057501_, _057502_, _057503_, _057504_, _057505_, _057506_, _057507_, _057508_, _057509_, _057510_, _057511_, _057512_, _057513_, _057514_, _057515_, _057516_, _057517_, _057518_, _057519_, _057520_, _057521_, _057522_, _057523_, _057524_, _057525_, _057526_, _057527_, _057528_, _057529_, _057530_, _057531_, _057532_, _057533_, _057534_, _057535_, _057536_, _057537_, _057538_, _057539_, _057540_, _057541_, _057542_, _057543_, _057544_, _057545_, _057546_, _057547_, _057548_, _057549_, _057550_, _057551_, _057552_, _057553_, _057554_, _057555_, _057556_, _057557_, _057558_, _057559_, _057560_, _057561_, _057562_, _057563_, _057564_, _057565_, _057566_, _057567_, _057568_, _057569_, _057570_, _057571_, _057572_, _057573_, _057574_, _057575_, _057576_, _057577_, _057578_, _057579_, _057580_, _057581_, _057582_, _057583_, _057584_, _057585_, _057586_, _057587_, _057588_, _057589_, _057590_, _057591_, _057592_, _057593_, _057594_, _057595_, _057596_, _057597_, _057598_, _057599_, _057600_, _057601_, _057602_, _057603_, _057604_, _057605_, _057606_, _057607_, _057608_, _057609_, _057610_, _057611_, _057612_, _057613_, _057614_, _057615_, _057616_, _057617_, _057618_, _057619_, _057620_, _057621_, _057622_, _057623_, _057624_, _057625_, _057626_, _057627_, _057628_, _057629_, _057630_, _057631_, _057632_, _057633_, _057634_, _057635_, _057636_, _057637_, _057638_, _057639_, _057640_, _057641_, _057642_, _057643_, _057644_, _057645_, _057646_, _057647_, _057648_, _057649_, _057650_, _057651_, _057652_, _057653_, _057654_, _057655_, _057656_, _057657_, _057658_, _057659_, _057660_, _057661_, _057662_, _057663_, _057664_, _057665_, _057666_, _057667_, _057668_, _057669_, _057670_, _057671_, _057672_, _057673_, _057674_, _057675_, _057676_, _057677_, _057678_, _057679_, _057680_, _057681_, _057682_, _057683_, _057684_, _057685_, _057686_, _057687_, _057688_, _057689_, _057690_, _057691_, _057692_, _057693_, _057694_, _057695_, _057696_, _057697_, _057698_, _057699_, _057700_, _057701_, _057702_, _057703_, _057704_, _057705_, _057706_, _057707_, _057708_, _057709_, _057710_, _057711_, _057712_, _057713_, _057714_, _057715_, _057716_, _057717_, _057718_, _057719_, _057720_, _057721_, _057722_, _057723_, _057724_, _057725_, _057726_, _057727_, _057728_, _057729_, _057730_, _057731_, _057732_, _057733_, _057734_, _057735_, _057736_, _057737_, _057738_, _057739_, _057740_, _057741_, _057742_, _057743_, _057744_, _057745_, _057746_, _057747_, _057748_, _057749_, _057750_, _057751_, _057752_, _057753_, _057754_, _057755_, _057756_, _057757_, _057758_, _057759_, _057760_, _057761_, _057762_, _057763_, _057764_, _057765_, _057766_, _057767_, _057768_, _057769_, _057770_, _057771_, _057772_, _057773_, _057774_, _057775_, _057776_, _057777_, _057778_, _057779_, _057780_, _057781_, _057782_, _057783_, _057784_, _057785_, _057786_, _057787_, _057788_, _057789_, _057790_, _057791_, _057792_, _057793_, _057794_, _057795_, _057796_, _057797_, _057798_, _057799_, _057800_, _057801_, _057802_, _057803_, _057804_, _057805_, _057806_, _057807_, _057808_, _057809_, _057810_, _057811_, _057812_, _057813_, _057814_, _057815_, _057816_, _057817_, _057818_, _057819_, _057820_, _057821_, _057822_, _057823_, _057824_, _057825_, _057826_, _057827_, _057828_, _057829_, _057830_, _057831_, _057832_, _057833_, _057834_, _057835_, _057836_, _057837_, _057838_, _057839_, _057840_, _057841_, _057842_, _057843_, _057844_, _057845_, _057846_, _057847_, _057848_, _057849_, _057850_, _057851_, _057852_, _057853_, _057854_, _057855_, _057856_, _057857_, _057858_, _057859_, _057860_, _057861_, _057862_, _057863_, _057864_, _057865_, _057866_, _057867_, _057868_, _057869_, _057870_, _057871_, _057872_, _057873_, _057874_, _057875_, _057876_, _057877_, _057878_, _057879_, _057880_, _057881_, _057882_, _057883_, _057884_, _057885_, _057886_, _057887_, _057888_, _057889_, _057890_, _057891_, _057892_, _057893_, _057894_, _057895_, _057896_, _057897_, _057898_, _057899_, _057900_, _057901_, _057902_, _057903_, _057904_, _057905_, _057906_, _057907_, _057908_, _057909_, _057910_, _057911_, _057912_, _057913_, _057914_, _057915_, _057916_, _057917_, _057918_, _057919_, _057920_, _057921_, _057922_, _057923_, _057924_, _057925_, _057926_, _057927_, _057928_, _057929_, _057930_, _057931_, _057932_, _057933_, _057934_, _057935_, _057936_, _057937_, _057938_, _057939_, _057940_, _057941_, _057942_, _057943_, _057944_, _057945_, _057946_, _057947_, _057948_, _057949_, _057950_, _057951_, _057952_, _057953_, _057954_, _057955_, _057956_, _057957_, _057958_, _057959_, _057960_, _057961_, _057962_, _057963_, _057964_, _057965_, _057966_, _057967_, _057968_, _057969_, _057970_, _057971_, _057972_, _057973_, _057974_, _057975_, _057976_, _057977_, _057978_, _057979_, _057980_, _057981_, _057982_, _057983_, _057984_, _057985_, _057986_, _057987_, _057988_, _057989_, _057990_, _057991_, _057992_, _057993_, _057994_, _057995_, _057996_, _057997_, _057998_, _057999_, _058000_, _058001_, _058002_, _058003_, _058004_, _058005_, _058006_, _058007_, _058008_, _058009_, _058010_, _058011_, _058012_, _058013_, _058014_, _058015_, _058016_, _058017_, _058018_, _058019_, _058020_, _058021_, _058022_, _058023_, _058024_, _058025_, _058026_, _058027_, _058028_, _058029_, _058030_, _058031_, _058032_, _058033_, _058034_, _058035_, _058036_, _058037_, _058038_, _058039_, _058040_, _058041_, _058042_, _058043_, _058044_, _058045_, _058046_, _058047_, _058048_, _058049_, _058050_, _058051_, _058052_, _058053_, _058054_, _058055_, _058056_, _058057_, _058058_, _058059_, _058060_, _058061_, _058062_, _058063_, _058064_, _058065_, _058066_, _058067_, _058068_, _058069_, _058070_, _058071_, _058072_, _058073_, _058074_, _058075_, _058076_, _058077_, _058078_, _058079_, _058080_, _058081_, _058082_, _058083_, _058084_, _058085_, _058086_, _058087_, _058088_, _058089_, _058090_, _058091_, _058092_, _058093_, _058094_, _058095_, _058096_, _058097_, _058098_, _058099_, _058100_, _058101_, _058102_, _058103_, _058104_, _058105_, _058106_, _058107_, _058108_, _058109_, _058110_, _058111_, _058112_, _058113_, _058114_, _058115_, _058116_, _058117_, _058118_, _058119_, _058120_, _058121_, _058122_, _058123_, _058124_, _058125_, _058126_, _058127_, _058128_, _058129_, _058130_, _058131_, _058132_, _058133_, _058134_, _058135_, _058136_, _058137_, _058138_, _058139_, _058140_, _058141_, _058142_, _058143_, _058144_, _058145_, _058146_, _058147_, _058148_, _058149_, _058150_, _058151_, _058152_, _058153_, _058154_, _058155_, _058156_, _058157_, _058158_, _058159_, _058160_, _058161_, _058162_, _058163_, _058164_, _058165_, _058166_, _058167_, _058168_, _058169_, _058170_, _058171_, _058172_, _058173_, _058174_, _058175_, _058176_, _058177_, _058178_, _058179_, _058180_, _058181_, _058182_, _058183_, _058184_, _058185_, _058186_, _058187_, _058188_, _058189_, _058190_, _058191_, _058192_, _058193_, _058194_, _058195_, _058196_, _058197_, _058198_, _058199_, _058200_, _058201_, _058202_, _058203_, _058204_, _058205_, _058206_, _058207_, _058208_, _058209_, _058210_, _058211_, _058212_, _058213_, _058214_, _058215_, _058216_, _058217_, _058218_, _058219_, _058220_, _058221_, _058222_, _058223_, _058224_, _058225_, _058226_, _058227_, _058228_, _058229_, _058230_, _058231_, _058232_, _058233_, _058234_, _058235_, _058236_, _058237_, _058238_, _058239_, _058240_, _058241_, _058242_, _058243_, _058244_, _058245_, _058246_, _058247_, _058248_, _058249_, _058250_, _058251_, _058252_, _058253_, _058254_, _058255_, _058256_, _058257_, _058258_, _058259_, _058260_, _058261_, _058262_, _058263_, _058264_, _058265_, _058266_, _058267_, _058268_, _058269_, _058270_, _058271_, _058272_, _058273_, _058274_, _058275_, _058276_, _058277_, _058278_, _058279_, _058280_, _058281_, _058282_, _058283_, _058284_, _058285_, _058286_, _058287_, _058288_, _058289_, _058290_, _058291_, _058292_, _058293_, _058294_, _058295_, _058296_, _058297_, _058298_, _058299_, _058300_, _058301_, _058302_, _058303_, _058304_, _058305_, _058306_, _058307_, _058308_, _058309_, _058310_, _058311_, _058312_, _058313_, _058314_, _058315_, _058316_, _058317_, _058318_, _058319_, _058320_, _058321_, _058322_, _058323_, _058324_, _058325_, _058326_, _058327_, _058328_, _058329_, _058330_, _058331_, _058332_, _058333_, _058334_, _058335_, _058336_, _058337_, _058338_, _058339_, _058340_, _058341_, _058342_, _058343_, _058344_, _058345_, _058346_, _058347_, _058348_, _058349_, _058350_, _058351_, _058352_, _058353_, _058354_, _058355_, _058356_, _058357_, _058358_, _058359_, _058360_, _058361_, _058362_, _058363_, _058364_, _058365_, _058366_, _058367_, _058368_, _058369_, _058370_, _058371_, _058372_, _058373_, _058374_, _058375_, _058376_, _058377_, _058378_, _058379_, _058380_, _058381_, _058382_, _058383_, _058384_, _058385_, _058386_, _058387_, _058388_, _058389_, _058390_, _058391_, _058392_, _058393_, _058394_, _058395_, _058396_, _058397_, _058398_, _058399_, _058400_, _058401_, _058402_, _058403_, _058404_, _058405_, _058406_, _058407_, _058408_, _058409_, _058410_, _058411_, _058412_, _058413_, _058414_, _058415_, _058416_, _058417_, _058418_, _058419_, _058420_, _058421_, _058422_, _058423_, _058424_, _058425_, _058426_, _058427_, _058428_, _058429_, _058430_, _058431_, _058432_, _058433_, _058434_, _058435_, _058436_, _058437_, _058438_, _058439_, _058440_, _058441_, _058442_, _058443_, _058444_, _058445_, _058446_, _058447_, _058448_, _058449_, _058450_, _058451_, _058452_, _058453_, _058454_, _058455_, _058456_, _058457_, _058458_, _058459_, _058460_, _058461_, _058462_, _058463_, _058464_, _058465_, _058466_, _058467_, _058468_, _058469_, _058470_, _058471_, _058472_, _058473_, _058474_, _058475_, _058476_, _058477_, _058478_, _058479_, _058480_, _058481_, _058482_, _058483_, _058484_, _058485_, _058486_, _058487_, _058488_, _058489_, _058490_, _058491_, _058492_, _058493_, _058494_, _058495_, _058496_, _058497_, _058498_, _058499_, _058500_, _058501_, _058502_, _058503_, _058504_, _058505_, _058506_, _058507_, _058508_, _058509_, _058510_, _058511_, _058512_, _058513_, _058514_, _058515_, _058516_, _058517_, _058518_, _058519_, _058520_, _058521_, _058522_, _058523_, _058524_, _058525_, _058526_, _058527_, _058528_, _058529_, _058530_, _058531_, _058532_, _058533_, _058534_, _058535_, _058536_, _058537_, _058538_, _058539_, _058540_, _058541_, _058542_, _058543_, _058544_, _058545_, _058546_, _058547_, _058548_, _058549_, _058550_, _058551_, _058552_, _058553_, _058554_, _058555_, _058556_, _058557_, _058558_, _058559_, _058560_, _058561_, _058562_, _058563_, _058564_, _058565_, _058566_, _058567_, _058568_, _058569_, _058570_, _058571_, _058572_, _058573_, _058574_, _058575_, _058576_, _058577_, _058578_, _058579_, _058580_, _058581_, _058582_, _058583_, _058584_, _058585_, _058586_, _058587_, _058588_, _058589_, _058590_, _058591_, _058592_, _058593_, _058594_, _058595_, _058596_, _058597_, _058598_, _058599_, _058600_, _058601_, _058602_, _058603_, _058604_, _058605_, _058606_, _058607_, _058608_, _058609_, _058610_, _058611_, _058612_, _058613_, _058614_, _058615_, _058616_, _058617_, _058618_, _058619_, _058620_, _058621_, _058622_, _058623_, _058624_, _058625_, _058626_, _058627_, _058628_, _058629_, _058630_, _058631_, _058632_, _058633_, _058634_, _058635_, _058636_, _058637_, _058638_, _058639_, _058640_, _058641_, _058642_, _058643_, _058644_, _058645_, _058646_, _058647_, _058648_, _058649_, _058650_, _058651_, _058652_, _058653_, _058654_, _058655_, _058656_, _058657_, _058658_, _058659_, _058660_, _058661_, _058662_, _058663_, _058664_, _058665_, _058666_, _058667_, _058668_, _058669_, _058670_, _058671_, _058672_, _058673_, _058674_, _058675_, _058676_, _058677_, _058678_, _058679_, _058680_, _058681_, _058682_, _058683_, _058684_, _058685_, _058686_, _058687_, _058688_, _058689_, _058690_, _058691_, _058692_, _058693_, _058694_, _058695_, _058696_, _058697_, _058698_, _058699_, _058700_, _058701_, _058702_, _058703_, _058704_, _058705_, _058706_, _058707_, _058708_, _058709_, _058710_, _058711_, _058712_, _058713_, _058714_, _058715_, _058716_, _058717_, _058718_, _058719_, _058720_, _058721_, _058722_, _058723_, _058724_, _058725_, _058726_, _058727_, _058728_, _058729_, _058730_, _058731_, _058732_, _058733_, _058734_, _058735_, _058736_, _058737_, _058738_, _058739_, _058740_, _058741_, _058742_, _058743_, _058744_, _058745_, _058746_, _058747_, _058748_, _058749_, _058750_, _058751_, _058752_, _058753_, _058754_, _058755_, _058756_, _058757_, _058758_, _058759_, _058760_, _058761_, _058762_, _058763_, _058764_, _058765_, _058766_, _058767_, _058768_, _058769_, _058770_, _058771_, _058772_, _058773_, _058774_, _058775_, _058776_, _058777_, _058778_, _058779_, _058780_, _058781_, _058782_, _058783_, _058784_, _058785_, _058786_, _058787_, _058788_, _058789_, _058790_, _058791_, _058792_, _058793_, _058794_, _058795_, _058796_, _058797_, _058798_, _058799_, _058800_, _058801_, _058802_, _058803_, _058804_, _058805_, _058806_, _058807_, _058808_, _058809_, _058810_, _058811_, _058812_, _058813_, _058814_, _058815_, _058816_, _058817_, _058818_, _058819_, _058820_, _058821_, _058822_, _058823_, _058824_, _058825_, _058826_, _058827_, _058828_, _058829_, _058830_, _058831_, _058832_, _058833_, _058834_, _058835_, _058836_, _058837_, _058838_, _058839_, _058840_, _058841_, _058842_, _058843_, _058844_, _058845_, _058846_, _058847_, _058848_, _058849_, _058850_, _058851_, _058852_, _058853_, _058854_, _058855_, _058856_, _058857_, _058858_, _058859_, _058860_, _058861_, _058862_, _058863_, _058864_, _058865_, _058866_, _058867_, _058868_, _058869_, _058870_, _058871_, _058872_, _058873_, _058874_, _058875_, _058876_, _058877_, _058878_, _058879_, _058880_, _058881_, _058882_, _058883_, _058884_, _058885_, _058886_, _058887_, _058888_, _058889_, _058890_, _058891_, _058892_, _058893_, _058894_, _058895_, _058896_, _058897_, _058898_, _058899_, _058900_, _058901_, _058902_, _058903_, _058904_, _058905_, _058906_, _058907_, _058908_, _058909_, _058910_, _058911_, _058912_, _058913_, _058914_, _058915_, _058916_, _058917_, _058918_, _058919_, _058920_, _058921_, _058922_, _058923_, _058924_, _058925_, _058926_, _058927_, _058928_, _058929_, _058930_, _058931_, _058932_, _058933_, _058934_, _058935_, _058936_, _058937_, _058938_, _058939_, _058940_, _058941_, _058942_, _058943_, _058944_, _058945_, _058946_, _058947_, _058948_, _058949_, _058950_, _058951_, _058952_, _058953_, _058954_, _058955_, _058956_, _058957_, _058958_, _058959_, _058960_, _058961_, _058962_, _058963_, _058964_, _058965_, _058966_, _058967_, _058968_, _058969_, _058970_, _058971_, _058972_, _058973_, _058974_, _058975_, _058976_, _058977_, _058978_, _058979_, _058980_, _058981_, _058982_, _058983_, _058984_, _058985_, _058986_, _058987_, _058988_, _058989_, _058990_, _058991_, _058992_, _058993_, _058994_, _058995_, _058996_, _058997_, _058998_, _058999_, _059000_, _059001_, _059002_, _059003_, _059004_, _059005_, _059006_, _059007_, _059008_, _059009_, _059010_, _059011_, _059012_, _059013_, _059014_, _059015_, _059016_, _059017_, _059018_, _059019_, _059020_, _059021_, _059022_, _059023_, _059024_, _059025_, _059026_, _059027_, _059028_, _059029_, _059030_, _059031_, _059032_, _059033_, _059034_, _059035_, _059036_, _059037_, _059038_, _059039_, _059040_, _059041_, _059042_, _059043_, _059044_, _059045_, _059046_, _059047_, _059048_, _059049_, _059050_, _059051_, _059052_, _059053_, _059054_, _059055_, _059056_, _059057_, _059058_, _059059_, _059060_, _059061_, _059062_, _059063_, _059064_, _059065_, _059066_, _059067_, _059068_, _059069_, _059070_, _059071_, _059072_, _059073_, _059074_, _059075_, _059076_, _059077_, _059078_, _059079_, _059080_, _059081_, _059082_, _059083_, _059084_, _059085_, _059086_, _059087_, _059088_, _059089_, _059090_, _059091_, _059092_, _059093_, _059094_, _059095_, _059096_, _059097_, _059098_, _059099_, _059100_, _059101_, _059102_, _059103_, _059104_, _059105_, _059106_, _059107_, _059108_, _059109_, _059110_, _059111_, _059112_, _059113_, _059114_, _059115_, _059116_, _059117_, _059118_, _059119_, _059120_, _059121_, _059122_, _059123_, _059124_, _059125_, _059126_, _059127_, _059128_, _059129_, _059130_, _059131_, _059132_, _059133_, _059134_, _059135_, _059136_, _059137_, _059138_, _059139_, _059140_, _059141_, _059142_, _059143_, _059144_, _059145_, _059146_, _059147_, _059148_, _059149_, _059150_, _059151_, _059152_, _059153_, _059154_, _059155_, _059156_, _059157_, _059158_, _059159_, _059160_, _059161_, _059162_, _059163_, _059164_, _059165_, _059166_, _059167_, _059168_, _059169_, _059170_, _059171_, _059172_, _059173_, _059174_, _059175_, _059176_, _059177_, _059178_, _059179_, _059180_, _059181_, _059182_, _059183_, _059184_, _059185_, _059186_, _059187_, _059188_, _059189_, _059190_, _059191_, _059192_, _059193_, _059194_, _059195_, _059196_, _059197_, _059198_, _059199_, _059200_, _059201_, _059202_, _059203_, _059204_, _059205_, _059206_, _059207_, _059208_, _059209_, _059210_, _059211_, _059212_, _059213_, _059214_, _059215_, _059216_, _059217_, _059218_, _059219_, _059220_, _059221_, _059222_, _059223_, _059224_, _059225_, _059226_, _059227_, _059228_, _059229_, _059230_, _059231_, _059232_, _059233_, _059234_, _059235_, _059236_, _059237_, _059238_, _059239_, _059240_, _059241_, _059242_, _059243_, _059244_, _059245_, _059246_, _059247_, _059248_, _059249_, _059250_, _059251_, _059252_, _059253_, _059254_, _059255_, _059256_, _059257_, _059258_, _059259_, _059260_, _059261_, _059262_, _059263_, _059264_, _059265_, _059266_, _059267_, _059268_, _059269_, _059270_, _059271_, _059272_, _059273_, _059274_, _059275_, _059276_, _059277_, _059278_, _059279_, _059280_, _059281_, _059282_, _059283_, _059284_, _059285_, _059286_, _059287_, _059288_, _059289_, _059290_, _059291_, _059292_, _059293_, _059294_, _059295_, _059296_, _059297_, _059298_, _059299_, _059300_, _059301_, _059302_, _059303_, _059304_, _059305_, _059306_, _059307_, _059308_, _059309_, _059310_, _059311_, _059312_, _059313_, _059314_, _059315_, _059316_, _059317_, _059318_, _059319_, _059320_, _059321_, _059322_, _059323_, _059324_, _059325_, _059326_, _059327_, _059328_, _059329_, _059330_, _059331_, _059332_, _059333_, _059334_, _059335_, _059336_, _059337_, _059338_, _059339_, _059340_, _059341_, _059342_, _059343_, _059344_, _059345_, _059346_, _059347_, _059348_, _059349_, _059350_, _059351_, _059352_, _059353_, _059354_, _059355_, _059356_, _059357_, _059358_, _059359_, _059360_, _059361_, _059362_, _059363_, _059364_, _059365_, _059366_, _059367_, _059368_, _059369_, _059370_, _059371_, _059372_, _059373_, _059374_, _059375_, _059376_, _059377_, _059378_, _059379_, _059380_, _059381_, _059382_, _059383_, _059384_, _059385_, _059386_, _059387_, _059388_, _059389_, _059390_, _059391_, _059392_, _059393_, _059394_, _059395_, _059396_, _059397_, _059398_, _059399_, _059400_, _059401_, _059402_, _059403_, _059404_, _059405_, _059406_, _059407_, _059408_, _059409_, _059410_, _059411_, _059412_, _059413_, _059414_, _059415_, _059416_, _059417_, _059418_, _059419_, _059420_, _059421_, _059422_, _059423_, _059424_, _059425_, _059426_, _059427_, _059428_, _059429_, _059430_, _059431_, _059432_, _059433_, _059434_, _059435_, _059436_, _059437_, _059438_, _059439_, _059440_, _059441_, _059442_, _059443_, _059444_, _059445_, _059446_, _059447_, _059448_, _059449_, _059450_, _059451_, _059452_, _059453_, _059454_, _059455_, _059456_, _059457_, _059458_, _059459_, _059460_, _059461_, _059462_, _059463_, _059464_, _059465_, _059466_, _059467_, _059468_, _059469_, _059470_, _059471_, _059472_, _059473_, _059474_, _059475_, _059476_, _059477_, _059478_, _059479_, _059480_, _059481_, _059482_, _059483_, _059484_, _059485_, _059486_, _059487_, _059488_, _059489_, _059490_, _059491_, _059492_, _059493_, _059494_, _059495_, _059496_, _059497_, _059498_, _059499_, _059500_, _059501_, _059502_, _059503_, _059504_, _059505_, _059506_, _059507_, _059508_, _059509_, _059510_, _059511_, _059512_, _059513_, _059514_, _059515_, _059516_, _059517_, _059518_, _059519_, _059520_, _059521_, _059522_, _059523_, _059524_, _059525_, _059526_, _059527_, _059528_, _059529_, _059530_, _059531_, _059532_, _059533_, _059534_, _059535_, _059536_, _059537_, _059538_, _059539_, _059540_, _059541_, _059542_, _059543_, _059544_, _059545_, _059546_, _059547_, _059548_, _059549_, _059550_, _059551_, _059552_, _059553_, _059554_, _059555_, _059556_, _059557_, _059558_, _059559_, _059560_, _059561_, _059562_, _059563_, _059564_, _059565_, _059566_, _059567_, _059568_, _059569_, _059570_, _059571_, _059572_, _059573_, _059574_, _059575_, _059576_, _059577_, _059578_, _059579_, _059580_, _059581_, _059582_, _059583_, _059584_, _059585_, _059586_, _059587_, _059588_, _059589_, _059590_, _059591_, _059592_, _059593_, _059594_, _059595_, _059596_, _059597_, _059598_, _059599_, _059600_, _059601_, _059602_, _059603_, _059604_, _059605_, _059606_, _059607_, _059608_, _059609_, _059610_, _059611_, _059612_, _059613_, _059614_, _059615_, _059616_, _059617_, _059618_, _059619_, _059620_, _059621_, _059622_, _059623_, _059624_, _059625_, _059626_, _059627_, _059628_, _059629_, _059630_, _059631_, _059632_, _059633_, _059634_, _059635_, _059636_, _059637_, _059638_, _059639_, _059640_, _059641_, _059642_, _059643_, _059644_, _059645_, _059646_, _059647_, _059648_, _059649_, _059650_, _059651_, _059652_, _059653_, _059654_, _059655_, _059656_, _059657_, _059658_, _059659_, _059660_, _059661_, _059662_, _059663_, _059664_, _059665_, _059666_, _059667_, _059668_, _059669_, _059670_, _059671_, _059672_, _059673_, _059674_, _059675_, _059676_, _059677_, _059678_, _059679_, _059680_, _059681_, _059682_, _059683_, _059684_, _059685_, _059686_, _059687_, _059688_, _059689_, _059690_, _059691_, _059692_, _059693_, _059694_, _059695_, _059696_, _059697_, _059698_, _059699_, _059700_, _059701_, _059702_, _059703_, _059704_, _059705_, _059706_, _059707_, _059708_, _059709_, _059710_, _059711_, _059712_, _059713_, _059714_, _059715_, _059716_, _059717_, _059718_, _059719_, _059720_, _059721_, _059722_, _059723_, _059724_, _059725_, _059726_, _059727_, _059728_, _059729_, _059730_, _059731_, _059732_, _059733_, _059734_, _059735_, _059736_, _059737_, _059738_, _059739_, _059740_, _059741_, _059742_, _059743_, _059744_, _059745_, _059746_, _059747_, _059748_, _059749_, _059750_, _059751_, _059752_, _059753_, _059754_, _059755_, _059756_, _059757_, _059758_, _059759_, _059760_, _059761_, _059762_, _059763_, _059764_, _059765_, _059766_, _059767_, _059768_, _059769_, _059770_, _059771_, _059772_, _059773_, _059774_, _059775_, _059776_, _059777_, _059778_, _059779_, _059780_, _059781_, _059782_, _059783_, _059784_, _059785_, _059786_, _059787_, _059788_, _059789_, _059790_, _059791_, _059792_, _059793_, _059794_, _059795_, _059796_, _059797_, _059798_, _059799_, _059800_, _059801_, _059802_, _059803_, _059804_, _059805_, _059806_, _059807_, _059808_, _059809_, _059810_, _059811_, _059812_, _059813_, _059814_, _059815_, _059816_, _059817_, _059818_, _059819_, _059820_, _059821_, _059822_, _059823_, _059824_, _059825_, _059826_, _059827_, _059828_, _059829_, _059830_, _059831_, _059832_, _059833_, _059834_, _059835_, _059836_, _059837_, _059838_, _059839_, _059840_, _059841_, _059842_, _059843_, _059844_, _059845_, _059846_, _059847_, _059848_, _059849_, _059850_, _059851_, _059852_, _059853_, _059854_, _059855_, _059856_, _059857_, _059858_, _059859_, _059860_, _059861_, _059862_, _059863_, _059864_, _059865_, _059866_, _059867_, _059868_, _059869_, _059870_, _059871_, _059872_, _059873_, _059874_, _059875_, _059876_, _059877_, _059878_, _059879_, _059880_, _059881_, _059882_, _059883_, _059884_, _059885_, _059886_, _059887_, _059888_, _059889_, _059890_, _059891_, _059892_, _059893_, _059894_, _059895_, _059896_, _059897_, _059898_, _059899_, _059900_, _059901_, _059902_, _059903_, _059904_, _059905_, _059906_, _059907_, _059908_, _059909_, _059910_, _059911_, _059912_, _059913_, _059914_, _059915_, _059916_, _059917_, _059918_, _059919_, _059920_, _059921_, _059922_, _059923_, _059924_, _059925_, _059926_, _059927_, _059928_, _059929_, _059930_, _059931_, _059932_, _059933_, _059934_, _059935_, _059936_, _059937_, _059938_, _059939_, _059940_, _059941_, _059942_, _059943_, _059944_, _059945_, _059946_, _059947_, _059948_, _059949_, _059950_, _059951_, _059952_, _059953_, _059954_, _059955_, _059956_, _059957_, _059958_, _059959_, _059960_, _059961_, _059962_, _059963_, _059964_, _059965_, _059966_, _059967_, _059968_, _059969_, _059970_, _059971_, _059972_, _059973_, _059974_, _059975_, _059976_, _059977_, _059978_, _059979_, _059980_, _059981_, _059982_, _059983_, _059984_, _059985_, _059986_, _059987_, _059988_, _059989_, _059990_, _059991_, _059992_, _059993_, _059994_, _059995_, _059996_, _059997_, _059998_, _059999_, _060000_, _060001_, _060002_, _060003_, _060004_, _060005_, _060006_, _060007_, _060008_, _060009_, _060010_, _060011_, _060012_, _060013_, _060014_, _060015_, _060016_, _060017_, _060018_, _060019_, _060020_, _060021_, _060022_, _060023_, _060024_, _060025_, _060026_, _060027_, _060028_, _060029_, _060030_, _060031_, _060032_, _060033_, _060034_, _060035_, _060036_, _060037_, _060038_, _060039_, _060040_, _060041_, _060042_, _060043_, _060044_, _060045_, _060046_, _060047_, _060048_, _060049_, _060050_, _060051_, _060052_, _060053_, _060054_, _060055_, _060056_, _060057_, _060058_, _060059_, _060060_, _060061_, _060062_, _060063_, _060064_, _060065_, _060066_, _060067_, _060068_, _060069_, _060070_, _060071_, _060072_, _060073_, _060074_, _060075_, _060076_, _060077_, _060078_, _060079_, _060080_, _060081_, _060082_, _060083_, _060084_, _060085_, _060086_, _060087_, _060088_, _060089_, _060090_, _060091_, _060092_, _060093_, _060094_, _060095_, _060096_, _060097_, _060098_, _060099_, _060100_, _060101_, _060102_, _060103_, _060104_, _060105_, _060106_, _060107_, _060108_, _060109_, _060110_, _060111_, _060112_, _060113_, _060114_, _060115_, _060116_, _060117_, _060118_, _060119_, _060120_, _060121_, _060122_, _060123_, _060124_, _060125_, _060126_, _060127_, _060128_, _060129_, _060130_, _060131_, _060132_, _060133_, _060134_, _060135_, _060136_, _060137_, _060138_, _060139_, _060140_, _060141_, _060142_, _060143_, _060144_, _060145_, _060146_, _060147_, _060148_, _060149_, _060150_, _060151_, _060152_, _060153_, _060154_, _060155_, _060156_, _060157_, _060158_, _060159_, _060160_, _060161_, _060162_, _060163_, _060164_, _060165_, _060166_, _060167_, _060168_, _060169_, _060170_, _060171_, _060172_, _060173_, _060174_, _060175_, _060176_, _060177_, _060178_, _060179_, _060180_, _060181_, _060182_, _060183_, _060184_, _060185_, _060186_, _060187_, _060188_, _060189_, _060190_, _060191_, _060192_, _060193_, _060194_, _060195_, _060196_, _060197_, _060198_, _060199_, _060200_, _060201_, _060202_, _060203_, _060204_, _060205_, _060206_, _060207_, _060208_, _060209_, _060210_, _060211_, _060212_, _060213_, _060214_, _060215_, _060216_, _060217_, _060218_, _060219_, _060220_, _060221_, _060222_, _060223_, _060224_, _060225_, _060226_, _060227_, _060228_, _060229_, _060230_, _060231_, _060232_, _060233_, _060234_, _060235_, _060236_, _060237_, _060238_, _060239_, _060240_, _060241_, _060242_, _060243_, _060244_, _060245_, _060246_, _060247_, _060248_, _060249_, _060250_, _060251_, _060252_, _060253_, _060254_, _060255_, _060256_, _060257_, _060258_, _060259_, _060260_, _060261_, _060262_, _060263_, _060264_, _060265_, _060266_, _060267_, _060268_, _060269_, _060270_, _060271_, _060272_, _060273_, _060274_, _060275_, _060276_, _060277_, _060278_, _060279_, _060280_, _060281_, _060282_, _060283_, _060284_, _060285_, _060286_, _060287_, _060288_, _060289_, _060290_, _060291_, _060292_, _060293_, _060294_, _060295_, _060296_, _060297_, _060298_, _060299_, _060300_, _060301_, _060302_, _060303_, _060304_, _060305_, _060306_, _060307_, _060308_, _060309_, _060310_, _060311_, _060312_, _060313_, _060314_, _060315_, _060316_, _060317_, _060318_, _060319_, _060320_, _060321_, _060322_, _060323_, _060324_, _060325_, _060326_, _060327_, _060328_, _060329_, _060330_, _060331_, _060332_, _060333_, _060334_, _060335_, _060336_, _060337_, _060338_, _060339_, _060340_, _060341_, _060342_, _060343_, _060344_, _060345_, _060346_, _060347_, _060348_, _060349_, _060350_, _060351_, _060352_, _060353_, _060354_, _060355_, _060356_, _060357_, _060358_, _060359_, _060360_, _060361_, _060362_, _060363_, _060364_, _060365_, _060366_, _060367_, _060368_, _060369_, _060370_, _060371_, _060372_, _060373_, _060374_, _060375_, _060376_, _060377_, _060378_, _060379_, _060380_, _060381_, _060382_, _060383_, _060384_, _060385_, _060386_, _060387_, _060388_, _060389_, _060390_, _060391_, _060392_, _060393_, _060394_, _060395_, _060396_, _060397_, _060398_, _060399_, _060400_, _060401_, _060402_, _060403_, _060404_, _060405_, _060406_, _060407_, _060408_, _060409_, _060410_, _060411_, _060412_, _060413_, _060414_, _060415_, _060416_, _060417_, _060418_, _060419_, _060420_, _060421_, _060422_, _060423_, _060424_, _060425_, _060426_, _060427_, _060428_, _060429_, _060430_, _060431_, _060432_, _060433_, _060434_, _060435_, _060436_, _060437_, _060438_, _060439_, _060440_, _060441_, _060442_, _060443_, _060444_, _060445_, _060446_, _060447_, _060448_, _060449_, _060450_, _060451_, _060452_, _060453_, _060454_, _060455_, _060456_, _060457_, _060458_, _060459_, _060460_, _060461_, _060462_, _060463_, _060464_, _060465_, _060466_, _060467_, _060468_, _060469_, _060470_, _060471_, _060472_, _060473_, _060474_, _060475_, _060476_, _060477_, _060478_, _060479_, _060480_, _060481_, _060482_, _060483_, _060484_, _060485_, _060486_, _060487_, _060488_, _060489_, _060490_, _060491_, _060492_, _060493_, _060494_, _060495_, _060496_, _060497_, _060498_, _060499_, _060500_, _060501_, _060502_, _060503_, _060504_, _060505_, _060506_, _060507_, _060508_, _060509_, _060510_, _060511_, _060512_, _060513_, _060514_, _060515_, _060516_, _060517_, _060518_, _060519_, _060520_, _060521_, _060522_, _060523_, _060524_, _060525_, _060526_, _060527_, _060528_, _060529_, _060530_, _060531_, _060532_, _060533_, _060534_, _060535_, _060536_, _060537_, _060538_, _060539_, _060540_, _060541_, _060542_, _060543_, _060544_, _060545_, _060546_, _060547_, _060548_, _060549_, _060550_, _060551_, _060552_, _060553_, _060554_, _060555_, _060556_, _060557_, _060558_, _060559_, _060560_, _060561_, _060562_, _060563_, _060564_, _060565_, _060566_, _060567_, _060568_, _060569_, _060570_, _060571_, _060572_, _060573_, _060574_, _060575_, _060576_, _060577_, _060578_, _060579_, _060580_, _060581_, _060582_, _060583_, _060584_, _060585_, _060586_, _060587_, _060588_, _060589_, _060590_, _060591_, _060592_, _060593_, _060594_, _060595_, _060596_, _060597_, _060598_, _060599_, _060600_, _060601_, _060602_, _060603_, _060604_, _060605_, _060606_, _060607_, _060608_, _060609_, _060610_, _060611_, _060612_, _060613_, _060614_, _060615_, _060616_, _060617_, _060618_, _060619_, _060620_, _060621_, _060622_, _060623_, _060624_, _060625_, _060626_, _060627_, _060628_, _060629_, _060630_, _060631_, _060632_, _060633_, _060634_, _060635_, _060636_, _060637_, _060638_, _060639_, _060640_, _060641_, _060642_, _060643_, _060644_, _060645_, _060646_, _060647_, _060648_, _060649_, _060650_, _060651_, _060652_, _060653_, _060654_, _060655_, _060656_, _060657_, _060658_, _060659_, _060660_, _060661_, _060662_, _060663_, _060664_, _060665_, _060666_, _060667_, _060668_, _060669_, _060670_, _060671_, _060672_, _060673_, _060674_, _060675_, _060676_, _060677_, _060678_, _060679_, _060680_, _060681_, _060682_, _060683_, _060684_, _060685_, _060686_, _060687_, _060688_, _060689_, _060690_, _060691_, _060692_, _060693_, _060694_, _060695_, _060696_, _060697_, _060698_, _060699_, _060700_, _060701_, _060702_, _060703_, _060704_, _060705_, _060706_, _060707_, _060708_, _060709_, _060710_, _060711_, _060712_, _060713_, _060714_, _060715_, _060716_, _060717_, _060718_, _060719_, _060720_, _060721_, _060722_, _060723_, _060724_, _060725_, _060726_, _060727_, _060728_, _060729_, _060730_, _060731_, _060732_, _060733_, _060734_, _060735_, _060736_, _060737_, _060738_, _060739_, _060740_, _060741_, _060742_, _060743_, _060744_, _060745_, _060746_, _060747_, _060748_, _060749_, _060750_, _060751_, _060752_, _060753_, _060754_, _060755_, _060756_, _060757_, _060758_, _060759_, _060760_, _060761_, _060762_, _060763_, _060764_, _060765_, _060766_, _060767_, _060768_, _060769_, _060770_, _060771_, _060772_, _060773_, _060774_, _060775_, _060776_, _060777_, _060778_, _060779_, _060780_, _060781_, _060782_, _060783_, _060784_, _060785_, _060786_, _060787_, _060788_, _060789_, _060790_, _060791_, _060792_, _060793_, _060794_, _060795_, _060796_, _060797_, _060798_, _060799_, _060800_, _060801_, _060802_, _060803_, _060804_, _060805_, _060806_, _060807_, _060808_, _060809_, _060810_, _060811_, _060812_, _060813_, _060814_, _060815_, _060816_, _060817_, _060818_, _060819_, _060820_, _060821_, _060822_, _060823_, _060824_, _060825_, _060826_, _060827_, _060828_, _060829_, _060830_, _060831_, _060832_, _060833_, _060834_, _060835_, _060836_, _060837_, _060838_, _060839_, _060840_, _060841_, _060842_, _060843_, _060844_, _060845_, _060846_, _060847_, _060848_, _060849_, _060850_, _060851_, _060852_, _060853_, _060854_, _060855_, _060856_, _060857_, _060858_, _060859_, _060860_, _060861_, _060862_, _060863_, _060864_, _060865_, _060866_, _060867_, _060868_, _060869_, _060870_, _060871_, _060872_, _060873_, _060874_, _060875_, _060876_, _060877_, _060878_, _060879_, _060880_, _060881_, _060882_, _060883_, _060884_, _060885_, _060886_, _060887_, _060888_, _060889_, _060890_, _060891_, _060892_, _060893_, _060894_, _060895_, _060896_, _060897_, _060898_, _060899_, _060900_, _060901_, _060902_, _060903_, _060904_, _060905_, _060906_, _060907_, _060908_, _060909_, _060910_, _060911_, _060912_, _060913_, _060914_, _060915_, _060916_, _060917_, _060918_, _060919_, _060920_, _060921_, _060922_, _060923_, _060924_, _060925_, _060926_, _060927_, _060928_, _060929_, _060930_, _060931_, _060932_, _060933_, _060934_, _060935_, _060936_, _060937_, _060938_, _060939_, _060940_, _060941_, _060942_, _060943_, _060944_, _060945_, _060946_, _060947_, _060948_, _060949_, _060950_, _060951_, _060952_, _060953_, _060954_, _060955_, _060956_, _060957_, _060958_, _060959_, _060960_, _060961_, _060962_, _060963_, _060964_, _060965_, _060966_, _060967_, _060968_, _060969_, _060970_, _060971_, _060972_, _060973_, _060974_, _060975_, _060976_, _060977_, _060978_, _060979_, _060980_, _060981_, _060982_, _060983_, _060984_, _060985_, _060986_, _060987_, _060988_, _060989_, _060990_, _060991_, _060992_, _060993_, _060994_, _060995_, _060996_, _060997_, _060998_, _060999_, _061000_, _061001_, _061002_, _061003_, _061004_, _061005_, _061006_, _061007_, _061008_, _061009_, _061010_, _061011_, _061012_, _061013_, _061014_, _061015_, _061016_, _061017_, _061018_, _061019_, _061020_, _061021_, _061022_, _061023_, _061024_, _061025_, _061026_, _061027_, _061028_, _061029_, _061030_, _061031_, _061032_, _061033_, _061034_, _061035_, _061036_, _061037_, _061038_, _061039_, _061040_, _061041_, _061042_, _061043_, _061044_, _061045_, _061046_, _061047_, _061048_, _061049_, _061050_, _061051_, _061052_, _061053_, _061054_, _061055_, _061056_, _061057_, _061058_, _061059_, _061060_, _061061_, _061062_, _061063_, _061064_, _061065_, _061066_, _061067_, _061068_, _061069_, _061070_, _061071_, _061072_, _061073_, _061074_, _061075_, _061076_, _061077_, _061078_, _061079_, _061080_, _061081_, _061082_, _061083_, _061084_, _061085_, _061086_, _061087_, _061088_, _061089_, _061090_, _061091_, _061092_, _061093_, _061094_, _061095_, _061096_, _061097_, _061098_, _061099_, _061100_, _061101_, _061102_, _061103_, _061104_, _061105_, _061106_, _061107_, _061108_, _061109_, _061110_, _061111_, _061112_, _061113_, _061114_, _061115_, _061116_, _061117_, _061118_, _061119_, _061120_, _061121_, _061122_, _061123_, _061124_, _061125_, _061126_, _061127_, _061128_, _061129_, _061130_, _061131_, _061132_, _061133_, _061134_, _061135_, _061136_, _061137_, _061138_, _061139_, _061140_, _061141_, _061142_, _061143_, _061144_, _061145_, _061146_, _061147_, _061148_, _061149_, _061150_, _061151_, _061152_, _061153_, _061154_, _061155_, _061156_, _061157_, _061158_, _061159_, _061160_, _061161_, _061162_, _061163_, _061164_, _061165_, _061166_, _061167_, _061168_, _061169_, _061170_, _061171_, _061172_, _061173_, _061174_, _061175_, _061176_, _061177_, _061178_, _061179_, _061180_, _061181_, _061182_, _061183_, _061184_, _061185_, _061186_, _061187_, _061188_, _061189_, _061190_, _061191_, _061192_, _061193_, _061194_, _061195_, _061196_, _061197_, _061198_, _061199_, _061200_, _061201_, _061202_, _061203_, _061204_, _061205_, _061206_, _061207_, _061208_, _061209_, _061210_, _061211_, _061212_, _061213_, _061214_, _061215_, _061216_, _061217_, _061218_, _061219_, _061220_, _061221_, _061222_, _061223_, _061224_, _061225_, _061226_, _061227_, _061228_, _061229_, _061230_, _061231_, _061232_, _061233_, _061234_, _061235_, _061236_, _061237_, _061238_, _061239_, _061240_, _061241_, _061242_, _061243_, _061244_, _061245_, _061246_, _061247_, _061248_, _061249_, _061250_, _061251_, _061252_, _061253_, _061254_, _061255_, _061256_, _061257_, _061258_, _061259_, _061260_, _061261_, _061262_, _061263_, _061264_, _061265_, _061266_, _061267_, _061268_, _061269_, _061270_, _061271_, _061272_, _061273_, _061274_, _061275_, _061276_, _061277_, _061278_, _061279_, _061280_, _061281_, _061282_, _061283_, _061284_, _061285_, _061286_, _061287_, _061288_, _061289_, _061290_, _061291_, _061292_, _061293_, _061294_, _061295_, _061296_, _061297_, _061298_, _061299_, _061300_, _061301_, _061302_, _061303_, _061304_, _061305_, _061306_, _061307_, _061308_, _061309_, _061310_, _061311_, _061312_, _061313_, _061314_, _061315_, _061316_, _061317_, _061318_, _061319_, _061320_, _061321_, _061322_, _061323_, _061324_, _061325_, _061326_, _061327_, _061328_, _061329_, _061330_, _061331_, _061332_, _061333_, _061334_, _061335_, _061336_, _061337_, _061338_, _061339_, _061340_, _061341_, _061342_, _061343_, _061344_, _061345_, _061346_, _061347_, _061348_, _061349_, _061350_, _061351_, _061352_, _061353_, _061354_, _061355_, _061356_, _061357_, _061358_, _061359_, _061360_, _061361_, _061362_, _061363_, _061364_, _061365_, _061366_, _061367_, _061368_, _061369_, _061370_, _061371_, _061372_, _061373_, _061374_, _061375_, _061376_, _061377_, _061378_, _061379_, _061380_, _061381_, _061382_, _061383_, _061384_, _061385_, _061386_, _061387_, _061388_, _061389_, _061390_, _061391_, _061392_, _061393_, _061394_, _061395_, _061396_, _061397_, _061398_, _061399_, _061400_, _061401_, _061402_, _061403_, _061404_, _061405_, _061406_, _061407_, _061408_, _061409_, _061410_, _061411_, _061412_, _061413_, _061414_, _061415_, _061416_, _061417_, _061418_, _061419_, _061420_, _061421_, _061422_, _061423_, _061424_, _061425_, _061426_, _061427_, _061428_, _061429_, _061430_, _061431_, _061432_, _061433_, _061434_, _061435_, _061436_, _061437_, _061438_, _061439_, _061440_, _061441_, _061442_, _061443_, _061444_, _061445_, _061446_, _061447_, _061448_, _061449_, _061450_, _061451_, _061452_, _061453_, _061454_, _061455_, _061456_, _061457_, _061458_, _061459_, _061460_, _061461_, _061462_, _061463_, _061464_, _061465_, _061466_, _061467_, _061468_, _061469_, _061470_, _061471_, _061472_, _061473_, _061474_, _061475_, _061476_, _061477_, _061478_, _061479_, _061480_, _061481_, _061482_, _061483_, _061484_, _061485_, _061486_, _061487_, _061488_, _061489_, _061490_, _061491_, _061492_, _061493_, _061494_, _061495_, _061496_, _061497_, _061498_, _061499_, _061500_, _061501_, _061502_, _061503_, _061504_, _061505_, _061506_, _061507_, _061508_, _061509_, _061510_, _061511_, _061512_, _061513_, _061514_, _061515_, _061516_, _061517_, _061518_, _061519_, _061520_, _061521_, _061522_, _061523_, _061524_, _061525_, _061526_, _061527_, _061528_, _061529_, _061530_, _061531_, _061532_, _061533_, _061534_, _061535_, _061536_, _061537_, _061538_, _061539_, _061540_, _061541_, _061542_, _061543_, _061544_, _061545_, _061546_, _061547_, _061548_, _061549_, _061550_, _061551_, _061552_, _061553_, _061554_, _061555_, _061556_, _061557_, _061558_, _061559_, _061560_, _061561_, _061562_, _061563_, _061564_, _061565_, _061566_, _061567_, _061568_, _061569_, _061570_, _061571_, _061572_, _061573_, _061574_, _061575_, _061576_, _061577_, _061578_, _061579_, _061580_, _061581_, _061582_, _061583_, _061584_, _061585_, _061586_, _061587_, _061588_, _061589_, _061590_, _061591_, _061592_, _061593_, _061594_, _061595_, _061596_, _061597_, _061598_, _061599_, _061600_, _061601_, _061602_, _061603_, _061604_, _061605_, _061606_, _061607_, _061608_, _061609_, _061610_, _061611_, _061612_, _061613_, _061614_, _061615_, _061616_, _061617_, _061618_, _061619_, _061620_, _061621_, _061622_, _061623_, _061624_, _061625_, _061626_, _061627_, _061628_, _061629_, _061630_, _061631_, _061632_, _061633_, _061634_, _061635_, _061636_, _061637_, _061638_, _061639_, _061640_, _061641_, _061642_, _061643_, _061644_, _061645_, _061646_, _061647_, _061648_, _061649_, _061650_, _061651_, _061652_, _061653_, _061654_, _061655_, _061656_, _061657_, _061658_, _061659_, _061660_, _061661_, _061662_, _061663_, _061664_, _061665_, _061666_, _061667_, _061668_, _061669_, _061670_, _061671_, _061672_, _061673_, _061674_, _061675_, _061676_, _061677_, _061678_, _061679_, _061680_, _061681_, _061682_, _061683_, _061684_, _061685_, _061686_, _061687_, _061688_, _061689_, _061690_, _061691_, _061692_, _061693_, _061694_, _061695_, _061696_, _061697_, _061698_, _061699_, _061700_, _061701_, _061702_, _061703_, _061704_, _061705_, _061706_, _061707_, _061708_, _061709_, _061710_, _061711_, _061712_, _061713_, _061714_, _061715_, _061716_, _061717_, _061718_, _061719_, _061720_, _061721_, _061722_, _061723_, _061724_, _061725_, _061726_, _061727_, _061728_, _061729_, _061730_, _061731_, _061732_, _061733_, _061734_, _061735_, _061736_, _061737_, _061738_, _061739_, _061740_, _061741_, _061742_, _061743_, _061744_, _061745_, _061746_, _061747_, _061748_, _061749_, _061750_, _061751_, _061752_, _061753_, _061754_, _061755_, _061756_, _061757_, _061758_, _061759_, _061760_, _061761_, _061762_, _061763_, _061764_, _061765_, _061766_, _061767_, _061768_, _061769_, _061770_, _061771_, _061772_, _061773_, _061774_, _061775_, _061776_, _061777_, _061778_, _061779_, _061780_, _061781_, _061782_, _061783_, _061784_, _061785_, _061786_, _061787_, _061788_, _061789_, _061790_, _061791_, _061792_, _061793_, _061794_, _061795_, _061796_, _061797_, _061798_, _061799_, _061800_, _061801_, _061802_, _061803_, _061804_, _061805_, _061806_, _061807_, _061808_, _061809_, _061810_, _061811_, _061812_, _061813_, _061814_, _061815_, _061816_, _061817_, _061818_, _061819_, _061820_, _061821_, _061822_, _061823_, _061824_, _061825_, _061826_, _061827_, _061828_, _061829_, _061830_, _061831_, _061832_, _061833_, _061834_, _061835_, _061836_, _061837_, _061838_, _061839_, _061840_, _061841_, _061842_, _061843_, _061844_, _061845_, _061846_, _061847_, _061848_, _061849_, _061850_, _061851_, _061852_, _061853_, _061854_, _061855_, _061856_, _061857_, _061858_, _061859_, _061860_, _061861_, _061862_, _061863_, _061864_, _061865_, _061866_, _061867_, _061868_, _061869_, _061870_, _061871_, _061872_, _061873_, _061874_, _061875_, _061876_, _061877_, _061878_, _061879_, _061880_, _061881_, _061882_, _061883_, _061884_, _061885_, _061886_, _061887_, _061888_, _061889_, _061890_, _061891_, _061892_, _061893_, _061894_, _061895_, _061896_, _061897_, _061898_, _061899_, _061900_, _061901_, _061902_, _061903_, _061904_, _061905_, _061906_, _061907_, _061908_, _061909_, _061910_, _061911_, _061912_, _061913_, _061914_, _061915_, _061916_, _061917_, _061918_, _061919_, _061920_, _061921_, _061922_, _061923_, _061924_, _061925_, _061926_, _061927_, _061928_, _061929_, _061930_, _061931_, _061932_, _061933_, _061934_, _061935_, _061936_, _061937_, _061938_, _061939_, _061940_, _061941_, _061942_, _061943_, _061944_, _061945_, _061946_, _061947_, _061948_, _061949_, _061950_, _061951_, _061952_, _061953_, _061954_, _061955_, _061956_, _061957_, _061958_, _061959_, _061960_, _061961_, _061962_, _061963_, _061964_, _061965_, _061966_, _061967_, _061968_, _061969_, _061970_, _061971_, _061972_, _061973_, _061974_, _061975_, _061976_, _061977_, _061978_, _061979_, _061980_, _061981_, _061982_, _061983_, _061984_, _061985_, _061986_, _061987_, _061988_, _061989_, _061990_, _061991_, _061992_, _061993_, _061994_, _061995_, _061996_, _061997_, _061998_, _061999_, _062000_, _062001_, _062002_, _062003_, _062004_, _062005_, _062006_, _062007_, _062008_, _062009_, _062010_, _062011_, _062012_, _062013_, _062014_, _062015_, _062016_, _062017_, _062018_, _062019_, _062020_, _062021_, _062022_, _062023_, _062024_, _062025_, _062026_, _062027_, _062028_, _062029_, _062030_, _062031_, _062032_, _062033_, _062034_, _062035_, _062036_, _062037_, _062038_, _062039_, _062040_, _062041_, _062042_, _062043_, _062044_, _062045_, _062046_, _062047_, _062048_, _062049_, _062050_, _062051_, _062052_, _062053_, _062054_, _062055_, _062056_, _062057_, _062058_, _062059_, _062060_, _062061_, _062062_, _062063_, _062064_, _062065_, _062066_, _062067_, _062068_, _062069_, _062070_, _062071_, _062072_, _062073_, _062074_, _062075_, _062076_, _062077_, _062078_, _062079_, _062080_, _062081_, _062082_, _062083_, _062084_, _062085_, _062086_, _062087_, _062088_, _062089_, _062090_, _062091_, _062092_, _062093_, _062094_, _062095_, _062096_, _062097_, _062098_, _062099_, _062100_, _062101_, _062102_, _062103_, _062104_, _062105_, _062106_, _062107_, _062108_, _062109_, _062110_, _062111_, _062112_, _062113_, _062114_, _062115_, _062116_, _062117_, _062118_, _062119_, _062120_, _062121_, _062122_, _062123_, _062124_, _062125_, _062126_, _062127_, _062128_, _062129_, _062130_, _062131_, _062132_, _062133_, _062134_, _062135_, _062136_, _062137_, _062138_, _062139_, _062140_, _062141_, _062142_, _062143_, _062144_, _062145_, _062146_, _062147_, _062148_, _062149_, _062150_, _062151_, _062152_, _062153_, _062154_, _062155_, _062156_, _062157_, _062158_, _062159_, _062160_, _062161_, _062162_, _062163_, _062164_, _062165_, _062166_, _062167_, _062168_, _062169_, _062170_, _062171_, _062172_, _062173_, _062174_, _062175_, _062176_, _062177_, _062178_, _062179_, _062180_, _062181_, _062182_, _062183_, _062184_, _062185_, _062186_, _062187_, _062188_, _062189_, _062190_, _062191_, _062192_, _062193_, _062194_, _062195_, _062196_, _062197_, _062198_, _062199_, _062200_, _062201_, _062202_, _062203_, _062204_, _062205_, _062206_, _062207_, _062208_, _062209_, _062210_, _062211_, _062212_, _062213_, _062214_, _062215_, _062216_, _062217_, _062218_, _062219_, _062220_, _062221_, _062222_, _062223_, _062224_, _062225_, _062226_, _062227_, _062228_, _062229_, _062230_, _062231_, _062232_, _062233_, _062234_, _062235_, _062236_, _062237_, _062238_, _062239_, _062240_, _062241_, _062242_, _062243_, _062244_, _062245_, _062246_, _062247_, _062248_, _062249_, _062250_, _062251_, _062252_, _062253_, _062254_, _062255_, _062256_, _062257_, _062258_, _062259_, _062260_, _062261_, _062262_, _062263_, _062264_, _062265_, _062266_, _062267_, _062268_, _062269_, _062270_, _062271_, _062272_, _062273_, _062274_, _062275_, _062276_, _062277_, _062278_, _062279_, _062280_, _062281_, _062282_, _062283_, _062284_, _062285_, _062286_, _062287_, _062288_, _062289_, _062290_, _062291_, _062292_, _062293_, _062294_, _062295_, _062296_, _062297_, _062298_, _062299_, _062300_, _062301_, _062302_, _062303_, _062304_, _062305_, _062306_, _062307_, _062308_, _062309_, _062310_, _062311_, _062312_, _062313_, _062314_, _062315_, _062316_, _062317_, _062318_, _062319_, _062320_, _062321_, _062322_, _062323_, _062324_, _062325_, _062326_, _062327_, _062328_, _062329_, _062330_, _062331_, _062332_, _062333_, _062334_, _062335_, _062336_, _062337_, _062338_, _062339_, _062340_, _062341_, _062342_, _062343_, _062344_, _062345_, _062346_, _062347_, _062348_, _062349_, _062350_, _062351_, _062352_, _062353_, _062354_, _062355_, _062356_, _062357_, _062358_, _062359_, _062360_, _062361_, _062362_, _062363_, _062364_, _062365_, _062366_, _062367_, _062368_, _062369_, _062370_, _062371_, _062372_, _062373_, _062374_, _062375_, _062376_, _062377_, _062378_, _062379_, _062380_, _062381_, _062382_, _062383_, _062384_, _062385_, _062386_, _062387_, _062388_, _062389_, _062390_, _062391_, _062392_, _062393_, _062394_, _062395_, _062396_, _062397_, _062398_, _062399_, _062400_, _062401_, _062402_, _062403_, _062404_, _062405_, _062406_, _062407_, _062408_, _062409_, _062410_, _062411_, _062412_, _062413_, _062414_, _062415_, _062416_, _062417_, _062418_, _062419_, _062420_, _062421_, _062422_, _062423_, _062424_, _062425_, _062426_, _062427_, _062428_, _062429_, _062430_, _062431_, _062432_, _062433_, _062434_, _062435_, _062436_, _062437_, _062438_, _062439_, _062440_, _062441_, _062442_, _062443_, _062444_, _062445_, _062446_, _062447_, _062448_, _062449_, _062450_, _062451_, _062452_, _062453_, _062454_, _062455_, _062456_, _062457_, _062458_, _062459_, _062460_, _062461_, _062462_, _062463_, _062464_, _062465_, _062466_, _062467_, _062468_, _062469_, _062470_, _062471_, _062472_, _062473_, _062474_, _062475_, _062476_, _062477_, _062478_, _062479_, _062480_, _062481_, _062482_, _062483_, _062484_, _062485_, _062486_, _062487_, _062488_, _062489_, _062490_, _062491_, _062492_, _062493_, _062494_, _062495_, _062496_, _062497_, _062498_, _062499_, _062500_, _062501_, _062502_, _062503_, _062504_, _062505_, _062506_, _062507_, _062508_, _062509_, _062510_, _062511_, _062512_, _062513_, _062514_, _062515_, _062516_, _062517_, _062518_, _062519_, _062520_, _062521_, _062522_, _062523_, _062524_, _062525_, _062526_, _062527_, _062528_, _062529_, _062530_, _062531_, _062532_, _062533_, _062534_, _062535_, _062536_, _062537_, _062538_, _062539_, _062540_, _062541_, _062542_, _062543_, _062544_, _062545_, _062546_, _062547_, _062548_, _062549_, _062550_, _062551_, _062552_, _062553_, _062554_, _062555_, _062556_, _062557_, _062558_, _062559_, _062560_, _062561_, _062562_, _062563_, _062564_, _062565_, _062566_, _062567_, _062568_, _062569_, _062570_, _062571_, _062572_, _062573_, _062574_, _062575_, _062576_, _062577_, _062578_, _062579_, _062580_, _062581_, _062582_, _062583_, _062584_, _062585_, _062586_, _062587_, _062588_, _062589_, _062590_, _062591_, _062592_, _062593_, _062594_, _062595_, _062596_, _062597_, _062598_, _062599_, _062600_, _062601_, _062602_, _062603_, _062604_, _062605_, _062606_, _062607_, _062608_, _062609_, _062610_, _062611_, _062612_, _062613_, _062614_, _062615_, _062616_, _062617_, _062618_, _062619_, _062620_, _062621_, _062622_, _062623_, _062624_, _062625_, _062626_, _062627_, _062628_, _062629_, _062630_, _062631_, _062632_, _062633_, _062634_, _062635_, _062636_, _062637_, _062638_, _062639_, _062640_, _062641_, _062642_, _062643_, _062644_, _062645_, _062646_, _062647_, _062648_, _062649_, _062650_, _062651_, _062652_, _062653_, _062654_, _062655_, _062656_, _062657_, _062658_, _062659_, _062660_, _062661_, _062662_, _062663_, _062664_, _062665_, _062666_, _062667_, _062668_, _062669_, _062670_, _062671_, _062672_, _062673_, _062674_, _062675_, _062676_, _062677_, _062678_, _062679_, _062680_, _062681_, _062682_, _062683_, _062684_, _062685_, _062686_, _062687_, _062688_, _062689_, _062690_, _062691_, _062692_, _062693_, _062694_, _062695_, _062696_, _062697_, _062698_, _062699_, _062700_, _062701_, _062702_, _062703_, _062704_, _062705_, _062706_, _062707_, _062708_, _062709_, _062710_, _062711_, _062712_, _062713_, _062714_, _062715_, _062716_, _062717_, _062718_, _062719_, _062720_, _062721_, _062722_, _062723_, _062724_, _062725_, _062726_, _062727_, _062728_, _062729_, _062730_, _062731_, _062732_, _062733_, _062734_, _062735_, _062736_, _062737_, _062738_, _062739_, _062740_, _062741_, _062742_, _062743_, _062744_, _062745_, _062746_, _062747_, _062748_, _062749_, _062750_, _062751_, _062752_, _062753_, _062754_, _062755_, _062756_, _062757_, _062758_, _062759_, _062760_, _062761_, _062762_, _062763_, _062764_, _062765_, _062766_, _062767_, _062768_, _062769_, _062770_, _062771_, _062772_, _062773_, _062774_, _062775_, _062776_, _062777_, _062778_, _062779_, _062780_, _062781_, _062782_, _062783_, _062784_, _062785_, _062786_, _062787_, _062788_, _062789_, _062790_, _062791_, _062792_, _062793_, _062794_, _062795_, _062796_, _062797_, _062798_, _062799_, _062800_, _062801_, _062802_, _062803_, _062804_, _062805_, _062806_, _062807_, _062808_, _062809_, _062810_, _062811_, _062812_, _062813_, _062814_, _062815_, _062816_, _062817_, _062818_, _062819_, _062820_, _062821_, _062822_, _062823_, _062824_, _062825_, _062826_, _062827_, _062828_, _062829_, _062830_, _062831_, _062832_, _062833_, _062834_, _062835_, _062836_, _062837_, _062838_, _062839_, _062840_, _062841_, _062842_, _062843_, _062844_, _062845_, _062846_, _062847_, _062848_, _062849_, _062850_, _062851_, _062852_, _062853_, _062854_, _062855_, _062856_, _062857_, _062858_, _062859_, _062860_, _062861_, _062862_, _062863_, _062864_, _062865_, _062866_, _062867_, _062868_, _062869_, _062870_, _062871_, _062872_, _062873_, _062874_, _062875_, _062876_, _062877_, _062878_, _062879_, _062880_, _062881_, _062882_, _062883_, _062884_, _062885_, _062886_, _062887_, _062888_, _062889_, _062890_, _062891_, _062892_, _062893_, _062894_, _062895_, _062896_, _062897_, _062898_, _062899_, _062900_, _062901_, _062902_, _062903_, _062904_, _062905_, _062906_, _062907_, _062908_, _062909_, _062910_, _062911_, _062912_, _062913_, _062914_, _062915_, _062916_, _062917_, _062918_, _062919_, _062920_, _062921_, _062922_, _062923_, _062924_, _062925_, _062926_, _062927_, _062928_, _062929_, _062930_, _062931_, _062932_, _062933_, _062934_, _062935_, _062936_, _062937_, _062938_, _062939_, _062940_, _062941_, _062942_, _062943_, _062944_, _062945_, _062946_, _062947_, _062948_, _062949_, _062950_, _062951_, _062952_, _062953_, _062954_, _062955_, _062956_, _062957_, _062958_, _062959_, _062960_, _062961_, _062962_, _062963_, _062964_, _062965_, _062966_, _062967_, _062968_, _062969_, _062970_, _062971_, _062972_, _062973_, _062974_, _062975_, _062976_, _062977_, _062978_, _062979_, _062980_, _062981_, _062982_, _062983_, _062984_, _062985_, _062986_, _062987_, _062988_, _062989_, _062990_, _062991_, _062992_, _062993_, _062994_, _062995_, _062996_, _062997_, _062998_, _062999_, _063000_, _063001_, _063002_, _063003_, _063004_, _063005_, _063006_, _063007_, _063008_, _063009_, _063010_, _063011_, _063012_, _063013_, _063014_, _063015_, _063016_, _063017_, _063018_, _063019_, _063020_, _063021_, _063022_, _063023_, _063024_, _063025_, _063026_, _063027_, _063028_, _063029_, _063030_, _063031_, _063032_, _063033_, _063034_, _063035_, _063036_, _063037_, _063038_, _063039_, _063040_, _063041_, _063042_, _063043_, _063044_, _063045_, _063046_, _063047_, _063048_, _063049_, _063050_, _063051_, _063052_, _063053_, _063054_, _063055_, _063056_, _063057_, _063058_, _063059_, _063060_, _063061_, _063062_, _063063_, _063064_, _063065_, _063066_, _063067_, _063068_, _063069_, _063070_, _063071_, _063072_, _063073_, _063074_, _063075_, _063076_, _063077_, _063078_, _063079_, _063080_, _063081_, _063082_, _063083_, _063084_, _063085_, _063086_, _063087_, _063088_, _063089_, _063090_, _063091_, _063092_, _063093_, _063094_, _063095_, _063096_, _063097_, _063098_, _063099_, _063100_, _063101_, _063102_, _063103_, _063104_, _063105_, _063106_, _063107_, _063108_, _063109_, _063110_, _063111_, _063112_, _063113_, _063114_, _063115_, _063116_, _063117_, _063118_, _063119_, _063120_, _063121_, _063122_, _063123_, _063124_, _063125_, _063126_, _063127_, _063128_, _063129_, _063130_, _063131_, _063132_, _063133_, _063134_, _063135_, _063136_, _063137_, _063138_, _063139_, _063140_, _063141_, _063142_, _063143_, _063144_, _063145_, _063146_, _063147_, _063148_, _063149_, _063150_, _063151_, _063152_, _063153_, _063154_, _063155_, _063156_, _063157_, _063158_, _063159_, _063160_, _063161_, _063162_, _063163_, _063164_, _063165_, _063166_, _063167_, _063168_, _063169_, _063170_, _063171_, _063172_, _063173_, _063174_, _063175_, _063176_, _063177_, _063178_, _063179_, _063180_, _063181_, _063182_, _063183_, _063184_, _063185_, _063186_, _063187_, _063188_, _063189_, _063190_, _063191_, _063192_, _063193_, _063194_, _063195_, _063196_, _063197_, _063198_, _063199_, _063200_, _063201_, _063202_, _063203_, _063204_, _063205_, _063206_, _063207_, _063208_, _063209_, _063210_, _063211_, _063212_, _063213_, _063214_, _063215_, _063216_, _063217_, _063218_, _063219_, _063220_, _063221_, _063222_, _063223_, _063224_, _063225_, _063226_, _063227_, _063228_, _063229_, _063230_, _063231_, _063232_, _063233_, _063234_, _063235_, _063236_, _063237_, _063238_, _063239_, _063240_, _063241_, _063242_, _063243_, _063244_, _063245_, _063246_, _063247_, _063248_, _063249_, _063250_, _063251_, _063252_, _063253_, _063254_, _063255_, _063256_, _063257_, _063258_, _063259_, _063260_, _063261_, _063262_, _063263_, _063264_, _063265_, _063266_, _063267_, _063268_, _063269_, _063270_, _063271_, _063272_, _063273_, _063274_, _063275_, _063276_, _063277_, _063278_, _063279_, _063280_, _063281_, _063282_, _063283_, _063284_, _063285_, _063286_, _063287_, _063288_, _063289_, _063290_, _063291_, _063292_, _063293_, _063294_, _063295_, _063296_, _063297_, _063298_, _063299_, _063300_, _063301_, _063302_, _063303_, _063304_, _063305_, _063306_, _063307_, _063308_, _063309_, _063310_, _063311_, _063312_, _063313_, _063314_, _063315_, _063316_, _063317_, _063318_, _063319_, _063320_, _063321_, _063322_, _063323_, _063324_, _063325_, _063326_, _063327_, _063328_, _063329_, _063330_, _063331_, _063332_, _063333_, _063334_, _063335_, _063336_, _063337_, _063338_, _063339_, _063340_, _063341_, _063342_, _063343_, _063344_, _063345_, _063346_, _063347_, _063348_, _063349_, _063350_, _063351_, _063352_, _063353_, _063354_, _063355_, _063356_, _063357_, _063358_, _063359_, _063360_, _063361_, _063362_, _063363_, _063364_, _063365_, _063366_, _063367_, _063368_, _063369_, _063370_, _063371_, _063372_, _063373_, _063374_, _063375_, _063376_, _063377_, _063378_, _063379_, _063380_, _063381_, _063382_, _063383_, _063384_, _063385_, _063386_, _063387_, _063388_, _063389_, _063390_, _063391_, _063392_, _063393_, _063394_, _063395_, _063396_, _063397_, _063398_, _063399_, _063400_, _063401_, _063402_, _063403_, _063404_, _063405_, _063406_, _063407_, _063408_, _063409_, _063410_, _063411_, _063412_, _063413_, _063414_, _063415_, _063416_, _063417_, _063418_, _063419_, _063420_, _063421_, _063422_, _063423_, _063424_, _063425_, _063426_, _063427_, _063428_, _063429_, _063430_, _063431_, _063432_, _063433_, _063434_, _063435_, _063436_, _063437_, _063438_, _063439_, _063440_, _063441_, _063442_, _063443_, _063444_, _063445_, _063446_, _063447_, _063448_, _063449_, _063450_, _063451_, _063452_, _063453_, _063454_, _063455_, _063456_, _063457_, _063458_, _063459_, _063460_, _063461_, _063462_, _063463_, _063464_, _063465_, _063466_, _063467_, _063468_, _063469_, _063470_, _063471_, _063472_, _063473_, _063474_, _063475_, _063476_, _063477_, _063478_, _063479_, _063480_, _063481_, _063482_, _063483_, _063484_, _063485_, _063486_, _063487_, _063488_, _063489_, _063490_, _063491_, _063492_, _063493_, _063494_, _063495_, _063496_, _063497_, _063498_, _063499_, _063500_, _063501_, _063502_, _063503_, _063504_, _063505_, _063506_, _063507_, _063508_, _063509_, _063510_, _063511_, _063512_, _063513_, _063514_, _063515_, _063516_, _063517_, _063518_, _063519_, _063520_, _063521_, _063522_, _063523_, _063524_, _063525_, _063526_, _063527_, _063528_, _063529_, _063530_, _063531_, _063532_, _063533_, _063534_, _063535_, _063536_, _063537_, _063538_, _063539_, _063540_, _063541_, _063542_, _063543_, _063544_, _063545_, _063546_, _063547_, _063548_, _063549_, _063550_, _063551_, _063552_, _063553_, _063554_, _063555_, _063556_, _063557_, _063558_, _063559_, _063560_, _063561_, _063562_, _063563_, _063564_, _063565_, _063566_, _063567_, _063568_, _063569_, _063570_, _063571_, _063572_, _063573_, _063574_, _063575_, _063576_, _063577_, _063578_, _063579_, _063580_, _063581_, _063582_, _063583_, _063584_, _063585_, _063586_, _063587_, _063588_, _063589_, _063590_, _063591_, _063592_, _063593_, _063594_, _063595_, _063596_, _063597_, _063598_, _063599_, _063600_, _063601_, _063602_, _063603_, _063604_, _063605_, _063606_, _063607_, _063608_, _063609_, _063610_, _063611_, _063612_, _063613_, _063614_, _063615_, _063616_, _063617_, _063618_, _063619_, _063620_, _063621_, _063622_, _063623_, _063624_, _063625_, _063626_, _063627_, _063628_, _063629_, _063630_, _063631_, _063632_, _063633_, _063634_, _063635_, _063636_, _063637_, _063638_, _063639_, _063640_, _063641_, _063642_, _063643_, _063644_, _063645_, _063646_, _063647_, _063648_, _063649_, _063650_, _063651_, _063652_, _063653_, _063654_, _063655_, _063656_, _063657_, _063658_, _063659_, _063660_, _063661_, _063662_, _063663_, _063664_, _063665_, _063666_, _063667_, _063668_, _063669_, _063670_, _063671_, _063672_, _063673_, _063674_, _063675_, _063676_, _063677_, _063678_, _063679_, _063680_, _063681_, _063682_, _063683_, _063684_, _063685_, _063686_, _063687_, _063688_, _063689_, _063690_, _063691_, _063692_, _063693_, _063694_, _063695_, _063696_, _063697_, _063698_, _063699_, _063700_, _063701_, _063702_, _063703_, _063704_, _063705_, _063706_, _063707_, _063708_, _063709_, _063710_, _063711_, _063712_, _063713_, _063714_, _063715_, _063716_, _063717_, _063718_, _063719_, _063720_, _063721_, _063722_, _063723_, _063724_, _063725_, _063726_, _063727_, _063728_, _063729_, _063730_, _063731_, _063732_, _063733_, _063734_, _063735_, _063736_, _063737_, _063738_, _063739_, _063740_, _063741_, _063742_, _063743_, _063744_, _063745_, _063746_, _063747_, _063748_, _063749_, _063750_, _063751_, _063752_, _063753_, _063754_, _063755_, _063756_, _063757_, _063758_, _063759_, _063760_, _063761_, _063762_, _063763_, _063764_, _063765_, _063766_, _063767_, _063768_, _063769_, _063770_, _063771_, _063772_, _063773_, _063774_, _063775_, _063776_, _063777_, _063778_, _063779_, _063780_, _063781_, _063782_, _063783_, _063784_, _063785_, _063786_, _063787_, _063788_, _063789_, _063790_, _063791_, _063792_, _063793_, _063794_, _063795_, _063796_, _063797_, _063798_, _063799_, _063800_, _063801_, _063802_, _063803_, _063804_, _063805_, _063806_, _063807_, _063808_, _063809_, _063810_, _063811_, _063812_, _063813_, _063814_, _063815_, _063816_, _063817_, _063818_, _063819_, _063820_, _063821_, _063822_, _063823_, _063824_, _063825_, _063826_, _063827_, _063828_, _063829_, _063830_, _063831_, _063832_, _063833_, _063834_, _063835_, _063836_, _063837_, _063838_, _063839_, _063840_, _063841_, _063842_, _063843_, _063844_, _063845_, _063846_, _063847_, _063848_, _063849_, _063850_, _063851_, _063852_, _063853_, _063854_, _063855_, _063856_, _063857_, _063858_, _063859_, _063860_, _063861_, _063862_, _063863_, _063864_, _063865_, _063866_, _063867_, _063868_, _063869_, _063870_, _063871_, _063872_, _063873_, _063874_, _063875_, _063876_, _063877_, _063878_, _063879_, _063880_, _063881_, _063882_, _063883_, _063884_, _063885_, _063886_, _063887_, _063888_, _063889_, _063890_, _063891_, _063892_, _063893_, _063894_, _063895_, _063896_, _063897_, _063898_, _063899_, _063900_, _063901_, _063902_, _063903_, _063904_, _063905_, _063906_, _063907_, _063908_, _063909_, _063910_, _063911_, _063912_, _063913_, _063914_, _063915_, _063916_, _063917_, _063918_, _063919_, _063920_, _063921_, _063922_, _063923_, _063924_, _063925_, _063926_, _063927_, _063928_, _063929_, _063930_, _063931_, _063932_, _063933_, _063934_, _063935_, _063936_, _063937_, _063938_, _063939_, _063940_, _063941_, _063942_, _063943_, _063944_, _063945_, _063946_, _063947_, _063948_, _063949_, _063950_, _063951_, _063952_, _063953_, _063954_, _063955_, _063956_, _063957_, _063958_, _063959_, _063960_, _063961_, _063962_, _063963_, _063964_, _063965_, _063966_, _063967_, _063968_, _063969_, _063970_, _063971_, _063972_, _063973_, _063974_, _063975_, _063976_, _063977_, _063978_, _063979_, _063980_, _063981_, _063982_, _063983_, _063984_, _063985_, _063986_, _063987_, _063988_, _063989_, _063990_, _063991_, _063992_, _063993_, _063994_, _063995_, _063996_, _063997_, _063998_, _063999_, _064000_, _064001_, _064002_, _064003_, _064004_, _064005_, _064006_, _064007_, _064008_, _064009_, _064010_, _064011_, _064012_, _064013_, _064014_, _064015_, _064016_, _064017_, _064018_, _064019_, _064020_, _064021_, _064022_, _064023_, _064024_, _064025_, _064026_, _064027_, _064028_, _064029_, _064030_, _064031_, _064032_, _064033_, _064034_, _064035_, _064036_, _064037_, _064038_, _064039_, _064040_, _064041_, _064042_, _064043_, _064044_, _064045_, _064046_, _064047_, _064048_, _064049_, _064050_, _064051_, _064052_, _064053_, _064054_, _064055_, _064056_, _064057_, _064058_, _064059_, _064060_, _064061_, _064062_, _064063_, _064064_, _064065_, _064066_, _064067_, _064068_, _064069_, _064070_, _064071_, _064072_, _064073_, _064074_, _064075_, _064076_, _064077_, _064078_, _064079_, _064080_, _064081_, _064082_, _064083_, _064084_, _064085_, _064086_, _064087_, _064088_, _064089_, _064090_, _064091_, _064092_, _064093_, _064094_, _064095_, _064096_, _064097_, _064098_, _064099_, _064100_, _064101_, _064102_, _064103_, _064104_, _064105_, _064106_, _064107_, _064108_, _064109_, _064110_, _064111_, _064112_, _064113_, _064114_, _064115_, _064116_, _064117_, _064118_, _064119_, _064120_, _064121_, _064122_, _064123_, _064124_, _064125_, _064126_, _064127_, _064128_, _064129_, _064130_, _064131_, _064132_, _064133_, _064134_, _064135_, _064136_, _064137_, _064138_, _064139_, _064140_, _064141_, _064142_, _064143_, _064144_, _064145_, _064146_, _064147_, _064148_, _064149_, _064150_, _064151_, _064152_, _064153_, _064154_, _064155_, _064156_, _064157_, _064158_, _064159_, _064160_, _064161_, _064162_, _064163_, _064164_, _064165_, _064166_, _064167_, _064168_, _064169_, _064170_, _064171_, _064172_, _064173_, _064174_, _064175_, _064176_, _064177_, _064178_, _064179_, _064180_, _064181_, _064182_, _064183_, _064184_, _064185_, _064186_, _064187_, _064188_, _064189_, _064190_, _064191_, _064192_, _064193_, _064194_, _064195_, _064196_, _064197_, _064198_, _064199_, _064200_, _064201_, _064202_, _064203_, _064204_, _064205_, _064206_, _064207_, _064208_, _064209_, _064210_, _064211_, _064212_, _064213_, _064214_, _064215_, _064216_, _064217_, _064218_, _064219_, _064220_, _064221_, _064222_, _064223_, _064224_, _064225_, _064226_, _064227_, _064228_, _064229_, _064230_, _064231_, _064232_, _064233_, _064234_, _064235_, _064236_, _064237_, _064238_, _064239_, _064240_, _064241_, _064242_, _064243_, _064244_, _064245_, _064246_, _064247_, _064248_, _064249_, _064250_, _064251_, _064252_, _064253_, _064254_, _064255_, _064256_, _064257_, _064258_, _064259_, _064260_, _064261_, _064262_, _064263_, _064264_, _064265_, _064266_, _064267_, _064268_, _064269_, _064270_, _064271_, _064272_, _064273_, _064274_, _064275_, _064276_, _064277_, _064278_, _064279_, _064280_, _064281_, _064282_, _064283_, _064284_, _064285_, _064286_, _064287_, _064288_, _064289_, _064290_, _064291_, _064292_, _064293_, _064294_, _064295_, _064296_, _064297_, _064298_, _064299_, _064300_, _064301_, _064302_, _064303_, _064304_, _064305_, _064306_, _064307_, _064308_, _064309_, _064310_, _064311_, _064312_, _064313_, _064314_, _064315_, _064316_, _064317_, _064318_, _064319_, _064320_, _064321_, _064322_, _064323_, _064324_, _064325_, _064326_, _064327_, _064328_, _064329_, _064330_, _064331_, _064332_, _064333_, _064334_, _064335_, _064336_, _064337_, _064338_, _064339_, _064340_, _064341_, _064342_, _064343_, _064344_, _064345_, _064346_, _064347_, _064348_, _064349_, _064350_, _064351_, _064352_, _064353_, _064354_, _064355_, _064356_, _064357_, _064358_, _064359_, _064360_, _064361_, _064362_, _064363_, _064364_, _064365_, _064366_, _064367_, _064368_, _064369_, _064370_, _064371_, _064372_, _064373_, _064374_, _064375_, _064376_, _064377_, _064378_, _064379_, _064380_, _064381_, _064382_, _064383_, _064384_, _064385_, _064386_, _064387_, _064388_, _064389_, _064390_, _064391_, _064392_, _064393_, _064394_, _064395_, _064396_, _064397_, _064398_, _064399_, _064400_, _064401_, _064402_, _064403_, _064404_, _064405_, _064406_, _064407_, _064408_, _064409_, _064410_, _064411_, _064412_, _064413_, _064414_, _064415_, _064416_, _064417_, _064418_, _064419_, _064420_, _064421_, _064422_, _064423_, _064424_, _064425_, _064426_, _064427_, _064428_, _064429_, _064430_, _064431_, _064432_, _064433_, _064434_, _064435_, _064436_, _064437_, _064438_, _064439_, _064440_, _064441_, _064442_, _064443_, _064444_, _064445_, _064446_, _064447_, _064448_, _064449_, _064450_, _064451_, _064452_, _064453_, _064454_, _064455_, _064456_, _064457_, _064458_, _064459_, _064460_, _064461_, _064462_, _064463_, _064464_, _064465_, _064466_, _064467_, _064468_, _064469_, _064470_, _064471_, _064472_, _064473_, _064474_, _064475_, _064476_, _064477_, _064478_, _064479_, _064480_, _064481_, _064482_, _064483_, _064484_, _064485_, _064486_, _064487_, _064488_, _064489_, _064490_, _064491_, _064492_, _064493_, _064494_, _064495_, _064496_, _064497_, _064498_, _064499_, _064500_, _064501_, _064502_, _064503_, _064504_, _064505_, _064506_, _064507_, _064508_, _064509_, _064510_, _064511_, _064512_, _064513_, _064514_, _064515_, _064516_, _064517_, _064518_, _064519_, _064520_, _064521_, _064522_, _064523_, _064524_, _064525_, _064526_, _064527_, _064528_, _064529_, _064530_, _064531_, _064532_, _064533_, _064534_, _064535_, _064536_, _064537_, _064538_, _064539_, _064540_, _064541_, _064542_, _064543_, _064544_, _064545_, _064546_, _064547_, _064548_, _064549_, _064550_, _064551_, _064552_, _064553_, _064554_, _064555_, _064556_, _064557_, _064558_, _064559_, _064560_, _064561_, _064562_, _064563_, _064564_, _064565_, _064566_, _064567_, _064568_, _064569_, _064570_, _064571_, _064572_, _064573_, _064574_, _064575_, _064576_, _064577_, _064578_, _064579_, _064580_, _064581_, _064582_, _064583_, _064584_, _064585_, _064586_, _064587_, _064588_, _064589_, _064590_, _064591_, _064592_, _064593_, _064594_, _064595_, _064596_, _064597_, _064598_, _064599_, _064600_, _064601_, _064602_, _064603_, _064604_, _064605_, _064606_, _064607_, _064608_, _064609_, _064610_, _064611_, _064612_, _064613_, _064614_, _064615_, _064616_, _064617_, _064618_, _064619_, _064620_, _064621_, _064622_, _064623_, _064624_, _064625_, _064626_, _064627_, _064628_, _064629_, _064630_, _064631_, _064632_, _064633_, _064634_, _064635_, _064636_, _064637_, _064638_, _064639_, _064640_, _064641_, _064642_, _064643_, _064644_, _064645_, _064646_, _064647_, _064648_, _064649_, _064650_, _064651_, _064652_, _064653_, _064654_, _064655_, _064656_, _064657_, _064658_, _064659_, _064660_, _064661_, _064662_, _064663_, _064664_, _064665_, _064666_, _064667_, _064668_, _064669_, _064670_, _064671_, _064672_, _064673_, _064674_, _064675_, _064676_, _064677_, _064678_, _064679_, _064680_, _064681_, _064682_, _064683_, _064684_, _064685_, _064686_, _064687_, _064688_, _064689_, _064690_, _064691_, _064692_, _064693_, _064694_, _064695_, _064696_, _064697_, _064698_, _064699_, _064700_, _064701_, _064702_, _064703_, _064704_, _064705_, _064706_, _064707_, _064708_, _064709_, _064710_, _064711_, _064712_, _064713_, _064714_, _064715_, _064716_, _064717_, _064718_, _064719_, _064720_, _064721_, _064722_, _064723_, _064724_, _064725_, _064726_, _064727_, _064728_, _064729_, _064730_, _064731_, _064732_, _064733_, _064734_, _064735_, _064736_, _064737_, _064738_, _064739_, _064740_, _064741_, _064742_, _064743_, _064744_, _064745_, _064746_, _064747_, _064748_, _064749_, _064750_, _064751_, _064752_, _064753_, _064754_, _064755_, _064756_, _064757_, _064758_, _064759_, _064760_, _064761_, _064762_, _064763_, _064764_, _064765_, _064766_, _064767_, _064768_, _064769_, _064770_, _064771_, _064772_, _064773_, _064774_, _064775_, _064776_, _064777_, _064778_, _064779_, _064780_, _064781_, _064782_, _064783_, _064784_, _064785_, _064786_, _064787_, _064788_, _064789_, _064790_, _064791_, _064792_, _064793_, _064794_, _064795_, _064796_, _064797_, _064798_, _064799_, _064800_, _064801_, _064802_, _064803_, _064804_, _064805_, _064806_, _064807_, _064808_, _064809_, _064810_, _064811_, _064812_, _064813_, _064814_, _064815_, _064816_, _064817_, _064818_, _064819_, _064820_, _064821_, _064822_, _064823_, _064824_, _064825_, _064826_, _064827_, _064828_, _064829_, _064830_, _064831_, _064832_, _064833_, _064834_, _064835_, _064836_, _064837_, _064838_, _064839_, _064840_, _064841_, _064842_, _064843_, _064844_, _064845_, _064846_, _064847_, _064848_, _064849_, _064850_, _064851_, _064852_, _064853_, _064854_, _064855_, _064856_, _064857_, _064858_, _064859_, _064860_, _064861_, _064862_, _064863_, _064864_, _064865_, _064866_, _064867_, _064868_, _064869_, _064870_, _064871_, _064872_, _064873_, _064874_, _064875_, _064876_, _064877_, _064878_, _064879_, _064880_, _064881_, _064882_, _064883_, _064884_, _064885_, _064886_, _064887_, _064888_, _064889_, _064890_, _064891_, _064892_, _064893_, _064894_, _064895_, _064896_, _064897_, _064898_, _064899_, _064900_, _064901_, _064902_, _064903_, _064904_, _064905_, _064906_, _064907_, _064908_, _064909_, _064910_, _064911_, _064912_, _064913_, _064914_, _064915_, _064916_, _064917_, _064918_, _064919_, _064920_, _064921_, _064922_, _064923_, _064924_, _064925_, _064926_, _064927_, _064928_, _064929_, _064930_, _064931_, _064932_, _064933_, _064934_, _064935_, _064936_, _064937_, _064938_, _064939_, _064940_, _064941_, _064942_, _064943_, _064944_, _064945_, _064946_, _064947_, _064948_, _064949_, _064950_, _064951_, _064952_, _064953_, _064954_, _064955_, _064956_, _064957_, _064958_, _064959_, _064960_, _064961_, _064962_, _064963_, _064964_, _064965_, _064966_, _064967_, _064968_, _064969_, _064970_, _064971_, _064972_, _064973_, _064974_, _064975_, _064976_, _064977_, _064978_, _064979_, _064980_, _064981_, _064982_, _064983_, _064984_, _064985_, _064986_, _064987_, _064988_, _064989_, _064990_, _064991_, _064992_, _064993_, _064994_, _064995_, _064996_, _064997_, _064998_, _064999_, _065000_, _065001_, _065002_, _065003_, _065004_, _065005_, _065006_, _065007_, _065008_, _065009_, _065010_, _065011_, _065012_, _065013_, _065014_, _065015_, _065016_, _065017_, _065018_, _065019_, _065020_, _065021_, _065022_, _065023_, _065024_, _065025_, _065026_, _065027_, _065028_, _065029_, _065030_, _065031_, _065032_, _065033_, _065034_, _065035_, _065036_, _065037_, _065038_, _065039_, _065040_, _065041_, _065042_, _065043_, _065044_, _065045_, _065046_, _065047_, _065048_, _065049_, _065050_, _065051_, _065052_, _065053_, _065054_, _065055_, _065056_, _065057_, _065058_, _065059_, _065060_, _065061_, _065062_, _065063_, _065064_, _065065_, _065066_, _065067_, _065068_, _065069_, _065070_, _065071_, _065072_, _065073_, _065074_, _065075_, _065076_, _065077_, _065078_, _065079_, _065080_, _065081_, _065082_, _065083_, _065084_, _065085_, _065086_, _065087_, _065088_, _065089_, _065090_, _065091_, _065092_, _065093_, _065094_, _065095_, _065096_, _065097_, _065098_, _065099_, _065100_, _065101_, _065102_, _065103_, _065104_, _065105_, _065106_, _065107_, _065108_, _065109_, _065110_, _065111_, _065112_, _065113_, _065114_, _065115_, _065116_, _065117_, _065118_, _065119_, _065120_, _065121_, _065122_, _065123_, _065124_, _065125_, _065126_, _065127_, _065128_, _065129_, _065130_, _065131_, _065132_, _065133_, _065134_, _065135_, _065136_, _065137_, _065138_, _065139_, _065140_, _065141_, _065142_, _065143_, _065144_, _065145_, _065146_, _065147_, _065148_, _065149_, _065150_, _065151_, _065152_, _065153_, _065154_, _065155_, _065156_, _065157_, _065158_, _065159_, _065160_, _065161_, _065162_, _065163_, _065164_, _065165_, _065166_, _065167_, _065168_, _065169_, _065170_, _065171_, _065172_, _065173_, _065174_, _065175_, _065176_, _065177_, _065178_, _065179_, _065180_, _065181_, _065182_, _065183_, _065184_, _065185_, _065186_, _065187_, _065188_, _065189_, _065190_, _065191_, _065192_, _065193_, _065194_, _065195_, _065196_, _065197_, _065198_, _065199_, _065200_, _065201_, _065202_, _065203_, _065204_, _065205_, _065206_, _065207_, _065208_, _065209_, _065210_, _065211_, _065212_, _065213_, _065214_, _065215_, _065216_, _065217_, _065218_, _065219_, _065220_, _065221_, _065222_, _065223_, _065224_, _065225_, _065226_, _065227_, _065228_, _065229_, _065230_, _065231_, _065232_, _065233_, _065234_, _065235_, _065236_, _065237_, _065238_, _065239_, _065240_, _065241_, _065242_, _065243_, _065244_, _065245_, _065246_, _065247_, _065248_, _065249_, _065250_, _065251_, _065252_, _065253_, _065254_, _065255_, _065256_, _065257_, _065258_, _065259_, _065260_, _065261_, _065262_, _065263_, _065264_, _065265_, _065266_, _065267_, _065268_, _065269_, _065270_, _065271_, _065272_, _065273_, _065274_, _065275_, _065276_, _065277_, _065278_, _065279_, _065280_, _065281_, _065282_, _065283_, _065284_, _065285_, _065286_, _065287_, _065288_, _065289_, _065290_, _065291_, _065292_, _065293_, _065294_, _065295_, _065296_, _065297_, _065298_, _065299_, _065300_, _065301_, _065302_, _065303_, _065304_, _065305_, _065306_, _065307_, _065308_, _065309_, _065310_, _065311_, _065312_, _065313_, _065314_, _065315_, _065316_, _065317_, _065318_, _065319_, _065320_, _065321_, _065322_, _065323_, _065324_, _065325_, _065326_, _065327_, _065328_, _065329_, _065330_, _065331_, _065332_, _065333_, _065334_, _065335_, _065336_, _065337_, _065338_, _065339_, _065340_, _065341_, _065342_, _065343_, _065344_, _065345_, _065346_, _065347_, _065348_, _065349_, _065350_, _065351_, _065352_, _065353_, _065354_, _065355_, _065356_, _065357_, _065358_, _065359_, _065360_, _065361_, _065362_, _065363_, _065364_, _065365_, _065366_, _065367_, _065368_, _065369_, _065370_, _065371_, _065372_, _065373_, _065374_, _065375_, _065376_, _065377_, _065378_, _065379_, _065380_, _065381_, _065382_, _065383_, _065384_, _065385_, _065386_, _065387_, _065388_, _065389_, _065390_, _065391_, _065392_, _065393_, _065394_, _065395_, _065396_, _065397_, _065398_, _065399_, _065400_, _065401_, _065402_, _065403_, _065404_, _065405_, _065406_, _065407_, _065408_, _065409_, _065410_, _065411_, _065412_, _065413_, _065414_, _065415_, _065416_, _065417_, _065418_, _065419_, _065420_, _065421_, _065422_, _065423_, _065424_, _065425_, _065426_, _065427_, _065428_, _065429_, _065430_, _065431_, _065432_, _065433_, _065434_, _065435_, _065436_, _065437_, _065438_, _065439_, _065440_, _065441_, _065442_, _065443_, _065444_, _065445_, _065446_, _065447_, _065448_, _065449_, _065450_, _065451_, _065452_, _065453_, _065454_, _065455_, _065456_, _065457_, _065458_, _065459_, _065460_, _065461_, _065462_, _065463_, _065464_, _065465_, _065466_, _065467_, _065468_, _065469_, _065470_, _065471_, _065472_, _065473_, _065474_, _065475_, _065476_, _065477_, _065478_, _065479_, _065480_, _065481_, _065482_, _065483_, _065484_, _065485_, _065486_, _065487_, _065488_, _065489_, _065490_, _065491_, _065492_, _065493_, _065494_, _065495_, _065496_, _065497_, _065498_, _065499_, _065500_, _065501_, _065502_, _065503_, _065504_, _065505_, _065506_, _065507_, _065508_, _065509_, _065510_, _065511_, _065512_, _065513_, _065514_, _065515_, _065516_, _065517_, _065518_, _065519_, _065520_, _065521_, _065522_, _065523_, _065524_, _065525_, _065526_, _065527_, _065528_, _065529_, _065530_, _065531_, _065532_, _065533_, _065534_, _065535_, _065536_, _065537_, _065538_, _065539_, _065540_, _065541_, _065542_, _065543_, _065544_, _065545_, _065546_, _065547_, _065548_, _065549_, _065550_, _065551_, _065552_, _065553_, _065554_, _065555_, _065556_, _065557_, _065558_, _065559_, _065560_, _065561_, _065562_, _065563_, _065564_, _065565_, _065566_, _065567_, _065568_, _065569_, _065570_, _065571_, _065572_, _065573_, _065574_, _065575_, _065576_, _065577_, _065578_, _065579_, _065580_, _065581_, _065582_, _065583_, _065584_, _065585_, _065586_, _065587_, _065588_, _065589_, _065590_, _065591_, _065592_, _065593_, _065594_, _065595_, _065596_, _065597_, _065598_, _065599_, _065600_, _065601_, _065602_, _065603_, _065604_, _065605_, _065606_, _065607_, _065608_, _065609_, _065610_, _065611_, _065612_, _065613_, _065614_, _065615_, _065616_, _065617_, _065618_, _065619_, _065620_, _065621_, _065622_, _065623_, _065624_, _065625_, _065626_, _065627_, _065628_, _065629_, _065630_, _065631_, _065632_, _065633_, _065634_, _065635_, _065636_, _065637_, _065638_, _065639_, _065640_, _065641_, _065642_, _065643_, _065644_, _065645_, _065646_, _065647_, _065648_, _065649_, _065650_, _065651_, _065652_, _065653_, _065654_, _065655_, _065656_, _065657_, _065658_, _065659_, _065660_, _065661_, _065662_, _065663_, _065664_, _065665_, _065666_, _065667_, _065668_, _065669_, _065670_, _065671_, _065672_, _065673_, _065674_, _065675_, _065676_, _065677_, _065678_, _065679_, _065680_, _065681_, _065682_, _065683_, _065684_, _065685_, _065686_, _065687_, _065688_, _065689_, _065690_, _065691_, _065692_, _065693_, _065694_, _065695_, _065696_, _065697_, _065698_, _065699_, _065700_, _065701_, _065702_, _065703_, _065704_, _065705_, _065706_, _065707_, _065708_, _065709_, _065710_, _065711_, _065712_, _065713_, _065714_, _065715_, _065716_, _065717_, _065718_, _065719_, _065720_, _065721_, _065722_, _065723_, _065724_, _065725_, _065726_, _065727_, _065728_, _065729_, _065730_, _065731_, _065732_, _065733_, _065734_, _065735_, _065736_, _065737_, _065738_, _065739_, _065740_, _065741_, _065742_, _065743_, _065744_, _065745_, _065746_, _065747_, _065748_, _065749_, _065750_, _065751_, _065752_, _065753_, _065754_, _065755_, _065756_, _065757_, _065758_, _065759_, _065760_, _065761_, _065762_, _065763_, _065764_, _065765_, _065766_, _065767_, _065768_, _065769_, _065770_, _065771_, _065772_, _065773_, _065774_, _065775_, _065776_, _065777_, _065778_, _065779_, _065780_, _065781_, _065782_, _065783_, _065784_, _065785_, _065786_, _065787_, _065788_, _065789_, _065790_, _065791_, _065792_, _065793_, _065794_, _065795_, _065796_, _065797_, _065798_, _065799_, _065800_, _065801_, _065802_, _065803_, _065804_, _065805_, _065806_, _065807_, _065808_, _065809_, _065810_, _065811_, _065812_, _065813_, _065814_, _065815_, _065816_, _065817_, _065818_, _065819_, _065820_, _065821_, _065822_, _065823_, _065824_, _065825_, _065826_, _065827_, _065828_, _065829_, _065830_, _065831_, _065832_, _065833_, _065834_, _065835_, _065836_, _065837_, _065838_, _065839_, _065840_, _065841_, _065842_, _065843_, _065844_, _065845_, _065846_, _065847_, _065848_, _065849_, _065850_, _065851_, _065852_, _065853_, _065854_, _065855_, _065856_, _065857_, _065858_, _065859_, _065860_, _065861_, _065862_, _065863_, _065864_, _065865_, _065866_, _065867_, _065868_, _065869_, _065870_, _065871_, _065872_, _065873_, _065874_, _065875_, _065876_, _065877_, _065878_, _065879_, _065880_, _065881_, _065882_, _065883_, _065884_, _065885_, _065886_, _065887_, _065888_, _065889_, _065890_, _065891_, _065892_, _065893_, _065894_, _065895_, _065896_, _065897_, _065898_, _065899_, _065900_, _065901_, _065902_, _065903_, _065904_, _065905_, _065906_, _065907_, _065908_, _065909_, _065910_, _065911_, _065912_, _065913_, _065914_, _065915_, _065916_, _065917_, _065918_, _065919_, _065920_, _065921_, _065922_, _065923_, _065924_, _065925_, _065926_, _065927_, _065928_, _065929_, _065930_, _065931_, _065932_, _065933_, _065934_, _065935_, _065936_, _065937_, _065938_, _065939_, _065940_, _065941_, _065942_, _065943_, _065944_, _065945_, _065946_, _065947_, _065948_, _065949_, _065950_, _065951_, _065952_, _065953_, _065954_, _065955_, _065956_, _065957_, _065958_, _065959_, _065960_, _065961_, _065962_, _065963_, _065964_, _065965_, _065966_, _065967_, _065968_, _065969_, _065970_, _065971_, _065972_, _065973_, _065974_, _065975_, _065976_, _065977_, _065978_, _065979_, _065980_, _065981_, _065982_, _065983_, _065984_, _065985_, _065986_, _065987_, _065988_, _065989_, _065990_, _065991_, _065992_, _065993_, _065994_, _065995_, _065996_, _065997_, _065998_, _065999_, _066000_, _066001_, _066002_, _066003_, _066004_, _066005_, _066006_, _066007_, _066008_, _066009_, _066010_, _066011_, _066012_, _066013_, _066014_, _066015_, _066016_, _066017_, _066018_, _066019_, _066020_, _066021_, _066022_, _066023_, _066024_, _066025_, _066026_, _066027_, _066028_, _066029_, _066030_, _066031_, _066032_, _066033_, _066034_, _066035_, _066036_, _066037_, _066038_, _066039_, _066040_, _066041_, _066042_, _066043_, _066044_, _066045_, _066046_, _066047_, _066048_, _066049_, _066050_, _066051_, _066052_, _066053_, _066054_, _066055_, _066056_, _066057_, _066058_, _066059_, _066060_, _066061_, _066062_, _066063_, _066064_, _066065_, _066066_, _066067_, _066068_, _066069_, _066070_, _066071_, _066072_, _066073_, _066074_, _066075_, _066076_, _066077_, _066078_, _066079_, _066080_, _066081_, _066082_, _066083_, _066084_, _066085_, _066086_, _066087_, _066088_, _066089_, _066090_, _066091_, _066092_, _066093_, _066094_, _066095_, _066096_, _066097_, _066098_, _066099_, _066100_, _066101_, _066102_, _066103_, _066104_, _066105_, _066106_, _066107_, _066108_, _066109_, _066110_, _066111_, _066112_, _066113_, _066114_, _066115_, _066116_, _066117_, _066118_, _066119_, _066120_, _066121_, _066122_, _066123_, _066124_, _066125_, _066126_, _066127_, _066128_, _066129_, _066130_, _066131_, _066132_, _066133_, _066134_, _066135_, _066136_, _066137_, _066138_, _066139_, _066140_, _066141_, _066142_, _066143_, _066144_, _066145_, _066146_, _066147_, _066148_, _066149_, _066150_, _066151_, _066152_, _066153_, _066154_, _066155_, _066156_, _066157_, _066158_, _066159_, _066160_, _066161_, _066162_, _066163_, _066164_, _066165_, _066166_, _066167_, _066168_, _066169_, _066170_, _066171_, _066172_, _066173_, _066174_, _066175_, _066176_, _066177_, _066178_, _066179_, _066180_, _066181_, _066182_, _066183_, _066184_, _066185_, _066186_, _066187_, _066188_, _066189_, _066190_, _066191_, _066192_, _066193_, _066194_, _066195_, _066196_, _066197_, _066198_, _066199_, _066200_, _066201_, _066202_, _066203_, _066204_, _066205_, _066206_, _066207_, _066208_, _066209_, _066210_, _066211_, _066212_, _066213_, _066214_, _066215_, _066216_, _066217_, _066218_, _066219_, _066220_, _066221_, _066222_, _066223_, _066224_, _066225_, _066226_, _066227_, _066228_, _066229_, _066230_, _066231_, _066232_, _066233_, _066234_, _066235_, _066236_, _066237_, _066238_, _066239_, _066240_, _066241_, _066242_, _066243_, _066244_, _066245_, _066246_, _066247_, _066248_, _066249_, _066250_, _066251_, _066252_, _066253_, _066254_, _066255_, _066256_, _066257_, _066258_, _066259_, _066260_, _066261_, _066262_, _066263_, _066264_, _066265_, _066266_, _066267_, _066268_, _066269_, _066270_, _066271_, _066272_, _066273_, _066274_, _066275_, _066276_, _066277_, _066278_, _066279_, _066280_, _066281_, _066282_, _066283_, _066284_, _066285_, _066286_, _066287_, _066288_, _066289_, _066290_, _066291_, _066292_, _066293_, _066294_, _066295_, _066296_, _066297_, _066298_, _066299_, _066300_, _066301_, _066302_, _066303_, _066304_, _066305_, _066306_, _066307_, _066308_, _066309_, _066310_, _066311_, _066312_, _066313_, _066314_, _066315_, _066316_, _066317_, _066318_, _066319_, _066320_, _066321_, _066322_, _066323_, _066324_, _066325_, _066326_, _066327_, _066328_, _066329_, _066330_, _066331_, _066332_, _066333_, _066334_, _066335_, _066336_, _066337_, _066338_, _066339_, _066340_, _066341_, _066342_, _066343_, _066344_, _066345_, _066346_, _066347_, _066348_, _066349_, _066350_, _066351_, _066352_, _066353_, _066354_, _066355_, _066356_, _066357_, _066358_, _066359_, _066360_, _066361_, _066362_, _066363_, _066364_, _066365_, _066366_, _066367_, _066368_, _066369_, _066370_, _066371_, _066372_, _066373_, _066374_, _066375_, _066376_, _066377_, _066378_, _066379_, _066380_, _066381_, _066382_, _066383_, _066384_, _066385_, _066386_, _066387_, _066388_, _066389_, _066390_, _066391_, _066392_, _066393_, _066394_, _066395_, _066396_, _066397_, _066398_, _066399_, _066400_, _066401_, _066402_, _066403_, _066404_, _066405_, _066406_, _066407_, _066408_, _066409_, _066410_, _066411_, _066412_, _066413_, _066414_, _066415_, _066416_, _066417_, _066418_, _066419_, _066420_, _066421_, _066422_, _066423_, _066424_, _066425_, _066426_, _066427_, _066428_, _066429_, _066430_, _066431_, _066432_, _066433_, _066434_, _066435_, _066436_, _066437_, _066438_, _066439_, _066440_, _066441_, _066442_, _066443_, _066444_, _066445_, _066446_, _066447_, _066448_, _066449_, _066450_, _066451_, _066452_, _066453_, _066454_, _066455_, _066456_, _066457_, _066458_, _066459_, _066460_, _066461_, _066462_, _066463_, _066464_, _066465_, _066466_, _066467_, _066468_, _066469_, _066470_, _066471_, _066472_, _066473_, _066474_, _066475_, _066476_, _066477_, _066478_, _066479_, _066480_, _066481_, _066482_, _066483_, _066484_, _066485_, _066486_, _066487_, _066488_, _066489_, _066490_, _066491_, _066492_, _066493_, _066494_, _066495_, _066496_, _066497_, _066498_, _066499_, _066500_, _066501_, _066502_, _066503_, _066504_, _066505_, _066506_, _066507_, _066508_, _066509_, _066510_, _066511_, _066512_, _066513_, _066514_, _066515_, _066516_, _066517_, _066518_, _066519_, _066520_, _066521_, _066522_, _066523_, _066524_, _066525_, _066526_, _066527_, _066528_, _066529_, _066530_, _066531_, _066532_, _066533_, _066534_, _066535_, _066536_, _066537_, _066538_, _066539_, _066540_, _066541_, _066542_, _066543_, _066544_, _066545_, _066546_, _066547_, _066548_, _066549_, _066550_, _066551_, _066552_, _066553_, _066554_, _066555_, _066556_, _066557_, _066558_, _066559_, _066560_, _066561_, _066562_, _066563_, _066564_, _066565_, _066566_, _066567_, _066568_, _066569_, _066570_, _066571_, _066572_, _066573_, _066574_, _066575_, _066576_, _066577_, _066578_, _066579_, _066580_, _066581_, _066582_, _066583_, _066584_, _066585_, _066586_, _066587_, _066588_, _066589_, _066590_, _066591_, _066592_, _066593_, _066594_, _066595_, _066596_, _066597_, _066598_, _066599_, _066600_, _066601_, _066602_, _066603_, _066604_, _066605_, _066606_, _066607_, _066608_, _066609_, _066610_, _066611_, _066612_, _066613_, _066614_, _066615_, _066616_, _066617_, _066618_, _066619_, _066620_, _066621_, _066622_, _066623_, _066624_, _066625_, _066626_, _066627_, _066628_, _066629_, _066630_, _066631_, _066632_, _066633_, _066634_, _066635_, _066636_, _066637_, _066638_, _066639_, _066640_, _066641_, _066642_, _066643_, _066644_, _066645_, _066646_, _066647_, _066648_, _066649_, _066650_, _066651_, _066652_, _066653_, _066654_, _066655_, _066656_, _066657_, _066658_, _066659_, _066660_, _066661_, _066662_, _066663_, _066664_, _066665_, _066666_, _066667_, _066668_, _066669_, _066670_, _066671_, _066672_, _066673_, _066674_, _066675_, _066676_, _066677_, _066678_, _066679_, _066680_, _066681_, _066682_, _066683_, _066684_, _066685_, _066686_, _066687_, _066688_, _066689_, _066690_, _066691_, _066692_, _066693_, _066694_, _066695_, _066696_, _066697_, _066698_, _066699_, _066700_, _066701_, _066702_, _066703_, _066704_, _066705_, _066706_, _066707_, _066708_, _066709_, _066710_, _066711_, _066712_, _066713_, _066714_, _066715_, _066716_, _066717_, _066718_, _066719_, _066720_, _066721_, _066722_, _066723_, _066724_, _066725_, _066726_, _066727_, _066728_, _066729_, _066730_, _066731_, _066732_, _066733_, _066734_, _066735_, _066736_, _066737_, _066738_, _066739_, _066740_, _066741_, _066742_, _066743_, _066744_, _066745_, _066746_, _066747_, _066748_, _066749_, _066750_, _066751_, _066752_, _066753_, _066754_, _066755_, _066756_, _066757_, _066758_, _066759_, _066760_, _066761_, _066762_, _066763_, _066764_, _066765_, _066766_, _066767_, _066768_, _066769_, _066770_, _066771_, _066772_, _066773_, _066774_, _066775_, _066776_, _066777_, _066778_, _066779_, _066780_, _066781_, _066782_, _066783_, _066784_, _066785_, _066786_, _066787_, _066788_, _066789_, _066790_, _066791_, _066792_, _066793_, _066794_, _066795_, _066796_, _066797_, _066798_, _066799_, _066800_, _066801_, _066802_, _066803_, _066804_, _066805_, _066806_, _066807_, _066808_, _066809_, _066810_, _066811_, _066812_, _066813_, _066814_, _066815_, _066816_, _066817_, _066818_, _066819_, _066820_, _066821_, _066822_, _066823_, _066824_, _066825_, _066826_, _066827_, _066828_, _066829_, _066830_, _066831_, _066832_, _066833_, _066834_, _066835_, _066836_, _066837_, _066838_, _066839_, _066840_, _066841_, _066842_, _066843_, _066844_, _066845_, _066846_, _066847_, _066848_, _066849_, _066850_, _066851_, _066852_, _066853_, _066854_, _066855_, _066856_, _066857_, _066858_, _066859_, _066860_, _066861_, _066862_, _066863_, _066864_, _066865_, _066866_, _066867_, _066868_, _066869_, _066870_, _066871_, _066872_, _066873_, _066874_, _066875_, _066876_, _066877_, _066878_, _066879_, _066880_, _066881_, _066882_, _066883_, _066884_, _066885_, _066886_, _066887_, _066888_, _066889_, _066890_, _066891_, _066892_, _066893_, _066894_, _066895_, _066896_, _066897_, _066898_, _066899_, _066900_, _066901_, _066902_, _066903_, _066904_, _066905_, _066906_, _066907_, _066908_, _066909_, _066910_, _066911_, _066912_, _066913_, _066914_, _066915_, _066916_, _066917_, _066918_, _066919_, _066920_, _066921_, _066922_, _066923_, _066924_, _066925_, _066926_, _066927_, _066928_, _066929_, _066930_, _066931_, _066932_, _066933_, _066934_, _066935_, _066936_, _066937_, _066938_, _066939_, _066940_, _066941_, _066942_, _066943_, _066944_, _066945_, _066946_, _066947_, _066948_, _066949_, _066950_, _066951_, _066952_, _066953_, _066954_, _066955_, _066956_, _066957_, _066958_, _066959_, _066960_, _066961_, _066962_, _066963_, _066964_, _066965_, _066966_, _066967_, _066968_, _066969_, _066970_, _066971_, _066972_, _066973_, _066974_, _066975_, _066976_, _066977_, _066978_, _066979_, _066980_, _066981_, _066982_, _066983_, _066984_, _066985_, _066986_, _066987_, _066988_, _066989_, _066990_, _066991_, _066992_, _066993_, _066994_, _066995_, _066996_, _066997_, _066998_, _066999_, _067000_, _067001_, _067002_, _067003_, _067004_, _067005_, _067006_, _067007_, _067008_, _067009_, _067010_, _067011_, _067012_, _067013_, _067014_, _067015_, _067016_, _067017_, _067018_, _067019_, _067020_, _067021_, _067022_, _067023_, _067024_, _067025_, _067026_, _067027_, _067028_, _067029_, _067030_, _067031_, _067032_, _067033_, _067034_, _067035_, _067036_, _067037_, _067038_, _067039_, _067040_, _067041_, _067042_, _067043_, _067044_, _067045_, _067046_, _067047_, _067048_, _067049_, _067050_, _067051_, _067052_, _067053_, _067054_, _067055_, _067056_, _067057_, _067058_, _067059_, _067060_, _067061_, _067062_, _067063_, _067064_, _067065_, _067066_, _067067_, _067068_, _067069_, _067070_, _067071_, _067072_, _067073_, _067074_, _067075_, _067076_, _067077_, _067078_, _067079_, _067080_, _067081_, _067082_, _067083_, _067084_, _067085_, _067086_, _067087_, _067088_, _067089_, _067090_, _067091_, _067092_, _067093_, _067094_, _067095_, _067096_, _067097_, _067098_, _067099_, _067100_, _067101_, _067102_, _067103_, _067104_, _067105_, _067106_, _067107_, _067108_, _067109_, _067110_, _067111_, _067112_, _067113_, _067114_, _067115_, _067116_, _067117_, _067118_, _067119_, _067120_, _067121_, _067122_, _067123_, _067124_, _067125_, _067126_, _067127_, _067128_, _067129_, _067130_, _067131_, _067132_, _067133_, _067134_, _067135_, _067136_, _067137_, _067138_, _067139_, _067140_, _067141_, _067142_, _067143_, _067144_, _067145_, _067146_, _067147_, _067148_, _067149_, _067150_, _067151_, _067152_, _067153_, _067154_, _067155_, _067156_, _067157_, _067158_, _067159_, _067160_, _067161_, _067162_, _067163_, _067164_, _067165_, _067166_, _067167_, _067168_, _067169_, _067170_, _067171_, _067172_, _067173_, _067174_, _067175_, _067176_, _067177_, _067178_, _067179_, _067180_, _067181_, _067182_, _067183_, _067184_, _067185_, _067186_, _067187_, _067188_, _067189_, _067190_, _067191_, _067192_, _067193_, _067194_, _067195_, _067196_, _067197_, _067198_, _067199_, _067200_, _067201_, _067202_, _067203_, _067204_, _067205_, _067206_, _067207_, _067208_, _067209_, _067210_, _067211_, _067212_, _067213_, _067214_, _067215_, _067216_, _067217_, _067218_, _067219_, _067220_, _067221_, _067222_, _067223_, _067224_, _067225_, _067226_, _067227_, _067228_, _067229_, _067230_, _067231_, _067232_, _067233_, _067234_, _067235_, _067236_, _067237_, _067238_, _067239_, _067240_, _067241_, _067242_, _067243_, _067244_, _067245_, _067246_, _067247_, _067248_, _067249_, _067250_, _067251_, _067252_, _067253_, _067254_, _067255_, _067256_, _067257_, _067258_, _067259_, _067260_, _067261_, _067262_, _067263_, _067264_, _067265_, _067266_, _067267_, _067268_, _067269_, _067270_, _067271_, _067272_, _067273_, _067274_, _067275_, _067276_, _067277_, _067278_, _067279_, _067280_, _067281_, _067282_, _067283_, _067284_, _067285_, _067286_, _067287_, _067288_, _067289_, _067290_, _067291_, _067292_, _067293_, _067294_, _067295_, _067296_, _067297_, _067298_, _067299_, _067300_, _067301_, _067302_, _067303_, _067304_, _067305_, _067306_, _067307_, _067308_, _067309_, _067310_, _067311_, _067312_, _067313_, _067314_, _067315_, _067316_, _067317_, _067318_, _067319_, _067320_, _067321_, _067322_, _067323_, _067324_, _067325_, _067326_, _067327_, _067328_, _067329_, _067330_, _067331_, _067332_, _067333_, _067334_, _067335_, _067336_, _067337_, _067338_, _067339_, _067340_, _067341_, _067342_, _067343_, _067344_, _067345_, _067346_, _067347_, _067348_, _067349_, _067350_, _067351_, _067352_, _067353_, _067354_, _067355_, _067356_, _067357_, _067358_, _067359_, _067360_, _067361_, _067362_, _067363_, _067364_, _067365_, _067366_, _067367_, _067368_, _067369_, _067370_, _067371_, _067372_, _067373_, _067374_, _067375_, _067376_, _067377_, _067378_, _067379_, _067380_, _067381_, _067382_, _067383_, _067384_, _067385_, _067386_, _067387_, _067388_, _067389_, _067390_, _067391_, _067392_, _067393_, _067394_, _067395_, _067396_, _067397_, _067398_, _067399_, _067400_, _067401_, _067402_, _067403_, _067404_, _067405_, _067406_, _067407_, _067408_, _067409_, _067410_, _067411_, _067412_, _067413_, _067414_, _067415_, _067416_, _067417_, _067418_, _067419_, _067420_, _067421_, _067422_, _067423_, _067424_, _067425_, _067426_, _067427_, _067428_, _067429_, _067430_, _067431_, _067432_, _067433_, _067434_, _067435_, _067436_, _067437_, _067438_, _067439_, _067440_, _067441_, _067442_, _067443_, _067444_, _067445_, _067446_, _067447_, _067448_, _067449_, _067450_, _067451_, _067452_, _067453_, _067454_, _067455_, _067456_, _067457_, _067458_, _067459_, _067460_, _067461_, _067462_, _067463_, _067464_, _067465_, _067466_, _067467_, _067468_, _067469_, _067470_, _067471_, _067472_, _067473_, _067474_, _067475_, _067476_, _067477_, _067478_, _067479_, _067480_, _067481_, _067482_, _067483_, _067484_, _067485_, _067486_, _067487_, _067488_, _067489_, _067490_, _067491_, _067492_, _067493_, _067494_, _067495_, _067496_, _067497_, _067498_, _067499_, _067500_, _067501_, _067502_, _067503_, _067504_, _067505_, _067506_, _067507_, _067508_, _067509_, _067510_, _067511_, _067512_, _067513_, _067514_, _067515_, _067516_, _067517_, _067518_, _067519_, _067520_, _067521_, _067522_, _067523_, _067524_, _067525_, _067526_, _067527_, _067528_, _067529_, _067530_, _067531_, _067532_, _067533_, _067534_, _067535_, _067536_, _067537_, _067538_, _067539_, _067540_, _067541_, _067542_, _067543_, _067544_, _067545_, _067546_, _067547_, _067548_, _067549_, _067550_, _067551_, _067552_, _067553_, _067554_, _067555_, _067556_, _067557_, _067558_, _067559_, _067560_, _067561_, _067562_, _067563_, _067564_, _067565_, _067566_, _067567_, _067568_, _067569_, _067570_, _067571_, _067572_, _067573_, _067574_, _067575_, _067576_, _067577_, _067578_, _067579_, _067580_, _067581_, _067582_, _067583_, _067584_, _067585_, _067586_, _067587_, _067588_, _067589_, _067590_, _067591_, _067592_, _067593_, _067594_, _067595_, _067596_, _067597_, _067598_, _067599_, _067600_, _067601_, _067602_, _067603_, _067604_, _067605_, _067606_, _067607_, _067608_, _067609_, _067610_, _067611_, _067612_, _067613_, _067614_, _067615_, _067616_, _067617_, _067618_, _067619_, _067620_, _067621_, _067622_, _067623_, _067624_, _067625_, _067626_, _067627_, _067628_, _067629_, _067630_, _067631_, _067632_, _067633_, _067634_, _067635_, _067636_, _067637_, _067638_, _067639_, _067640_, _067641_, _067642_, _067643_, _067644_, _067645_, _067646_, _067647_, _067648_, _067649_, _067650_, _067651_, _067652_, _067653_, _067654_, _067655_, _067656_, _067657_, _067658_, _067659_, _067660_, _067661_, _067662_, _067663_, _067664_, _067665_, _067666_, _067667_, _067668_, _067669_, _067670_, _067671_, _067672_, _067673_, _067674_, _067675_, _067676_, _067677_, _067678_, _067679_, _067680_, _067681_, _067682_, _067683_, _067684_, _067685_, _067686_, _067687_, _067688_, _067689_, _067690_, _067691_, _067692_, _067693_, _067694_, _067695_, _067696_, _067697_, _067698_, _067699_, _067700_, _067701_, _067702_, _067703_, _067704_, _067705_, _067706_, _067707_, _067708_, _067709_, _067710_, _067711_, _067712_, _067713_, _067714_, _067715_, _067716_, _067717_, _067718_, _067719_, _067720_, _067721_, _067722_, _067723_, _067724_, _067725_, _067726_, _067727_, _067728_, _067729_, _067730_, _067731_, _067732_, _067733_, _067734_, _067735_, _067736_, _067737_, _067738_, _067739_, _067740_, _067741_, _067742_, _067743_, _067744_, _067745_, _067746_, _067747_, _067748_, _067749_, _067750_, _067751_, _067752_, _067753_, _067754_, _067755_, _067756_, _067757_, _067758_, _067759_, _067760_, _067761_, _067762_, _067763_, _067764_, _067765_, _067766_, _067767_, _067768_, _067769_, _067770_, _067771_, _067772_, _067773_, _067774_, _067775_, _067776_, _067777_, _067778_, _067779_, _067780_, _067781_, _067782_, _067783_, _067784_, _067785_, _067786_, _067787_, _067788_, _067789_, _067790_, _067791_, _067792_, _067793_, _067794_, _067795_, _067796_, _067797_, _067798_, _067799_, _067800_, _067801_, _067802_, _067803_, _067804_, _067805_, _067806_, _067807_, _067808_, _067809_, _067810_, _067811_, _067812_, _067813_, _067814_, _067815_, _067816_, _067817_, _067818_, _067819_, _067820_, _067821_, _067822_, _067823_, _067824_, _067825_, _067826_, _067827_, _067828_, _067829_, _067830_, _067831_, _067832_, _067833_, _067834_, _067835_, _067836_, _067837_, _067838_, _067839_, _067840_, _067841_, _067842_, _067843_, _067844_, _067845_, _067846_, _067847_, _067848_, _067849_, _067850_, _067851_, _067852_, _067853_, _067854_, _067855_, _067856_, _067857_, _067858_, _067859_, _067860_, _067861_, _067862_, _067863_, _067864_, _067865_, _067866_, _067867_, _067868_, _067869_, _067870_, _067871_, _067872_, _067873_, _067874_, _067875_, _067876_, _067877_, _067878_, _067879_, _067880_, _067881_, _067882_, _067883_, _067884_, _067885_, _067886_, _067887_, _067888_, _067889_, _067890_, _067891_, _067892_, _067893_, _067894_, _067895_, _067896_, _067897_, _067898_, _067899_, _067900_, _067901_, _067902_, _067903_, _067904_, _067905_, _067906_, _067907_, _067908_, _067909_, _067910_, _067911_, _067912_, _067913_, _067914_, _067915_, _067916_, _067917_, _067918_, _067919_, _067920_, _067921_, _067922_, _067923_, _067924_, _067925_, _067926_, _067927_, _067928_, _067929_, _067930_, _067931_, _067932_, _067933_, _067934_, _067935_, _067936_, _067937_, _067938_, _067939_, _067940_, _067941_, _067942_, _067943_, _067944_, _067945_, _067946_, _067947_, _067948_, _067949_, _067950_, _067951_, _067952_, _067953_, _067954_, _067955_, _067956_, _067957_, _067958_, _067959_, _067960_, _067961_, _067962_, _067963_, _067964_, _067965_, _067966_, _067967_, _067968_, _067969_, _067970_, _067971_, _067972_, _067973_, _067974_, _067975_, _067976_, _067977_, _067978_, _067979_, _067980_, _067981_, _067982_, _067983_, _067984_, _067985_, _067986_, _067987_, _067988_, _067989_, _067990_, _067991_, _067992_, _067993_, _067994_, _067995_, _067996_, _067997_, _067998_, _067999_, _068000_, _068001_, _068002_, _068003_, _068004_, _068005_, _068006_, _068007_, _068008_, _068009_, _068010_, _068011_, _068012_, _068013_, _068014_, _068015_, _068016_, _068017_, _068018_, _068019_, _068020_, _068021_, _068022_, _068023_, _068024_, _068025_, _068026_, _068027_, _068028_, _068029_, _068030_, _068031_, _068032_, _068033_, _068034_, _068035_, _068036_, _068037_, _068038_, _068039_, _068040_, _068041_, _068042_, _068043_, _068044_, _068045_, _068046_, _068047_, _068048_, _068049_, _068050_, _068051_, _068052_, _068053_, _068054_, _068055_, _068056_, _068057_, _068058_, _068059_, _068060_, _068061_, _068062_, _068063_, _068064_, _068065_, _068066_, _068067_, _068068_, _068069_, _068070_, _068071_, _068072_, _068073_, _068074_, _068075_, _068076_, _068077_, _068078_, _068079_, _068080_, _068081_, _068082_, _068083_, _068084_, _068085_, _068086_, _068087_, _068088_, _068089_, _068090_, _068091_, _068092_, _068093_, _068094_, _068095_, _068096_, _068097_, _068098_, _068099_, _068100_, _068101_, _068102_, _068103_, _068104_, _068105_, _068106_, _068107_, _068108_, _068109_, _068110_, _068111_, _068112_, _068113_, _068114_, _068115_, _068116_, _068117_, _068118_, _068119_, _068120_, _068121_, _068122_, _068123_, _068124_, _068125_, _068126_, _068127_, _068128_, _068129_, _068130_, _068131_, _068132_, _068133_, _068134_, _068135_, _068136_, _068137_, _068138_, _068139_, _068140_, _068141_, _068142_, _068143_, _068144_, _068145_, _068146_, _068147_, _068148_, _068149_, _068150_, _068151_, _068152_, _068153_, _068154_, _068155_, _068156_, _068157_, _068158_, _068159_, _068160_, _068161_, _068162_, _068163_, _068164_, _068165_, _068166_, _068167_, _068168_, _068169_, _068170_, _068171_, _068172_, _068173_, _068174_, _068175_, _068176_, _068177_, _068178_, _068179_, _068180_, _068181_, _068182_, _068183_, _068184_, _068185_, _068186_, _068187_, _068188_, _068189_, _068190_, _068191_, _068192_, _068193_, _068194_, _068195_, _068196_, _068197_, _068198_, _068199_, _068200_, _068201_, _068202_, _068203_, _068204_, _068205_, _068206_, _068207_, _068208_, _068209_, _068210_, _068211_, _068212_, _068213_, _068214_, _068215_, _068216_, _068217_, _068218_, _068219_, _068220_, _068221_, _068222_, _068223_, _068224_, _068225_, _068226_, _068227_, _068228_, _068229_, _068230_, _068231_, _068232_, _068233_, _068234_, _068235_, _068236_, _068237_, _068238_, _068239_, _068240_, _068241_, _068242_, _068243_, _068244_, _068245_, _068246_, _068247_, _068248_, _068249_, _068250_, _068251_, _068252_, _068253_, _068254_, _068255_, _068256_, _068257_, _068258_, _068259_, _068260_, _068261_, _068262_, _068263_, _068264_, _068265_, _068266_, _068267_, _068268_, _068269_, _068270_, _068271_, _068272_, _068273_, _068274_, _068275_, _068276_, _068277_, _068278_, _068279_, _068280_, _068281_, _068282_, _068283_, _068284_, _068285_, _068286_, _068287_, _068288_, _068289_, _068290_, _068291_, _068292_, _068293_, _068294_, _068295_, _068296_, _068297_, _068298_, _068299_, _068300_, _068301_, _068302_, _068303_, _068304_, _068305_, _068306_, _068307_, _068308_, _068309_, _068310_, _068311_, _068312_, _068313_, _068314_, _068315_, _068316_, _068317_, _068318_, _068319_, _068320_, _068321_, _068322_, _068323_, _068324_, _068325_, _068326_, _068327_, _068328_, _068329_, _068330_, _068331_, _068332_, _068333_, _068334_, _068335_, _068336_, _068337_, _068338_, _068339_, _068340_, _068341_, _068342_, _068343_, _068344_, _068345_, _068346_, _068347_, _068348_, _068349_, _068350_, _068351_, _068352_, _068353_, _068354_, _068355_, _068356_, _068357_, _068358_, _068359_, _068360_, _068361_, _068362_, _068363_, _068364_, _068365_, _068366_, _068367_, _068368_, _068369_, _068370_, _068371_, _068372_, _068373_, _068374_, _068375_, _068376_, _068377_, _068378_, _068379_, _068380_, _068381_, _068382_, _068383_, _068384_, _068385_, _068386_, _068387_, _068388_, _068389_, _068390_, _068391_, _068392_, _068393_, _068394_, _068395_, _068396_, _068397_, _068398_, _068399_, _068400_, _068401_, _068402_, _068403_, _068404_, _068405_, _068406_, _068407_, _068408_, _068409_, _068410_, _068411_, _068412_, _068413_, _068414_, _068415_, _068416_, _068417_, _068418_, _068419_, _068420_, _068421_, _068422_, _068423_, _068424_, _068425_, _068426_, _068427_, _068428_, _068429_, _068430_, _068431_, _068432_, _068433_, _068434_, _068435_, _068436_, _068437_, _068438_, _068439_, _068440_, _068441_, _068442_, _068443_, _068444_, _068445_, _068446_, _068447_, _068448_, _068449_, _068450_, _068451_, _068452_, _068453_, _068454_, _068455_, _068456_, _068457_, _068458_, _068459_, _068460_, _068461_, _068462_, _068463_, _068464_, _068465_, _068466_, _068467_, _068468_, _068469_, _068470_, _068471_, _068472_, _068473_, _068474_, _068475_, _068476_, _068477_, _068478_, _068479_, _068480_, _068481_, _068482_, _068483_, _068484_, _068485_, _068486_, _068487_, _068488_, _068489_, _068490_, _068491_, _068492_, _068493_, _068494_, _068495_, _068496_, _068497_, _068498_, _068499_, _068500_, _068501_, _068502_, _068503_, _068504_, _068505_, _068506_, _068507_, _068508_, _068509_, _068510_, _068511_, _068512_, _068513_, _068514_, _068515_, _068516_, _068517_, _068518_, _068519_, _068520_, _068521_, _068522_, _068523_, _068524_, _068525_, _068526_, _068527_, _068528_, _068529_, _068530_, _068531_, _068532_, _068533_, _068534_, _068535_, _068536_, _068537_, _068538_, _068539_, _068540_, _068541_, _068542_, _068543_, _068544_, _068545_, _068546_, _068547_, _068548_, _068549_, _068550_, _068551_, _068552_, _068553_, _068554_, _068555_, _068556_, _068557_, _068558_, _068559_, _068560_, _068561_, _068562_, _068563_, _068564_, _068565_, _068566_, _068567_, _068568_, _068569_, _068570_, _068571_, _068572_, _068573_, _068574_, _068575_, _068576_, _068577_, _068578_, _068579_, _068580_, _068581_, _068582_, _068583_, _068584_, _068585_, _068586_, _068587_, _068588_, _068589_, _068590_, _068591_, _068592_, _068593_, _068594_, _068595_, _068596_, _068597_, _068598_, _068599_, _068600_, _068601_, _068602_, _068603_, _068604_, _068605_, _068606_, _068607_, _068608_, _068609_, _068610_, _068611_, _068612_, _068613_, _068614_, _068615_, _068616_, _068617_, _068618_, _068619_, _068620_, _068621_, _068622_, _068623_, _068624_, _068625_, _068626_, _068627_, _068628_, _068629_, _068630_, _068631_, _068632_, _068633_, _068634_, _068635_, _068636_, _068637_, _068638_, _068639_, _068640_, _068641_, _068642_, _068643_, _068644_, _068645_, _068646_, _068647_, _068648_, _068649_, _068650_, _068651_, _068652_, _068653_, _068654_, _068655_, _068656_, _068657_, _068658_, _068659_, _068660_, _068661_, _068662_, _068663_, _068664_, _068665_, _068666_, _068667_, _068668_, _068669_, _068670_, _068671_, _068672_, _068673_, _068674_, _068675_, _068676_, _068677_, _068678_, _068679_, _068680_, _068681_, _068682_, _068683_, _068684_, _068685_, _068686_, _068687_, _068688_, _068689_, _068690_, _068691_, _068692_, _068693_, _068694_, _068695_, _068696_, _068697_, _068698_, _068699_, _068700_, _068701_, _068702_, _068703_, _068704_, _068705_, _068706_, _068707_, _068708_, _068709_, _068710_, _068711_, _068712_, _068713_, _068714_, _068715_, _068716_, _068717_, _068718_, _068719_, _068720_, _068721_, _068722_, _068723_, _068724_, _068725_, _068726_, _068727_, _068728_, _068729_, _068730_, _068731_, _068732_, _068733_, _068734_, _068735_, _068736_, _068737_, _068738_, _068739_, _068740_, _068741_, _068742_, _068743_, _068744_, _068745_, _068746_, _068747_, _068748_, _068749_, _068750_, _068751_, _068752_, _068753_, _068754_, _068755_, _068756_, _068757_, _068758_, _068759_, _068760_, _068761_, _068762_, _068763_, _068764_, _068765_, _068766_, _068767_, _068768_, _068769_, _068770_, _068771_, _068772_, _068773_, _068774_, _068775_, _068776_, _068777_, _068778_, _068779_, _068780_, _068781_, _068782_, _068783_, _068784_, _068785_, _068786_, _068787_, _068788_, _068789_, _068790_, _068791_, _068792_, _068793_, _068794_, _068795_, _068796_, _068797_, _068798_, _068799_, _068800_, _068801_, _068802_, _068803_, _068804_, _068805_, _068806_, _068807_, _068808_, _068809_, _068810_, _068811_, _068812_, _068813_, _068814_, _068815_, _068816_, _068817_, _068818_, _068819_, _068820_, _068821_, _068822_, _068823_, _068824_, _068825_, _068826_, _068827_, _068828_, _068829_, _068830_, _068831_, _068832_, _068833_, _068834_, _068835_, _068836_, _068837_, _068838_, _068839_, _068840_, _068841_, _068842_, _068843_, _068844_, _068845_, _068846_, _068847_, _068848_, _068849_, _068850_, _068851_, _068852_, _068853_, _068854_, _068855_, _068856_, _068857_, _068858_, _068859_, _068860_, _068861_, _068862_, _068863_, _068864_, _068865_, _068866_, _068867_, _068868_, _068869_, _068870_, _068871_, _068872_, _068873_, _068874_, _068875_, _068876_, _068877_, _068878_, _068879_, _068880_, _068881_, _068882_, _068883_, _068884_, _068885_, _068886_, _068887_, _068888_, _068889_, _068890_, _068891_, _068892_, _068893_, _068894_, _068895_, _068896_, _068897_, _068898_, _068899_, _068900_, _068901_, _068902_, _068903_, _068904_, _068905_, _068906_, _068907_, _068908_, _068909_, _068910_, _068911_, _068912_, _068913_, _068914_, _068915_, _068916_, _068917_, _068918_, _068919_, _068920_, _068921_, _068922_, _068923_, _068924_, _068925_, _068926_, _068927_, _068928_, _068929_, _068930_, _068931_, _068932_, _068933_, _068934_, _068935_, _068936_, _068937_, _068938_, _068939_, _068940_, _068941_, _068942_, _068943_, _068944_, _068945_, _068946_, _068947_, _068948_, _068949_, _068950_, _068951_, _068952_, _068953_, _068954_, _068955_, _068956_, _068957_, _068958_, _068959_, _068960_, _068961_, _068962_, _068963_, _068964_, _068965_, _068966_, _068967_, _068968_, _068969_, _068970_, _068971_, _068972_, _068973_, _068974_, _068975_, _068976_, _068977_, _068978_, _068979_, _068980_, _068981_, _068982_, _068983_, _068984_, _068985_, _068986_, _068987_, _068988_, _068989_, _068990_, _068991_, _068992_, _068993_, _068994_, _068995_, _068996_, _068997_, _068998_, _068999_, _069000_, _069001_, _069002_, _069003_, _069004_, _069005_, _069006_, _069007_, _069008_, _069009_, _069010_, _069011_, _069012_, _069013_, _069014_, _069015_, _069016_, _069017_, _069018_, _069019_, _069020_, _069021_, _069022_, _069023_, _069024_, _069025_, _069026_, _069027_, _069028_, _069029_, _069030_, _069031_, _069032_, _069033_, _069034_, _069035_, _069036_, _069037_, _069038_, _069039_, _069040_, _069041_, _069042_, _069043_, _069044_, _069045_, _069046_, _069047_, _069048_, _069049_, _069050_, _069051_, _069052_, _069053_, _069054_, _069055_, _069056_, _069057_, _069058_, _069059_, _069060_, _069061_, _069062_, _069063_, _069064_, _069065_, _069066_, _069067_, _069068_, _069069_, _069070_, _069071_, _069072_, _069073_, _069074_, _069075_, _069076_, _069077_, _069078_, _069079_, _069080_, _069081_, _069082_, _069083_, _069084_, _069085_, _069086_, _069087_, _069088_, _069089_, _069090_, _069091_, _069092_, _069093_, _069094_, _069095_, _069096_, _069097_, _069098_, _069099_, _069100_, _069101_, _069102_, _069103_, _069104_, _069105_, _069106_, _069107_, _069108_, _069109_, _069110_, _069111_, _069112_, _069113_, _069114_, _069115_, _069116_, _069117_, _069118_, _069119_, _069120_, _069121_, _069122_, _069123_, _069124_, _069125_, _069126_, _069127_, _069128_, _069129_, _069130_, _069131_, _069132_, _069133_, _069134_, _069135_, _069136_, _069137_, _069138_, _069139_, _069140_, _069141_, _069142_, _069143_, _069144_, _069145_, _069146_, _069147_, _069148_, _069149_, _069150_, _069151_, _069152_, _069153_, _069154_, _069155_, _069156_, _069157_, _069158_, _069159_, _069160_, _069161_, _069162_, _069163_, _069164_, _069165_, _069166_, _069167_, _069168_, _069169_, _069170_, _069171_, _069172_, _069173_, _069174_, _069175_, _069176_, _069177_, _069178_, _069179_, _069180_, _069181_, _069182_, _069183_, _069184_, _069185_, _069186_, _069187_, _069188_, _069189_, _069190_, _069191_, _069192_, _069193_, _069194_, _069195_, _069196_, _069197_, _069198_, _069199_, _069200_, _069201_, _069202_, _069203_, _069204_, _069205_, _069206_, _069207_, _069208_, _069209_, _069210_, _069211_, _069212_, _069213_, _069214_, _069215_, _069216_, _069217_, _069218_, _069219_, _069220_, _069221_, _069222_, _069223_, _069224_, _069225_, _069226_, _069227_, _069228_, _069229_, _069230_, _069231_, _069232_, _069233_, _069234_, _069235_, _069236_, _069237_, _069238_, _069239_, _069240_, _069241_, _069242_, _069243_, _069244_, _069245_, _069246_, _069247_, _069248_, _069249_, _069250_, _069251_, _069252_, _069253_, _069254_, _069255_, _069256_, _069257_, _069258_, _069259_, _069260_, _069261_, _069262_, _069263_, _069264_, _069265_, _069266_, _069267_, _069268_, _069269_, _069270_, _069271_, _069272_, _069273_, _069274_, _069275_, _069276_, _069277_, _069278_, _069279_, _069280_, _069281_, _069282_, _069283_, _069284_, _069285_, _069286_, _069287_, _069288_, _069289_, _069290_, _069291_, _069292_, _069293_, _069294_, _069295_, _069296_, _069297_, _069298_, _069299_, _069300_, _069301_, _069302_, _069303_, _069304_, _069305_, _069306_, _069307_, _069308_, _069309_, _069310_, _069311_, _069312_, _069313_, _069314_, _069315_, _069316_, _069317_, _069318_, _069319_, _069320_, _069321_, _069322_, _069323_, _069324_, _069325_, _069326_, _069327_, _069328_, _069329_, _069330_, _069331_, _069332_, _069333_, _069334_, _069335_, _069336_, _069337_, _069338_, _069339_, _069340_, _069341_, _069342_, _069343_, _069344_, _069345_, _069346_, _069347_, _069348_, _069349_, _069350_, _069351_, _069352_, _069353_, _069354_, _069355_, _069356_, _069357_, _069358_, _069359_, _069360_, _069361_, _069362_, _069363_, _069364_, _069365_, _069366_, _069367_, _069368_, _069369_, _069370_, _069371_, _069372_, _069373_, _069374_, _069375_, _069376_, _069377_, _069378_, _069379_, _069380_, _069381_, _069382_, _069383_, _069384_, _069385_, _069386_, _069387_, _069388_, _069389_, _069390_, _069391_, _069392_, _069393_, _069394_, _069395_, _069396_, _069397_, _069398_, _069399_, _069400_, _069401_, _069402_, _069403_, _069404_, _069405_, _069406_, _069407_, _069408_, _069409_, _069410_, _069411_, _069412_, _069413_, _069414_, _069415_, _069416_, _069417_, _069418_, _069419_, _069420_, _069421_, _069422_, _069423_, _069424_, _069425_, _069426_, _069427_, _069428_, _069429_, _069430_, _069431_, _069432_, _069433_, _069434_, _069435_, _069436_, _069437_, _069438_, _069439_, _069440_, _069441_, _069442_, _069443_, _069444_, _069445_, _069446_, _069447_, _069448_, _069449_, _069450_, _069451_, _069452_, _069453_, _069454_, _069455_, _069456_, _069457_, _069458_, _069459_, _069460_, _069461_, _069462_, _069463_, _069464_, _069465_, _069466_, _069467_, _069468_, _069469_, _069470_, _069471_, _069472_, _069473_, _069474_, _069475_, _069476_, _069477_, _069478_, _069479_, _069480_, _069481_, _069482_, _069483_, _069484_, _069485_, _069486_, _069487_, _069488_, _069489_, _069490_, _069491_, _069492_, _069493_, _069494_, _069495_, _069496_, _069497_, _069498_, _069499_, _069500_, _069501_, _069502_, _069503_, _069504_, _069505_, _069506_, _069507_, _069508_, _069509_, _069510_, _069511_, _069512_, _069513_, _069514_, _069515_, _069516_, _069517_, _069518_, _069519_, _069520_, _069521_, _069522_, _069523_, _069524_, _069525_, _069526_, _069527_, _069528_, _069529_, _069530_, _069531_, _069532_, _069533_, _069534_, _069535_, _069536_, _069537_, _069538_, _069539_, _069540_, _069541_, _069542_, _069543_, _069544_, _069545_, _069546_, _069547_, _069548_, _069549_, _069550_, _069551_, _069552_, _069553_, _069554_, _069555_, _069556_, _069557_, _069558_, _069559_, _069560_, _069561_, _069562_, _069563_, _069564_, _069565_, _069566_, _069567_, _069568_, _069569_, _069570_, _069571_, _069572_, _069573_, _069574_, _069575_, _069576_, _069577_, _069578_, _069579_, _069580_, _069581_, _069582_, _069583_, _069584_, _069585_, _069586_, _069587_, _069588_, _069589_, _069590_, _069591_, _069592_, _069593_, _069594_, _069595_, _069596_, _069597_, _069598_, _069599_, _069600_, _069601_, _069602_, _069603_, _069604_, _069605_, _069606_, _069607_, _069608_, _069609_, _069610_, _069611_, _069612_, _069613_, _069614_, _069615_, _069616_, _069617_, _069618_, _069619_, _069620_, _069621_, _069622_, _069623_, _069624_, _069625_, _069626_, _069627_, _069628_, _069629_, _069630_, _069631_, _069632_, _069633_, _069634_, _069635_, _069636_, _069637_, _069638_, _069639_, _069640_, _069641_, _069642_, _069643_, _069644_, _069645_, _069646_, _069647_, _069648_, _069649_, _069650_, _069651_, _069652_, _069653_, _069654_, _069655_, _069656_, _069657_, _069658_, _069659_, _069660_, _069661_, _069662_, _069663_, _069664_, _069665_, _069666_, _069667_, _069668_, _069669_, _069670_, _069671_, _069672_, _069673_, _069674_, _069675_, _069676_, _069677_, _069678_, _069679_, _069680_, _069681_, _069682_, _069683_, _069684_, _069685_, _069686_, _069687_, _069688_, _069689_, _069690_, _069691_, _069692_, _069693_, _069694_, _069695_, _069696_, _069697_, _069698_, _069699_, _069700_, _069701_, _069702_, _069703_, _069704_, _069705_, _069706_, _069707_, _069708_, _069709_, _069710_, _069711_, _069712_, _069713_, _069714_, _069715_, _069716_, _069717_, _069718_, _069719_, _069720_, _069721_, _069722_, _069723_, _069724_, _069725_, _069726_, _069727_, _069728_, _069729_, _069730_, _069731_, _069732_, _069733_, _069734_, _069735_, _069736_, _069737_, _069738_, _069739_, _069740_, _069741_, _069742_, _069743_, _069744_, _069745_, _069746_, _069747_, _069748_, _069749_, _069750_, _069751_, _069752_, _069753_, _069754_, _069755_, _069756_, _069757_, _069758_, _069759_, _069760_, _069761_, _069762_, _069763_, _069764_, _069765_, _069766_, _069767_, _069768_, _069769_, _069770_, _069771_, _069772_, _069773_, _069774_, _069775_, _069776_, _069777_, _069778_, _069779_, _069780_, _069781_, _069782_, _069783_, _069784_, _069785_, _069786_, _069787_, _069788_, _069789_, _069790_, _069791_, _069792_, _069793_, _069794_, _069795_, _069796_, _069797_, _069798_, _069799_, _069800_, _069801_, _069802_, _069803_, _069804_, _069805_, _069806_, _069807_, _069808_, _069809_, _069810_, _069811_, _069812_, _069813_, _069814_, _069815_, _069816_, _069817_, _069818_, _069819_, _069820_, _069821_, _069822_, _069823_, _069824_, _069825_, _069826_, _069827_, _069828_, _069829_, _069830_, _069831_, _069832_, _069833_, _069834_, _069835_, _069836_, _069837_, _069838_, _069839_, _069840_, _069841_, _069842_, _069843_, _069844_, _069845_, _069846_, _069847_, _069848_, _069849_, _069850_, _069851_, _069852_, _069853_, _069854_, _069855_, _069856_, _069857_, _069858_, _069859_, _069860_, _069861_, _069862_, _069863_, _069864_, _069865_, _069866_, _069867_, _069868_, _069869_, _069870_, _069871_, _069872_, _069873_, _069874_, _069875_, _069876_, _069877_, _069878_, _069879_, _069880_, _069881_, _069882_, _069883_, _069884_, _069885_, _069886_, _069887_, _069888_, _069889_, _069890_, _069891_, _069892_, _069893_, _069894_, _069895_, _069896_, _069897_, _069898_, _069899_, _069900_, _069901_, _069902_, _069903_, _069904_, _069905_, _069906_, _069907_, _069908_, _069909_, _069910_, _069911_, _069912_, _069913_, _069914_, _069915_, _069916_, _069917_, _069918_, _069919_, _069920_, _069921_, _069922_, _069923_, _069924_, _069925_, _069926_, _069927_, _069928_, _069929_, _069930_, _069931_, _069932_, _069933_, _069934_, _069935_, _069936_, _069937_, _069938_, _069939_, _069940_, _069941_, _069942_, _069943_, _069944_, _069945_, _069946_, _069947_, _069948_, _069949_, _069950_, _069951_, _069952_, _069953_, _069954_, _069955_, _069956_, _069957_, _069958_, _069959_, _069960_, _069961_, _069962_, _069963_, _069964_, _069965_, _069966_, _069967_, _069968_, _069969_, _069970_, _069971_, _069972_, _069973_, _069974_, _069975_, _069976_, _069977_, _069978_, _069979_, _069980_, _069981_, _069982_, _069983_, _069984_, _069985_, _069986_, _069987_, _069988_, _069989_, _069990_, _069991_, _069992_, _069993_, _069994_, _069995_, _069996_, _069997_, _069998_, _069999_, _070000_, _070001_, _070002_, _070003_, _070004_, _070005_, _070006_, _070007_, _070008_, _070009_, _070010_, _070011_, _070012_, _070013_, _070014_, _070015_, _070016_, _070017_, _070018_, _070019_, _070020_, _070021_, _070022_, _070023_, _070024_, _070025_, _070026_, _070027_, _070028_, _070029_, _070030_, _070031_, _070032_, _070033_, _070034_, _070035_, _070036_, _070037_, _070038_, _070039_, _070040_, _070041_, _070042_, _070043_, _070044_, _070045_, _070046_, _070047_, _070048_, _070049_, _070050_, _070051_, _070052_, _070053_, _070054_, _070055_, _070056_, _070057_, _070058_, _070059_, _070060_, _070061_, _070062_, _070063_, _070064_, _070065_, _070066_, _070067_, _070068_, _070069_, _070070_, _070071_, _070072_, _070073_, _070074_, _070075_, _070076_, _070077_, _070078_, _070079_, _070080_, _070081_, _070082_, _070083_, _070084_, _070085_, _070086_, _070087_, _070088_, _070089_, _070090_, _070091_, _070092_, _070093_, _070094_, _070095_, _070096_, _070097_, _070098_, _070099_, _070100_, _070101_, _070102_, _070103_, _070104_, _070105_, _070106_, _070107_, _070108_, _070109_, _070110_, _070111_, _070112_, _070113_, _070114_, _070115_, _070116_, _070117_, _070118_, _070119_, _070120_, _070121_, _070122_, _070123_, _070124_, _070125_, _070126_, _070127_, _070128_, _070129_, _070130_, _070131_, _070132_, _070133_, _070134_, _070135_, _070136_, _070137_, _070138_, _070139_, _070140_, _070141_, _070142_, _070143_, _070144_, _070145_, _070146_, _070147_, _070148_, _070149_, _070150_, _070151_, _070152_, _070153_, _070154_, _070155_, _070156_, _070157_, _070158_, _070159_, _070160_, _070161_, _070162_, _070163_, _070164_, _070165_, _070166_, _070167_, _070168_, _070169_, _070170_, _070171_, _070172_, _070173_, _070174_, _070175_, _070176_, _070177_, _070178_, _070179_, _070180_, _070181_, _070182_, _070183_, _070184_, _070185_, _070186_, _070187_, _070188_, _070189_, _070190_, _070191_, _070192_, _070193_, _070194_, _070195_, _070196_, _070197_, _070198_, _070199_, _070200_, _070201_, _070202_, _070203_, _070204_, _070205_, _070206_, _070207_, _070208_, _070209_, _070210_, _070211_, _070212_, _070213_, _070214_, _070215_, _070216_, _070217_, _070218_, _070219_, _070220_, _070221_, _070222_, _070223_, _070224_, _070225_, _070226_, _070227_, _070228_, _070229_, _070230_, _070231_, _070232_, _070233_, _070234_, _070235_, _070236_, _070237_, _070238_, _070239_, _070240_, _070241_, _070242_, _070243_, _070244_, _070245_, _070246_, _070247_, _070248_, _070249_, _070250_, _070251_, _070252_, _070253_, _070254_, _070255_, _070256_, _070257_, _070258_, _070259_, _070260_, _070261_, _070262_, _070263_, _070264_, _070265_, _070266_, _070267_, _070268_, _070269_, _070270_, _070271_, _070272_, _070273_, _070274_, _070275_, _070276_, _070277_, _070278_, _070279_, _070280_, _070281_, _070282_, _070283_, _070284_, _070285_, _070286_, _070287_, _070288_, _070289_, _070290_, _070291_, _070292_, _070293_, _070294_, _070295_, _070296_, _070297_, _070298_, _070299_, _070300_, _070301_, _070302_, _070303_, _070304_, _070305_, _070306_, _070307_, _070308_, _070309_, _070310_, _070311_, _070312_, _070313_, _070314_, _070315_, _070316_, _070317_, _070318_, _070319_, _070320_, _070321_, _070322_, _070323_, _070324_, _070325_, _070326_, _070327_, _070328_, _070329_, _070330_, _070331_, _070332_, _070333_, _070334_, _070335_, _070336_, _070337_, _070338_, _070339_, _070340_, _070341_, _070342_, _070343_, _070344_, _070345_, _070346_, _070347_, _070348_, _070349_, _070350_, _070351_, _070352_, _070353_, _070354_, _070355_, _070356_, _070357_, _070358_, _070359_, _070360_, _070361_, _070362_, _070363_, _070364_, _070365_, _070366_, _070367_, _070368_, _070369_, _070370_, _070371_, _070372_, _070373_, _070374_, _070375_, _070376_, _070377_, _070378_, _070379_, _070380_, _070381_, _070382_, _070383_, _070384_, _070385_, _070386_, _070387_, _070388_, _070389_, _070390_, _070391_, _070392_, _070393_, _070394_, _070395_, _070396_, _070397_, _070398_, _070399_, _070400_, _070401_, _070402_, _070403_, _070404_, _070405_, _070406_, _070407_, _070408_, _070409_, _070410_, _070411_, _070412_, _070413_, _070414_, _070415_, _070416_, _070417_, _070418_, _070419_, _070420_, _070421_, _070422_, _070423_, _070424_, _070425_, _070426_, _070427_, _070428_, _070429_, _070430_, _070431_, _070432_, _070433_, _070434_, _070435_, _070436_, _070437_, _070438_, _070439_, _070440_, _070441_, _070442_, _070443_, _070444_, _070445_, _070446_, _070447_, _070448_, _070449_, _070450_, _070451_, _070452_, _070453_, _070454_, _070455_, _070456_, _070457_, _070458_, _070459_, _070460_, _070461_, _070462_, _070463_, _070464_, _070465_, _070466_, _070467_, _070468_, _070469_, _070470_, _070471_, _070472_, _070473_, _070474_, _070475_, _070476_, _070477_, _070478_, _070479_, _070480_, _070481_, _070482_, _070483_, _070484_, _070485_, _070486_, _070487_, _070488_, _070489_, _070490_, _070491_, _070492_, _070493_, _070494_, _070495_, _070496_, _070497_, _070498_, _070499_, _070500_, _070501_, _070502_, _070503_, _070504_, _070505_, _070506_, _070507_, _070508_, _070509_, _070510_, _070511_, _070512_, _070513_, _070514_, _070515_, _070516_, _070517_, _070518_, _070519_, _070520_, _070521_, _070522_, _070523_, _070524_, _070525_, _070526_, _070527_, _070528_, _070529_, _070530_, _070531_, _070532_, _070533_, _070534_, _070535_, _070536_, _070537_, _070538_, _070539_, _070540_, _070541_, _070542_, _070543_, _070544_, _070545_, _070546_, _070547_, _070548_, _070549_, _070550_, _070551_, _070552_, _070553_, _070554_, _070555_, _070556_, _070557_, _070558_, _070559_, _070560_, _070561_, _070562_, _070563_, _070564_, _070565_, _070566_, _070567_, _070568_, _070569_, _070570_, _070571_, _070572_, _070573_, _070574_, _070575_, _070576_, _070577_, _070578_, _070579_, _070580_, _070581_, _070582_, _070583_, _070584_, _070585_, _070586_, _070587_, _070588_, _070589_, _070590_, _070591_, _070592_, _070593_, _070594_, _070595_, _070596_, _070597_, _070598_, _070599_, _070600_, _070601_, _070602_, _070603_, _070604_, _070605_, _070606_, _070607_, _070608_, _070609_, _070610_, _070611_, _070612_, _070613_, _070614_, _070615_, _070616_, _070617_, _070618_, _070619_, _070620_, _070621_, _070622_, _070623_, _070624_, _070625_, _070626_, _070627_, _070628_, _070629_, _070630_, _070631_, _070632_, _070633_, _070634_, _070635_, _070636_, _070637_, _070638_, _070639_, _070640_, _070641_, _070642_, _070643_, _070644_, _070645_, _070646_, _070647_, _070648_, _070649_, _070650_, _070651_, _070652_, _070653_, _070654_, _070655_, _070656_, _070657_, _070658_, _070659_, _070660_, _070661_, _070662_, _070663_, _070664_, _070665_, _070666_, _070667_, _070668_, _070669_, _070670_, _070671_, _070672_, _070673_, _070674_, _070675_, _070676_, _070677_, _070678_, _070679_, _070680_, _070681_, _070682_, _070683_, _070684_, _070685_, _070686_, _070687_, _070688_, _070689_, _070690_, _070691_, _070692_, _070693_, _070694_, _070695_, _070696_, _070697_, _070698_, _070699_, _070700_, _070701_, _070702_, _070703_, _070704_, _070705_, _070706_, _070707_, _070708_, _070709_, _070710_, _070711_, _070712_, _070713_, _070714_, _070715_, _070716_, _070717_, _070718_, _070719_, _070720_, _070721_, _070722_, _070723_, _070724_, _070725_, _070726_, _070727_, _070728_, _070729_, _070730_, _070731_, _070732_, _070733_, _070734_, _070735_, _070736_, _070737_, _070738_, _070739_, _070740_, _070741_, _070742_, _070743_, _070744_, _070745_, _070746_, _070747_, _070748_, _070749_, _070750_, _070751_, _070752_, _070753_, _070754_, _070755_, _070756_, _070757_, _070758_, _070759_, _070760_, _070761_, _070762_, _070763_, _070764_, _070765_, _070766_, _070767_, _070768_, _070769_, _070770_, _070771_, _070772_, _070773_, _070774_, _070775_, _070776_, _070777_, _070778_, _070779_, _070780_, _070781_, _070782_, _070783_, _070784_, _070785_, _070786_, _070787_, _070788_, _070789_, _070790_, _070791_, _070792_, _070793_, _070794_, _070795_, _070796_, _070797_, _070798_, _070799_, _070800_, _070801_, _070802_, _070803_, _070804_, _070805_, _070806_, _070807_, _070808_, _070809_, _070810_, _070811_, _070812_, _070813_, _070814_, _070815_, _070816_, _070817_, _070818_, _070819_, _070820_, _070821_, _070822_, _070823_, _070824_, _070825_, _070826_, _070827_, _070828_, _070829_, _070830_, _070831_, _070832_, _070833_, _070834_, _070835_, _070836_, _070837_, _070838_, _070839_, _070840_, _070841_, _070842_, _070843_, _070844_, _070845_, _070846_, _070847_, _070848_, _070849_, _070850_, _070851_, _070852_, _070853_, _070854_, _070855_, _070856_, _070857_, _070858_, _070859_, _070860_, _070861_, _070862_, _070863_, _070864_, _070865_, _070866_, _070867_, _070868_, _070869_, _070870_, _070871_, _070872_, _070873_, _070874_, _070875_, _070876_, _070877_, _070878_, _070879_, _070880_, _070881_, _070882_, _070883_, _070884_, _070885_, _070886_, _070887_, _070888_, _070889_, _070890_, _070891_, _070892_, _070893_, _070894_, _070895_, _070896_, _070897_, _070898_, _070899_, _070900_, _070901_, _070902_, _070903_, _070904_, _070905_, _070906_, _070907_, _070908_, _070909_, _070910_, _070911_, _070912_, _070913_, _070914_, _070915_, _070916_, _070917_, _070918_, _070919_, _070920_, _070921_, _070922_, _070923_, _070924_, _070925_, _070926_, _070927_, _070928_, _070929_, _070930_, _070931_, _070932_, _070933_, _070934_, _070935_, _070936_, _070937_, _070938_, _070939_, _070940_, _070941_, _070942_, _070943_, _070944_, _070945_, _070946_, _070947_, _070948_, _070949_, _070950_, _070951_, _070952_, _070953_, _070954_, _070955_, _070956_, _070957_, _070958_, _070959_, _070960_, _070961_, _070962_, _070963_, _070964_, _070965_, _070966_, _070967_, _070968_, _070969_, _070970_, _070971_, _070972_, _070973_, _070974_, _070975_, _070976_, _070977_, _070978_, _070979_, _070980_, _070981_, _070982_, _070983_, _070984_, _070985_, _070986_, _070987_, _070988_, _070989_, _070990_, _070991_, _070992_, _070993_, _070994_, _070995_, _070996_, _070997_, _070998_, _070999_, _071000_, _071001_, _071002_, _071003_, _071004_, _071005_, _071006_, _071007_, _071008_, _071009_, _071010_, _071011_, _071012_, _071013_, _071014_, _071015_, _071016_, _071017_, _071018_, _071019_, _071020_, _071021_, _071022_, _071023_, _071024_, _071025_, _071026_, _071027_, _071028_, _071029_, _071030_, _071031_, _071032_, _071033_, _071034_, _071035_, _071036_, _071037_, _071038_, _071039_, _071040_, _071041_, _071042_, _071043_, _071044_, _071045_, _071046_, _071047_, _071048_, _071049_, _071050_, _071051_, _071052_, _071053_, _071054_, _071055_, _071056_, _071057_, _071058_, _071059_, _071060_, _071061_, _071062_, _071063_, _071064_, _071065_, _071066_, _071067_, _071068_, _071069_, _071070_, _071071_, _071072_, _071073_, _071074_, _071075_, _071076_, _071077_, _071078_, _071079_, _071080_, _071081_, _071082_, _071083_, _071084_, _071085_, _071086_, _071087_, _071088_, _071089_, _071090_, _071091_, _071092_, _071093_, _071094_, _071095_, _071096_, _071097_, _071098_, _071099_, _071100_, _071101_, _071102_, _071103_, _071104_, _071105_, _071106_, _071107_, _071108_, _071109_, _071110_, _071111_, _071112_, _071113_, _071114_, _071115_, _071116_, _071117_, _071118_, _071119_, _071120_, _071121_, _071122_, _071123_, _071124_, _071125_, _071126_, _071127_, _071128_, _071129_, _071130_, _071131_, _071132_, _071133_, _071134_, _071135_, _071136_, _071137_, _071138_, _071139_, _071140_, _071141_, _071142_, _071143_, _071144_, _071145_, _071146_, _071147_, _071148_, _071149_, _071150_, _071151_, _071152_, _071153_, _071154_, _071155_, _071156_, _071157_, _071158_, _071159_, _071160_, _071161_, _071162_, _071163_, _071164_, _071165_, _071166_, _071167_, _071168_, _071169_, _071170_, _071171_, _071172_, _071173_, _071174_, _071175_, _071176_, _071177_, _071178_, _071179_, _071180_, _071181_, _071182_, _071183_, _071184_, _071185_, _071186_, _071187_, _071188_, _071189_, _071190_, _071191_, _071192_, _071193_, _071194_, _071195_, _071196_, _071197_, _071198_, _071199_, _071200_, _071201_, _071202_, _071203_, _071204_, _071205_, _071206_, _071207_, _071208_, _071209_, _071210_, _071211_, _071212_, _071213_, _071214_, _071215_, _071216_, _071217_, _071218_, _071219_, _071220_, _071221_, _071222_, _071223_, _071224_, _071225_, _071226_, _071227_, _071228_, _071229_, _071230_, _071231_, _071232_, _071233_, _071234_, _071235_, _071236_, _071237_, _071238_, _071239_, _071240_, _071241_, _071242_, _071243_, _071244_, _071245_, _071246_, _071247_, _071248_, _071249_, _071250_, _071251_, _071252_, _071253_, _071254_, _071255_, _071256_, _071257_, _071258_, _071259_, _071260_, _071261_, _071262_, _071263_, _071264_, _071265_, _071266_, _071267_, _071268_, _071269_, _071270_, _071271_, _071272_, _071273_, _071274_, _071275_, _071276_, _071277_, _071278_, _071279_, _071280_, _071281_, _071282_, _071283_, _071284_, _071285_, _071286_, _071287_, _071288_, _071289_, _071290_, _071291_, _071292_, _071293_, _071294_, _071295_, _071296_, _071297_, _071298_, _071299_, _071300_, _071301_, _071302_, _071303_, _071304_, _071305_, _071306_, _071307_, _071308_, _071309_, _071310_, _071311_, _071312_, _071313_, _071314_, _071315_, _071316_, _071317_, _071318_, _071319_, _071320_, _071321_, _071322_, _071323_, _071324_, _071325_, _071326_, _071327_, _071328_, _071329_, _071330_, _071331_, _071332_, _071333_, _071334_, _071335_, _071336_, _071337_, _071338_, _071339_, _071340_, _071341_, _071342_, _071343_, _071344_, _071345_, _071346_, _071347_, _071348_, _071349_, _071350_, _071351_, _071352_, _071353_, _071354_, _071355_, _071356_, _071357_, _071358_, _071359_, _071360_, _071361_, _071362_, _071363_, _071364_, _071365_, _071366_, _071367_, _071368_, _071369_, _071370_, _071371_, _071372_, _071373_, _071374_, _071375_, _071376_, _071377_, _071378_, _071379_, _071380_, _071381_, _071382_, _071383_, _071384_, _071385_, _071386_, _071387_, _071388_, _071389_, _071390_, _071391_, _071392_, _071393_, _071394_, _071395_, _071396_, _071397_, _071398_, _071399_, _071400_, _071401_, _071402_, _071403_, _071404_, _071405_, _071406_, _071407_, _071408_, _071409_, _071410_, _071411_, _071412_, _071413_, _071414_, _071415_, _071416_, _071417_, _071418_, _071419_, _071420_, _071421_, _071422_, _071423_, _071424_, _071425_, _071426_, _071427_, _071428_, _071429_, _071430_, _071431_, _071432_, _071433_, _071434_, _071435_, _071436_, _071437_, _071438_, _071439_, _071440_, _071441_, _071442_, _071443_, _071444_, _071445_, _071446_, _071447_, _071448_, _071449_, _071450_, _071451_, _071452_, _071453_, _071454_, _071455_, _071456_, _071457_, _071458_, _071459_, _071460_, _071461_, _071462_, _071463_, _071464_, _071465_, _071466_, _071467_, _071468_, _071469_, _071470_, _071471_, _071472_, _071473_, _071474_, _071475_, _071476_, _071477_, _071478_, _071479_, _071480_, _071481_, _071482_, _071483_, _071484_, _071485_, _071486_, _071487_, _071488_, _071489_, _071490_, _071491_, _071492_, _071493_, _071494_, _071495_, _071496_, _071497_, _071498_, _071499_, _071500_, _071501_, _071502_, _071503_, _071504_, _071505_, _071506_, _071507_, _071508_, _071509_, _071510_, _071511_, _071512_, _071513_, _071514_, _071515_, _071516_, _071517_, _071518_, _071519_, _071520_, _071521_, _071522_, _071523_, _071524_, _071525_, _071526_, _071527_, _071528_, _071529_, _071530_, _071531_, _071532_, _071533_, _071534_, _071535_, _071536_, _071537_, _071538_, _071539_, _071540_, _071541_, _071542_, _071543_, _071544_, _071545_, _071546_, _071547_, _071548_, _071549_, _071550_, _071551_, _071552_, _071553_, _071554_, _071555_, _071556_, _071557_, _071558_, _071559_, _071560_, _071561_, _071562_, _071563_, _071564_, _071565_, _071566_, _071567_, _071568_, _071569_, _071570_, _071571_, _071572_, _071573_, _071574_, _071575_, _071576_, _071577_, _071578_, _071579_, _071580_, _071581_, _071582_, _071583_, _071584_, _071585_, _071586_, _071587_, _071588_, _071589_, _071590_, _071591_, _071592_, _071593_, _071594_, _071595_, _071596_, _071597_, _071598_, _071599_, _071600_, _071601_, _071602_, _071603_, _071604_, _071605_, _071606_, _071607_, _071608_, _071609_, _071610_, _071611_, _071612_, _071613_, _071614_, _071615_, _071616_, _071617_, _071618_, _071619_, _071620_, _071621_, _071622_, _071623_, _071624_, _071625_, _071626_, _071627_, _071628_, _071629_, _071630_, _071631_, _071632_, _071633_, _071634_, _071635_, _071636_, _071637_, _071638_, _071639_, _071640_, _071641_, _071642_, _071643_, _071644_, _071645_, _071646_, _071647_, _071648_, _071649_, _071650_, _071651_, _071652_, _071653_, _071654_, _071655_, _071656_, _071657_, _071658_, _071659_, _071660_, _071661_, _071662_, _071663_, _071664_, _071665_, _071666_, _071667_, _071668_, _071669_, _071670_, _071671_, _071672_, _071673_, _071674_, _071675_, _071676_, _071677_, _071678_, _071679_, _071680_, _071681_, _071682_, _071683_, _071684_, _071685_, _071686_, _071687_, _071688_, _071689_, _071690_, _071691_, _071692_, _071693_, _071694_, _071695_, _071696_, _071697_, _071698_, _071699_, _071700_, _071701_, _071702_, _071703_, _071704_, _071705_, _071706_, _071707_, _071708_, _071709_, _071710_, _071711_, _071712_, _071713_, _071714_, _071715_, _071716_, _071717_, _071718_, _071719_, _071720_, _071721_, _071722_, _071723_, _071724_, _071725_, _071726_, _071727_, _071728_, _071729_, _071730_, _071731_, _071732_, _071733_, _071734_, _071735_, _071736_, _071737_, _071738_, _071739_, _071740_, _071741_, _071742_, _071743_, _071744_, _071745_, _071746_, _071747_, _071748_, _071749_, _071750_, _071751_, _071752_, _071753_, _071754_, _071755_, _071756_, _071757_, _071758_, _071759_, _071760_, _071761_, _071762_, _071763_, _071764_, _071765_, _071766_, _071767_, _071768_, _071769_, _071770_, _071771_, _071772_, _071773_, _071774_, _071775_, _071776_, _071777_, _071778_, _071779_, _071780_, _071781_, _071782_, _071783_, _071784_, _071785_, _071786_, _071787_, _071788_, _071789_, _071790_, _071791_, _071792_, _071793_, _071794_, _071795_, _071796_, _071797_, _071798_, _071799_, _071800_, _071801_, _071802_, _071803_, _071804_, _071805_, _071806_, _071807_, _071808_, _071809_, _071810_, _071811_, _071812_, _071813_, _071814_, _071815_, _071816_, _071817_, _071818_, _071819_, _071820_, _071821_, _071822_, _071823_, _071824_, _071825_, _071826_, _071827_, _071828_, _071829_, _071830_, _071831_, _071832_, _071833_, _071834_, _071835_, _071836_, _071837_, _071838_, _071839_, _071840_, _071841_, _071842_, _071843_, _071844_, _071845_, _071846_, _071847_, _071848_, _071849_, _071850_, _071851_, _071852_, _071853_, _071854_, _071855_, _071856_, _071857_, _071858_, _071859_, _071860_, _071861_, _071862_, _071863_, _071864_, _071865_, _071866_, _071867_, _071868_, _071869_, _071870_, _071871_, _071872_, _071873_, _071874_, _071875_, _071876_, _071877_, _071878_, _071879_, _071880_, _071881_, _071882_, _071883_, _071884_, _071885_, _071886_, _071887_, _071888_, _071889_, _071890_, _071891_, _071892_, _071893_, _071894_, _071895_, _071896_, _071897_, _071898_, _071899_, _071900_, _071901_, _071902_, _071903_, _071904_, _071905_, _071906_, _071907_, _071908_, _071909_, _071910_, _071911_, _071912_, _071913_, _071914_, _071915_, _071916_, _071917_, _071918_, _071919_, _071920_, _071921_, _071922_, _071923_, _071924_, _071925_, _071926_, _071927_, _071928_, _071929_, _071930_, _071931_, _071932_, _071933_, _071934_, _071935_, _071936_, _071937_, _071938_, _071939_, _071940_, _071941_, _071942_, _071943_, _071944_, _071945_, _071946_, _071947_, _071948_, _071949_, _071950_, _071951_, _071952_, _071953_, _071954_, _071955_, _071956_, _071957_, _071958_, _071959_, _071960_, _071961_, _071962_, _071963_, _071964_, _071965_, _071966_, _071967_, _071968_, _071969_, _071970_, _071971_, _071972_, _071973_, _071974_, _071975_, _071976_, _071977_, _071978_, _071979_, _071980_, _071981_, _071982_, _071983_, _071984_, _071985_, _071986_, _071987_, _071988_, _071989_, _071990_, _071991_, _071992_, _071993_, _071994_, _071995_, _071996_, _071997_, _071998_, _071999_, _072000_, _072001_, _072002_, _072003_, _072004_, _072005_, _072006_, _072007_, _072008_, _072009_, _072010_, _072011_, _072012_, _072013_, _072014_, _072015_, _072016_, _072017_, _072018_, _072019_, _072020_, _072021_, _072022_, _072023_, _072024_, _072025_, _072026_, _072027_, _072028_, _072029_, _072030_, _072031_, _072032_, _072033_, _072034_, _072035_, _072036_, _072037_, _072038_, _072039_, _072040_, _072041_, _072042_, _072043_, _072044_, _072045_, _072046_, _072047_, _072048_, _072049_, _072050_, _072051_, _072052_, _072053_, _072054_, _072055_, _072056_, _072057_, _072058_, _072059_, _072060_, _072061_, _072062_, _072063_, _072064_, _072065_, _072066_, _072067_, _072068_, _072069_, _072070_, _072071_, _072072_, _072073_, _072074_, _072075_, _072076_, _072077_, _072078_, _072079_, _072080_, _072081_, _072082_, _072083_, _072084_, _072085_, _072086_, _072087_, _072088_, _072089_, _072090_, _072091_, _072092_, _072093_, _072094_, _072095_, _072096_, _072097_, _072098_, _072099_, _072100_, _072101_, _072102_, _072103_, _072104_, _072105_, _072106_, _072107_, _072108_, _072109_, _072110_, _072111_, _072112_, _072113_, _072114_, _072115_, _072116_, _072117_, _072118_, _072119_, _072120_, _072121_, _072122_, _072123_, _072124_, _072125_, _072126_, _072127_, _072128_, _072129_, _072130_, _072131_, _072132_, _072133_, _072134_, _072135_, _072136_, _072137_, _072138_, _072139_, _072140_, _072141_, _072142_, _072143_, _072144_, _072145_, _072146_, _072147_, _072148_, _072149_, _072150_, _072151_, _072152_, _072153_, _072154_, _072155_, _072156_, _072157_, _072158_, _072159_, _072160_, _072161_, _072162_, _072163_, _072164_, _072165_, _072166_, _072167_, _072168_, _072169_, _072170_, _072171_, _072172_, _072173_, _072174_, _072175_, _072176_, _072177_, _072178_, _072179_, _072180_, _072181_, _072182_, _072183_, _072184_, _072185_, _072186_, _072187_, _072188_, _072189_, _072190_, _072191_, _072192_, _072193_, _072194_, _072195_, _072196_, _072197_, _072198_, _072199_, _072200_, _072201_, _072202_, _072203_, _072204_, _072205_, _072206_, _072207_, _072208_, _072209_, _072210_, _072211_, _072212_, _072213_, _072214_, _072215_, _072216_, _072217_, _072218_, _072219_, _072220_, _072221_, _072222_, _072223_, _072224_, _072225_, _072226_, _072227_, _072228_, _072229_, _072230_, _072231_, _072232_, _072233_, _072234_, _072235_, _072236_, _072237_, _072238_, _072239_, _072240_, _072241_, _072242_, _072243_, _072244_, _072245_, _072246_, _072247_, _072248_, _072249_, _072250_, _072251_, _072252_, _072253_, _072254_, _072255_, _072256_, _072257_, _072258_, _072259_, _072260_, _072261_, _072262_, _072263_, _072264_, _072265_, _072266_, _072267_, _072268_, _072269_, _072270_, _072271_, _072272_, _072273_, _072274_, _072275_, _072276_, _072277_, _072278_, _072279_, _072280_, _072281_, _072282_, _072283_, _072284_, _072285_, _072286_, _072287_, _072288_, _072289_, _072290_, _072291_, _072292_, _072293_, _072294_, _072295_, _072296_, _072297_, _072298_, _072299_, _072300_, _072301_, _072302_, _072303_, _072304_, _072305_, _072306_, _072307_, _072308_, _072309_, _072310_, _072311_, _072312_, _072313_, _072314_, _072315_, _072316_, _072317_, _072318_, _072319_, _072320_, _072321_, _072322_, _072323_, _072324_, _072325_, _072326_, _072327_, _072328_, _072329_, _072330_, _072331_, _072332_, _072333_, _072334_, _072335_, _072336_, _072337_, _072338_, _072339_, _072340_, _072341_, _072342_, _072343_, _072344_, _072345_, _072346_, _072347_, _072348_, _072349_, _072350_, _072351_, _072352_, _072353_, _072354_, _072355_, _072356_, _072357_, _072358_, _072359_, _072360_, _072361_, _072362_, _072363_, _072364_, _072365_, _072366_, _072367_, _072368_, _072369_, _072370_, _072371_, _072372_, _072373_, _072374_, _072375_, _072376_, _072377_, _072378_, _072379_, _072380_, _072381_, _072382_, _072383_, _072384_, _072385_, _072386_, _072387_, _072388_, _072389_, _072390_, _072391_, _072392_, _072393_, _072394_, _072395_, _072396_, _072397_, _072398_, _072399_, _072400_, _072401_, _072402_, _072403_, _072404_, _072405_, _072406_, _072407_, _072408_, _072409_, _072410_, _072411_, _072412_, _072413_, _072414_, _072415_, _072416_, _072417_, _072418_, _072419_, _072420_, _072421_, _072422_, _072423_, _072424_, _072425_, _072426_, _072427_, _072428_, _072429_, _072430_, _072431_, _072432_, _072433_, _072434_, _072435_, _072436_, _072437_, _072438_, _072439_, _072440_, _072441_, _072442_, _072443_, _072444_, _072445_, _072446_, _072447_, _072448_, _072449_, _072450_, _072451_, _072452_, _072453_, _072454_, _072455_, _072456_, _072457_, _072458_, _072459_, _072460_, _072461_, _072462_, _072463_, _072464_, _072465_, _072466_, _072467_, _072468_, _072469_, _072470_, _072471_, _072472_, _072473_, _072474_, _072475_, _072476_, _072477_, _072478_, _072479_, _072480_, _072481_, _072482_, _072483_, _072484_, _072485_, _072486_, _072487_, _072488_, _072489_, _072490_, _072491_, _072492_, _072493_, _072494_, _072495_, _072496_, _072497_, _072498_, _072499_, _072500_, _072501_, _072502_, _072503_, _072504_, _072505_, _072506_, _072507_, _072508_, _072509_, _072510_, _072511_, _072512_, _072513_, _072514_, _072515_, _072516_, _072517_, _072518_, _072519_, _072520_, _072521_, _072522_, _072523_, _072524_, _072525_, _072526_, _072527_, _072528_, _072529_, _072530_, _072531_, _072532_, _072533_, _072534_, _072535_, _072536_, _072537_, _072538_, _072539_, _072540_, _072541_, _072542_, _072543_, _072544_, _072545_, _072546_, _072547_, _072548_, _072549_, _072550_, _072551_, _072552_, _072553_, _072554_, _072555_, _072556_, _072557_, _072558_, _072559_, _072560_, _072561_, _072562_, _072563_, _072564_, _072565_, _072566_, _072567_, _072568_, _072569_, _072570_, _072571_, _072572_, _072573_, _072574_, _072575_, _072576_, _072577_, _072578_, _072579_, _072580_, _072581_, _072582_, _072583_, _072584_, _072585_, _072586_, _072587_, _072588_, _072589_, _072590_, _072591_, _072592_, _072593_, _072594_, _072595_, _072596_, _072597_, _072598_, _072599_, _072600_, _072601_, _072602_, _072603_, _072604_, _072605_, _072606_, _072607_, _072608_, _072609_, _072610_, _072611_, _072612_, _072613_, _072614_, _072615_, _072616_, _072617_, _072618_, _072619_, _072620_, _072621_, _072622_, _072623_, _072624_, _072625_, _072626_, _072627_, _072628_, _072629_, _072630_, _072631_, _072632_, _072633_, _072634_, _072635_, _072636_, _072637_, _072638_, _072639_, _072640_, _072641_, _072642_, _072643_, _072644_, _072645_, _072646_, _072647_, _072648_, _072649_, _072650_, _072651_, _072652_, _072653_, _072654_, _072655_, _072656_, _072657_, _072658_, _072659_, _072660_, _072661_, _072662_, _072663_, _072664_, _072665_, _072666_, _072667_, _072668_, _072669_, _072670_, _072671_, _072672_, _072673_, _072674_, _072675_, _072676_, _072677_, _072678_, _072679_, _072680_, _072681_, _072682_, _072683_, _072684_, _072685_, _072686_, _072687_, _072688_, _072689_, _072690_, _072691_, _072692_, _072693_, _072694_, _072695_, _072696_, _072697_, _072698_, _072699_, _072700_, _072701_, _072702_, _072703_, _072704_, _072705_, _072706_, _072707_, _072708_, _072709_, _072710_, _072711_, _072712_, _072713_, _072714_, _072715_, _072716_, _072717_, _072718_, _072719_, _072720_, _072721_, _072722_, _072723_, _072724_, _072725_, _072726_, _072727_, _072728_, _072729_, _072730_, _072731_, _072732_, _072733_, _072734_, _072735_, _072736_, _072737_, _072738_, _072739_, _072740_, _072741_, _072742_, _072743_, _072744_, _072745_, _072746_, _072747_, _072748_, _072749_, _072750_, _072751_, _072752_, _072753_, _072754_, _072755_, _072756_, _072757_, _072758_, _072759_, _072760_, _072761_, _072762_, _072763_, _072764_, _072765_, _072766_, _072767_, _072768_, _072769_, _072770_, _072771_, _072772_, _072773_, _072774_, _072775_, _072776_, _072777_, _072778_, _072779_, _072780_, _072781_, _072782_, _072783_, _072784_, _072785_, _072786_, _072787_, _072788_, _072789_, _072790_, _072791_, _072792_, _072793_, _072794_, _072795_, _072796_, _072797_, _072798_, _072799_, _072800_, _072801_, _072802_, _072803_, _072804_, _072805_, _072806_, _072807_, _072808_, _072809_, _072810_, _072811_, _072812_, _072813_, _072814_, _072815_, _072816_, _072817_, _072818_, _072819_, _072820_, _072821_, _072822_, _072823_, _072824_, _072825_, _072826_, _072827_, _072828_, _072829_, _072830_, _072831_, _072832_, _072833_, _072834_, _072835_, _072836_, _072837_, _072838_, _072839_, _072840_, _072841_, _072842_, _072843_, _072844_, _072845_, _072846_, _072847_, _072848_, _072849_, _072850_, _072851_, _072852_, _072853_, _072854_, _072855_, _072856_, _072857_, _072858_, _072859_, _072860_, _072861_, _072862_, _072863_, _072864_, _072865_, _072866_, _072867_, _072868_, _072869_, _072870_, _072871_, _072872_, _072873_, _072874_, _072875_, _072876_, _072877_, _072878_, _072879_, _072880_, _072881_, _072882_, _072883_, _072884_, _072885_, _072886_, _072887_, _072888_, _072889_, _072890_, _072891_, _072892_, _072893_, _072894_, _072895_, _072896_, _072897_, _072898_, _072899_, _072900_, _072901_, _072902_, _072903_, _072904_, _072905_, _072906_, _072907_, _072908_, _072909_, _072910_, _072911_, _072912_, _072913_, _072914_, _072915_, _072916_, _072917_, _072918_, _072919_, _072920_, _072921_, _072922_, _072923_, _072924_, _072925_, _072926_, _072927_, _072928_, _072929_, _072930_, _072931_, _072932_, _072933_, _072934_, _072935_, _072936_, _072937_, _072938_, _072939_, _072940_, _072941_, _072942_, _072943_, _072944_, _072945_, _072946_, _072947_, _072948_, _072949_, _072950_, _072951_, _072952_, _072953_, _072954_, _072955_, _072956_, _072957_, _072958_, _072959_, _072960_, _072961_, _072962_, _072963_, _072964_, _072965_, _072966_, _072967_, _072968_, _072969_, _072970_, _072971_, _072972_, _072973_, _072974_, _072975_, _072976_, _072977_, _072978_, _072979_, _072980_, _072981_, _072982_, _072983_, _072984_, _072985_, _072986_, _072987_, _072988_, _072989_, _072990_, _072991_, _072992_, _072993_, _072994_, _072995_, _072996_, _072997_, _072998_, _072999_, _073000_, _073001_, _073002_, _073003_, _073004_, _073005_, _073006_, _073007_, _073008_, _073009_, _073010_, _073011_, _073012_, _073013_, _073014_, _073015_, _073016_, _073017_, _073018_, _073019_, _073020_, _073021_, _073022_, _073023_, _073024_, _073025_, _073026_, _073027_, _073028_, _073029_, _073030_, _073031_, _073032_, _073033_, _073034_, _073035_, _073036_, _073037_, _073038_, _073039_, _073040_, _073041_, _073042_, _073043_, _073044_, _073045_, _073046_, _073047_, _073048_, _073049_, _073050_, _073051_, _073052_, _073053_, _073054_, _073055_, _073056_, _073057_, _073058_, _073059_, _073060_, _073061_, _073062_, _073063_, _073064_, _073065_, _073066_, _073067_, _073068_, _073069_, _073070_, _073071_, _073072_, _073073_, _073074_, _073075_, _073076_, _073077_, _073078_, _073079_, _073080_, _073081_, _073082_, _073083_, _073084_, _073085_, _073086_, _073087_, _073088_, _073089_, _073090_, _073091_, _073092_, _073093_, _073094_, _073095_, _073096_, _073097_, _073098_, _073099_, _073100_, _073101_, _073102_, _073103_, _073104_, _073105_, _073106_, _073107_, _073108_, _073109_, _073110_, _073111_, _073112_, _073113_, _073114_, _073115_, _073116_, _073117_, _073118_, _073119_, _073120_, _073121_, _073122_, _073123_, _073124_, _073125_, _073126_, _073127_, _073128_, _073129_, _073130_, _073131_, _073132_, _073133_, _073134_, _073135_, _073136_, _073137_, _073138_, _073139_, _073140_, _073141_, _073142_, _073143_, _073144_, _073145_, _073146_, _073147_, _073148_, _073149_, _073150_, _073151_, _073152_, _073153_, _073154_, _073155_, _073156_, _073157_, _073158_, _073159_, _073160_, _073161_, _073162_, _073163_, _073164_, _073165_, _073166_, _073167_, _073168_, _073169_, _073170_, _073171_, _073172_, _073173_, _073174_, _073175_, _073176_, _073177_, _073178_, _073179_, _073180_, _073181_, _073182_, _073183_, _073184_, _073185_, _073186_, _073187_, _073188_, _073189_, _073190_, _073191_, _073192_, _073193_, _073194_, _073195_, _073196_, _073197_, _073198_, _073199_, _073200_, _073201_, _073202_, _073203_, _073204_, _073205_, _073206_, _073207_, _073208_, _073209_, _073210_, _073211_, _073212_, _073213_, _073214_, _073215_, _073216_, _073217_, _073218_, _073219_, _073220_, _073221_, _073222_, _073223_, _073224_, _073225_, _073226_, _073227_, _073228_, _073229_, _073230_, _073231_, _073232_, _073233_, _073234_, _073235_, _073236_, _073237_, _073238_, _073239_, _073240_, _073241_, _073242_, _073243_, _073244_, _073245_, _073246_, _073247_, _073248_, _073249_, _073250_, _073251_, _073252_, _073253_, _073254_, _073255_, _073256_, _073257_, _073258_, _073259_, _073260_, _073261_, _073262_, _073263_, _073264_, _073265_, _073266_, _073267_, _073268_, _073269_, _073270_, _073271_, _073272_, _073273_, _073274_, _073275_, _073276_, _073277_, _073278_, _073279_, _073280_, _073281_, _073282_, _073283_, _073284_, _073285_, _073286_, _073287_, _073288_, _073289_, _073290_, _073291_, _073292_, _073293_, _073294_, _073295_, _073296_, _073297_, _073298_, _073299_, _073300_, _073301_, _073302_, _073303_, _073304_, _073305_, _073306_, _073307_, _073308_, _073309_, _073310_, _073311_, _073312_, _073313_, _073314_, _073315_, _073316_, _073317_, _073318_, _073319_, _073320_, _073321_, _073322_, _073323_, _073324_, _073325_, _073326_, _073327_, _073328_, _073329_, _073330_, _073331_, _073332_, _073333_, _073334_, _073335_, _073336_, _073337_, _073338_, _073339_, _073340_, _073341_, _073342_, _073343_, _073344_, _073345_, _073346_, _073347_, _073348_, _073349_, _073350_, _073351_, _073352_, _073353_, _073354_, _073355_, _073356_, _073357_, _073358_, _073359_, _073360_, _073361_, _073362_, _073363_, _073364_, _073365_, _073366_, _073367_, _073368_, _073369_, _073370_, _073371_, _073372_, _073373_, _073374_, _073375_, _073376_, _073377_, _073378_, _073379_, _073380_, _073381_, _073382_, _073383_, _073384_, _073385_, _073386_, _073387_, _073388_, _073389_, _073390_, _073391_, _073392_, _073393_, _073394_, _073395_, _073396_, _073397_, _073398_, _073399_, _073400_, _073401_, _073402_, _073403_, _073404_, _073405_, _073406_, _073407_, _073408_, _073409_, _073410_, _073411_, _073412_, _073413_, _073414_, _073415_, _073416_, _073417_, _073418_, _073419_, _073420_, _073421_, _073422_, _073423_, _073424_, _073425_, _073426_, _073427_, _073428_, _073429_, _073430_, _073431_, _073432_, _073433_, _073434_, _073435_, _073436_, _073437_, _073438_, _073439_, _073440_, _073441_, _073442_, _073443_, _073444_, _073445_, _073446_, _073447_, _073448_, _073449_, _073450_, _073451_, _073452_, _073453_, _073454_, _073455_, _073456_, _073457_, _073458_, _073459_, _073460_, _073461_, _073462_, _073463_, _073464_, _073465_, _073466_, _073467_, _073468_, _073469_, _073470_, _073471_, _073472_, _073473_, _073474_, _073475_, _073476_, _073477_, _073478_, _073479_, _073480_, _073481_, _073482_, _073483_, _073484_, _073485_, _073486_, _073487_, _073488_, _073489_, _073490_, _073491_, _073492_, _073493_, _073494_, _073495_, _073496_, _073497_, _073498_, _073499_, _073500_, _073501_, _073502_, _073503_, _073504_, _073505_, _073506_, _073507_, _073508_, _073509_, _073510_, _073511_, _073512_, _073513_, _073514_, _073515_, _073516_, _073517_, _073518_, _073519_, _073520_, _073521_, _073522_, _073523_, _073524_, _073525_, _073526_, _073527_, _073528_, _073529_, _073530_, _073531_, _073532_, _073533_, _073534_, _073535_, _073536_, _073537_, _073538_, _073539_, _073540_, _073541_, _073542_, _073543_, _073544_, _073545_, _073546_, _073547_, _073548_, _073549_, _073550_, _073551_, _073552_, _073553_, _073554_, _073555_, _073556_, _073557_, _073558_, _073559_, _073560_, _073561_, _073562_, _073563_, _073564_, _073565_, _073566_, _073567_, _073568_, _073569_, _073570_, _073571_, _073572_, _073573_, _073574_, _073575_, _073576_, _073577_, _073578_, _073579_, _073580_, _073581_, _073582_, _073583_, _073584_, _073585_, _073586_, _073587_, _073588_, _073589_, _073590_, _073591_, _073592_, _073593_, _073594_, _073595_, _073596_, _073597_, _073598_, _073599_, _073600_, _073601_, _073602_, _073603_, _073604_, _073605_, _073606_, _073607_, _073608_, _073609_, _073610_, _073611_, _073612_, _073613_, _073614_, _073615_, _073616_, _073617_, _073618_, _073619_, _073620_, _073621_, _073622_, _073623_, _073624_, _073625_, _073626_, _073627_, _073628_, _073629_, _073630_, _073631_, _073632_, _073633_, _073634_, _073635_, _073636_, _073637_, _073638_, _073639_, _073640_, _073641_, _073642_, _073643_, _073644_, _073645_, _073646_, _073647_, _073648_, _073649_, _073650_, _073651_, _073652_, _073653_, _073654_, _073655_, _073656_, _073657_, _073658_, _073659_, _073660_, _073661_, _073662_, _073663_, _073664_, _073665_, _073666_, _073667_, _073668_, _073669_, _073670_, _073671_, _073672_, _073673_, _073674_, _073675_, _073676_, _073677_, _073678_, _073679_, _073680_, _073681_, _073682_, _073683_, _073684_, _073685_, _073686_, _073687_, _073688_, _073689_, _073690_, _073691_, _073692_, _073693_, _073694_, _073695_, _073696_, _073697_, _073698_, _073699_, _073700_, _073701_, _073702_, _073703_, _073704_, _073705_, _073706_, _073707_, _073708_, _073709_, _073710_, _073711_, _073712_, _073713_, _073714_, _073715_, _073716_, _073717_, _073718_, _073719_, _073720_, _073721_, _073722_, _073723_, _073724_, _073725_, _073726_, _073727_, _073728_, _073729_, _073730_, _073731_, _073732_, _073733_, _073734_, _073735_, _073736_, _073737_, _073738_, _073739_, _073740_, _073741_, _073742_, _073743_, _073744_, _073745_, _073746_, _073747_, _073748_, _073749_, _073750_, _073751_, _073752_, _073753_, _073754_, _073755_, _073756_, _073757_, _073758_, _073759_, _073760_, _073761_, _073762_, _073763_, _073764_, _073765_, _073766_, _073767_, _073768_, _073769_, _073770_, _073771_, _073772_, _073773_, _073774_, _073775_, _073776_, _073777_, _073778_, _073779_, _073780_, _073781_, _073782_, _073783_, _073784_, _073785_, _073786_, _073787_, _073788_, _073789_, _073790_, _073791_, _073792_, _073793_, _073794_, _073795_, _073796_, _073797_, _073798_, _073799_, _073800_, _073801_, _073802_, _073803_, _073804_, _073805_, _073806_, _073807_, _073808_, _073809_, _073810_, _073811_, _073812_, _073813_, _073814_, _073815_, _073816_, _073817_, _073818_, _073819_, _073820_, _073821_, _073822_, _073823_, _073824_, _073825_, _073826_, _073827_, _073828_, _073829_, _073830_, _073831_, _073832_, _073833_, _073834_, _073835_, _073836_, _073837_, _073838_, _073839_, _073840_, _073841_, _073842_, _073843_, _073844_, _073845_, _073846_, _073847_, _073848_, _073849_, _073850_, _073851_, _073852_, _073853_, _073854_, _073855_, _073856_, _073857_, _073858_, _073859_, _073860_, _073861_, _073862_, _073863_, _073864_, _073865_, _073866_, _073867_, _073868_, _073869_, _073870_, _073871_, _073872_, _073873_, _073874_, _073875_, _073876_, _073877_, _073878_, _073879_, _073880_, _073881_, _073882_, _073883_, _073884_, _073885_, _073886_, _073887_, _073888_, _073889_, _073890_, _073891_, _073892_, _073893_, _073894_, _073895_, _073896_, _073897_, _073898_, _073899_, _073900_, _073901_, _073902_, _073903_, _073904_, _073905_, _073906_, _073907_, _073908_, _073909_, _073910_, _073911_, _073912_, _073913_, _073914_, _073915_, _073916_, _073917_, _073918_, _073919_, _073920_, _073921_, _073922_, _073923_, _073924_, _073925_, _073926_, _073927_, _073928_, _073929_, _073930_, _073931_, _073932_, _073933_, _073934_, _073935_, _073936_, _073937_, _073938_, _073939_, _073940_, _073941_, _073942_, _073943_, _073944_, _073945_, _073946_, _073947_, _073948_, _073949_, _073950_, _073951_, _073952_, _073953_, _073954_, _073955_, _073956_, _073957_, _073958_, _073959_, _073960_, _073961_, _073962_, _073963_, _073964_, _073965_, _073966_, _073967_, _073968_, _073969_, _073970_, _073971_, _073972_, _073973_, _073974_, _073975_, _073976_, _073977_, _073978_, _073979_, _073980_, _073981_, _073982_, _073983_, _073984_, _073985_, _073986_, _073987_, _073988_, _073989_, _073990_, _073991_, _073992_, _073993_, _073994_, _073995_, _073996_, _073997_, _073998_, _073999_, _074000_, _074001_, _074002_, _074003_, _074004_, _074005_, _074006_, _074007_, _074008_, _074009_, _074010_, _074011_, _074012_, _074013_, _074014_, _074015_, _074016_, _074017_, _074018_, _074019_, _074020_, _074021_, _074022_, _074023_, _074024_, _074025_, _074026_, _074027_, _074028_, _074029_, _074030_, _074031_, _074032_, _074033_, _074034_, _074035_, _074036_, _074037_, _074038_, _074039_, _074040_, _074041_, _074042_, _074043_, _074044_, _074045_, _074046_, _074047_, _074048_, _074049_, _074050_, _074051_, _074052_, _074053_, _074054_, _074055_, _074056_, _074057_, _074058_, _074059_, _074060_, _074061_, _074062_, _074063_, _074064_, _074065_, _074066_, _074067_, _074068_, _074069_, _074070_, _074071_, _074072_, _074073_, _074074_, _074075_, _074076_, _074077_, _074078_, _074079_, _074080_, _074081_, _074082_, _074083_, _074084_, _074085_, _074086_, _074087_, _074088_, _074089_, _074090_, _074091_, _074092_, _074093_, _074094_, _074095_, _074096_, _074097_, _074098_, _074099_, _074100_, _074101_, _074102_, _074103_, _074104_, _074105_, _074106_, _074107_, _074108_, _074109_, _074110_, _074111_, _074112_, _074113_, _074114_, _074115_, _074116_, _074117_, _074118_, _074119_, _074120_, _074121_, _074122_, _074123_, _074124_, _074125_, _074126_, _074127_, _074128_, _074129_, _074130_, _074131_, _074132_, _074133_, _074134_, _074135_, _074136_, _074137_, _074138_, _074139_, _074140_, _074141_, _074142_, _074143_, _074144_, _074145_, _074146_, _074147_, _074148_, _074149_, _074150_, _074151_, _074152_, _074153_, _074154_, _074155_, _074156_, _074157_, _074158_, _074159_, _074160_, _074161_, _074162_, _074163_, _074164_, _074165_, _074166_, _074167_, _074168_, _074169_, _074170_, _074171_, _074172_, _074173_, _074174_, _074175_, _074176_, _074177_, _074178_, _074179_, _074180_, _074181_, _074182_, _074183_, _074184_, _074185_, _074186_, _074187_, _074188_, _074189_, _074190_, _074191_, _074192_, _074193_, _074194_, _074195_, _074196_, _074197_, _074198_, _074199_, _074200_, _074201_, _074202_, _074203_, _074204_, _074205_, _074206_, _074207_, _074208_, _074209_, _074210_, _074211_, _074212_, _074213_, _074214_, _074215_, _074216_, _074217_, _074218_, _074219_, _074220_, _074221_, _074222_, _074223_, _074224_, _074225_, _074226_, _074227_, _074228_, _074229_, _074230_, _074231_, _074232_, _074233_, _074234_, _074235_, _074236_, _074237_, _074238_, _074239_, _074240_, _074241_, _074242_, _074243_, _074244_, _074245_, _074246_, _074247_, _074248_, _074249_, _074250_, _074251_, _074252_, _074253_, _074254_, _074255_, _074256_, _074257_, _074258_, _074259_, _074260_, _074261_, _074262_, _074263_, _074264_, _074265_, _074266_, _074267_, _074268_, _074269_, _074270_, _074271_, _074272_, _074273_, _074274_, _074275_, _074276_, _074277_, _074278_, _074279_, _074280_, _074281_, _074282_, _074283_, _074284_, _074285_, _074286_, _074287_, _074288_, _074289_, _074290_, _074291_, _074292_, _074293_, _074294_, _074295_, _074296_, _074297_, _074298_, _074299_, _074300_, _074301_, _074302_, _074303_, _074304_, _074305_, _074306_, _074307_, _074308_, _074309_, _074310_, _074311_, _074312_, _074313_, _074314_, _074315_, _074316_, _074317_, _074318_, _074319_, _074320_, _074321_, _074322_, _074323_, _074324_, _074325_, _074326_, _074327_, _074328_, _074329_, _074330_, _074331_, _074332_, _074333_, _074334_, _074335_, _074336_, _074337_, _074338_, _074339_, _074340_, _074341_, _074342_, _074343_, _074344_, _074345_, _074346_, _074347_, _074348_, _074349_, _074350_, _074351_, _074352_, _074353_, _074354_, _074355_, _074356_, _074357_, _074358_, _074359_, _074360_, _074361_, _074362_, _074363_, _074364_, _074365_, _074366_, _074367_, _074368_, _074369_, _074370_, _074371_, _074372_, _074373_, _074374_, _074375_, _074376_, _074377_, _074378_, _074379_, _074380_, _074381_, _074382_, _074383_, _074384_, _074385_, _074386_, _074387_, _074388_, _074389_, _074390_, _074391_, _074392_, _074393_, _074394_, _074395_, _074396_, _074397_, _074398_, _074399_, _074400_, _074401_, _074402_, _074403_, _074404_, _074405_, _074406_, _074407_, _074408_, _074409_, _074410_, _074411_, _074412_, _074413_, _074414_, _074415_, _074416_, _074417_, _074418_, _074419_, _074420_, _074421_, _074422_, _074423_, _074424_, _074425_, _074426_, _074427_, _074428_, _074429_, _074430_, _074431_, _074432_, _074433_, _074434_, _074435_, _074436_, _074437_, _074438_, _074439_, _074440_, _074441_, _074442_, _074443_, _074444_, _074445_, _074446_, _074447_, _074448_, _074449_, _074450_, _074451_, _074452_, _074453_, _074454_, _074455_, _074456_, _074457_, _074458_, _074459_, _074460_, _074461_, _074462_, _074463_, _074464_, _074465_, _074466_, _074467_, _074468_, _074469_, _074470_, _074471_, _074472_, _074473_, _074474_, _074475_, _074476_, _074477_, _074478_, _074479_, _074480_, _074481_, _074482_, _074483_, _074484_, _074485_, _074486_, _074487_, _074488_, _074489_, _074490_, _074491_, _074492_, _074493_, _074494_, _074495_, _074496_, _074497_, _074498_, _074499_, _074500_, _074501_, _074502_, _074503_, _074504_, _074505_, _074506_, _074507_, _074508_, _074509_, _074510_, _074511_, _074512_, _074513_, _074514_, _074515_, _074516_, _074517_, _074518_, _074519_, _074520_, _074521_, _074522_, _074523_, _074524_, _074525_, _074526_, _074527_, _074528_, _074529_, _074530_, _074531_, _074532_, _074533_, _074534_, _074535_, _074536_, _074537_, _074538_, _074539_, _074540_, _074541_, _074542_, _074543_, _074544_, _074545_, _074546_, _074547_, _074548_, _074549_, _074550_, _074551_, _074552_, _074553_, _074554_, _074555_, _074556_, _074557_, _074558_, _074559_, _074560_, _074561_, _074562_, _074563_, _074564_, _074565_, _074566_, _074567_, _074568_, _074569_, _074570_, _074571_, _074572_, _074573_, _074574_, _074575_, _074576_, _074577_, _074578_, _074579_, _074580_, _074581_, _074582_, _074583_, _074584_, _074585_, _074586_, _074587_, _074588_, _074589_, _074590_, _074591_, _074592_, _074593_, _074594_, _074595_, _074596_, _074597_, _074598_, _074599_, _074600_, _074601_, _074602_, _074603_, _074604_, _074605_, _074606_, _074607_, _074608_, _074609_, _074610_, _074611_, _074612_, _074613_, _074614_, _074615_, _074616_, _074617_, _074618_, _074619_, _074620_, _074621_, _074622_, _074623_, _074624_, _074625_, _074626_, _074627_, _074628_, _074629_, _074630_, _074631_, _074632_, _074633_, _074634_, _074635_, _074636_, _074637_, _074638_, _074639_, _074640_, _074641_, _074642_, _074643_, _074644_, _074645_, _074646_, _074647_, _074648_, _074649_, _074650_, _074651_, _074652_, _074653_, _074654_, _074655_, _074656_, _074657_, _074658_, _074659_, _074660_, _074661_, _074662_, _074663_, _074664_, _074665_, _074666_, _074667_, _074668_, _074669_, _074670_, _074671_, _074672_, _074673_, _074674_, _074675_, _074676_, _074677_, _074678_, _074679_, _074680_, _074681_, _074682_, _074683_, _074684_, _074685_, _074686_, _074687_, _074688_, _074689_, _074690_, _074691_, _074692_, _074693_, _074694_, _074695_, _074696_, _074697_, _074698_, _074699_, _074700_, _074701_, _074702_, _074703_, _074704_, _074705_, _074706_, _074707_, _074708_, _074709_, _074710_, _074711_, _074712_, _074713_, _074714_, _074715_, _074716_, _074717_, _074718_, _074719_, _074720_, _074721_, _074722_, _074723_, _074724_, _074725_, _074726_, _074727_, _074728_, _074729_, _074730_, _074731_, _074732_, _074733_, _074734_, _074735_, _074736_, _074737_, _074738_, _074739_, _074740_, _074741_, _074742_, _074743_, _074744_, _074745_, _074746_, _074747_, _074748_, _074749_, _074750_, _074751_, _074752_, _074753_, _074754_, _074755_, _074756_, _074757_, _074758_, _074759_, _074760_, _074761_, _074762_, _074763_, _074764_, _074765_, _074766_, _074767_, _074768_, _074769_, _074770_, _074771_, _074772_, _074773_, _074774_, _074775_, _074776_, _074777_, _074778_, _074779_, _074780_, _074781_, _074782_, _074783_, _074784_, _074785_, _074786_, _074787_, _074788_, _074789_, _074790_, _074791_, _074792_, _074793_, _074794_, _074795_, _074796_, _074797_, _074798_, _074799_, _074800_, _074801_, _074802_, _074803_, _074804_, _074805_, _074806_, _074807_, _074808_, _074809_, _074810_, _074811_, _074812_, _074813_, _074814_, _074815_, _074816_, _074817_, _074818_, _074819_, _074820_, _074821_, _074822_, _074823_, _074824_, _074825_, _074826_, _074827_, _074828_, _074829_, _074830_, _074831_, _074832_, _074833_, _074834_, _074835_, _074836_, _074837_, _074838_, _074839_, _074840_, _074841_, _074842_, _074843_, _074844_, _074845_, _074846_, _074847_, _074848_, _074849_, _074850_, _074851_, _074852_, _074853_, _074854_, _074855_, _074856_, _074857_, _074858_, _074859_, _074860_, _074861_, _074862_, _074863_, _074864_, _074865_, _074866_, _074867_, _074868_, _074869_, _074870_, _074871_, _074872_, _074873_, _074874_, _074875_, _074876_, _074877_, _074878_, _074879_, _074880_, _074881_, _074882_, _074883_, _074884_, _074885_, _074886_, _074887_, _074888_, _074889_, _074890_, _074891_, _074892_, _074893_, _074894_, _074895_, _074896_, _074897_, _074898_, _074899_, _074900_, _074901_, _074902_, _074903_, _074904_, _074905_, _074906_, _074907_, _074908_, _074909_, _074910_, _074911_, _074912_, _074913_, _074914_, _074915_, _074916_, _074917_, _074918_, _074919_, _074920_, _074921_, _074922_, _074923_, _074924_, _074925_, _074926_, _074927_, _074928_, _074929_, _074930_, _074931_, _074932_, _074933_, _074934_, _074935_, _074936_, _074937_, _074938_, _074939_, _074940_, _074941_, _074942_, _074943_, _074944_, _074945_, _074946_, _074947_, _074948_, _074949_, _074950_, _074951_, _074952_, _074953_, _074954_, _074955_, _074956_, _074957_, _074958_, _074959_, _074960_, _074961_, _074962_, _074963_, _074964_, _074965_, _074966_, _074967_, _074968_, _074969_, _074970_, _074971_, _074972_, _074973_, _074974_, _074975_, _074976_, _074977_, _074978_, _074979_, _074980_, _074981_, _074982_, _074983_, _074984_, _074985_, _074986_, _074987_, _074988_, _074989_, _074990_, _074991_, _074992_, _074993_, _074994_, _074995_, _074996_, _074997_, _074998_, _074999_, _075000_, _075001_, _075002_, _075003_, _075004_, _075005_, _075006_, _075007_, _075008_, _075009_, _075010_, _075011_, _075012_, _075013_, _075014_, _075015_, _075016_, _075017_, _075018_, _075019_, _075020_, _075021_, _075022_, _075023_, _075024_, _075025_, _075026_, _075027_, _075028_, _075029_, _075030_, _075031_, _075032_, _075033_, _075034_, _075035_, _075036_, _075037_, _075038_, _075039_, _075040_, _075041_, _075042_, _075043_, _075044_, _075045_, _075046_, _075047_, _075048_, _075049_, _075050_, _075051_, _075052_, _075053_, _075054_, _075055_, _075056_, _075057_, _075058_, _075059_, _075060_, _075061_, _075062_, _075063_, _075064_, _075065_, _075066_, _075067_, _075068_, _075069_, _075070_, _075071_, _075072_, _075073_, _075074_, _075075_, _075076_, _075077_, _075078_, _075079_, _075080_, _075081_, _075082_, _075083_, _075084_, _075085_, _075086_, _075087_, _075088_, _075089_, _075090_, _075091_, _075092_, _075093_, _075094_, _075095_, _075096_, _075097_, _075098_, _075099_, _075100_, _075101_, _075102_, _075103_, _075104_, _075105_, _075106_, _075107_, _075108_, _075109_, _075110_, _075111_, _075112_, _075113_, _075114_, _075115_, _075116_, _075117_, _075118_, _075119_, _075120_, _075121_, _075122_, _075123_, _075124_, _075125_, _075126_, _075127_, _075128_, _075129_, _075130_, _075131_, _075132_, _075133_, _075134_, _075135_, _075136_, _075137_, _075138_, _075139_, _075140_, _075141_, _075142_, _075143_, _075144_, _075145_, _075146_, _075147_, _075148_, _075149_, _075150_, _075151_, _075152_, _075153_, _075154_, _075155_, _075156_, _075157_, _075158_, _075159_, _075160_, _075161_, _075162_, _075163_, _075164_, _075165_, _075166_, _075167_, _075168_, _075169_, _075170_, _075171_, _075172_, _075173_, _075174_, _075175_, _075176_, _075177_, _075178_, _075179_, _075180_, _075181_, _075182_, _075183_, _075184_, _075185_, _075186_, _075187_, _075188_, _075189_, _075190_, _075191_, _075192_, _075193_, _075194_, _075195_, _075196_, _075197_, _075198_, _075199_, _075200_, _075201_, _075202_, _075203_, _075204_, _075205_, _075206_, _075207_, _075208_, _075209_, _075210_, _075211_, _075212_, _075213_, _075214_, _075215_, _075216_, _075217_, _075218_, _075219_, _075220_, _075221_, _075222_, _075223_, _075224_, _075225_, _075226_, _075227_, _075228_, _075229_, _075230_, _075231_, _075232_, _075233_, _075234_, _075235_, _075236_, _075237_, _075238_, _075239_, _075240_, _075241_, _075242_, _075243_, _075244_, _075245_, _075246_, _075247_, _075248_, _075249_, _075250_, _075251_, _075252_, _075253_, _075254_, _075255_, _075256_, _075257_, _075258_, _075259_, _075260_, _075261_, _075262_, _075263_, _075264_, _075265_, _075266_, _075267_, _075268_, _075269_, _075270_, _075271_, _075272_, _075273_, _075274_, _075275_, _075276_, _075277_, _075278_, _075279_, _075280_, _075281_, _075282_, _075283_, _075284_, _075285_, _075286_, _075287_, _075288_, _075289_, _075290_, _075291_, _075292_, _075293_, _075294_, _075295_, _075296_, _075297_, _075298_, _075299_, _075300_, _075301_, _075302_, _075303_, _075304_, _075305_, _075306_, _075307_, _075308_, _075309_, _075310_, _075311_, _075312_, _075313_, _075314_, _075315_, _075316_, _075317_, _075318_, _075319_, _075320_, _075321_, _075322_, _075323_, _075324_, _075325_, _075326_, _075327_, _075328_, _075329_, _075330_, _075331_, _075332_, _075333_, _075334_, _075335_, _075336_, _075337_, _075338_, _075339_, _075340_, _075341_, _075342_, _075343_, _075344_, _075345_, _075346_, _075347_, _075348_, _075349_, _075350_, _075351_, _075352_, _075353_, _075354_, _075355_, _075356_, _075357_, _075358_, _075359_, _075360_, _075361_, _075362_, _075363_, _075364_, _075365_, _075366_, _075367_, _075368_, _075369_, _075370_, _075371_, _075372_, _075373_, _075374_, _075375_, _075376_, _075377_, _075378_, _075379_, _075380_, _075381_, _075382_, _075383_, _075384_, _075385_, _075386_, _075387_, _075388_, _075389_, _075390_, _075391_, _075392_, _075393_, _075394_, _075395_, _075396_, _075397_, _075398_, _075399_, _075400_, _075401_, _075402_, _075403_, _075404_, _075405_, _075406_, _075407_, _075408_, _075409_, _075410_, _075411_, _075412_, _075413_, _075414_, _075415_, _075416_, _075417_, _075418_, _075419_, _075420_, _075421_, _075422_, _075423_, _075424_, _075425_, _075426_, _075427_, _075428_, _075429_, _075430_, _075431_, _075432_, _075433_, _075434_, _075435_, _075436_, _075437_, _075438_, _075439_, _075440_, _075441_, _075442_, _075443_, _075444_, _075445_, _075446_, _075447_, _075448_, _075449_, _075450_, _075451_, _075452_, _075453_, _075454_, _075455_, _075456_, _075457_, _075458_, _075459_, _075460_, _075461_, _075462_, _075463_, _075464_, _075465_, _075466_, _075467_, _075468_, _075469_, _075470_, _075471_, _075472_, _075473_, _075474_, _075475_, _075476_, _075477_, _075478_, _075479_, _075480_, _075481_, _075482_, _075483_, _075484_, _075485_, _075486_, _075487_, _075488_, _075489_, _075490_, _075491_, _075492_, _075493_, _075494_, _075495_, _075496_, _075497_, _075498_, _075499_, _075500_, _075501_, _075502_, _075503_, _075504_, _075505_, _075506_, _075507_, _075508_, _075509_, _075510_, _075511_, _075512_, _075513_, _075514_, _075515_, _075516_, _075517_, _075518_, _075519_, _075520_, _075521_, _075522_, _075523_, _075524_, _075525_, _075526_, _075527_, _075528_, _075529_, _075530_, _075531_, _075532_, _075533_, _075534_, _075535_, _075536_, _075537_, _075538_, _075539_, _075540_, _075541_, _075542_, _075543_, _075544_, _075545_, _075546_, _075547_, _075548_, _075549_, _075550_, _075551_, _075552_, _075553_, _075554_, _075555_, _075556_, _075557_, _075558_, _075559_, _075560_, _075561_, _075562_, _075563_, _075564_, _075565_, _075566_, _075567_, _075568_, _075569_, _075570_, _075571_, _075572_, _075573_, _075574_, _075575_, _075576_, _075577_, _075578_, _075579_, _075580_, _075581_, _075582_, _075583_, _075584_, _075585_, _075586_, _075587_, _075588_, _075589_, _075590_, _075591_, _075592_, _075593_, _075594_, _075595_, _075596_, _075597_, _075598_, _075599_, _075600_, _075601_, _075602_, _075603_, _075604_, _075605_, _075606_, _075607_, _075608_, _075609_, _075610_, _075611_, _075612_, _075613_, _075614_, _075615_, _075616_, _075617_, _075618_, _075619_, _075620_, _075621_, _075622_, _075623_, _075624_, _075625_, _075626_, _075627_, _075628_, _075629_, _075630_, _075631_, _075632_, _075633_, _075634_, _075635_, _075636_, _075637_, _075638_, _075639_, _075640_, _075641_, _075642_, _075643_, _075644_, _075645_, _075646_, _075647_, _075648_, _075649_, _075650_, _075651_, _075652_, _075653_, _075654_, _075655_, _075656_, _075657_, _075658_, _075659_, _075660_, _075661_, _075662_, _075663_, _075664_, _075665_, _075666_, _075667_, _075668_, _075669_, _075670_, _075671_, _075672_, _075673_, _075674_, _075675_, _075676_, _075677_, _075678_, _075679_, _075680_, _075681_, _075682_, _075683_, _075684_, _075685_, _075686_, _075687_, _075688_, _075689_, _075690_, _075691_, _075692_, _075693_, _075694_, _075695_, _075696_, _075697_, _075698_, _075699_, _075700_, _075701_, _075702_, _075703_, _075704_, _075705_, _075706_, _075707_, _075708_, _075709_, _075710_, _075711_, _075712_, _075713_, _075714_, _075715_, _075716_, _075717_, _075718_, _075719_, _075720_, _075721_, _075722_, _075723_, _075724_, _075725_, _075726_, _075727_, _075728_, _075729_, _075730_, _075731_, _075732_, _075733_, _075734_, _075735_, _075736_, _075737_, _075738_, _075739_, _075740_, _075741_, _075742_, _075743_, _075744_, _075745_, _075746_, _075747_, _075748_, _075749_, _075750_, _075751_, _075752_, _075753_, _075754_, _075755_, _075756_, _075757_, _075758_, _075759_, _075760_, _075761_, _075762_, _075763_, _075764_, _075765_, _075766_, _075767_, _075768_, _075769_, _075770_, _075771_, _075772_, _075773_, _075774_, _075775_, _075776_, _075777_, _075778_, _075779_, _075780_, _075781_, _075782_, _075783_, _075784_, _075785_, _075786_, _075787_, _075788_, _075789_, _075790_, _075791_, _075792_, _075793_, _075794_, _075795_, _075796_, _075797_, _075798_, _075799_, _075800_, _075801_, _075802_, _075803_, _075804_, _075805_, _075806_, _075807_, _075808_, _075809_, _075810_, _075811_, _075812_, _075813_, _075814_, _075815_, _075816_, _075817_, _075818_, _075819_, _075820_, _075821_, _075822_, _075823_, _075824_, _075825_, _075826_, _075827_, _075828_, _075829_, _075830_, _075831_, _075832_, _075833_, _075834_, _075835_, _075836_, _075837_, _075838_, _075839_, _075840_, _075841_, _075842_, _075843_, _075844_, _075845_, _075846_, _075847_, _075848_, _075849_, _075850_, _075851_, _075852_, _075853_, _075854_, _075855_, _075856_, _075857_, _075858_, _075859_, _075860_, _075861_, _075862_, _075863_, _075864_, _075865_, _075866_, _075867_, _075868_, _075869_, _075870_, _075871_, _075872_, _075873_, _075874_, _075875_, _075876_, _075877_, _075878_, _075879_, _075880_, _075881_, _075882_, _075883_, _075884_, _075885_, _075886_, _075887_, _075888_, _075889_, _075890_, _075891_, _075892_, _075893_, _075894_, _075895_, _075896_, _075897_, _075898_, _075899_, _075900_, _075901_, _075902_, _075903_, _075904_, _075905_, _075906_, _075907_, _075908_, _075909_, _075910_, _075911_, _075912_, _075913_, _075914_, _075915_, _075916_, _075917_, _075918_, _075919_, _075920_, _075921_, _075922_, _075923_, _075924_, _075925_, _075926_, _075927_, _075928_, _075929_, _075930_, _075931_, _075932_, _075933_, _075934_, _075935_, _075936_, _075937_, _075938_, _075939_, _075940_, _075941_, _075942_, _075943_, _075944_, _075945_, _075946_, _075947_, _075948_, _075949_, _075950_, _075951_, _075952_, _075953_, _075954_, _075955_, _075956_, _075957_, _075958_, _075959_, _075960_, _075961_, _075962_, _075963_, _075964_, _075965_, _075966_, _075967_, _075968_, _075969_, _075970_, _075971_, _075972_, _075973_, _075974_, _075975_, _075976_, _075977_, _075978_, _075979_, _075980_, _075981_, _075982_, _075983_, _075984_, _075985_, _075986_, _075987_, _075988_, _075989_, _075990_, _075991_, _075992_, _075993_, _075994_, _075995_, _075996_, _075997_, _075998_, _075999_, _076000_, _076001_, _076002_, _076003_, _076004_, _076005_, _076006_, _076007_, _076008_, _076009_, _076010_, _076011_, _076012_, _076013_, _076014_, _076015_, _076016_, _076017_, _076018_, _076019_, _076020_, _076021_, _076022_, _076023_, _076024_, _076025_, _076026_, _076027_, _076028_, _076029_, _076030_, _076031_, _076032_, _076033_, _076034_, _076035_, _076036_, _076037_, _076038_, _076039_, _076040_, _076041_, _076042_, _076043_, _076044_, _076045_, _076046_, _076047_, _076048_, _076049_, _076050_, _076051_, _076052_, _076053_, _076054_, _076055_, _076056_, _076057_, _076058_, _076059_, _076060_, _076061_, _076062_, _076063_, _076064_, _076065_, _076066_, _076067_, _076068_, _076069_, _076070_, _076071_, _076072_, _076073_, _076074_, _076075_, _076076_, _076077_, _076078_, _076079_, _076080_, _076081_, _076082_, _076083_, _076084_, _076085_, _076086_, _076087_, _076088_, _076089_, _076090_, _076091_, _076092_, _076093_, _076094_, _076095_, _076096_, _076097_, _076098_, _076099_, _076100_, _076101_, _076102_, _076103_, _076104_, _076105_, _076106_, _076107_, _076108_, _076109_, _076110_, _076111_, _076112_, _076113_, _076114_, _076115_, _076116_, _076117_, _076118_, _076119_, _076120_, _076121_, _076122_, _076123_, _076124_, _076125_, _076126_, _076127_, _076128_, _076129_, _076130_, _076131_, _076132_, _076133_, _076134_, _076135_, _076136_, _076137_, _076138_, _076139_, _076140_, _076141_, _076142_, _076143_, _076144_, _076145_, _076146_, _076147_, _076148_, _076149_, _076150_, _076151_, _076152_, _076153_, _076154_, _076155_, _076156_, _076157_, _076158_, _076159_, _076160_, _076161_, _076162_, _076163_, _076164_, _076165_, _076166_, _076167_, _076168_, _076169_, _076170_, _076171_, _076172_, _076173_, _076174_, _076175_, _076176_, _076177_, _076178_, _076179_, _076180_, _076181_, _076182_, _076183_, _076184_, _076185_, _076186_, _076187_, _076188_, _076189_, _076190_, _076191_, _076192_, _076193_, _076194_, _076195_, _076196_, _076197_, _076198_, _076199_, _076200_, _076201_, _076202_, _076203_, _076204_, _076205_, _076206_, _076207_, _076208_, _076209_, _076210_, _076211_, _076212_, _076213_, _076214_, _076215_, _076216_, _076217_, _076218_, _076219_, _076220_, _076221_, _076222_, _076223_, _076224_, _076225_, _076226_, _076227_, _076228_, _076229_, _076230_, _076231_, _076232_, _076233_, _076234_, _076235_, _076236_, _076237_, _076238_, _076239_, _076240_, _076241_, _076242_, _076243_, _076244_, _076245_, _076246_, _076247_, _076248_, _076249_, _076250_, _076251_, _076252_, _076253_, _076254_, _076255_, _076256_, _076257_, _076258_, _076259_, _076260_, _076261_, _076262_, _076263_, _076264_, _076265_, _076266_, _076267_, _076268_, _076269_, _076270_, _076271_, _076272_, _076273_, _076274_, _076275_, _076276_, _076277_, _076278_, _076279_, _076280_, _076281_, _076282_, _076283_, _076284_, _076285_, _076286_, _076287_, _076288_, _076289_, _076290_, _076291_, _076292_, _076293_, _076294_, _076295_, _076296_, _076297_, _076298_, _076299_, _076300_, _076301_, _076302_, _076303_, _076304_, _076305_, _076306_, _076307_, _076308_, _076309_, _076310_, _076311_, _076312_, _076313_, _076314_, _076315_, _076316_, _076317_, _076318_, _076319_, _076320_, _076321_, _076322_, _076323_, _076324_, _076325_, _076326_, _076327_, _076328_, _076329_, _076330_, _076331_, _076332_, _076333_, _076334_, _076335_, _076336_, _076337_, _076338_, _076339_, _076340_, _076341_, _076342_, _076343_, _076344_, _076345_, _076346_, _076347_, _076348_, _076349_, _076350_, _076351_, _076352_, _076353_, _076354_, _076355_, _076356_, _076357_, _076358_, _076359_, _076360_, _076361_, _076362_, _076363_, _076364_, _076365_, _076366_, _076367_, _076368_, _076369_, _076370_, _076371_, _076372_, _076373_, _076374_, _076375_, _076376_, _076377_, _076378_, _076379_, _076380_, _076381_, _076382_, _076383_, _076384_, _076385_, _076386_, _076387_, _076388_, _076389_, _076390_, _076391_, _076392_, _076393_, _076394_, _076395_, _076396_, _076397_, _076398_, _076399_, _076400_, _076401_, _076402_, _076403_, _076404_, _076405_, _076406_, _076407_, _076408_, _076409_, _076410_, _076411_, _076412_, _076413_, _076414_, _076415_, _076416_, _076417_, _076418_, _076419_, _076420_, _076421_, _076422_, _076423_, _076424_, _076425_, _076426_, _076427_, _076428_, _076429_, _076430_, _076431_, _076432_, _076433_, _076434_, _076435_, _076436_, _076437_, _076438_, _076439_, _076440_, _076441_, _076442_, _076443_, _076444_, _076445_, _076446_, _076447_, _076448_, _076449_, _076450_, _076451_, _076452_, _076453_, _076454_, _076455_, _076456_, _076457_, _076458_, _076459_, _076460_, _076461_, _076462_, _076463_, _076464_, _076465_, _076466_, _076467_, _076468_, _076469_, _076470_, _076471_, _076472_, _076473_, _076474_, _076475_, _076476_, _076477_, _076478_, _076479_, _076480_, _076481_, _076482_, _076483_, _076484_, _076485_, _076486_, _076487_, _076488_, _076489_, _076490_, _076491_, _076492_, _076493_, _076494_, _076495_, _076496_, _076497_, _076498_, _076499_, _076500_, _076501_, _076502_, _076503_, _076504_, _076505_, _076506_, _076507_, _076508_, _076509_, _076510_, _076511_, _076512_, _076513_, _076514_, _076515_, _076516_, _076517_, _076518_, _076519_, _076520_, _076521_, _076522_, _076523_, _076524_, _076525_, _076526_, _076527_, _076528_, _076529_, _076530_, _076531_, _076532_, _076533_, _076534_, _076535_, _076536_, _076537_, _076538_, _076539_, _076540_, _076541_, _076542_, _076543_, _076544_, _076545_, _076546_, _076547_, _076548_, _076549_, _076550_, _076551_, _076552_, _076553_, _076554_, _076555_, _076556_, _076557_, _076558_, _076559_, _076560_, _076561_, _076562_, _076563_, _076564_, _076565_, _076566_, _076567_, _076568_, _076569_, _076570_, _076571_, _076572_, _076573_, _076574_, _076575_, _076576_, _076577_, _076578_, _076579_, _076580_, _076581_, _076582_, _076583_, _076584_, _076585_, _076586_, _076587_, _076588_, _076589_, _076590_, _076591_, _076592_, _076593_, _076594_, _076595_, _076596_, _076597_, _076598_, _076599_, _076600_, _076601_, _076602_, _076603_, _076604_, _076605_, _076606_, _076607_, _076608_, _076609_, _076610_, _076611_, _076612_, _076613_, _076614_, _076615_, _076616_, _076617_, _076618_, _076619_, _076620_, _076621_, _076622_, _076623_, _076624_, _076625_, _076626_, _076627_, _076628_, _076629_, _076630_, _076631_, _076632_, _076633_, _076634_, _076635_, _076636_, _076637_, _076638_, _076639_, _076640_, _076641_, _076642_, _076643_, _076644_, _076645_, _076646_, _076647_, _076648_, _076649_, _076650_, _076651_, _076652_, _076653_, _076654_, _076655_, _076656_, _076657_, _076658_, _076659_, _076660_, _076661_, _076662_, _076663_, _076664_, _076665_, _076666_, _076667_, _076668_, _076669_, _076670_, _076671_, _076672_, _076673_, _076674_, _076675_, _076676_, _076677_, _076678_, _076679_, _076680_, _076681_, _076682_, _076683_, _076684_, _076685_, _076686_, _076687_, _076688_, _076689_, _076690_, _076691_, _076692_, _076693_, _076694_, _076695_, _076696_, _076697_, _076698_, _076699_, _076700_, _076701_, _076702_, _076703_, _076704_, _076705_, _076706_, _076707_, _076708_, _076709_, _076710_, _076711_, _076712_, _076713_, _076714_, _076715_, _076716_, _076717_, _076718_, _076719_, _076720_, _076721_, _076722_, _076723_, _076724_, _076725_, _076726_, _076727_, _076728_, _076729_, _076730_, _076731_, _076732_, _076733_, _076734_, _076735_, _076736_, _076737_, _076738_, _076739_, _076740_, _076741_, _076742_, _076743_, _076744_, _076745_, _076746_, _076747_, _076748_, _076749_, _076750_, _076751_, _076752_, _076753_, _076754_, _076755_, _076756_, _076757_, _076758_, _076759_, _076760_, _076761_, _076762_, _076763_, _076764_, _076765_, _076766_, _076767_, _076768_, _076769_, _076770_, _076771_, _076772_, _076773_, _076774_, _076775_, _076776_, _076777_, _076778_, _076779_, _076780_, _076781_, _076782_, _076783_, _076784_, _076785_, _076786_, _076787_, _076788_, _076789_, _076790_, _076791_, _076792_, _076793_, _076794_, _076795_, _076796_, _076797_, _076798_, _076799_, _076800_, _076801_, _076802_, _076803_, _076804_, _076805_, _076806_, _076807_, _076808_, _076809_, _076810_, _076811_, _076812_, _076813_, _076814_, _076815_, _076816_, _076817_, _076818_, _076819_, _076820_, _076821_, _076822_, _076823_, _076824_, _076825_, _076826_, _076827_, _076828_, _076829_, _076830_, _076831_, _076832_, _076833_, _076834_, _076835_, _076836_, _076837_, _076838_, _076839_, _076840_, _076841_, _076842_, _076843_, _076844_, _076845_, _076846_, _076847_, _076848_, _076849_, _076850_, _076851_, _076852_, _076853_, _076854_, _076855_, _076856_, _076857_, _076858_, _076859_, _076860_, _076861_, _076862_, _076863_, _076864_, _076865_, _076866_, _076867_, _076868_, _076869_, _076870_, _076871_, _076872_, _076873_, _076874_, _076875_, _076876_, _076877_, _076878_, _076879_, _076880_, _076881_, _076882_, _076883_, _076884_, _076885_, _076886_, _076887_, _076888_, _076889_, _076890_, _076891_, _076892_, _076893_, _076894_, _076895_, _076896_, _076897_, _076898_, _076899_, _076900_, _076901_, _076902_, _076903_, _076904_, _076905_, _076906_, _076907_, _076908_, _076909_, _076910_, _076911_, _076912_, _076913_, _076914_, _076915_, _076916_, _076917_, _076918_, _076919_, _076920_, _076921_, _076922_, _076923_, _076924_, _076925_, _076926_, _076927_, _076928_, _076929_, _076930_, _076931_, _076932_, _076933_, _076934_, _076935_, _076936_, _076937_, _076938_, _076939_, _076940_, _076941_, _076942_, _076943_, _076944_, _076945_, _076946_, _076947_, _076948_, _076949_, _076950_, _076951_, _076952_, _076953_, _076954_, _076955_, _076956_, _076957_, _076958_, _076959_, _076960_, _076961_, _076962_, _076963_, _076964_, _076965_, _076966_, _076967_, _076968_, _076969_, _076970_, _076971_, _076972_, _076973_, _076974_, _076975_, _076976_, _076977_, _076978_, _076979_, _076980_, _076981_, _076982_, _076983_, _076984_, _076985_, _076986_, _076987_, _076988_, _076989_, _076990_, _076991_, _076992_, _076993_, _076994_, _076995_, _076996_, _076997_, _076998_, _076999_, _077000_, _077001_, _077002_, _077003_, _077004_, _077005_, _077006_, _077007_, _077008_, _077009_, _077010_, _077011_, _077012_, _077013_, _077014_, _077015_, _077016_, _077017_, _077018_, _077019_, _077020_, _077021_, _077022_, _077023_, _077024_, _077025_, _077026_, _077027_, _077028_, _077029_, _077030_, _077031_, _077032_, _077033_, _077034_, _077035_, _077036_, _077037_, _077038_, _077039_, _077040_, _077041_, _077042_, _077043_, _077044_, _077045_, _077046_, _077047_, _077048_, _077049_, _077050_, _077051_, _077052_, _077053_, _077054_, _077055_, _077056_, _077057_, _077058_, _077059_, _077060_, _077061_, _077062_, _077063_, _077064_, _077065_, _077066_, _077067_, _077068_, _077069_, _077070_, _077071_, _077072_, _077073_, _077074_, _077075_, _077076_, _077077_, _077078_, _077079_, _077080_, _077081_, _077082_, _077083_, _077084_, _077085_, _077086_, _077087_, _077088_, _077089_, _077090_, _077091_, _077092_, _077093_, _077094_, _077095_, _077096_, _077097_, _077098_, _077099_, _077100_, _077101_, _077102_, _077103_, _077104_, _077105_, _077106_, _077107_, _077108_, _077109_, _077110_, _077111_, _077112_, _077113_, _077114_, _077115_, _077116_, _077117_, _077118_, _077119_, _077120_, _077121_, _077122_, _077123_, _077124_, _077125_, _077126_, _077127_, _077128_, _077129_, _077130_, _077131_, _077132_, _077133_, _077134_, _077135_, _077136_, _077137_, _077138_, _077139_, _077140_, _077141_, _077142_, _077143_, _077144_, _077145_, _077146_, _077147_, _077148_, _077149_, _077150_, _077151_, _077152_, _077153_, _077154_, _077155_, _077156_, _077157_, _077158_, _077159_, _077160_, _077161_, _077162_, _077163_, _077164_, _077165_, _077166_, _077167_, _077168_, _077169_, _077170_, _077171_, _077172_, _077173_, _077174_, _077175_, _077176_, _077177_, _077178_, _077179_, _077180_, _077181_, _077182_, _077183_, _077184_, _077185_, _077186_, _077187_, _077188_, _077189_, _077190_, _077191_, _077192_, _077193_, _077194_, _077195_, _077196_, _077197_, _077198_, _077199_, _077200_, _077201_, _077202_, _077203_, _077204_, _077205_, _077206_, _077207_, _077208_, _077209_, _077210_, _077211_, _077212_, _077213_, _077214_, _077215_, _077216_, _077217_, _077218_, _077219_, _077220_, _077221_, _077222_, _077223_, _077224_, _077225_, _077226_, _077227_, _077228_, _077229_, _077230_, _077231_, _077232_, _077233_, _077234_, _077235_, _077236_, _077237_, _077238_, _077239_, _077240_, _077241_, _077242_, _077243_, _077244_, _077245_, _077246_, _077247_, _077248_, _077249_, _077250_, _077251_, _077252_, _077253_, _077254_, _077255_, _077256_, _077257_, _077258_, _077259_, _077260_, _077261_, _077262_, _077263_, _077264_, _077265_, _077266_, _077267_, _077268_, _077269_, _077270_, _077271_, _077272_, _077273_, _077274_, _077275_, _077276_, _077277_, _077278_, _077279_, _077280_, _077281_, _077282_, _077283_, _077284_, _077285_, _077286_, _077287_, _077288_, _077289_, _077290_, _077291_, _077292_, _077293_, _077294_, _077295_, _077296_, _077297_, _077298_, _077299_, _077300_, _077301_, _077302_, _077303_, _077304_, _077305_, _077306_, _077307_, _077308_, _077309_, _077310_, _077311_, _077312_, _077313_, _077314_, _077315_, _077316_, _077317_, _077318_, _077319_, _077320_, _077321_, _077322_, _077323_, _077324_, _077325_, _077326_, _077327_, _077328_, _077329_, _077330_, _077331_, _077332_, _077333_, _077334_, _077335_, _077336_, _077337_, _077338_, _077339_, _077340_, _077341_, _077342_, _077343_, _077344_, _077345_, _077346_, _077347_, _077348_, _077349_, _077350_, _077351_, _077352_, _077353_, _077354_, _077355_, _077356_, _077357_, _077358_, _077359_, _077360_, _077361_, _077362_, _077363_, _077364_, _077365_, _077366_, _077367_, _077368_, _077369_, _077370_, _077371_, _077372_, _077373_, _077374_, _077375_, _077376_, _077377_, _077378_, _077379_, _077380_, _077381_, _077382_, _077383_, _077384_, _077385_, _077386_, _077387_, _077388_, _077389_, _077390_, _077391_, _077392_, _077393_, _077394_, _077395_, _077396_, _077397_, _077398_, _077399_, _077400_, _077401_, _077402_, _077403_, _077404_, _077405_, _077406_, _077407_, _077408_, _077409_, _077410_, _077411_, _077412_, _077413_, _077414_, _077415_, _077416_, _077417_, _077418_, _077419_, _077420_, _077421_, _077422_, _077423_, _077424_, _077425_, _077426_, _077427_, _077428_, _077429_, _077430_, _077431_, _077432_, _077433_, _077434_, _077435_, _077436_, _077437_, _077438_, _077439_, _077440_, _077441_, _077442_, _077443_, _077444_, _077445_, _077446_, _077447_, _077448_, _077449_, _077450_, _077451_, _077452_, _077453_, _077454_, _077455_, _077456_, _077457_, _077458_, _077459_, _077460_, _077461_, _077462_, _077463_, _077464_, _077465_, _077466_, _077467_, _077468_, _077469_, _077470_, _077471_, _077472_, _077473_, _077474_, _077475_, _077476_, _077477_, _077478_, _077479_, _077480_, _077481_, _077482_, _077483_, _077484_, _077485_, _077486_, _077487_, _077488_, _077489_, _077490_, _077491_, _077492_, _077493_, _077494_, _077495_, _077496_, _077497_, _077498_, _077499_, _077500_, _077501_, _077502_, _077503_, _077504_, _077505_, _077506_, _077507_, _077508_, _077509_, _077510_, _077511_, _077512_, _077513_, _077514_, _077515_, _077516_, _077517_, _077518_, _077519_, _077520_, _077521_, _077522_, _077523_, _077524_, _077525_, _077526_, _077527_, _077528_, _077529_, _077530_, _077531_, _077532_, _077533_, _077534_, _077535_, _077536_, _077537_, _077538_, _077539_, _077540_, _077541_, _077542_, _077543_, _077544_, _077545_, _077546_, _077547_, _077548_, _077549_, _077550_, _077551_, _077552_, _077553_, _077554_, _077555_, _077556_, _077557_, _077558_, _077559_, _077560_, _077561_, _077562_, _077563_, _077564_, _077565_, _077566_, _077567_, _077568_, _077569_, _077570_, _077571_, _077572_, _077573_, _077574_, _077575_, _077576_, _077577_, _077578_, _077579_, _077580_, _077581_, _077582_, _077583_, _077584_, _077585_, _077586_, _077587_, _077588_, _077589_, _077590_, _077591_, _077592_, _077593_, _077594_, _077595_, _077596_, _077597_, _077598_, _077599_, _077600_, _077601_, _077602_, _077603_, _077604_, _077605_, _077606_, _077607_, _077608_, _077609_, _077610_, _077611_, _077612_, _077613_, _077614_, _077615_, _077616_, _077617_, _077618_, _077619_, _077620_, _077621_, _077622_, _077623_, _077624_, _077625_, _077626_, _077627_, _077628_, _077629_, _077630_, _077631_, _077632_, _077633_, _077634_, _077635_, _077636_, _077637_, _077638_, _077639_, _077640_, _077641_, _077642_, _077643_, _077644_, _077645_, _077646_, _077647_, _077648_, _077649_, _077650_, _077651_, _077652_, _077653_, _077654_, _077655_, _077656_, _077657_, _077658_, _077659_, _077660_, _077661_, _077662_, _077663_, _077664_, _077665_, _077666_, _077667_, _077668_, _077669_, _077670_, _077671_, _077672_, _077673_, _077674_, _077675_, _077676_, _077677_, _077678_, _077679_, _077680_, _077681_, _077682_, _077683_, _077684_, _077685_, _077686_, _077687_, _077688_, _077689_, _077690_, _077691_, _077692_, _077693_, _077694_, _077695_, _077696_, _077697_, _077698_, _077699_, _077700_, _077701_, _077702_, _077703_, _077704_, _077705_, _077706_, _077707_, _077708_, _077709_, _077710_, _077711_, _077712_, _077713_, _077714_, _077715_, _077716_, _077717_, _077718_, _077719_, _077720_, _077721_, _077722_, _077723_, _077724_, _077725_, _077726_, _077727_, _077728_, _077729_, _077730_, _077731_, _077732_, _077733_, _077734_, _077735_, _077736_, _077737_, _077738_, _077739_, _077740_, _077741_, _077742_, _077743_, _077744_, _077745_, _077746_, _077747_, _077748_, _077749_, _077750_, _077751_, _077752_, _077753_, _077754_, _077755_, _077756_, _077757_, _077758_, _077759_, _077760_, _077761_, _077762_, _077763_, _077764_, _077765_, _077766_, _077767_, _077768_, _077769_, _077770_, _077771_, _077772_, _077773_, _077774_, _077775_, _077776_, _077777_, _077778_, _077779_, _077780_, _077781_, _077782_, _077783_, _077784_, _077785_, _077786_, _077787_, _077788_, _077789_, _077790_, _077791_, _077792_, _077793_, _077794_, _077795_, _077796_, _077797_, _077798_, _077799_, _077800_, _077801_, _077802_, _077803_, _077804_, _077805_, _077806_, _077807_, _077808_, _077809_, _077810_, _077811_, _077812_, _077813_, _077814_, _077815_, _077816_, _077817_, _077818_, _077819_, _077820_, _077821_, _077822_, _077823_, _077824_, _077825_, _077826_, _077827_, _077828_, _077829_, _077830_, _077831_, _077832_, _077833_, _077834_, _077835_, _077836_, _077837_, _077838_, _077839_, _077840_, _077841_, _077842_, _077843_, _077844_, _077845_, _077846_, _077847_, _077848_, _077849_, _077850_, _077851_, _077852_, _077853_, _077854_, _077855_, _077856_, _077857_, _077858_, _077859_, _077860_, _077861_, _077862_, _077863_, _077864_, _077865_, _077866_, _077867_, _077868_, _077869_, _077870_, _077871_, _077872_, _077873_, _077874_, _077875_, _077876_, _077877_, _077878_, _077879_, _077880_, _077881_, _077882_, _077883_, _077884_, _077885_, _077886_, _077887_, _077888_, _077889_, _077890_, _077891_, _077892_, _077893_, _077894_, _077895_, _077896_, _077897_, _077898_, _077899_, _077900_, _077901_, _077902_, _077903_, _077904_, _077905_, _077906_, _077907_, _077908_, _077909_, _077910_, _077911_, _077912_, _077913_, _077914_, _077915_, _077916_, _077917_, _077918_, _077919_, _077920_, _077921_, _077922_, _077923_, _077924_, _077925_, _077926_, _077927_, _077928_, _077929_, _077930_, _077931_, _077932_, _077933_, _077934_, _077935_, _077936_, _077937_, _077938_, _077939_, _077940_, _077941_, _077942_, _077943_, _077944_, _077945_, _077946_, _077947_, _077948_, _077949_, _077950_, _077951_, _077952_, _077953_, _077954_, _077955_, _077956_, _077957_, _077958_, _077959_, _077960_, _077961_, _077962_, _077963_, _077964_, _077965_, _077966_, _077967_, _077968_, _077969_, _077970_, _077971_, _077972_, _077973_, _077974_, _077975_, _077976_, _077977_, _077978_, _077979_, _077980_, _077981_, _077982_, _077983_, _077984_, _077985_, _077986_, _077987_, _077988_, _077989_, _077990_, _077991_, _077992_, _077993_, _077994_, _077995_, _077996_, _077997_, _077998_, _077999_, _078000_, _078001_, _078002_, _078003_, _078004_, _078005_, _078006_, _078007_, _078008_, _078009_, _078010_, _078011_, _078012_, _078013_, _078014_, _078015_, _078016_, _078017_, _078018_, _078019_, _078020_, _078021_, _078022_, _078023_, _078024_, _078025_, _078026_, _078027_, _078028_, _078029_, _078030_, _078031_, _078032_, _078033_, _078034_, _078035_, _078036_, _078037_, _078038_, _078039_, _078040_, _078041_, _078042_, _078043_, _078044_, _078045_, _078046_, _078047_, _078048_, _078049_, _078050_, _078051_, _078052_, _078053_, _078054_, _078055_, _078056_, _078057_, _078058_, _078059_, _078060_, _078061_, _078062_, _078063_, _078064_, _078065_, _078066_, _078067_, _078068_, _078069_, _078070_, _078071_, _078072_, _078073_, _078074_, _078075_, _078076_, _078077_, _078078_, _078079_, _078080_, _078081_, _078082_, _078083_, _078084_, _078085_, _078086_, _078087_, _078088_, _078089_, _078090_, _078091_, _078092_, _078093_, _078094_, _078095_, _078096_, _078097_, _078098_, _078099_, _078100_, _078101_, _078102_, _078103_, _078104_, _078105_, _078106_, _078107_, _078108_, _078109_, _078110_, _078111_, _078112_, _078113_, _078114_, _078115_, _078116_, _078117_, _078118_, _078119_, _078120_, _078121_, _078122_, _078123_, _078124_, _078125_, _078126_, _078127_, _078128_, _078129_, _078130_, _078131_, _078132_, _078133_, _078134_, _078135_, _078136_, _078137_, _078138_, _078139_, _078140_, _078141_, _078142_, _078143_, _078144_, _078145_, _078146_, _078147_, _078148_, _078149_, _078150_, _078151_, _078152_, _078153_, _078154_, _078155_, _078156_, _078157_, _078158_, _078159_, _078160_, _078161_, _078162_, _078163_, _078164_, _078165_, _078166_, _078167_, _078168_, _078169_, _078170_, _078171_, _078172_, _078173_, _078174_, _078175_, _078176_, _078177_, _078178_, _078179_, _078180_, _078181_, _078182_, _078183_, _078184_, _078185_, _078186_, _078187_, _078188_, _078189_, _078190_, _078191_, _078192_, _078193_, _078194_, _078195_, _078196_, _078197_, _078198_, _078199_, _078200_, _078201_, _078202_, _078203_, _078204_, _078205_, _078206_, _078207_, _078208_, _078209_, _078210_, _078211_, _078212_, _078213_, _078214_, _078215_, _078216_, _078217_, _078218_, _078219_, _078220_, _078221_, _078222_, _078223_, _078224_, _078225_, _078226_, _078227_, _078228_, _078229_, _078230_, _078231_, _078232_, _078233_, _078234_, _078235_, _078236_, _078237_, _078238_, _078239_, _078240_, _078241_, _078242_, _078243_, _078244_, _078245_, _078246_, _078247_, _078248_, _078249_, _078250_, _078251_, _078252_, _078253_, _078254_, _078255_, _078256_, _078257_, _078258_, _078259_, _078260_, _078261_, _078262_, _078263_, _078264_, _078265_, _078266_, _078267_, _078268_, _078269_, _078270_, _078271_, _078272_, _078273_, _078274_, _078275_, _078276_, _078277_, _078278_, _078279_, _078280_, _078281_, _078282_, _078283_, _078284_, _078285_, _078286_, _078287_, _078288_, _078289_, _078290_, _078291_, _078292_, _078293_, _078294_, _078295_, _078296_, _078297_, _078298_, _078299_, _078300_, _078301_, _078302_, _078303_, _078304_, _078305_, _078306_, _078307_, _078308_, _078309_, _078310_, _078311_, _078312_, _078313_, _078314_, _078315_, _078316_, _078317_, _078318_, _078319_, _078320_, _078321_, _078322_, _078323_, _078324_, _078325_, _078326_, _078327_, _078328_, _078329_, _078330_, _078331_, _078332_, _078333_, _078334_, _078335_, _078336_, _078337_, _078338_, _078339_, _078340_, _078341_, _078342_, _078343_, _078344_, _078345_, _078346_, _078347_, _078348_, _078349_, _078350_, _078351_, _078352_, _078353_, _078354_, _078355_, _078356_, _078357_, _078358_, _078359_, _078360_, _078361_, _078362_, _078363_, _078364_, _078365_, _078366_, _078367_, _078368_, _078369_, _078370_, _078371_, _078372_, _078373_, _078374_, _078375_, _078376_, _078377_, _078378_, _078379_, _078380_, _078381_, _078382_, _078383_, _078384_, _078385_, _078386_, _078387_, _078388_, _078389_, _078390_, _078391_, _078392_, _078393_, _078394_, _078395_, _078396_, _078397_, _078398_, _078399_, _078400_, _078401_, _078402_, _078403_, _078404_, _078405_, _078406_, _078407_, _078408_, _078409_, _078410_, _078411_, _078412_, _078413_, _078414_, _078415_, _078416_, _078417_, _078418_, _078419_, _078420_, _078421_, _078422_, _078423_, _078424_, _078425_, _078426_, _078427_, _078428_, _078429_, _078430_, _078431_, _078432_, _078433_, _078434_, _078435_, _078436_, _078437_, _078438_, _078439_, _078440_, _078441_, _078442_, _078443_, _078444_, _078445_, _078446_, _078447_, _078448_, _078449_, _078450_, _078451_, _078452_, _078453_, _078454_, _078455_, _078456_, _078457_, _078458_, _078459_, _078460_, _078461_, _078462_, _078463_, _078464_, _078465_, _078466_, _078467_, _078468_, _078469_, _078470_, _078471_, _078472_, _078473_, _078474_, _078475_, _078476_, _078477_, _078478_, _078479_, _078480_, _078481_, _078482_, _078483_, _078484_, _078485_, _078486_, _078487_, _078488_, _078489_, _078490_, _078491_, _078492_, _078493_, _078494_, _078495_, _078496_, _078497_, _078498_, _078499_, _078500_, _078501_, _078502_, _078503_, _078504_, _078505_, _078506_, _078507_, _078508_, _078509_, _078510_, _078511_, _078512_, _078513_, _078514_, _078515_, _078516_, _078517_, _078518_, _078519_, _078520_, _078521_, _078522_, _078523_, _078524_, _078525_, _078526_, _078527_, _078528_, _078529_, _078530_, _078531_, _078532_, _078533_, _078534_, _078535_, _078536_, _078537_, _078538_, _078539_, _078540_, _078541_, _078542_, _078543_, _078544_, _078545_, _078546_, _078547_, _078548_, _078549_, _078550_, _078551_, _078552_, _078553_, _078554_, _078555_, _078556_, _078557_, _078558_, _078559_, _078560_, _078561_, _078562_, _078563_, _078564_, _078565_, _078566_, _078567_, _078568_, _078569_, _078570_, _078571_, _078572_, _078573_, _078574_, _078575_, _078576_, _078577_, _078578_, _078579_, _078580_, _078581_, _078582_, _078583_, _078584_, _078585_, _078586_, _078587_, _078588_, _078589_, _078590_, _078591_, _078592_, _078593_, _078594_, _078595_, _078596_, _078597_, _078598_, _078599_, _078600_, _078601_, _078602_, _078603_, _078604_, _078605_, _078606_, _078607_, _078608_, _078609_, _078610_, _078611_, _078612_, _078613_, _078614_, _078615_, _078616_, _078617_, _078618_, _078619_, _078620_, _078621_, _078622_, _078623_, _078624_, _078625_, _078626_, _078627_, _078628_, _078629_, _078630_, _078631_, _078632_, _078633_, _078634_, _078635_, _078636_, _078637_, _078638_, _078639_, _078640_, _078641_, _078642_, _078643_, _078644_, _078645_, _078646_, _078647_, _078648_, _078649_, _078650_, _078651_, _078652_, _078653_, _078654_, _078655_, _078656_, _078657_, _078658_, _078659_, _078660_, _078661_, _078662_, _078663_, _078664_, _078665_, _078666_, _078667_, _078668_, _078669_, _078670_, _078671_, _078672_, _078673_, _078674_, _078675_, _078676_, _078677_, _078678_, _078679_, _078680_, _078681_, _078682_, _078683_, _078684_, _078685_, _078686_, _078687_, _078688_, _078689_, _078690_, _078691_, _078692_, _078693_, _078694_, _078695_, _078696_, _078697_, _078698_, _078699_, _078700_, _078701_, _078702_, _078703_, _078704_, _078705_, _078706_, _078707_, _078708_, _078709_, _078710_, _078711_, _078712_, _078713_, _078714_, _078715_, _078716_, _078717_, _078718_, _078719_, _078720_, _078721_, _078722_, _078723_, _078724_, _078725_, _078726_, _078727_, _078728_, _078729_, _078730_, _078731_, _078732_, _078733_, _078734_, _078735_, _078736_, _078737_, _078738_, _078739_, _078740_, _078741_, _078742_, _078743_, _078744_, _078745_, _078746_, _078747_, _078748_, _078749_, _078750_, _078751_, _078752_, _078753_, _078754_, _078755_, _078756_, _078757_, _078758_, _078759_, _078760_, _078761_, _078762_, _078763_, _078764_, _078765_, _078766_, _078767_, _078768_, _078769_, _078770_, _078771_, _078772_, _078773_, _078774_, _078775_, _078776_, _078777_, _078778_, _078779_, _078780_, _078781_, _078782_, _078783_, _078784_, _078785_, _078786_, _078787_, _078788_, _078789_, _078790_, _078791_, _078792_, _078793_, _078794_, _078795_, _078796_, _078797_, _078798_, _078799_, _078800_, _078801_, _078802_, _078803_, _078804_, _078805_, _078806_, _078807_, _078808_, _078809_, _078810_, _078811_, _078812_, _078813_, _078814_, _078815_, _078816_, _078817_, _078818_, _078819_, _078820_, _078821_, _078822_, _078823_, _078824_, _078825_, _078826_, _078827_, _078828_, _078829_, _078830_, _078831_, _078832_, _078833_, _078834_, _078835_, _078836_, _078837_, _078838_, _078839_, _078840_, _078841_, _078842_, _078843_, _078844_, _078845_, _078846_, _078847_, _078848_, _078849_, _078850_, _078851_, _078852_, _078853_, _078854_, _078855_, _078856_, _078857_, _078858_, _078859_, _078860_, _078861_, _078862_, _078863_, _078864_, _078865_, _078866_, _078867_, _078868_, _078869_, _078870_, _078871_, _078872_, _078873_, _078874_, _078875_, _078876_, _078877_, _078878_, _078879_, _078880_, _078881_, _078882_, _078883_, _078884_, _078885_, _078886_, _078887_, _078888_, _078889_, _078890_, _078891_, _078892_, _078893_, _078894_, _078895_, _078896_, _078897_, _078898_, _078899_, _078900_, _078901_, _078902_, _078903_, _078904_, _078905_, _078906_, _078907_, _078908_, _078909_, _078910_, _078911_, _078912_, _078913_, _078914_, _078915_, _078916_, _078917_, _078918_, _078919_, _078920_, _078921_, _078922_, _078923_, _078924_, _078925_, _078926_, _078927_, _078928_, _078929_, _078930_, _078931_, _078932_, _078933_, _078934_, _078935_, _078936_, _078937_, _078938_, _078939_, _078940_, _078941_, _078942_, _078943_, _078944_, _078945_, _078946_, _078947_, _078948_, _078949_, _078950_, _078951_, _078952_, _078953_, _078954_, _078955_, _078956_, _078957_, _078958_, _078959_, _078960_, _078961_, _078962_, _078963_, _078964_, _078965_, _078966_, _078967_, _078968_, _078969_, _078970_, _078971_, _078972_, _078973_, _078974_, _078975_, _078976_, _078977_, _078978_, _078979_, _078980_, _078981_, _078982_, _078983_, _078984_, _078985_, _078986_, _078987_, _078988_, _078989_, _078990_, _078991_, _078992_, _078993_, _078994_, _078995_, _078996_, _078997_, _078998_, _078999_, _079000_, _079001_, _079002_, _079003_, _079004_, _079005_, _079006_, _079007_, _079008_, _079009_, _079010_, _079011_, _079012_, _079013_, _079014_, _079015_, _079016_, _079017_, _079018_, _079019_, _079020_, _079021_, _079022_, _079023_, _079024_, _079025_, _079026_, _079027_, _079028_, _079029_, _079030_, _079031_, _079032_, _079033_, _079034_, _079035_, _079036_, _079037_, _079038_, _079039_, _079040_, _079041_, _079042_, _079043_, _079044_, _079045_, _079046_, _079047_, _079048_, _079049_, _079050_, _079051_, _079052_, _079053_, _079054_, _079055_, _079056_, _079057_, _079058_, _079059_, _079060_, _079061_, _079062_, _079063_, _079064_, _079065_, _079066_, _079067_, _079068_, _079069_, _079070_, _079071_, _079072_, _079073_, _079074_, _079075_, _079076_, _079077_, _079078_, _079079_, _079080_, _079081_, _079082_, _079083_, _079084_, _079085_, _079086_, _079087_, _079088_, _079089_, _079090_, _079091_, _079092_, _079093_, _079094_, _079095_, _079096_, _079097_, _079098_, _079099_, _079100_, _079101_, _079102_, _079103_, _079104_, _079105_, _079106_, _079107_, _079108_, _079109_, _079110_, _079111_, _079112_, _079113_, _079114_, _079115_, _079116_, _079117_, _079118_, _079119_, _079120_, _079121_, _079122_, _079123_, _079124_, _079125_, _079126_, _079127_, _079128_, _079129_, _079130_, _079131_, _079132_, _079133_, _079134_, _079135_, _079136_, _079137_, _079138_, _079139_, _079140_, _079141_, _079142_, _079143_, _079144_, _079145_, _079146_, _079147_, _079148_, _079149_, _079150_, _079151_, _079152_, _079153_, _079154_, _079155_, _079156_, _079157_, _079158_, _079159_, _079160_, _079161_, _079162_, _079163_, _079164_, _079165_, _079166_, _079167_, _079168_, _079169_, _079170_, _079171_, _079172_, _079173_, _079174_, _079175_, _079176_, _079177_, _079178_, _079179_, _079180_, _079181_, _079182_, _079183_, _079184_, _079185_, _079186_, _079187_, _079188_, _079189_, _079190_, _079191_, _079192_, _079193_, _079194_, _079195_, _079196_, _079197_, _079198_, _079199_, _079200_, _079201_, _079202_, _079203_, _079204_, _079205_, _079206_, _079207_, _079208_, _079209_, _079210_, _079211_, _079212_, _079213_, _079214_, _079215_, _079216_, _079217_, _079218_, _079219_, _079220_, _079221_, _079222_, _079223_, _079224_, _079225_, _079226_, _079227_, _079228_, _079229_, _079230_, _079231_, _079232_, _079233_, _079234_, _079235_, _079236_, _079237_, _079238_, _079239_, _079240_, _079241_, _079242_, _079243_, _079244_, _079245_, _079246_, _079247_, _079248_, _079249_, _079250_, _079251_, _079252_, _079253_, _079254_, _079255_, _079256_, _079257_, _079258_, _079259_, _079260_, _079261_, _079262_, _079263_, _079264_, _079265_, _079266_, _079267_, _079268_, _079269_, _079270_, _079271_, _079272_, _079273_, _079274_, _079275_, _079276_, _079277_, _079278_, _079279_, _079280_, _079281_, _079282_, _079283_, _079284_, _079285_, _079286_, _079287_, _079288_, _079289_, _079290_, _079291_, _079292_, _079293_, _079294_, _079295_, _079296_, _079297_, _079298_, _079299_, _079300_, _079301_, _079302_, _079303_, _079304_, _079305_, _079306_, _079307_, _079308_, _079309_, _079310_, _079311_, _079312_, _079313_, _079314_, _079315_, _079316_, _079317_, _079318_, _079319_, _079320_, _079321_, _079322_, _079323_, _079324_, _079325_, _079326_, _079327_, _079328_, _079329_, _079330_, _079331_, _079332_, _079333_, _079334_, _079335_, _079336_, _079337_, _079338_, _079339_, _079340_, _079341_, _079342_, _079343_, _079344_, _079345_, _079346_, _079347_, _079348_, _079349_, _079350_, _079351_, _079352_, _079353_, _079354_, _079355_, _079356_, _079357_, _079358_, _079359_, _079360_, _079361_, _079362_, _079363_, _079364_, _079365_, _079366_, _079367_, _079368_, _079369_, _079370_, _079371_, _079372_, _079373_, _079374_, _079375_, _079376_, _079377_, _079378_, _079379_, _079380_, _079381_, _079382_, _079383_, _079384_, _079385_, _079386_, _079387_, _079388_, _079389_, _079390_, _079391_, _079392_, _079393_, _079394_, _079395_, _079396_, _079397_, _079398_, _079399_, _079400_, _079401_, _079402_, _079403_, _079404_, _079405_, _079406_, _079407_, _079408_, _079409_, _079410_, _079411_, _079412_, _079413_, _079414_, _079415_, _079416_, _079417_, _079418_, _079419_, _079420_, _079421_, _079422_, _079423_, _079424_, _079425_, _079426_, _079427_, _079428_, _079429_, _079430_, _079431_, _079432_, _079433_, _079434_, _079435_, _079436_, _079437_, _079438_, _079439_, _079440_, _079441_, _079442_, _079443_, _079444_, _079445_, _079446_, _079447_, _079448_, _079449_, _079450_, _079451_, _079452_, _079453_, _079454_, _079455_, _079456_, _079457_, _079458_, _079459_, _079460_, _079461_, _079462_, _079463_, _079464_, _079465_, _079466_, _079467_, _079468_, _079469_, _079470_, _079471_, _079472_, _079473_, _079474_, _079475_, _079476_, _079477_, _079478_, _079479_, _079480_, _079481_, _079482_, _079483_, _079484_, _079485_, _079486_, _079487_, _079488_, _079489_, _079490_, _079491_, _079492_, _079493_, _079494_, _079495_, _079496_, _079497_, _079498_, _079499_, _079500_, _079501_, _079502_, _079503_, _079504_, _079505_, _079506_, _079507_, _079508_, _079509_, _079510_, _079511_, _079512_, _079513_, _079514_, _079515_, _079516_, _079517_, _079518_, _079519_, _079520_, _079521_, _079522_, _079523_, _079524_, _079525_, _079526_, _079527_, _079528_, _079529_, _079530_, _079531_, _079532_, _079533_, _079534_, _079535_, _079536_, _079537_, _079538_, _079539_, _079540_, _079541_, _079542_, _079543_, _079544_, _079545_, _079546_, _079547_, _079548_, _079549_, _079550_, _079551_, _079552_, _079553_, _079554_, _079555_, _079556_, _079557_, _079558_, _079559_, _079560_, _079561_, _079562_, _079563_, _079564_, _079565_, _079566_, _079567_, _079568_, _079569_, _079570_, _079571_, _079572_, _079573_, _079574_, _079575_, _079576_, _079577_, _079578_, _079579_, _079580_, _079581_, _079582_, _079583_, _079584_, _079585_, _079586_, _079587_, _079588_, _079589_, _079590_, _079591_, _079592_, _079593_, _079594_, _079595_, _079596_, _079597_, _079598_, _079599_, _079600_, _079601_, _079602_, _079603_, _079604_, _079605_, _079606_, _079607_, _079608_, _079609_, _079610_, _079611_, _079612_, _079613_, _079614_, _079615_, _079616_, _079617_, _079618_, _079619_, _079620_, _079621_, _079622_, _079623_, _079624_, _079625_, _079626_, _079627_, _079628_, _079629_, _079630_, _079631_, _079632_, _079633_, _079634_, _079635_, _079636_, _079637_, _079638_, _079639_, _079640_, _079641_, _079642_, _079643_, _079644_, _079645_, _079646_, _079647_, _079648_, _079649_, _079650_, _079651_, _079652_, _079653_, _079654_, _079655_, _079656_, _079657_, _079658_, _079659_, _079660_, _079661_, _079662_, _079663_, _079664_, _079665_, _079666_, _079667_, _079668_, _079669_, _079670_, _079671_, _079672_, _079673_, _079674_, _079675_, _079676_, _079677_, _079678_, _079679_, _079680_, _079681_, _079682_, _079683_, _079684_, _079685_, _079686_, _079687_, _079688_, _079689_, _079690_, _079691_, _079692_, _079693_, _079694_, _079695_, _079696_, _079697_, _079698_, _079699_, _079700_, _079701_, _079702_, _079703_, _079704_, _079705_, _079706_, _079707_, _079708_, _079709_, _079710_, _079711_, _079712_, _079713_, _079714_, _079715_, _079716_, _079717_, _079718_, _079719_, _079720_, _079721_, _079722_, _079723_, _079724_, _079725_, _079726_, _079727_, _079728_, _079729_, _079730_, _079731_, _079732_, _079733_, _079734_, _079735_, _079736_, _079737_, _079738_, _079739_, _079740_, _079741_, _079742_, _079743_, _079744_, _079745_, _079746_, _079747_, _079748_, _079749_, _079750_, _079751_, _079752_, _079753_, _079754_, _079755_, _079756_, _079757_, _079758_, _079759_, _079760_, _079761_, _079762_, _079763_, _079764_, _079765_, _079766_, _079767_, _079768_, _079769_, _079770_, _079771_, _079772_, _079773_, _079774_, _079775_, _079776_, _079777_, _079778_, _079779_, _079780_, _079781_, _079782_, _079783_, _079784_, _079785_, _079786_, _079787_, _079788_, _079789_, _079790_, _079791_, _079792_, _079793_, _079794_, _079795_, _079796_, _079797_, _079798_, _079799_, _079800_, _079801_, _079802_, _079803_, _079804_, _079805_, _079806_, _079807_, _079808_, _079809_, _079810_, _079811_, _079812_, _079813_, _079814_, _079815_, _079816_, _079817_, _079818_, _079819_, _079820_, _079821_, _079822_, _079823_, _079824_, _079825_, _079826_, _079827_, _079828_, _079829_, _079830_, _079831_, _079832_, _079833_, _079834_, _079835_, _079836_, _079837_, _079838_, _079839_, _079840_, _079841_, _079842_, _079843_, _079844_, _079845_, _079846_, _079847_, _079848_, _079849_, _079850_, _079851_, _079852_, _079853_, _079854_, _079855_, _079856_, _079857_, _079858_, _079859_, _079860_, _079861_, _079862_, _079863_, _079864_, _079865_, _079866_, _079867_, _079868_, _079869_, _079870_, _079871_, _079872_, _079873_, _079874_, _079875_, _079876_, _079877_, _079878_, _079879_, _079880_, _079881_, _079882_, _079883_, _079884_, _079885_, _079886_, _079887_, _079888_, _079889_, _079890_, _079891_, _079892_, _079893_, _079894_, _079895_, _079896_, _079897_, _079898_, _079899_, _079900_, _079901_, _079902_, _079903_, _079904_, _079905_, _079906_, _079907_, _079908_, _079909_, _079910_, _079911_, _079912_, _079913_, _079914_, _079915_, _079916_, _079917_, _079918_, _079919_, _079920_, _079921_, _079922_, _079923_, _079924_, _079925_, _079926_, _079927_, _079928_, _079929_, _079930_, _079931_, _079932_, _079933_, _079934_, _079935_, _079936_, _079937_, _079938_, _079939_, _079940_, _079941_, _079942_, _079943_, _079944_, _079945_, _079946_, _079947_, _079948_, _079949_, _079950_, _079951_, _079952_, _079953_, _079954_, _079955_, _079956_, _079957_, _079958_, _079959_, _079960_, _079961_, _079962_, _079963_, _079964_, _079965_, _079966_, _079967_, _079968_, _079969_, _079970_, _079971_, _079972_, _079973_, _079974_, _079975_, _079976_, _079977_, _079978_, _079979_, _079980_, _079981_, _079982_, _079983_, _079984_, _079985_, _079986_, _079987_, _079988_, _079989_, _079990_, _079991_, _079992_, _079993_, _079994_, _079995_, _079996_, _079997_, _079998_, _079999_, _080000_, _080001_, _080002_, _080003_, _080004_, _080005_, _080006_, _080007_, _080008_, _080009_, _080010_, _080011_, _080012_, _080013_, _080014_, _080015_, _080016_, _080017_, _080018_, _080019_, _080020_, _080021_, _080022_, _080023_, _080024_, _080025_, _080026_, _080027_, _080028_, _080029_, _080030_, _080031_, _080032_, _080033_, _080034_, _080035_, _080036_, _080037_, _080038_, _080039_, _080040_, _080041_, _080042_, _080043_, _080044_, _080045_, _080046_, _080047_, _080048_, _080049_, _080050_, _080051_, _080052_, _080053_, _080054_, _080055_, _080056_, _080057_, _080058_, _080059_, _080060_, _080061_, _080062_, _080063_, _080064_, _080065_, _080066_, _080067_, _080068_, _080069_, _080070_, _080071_, _080072_, _080073_, _080074_, _080075_, _080076_, _080077_, _080078_, _080079_, _080080_, _080081_, _080082_, _080083_, _080084_, _080085_, _080086_, _080087_, _080088_, _080089_, _080090_, _080091_, _080092_, _080093_, _080094_, _080095_, _080096_, _080097_, _080098_, _080099_, _080100_, _080101_, _080102_, _080103_, _080104_, _080105_, _080106_, _080107_, _080108_, _080109_, _080110_, _080111_, _080112_, _080113_, _080114_, _080115_, _080116_, _080117_, _080118_, _080119_, _080120_, _080121_, _080122_, _080123_, _080124_, _080125_, _080126_, _080127_, _080128_, _080129_, _080130_, _080131_, _080132_, _080133_, _080134_, _080135_, _080136_, _080137_, _080138_, _080139_, _080140_, _080141_, _080142_, _080143_, _080144_, _080145_, _080146_, _080147_, _080148_, _080149_, _080150_, _080151_, _080152_, _080153_, _080154_, _080155_, _080156_, _080157_, _080158_, _080159_, _080160_, _080161_, _080162_, _080163_, _080164_, _080165_, _080166_, _080167_, _080168_, _080169_, _080170_, _080171_, _080172_, _080173_, _080174_, _080175_, _080176_, _080177_, _080178_, _080179_, _080180_, _080181_, _080182_, _080183_, _080184_, _080185_, _080186_, _080187_, _080188_, _080189_, _080190_, _080191_, _080192_, _080193_, _080194_, _080195_, _080196_, _080197_, _080198_, _080199_, _080200_, _080201_, _080202_, _080203_, _080204_, _080205_, _080206_, _080207_, _080208_, _080209_, _080210_, _080211_, _080212_, _080213_, _080214_, _080215_, _080216_, _080217_, _080218_, _080219_, _080220_, _080221_, _080222_, _080223_, _080224_, _080225_, _080226_, _080227_, _080228_, _080229_, _080230_, _080231_, _080232_, _080233_, _080234_, _080235_, _080236_, _080237_, _080238_, _080239_, _080240_, _080241_, _080242_, _080243_, _080244_, _080245_, _080246_, _080247_, _080248_, _080249_, _080250_, _080251_, _080252_, _080253_, _080254_, _080255_, _080256_, _080257_, _080258_, _080259_, _080260_, _080261_, _080262_, _080263_, _080264_, _080265_, _080266_, _080267_, _080268_, _080269_, _080270_, _080271_, _080272_, _080273_, _080274_, _080275_, _080276_, _080277_, _080278_, _080279_, _080280_, _080281_, _080282_, _080283_, _080284_, _080285_, _080286_, _080287_, _080288_, _080289_, _080290_, _080291_, _080292_, _080293_, _080294_, _080295_, _080296_, _080297_, _080298_, _080299_, _080300_, _080301_, _080302_, _080303_, _080304_, _080305_, _080306_, _080307_, _080308_, _080309_, _080310_, _080311_, _080312_, _080313_, _080314_, _080315_, _080316_, _080317_, _080318_, _080319_, _080320_, _080321_, _080322_, _080323_, _080324_, _080325_, _080326_, _080327_, _080328_, _080329_, _080330_, _080331_, _080332_, _080333_, _080334_, _080335_, _080336_, _080337_, _080338_, _080339_, _080340_, _080341_, _080342_, _080343_, _080344_, _080345_, _080346_, _080347_, _080348_, _080349_, _080350_, _080351_, _080352_, _080353_, _080354_, _080355_, _080356_, _080357_, _080358_, _080359_, _080360_, _080361_, _080362_, _080363_, _080364_, _080365_, _080366_, _080367_, _080368_, _080369_, _080370_, _080371_, _080372_, _080373_, _080374_, _080375_, _080376_, _080377_, _080378_, _080379_, _080380_, _080381_, _080382_, _080383_, _080384_, _080385_, _080386_, _080387_, _080388_, _080389_, _080390_, _080391_, _080392_, _080393_, _080394_, _080395_, _080396_, _080397_, _080398_, _080399_, _080400_, _080401_, _080402_, _080403_, _080404_, _080405_, _080406_, _080407_, _080408_, _080409_, _080410_, _080411_, _080412_, _080413_, _080414_, _080415_, _080416_, _080417_, _080418_, _080419_, _080420_, _080421_, _080422_, _080423_, _080424_, _080425_, _080426_, _080427_, _080428_, _080429_, _080430_, _080431_, _080432_, _080433_, _080434_, _080435_, _080436_, _080437_, _080438_, _080439_, _080440_, _080441_, _080442_, _080443_, _080444_, _080445_, _080446_, _080447_, _080448_, _080449_, _080450_, _080451_, _080452_, _080453_, _080454_, _080455_, _080456_, _080457_, _080458_, _080459_, _080460_, _080461_, _080462_, _080463_, _080464_, _080465_, _080466_, _080467_, _080468_, _080469_, _080470_, _080471_, _080472_, _080473_, _080474_, _080475_, _080476_, _080477_, _080478_, _080479_, _080480_, _080481_, _080482_, _080483_, _080484_, _080485_, _080486_, _080487_, _080488_, _080489_, _080490_, _080491_, _080492_, _080493_, _080494_, _080495_, _080496_, _080497_, _080498_, _080499_, _080500_, _080501_, _080502_, _080503_, _080504_, _080505_, _080506_, _080507_, _080508_, _080509_, _080510_, _080511_, _080512_, _080513_, _080514_, _080515_, _080516_, _080517_, _080518_, _080519_, _080520_, _080521_, _080522_, _080523_, _080524_, _080525_, _080526_, _080527_, _080528_, _080529_, _080530_, _080531_, _080532_, _080533_, _080534_, _080535_, _080536_, _080537_, _080538_, _080539_, _080540_, _080541_, _080542_, _080543_, _080544_, _080545_, _080546_, _080547_, _080548_, _080549_, _080550_, _080551_, _080552_, _080553_, _080554_, _080555_, _080556_, _080557_, _080558_, _080559_, _080560_, _080561_, _080562_, _080563_, _080564_, _080565_, _080566_, _080567_, _080568_, _080569_, _080570_, _080571_, _080572_, _080573_, _080574_, _080575_, _080576_, _080577_, _080578_, _080579_, _080580_, _080581_, _080582_, _080583_, _080584_, _080585_, _080586_, _080587_, _080588_, _080589_, _080590_, _080591_, _080592_, _080593_, _080594_, _080595_, _080596_, _080597_, _080598_, _080599_, _080600_, _080601_, _080602_, _080603_, _080604_, _080605_, _080606_, _080607_, _080608_, _080609_, _080610_, _080611_, _080612_, _080613_, _080614_, _080615_, _080616_, _080617_, _080618_, _080619_, _080620_, _080621_, _080622_, _080623_, _080624_, _080625_, _080626_, _080627_, _080628_, _080629_, _080630_, _080631_, _080632_, _080633_, _080634_, _080635_, _080636_, _080637_, _080638_, _080639_, _080640_, _080641_, _080642_, _080643_, _080644_, _080645_, _080646_, _080647_, _080648_, _080649_, _080650_, _080651_, _080652_, _080653_, _080654_, _080655_, _080656_, _080657_, _080658_, _080659_, _080660_, _080661_, _080662_, _080663_, _080664_, _080665_, _080666_, _080667_, _080668_, _080669_, _080670_, _080671_, _080672_, _080673_, _080674_, _080675_, _080676_, _080677_, _080678_, _080679_, _080680_, _080681_, _080682_, _080683_, _080684_, _080685_, _080686_, _080687_, _080688_, _080689_, _080690_, _080691_, _080692_, _080693_, _080694_, _080695_, _080696_, _080697_, _080698_, _080699_, _080700_, _080701_, _080702_, _080703_, _080704_, _080705_, _080706_, _080707_, _080708_, _080709_, _080710_, _080711_, _080712_, _080713_, _080714_, _080715_, _080716_, _080717_, _080718_, _080719_, _080720_, _080721_, _080722_, _080723_, _080724_, _080725_, _080726_, _080727_, _080728_, _080729_, _080730_, _080731_, _080732_, _080733_, _080734_, _080735_, _080736_, _080737_, _080738_, _080739_, _080740_, _080741_, _080742_, _080743_, _080744_, _080745_, _080746_, _080747_, _080748_, _080749_, _080750_, _080751_, _080752_, _080753_, _080754_, _080755_, _080756_, _080757_, _080758_, _080759_, _080760_, _080761_, _080762_, _080763_, _080764_, _080765_, _080766_, _080767_, _080768_, _080769_, _080770_, _080771_, _080772_, _080773_, _080774_, _080775_, _080776_, _080777_, _080778_, _080779_, _080780_, _080781_, _080782_, _080783_, _080784_, _080785_, _080786_, _080787_, _080788_, _080789_, _080790_, _080791_, _080792_, _080793_, _080794_, _080795_, _080796_, _080797_, _080798_, _080799_, _080800_, _080801_, _080802_, _080803_, _080804_, _080805_, _080806_, _080807_, _080808_, _080809_, _080810_, _080811_, _080812_, _080813_, _080814_, _080815_, _080816_, _080817_, _080818_, _080819_, _080820_, _080821_, _080822_, _080823_, _080824_, _080825_, _080826_, _080827_, _080828_, _080829_, _080830_, _080831_, _080832_, _080833_, _080834_, _080835_, _080836_, _080837_, _080838_, _080839_, _080840_, _080841_, _080842_, _080843_, _080844_, _080845_, _080846_, _080847_, _080848_, _080849_, _080850_, _080851_, _080852_, _080853_, _080854_, _080855_, _080856_, _080857_, _080858_, _080859_, _080860_, _080861_, _080862_, _080863_, _080864_, _080865_, _080866_, _080867_, _080868_, _080869_, _080870_, _080871_, _080872_, _080873_, _080874_, _080875_, _080876_, _080877_, _080878_, _080879_, _080880_, _080881_, _080882_, _080883_, _080884_, _080885_, _080886_, _080887_, _080888_, _080889_, _080890_, _080891_, _080892_, _080893_, _080894_, _080895_, _080896_, _080897_, _080898_, _080899_, _080900_, _080901_, _080902_, _080903_, _080904_, _080905_, _080906_, _080907_, _080908_, _080909_, _080910_, _080911_, _080912_, _080913_, _080914_, _080915_, _080916_, _080917_, _080918_, _080919_, _080920_, _080921_, _080922_, _080923_, _080924_, _080925_, _080926_, _080927_, _080928_, _080929_, _080930_, _080931_, _080932_, _080933_, _080934_, _080935_, _080936_, _080937_, _080938_, _080939_, _080940_, _080941_, _080942_, _080943_, _080944_, _080945_, _080946_, _080947_, _080948_, _080949_, _080950_, _080951_, _080952_, _080953_, _080954_, _080955_, _080956_, _080957_, _080958_, _080959_, _080960_, _080961_, _080962_, _080963_, _080964_, _080965_, _080966_, _080967_, _080968_, _080969_, _080970_, _080971_, _080972_, _080973_, _080974_, _080975_, _080976_, _080977_, _080978_, _080979_, _080980_, _080981_, _080982_, _080983_, _080984_, _080985_, _080986_, _080987_, _080988_, _080989_, _080990_, _080991_, _080992_, _080993_, _080994_, _080995_, _080996_, _080997_, _080998_, _080999_, _081000_, _081001_, _081002_, _081003_, _081004_, _081005_, _081006_, _081007_, _081008_, _081009_, _081010_, _081011_, _081012_, _081013_, _081014_, _081015_, _081016_, _081017_, _081018_, _081019_, _081020_, _081021_, _081022_, _081023_, _081024_, _081025_, _081026_, _081027_, _081028_, _081029_, _081030_, _081031_, _081032_, _081033_, _081034_, _081035_, _081036_, _081037_, _081038_, _081039_, _081040_, _081041_, _081042_, _081043_, _081044_, _081045_, _081046_, _081047_, _081048_, _081049_, _081050_, _081051_, _081052_, _081053_, _081054_, _081055_, _081056_, _081057_, _081058_, _081059_, _081060_, _081061_, _081062_, _081063_, _081064_, _081065_, _081066_, _081067_, _081068_, _081069_, _081070_, _081071_, _081072_, _081073_, _081074_, _081075_, _081076_, _081077_, _081078_, _081079_, _081080_, _081081_, _081082_, _081083_, _081084_, _081085_, _081086_, _081087_, _081088_, _081089_, _081090_, _081091_, _081092_, _081093_, _081094_, _081095_, _081096_, _081097_, _081098_, _081099_, _081100_, _081101_, _081102_, _081103_, _081104_, _081105_, _081106_, _081107_, _081108_, _081109_, _081110_, _081111_, _081112_, _081113_, _081114_, _081115_, _081116_, _081117_, _081118_, _081119_, _081120_, _081121_, _081122_, _081123_, _081124_, _081125_, _081126_, _081127_, _081128_, _081129_, _081130_, _081131_, _081132_, _081133_, _081134_, _081135_, _081136_, _081137_, _081138_, _081139_, _081140_, _081141_, _081142_, _081143_, _081144_, _081145_, _081146_, _081147_, _081148_, _081149_, _081150_, _081151_, _081152_, _081153_, _081154_, _081155_, _081156_, _081157_, _081158_, _081159_, _081160_, _081161_, _081162_, _081163_, _081164_, _081165_, _081166_, _081167_, _081168_, _081169_, _081170_, _081171_, _081172_, _081173_, _081174_, _081175_, _081176_, _081177_, _081178_, _081179_, _081180_, _081181_, _081182_, _081183_, _081184_, _081185_, _081186_, _081187_, _081188_, _081189_, _081190_, _081191_, _081192_, _081193_, _081194_, _081195_, _081196_, _081197_, _081198_, _081199_, _081200_, _081201_, _081202_, _081203_, _081204_, _081205_, _081206_, _081207_, _081208_, _081209_, _081210_, _081211_, _081212_, _081213_, _081214_, _081215_, _081216_, _081217_, _081218_, _081219_, _081220_, _081221_, _081222_, _081223_, _081224_, _081225_, _081226_, _081227_, _081228_, _081229_, _081230_, _081231_, _081232_, _081233_, _081234_, _081235_, _081236_, _081237_, _081238_, _081239_, _081240_, _081241_, _081242_, _081243_, _081244_, _081245_, _081246_, _081247_, _081248_, _081249_, _081250_, _081251_, _081252_, _081253_, _081254_, _081255_, _081256_, _081257_, _081258_, _081259_, _081260_, _081261_, _081262_, _081263_, _081264_, _081265_, _081266_, _081267_, _081268_, _081269_, _081270_, _081271_, _081272_, _081273_, _081274_, _081275_, _081276_, _081277_, _081278_, _081279_, _081280_, _081281_, _081282_, _081283_, _081284_, _081285_, _081286_, _081287_, _081288_, _081289_, _081290_, _081291_, _081292_, _081293_, _081294_, _081295_, _081296_, _081297_, _081298_, _081299_, _081300_, _081301_, _081302_, _081303_, _081304_, _081305_, _081306_, _081307_, _081308_, _081309_, _081310_, _081311_, _081312_, _081313_, _081314_, _081315_, _081316_, _081317_, _081318_, _081319_, _081320_, _081321_, _081322_, _081323_, _081324_, _081325_, _081326_, _081327_, _081328_, _081329_, _081330_, _081331_, _081332_, _081333_, _081334_, _081335_, _081336_, _081337_, _081338_, _081339_, _081340_, _081341_, _081342_, _081343_, _081344_, _081345_, _081346_, _081347_, _081348_, _081349_, _081350_, _081351_, _081352_, _081353_, _081354_, _081355_, _081356_, _081357_, _081358_, _081359_, _081360_, _081361_, _081362_, _081363_, _081364_, _081365_, _081366_, _081367_, _081368_, _081369_, _081370_, _081371_, _081372_, _081373_, _081374_, _081375_, _081376_, _081377_, _081378_, _081379_, _081380_, _081381_, _081382_, _081383_, _081384_, _081385_, _081386_, _081387_, _081388_, _081389_, _081390_, _081391_, _081392_, _081393_, _081394_, _081395_, _081396_, _081397_, _081398_, _081399_, _081400_, _081401_, _081402_, _081403_, _081404_, _081405_, _081406_, _081407_, _081408_, _081409_, _081410_, _081411_, _081412_, _081413_, _081414_, _081415_, _081416_, _081417_, _081418_, _081419_, _081420_, _081421_, _081422_, _081423_, _081424_, _081425_, _081426_, _081427_, _081428_, _081429_, _081430_, _081431_, _081432_, _081433_, _081434_, _081435_, _081436_, _081437_, _081438_, _081439_, _081440_, _081441_, _081442_, _081443_, _081444_, _081445_, _081446_, _081447_, _081448_, _081449_, _081450_, _081451_, _081452_, _081453_, _081454_, _081455_, _081456_, _081457_, _081458_, _081459_, _081460_, _081461_, _081462_, _081463_, _081464_, _081465_, _081466_, _081467_, _081468_, _081469_, _081470_, _081471_, _081472_, _081473_, _081474_, _081475_, _081476_, _081477_, _081478_, _081479_, _081480_, _081481_, _081482_, _081483_, _081484_, _081485_, _081486_, _081487_, _081488_, _081489_, _081490_, _081491_, _081492_, _081493_, _081494_, _081495_, _081496_, _081497_, _081498_, _081499_, _081500_, _081501_, _081502_, _081503_, _081504_, _081505_, _081506_, _081507_, _081508_, _081509_, _081510_, _081511_, _081512_, _081513_, _081514_, _081515_, _081516_, _081517_, _081518_, _081519_, _081520_, _081521_, _081522_, _081523_, _081524_, _081525_, _081526_, _081527_, _081528_, _081529_, _081530_, _081531_, _081532_, _081533_, _081534_, _081535_, _081536_, _081537_, _081538_, _081539_, _081540_, _081541_, _081542_, _081543_, _081544_, _081545_, _081546_, _081547_, _081548_, _081549_, _081550_, _081551_, _081552_, _081553_, _081554_, _081555_, _081556_, _081557_, _081558_, _081559_, _081560_, _081561_, _081562_, _081563_, _081564_, _081565_, _081566_, _081567_, _081568_, _081569_, _081570_, _081571_, _081572_, _081573_, _081574_, _081575_, _081576_, _081577_, _081578_, _081579_, _081580_, _081581_, _081582_, _081583_, _081584_, _081585_, _081586_, _081587_, _081588_, _081589_, _081590_, _081591_, _081592_, _081593_, _081594_, _081595_, _081596_, _081597_, _081598_, _081599_, _081600_, _081601_, _081602_, _081603_, _081604_, _081605_, _081606_, _081607_, _081608_, _081609_, _081610_, _081611_, _081612_, _081613_, _081614_, _081615_, _081616_, _081617_, _081618_, _081619_, _081620_, _081621_, _081622_, _081623_, _081624_, _081625_, _081626_, _081627_, _081628_, _081629_, _081630_, _081631_, _081632_, _081633_, _081634_, _081635_, _081636_, _081637_, _081638_, _081639_, _081640_, _081641_, _081642_, _081643_, _081644_, _081645_, _081646_, _081647_, _081648_, _081649_, _081650_, _081651_, _081652_, _081653_, _081654_, _081655_, _081656_, _081657_, _081658_, _081659_, _081660_, _081661_, _081662_, _081663_, _081664_, _081665_, _081666_, _081667_, _081668_, _081669_, _081670_, _081671_, _081672_, _081673_, _081674_, _081675_, _081676_, _081677_, _081678_, _081679_, _081680_, _081681_, _081682_, _081683_, _081684_, _081685_, _081686_, _081687_, _081688_, _081689_, _081690_, _081691_, _081692_, _081693_, _081694_, _081695_, _081696_, _081697_, _081698_, _081699_, _081700_, _081701_, _081702_, _081703_, _081704_, _081705_, _081706_, _081707_, _081708_, _081709_, _081710_, _081711_, _081712_, _081713_, _081714_, _081715_, _081716_, _081717_, _081718_, _081719_, _081720_, _081721_, _081722_, _081723_, _081724_, _081725_, _081726_, _081727_, _081728_, _081729_, _081730_, _081731_, _081732_, _081733_, _081734_, _081735_, _081736_, _081737_, _081738_, _081739_, _081740_, _081741_, _081742_, _081743_, _081744_, _081745_, _081746_, _081747_, _081748_, _081749_, _081750_, _081751_, _081752_, _081753_, _081754_, _081755_, _081756_, _081757_, _081758_, _081759_, _081760_, _081761_, _081762_, _081763_, _081764_, _081765_, _081766_, _081767_, _081768_, _081769_, _081770_, _081771_, _081772_, _081773_, _081774_, _081775_, _081776_, _081777_, _081778_, _081779_, _081780_, _081781_, _081782_, _081783_, _081784_, _081785_, _081786_, _081787_, _081788_, _081789_, _081790_, _081791_, _081792_, _081793_, _081794_, _081795_, _081796_, _081797_, _081798_, _081799_, _081800_, _081801_, _081802_, _081803_, _081804_, _081805_, _081806_, _081807_, _081808_, _081809_, _081810_, _081811_, _081812_, _081813_, _081814_, _081815_, _081816_, _081817_, _081818_, _081819_, _081820_, _081821_, _081822_, _081823_, _081824_, _081825_, _081826_, _081827_, _081828_, _081829_, _081830_, _081831_, _081832_, _081833_, _081834_, _081835_, _081836_, _081837_, _081838_, _081839_, _081840_, _081841_, _081842_, _081843_, _081844_, _081845_, _081846_, _081847_, _081848_, _081849_, _081850_, _081851_, _081852_, _081853_, _081854_, _081855_, _081856_, _081857_, _081858_, _081859_, _081860_, _081861_, _081862_, _081863_, _081864_, _081865_, _081866_, _081867_, _081868_, _081869_, _081870_, _081871_, _081872_, _081873_, _081874_, _081875_, _081876_, _081877_, _081878_, _081879_, _081880_, _081881_, _081882_, _081883_, _081884_, _081885_, _081886_, _081887_, _081888_, _081889_, _081890_, _081891_, _081892_, _081893_, _081894_, _081895_, _081896_, _081897_, _081898_, _081899_, _081900_, _081901_, _081902_, _081903_, _081904_, _081905_, _081906_, _081907_, _081908_, _081909_, _081910_, _081911_, _081912_, _081913_, _081914_, _081915_, _081916_, _081917_, _081918_, _081919_, _081920_, _081921_, _081922_, _081923_, _081924_, _081925_, _081926_, _081927_, _081928_, _081929_, _081930_, _081931_, _081932_, _081933_, _081934_, _081935_, _081936_, _081937_, _081938_, _081939_, _081940_, _081941_, _081942_, _081943_, _081944_, _081945_, _081946_, _081947_, _081948_, _081949_, _081950_, _081951_, _081952_, _081953_, _081954_, _081955_, _081956_, _081957_, _081958_, _081959_, _081960_, _081961_, _081962_, _081963_, _081964_, _081965_, _081966_, _081967_, _081968_, _081969_, _081970_, _081971_, _081972_, _081973_, _081974_, _081975_, _081976_, _081977_, _081978_, _081979_, _081980_, _081981_, _081982_, _081983_, _081984_, _081985_, _081986_, _081987_, _081988_, _081989_, _081990_, _081991_, _081992_, _081993_, _081994_, _081995_, _081996_, _081997_, _081998_, _081999_, _082000_, _082001_, _082002_, _082003_, _082004_, _082005_, _082006_, _082007_, _082008_, _082009_, _082010_, _082011_, _082012_, _082013_, _082014_, _082015_, _082016_, _082017_, _082018_, _082019_, _082020_, _082021_, _082022_, _082023_, _082024_, _082025_, _082026_, _082027_, _082028_, _082029_, _082030_, _082031_, _082032_, _082033_, _082034_, _082035_, _082036_, _082037_, _082038_, _082039_, _082040_, _082041_, _082042_, _082043_, _082044_, _082045_, _082046_, _082047_, _082048_, _082049_, _082050_, _082051_, _082052_, _082053_, _082054_, _082055_, _082056_, _082057_, _082058_, _082059_, _082060_, _082061_, _082062_, _082063_, _082064_, _082065_, _082066_, _082067_, _082068_, _082069_, _082070_, _082071_, _082072_, _082073_, _082074_, _082075_, _082076_, _082077_, _082078_, _082079_, _082080_, _082081_, _082082_, _082083_, _082084_, _082085_, _082086_, _082087_, _082088_, _082089_, _082090_, _082091_, _082092_, _082093_, _082094_, _082095_, _082096_, _082097_, _082098_, _082099_, _082100_, _082101_, _082102_, _082103_, _082104_, _082105_, _082106_, _082107_, _082108_, _082109_, _082110_, _082111_, _082112_, _082113_, _082114_, _082115_, _082116_, _082117_, _082118_, _082119_, _082120_, _082121_, _082122_, _082123_, _082124_, _082125_, _082126_, _082127_, _082128_, _082129_, _082130_, _082131_, _082132_, _082133_, _082134_, _082135_, _082136_, _082137_, _082138_, _082139_, _082140_, _082141_, _082142_, _082143_, _082144_, _082145_, _082146_, _082147_, _082148_, _082149_, _082150_, _082151_, _082152_, _082153_, _082154_, _082155_, _082156_, _082157_, _082158_, _082159_, _082160_, _082161_, _082162_, _082163_, _082164_, _082165_, _082166_, _082167_, _082168_, _082169_, _082170_, _082171_, _082172_, _082173_, _082174_, _082175_, _082176_, _082177_, _082178_, _082179_, _082180_, _082181_, _082182_, _082183_, _082184_, _082185_, _082186_, _082187_, _082188_, _082189_, _082190_, _082191_, _082192_, _082193_, _082194_, _082195_, _082196_, _082197_, _082198_, _082199_, _082200_, _082201_, _082202_, _082203_, _082204_, _082205_, _082206_, _082207_, _082208_, _082209_, _082210_, _082211_, _082212_, _082213_, _082214_, _082215_, _082216_, _082217_, _082218_, _082219_, _082220_, _082221_, _082222_, _082223_, _082224_, _082225_, _082226_, _082227_, _082228_, _082229_, _082230_, _082231_, _082232_, _082233_, _082234_, _082235_, _082236_, _082237_, _082238_, _082239_, _082240_, _082241_, _082242_, _082243_, _082244_, _082245_, _082246_, _082247_, _082248_, _082249_, _082250_, _082251_, _082252_, _082253_, _082254_, _082255_, _082256_, _082257_, _082258_, _082259_, _082260_, _082261_, _082262_, _082263_, _082264_, _082265_, _082266_, _082267_, _082268_, _082269_, _082270_, _082271_, _082272_, _082273_, _082274_, _082275_, _082276_, _082277_, _082278_, _082279_, _082280_, _082281_, _082282_, _082283_, _082284_, _082285_, _082286_, _082287_, _082288_, _082289_, _082290_, _082291_, _082292_, _082293_, _082294_, _082295_, _082296_, _082297_, _082298_, _082299_, _082300_, _082301_, _082302_, _082303_, _082304_, _082305_, _082306_, _082307_, _082308_, _082309_, _082310_, _082311_, _082312_, _082313_, _082314_, _082315_, _082316_, _082317_, _082318_, _082319_, _082320_, _082321_, _082322_, _082323_, _082324_, _082325_, _082326_, _082327_, _082328_, _082329_, _082330_, _082331_, _082332_, _082333_, _082334_, _082335_, _082336_, _082337_, _082338_, _082339_, _082340_, _082341_, _082342_, _082343_, _082344_, _082345_, _082346_, _082347_, _082348_, _082349_, _082350_, _082351_, _082352_, _082353_, _082354_, _082355_, _082356_, _082357_, _082358_, _082359_, _082360_, _082361_, _082362_, _082363_, _082364_, _082365_, _082366_, _082367_, _082368_, _082369_, _082370_, _082371_, _082372_, _082373_, _082374_, _082375_, _082376_, _082377_, _082378_, _082379_, _082380_, _082381_, _082382_, _082383_, _082384_, _082385_, _082386_, _082387_, _082388_, _082389_, _082390_, _082391_, _082392_, _082393_, _082394_, _082395_, _082396_, _082397_, _082398_, _082399_, _082400_, _082401_, _082402_, _082403_, _082404_, _082405_, _082406_, _082407_, _082408_, _082409_, _082410_, _082411_, _082412_, _082413_, _082414_, _082415_, _082416_, _082417_, _082418_, _082419_, _082420_, _082421_, _082422_, _082423_, _082424_, _082425_, _082426_, _082427_, _082428_, _082429_, _082430_, _082431_, _082432_, _082433_, _082434_, _082435_, _082436_, _082437_, _082438_, _082439_, _082440_, _082441_, _082442_, _082443_, _082444_, _082445_, _082446_, _082447_, _082448_, _082449_, _082450_, _082451_, _082452_, _082453_, _082454_, _082455_, _082456_, _082457_, _082458_, _082459_, _082460_, _082461_, _082462_, _082463_, _082464_, _082465_, _082466_, _082467_, _082468_, _082469_, _082470_, _082471_, _082472_, _082473_, _082474_, _082475_, _082476_, _082477_, _082478_, _082479_, _082480_, _082481_, _082482_, _082483_, _082484_, _082485_, _082486_, _082487_, _082488_, _082489_, _082490_, _082491_, _082492_, _082493_, _082494_, _082495_, _082496_, _082497_, _082498_, _082499_, _082500_, _082501_, _082502_, _082503_, _082504_, _082505_, _082506_, _082507_, _082508_, _082509_, _082510_, _082511_, _082512_, _082513_, _082514_, _082515_, _082516_, _082517_, _082518_, _082519_, _082520_, _082521_, _082522_, _082523_, _082524_, _082525_, _082526_, _082527_, _082528_, _082529_, _082530_, _082531_, _082532_, _082533_, _082534_, _082535_, _082536_, _082537_, _082538_, _082539_, _082540_, _082541_, _082542_, _082543_, _082544_, _082545_, _082546_, _082547_, _082548_, _082549_, _082550_, _082551_, _082552_, _082553_, _082554_, _082555_, _082556_, _082557_, _082558_, _082559_, _082560_, _082561_, _082562_, _082563_, _082564_, _082565_, _082566_, _082567_, _082568_, _082569_, _082570_, _082571_, _082572_, _082573_, _082574_, _082575_, _082576_, _082577_, _082578_, _082579_, _082580_, _082581_, _082582_, _082583_, _082584_, _082585_, _082586_, _082587_, _082588_, _082589_, _082590_, _082591_, _082592_, _082593_, _082594_, _082595_, _082596_, _082597_, _082598_, _082599_, _082600_, _082601_, _082602_, _082603_, _082604_, _082605_, _082606_, _082607_, _082608_, _082609_, _082610_, _082611_, _082612_, _082613_, _082614_, _082615_, _082616_, _082617_, _082618_, _082619_, _082620_, _082621_, _082622_, _082623_, _082624_, _082625_, _082626_, _082627_, _082628_, _082629_, _082630_, _082631_, _082632_, _082633_, _082634_, _082635_, _082636_, _082637_, _082638_, _082639_, _082640_, _082641_, _082642_, _082643_, _082644_, _082645_, _082646_, _082647_, _082648_, _082649_, _082650_, _082651_, _082652_, _082653_, _082654_, _082655_, _082656_, _082657_, _082658_, _082659_, _082660_, _082661_, _082662_, _082663_, _082664_, _082665_, _082666_, _082667_, _082668_, _082669_, _082670_, _082671_, _082672_, _082673_, _082674_, _082675_, _082676_, _082677_, _082678_, _082679_, _082680_, _082681_, _082682_, _082683_, _082684_, _082685_, _082686_, _082687_, _082688_, _082689_, _082690_, _082691_, _082692_, _082693_, _082694_, _082695_, _082696_, _082697_, _082698_, _082699_, _082700_, _082701_, _082702_, _082703_, _082704_, _082705_, _082706_, _082707_, _082708_, _082709_, _082710_, _082711_, _082712_, _082713_, _082714_, _082715_, _082716_, _082717_, _082718_, _082719_, _082720_, _082721_, _082722_, _082723_, _082724_, _082725_, _082726_, _082727_, _082728_, _082729_, _082730_, _082731_, _082732_, _082733_, _082734_, _082735_, _082736_, _082737_, _082738_, _082739_, _082740_, _082741_, _082742_, _082743_, _082744_, _082745_, _082746_, _082747_, _082748_, _082749_, _082750_, _082751_, _082752_, _082753_, _082754_, _082755_, _082756_, _082757_, _082758_, _082759_, _082760_, _082761_, _082762_, _082763_, _082764_, _082765_, _082766_, _082767_, _082768_, _082769_, _082770_, _082771_, _082772_, _082773_, _082774_, _082775_, _082776_, _082777_, _082778_, _082779_, _082780_, _082781_, _082782_, _082783_, _082784_, _082785_, _082786_, _082787_, _082788_, _082789_, _082790_, _082791_, _082792_, _082793_, _082794_, _082795_, _082796_, _082797_, _082798_, _082799_, _082800_, _082801_, _082802_, _082803_, _082804_, _082805_, _082806_, _082807_, _082808_, _082809_, _082810_, _082811_, _082812_, _082813_, _082814_, _082815_, _082816_, _082817_, _082818_, _082819_, _082820_, _082821_, _082822_, _082823_, _082824_, _082825_, _082826_, _082827_, _082828_, _082829_, _082830_, _082831_, _082832_, _082833_, _082834_, _082835_, _082836_, _082837_, _082838_, _082839_, _082840_, _082841_, _082842_, _082843_, _082844_, _082845_, _082846_, _082847_, _082848_, _082849_, _082850_, _082851_, _082852_, _082853_, _082854_, _082855_, _082856_, _082857_, _082858_, _082859_, _082860_, _082861_, _082862_, _082863_, _082864_, _082865_, _082866_, _082867_, _082868_, _082869_, _082870_, _082871_, _082872_, _082873_, _082874_, _082875_, _082876_, _082877_, _082878_, _082879_, _082880_, _082881_, _082882_, _082883_, _082884_, _082885_, _082886_, _082887_, _082888_, _082889_, _082890_, _082891_, _082892_, _082893_, _082894_, _082895_, _082896_, _082897_, _082898_, _082899_, _082900_, _082901_, _082902_, _082903_, _082904_, _082905_, _082906_, _082907_, _082908_, _082909_, _082910_, _082911_, _082912_, _082913_, _082914_, _082915_, _082916_, _082917_, _082918_, _082919_, _082920_, _082921_, _082922_, _082923_, _082924_, _082925_, _082926_, _082927_, _082928_, _082929_, _082930_, _082931_, _082932_, _082933_, _082934_, _082935_, _082936_, _082937_, _082938_, _082939_, _082940_, _082941_, _082942_, _082943_, _082944_, _082945_, _082946_, _082947_, _082948_, _082949_, _082950_, _082951_, _082952_, _082953_, _082954_, _082955_, _082956_, _082957_, _082958_, _082959_, _082960_, _082961_, _082962_, _082963_, _082964_, _082965_, _082966_, _082967_, _082968_, _082969_, _082970_, _082971_, _082972_, _082973_, _082974_, _082975_, _082976_, _082977_, _082978_, _082979_, _082980_, _082981_, _082982_, _082983_, _082984_, _082985_, _082986_, _082987_, _082988_, _082989_, _082990_, _082991_, _082992_, _082993_, _082994_, _082995_, _082996_, _082997_, _082998_, _082999_, _083000_, _083001_, _083002_, _083003_, _083004_, _083005_, _083006_, _083007_, _083008_, _083009_, _083010_, _083011_, _083012_, _083013_, _083014_, _083015_, _083016_, _083017_, _083018_, _083019_, _083020_, _083021_, _083022_, _083023_, _083024_, _083025_, _083026_, _083027_, _083028_, _083029_, _083030_, _083031_, _083032_, _083033_, _083034_, _083035_, _083036_, _083037_, _083038_, _083039_, _083040_, _083041_, _083042_, _083043_, _083044_, _083045_, _083046_, _083047_, _083048_, _083049_, _083050_, _083051_, _083052_, _083053_, _083054_, _083055_, _083056_, _083057_, _083058_, _083059_, _083060_, _083061_, _083062_, _083063_, _083064_, _083065_, _083066_, _083067_, _083068_, _083069_, _083070_, _083071_, _083072_, _083073_, _083074_, _083075_, _083076_, _083077_, _083078_, _083079_, _083080_, _083081_, _083082_, _083083_, _083084_, _083085_, _083086_, _083087_, _083088_, _083089_, _083090_, _083091_, _083092_, _083093_, _083094_, _083095_, _083096_, _083097_, _083098_, _083099_, _083100_, _083101_, _083102_, _083103_, _083104_, _083105_, _083106_, _083107_, _083108_, _083109_, _083110_, _083111_, _083112_, _083113_, _083114_, _083115_, _083116_, _083117_, _083118_, _083119_, _083120_, _083121_, _083122_, _083123_, _083124_, _083125_, _083126_, _083127_, _083128_, _083129_, _083130_, _083131_, _083132_, _083133_, _083134_, _083135_, _083136_, _083137_, _083138_, _083139_, _083140_, _083141_, _083142_, _083143_, _083144_, _083145_, _083146_, _083147_, _083148_, _083149_, _083150_, _083151_, _083152_, _083153_, _083154_, _083155_, _083156_, _083157_, _083158_, _083159_, _083160_, _083161_, _083162_, _083163_, _083164_, _083165_, _083166_, _083167_, _083168_, _083169_, _083170_, _083171_, _083172_, _083173_, _083174_, _083175_, _083176_, _083177_, _083178_, _083179_, _083180_, _083181_, _083182_, _083183_, _083184_, _083185_, _083186_, _083187_, _083188_, _083189_, _083190_, _083191_, _083192_, _083193_, _083194_, _083195_, _083196_, _083197_, _083198_, _083199_, _083200_, _083201_, _083202_, _083203_, _083204_, _083205_, _083206_, _083207_, _083208_, _083209_, _083210_, _083211_, _083212_, _083213_, _083214_, _083215_, _083216_, _083217_, _083218_, _083219_, _083220_, _083221_, _083222_, _083223_, _083224_, _083225_, _083226_, _083227_, _083228_, _083229_, _083230_, _083231_, _083232_, _083233_, _083234_, _083235_, _083236_, _083237_, _083238_, _083239_, _083240_, _083241_, _083242_, _083243_, _083244_, _083245_, _083246_, _083247_, _083248_, _083249_, _083250_, _083251_, _083252_, _083253_, _083254_, _083255_, _083256_, _083257_, _083258_, _083259_, _083260_, _083261_, _083262_, _083263_, _083264_, _083265_, _083266_, _083267_, _083268_, _083269_, _083270_, _083271_, _083272_, _083273_, _083274_, _083275_, _083276_, _083277_, _083278_, _083279_, _083280_, _083281_, _083282_, _083283_, _083284_, _083285_, _083286_, _083287_, _083288_, _083289_, _083290_, _083291_, _083292_, _083293_, _083294_, _083295_, _083296_, _083297_, _083298_, _083299_, _083300_, _083301_, _083302_, _083303_, _083304_, _083305_, _083306_, _083307_, _083308_, _083309_, _083310_, _083311_, _083312_, _083313_, _083314_, _083315_, _083316_, _083317_, _083318_, _083319_, _083320_, _083321_, _083322_, _083323_, _083324_, _083325_, _083326_, _083327_, _083328_, _083329_, _083330_, _083331_, _083332_, _083333_, _083334_, _083335_, _083336_, _083337_, _083338_, _083339_, _083340_, _083341_, _083342_, _083343_, _083344_, _083345_, _083346_, _083347_, _083348_, _083349_, _083350_, _083351_, _083352_, _083353_, _083354_, _083355_, _083356_, _083357_, _083358_, _083359_, _083360_, _083361_, _083362_, _083363_, _083364_, _083365_, _083366_, _083367_, _083368_, _083369_, _083370_, _083371_, _083372_, _083373_, _083374_, _083375_, _083376_, _083377_, _083378_, _083379_, _083380_, _083381_, _083382_, _083383_, _083384_, _083385_, _083386_, _083387_, _083388_, _083389_, _083390_, _083391_, _083392_, _083393_, _083394_, _083395_, _083396_, _083397_, _083398_, _083399_, _083400_, _083401_, _083402_, _083403_, _083404_, _083405_, _083406_, _083407_, _083408_, _083409_, _083410_, _083411_, _083412_, _083413_, _083414_, _083415_, _083416_, _083417_, _083418_, _083419_, _083420_, _083421_, _083422_, _083423_, _083424_, _083425_, _083426_, _083427_, _083428_, _083429_, _083430_, _083431_, _083432_, _083433_, _083434_, _083435_, _083436_, _083437_, _083438_, _083439_, _083440_, _083441_, _083442_, _083443_, _083444_, _083445_, _083446_, _083447_, _083448_, _083449_, _083450_, _083451_, _083452_, _083453_, _083454_, _083455_, _083456_, _083457_, _083458_, _083459_, _083460_, _083461_, _083462_, _083463_, _083464_, _083465_, _083466_, _083467_, _083468_, _083469_, _083470_, _083471_, _083472_, _083473_, _083474_, _083475_, _083476_, _083477_, _083478_, _083479_, _083480_, _083481_, _083482_, _083483_, _083484_, _083485_, _083486_, _083487_, _083488_, _083489_, _083490_, _083491_, _083492_, _083493_, _083494_, _083495_, _083496_, _083497_, _083498_, _083499_, _083500_, _083501_, _083502_, _083503_, _083504_, _083505_, _083506_, _083507_, _083508_, _083509_, _083510_, _083511_, _083512_, _083513_, _083514_, _083515_, _083516_, _083517_, _083518_, _083519_, _083520_, _083521_, _083522_, _083523_, _083524_, _083525_, _083526_, _083527_, _083528_, _083529_, _083530_, _083531_, _083532_, _083533_, _083534_, _083535_, _083536_, _083537_, _083538_, _083539_, _083540_, _083541_, _083542_, _083543_, _083544_, _083545_, _083546_, _083547_, _083548_, _083549_, _083550_, _083551_, _083552_, _083553_, _083554_, _083555_, _083556_, _083557_, _083558_, _083559_, _083560_, _083561_, _083562_, _083563_, _083564_, _083565_, _083566_, _083567_, _083568_, _083569_, _083570_, _083571_, _083572_, _083573_, _083574_, _083575_, _083576_, _083577_, _083578_, _083579_, _083580_, _083581_, _083582_, _083583_, _083584_, _083585_, _083586_, _083587_, _083588_, _083589_, _083590_, _083591_, _083592_, _083593_, _083594_, _083595_, _083596_, _083597_, _083598_, _083599_, _083600_, _083601_, _083602_, _083603_, _083604_, _083605_, _083606_, _083607_, _083608_, _083609_, _083610_, _083611_, _083612_, _083613_, _083614_, _083615_, _083616_, _083617_, _083618_, _083619_, _083620_, _083621_, _083622_, _083623_, _083624_, _083625_, _083626_, _083627_, _083628_, _083629_, _083630_, _083631_, _083632_, _083633_, _083634_, _083635_, _083636_, _083637_, _083638_, _083639_, _083640_, _083641_, _083642_, _083643_, _083644_, _083645_, _083646_, _083647_, _083648_, _083649_, _083650_, _083651_, _083652_, _083653_, _083654_, _083655_, _083656_, _083657_, _083658_, _083659_, _083660_, _083661_, _083662_, _083663_, _083664_, _083665_, _083666_, _083667_, _083668_, _083669_, _083670_, _083671_, _083672_, _083673_, _083674_, _083675_, _083676_, _083677_, _083678_, _083679_, _083680_, _083681_, _083682_, _083683_, _083684_, _083685_, _083686_, _083687_, _083688_, _083689_, _083690_, _083691_, _083692_, _083693_, _083694_, _083695_, _083696_, _083697_, _083698_, _083699_, _083700_, _083701_, _083702_, _083703_, _083704_, _083705_, _083706_, _083707_, _083708_, _083709_, _083710_, _083711_, _083712_, _083713_, _083714_, _083715_, _083716_, _083717_, _083718_, _083719_, _083720_, _083721_, _083722_, _083723_, _083724_, _083725_, _083726_, _083727_, _083728_, _083729_, _083730_, _083731_, _083732_, _083733_, _083734_, _083735_, _083736_, _083737_, _083738_, _083739_, _083740_, _083741_, _083742_, _083743_, _083744_, _083745_, _083746_, _083747_, _083748_, _083749_, _083750_, _083751_, _083752_, _083753_, _083754_, _083755_, _083756_, _083757_, _083758_, _083759_, _083760_, _083761_, _083762_, _083763_, _083764_, _083765_, _083766_, _083767_, _083768_, _083769_, _083770_, _083771_, _083772_, _083773_, _083774_, _083775_, _083776_, _083777_, _083778_, _083779_, _083780_, _083781_, _083782_, _083783_, _083784_, _083785_, _083786_, _083787_, _083788_, _083789_, _083790_, _083791_, _083792_, _083793_, _083794_, _083795_, _083796_, _083797_, _083798_, _083799_, _083800_, _083801_, _083802_, _083803_, _083804_, _083805_, _083806_, _083807_, _083808_, _083809_, _083810_, _083811_, _083812_, _083813_, _083814_, _083815_, _083816_, _083817_, _083818_, _083819_, _083820_, _083821_, _083822_, _083823_, _083824_, _083825_, _083826_, _083827_, _083828_, _083829_, _083830_, _083831_, _083832_, _083833_, _083834_, _083835_, _083836_, _083837_, _083838_, _083839_, _083840_, _083841_, _083842_, _083843_, _083844_, _083845_, _083846_, _083847_, _083848_, _083849_, _083850_, _083851_, _083852_, _083853_, _083854_, _083855_, _083856_, _083857_, _083858_, _083859_, _083860_, _083861_, _083862_, _083863_, _083864_, _083865_, _083866_, _083867_, _083868_, _083869_, _083870_, _083871_, _083872_, _083873_, _083874_, _083875_, _083876_, _083877_, _083878_, _083879_, _083880_, _083881_, _083882_, _083883_, _083884_, _083885_, _083886_, _083887_, _083888_, _083889_, _083890_, _083891_, _083892_, _083893_, _083894_, _083895_, _083896_, _083897_, _083898_, _083899_, _083900_, _083901_, _083902_, _083903_, _083904_, _083905_, _083906_, _083907_, _083908_, _083909_, _083910_, _083911_, _083912_, _083913_, _083914_, _083915_, _083916_, _083917_, _083918_, _083919_, _083920_, _083921_, _083922_, _083923_, _083924_, _083925_, _083926_, _083927_, _083928_, _083929_, _083930_, _083931_, _083932_, _083933_, _083934_, _083935_, _083936_, _083937_, _083938_, _083939_, _083940_, _083941_, _083942_, _083943_, _083944_, _083945_, _083946_, _083947_, _083948_, _083949_, _083950_, _083951_, _083952_, _083953_, _083954_, _083955_, _083956_, _083957_, _083958_, _083959_, _083960_, _083961_, _083962_, _083963_, _083964_, _083965_, _083966_, _083967_, _083968_, _083969_, _083970_, _083971_, _083972_, _083973_, _083974_, _083975_, _083976_, _083977_, _083978_, _083979_, _083980_, _083981_, _083982_, _083983_, _083984_, _083985_, _083986_, _083987_, _083988_, _083989_, _083990_, _083991_, _083992_, _083993_, _083994_, _083995_, _083996_, _083997_, _083998_, _083999_, _084000_, _084001_, _084002_, _084003_, _084004_, _084005_, _084006_, _084007_, _084008_, _084009_, _084010_, _084011_, _084012_, _084013_, _084014_, _084015_, _084016_, _084017_, _084018_, _084019_, _084020_, _084021_, _084022_, _084023_, _084024_, _084025_, _084026_, _084027_, _084028_, _084029_, _084030_, _084031_, _084032_, _084033_, _084034_, _084035_, _084036_, _084037_, _084038_, _084039_, _084040_, _084041_, _084042_, _084043_, _084044_, _084045_, _084046_, _084047_, _084048_, _084049_, _084050_, _084051_, _084052_, _084053_, _084054_, _084055_, _084056_, _084057_, _084058_, _084059_, _084060_, _084061_, _084062_, _084063_, _084064_, _084065_, _084066_, _084067_, _084068_, _084069_, _084070_, _084071_, _084072_, _084073_, _084074_, _084075_, _084076_, _084077_, _084078_, _084079_, _084080_, _084081_, _084082_, _084083_, _084084_, _084085_, _084086_, _084087_, _084088_, _084089_, _084090_, _084091_, _084092_, _084093_, _084094_, _084095_, _084096_, _084097_, _084098_, _084099_, _084100_, _084101_, _084102_, _084103_, _084104_, _084105_, _084106_, _084107_, _084108_, _084109_, _084110_, _084111_, _084112_, _084113_, _084114_, _084115_, _084116_, _084117_, _084118_, _084119_, _084120_, _084121_, _084122_, _084123_, _084124_, _084125_, _084126_, _084127_, _084128_, _084129_, _084130_, _084131_, _084132_, _084133_, _084134_, _084135_, _084136_, _084137_, _084138_, _084139_, _084140_, _084141_, _084142_, _084143_, _084144_, _084145_, _084146_, _084147_, _084148_, _084149_, _084150_, _084151_, _084152_, _084153_, _084154_, _084155_, _084156_, _084157_, _084158_, _084159_, _084160_, _084161_, _084162_, _084163_, _084164_, _084165_, _084166_, _084167_, _084168_, _084169_, _084170_, _084171_, _084172_, _084173_, _084174_, _084175_, _084176_, _084177_, _084178_, _084179_, _084180_, _084181_, _084182_, _084183_, _084184_, _084185_, _084186_, _084187_, _084188_, _084189_, _084190_, _084191_, _084192_, _084193_, _084194_, _084195_, _084196_, _084197_, _084198_, _084199_, _084200_, _084201_, _084202_, _084203_, _084204_, _084205_, _084206_, _084207_, _084208_, _084209_, _084210_, _084211_, _084212_, _084213_, _084214_, _084215_, _084216_, _084217_, _084218_, _084219_, _084220_, _084221_, _084222_, _084223_, _084224_, _084225_, _084226_, _084227_, _084228_, _084229_, _084230_, _084231_, _084232_, _084233_, _084234_, _084235_, _084236_, _084237_, _084238_, _084239_, _084240_, _084241_, _084242_, _084243_, _084244_, _084245_, _084246_, _084247_, _084248_, _084249_, _084250_, _084251_, _084252_, _084253_, _084254_, _084255_, _084256_, _084257_, _084258_, _084259_, _084260_, _084261_, _084262_, _084263_, _084264_, _084265_, _084266_, _084267_, _084268_, _084269_, _084270_, _084271_, _084272_, _084273_, _084274_, _084275_, _084276_, _084277_, _084278_, _084279_, _084280_, _084281_, _084282_, _084283_, _084284_, _084285_, _084286_, _084287_, _084288_, _084289_, _084290_, _084291_, _084292_, _084293_, _084294_, _084295_, _084296_, _084297_, _084298_, _084299_, _084300_, _084301_, _084302_, _084303_, _084304_, _084305_, _084306_, _084307_, _084308_, _084309_, _084310_, _084311_, _084312_, _084313_, _084314_, _084315_, _084316_, _084317_, _084318_, _084319_, _084320_, _084321_, _084322_, _084323_, _084324_, _084325_, _084326_, _084327_, _084328_, _084329_, _084330_, _084331_, _084332_, _084333_, _084334_, _084335_, _084336_, _084337_, _084338_, _084339_, _084340_, _084341_, _084342_, _084343_, _084344_, _084345_, _084346_, _084347_, _084348_, _084349_, _084350_, _084351_, _084352_, _084353_, _084354_, _084355_, _084356_, _084357_, _084358_, _084359_, _084360_, _084361_, _084362_, _084363_, _084364_, _084365_, _084366_, _084367_, _084368_, _084369_, _084370_, _084371_, _084372_, _084373_, _084374_, _084375_, _084376_, _084377_, _084378_, _084379_, _084380_, _084381_, _084382_, _084383_, _084384_, _084385_, _084386_, _084387_, _084388_, _084389_, _084390_, _084391_, _084392_, _084393_, _084394_, _084395_, _084396_, _084397_, _084398_, _084399_, _084400_, _084401_, _084402_, _084403_, _084404_, _084405_, _084406_, _084407_, _084408_, _084409_, _084410_, _084411_, _084412_, _084413_, _084414_, _084415_, _084416_, _084417_, _084418_, _084419_, _084420_, _084421_, _084422_, _084423_, _084424_, _084425_, _084426_, _084427_, _084428_, _084429_, _084430_, _084431_, _084432_, _084433_, _084434_, _084435_, _084436_, _084437_, _084438_, _084439_, _084440_, _084441_, _084442_, _084443_, _084444_, _084445_, _084446_, _084447_, _084448_, _084449_, _084450_, _084451_, _084452_, _084453_, _084454_, _084455_, _084456_, _084457_, _084458_, _084459_, _084460_, _084461_, _084462_, _084463_, _084464_, _084465_, _084466_, _084467_, _084468_, _084469_, _084470_, _084471_, _084472_, _084473_, _084474_, _084475_, _084476_, _084477_, _084478_, _084479_, _084480_, _084481_, _084482_, _084483_, _084484_, _084485_, _084486_, _084487_, _084488_, _084489_, _084490_, _084491_, _084492_, _084493_, _084494_, _084495_, _084496_, _084497_, _084498_, _084499_, _084500_, _084501_, _084502_, _084503_, _084504_, _084505_, _084506_, _084507_, _084508_, _084509_, _084510_, _084511_, _084512_, _084513_, _084514_, _084515_, _084516_, _084517_, _084518_, _084519_, _084520_, _084521_, _084522_, _084523_, _084524_, _084525_, _084526_, _084527_, _084528_, _084529_, _084530_, _084531_, _084532_, _084533_, _084534_, _084535_, _084536_, _084537_, _084538_, _084539_, _084540_, _084541_, _084542_, _084543_, _084544_, _084545_, _084546_, _084547_, _084548_, _084549_, _084550_, _084551_, _084552_, _084553_, _084554_, _084555_, _084556_, _084557_, _084558_, _084559_, _084560_, _084561_, _084562_, _084563_, _084564_, _084565_, _084566_, _084567_, _084568_, _084569_, _084570_, _084571_, _084572_, _084573_, _084574_, _084575_, _084576_, _084577_, _084578_, _084579_, _084580_, _084581_, _084582_, _084583_, _084584_, _084585_, _084586_, _084587_, _084588_, _084589_, _084590_, _084591_, _084592_, _084593_, _084594_, _084595_, _084596_, _084597_, _084598_, _084599_, _084600_, _084601_, _084602_, _084603_, _084604_, _084605_, _084606_, _084607_, _084608_, _084609_, _084610_, _084611_, _084612_, _084613_, _084614_, _084615_, _084616_, _084617_, _084618_, _084619_, _084620_, _084621_, _084622_, _084623_, _084624_, _084625_, _084626_, _084627_, _084628_, _084629_, _084630_, _084631_, _084632_, _084633_, _084634_, _084635_, _084636_, _084637_, _084638_, _084639_, _084640_, _084641_, _084642_, _084643_, _084644_, _084645_, _084646_, _084647_, _084648_, _084649_, _084650_, _084651_, _084652_, _084653_, _084654_, _084655_, _084656_, _084657_, _084658_, _084659_, _084660_, _084661_, _084662_, _084663_, _084664_, _084665_, _084666_, _084667_, _084668_, _084669_, _084670_, _084671_, _084672_, _084673_, _084674_, _084675_, _084676_, _084677_, _084678_, _084679_, _084680_, _084681_, _084682_, _084683_, _084684_, _084685_, _084686_, _084687_, _084688_, _084689_, _084690_, _084691_, _084692_, _084693_, _084694_, _084695_, _084696_, _084697_, _084698_, _084699_, _084700_, _084701_, _084702_, _084703_, _084704_, _084705_, _084706_, _084707_, _084708_, _084709_, _084710_, _084711_, _084712_, _084713_, _084714_, _084715_, _084716_, _084717_, _084718_, _084719_, _084720_, _084721_, _084722_, _084723_, _084724_, _084725_, _084726_, _084727_, _084728_, _084729_, _084730_, _084731_, _084732_, _084733_, _084734_, _084735_, _084736_, _084737_, _084738_, _084739_, _084740_, _084741_, _084742_, _084743_, _084744_, _084745_, _084746_, _084747_, _084748_, _084749_, _084750_, _084751_, _084752_, _084753_, _084754_, _084755_, _084756_, _084757_, _084758_, _084759_, _084760_, _084761_, _084762_, _084763_, _084764_, _084765_, _084766_, _084767_, _084768_, _084769_, _084770_, _084771_, _084772_, _084773_, _084774_, _084775_, _084776_, _084777_, _084778_, _084779_, _084780_, _084781_, _084782_, _084783_, _084784_, _084785_, _084786_, _084787_, _084788_, _084789_, _084790_, _084791_, _084792_, _084793_, _084794_, _084795_, _084796_, _084797_, _084798_, _084799_, _084800_, _084801_, _084802_, _084803_, _084804_, _084805_, _084806_, _084807_, _084808_, _084809_, _084810_, _084811_, _084812_, _084813_, _084814_, _084815_, _084816_, _084817_, _084818_, _084819_, _084820_, _084821_, _084822_, _084823_, _084824_, _084825_, _084826_, _084827_, _084828_, _084829_, _084830_, _084831_, _084832_, _084833_, _084834_, _084835_, _084836_, _084837_, _084838_, _084839_, _084840_, _084841_, _084842_, _084843_, _084844_, _084845_, _084846_, _084847_, _084848_, _084849_, _084850_, _084851_, _084852_, _084853_, _084854_, _084855_, _084856_, _084857_, _084858_, _084859_, _084860_, _084861_, _084862_, _084863_, _084864_, _084865_, _084866_, _084867_, _084868_, _084869_, _084870_, _084871_, _084872_, _084873_, _084874_, _084875_, _084876_, _084877_, _084878_, _084879_, _084880_, _084881_, _084882_, _084883_, _084884_, _084885_, _084886_, _084887_, _084888_, _084889_, _084890_, _084891_, _084892_, _084893_, _084894_, _084895_, _084896_, _084897_, _084898_, _084899_, _084900_, _084901_, _084902_, _084903_, _084904_, _084905_, _084906_, _084907_, _084908_, _084909_, _084910_, _084911_, _084912_, _084913_, _084914_, _084915_, _084916_, _084917_, _084918_, _084919_, _084920_, _084921_, _084922_, _084923_, _084924_, _084925_, _084926_, _084927_, _084928_, _084929_, _084930_, _084931_, _084932_, _084933_, _084934_, _084935_, _084936_, _084937_, _084938_, _084939_, _084940_, _084941_, _084942_, _084943_, _084944_, _084945_, _084946_, _084947_, _084948_, _084949_, _084950_, _084951_, _084952_, _084953_, _084954_, _084955_, _084956_, _084957_, _084958_, _084959_, _084960_, _084961_, _084962_, _084963_, _084964_, _084965_, _084966_, _084967_, _084968_, _084969_, _084970_, _084971_, _084972_, _084973_, _084974_, _084975_, _084976_, _084977_, _084978_, _084979_, _084980_, _084981_, _084982_, _084983_, _084984_, _084985_, _084986_, _084987_, _084988_, _084989_, _084990_, _084991_, _084992_, _084993_, _084994_, _084995_, _084996_, _084997_, _084998_, _084999_, _085000_, _085001_, _085002_, _085003_, _085004_, _085005_, _085006_, _085007_, _085008_, _085009_, _085010_, _085011_, _085012_, _085013_, _085014_, _085015_, _085016_, _085017_, _085018_, _085019_, _085020_, _085021_, _085022_, _085023_, _085024_, _085025_, _085026_, _085027_, _085028_, _085029_, _085030_, _085031_, _085032_, _085033_, _085034_, _085035_, _085036_, _085037_, _085038_, _085039_, _085040_, _085041_, _085042_, _085043_, _085044_, _085045_, _085046_, _085047_, _085048_, _085049_, _085050_, _085051_, _085052_, _085053_, _085054_, _085055_, _085056_, _085057_, _085058_, _085059_, _085060_, _085061_, _085062_, _085063_, _085064_, _085065_, _085066_, _085067_, _085068_, _085069_, _085070_, _085071_, _085072_, _085073_, _085074_, _085075_, _085076_, _085077_, _085078_, _085079_, _085080_, _085081_, _085082_, _085083_, _085084_, _085085_, _085086_, _085087_, _085088_, _085089_, _085090_, _085091_, _085092_, _085093_, _085094_, _085095_, _085096_, _085097_, _085098_, _085099_, _085100_, _085101_, _085102_, _085103_, _085104_, _085105_, _085106_, _085107_, _085108_, _085109_, _085110_, _085111_, _085112_, _085113_, _085114_, _085115_, _085116_, _085117_, _085118_, _085119_, _085120_, _085121_, _085122_, _085123_, _085124_, _085125_, _085126_, _085127_, _085128_, _085129_, _085130_, _085131_, _085132_, _085133_, _085134_, _085135_, _085136_, _085137_, _085138_, _085139_, _085140_, _085141_, _085142_, _085143_, _085144_, _085145_, _085146_, _085147_, _085148_, _085149_, _085150_, _085151_, _085152_, _085153_, _085154_, _085155_, _085156_, _085157_, _085158_, _085159_, _085160_, _085161_, _085162_, _085163_, _085164_, _085165_, _085166_, _085167_, _085168_, _085169_, _085170_, _085171_, _085172_, _085173_, _085174_, _085175_, _085176_, _085177_, _085178_, _085179_, _085180_, _085181_, _085182_, _085183_, _085184_, _085185_, _085186_, _085187_, _085188_, _085189_, _085190_, _085191_, _085192_, _085193_, _085194_, _085195_, _085196_, _085197_, _085198_, _085199_, _085200_, _085201_, _085202_, _085203_, _085204_, _085205_, _085206_, _085207_, _085208_, _085209_, _085210_, _085211_, _085212_, _085213_, _085214_, _085215_, _085216_, _085217_, _085218_, _085219_, _085220_, _085221_, _085222_, _085223_, _085224_, _085225_, _085226_, _085227_, _085228_, _085229_, _085230_, _085231_, _085232_, _085233_, _085234_, _085235_, _085236_, _085237_, _085238_, _085239_, _085240_, _085241_, _085242_, _085243_, _085244_, _085245_, _085246_, _085247_, _085248_, _085249_, _085250_, _085251_, _085252_, _085253_, _085254_, _085255_, _085256_, _085257_, _085258_, _085259_, _085260_, _085261_, _085262_, _085263_, _085264_, _085265_, _085266_, _085267_, _085268_, _085269_, _085270_, _085271_, _085272_, _085273_, _085274_, _085275_, _085276_, _085277_, _085278_, _085279_, _085280_, _085281_, _085282_, _085283_, _085284_, _085285_, _085286_, _085287_, _085288_, _085289_, _085290_, _085291_, _085292_, _085293_, _085294_, _085295_, _085296_, _085297_, _085298_, _085299_, _085300_, _085301_, _085302_, _085303_, _085304_, _085305_, _085306_, _085307_, _085308_, _085309_, _085310_, _085311_, _085312_, _085313_, _085314_, _085315_, _085316_, _085317_, _085318_, _085319_, _085320_, _085321_, _085322_, _085323_, _085324_, _085325_, _085326_, _085327_, _085328_, _085329_, _085330_, _085331_, _085332_, _085333_, _085334_, _085335_, _085336_, _085337_, _085338_, _085339_, _085340_, _085341_, _085342_, _085343_, _085344_, _085345_, _085346_, _085347_, _085348_, _085349_, _085350_, _085351_, _085352_, _085353_, _085354_, _085355_, _085356_, _085357_, _085358_, _085359_, _085360_, _085361_, _085362_, _085363_, _085364_, _085365_, _085366_, _085367_, _085368_, _085369_, _085370_, _085371_, _085372_, _085373_, _085374_, _085375_, _085376_, _085377_, _085378_, _085379_, _085380_, _085381_, _085382_, _085383_, _085384_, _085385_, _085386_, _085387_, _085388_, _085389_, _085390_, _085391_, _085392_, _085393_, _085394_, _085395_, _085396_, _085397_, _085398_, _085399_, _085400_, _085401_, _085402_, _085403_, _085404_, _085405_, _085406_, _085407_, _085408_, _085409_, _085410_, _085411_, _085412_, _085413_, _085414_, _085415_, _085416_, _085417_, _085418_, _085419_, _085420_, _085421_, _085422_, _085423_, _085424_, _085425_, _085426_, _085427_, _085428_, _085429_, _085430_, _085431_, _085432_, _085433_, _085434_, _085435_, _085436_, _085437_, _085438_, _085439_, _085440_, _085441_, _085442_, _085443_, _085444_, _085445_, _085446_, _085447_, _085448_, _085449_, _085450_, _085451_, _085452_, _085453_, _085454_, _085455_, _085456_, _085457_, _085458_, _085459_, _085460_, _085461_, _085462_, _085463_, _085464_, _085465_, _085466_, _085467_, _085468_, _085469_, _085470_, _085471_, _085472_, _085473_, _085474_, _085475_, _085476_, _085477_, _085478_, _085479_, _085480_, _085481_, _085482_, _085483_, _085484_, _085485_, _085486_, _085487_, _085488_, _085489_, _085490_, _085491_, _085492_, _085493_, _085494_, _085495_, _085496_, _085497_, _085498_, _085499_, _085500_, _085501_, _085502_, _085503_, _085504_, _085505_, _085506_, _085507_, _085508_, _085509_, _085510_, _085511_, _085512_, _085513_, _085514_, _085515_, _085516_, _085517_, _085518_, _085519_, _085520_, _085521_, _085522_, _085523_, _085524_, _085525_, _085526_, _085527_, _085528_, _085529_, _085530_, _085531_, _085532_, _085533_, _085534_, _085535_, _085536_, _085537_, _085538_, _085539_, _085540_, _085541_, _085542_, _085543_, _085544_, _085545_, _085546_, _085547_, _085548_, _085549_, _085550_, _085551_, _085552_, _085553_, _085554_, _085555_, _085556_, _085557_, _085558_, _085559_, _085560_, _085561_, _085562_, _085563_, _085564_, _085565_, _085566_, _085567_, _085568_, _085569_, _085570_, _085571_, _085572_, _085573_, _085574_, _085575_, _085576_, _085577_, _085578_, _085579_, _085580_, _085581_, _085582_, _085583_, _085584_, _085585_, _085586_, _085587_, _085588_, _085589_, _085590_, _085591_, _085592_, _085593_, _085594_, _085595_, _085596_, _085597_, _085598_, _085599_, _085600_, _085601_, _085602_, _085603_, _085604_, _085605_, _085606_, _085607_, _085608_, _085609_, _085610_, _085611_, _085612_, _085613_, _085614_, _085615_, _085616_, _085617_, _085618_, _085619_, _085620_, _085621_, _085622_, _085623_, _085624_, _085625_, _085626_, _085627_, _085628_, _085629_, _085630_, _085631_, _085632_, _085633_, _085634_, _085635_, _085636_, _085637_, _085638_, _085639_, _085640_, _085641_, _085642_, _085643_, _085644_, _085645_, _085646_, _085647_, _085648_, _085649_, _085650_, _085651_, _085652_, _085653_, _085654_, _085655_, _085656_, _085657_, _085658_, _085659_, _085660_, _085661_, _085662_, _085663_, _085664_, _085665_, _085666_, _085667_, _085668_, _085669_, _085670_, _085671_, _085672_, _085673_, _085674_, _085675_, _085676_, _085677_, _085678_, _085679_, _085680_, _085681_, _085682_, _085683_, _085684_, _085685_, _085686_, _085687_, _085688_, _085689_, _085690_, _085691_, _085692_, _085693_, _085694_, _085695_, _085696_, _085697_, _085698_, _085699_, _085700_, _085701_, _085702_, _085703_, _085704_, _085705_, _085706_, _085707_, _085708_, _085709_, _085710_, _085711_, _085712_, _085713_, _085714_, _085715_, _085716_, _085717_, _085718_, _085719_, _085720_, _085721_, _085722_, _085723_, _085724_, _085725_, _085726_, _085727_, _085728_, _085729_, _085730_, _085731_, _085732_, _085733_, _085734_, _085735_, _085736_, _085737_, _085738_, _085739_, _085740_, _085741_, _085742_, _085743_, _085744_, _085745_, _085746_, _085747_, _085748_, _085749_, _085750_, _085751_, _085752_, _085753_, _085754_, _085755_, _085756_, _085757_, _085758_, _085759_, _085760_, _085761_, _085762_, _085763_, _085764_, _085765_, _085766_, _085767_, _085768_, _085769_, _085770_, _085771_, _085772_, _085773_, _085774_, _085775_, _085776_, _085777_, _085778_, _085779_, _085780_, _085781_, _085782_, _085783_, _085784_, _085785_, _085786_, _085787_, _085788_, _085789_, _085790_, _085791_, _085792_, _085793_, _085794_, _085795_, _085796_, _085797_, _085798_, _085799_, _085800_, _085801_, _085802_, _085803_, _085804_, _085805_, _085806_, _085807_, _085808_, _085809_, _085810_, _085811_, _085812_, _085813_, _085814_, _085815_, _085816_, _085817_, _085818_, _085819_, _085820_, _085821_, _085822_, _085823_, _085824_, _085825_, _085826_, _085827_, _085828_, _085829_, _085830_, _085831_, _085832_, _085833_, _085834_, _085835_, _085836_, _085837_, _085838_, _085839_, _085840_, _085841_, _085842_, _085843_, _085844_, _085845_, _085846_, _085847_, _085848_, _085849_, _085850_, _085851_, _085852_, _085853_, _085854_, _085855_, _085856_, _085857_, _085858_, _085859_, _085860_, _085861_, _085862_, _085863_, _085864_, _085865_, _085866_, _085867_, _085868_, _085869_, _085870_, _085871_, _085872_, _085873_, _085874_, _085875_, _085876_, _085877_, _085878_, _085879_, _085880_, _085881_, _085882_, _085883_, _085884_, _085885_, _085886_, _085887_, _085888_, _085889_, _085890_, _085891_, _085892_, _085893_, _085894_, _085895_, _085896_, _085897_, _085898_, _085899_, _085900_, _085901_, _085902_, _085903_, _085904_, _085905_, _085906_, _085907_, _085908_, _085909_, _085910_, _085911_, _085912_, _085913_, _085914_, _085915_, _085916_, _085917_, _085918_, _085919_, _085920_, _085921_, _085922_, _085923_, _085924_, _085925_, _085926_, _085927_, _085928_, _085929_, _085930_, _085931_, _085932_, _085933_, _085934_, _085935_, _085936_, _085937_, _085938_, _085939_, _085940_, _085941_, _085942_, _085943_, _085944_, _085945_, _085946_, _085947_, _085948_, _085949_, _085950_, _085951_, _085952_, _085953_, _085954_, _085955_, _085956_, _085957_, _085958_, _085959_, _085960_, _085961_, _085962_, _085963_, _085964_, _085965_, _085966_, _085967_, _085968_, _085969_, _085970_, _085971_, _085972_, _085973_, _085974_, _085975_, _085976_, _085977_, _085978_, _085979_, _085980_, _085981_, _085982_, _085983_, _085984_, _085985_, _085986_, _085987_, _085988_, _085989_, _085990_, _085991_, _085992_, _085993_, _085994_, _085995_, _085996_, _085997_, _085998_, _085999_, _086000_, _086001_, _086002_, _086003_, _086004_, _086005_, _086006_, _086007_, _086008_, _086009_, _086010_, _086011_, _086012_, _086013_, _086014_, _086015_, _086016_, _086017_, _086018_, _086019_, _086020_, _086021_, _086022_, _086023_, _086024_, _086025_, _086026_, _086027_, _086028_, _086029_, _086030_, _086031_, _086032_, _086033_, _086034_, _086035_, _086036_, _086037_, _086038_, _086039_, _086040_, _086041_, _086042_, _086043_, _086044_, _086045_, _086046_, _086047_, _086048_, _086049_, _086050_, _086051_, _086052_, _086053_, _086054_, _086055_, _086056_, _086057_, _086058_, _086059_, _086060_, _086061_, _086062_, _086063_, _086064_, _086065_, _086066_, _086067_, _086068_, _086069_, _086070_, _086071_, _086072_, _086073_, _086074_, _086075_, _086076_, _086077_, _086078_, _086079_, _086080_, _086081_, _086082_, _086083_, _086084_, _086085_, _086086_, _086087_, _086088_, _086089_, _086090_, _086091_, _086092_, _086093_, _086094_, _086095_, _086096_, _086097_, _086098_, _086099_, _086100_, _086101_, _086102_, _086103_, _086104_, _086105_, _086106_, _086107_, _086108_, _086109_, _086110_, _086111_, _086112_, _086113_, _086114_, _086115_, _086116_, _086117_, _086118_, _086119_, _086120_, _086121_, _086122_, _086123_, _086124_, _086125_, _086126_, _086127_, _086128_, _086129_, _086130_, _086131_, _086132_, _086133_, _086134_, _086135_, _086136_, _086137_, _086138_, _086139_, _086140_, _086141_, _086142_, _086143_, _086144_, _086145_, _086146_, _086147_, _086148_, _086149_, _086150_, _086151_, _086152_, _086153_, _086154_, _086155_, _086156_, _086157_, _086158_, _086159_, _086160_, _086161_, _086162_, _086163_, _086164_, _086165_, _086166_, _086167_, _086168_, _086169_, _086170_, _086171_, _086172_, _086173_, _086174_, _086175_, _086176_, _086177_, _086178_, _086179_, _086180_, _086181_, _086182_, _086183_, _086184_, _086185_, _086186_, _086187_, _086188_, _086189_, _086190_, _086191_, _086192_, _086193_, _086194_, _086195_, _086196_, _086197_, _086198_, _086199_, _086200_, _086201_, _086202_, _086203_, _086204_, _086205_, _086206_, _086207_, _086208_, _086209_, _086210_, _086211_, _086212_, _086213_, _086214_, _086215_, _086216_, _086217_, _086218_, _086219_, _086220_, _086221_, _086222_, _086223_, _086224_, _086225_, _086226_, _086227_, _086228_, _086229_, _086230_, _086231_, _086232_, _086233_, _086234_, _086235_, _086236_, _086237_, _086238_, _086239_, _086240_, _086241_, _086242_, _086243_, _086244_, _086245_, _086246_, _086247_, _086248_, _086249_, _086250_, _086251_, _086252_, _086253_, _086254_, _086255_, _086256_, _086257_, _086258_, _086259_, _086260_, _086261_, _086262_, _086263_, _086264_, _086265_, _086266_, _086267_, _086268_, _086269_, _086270_, _086271_, _086272_, _086273_, _086274_, _086275_, _086276_, _086277_, _086278_, _086279_, _086280_, _086281_, _086282_, _086283_, _086284_, _086285_, _086286_, _086287_, _086288_, _086289_, _086290_, _086291_, _086292_, _086293_, _086294_, _086295_, _086296_, _086297_, _086298_, _086299_, _086300_, _086301_, _086302_, _086303_, _086304_, _086305_, _086306_, _086307_, _086308_, _086309_, _086310_, _086311_, _086312_, _086313_, _086314_, _086315_, _086316_, _086317_, _086318_, _086319_, _086320_, _086321_, _086322_, _086323_, _086324_, _086325_, _086326_, _086327_, _086328_, _086329_, _086330_, _086331_, _086332_, _086333_, _086334_, _086335_, _086336_, _086337_, _086338_, _086339_, _086340_, _086341_, _086342_, _086343_, _086344_, _086345_, _086346_, _086347_, _086348_, _086349_, _086350_, _086351_, _086352_, _086353_, _086354_, _086355_, _086356_, _086357_, _086358_, _086359_, _086360_, _086361_, _086362_, _086363_, _086364_, _086365_, _086366_, _086367_, _086368_, _086369_, _086370_, _086371_, _086372_, _086373_, _086374_, _086375_, _086376_, _086377_, _086378_, _086379_, _086380_, _086381_, _086382_, _086383_, _086384_, _086385_, _086386_, _086387_, _086388_, _086389_, _086390_, _086391_, _086392_, _086393_, _086394_, _086395_, _086396_, _086397_, _086398_, _086399_, _086400_, _086401_, _086402_, _086403_, _086404_, _086405_, _086406_, _086407_, _086408_, _086409_, _086410_, _086411_, _086412_, _086413_, _086414_, _086415_, _086416_, _086417_, _086418_, _086419_, _086420_, _086421_, _086422_, _086423_, _086424_, _086425_, _086426_, _086427_, _086428_, _086429_, _086430_, _086431_, _086432_, _086433_, _086434_, _086435_, _086436_, _086437_, _086438_, _086439_, _086440_, _086441_, _086442_, _086443_, _086444_, _086445_, _086446_, _086447_, _086448_, _086449_, _086450_, _086451_, _086452_, _086453_, _086454_, _086455_, _086456_, _086457_, _086458_, _086459_, _086460_, _086461_, _086462_, _086463_, _086464_, _086465_, _086466_, _086467_, _086468_, _086469_, _086470_, _086471_, _086472_, _086473_, _086474_, _086475_, _086476_, _086477_, _086478_, _086479_, _086480_, _086481_, _086482_, _086483_, _086484_, _086485_, _086486_, _086487_, _086488_, _086489_, _086490_, _086491_, _086492_, _086493_, _086494_, _086495_, _086496_, _086497_, _086498_, _086499_, _086500_, _086501_, _086502_, _086503_, _086504_, _086505_, _086506_, _086507_, _086508_, _086509_, _086510_, _086511_, _086512_, _086513_, _086514_, _086515_, _086516_, _086517_, _086518_, _086519_, _086520_, _086521_, _086522_, _086523_, _086524_, _086525_, _086526_, _086527_, _086528_, _086529_, _086530_, _086531_, _086532_, _086533_, _086534_, _086535_, _086536_, _086537_, _086538_, _086539_, _086540_, _086541_, _086542_, _086543_, _086544_, _086545_, _086546_, _086547_, _086548_, _086549_, _086550_, _086551_, _086552_, _086553_, _086554_, _086555_, _086556_, _086557_, _086558_, _086559_, _086560_, _086561_, _086562_, _086563_, _086564_, _086565_, _086566_, _086567_, _086568_, _086569_, _086570_, _086571_, _086572_, _086573_, _086574_, _086575_, _086576_, _086577_, _086578_, _086579_, _086580_, _086581_, _086582_, _086583_, _086584_, _086585_, _086586_, _086587_, _086588_, _086589_, _086590_, _086591_, _086592_, _086593_, _086594_, _086595_, _086596_, _086597_, _086598_, _086599_, _086600_, _086601_, _086602_, _086603_, _086604_, _086605_, _086606_, _086607_, _086608_, _086609_, _086610_, _086611_, _086612_, _086613_, _086614_, _086615_, _086616_, _086617_, _086618_, _086619_, _086620_, _086621_, _086622_, _086623_, _086624_, _086625_, _086626_, _086627_, _086628_, _086629_, _086630_, _086631_, _086632_, _086633_, _086634_, _086635_, _086636_, _086637_, _086638_, _086639_, _086640_, _086641_, _086642_, _086643_, _086644_, _086645_, _086646_, _086647_, _086648_, _086649_, _086650_, _086651_, _086652_, _086653_, _086654_, _086655_, _086656_, _086657_, _086658_, _086659_, _086660_, _086661_, _086662_, _086663_, _086664_, _086665_, _086666_, _086667_, _086668_, _086669_, _086670_, _086671_, _086672_, _086673_, _086674_, _086675_, _086676_, _086677_, _086678_, _086679_, _086680_, _086681_, _086682_, _086683_, _086684_, _086685_, _086686_, _086687_, _086688_, _086689_, _086690_, _086691_, _086692_, _086693_, _086694_, _086695_, _086696_, _086697_, _086698_, _086699_, _086700_, _086701_, _086702_, _086703_, _086704_, _086705_, _086706_, _086707_, _086708_, _086709_, _086710_, _086711_, _086712_, _086713_, _086714_, _086715_, _086716_, _086717_, _086718_, _086719_, _086720_, _086721_, _086722_, _086723_, _086724_, _086725_, _086726_, _086727_, _086728_, _086729_, _086730_, _086731_, _086732_, _086733_, _086734_, _086735_, _086736_, _086737_, _086738_, _086739_, _086740_, _086741_, _086742_, _086743_, _086744_, _086745_, _086746_, _086747_, _086748_, _086749_, _086750_, _086751_, _086752_, _086753_, _086754_, _086755_, _086756_, _086757_, _086758_, _086759_, _086760_, _086761_, _086762_, _086763_, _086764_, _086765_, _086766_, _086767_, _086768_, _086769_, _086770_, _086771_, _086772_, _086773_, _086774_, _086775_, _086776_, _086777_, _086778_, _086779_, _086780_, _086781_, _086782_, _086783_, _086784_, _086785_, _086786_, _086787_, _086788_, _086789_, _086790_, _086791_, _086792_, _086793_, _086794_, _086795_, _086796_, _086797_, _086798_, _086799_, _086800_, _086801_, _086802_, _086803_, _086804_, _086805_, _086806_, _086807_, _086808_, _086809_, _086810_, _086811_, _086812_, _086813_, _086814_, _086815_, _086816_, _086817_, _086818_, _086819_, _086820_, _086821_, _086822_, _086823_, _086824_, _086825_, _086826_, _086827_, _086828_, _086829_, _086830_, _086831_, _086832_, _086833_, _086834_, _086835_, _086836_, _086837_, _086838_, _086839_, _086840_, _086841_, _086842_, _086843_, _086844_, _086845_, _086846_, _086847_, _086848_, _086849_, _086850_, _086851_, _086852_, _086853_, _086854_, _086855_, _086856_, _086857_, _086858_, _086859_, _086860_, _086861_, _086862_, _086863_, _086864_, _086865_, _086866_, _086867_, _086868_, _086869_, _086870_, _086871_, _086872_, _086873_, _086874_, _086875_, _086876_, _086877_, _086878_, _086879_, _086880_, _086881_, _086882_, _086883_, _086884_, _086885_, _086886_, _086887_, _086888_, _086889_, _086890_, _086891_, _086892_, _086893_, _086894_, _086895_, _086896_, _086897_, _086898_, _086899_, _086900_, _086901_, _086902_, _086903_, _086904_, _086905_, _086906_, _086907_, _086908_, _086909_, _086910_, _086911_, _086912_, _086913_, _086914_, _086915_, _086916_, _086917_, _086918_, _086919_, _086920_, _086921_, _086922_, _086923_, _086924_, _086925_, _086926_, _086927_, _086928_, _086929_, _086930_, _086931_, _086932_, _086933_, _086934_, _086935_, _086936_, _086937_, _086938_, _086939_, _086940_, _086941_, _086942_, _086943_, _086944_, _086945_, _086946_, _086947_, _086948_, _086949_, _086950_, _086951_, _086952_, _086953_, _086954_, _086955_, _086956_, _086957_, _086958_, _086959_, _086960_, _086961_, _086962_, _086963_, _086964_, _086965_, _086966_, _086967_, _086968_, _086969_, _086970_, _086971_, _086972_, _086973_, _086974_, _086975_, _086976_, _086977_, _086978_, _086979_, _086980_, _086981_, _086982_, _086983_, _086984_, _086985_, _086986_, _086987_, _086988_, _086989_, _086990_, _086991_, _086992_, _086993_, _086994_, _086995_, _086996_, _086997_, _086998_, _086999_, _087000_, _087001_, _087002_, _087003_, _087004_, _087005_, _087006_, _087007_, _087008_, _087009_, _087010_, _087011_, _087012_, _087013_, _087014_, _087015_, _087016_, _087017_, _087018_, _087019_, _087020_, _087021_, _087022_, _087023_, _087024_, _087025_, _087026_, _087027_, _087028_, _087029_, _087030_, _087031_, _087032_, _087033_, _087034_, _087035_, _087036_, _087037_, _087038_, _087039_, _087040_, _087041_, _087042_, _087043_, _087044_, _087045_, _087046_, _087047_, _087048_, _087049_, _087050_, _087051_, _087052_, _087053_, _087054_, _087055_, _087056_, _087057_, _087058_, _087059_, _087060_, _087061_, _087062_, _087063_, _087064_, _087065_, _087066_, _087067_, _087068_, _087069_, _087070_, _087071_, _087072_, _087073_, _087074_, _087075_, _087076_, _087077_, _087078_, _087079_, _087080_, _087081_, _087082_, _087083_, _087084_, _087085_, _087086_, _087087_, _087088_, _087089_, _087090_, _087091_, _087092_, _087093_, _087094_, _087095_, _087096_, _087097_, _087098_, _087099_, _087100_, _087101_, _087102_, _087103_, _087104_, _087105_, _087106_, _087107_, _087108_, _087109_, _087110_, _087111_, _087112_, _087113_, _087114_, _087115_, _087116_, _087117_, _087118_, _087119_, _087120_, _087121_, _087122_, _087123_, _087124_, _087125_, _087126_, _087127_, _087128_, _087129_, _087130_, _087131_, _087132_, _087133_, _087134_, _087135_, _087136_, _087137_, _087138_, _087139_, _087140_, _087141_, _087142_, _087143_, _087144_, _087145_, _087146_, _087147_, _087148_, _087149_, _087150_, _087151_, _087152_, _087153_, _087154_, _087155_, _087156_, _087157_, _087158_, _087159_, _087160_, _087161_, _087162_, _087163_, _087164_, _087165_, _087166_, _087167_, _087168_, _087169_, _087170_, _087171_, _087172_, _087173_, _087174_, _087175_, _087176_, _087177_, _087178_, _087179_, _087180_, _087181_, _087182_, _087183_, _087184_, _087185_, _087186_, _087187_, _087188_, _087189_, _087190_, _087191_, _087192_, _087193_, _087194_, _087195_, _087196_, _087197_, _087198_, _087199_, _087200_, _087201_, _087202_, _087203_, _087204_, _087205_, _087206_, _087207_, _087208_, _087209_, _087210_, _087211_, _087212_, _087213_, _087214_, _087215_, _087216_, _087217_, _087218_, _087219_, _087220_, _087221_, _087222_, _087223_, _087224_, _087225_, _087226_, _087227_, _087228_, _087229_, _087230_, _087231_, _087232_, _087233_, _087234_, _087235_, _087236_, _087237_, _087238_, _087239_, _087240_, _087241_, _087242_, _087243_, _087244_, _087245_, _087246_, _087247_, _087248_, _087249_, _087250_, _087251_, _087252_, _087253_, _087254_, _087255_, _087256_, _087257_, _087258_, _087259_, _087260_, _087261_, _087262_, _087263_, _087264_, _087265_, _087266_, _087267_, _087268_, _087269_, _087270_, _087271_, _087272_, _087273_, _087274_, _087275_, _087276_, _087277_, _087278_, _087279_, _087280_, _087281_, _087282_, _087283_, _087284_, _087285_, _087286_, _087287_, _087288_, _087289_, _087290_, _087291_, _087292_, _087293_, _087294_, _087295_, _087296_, _087297_, _087298_, _087299_, _087300_, _087301_, _087302_, _087303_, _087304_, _087305_, _087306_, _087307_, _087308_, _087309_, _087310_, _087311_, _087312_, _087313_, _087314_, _087315_, _087316_, _087317_, _087318_, _087319_, _087320_, _087321_, _087322_, _087323_, _087324_, _087325_, _087326_, _087327_, _087328_, _087329_, _087330_, _087331_, _087332_, _087333_, _087334_, _087335_, _087336_, _087337_, _087338_, _087339_, _087340_, _087341_, _087342_, _087343_, _087344_, _087345_, _087346_, _087347_, _087348_, _087349_, _087350_, _087351_, _087352_, _087353_, _087354_, _087355_, _087356_, _087357_, _087358_, _087359_, _087360_, _087361_, _087362_, _087363_, _087364_, _087365_, _087366_, _087367_, _087368_, _087369_, _087370_, _087371_, _087372_, _087373_, _087374_, _087375_, _087376_, _087377_, _087378_, _087379_, _087380_, _087381_, _087382_, _087383_, _087384_, _087385_, _087386_, _087387_, _087388_, _087389_, _087390_, _087391_, _087392_, _087393_, _087394_, _087395_, _087396_, _087397_, _087398_, _087399_, _087400_, _087401_, _087402_, _087403_, _087404_, _087405_, _087406_, _087407_, _087408_, _087409_, _087410_, _087411_, _087412_, _087413_, _087414_, _087415_, _087416_, _087417_, _087418_, _087419_, _087420_, _087421_, _087422_, _087423_, _087424_, _087425_, _087426_, _087427_, _087428_, _087429_, _087430_, _087431_, _087432_, _087433_, _087434_, _087435_, _087436_, _087437_, _087438_, _087439_, _087440_, _087441_, _087442_, _087443_, _087444_, _087445_, _087446_, _087447_, _087448_, _087449_, _087450_, _087451_, _087452_, _087453_, _087454_, _087455_, _087456_, _087457_, _087458_, _087459_, _087460_, _087461_, _087462_, _087463_, _087464_, _087465_, _087466_, _087467_, _087468_, _087469_, _087470_, _087471_, _087472_, _087473_, _087474_, _087475_, _087476_, _087477_, _087478_, _087479_, _087480_, _087481_, _087482_, _087483_, _087484_, _087485_, _087486_, _087487_, _087488_, _087489_, _087490_, _087491_, _087492_, _087493_, _087494_, _087495_, _087496_, _087497_, _087498_, _087499_, _087500_, _087501_, _087502_, _087503_, _087504_, _087505_, _087506_, _087507_, _087508_, _087509_, _087510_, _087511_, _087512_, _087513_, _087514_, _087515_, _087516_, _087517_, _087518_, _087519_, _087520_, _087521_, _087522_, _087523_, _087524_, _087525_, _087526_, _087527_, _087528_, _087529_, _087530_, _087531_, _087532_, _087533_, _087534_, _087535_, _087536_, _087537_, _087538_, _087539_, _087540_, _087541_, _087542_, _087543_, _087544_, _087545_, _087546_, _087547_, _087548_, _087549_, _087550_, _087551_, _087552_, _087553_, _087554_, _087555_, _087556_, _087557_, _087558_, _087559_, _087560_, _087561_, _087562_, _087563_, _087564_, _087565_, _087566_, _087567_, _087568_, _087569_, _087570_, _087571_, _087572_, _087573_, _087574_, _087575_, _087576_, _087577_, _087578_, _087579_, _087580_, _087581_, _087582_, _087583_, _087584_, _087585_, _087586_, _087587_, _087588_, _087589_, _087590_, _087591_, _087592_, _087593_, _087594_, _087595_, _087596_, _087597_, _087598_, _087599_, _087600_, _087601_, _087602_, _087603_, _087604_, _087605_, _087606_, _087607_, _087608_, _087609_, _087610_, _087611_, _087612_, _087613_, _087614_, _087615_, _087616_, _087617_, _087618_, _087619_, _087620_, _087621_, _087622_, _087623_, _087624_, _087625_, _087626_, _087627_, _087628_, _087629_, _087630_, _087631_, _087632_, _087633_, _087634_, _087635_, _087636_, _087637_, _087638_, _087639_, _087640_, _087641_, _087642_, _087643_, _087644_, _087645_, _087646_, _087647_, _087648_, _087649_, _087650_, _087651_, _087652_, _087653_, _087654_, _087655_, _087656_, _087657_, _087658_, _087659_, _087660_, _087661_, _087662_, _087663_, _087664_, _087665_, _087666_, _087667_, _087668_, _087669_, _087670_, _087671_, _087672_, _087673_, _087674_, _087675_, _087676_, _087677_, _087678_, _087679_, _087680_, _087681_, _087682_, _087683_, _087684_, _087685_, _087686_, _087687_, _087688_, _087689_, _087690_, _087691_, _087692_, _087693_, _087694_, _087695_, _087696_, _087697_, _087698_, _087699_, _087700_, _087701_, _087702_, _087703_, _087704_, _087705_, _087706_, _087707_, _087708_, _087709_, _087710_, _087711_, _087712_, _087713_, _087714_, _087715_, _087716_, _087717_, _087718_, _087719_, _087720_, _087721_, _087722_, _087723_, _087724_, _087725_, _087726_, _087727_, _087728_, _087729_, _087730_, _087731_, _087732_, _087733_, _087734_, _087735_, _087736_, _087737_, _087738_, _087739_, _087740_, _087741_, _087742_, _087743_, _087744_, _087745_, _087746_, _087747_, _087748_, _087749_, _087750_, _087751_, _087752_, _087753_, _087754_, _087755_, _087756_, _087757_, _087758_, _087759_, _087760_, _087761_, _087762_, _087763_, _087764_, _087765_, _087766_, _087767_, _087768_, _087769_, _087770_, _087771_, _087772_, _087773_, _087774_, _087775_, _087776_, _087777_, _087778_, _087779_, _087780_, _087781_, _087782_, _087783_, _087784_, _087785_, _087786_, _087787_, _087788_, _087789_, _087790_, _087791_, _087792_, _087793_, _087794_, _087795_, _087796_, _087797_, _087798_, _087799_, _087800_, _087801_, _087802_, _087803_, _087804_, _087805_, _087806_, _087807_, _087808_, _087809_, _087810_, _087811_, _087812_, _087813_, _087814_, _087815_, _087816_, _087817_, _087818_, _087819_, _087820_, _087821_, _087822_, _087823_, _087824_, _087825_, _087826_, _087827_, _087828_, _087829_, _087830_, _087831_, _087832_, _087833_, _087834_, _087835_, _087836_, _087837_, _087838_, _087839_, _087840_, _087841_, _087842_, _087843_, _087844_, _087845_, _087846_, _087847_, _087848_, _087849_, _087850_, _087851_, _087852_, _087853_, _087854_, _087855_, _087856_, _087857_, _087858_, _087859_, _087860_, _087861_, _087862_, _087863_, _087864_, _087865_, _087866_, _087867_, _087868_, _087869_, _087870_, _087871_, _087872_, _087873_, _087874_, _087875_, _087876_, _087877_, _087878_, _087879_, _087880_, _087881_, _087882_, _087883_, _087884_, _087885_, _087886_, _087887_, _087888_, _087889_, _087890_, _087891_, _087892_, _087893_, _087894_, _087895_, _087896_, _087897_, _087898_, _087899_, _087900_, _087901_, _087902_, _087903_, _087904_, _087905_, _087906_, _087907_, _087908_, _087909_, _087910_, _087911_, _087912_, _087913_, _087914_, _087915_, _087916_, _087917_, _087918_, _087919_, _087920_, _087921_, _087922_, _087923_, _087924_, _087925_, _087926_, _087927_, _087928_, _087929_, _087930_, _087931_, _087932_, _087933_, _087934_, _087935_, _087936_, _087937_, _087938_, _087939_, _087940_, _087941_, _087942_, _087943_, _087944_, _087945_, _087946_, _087947_, _087948_, _087949_, _087950_, _087951_, _087952_, _087953_, _087954_, _087955_, _087956_, _087957_, _087958_, _087959_, _087960_, _087961_, _087962_, _087963_, _087964_, _087965_, _087966_, _087967_, _087968_, _087969_, _087970_, _087971_, _087972_, _087973_, _087974_, _087975_, _087976_, _087977_, _087978_, _087979_, _087980_, _087981_, _087982_, _087983_, _087984_, _087985_, _087986_, _087987_, _087988_, _087989_, _087990_, _087991_, _087992_, _087993_, _087994_, _087995_, _087996_, _087997_, _087998_, _087999_, _088000_, _088001_, _088002_, _088003_, _088004_, _088005_, _088006_, _088007_, _088008_, _088009_, _088010_, _088011_, _088012_, _088013_, _088014_, _088015_, _088016_, _088017_, _088018_, _088019_, _088020_, _088021_, _088022_, _088023_, _088024_, _088025_, _088026_, _088027_, _088028_, _088029_, _088030_, _088031_, _088032_, _088033_, _088034_, _088035_, _088036_, _088037_, _088038_, _088039_, _088040_, _088041_, _088042_, _088043_, _088044_, _088045_, _088046_, _088047_, _088048_, _088049_, _088050_, _088051_, _088052_, _088053_, _088054_, _088055_, _088056_, _088057_, _088058_, _088059_, _088060_, _088061_, _088062_, _088063_, _088064_, _088065_, _088066_, _088067_, _088068_, _088069_, _088070_, _088071_, _088072_, _088073_, _088074_, _088075_, _088076_, _088077_, _088078_, _088079_, _088080_, _088081_, _088082_, _088083_, _088084_, _088085_, _088086_, _088087_, _088088_, _088089_, _088090_, _088091_, _088092_, _088093_, _088094_, _088095_, _088096_, _088097_, _088098_, _088099_, _088100_, _088101_, _088102_, _088103_, _088104_, _088105_, _088106_, _088107_, _088108_, _088109_, _088110_, _088111_, _088112_, _088113_, _088114_, _088115_, _088116_, _088117_, _088118_, _088119_, _088120_, _088121_, _088122_, _088123_, _088124_, _088125_, _088126_, _088127_, _088128_, _088129_, _088130_, _088131_, _088132_, _088133_, _088134_, _088135_, _088136_, _088137_, _088138_, _088139_, _088140_, _088141_, _088142_, _088143_, _088144_, _088145_, _088146_, _088147_, _088148_, _088149_, _088150_, _088151_, _088152_, _088153_, _088154_, _088155_, _088156_, _088157_, _088158_, _088159_, _088160_, _088161_, _088162_, _088163_, _088164_, _088165_, _088166_, _088167_, _088168_, _088169_, _088170_, _088171_, _088172_, _088173_, _088174_, _088175_, _088176_, _088177_, _088178_, _088179_, _088180_, _088181_, _088182_, _088183_, _088184_, _088185_, _088186_, _088187_, _088188_, _088189_, _088190_, _088191_, _088192_, _088193_, _088194_, _088195_, _088196_, _088197_, _088198_, _088199_, _088200_, _088201_, _088202_, _088203_, _088204_, _088205_, _088206_, _088207_, _088208_, _088209_, _088210_, _088211_, _088212_, _088213_, _088214_, _088215_, _088216_, _088217_, _088218_, _088219_, _088220_, _088221_, _088222_, _088223_, _088224_, _088225_, _088226_, _088227_, _088228_, _088229_, _088230_, _088231_, _088232_, _088233_, _088234_, _088235_, _088236_, _088237_, _088238_, _088239_, _088240_, _088241_, _088242_, _088243_, _088244_, _088245_, _088246_, _088247_, _088248_, _088249_, _088250_, _088251_, _088252_, _088253_, _088254_, _088255_, _088256_, _088257_, _088258_, _088259_, _088260_, _088261_, _088262_, _088263_, _088264_, _088265_, _088266_, _088267_, _088268_, _088269_, _088270_, _088271_, _088272_, _088273_, _088274_, _088275_, _088276_, _088277_, _088278_, _088279_, _088280_, _088281_, _088282_, _088283_, _088284_, _088285_, _088286_, _088287_, _088288_, _088289_, _088290_, _088291_, _088292_, _088293_, _088294_, _088295_, _088296_, _088297_, _088298_, _088299_, _088300_, _088301_, _088302_, _088303_, _088304_, _088305_, _088306_, _088307_, _088308_, _088309_, _088310_, _088311_, _088312_, _088313_, _088314_, _088315_, _088316_, _088317_, _088318_, _088319_, _088320_, _088321_, _088322_, _088323_, _088324_, _088325_, _088326_, _088327_, _088328_, _088329_, _088330_, _088331_, _088332_, _088333_, _088334_, _088335_, _088336_, _088337_, _088338_, _088339_, _088340_, _088341_, _088342_, _088343_, _088344_, _088345_, _088346_, _088347_, _088348_, _088349_, _088350_, _088351_, _088352_, _088353_, _088354_, _088355_, _088356_, _088357_, _088358_, _088359_, _088360_, _088361_, _088362_, _088363_, _088364_, _088365_, _088366_, _088367_, _088368_, _088369_, _088370_, _088371_, _088372_, _088373_, _088374_, _088375_, _088376_, _088377_, _088378_, _088379_, _088380_, _088381_, _088382_, _088383_, _088384_, _088385_, _088386_, _088387_, _088388_, _088389_, _088390_, _088391_, _088392_, _088393_, _088394_, _088395_, _088396_, _088397_, _088398_, _088399_, _088400_, _088401_, _088402_, _088403_, _088404_, _088405_, _088406_, _088407_, _088408_, _088409_, _088410_, _088411_, _088412_, _088413_, _088414_, _088415_, _088416_, _088417_, _088418_, _088419_, _088420_, _088421_, _088422_, _088423_, _088424_, _088425_, _088426_, _088427_, _088428_, _088429_, _088430_, _088431_, _088432_, _088433_, _088434_, _088435_, _088436_, _088437_, _088438_, _088439_, _088440_, _088441_, _088442_, _088443_, _088444_, _088445_, _088446_, _088447_, _088448_, _088449_, _088450_, _088451_, _088452_, _088453_, _088454_, _088455_, _088456_, _088457_, _088458_, _088459_, _088460_, _088461_, _088462_, _088463_, _088464_, _088465_, _088466_, _088467_, _088468_, _088469_, _088470_, _088471_, _088472_, _088473_, _088474_, _088475_, _088476_, _088477_, _088478_, _088479_, _088480_, _088481_, _088482_, _088483_, _088484_, _088485_, _088486_, _088487_, _088488_, _088489_, _088490_, _088491_, _088492_, _088493_, _088494_, _088495_, _088496_, _088497_, _088498_, _088499_, _088500_, _088501_, _088502_, _088503_, _088504_, _088505_, _088506_, _088507_, _088508_, _088509_, _088510_, _088511_, _088512_, _088513_, _088514_, _088515_, _088516_, _088517_, _088518_, _088519_, _088520_, _088521_, _088522_, _088523_, _088524_, _088525_, _088526_, _088527_, _088528_, _088529_, _088530_, _088531_, _088532_, _088533_, _088534_, _088535_, _088536_, _088537_, _088538_, _088539_, _088540_, _088541_, _088542_, _088543_, _088544_, _088545_, _088546_, _088547_, _088548_, _088549_, _088550_, _088551_, _088552_, _088553_, _088554_, _088555_, _088556_, _088557_, _088558_, _088559_, _088560_, _088561_, _088562_, _088563_, _088564_, _088565_, _088566_, _088567_, _088568_, _088569_, _088570_, _088571_, _088572_, _088573_, _088574_, _088575_, _088576_, _088577_, _088578_, _088579_, _088580_, _088581_, _088582_, _088583_, _088584_, _088585_, _088586_, _088587_, _088588_, _088589_, _088590_, _088591_, _088592_, _088593_, _088594_, _088595_, _088596_, _088597_, _088598_, _088599_, _088600_, _088601_, _088602_, _088603_, _088604_, _088605_, _088606_, _088607_, _088608_, _088609_, _088610_, _088611_, _088612_, _088613_, _088614_, _088615_, _088616_, _088617_, _088618_, _088619_, _088620_, _088621_, _088622_, _088623_, _088624_, _088625_, _088626_, _088627_, _088628_, _088629_, _088630_, _088631_, _088632_, _088633_, _088634_, _088635_, _088636_, _088637_, _088638_, _088639_, _088640_, _088641_, _088642_, _088643_, _088644_, _088645_, _088646_, _088647_, _088648_, _088649_, _088650_, _088651_, _088652_, _088653_, _088654_, _088655_, _088656_, _088657_, _088658_, _088659_, _088660_, _088661_, _088662_, _088663_, _088664_, _088665_, _088666_, _088667_, _088668_, _088669_, _088670_, _088671_, _088672_, _088673_, _088674_, _088675_, _088676_, _088677_, _088678_, _088679_, _088680_, _088681_, _088682_, _088683_, _088684_, _088685_, _088686_, _088687_, _088688_, _088689_, _088690_, _088691_, _088692_, _088693_, _088694_, _088695_, _088696_, _088697_, _088698_, _088699_, _088700_, _088701_, _088702_, _088703_, _088704_, _088705_, _088706_, _088707_, _088708_, _088709_, _088710_, _088711_, _088712_, _088713_, _088714_, _088715_, _088716_, _088717_, _088718_, _088719_, _088720_, _088721_, _088722_, _088723_, _088724_, _088725_, _088726_, _088727_, _088728_, _088729_, _088730_, _088731_, _088732_, _088733_, _088734_, _088735_, _088736_, _088737_, _088738_, _088739_, _088740_, _088741_, _088742_, _088743_, _088744_, _088745_, _088746_, _088747_, _088748_, _088749_, _088750_, _088751_, _088752_, _088753_, _088754_, _088755_, _088756_, _088757_, _088758_, _088759_, _088760_, _088761_, _088762_, _088763_, _088764_, _088765_, _088766_, _088767_, _088768_, _088769_, _088770_, _088771_, _088772_, _088773_, _088774_, _088775_, _088776_, _088777_, _088778_, _088779_, _088780_, _088781_, _088782_, _088783_, _088784_, _088785_, _088786_, _088787_, _088788_, _088789_, _088790_, _088791_, _088792_, _088793_, _088794_, _088795_, _088796_, _088797_, _088798_, _088799_, _088800_, _088801_, _088802_, _088803_, _088804_, _088805_, _088806_, _088807_, _088808_, _088809_, _088810_, _088811_, _088812_, _088813_, _088814_, _088815_, _088816_, _088817_, _088818_, _088819_, _088820_, _088821_, _088822_, _088823_, _088824_, _088825_, _088826_, _088827_, _088828_, _088829_, _088830_, _088831_, _088832_, _088833_, _088834_, _088835_, _088836_, _088837_, _088838_, _088839_, _088840_, _088841_, _088842_, _088843_, _088844_, _088845_, _088846_, _088847_, _088848_, _088849_, _088850_, _088851_, _088852_, _088853_, _088854_, _088855_, _088856_, _088857_, _088858_, _088859_, _088860_, _088861_, _088862_, _088863_, _088864_, _088865_, _088866_, _088867_, _088868_, _088869_, _088870_, _088871_, _088872_, _088873_, _088874_, _088875_, _088876_, _088877_, _088878_, _088879_, _088880_, _088881_, _088882_, _088883_, _088884_, _088885_, _088886_, _088887_, _088888_, _088889_, _088890_, _088891_, _088892_, _088893_, _088894_, _088895_, _088896_, _088897_, _088898_, _088899_, _088900_, _088901_, _088902_, _088903_, _088904_, _088905_, _088906_, _088907_, _088908_, _088909_, _088910_, _088911_, _088912_, _088913_, _088914_, _088915_, _088916_, _088917_, _088918_, _088919_, _088920_, _088921_, _088922_, _088923_, _088924_, _088925_, _088926_, _088927_, _088928_, _088929_, _088930_, _088931_, _088932_, _088933_, _088934_, _088935_, _088936_, _088937_, _088938_, _088939_, _088940_, _088941_, _088942_, _088943_, _088944_, _088945_, _088946_, _088947_, _088948_, _088949_, _088950_, _088951_, _088952_, _088953_, _088954_, _088955_, _088956_, _088957_, _088958_, _088959_, _088960_, _088961_, _088962_, _088963_, _088964_, _088965_, _088966_, _088967_, _088968_, _088969_, _088970_, _088971_, _088972_, _088973_, _088974_, _088975_, _088976_, _088977_, _088978_, _088979_, _088980_, _088981_, _088982_, _088983_, _088984_, _088985_, _088986_, _088987_, _088988_, _088989_, _088990_, _088991_, _088992_, _088993_, _088994_, _088995_, _088996_, _088997_, _088998_, _088999_, _089000_, _089001_, _089002_, _089003_, _089004_, _089005_, _089006_, _089007_, _089008_, _089009_, _089010_, _089011_, _089012_, _089013_, _089014_, _089015_, _089016_, _089017_, _089018_, _089019_, _089020_, _089021_, _089022_, _089023_, _089024_, _089025_, _089026_, _089027_, _089028_, _089029_, _089030_, _089031_, _089032_, _089033_, _089034_, _089035_, _089036_, _089037_, _089038_, _089039_, _089040_, _089041_, _089042_, _089043_, _089044_, _089045_, _089046_, _089047_, _089048_, _089049_, _089050_, _089051_, _089052_, _089053_, _089054_, _089055_, _089056_, _089057_, _089058_, _089059_, _089060_, _089061_, _089062_, _089063_, _089064_, _089065_, _089066_, _089067_, _089068_, _089069_, _089070_, _089071_, _089072_, _089073_, _089074_, _089075_, _089076_, _089077_, _089078_, _089079_, _089080_, _089081_, _089082_, _089083_, _089084_, _089085_, _089086_, _089087_, _089088_, _089089_, _089090_, _089091_, _089092_, _089093_, _089094_, _089095_, _089096_, _089097_, _089098_, _089099_, _089100_, _089101_, _089102_, _089103_, _089104_, _089105_, _089106_, _089107_, _089108_, _089109_, _089110_, _089111_, _089112_, _089113_, _089114_, _089115_, _089116_, _089117_, _089118_, _089119_, _089120_, _089121_, _089122_, _089123_, _089124_, _089125_, _089126_, _089127_, _089128_, _089129_, _089130_, _089131_, _089132_, _089133_, _089134_, _089135_, _089136_, _089137_, _089138_, _089139_, _089140_, _089141_, _089142_, _089143_, _089144_, _089145_, _089146_, _089147_, _089148_, _089149_, _089150_, _089151_, _089152_, _089153_, _089154_, _089155_, _089156_, _089157_, _089158_, _089159_, _089160_, _089161_, _089162_, _089163_, _089164_, _089165_, _089166_, _089167_, _089168_, _089169_, _089170_, _089171_, _089172_, _089173_, _089174_, _089175_, _089176_, _089177_, _089178_, _089179_, _089180_, _089181_, _089182_, _089183_, _089184_, _089185_, _089186_, _089187_, _089188_, _089189_, _089190_, _089191_, _089192_, _089193_, _089194_, _089195_, _089196_, _089197_, _089198_, _089199_, _089200_, _089201_, _089202_, _089203_, _089204_, _089205_, _089206_, _089207_, _089208_, _089209_, _089210_, _089211_, _089212_, _089213_, _089214_, _089215_, _089216_, _089217_, _089218_, _089219_, _089220_, _089221_, _089222_, _089223_, _089224_, _089225_, _089226_, _089227_, _089228_, _089229_, _089230_, _089231_, _089232_, _089233_, _089234_, _089235_, _089236_, _089237_, _089238_, _089239_, _089240_, _089241_, _089242_, _089243_, _089244_, _089245_, _089246_, _089247_, _089248_, _089249_, _089250_, _089251_, _089252_, _089253_, _089254_, _089255_, _089256_, _089257_, _089258_, _089259_, _089260_, _089261_, _089262_, _089263_, _089264_, _089265_, _089266_, _089267_, _089268_, _089269_, _089270_, _089271_, _089272_, _089273_, _089274_, _089275_, _089276_, _089277_, _089278_, _089279_, _089280_, _089281_, _089282_, _089283_, _089284_, _089285_, _089286_, _089287_, _089288_, _089289_, _089290_, _089291_, _089292_, _089293_, _089294_, _089295_, _089296_, _089297_, _089298_, _089299_, _089300_, _089301_, _089302_, _089303_, _089304_, _089305_, _089306_, _089307_, _089308_, _089309_, _089310_, _089311_, _089312_, _089313_, _089314_, _089315_, _089316_, _089317_, _089318_, _089319_, _089320_, _089321_, _089322_, _089323_, _089324_, _089325_, _089326_, _089327_, _089328_, _089329_, _089330_, _089331_, _089332_, _089333_, _089334_, _089335_, _089336_, _089337_, _089338_, _089339_, _089340_, _089341_, _089342_, _089343_, _089344_, _089345_, _089346_, _089347_, _089348_, _089349_, _089350_, _089351_, _089352_, _089353_, _089354_, _089355_, _089356_, _089357_, _089358_, _089359_, _089360_, _089361_, _089362_, _089363_, _089364_, _089365_, _089366_, _089367_, _089368_, _089369_, _089370_, _089371_, _089372_, _089373_, _089374_, _089375_, _089376_, _089377_, _089378_, _089379_, _089380_, _089381_, _089382_, _089383_, _089384_, _089385_, _089386_, _089387_, _089388_, _089389_, _089390_, _089391_, _089392_, _089393_, _089394_, _089395_, _089396_, _089397_, _089398_, _089399_, _089400_, _089401_, _089402_, _089403_, _089404_, _089405_, _089406_, _089407_, _089408_, _089409_, _089410_, _089411_, _089412_, _089413_, _089414_, _089415_, _089416_, _089417_, _089418_, _089419_, _089420_, _089421_, _089422_, _089423_, _089424_, _089425_, _089426_, _089427_, _089428_, _089429_, _089430_, _089431_, _089432_, _089433_, _089434_, _089435_, _089436_, _089437_, _089438_, _089439_, _089440_, _089441_, _089442_, _089443_, _089444_, _089445_, _089446_, _089447_, _089448_, _089449_, _089450_, _089451_, _089452_, _089453_, _089454_, _089455_, _089456_, _089457_, _089458_, _089459_, _089460_, _089461_, _089462_, _089463_, _089464_, _089465_, _089466_, _089467_, _089468_, _089469_, _089470_, _089471_, _089472_, _089473_, _089474_, _089475_, _089476_, _089477_, _089478_, _089479_, _089480_, _089481_, _089482_, _089483_, _089484_, _089485_, _089486_, _089487_, _089488_, _089489_, _089490_, _089491_, _089492_, _089493_, _089494_, _089495_, _089496_, _089497_, _089498_, _089499_, _089500_, _089501_, _089502_, _089503_, _089504_, _089505_, _089506_, _089507_, _089508_, _089509_, _089510_, _089511_, _089512_, _089513_, _089514_, _089515_, _089516_, _089517_, _089518_, _089519_, _089520_, _089521_, _089522_, _089523_, _089524_, _089525_, _089526_, _089527_, _089528_, _089529_, _089530_, _089531_, _089532_, _089533_, _089534_, _089535_, _089536_, _089537_, _089538_, _089539_, _089540_, _089541_, _089542_, _089543_, _089544_, _089545_, _089546_, _089547_, _089548_, _089549_, _089550_, _089551_, _089552_, _089553_, _089554_, _089555_, _089556_, _089557_, _089558_, _089559_, _089560_, _089561_, _089562_, _089563_, _089564_, _089565_, _089566_, _089567_, _089568_, _089569_, _089570_, _089571_, _089572_, _089573_, _089574_, _089575_, _089576_, _089577_, _089578_, _089579_, _089580_, _089581_, _089582_, _089583_, _089584_, _089585_, _089586_, _089587_, _089588_, _089589_, _089590_, _089591_, _089592_, _089593_, _089594_, _089595_, _089596_, _089597_, _089598_, _089599_, _089600_, _089601_, _089602_, _089603_, _089604_, _089605_, _089606_, _089607_, _089608_, _089609_, _089610_, _089611_, _089612_, _089613_, _089614_, _089615_, _089616_, _089617_, _089618_, _089619_, _089620_, _089621_, _089622_, _089623_, _089624_, _089625_, _089626_, _089627_, _089628_, _089629_, _089630_, _089631_, _089632_, _089633_, _089634_, _089635_, _089636_, _089637_, _089638_, _089639_, _089640_, _089641_, _089642_, _089643_, _089644_, _089645_, _089646_, _089647_, _089648_, _089649_, _089650_, _089651_, _089652_, _089653_, _089654_, _089655_, _089656_, _089657_, _089658_, _089659_, _089660_, _089661_, _089662_, _089663_, _089664_, _089665_, _089666_, _089667_, _089668_, _089669_, _089670_, _089671_, _089672_, _089673_, _089674_, _089675_, _089676_, _089677_, _089678_, _089679_, _089680_, _089681_, _089682_, _089683_, _089684_, _089685_, _089686_, _089687_, _089688_, _089689_, _089690_, _089691_, _089692_, _089693_, _089694_, _089695_, _089696_, _089697_, _089698_, _089699_, _089700_, _089701_, _089702_, _089703_, _089704_, _089705_, _089706_, _089707_, _089708_, _089709_, _089710_, _089711_, _089712_, _089713_, _089714_, _089715_, _089716_, _089717_, _089718_, _089719_, _089720_, _089721_, _089722_, _089723_, _089724_, _089725_, _089726_, _089727_, _089728_, _089729_, _089730_, _089731_, _089732_, _089733_, _089734_, _089735_, _089736_, _089737_, _089738_, _089739_, _089740_, _089741_, _089742_, _089743_, _089744_, _089745_, _089746_, _089747_, _089748_, _089749_, _089750_, _089751_, _089752_, _089753_, _089754_, _089755_, _089756_, _089757_, _089758_, _089759_, _089760_, _089761_, _089762_, _089763_, _089764_, _089765_, _089766_, _089767_, _089768_, _089769_, _089770_, _089771_, _089772_, _089773_, _089774_, _089775_, _089776_, _089777_, _089778_, _089779_, _089780_, _089781_, _089782_, _089783_, _089784_, _089785_, _089786_, _089787_, _089788_, _089789_, _089790_, _089791_, _089792_, _089793_, _089794_, _089795_, _089796_, _089797_, _089798_, _089799_, _089800_, _089801_, _089802_, _089803_, _089804_, _089805_, _089806_, _089807_, _089808_, _089809_, _089810_, _089811_, _089812_, _089813_, _089814_, _089815_, _089816_, _089817_, _089818_, _089819_, _089820_, _089821_, _089822_, _089823_, _089824_, _089825_, _089826_, _089827_, _089828_, _089829_, _089830_, _089831_, _089832_, _089833_, _089834_, _089835_, _089836_, _089837_, _089838_, _089839_, _089840_, _089841_, _089842_, _089843_, _089844_, _089845_, _089846_, _089847_, _089848_, _089849_, _089850_, _089851_, _089852_, _089853_, _089854_, _089855_, _089856_, _089857_, _089858_, _089859_, _089860_, _089861_, _089862_, _089863_, _089864_, _089865_, _089866_, _089867_, _089868_, _089869_, _089870_, _089871_, _089872_, _089873_, _089874_, _089875_, _089876_, _089877_, _089878_, _089879_, _089880_, _089881_, _089882_, _089883_, _089884_, _089885_, _089886_, _089887_, _089888_, _089889_, _089890_, _089891_, _089892_, _089893_, _089894_, _089895_, _089896_, _089897_, _089898_, _089899_, _089900_, _089901_, _089902_, _089903_, _089904_, _089905_, _089906_, _089907_, _089908_, _089909_, _089910_, _089911_, _089912_, _089913_, _089914_, _089915_, _089916_, _089917_, _089918_, _089919_, _089920_, _089921_, _089922_, _089923_, _089924_, _089925_, _089926_, _089927_, _089928_, _089929_, _089930_, _089931_, _089932_, _089933_, _089934_, _089935_, _089936_, _089937_, _089938_, _089939_, _089940_, _089941_, _089942_, _089943_, _089944_, _089945_, _089946_, _089947_, _089948_, _089949_, _089950_, _089951_, _089952_, _089953_, _089954_, _089955_, _089956_, _089957_, _089958_, _089959_, _089960_, _089961_, _089962_, _089963_, _089964_, _089965_, _089966_, _089967_, _089968_, _089969_, _089970_, _089971_, _089972_, _089973_, _089974_, _089975_, _089976_, _089977_, _089978_, _089979_, _089980_, _089981_, _089982_, _089983_, _089984_, _089985_, _089986_, _089987_, _089988_, _089989_, _089990_, _089991_, _089992_, _089993_, _089994_, _089995_, _089996_, _089997_, _089998_, _089999_, _090000_, _090001_, _090002_, _090003_, _090004_, _090005_, _090006_, _090007_, _090008_, _090009_, _090010_, _090011_, _090012_, _090013_, _090014_, _090015_, _090016_, _090017_, _090018_, _090019_, _090020_, _090021_, _090022_, _090023_, _090024_, _090025_, _090026_, _090027_, _090028_, _090029_, _090030_, _090031_, _090032_, _090033_, _090034_, _090035_, _090036_, _090037_, _090038_, _090039_, _090040_, _090041_, _090042_, _090043_, _090044_, _090045_, _090046_, _090047_, _090048_, _090049_, _090050_, _090051_, _090052_, _090053_, _090054_, _090055_, _090056_, _090057_, _090058_, _090059_, _090060_, _090061_, _090062_, _090063_, _090064_, _090065_, _090066_, _090067_, _090068_, _090069_, _090070_, _090071_, _090072_, _090073_, _090074_, _090075_, _090076_, _090077_, _090078_, _090079_, _090080_, _090081_, _090082_, _090083_, _090084_, _090085_, _090086_, _090087_, _090088_, _090089_, _090090_, _090091_, _090092_, _090093_, _090094_, _090095_, _090096_, _090097_, _090098_, _090099_, _090100_, _090101_, _090102_, _090103_, _090104_, _090105_, _090106_, _090107_, _090108_, _090109_, _090110_, _090111_, _090112_, _090113_, _090114_, _090115_, _090116_, _090117_, _090118_, _090119_, _090120_, _090121_, _090122_, _090123_, _090124_, _090125_, _090126_, _090127_, _090128_, _090129_, _090130_, _090131_, _090132_, _090133_, _090134_, _090135_, _090136_, _090137_, _090138_, _090139_, _090140_, _090141_, _090142_, _090143_, _090144_, _090145_, _090146_, _090147_, _090148_, _090149_, _090150_, _090151_, _090152_, _090153_, _090154_, _090155_, _090156_, _090157_, _090158_, _090159_, _090160_, _090161_, _090162_, _090163_, _090164_, _090165_, _090166_, _090167_, _090168_, _090169_, _090170_, _090171_, _090172_, _090173_, _090174_, _090175_, _090176_, _090177_, _090178_, _090179_, _090180_, _090181_, _090182_, _090183_, _090184_, _090185_, _090186_, _090187_, _090188_, _090189_, _090190_, _090191_, _090192_, _090193_, _090194_, _090195_, _090196_, _090197_, _090198_, _090199_, _090200_, _090201_, _090202_, _090203_, _090204_, _090205_, _090206_, _090207_, _090208_, _090209_, _090210_, _090211_, _090212_, _090213_, _090214_, _090215_, _090216_, _090217_, _090218_, _090219_, _090220_, _090221_, _090222_, _090223_, _090224_, _090225_, _090226_, _090227_, _090228_, _090229_, _090230_, _090231_, _090232_, _090233_, _090234_, _090235_, _090236_, _090237_, _090238_, _090239_, _090240_, _090241_, _090242_, _090243_, _090244_, _090245_, _090246_, _090247_, _090248_, _090249_, _090250_, _090251_, _090252_, _090253_, _090254_, _090255_, _090256_, _090257_, _090258_, _090259_, _090260_, _090261_, _090262_, _090263_, _090264_, _090265_, _090266_, _090267_, _090268_, _090269_, _090270_, _090271_, _090272_, _090273_, _090274_, _090275_, _090276_, _090277_, _090278_, _090279_, _090280_, _090281_, _090282_, _090283_, _090284_, _090285_, _090286_, _090287_, _090288_, _090289_, _090290_, _090291_, _090292_, _090293_, _090294_, _090295_, _090296_, _090297_, _090298_, _090299_, _090300_, _090301_, _090302_, _090303_, _090304_, _090305_, _090306_, _090307_, _090308_, _090309_, _090310_, _090311_, _090312_, _090313_, _090314_, _090315_, _090316_, _090317_, _090318_, _090319_, _090320_, _090321_, _090322_, _090323_, _090324_, _090325_, _090326_, _090327_, _090328_, _090329_, _090330_, _090331_, _090332_, _090333_, _090334_, _090335_, _090336_, _090337_, _090338_, _090339_, _090340_, _090341_, _090342_, _090343_, _090344_, _090345_, _090346_, _090347_, _090348_, _090349_, _090350_, _090351_, _090352_, _090353_, _090354_, _090355_, _090356_, _090357_, _090358_, _090359_, _090360_, _090361_, _090362_, _090363_, _090364_, _090365_, _090366_, _090367_, _090368_, _090369_, _090370_, _090371_, _090372_, _090373_, _090374_, _090375_, _090376_, _090377_, _090378_, _090379_, _090380_, _090381_, _090382_, _090383_, _090384_, _090385_, _090386_, _090387_, _090388_, _090389_, _090390_, _090391_, _090392_, _090393_, _090394_, _090395_, _090396_, _090397_, _090398_, _090399_, _090400_, _090401_, _090402_, _090403_, _090404_, _090405_, _090406_, _090407_, _090408_, _090409_, _090410_, _090411_, _090412_, _090413_, _090414_, _090415_, _090416_, _090417_, _090418_, _090419_, _090420_, _090421_, _090422_, _090423_, _090424_, _090425_, _090426_, _090427_, _090428_, _090429_, _090430_, _090431_, _090432_, _090433_, _090434_, _090435_, _090436_, _090437_, _090438_, _090439_, _090440_, _090441_, _090442_, _090443_, _090444_, _090445_, _090446_, _090447_, _090448_, _090449_, _090450_, _090451_, _090452_, _090453_, _090454_, _090455_, _090456_, _090457_, _090458_, _090459_, _090460_, _090461_, _090462_, _090463_, _090464_, _090465_, _090466_, _090467_, _090468_, _090469_, _090470_, _090471_, _090472_, _090473_, _090474_, _090475_, _090476_, _090477_, _090478_, _090479_, _090480_, _090481_, _090482_, _090483_, _090484_, _090485_, _090486_, _090487_, _090488_, _090489_, _090490_, _090491_, _090492_, _090493_, _090494_, _090495_, _090496_, _090497_, _090498_, _090499_, _090500_, _090501_, _090502_, _090503_, _090504_, _090505_, _090506_, _090507_, _090508_, _090509_, _090510_, _090511_, _090512_, _090513_, _090514_, _090515_, _090516_, _090517_, _090518_, _090519_, _090520_, _090521_, _090522_, _090523_, _090524_, _090525_, _090526_, _090527_, _090528_, _090529_, _090530_, _090531_, _090532_, _090533_, _090534_, _090535_, _090536_, _090537_, _090538_, _090539_, _090540_, _090541_, _090542_, _090543_, _090544_, _090545_, _090546_, _090547_, _090548_, _090549_, _090550_, _090551_, _090552_, _090553_, _090554_, _090555_, _090556_, _090557_, _090558_, _090559_, _090560_, _090561_, _090562_, _090563_, _090564_, _090565_, _090566_, _090567_, _090568_, _090569_, _090570_, _090571_, _090572_, _090573_, _090574_, _090575_, _090576_, _090577_, _090578_, _090579_, _090580_, _090581_, _090582_, _090583_, _090584_, _090585_, _090586_, _090587_, _090588_, _090589_, _090590_, _090591_, _090592_, _090593_, _090594_, _090595_, _090596_, _090597_, _090598_, _090599_, _090600_, _090601_, _090602_, _090603_, _090604_, _090605_, _090606_, _090607_, _090608_, _090609_, _090610_, _090611_, _090612_, _090613_, _090614_, _090615_, _090616_, _090617_, _090618_, _090619_, _090620_, _090621_, _090622_, _090623_, _090624_, _090625_, _090626_, _090627_, _090628_, _090629_, _090630_, _090631_, _090632_, _090633_, _090634_, _090635_, _090636_, _090637_, _090638_, _090639_, _090640_, _090641_, _090642_, _090643_, _090644_, _090645_, _090646_, _090647_, _090648_, _090649_, _090650_, _090651_, _090652_, _090653_, _090654_, _090655_, _090656_, _090657_, _090658_, _090659_, _090660_, _090661_, _090662_, _090663_, _090664_, _090665_, _090666_, _090667_, _090668_, _090669_, _090670_, _090671_, _090672_, _090673_, _090674_, _090675_, _090676_, _090677_, _090678_, _090679_, _090680_, _090681_, _090682_, _090683_, _090684_, _090685_, _090686_, _090687_, _090688_, _090689_, _090690_, _090691_, _090692_, _090693_, _090694_, _090695_, _090696_, _090697_, _090698_, _090699_, _090700_, _090701_, _090702_, _090703_, _090704_, _090705_, _090706_, _090707_, _090708_, _090709_, _090710_, _090711_, _090712_, _090713_, _090714_, _090715_, _090716_, _090717_, _090718_, _090719_, _090720_, _090721_, _090722_, _090723_, _090724_, _090725_, _090726_, _090727_, _090728_, _090729_, _090730_, _090731_, _090732_, _090733_, _090734_, _090735_, _090736_, _090737_, _090738_, _090739_, _090740_, _090741_, _090742_, _090743_, _090744_, _090745_, _090746_, _090747_, _090748_, _090749_, _090750_, _090751_, _090752_, _090753_, _090754_, _090755_, _090756_, _090757_, _090758_, _090759_, _090760_, _090761_, _090762_, _090763_, _090764_, _090765_, _090766_, _090767_, _090768_, _090769_, _090770_, _090771_, _090772_, _090773_, _090774_, _090775_, _090776_, _090777_, _090778_, _090779_, _090780_, _090781_, _090782_, _090783_, _090784_, _090785_, _090786_, _090787_, _090788_, _090789_, _090790_, _090791_, _090792_, _090793_, _090794_, _090795_, _090796_, _090797_, _090798_, _090799_, _090800_, _090801_, _090802_, _090803_, _090804_, _090805_, _090806_, _090807_, _090808_, _090809_, _090810_, _090811_, _090812_, _090813_, _090814_, _090815_, _090816_, _090817_, _090818_, _090819_, _090820_, _090821_, _090822_, _090823_, _090824_, _090825_, _090826_, _090827_, _090828_, _090829_, _090830_, _090831_, _090832_, _090833_, _090834_, _090835_, _090836_, _090837_, _090838_, _090839_, _090840_, _090841_, _090842_, _090843_, _090844_, _090845_, _090846_, _090847_, _090848_, _090849_, _090850_, _090851_, _090852_, _090853_, _090854_, _090855_, _090856_, _090857_, _090858_, _090859_, _090860_, _090861_, _090862_, _090863_, _090864_, _090865_, _090866_, _090867_, _090868_, _090869_, _090870_, _090871_, _090872_, _090873_, _090874_, _090875_, _090876_, _090877_, _090878_, _090879_, _090880_, _090881_, _090882_, _090883_, _090884_, _090885_, _090886_, _090887_, _090888_, _090889_, _090890_, _090891_, _090892_, _090893_, _090894_, _090895_, _090896_, _090897_, _090898_, _090899_, _090900_, _090901_, _090902_, _090903_, _090904_, _090905_, _090906_, _090907_, _090908_, _090909_, _090910_, _090911_, _090912_, _090913_, _090914_, _090915_, _090916_, _090917_, _090918_, _090919_, _090920_, _090921_, _090922_, _090923_, _090924_, _090925_, _090926_, _090927_, _090928_, _090929_, _090930_, _090931_, _090932_, _090933_, _090934_, _090935_, _090936_, _090937_, _090938_, _090939_, _090940_, _090941_, _090942_, _090943_, _090944_, _090945_, _090946_, _090947_, _090948_, _090949_, _090950_, _090951_, _090952_, _090953_, _090954_, _090955_, _090956_, _090957_, _090958_, _090959_, _090960_, _090961_, _090962_, _090963_, _090964_, _090965_, _090966_, _090967_, _090968_, _090969_, _090970_, _090971_, _090972_, _090973_, _090974_, _090975_, _090976_, _090977_, _090978_, _090979_, _090980_, _090981_, _090982_, _090983_, _090984_, _090985_, _090986_, _090987_, _090988_, _090989_, _090990_, _090991_, _090992_, _090993_, _090994_, _090995_, _090996_, _090997_, _090998_, _090999_, _091000_, _091001_, _091002_, _091003_, _091004_, _091005_, _091006_, _091007_, _091008_, _091009_, _091010_, _091011_, _091012_, _091013_, _091014_, _091015_, _091016_, _091017_, _091018_, _091019_, _091020_, _091021_, _091022_, _091023_, _091024_, _091025_, _091026_, _091027_, _091028_, _091029_, _091030_, _091031_, _091032_, _091033_, _091034_, _091035_, _091036_, _091037_, _091038_, _091039_, _091040_, _091041_, _091042_, _091043_, _091044_, _091045_, _091046_, _091047_, _091048_, _091049_, _091050_, _091051_, _091052_, _091053_, _091054_, _091055_, _091056_, _091057_, _091058_, _091059_, _091060_, _091061_, _091062_, _091063_, _091064_, _091065_, _091066_, _091067_, _091068_, _091069_, _091070_, _091071_, _091072_, _091073_, _091074_, _091075_, _091076_, _091077_, _091078_, _091079_, _091080_, _091081_, _091082_, _091083_, _091084_, _091085_, _091086_, _091087_, _091088_, _091089_, _091090_, _091091_, _091092_, _091093_, _091094_, _091095_, _091096_, _091097_, _091098_, _091099_, _091100_, _091101_, _091102_, _091103_, _091104_, _091105_, _091106_, _091107_, _091108_, _091109_, _091110_, _091111_, _091112_, _091113_, _091114_, _091115_, _091116_, _091117_, _091118_, _091119_, _091120_, _091121_, _091122_, _091123_, _091124_, _091125_, _091126_, _091127_, _091128_, _091129_, _091130_, _091131_, _091132_, _091133_, _091134_, _091135_, _091136_, _091137_, _091138_, _091139_, _091140_, _091141_, _091142_, _091143_, _091144_, _091145_, _091146_, _091147_, _091148_, _091149_, _091150_, _091151_, _091152_, _091153_, _091154_, _091155_, _091156_, _091157_, _091158_, _091159_, _091160_, _091161_, _091162_, _091163_, _091164_, _091165_, _091166_, _091167_, _091168_, _091169_, _091170_, _091171_, _091172_, _091173_, _091174_, _091175_, _091176_, _091177_, _091178_, _091179_, _091180_, _091181_, _091182_, _091183_, _091184_, _091185_, _091186_, _091187_, _091188_, _091189_, _091190_, _091191_, _091192_, _091193_, _091194_, _091195_, _091196_, _091197_, _091198_, _091199_, _091200_, _091201_, _091202_, _091203_, _091204_, _091205_, _091206_, _091207_, _091208_, _091209_, _091210_, _091211_, _091212_, _091213_, _091214_, _091215_, _091216_, _091217_, _091218_, _091219_, _091220_, _091221_, _091222_, _091223_, _091224_, _091225_, _091226_, _091227_, _091228_, _091229_, _091230_, _091231_, _091232_, _091233_, _091234_, _091235_, _091236_, _091237_, _091238_, _091239_, _091240_, _091241_, _091242_, _091243_, _091244_, _091245_, _091246_, _091247_, _091248_, _091249_, _091250_, _091251_, _091252_, _091253_, _091254_, _091255_, _091256_, _091257_, _091258_, _091259_, _091260_, _091261_, _091262_, _091263_, _091264_, _091265_, _091266_, _091267_, _091268_, _091269_, _091270_, _091271_, _091272_, _091273_, _091274_, _091275_, _091276_, _091277_, _091278_, _091279_, _091280_, _091281_, _091282_, _091283_, _091284_, _091285_, _091286_, _091287_, _091288_, _091289_, _091290_, _091291_, _091292_, _091293_, _091294_, _091295_, _091296_, _091297_, _091298_, _091299_, _091300_, _091301_, _091302_, _091303_, _091304_, _091305_, _091306_, _091307_, _091308_, _091309_, _091310_, _091311_, _091312_, _091313_, _091314_, _091315_, _091316_, _091317_, _091318_, _091319_, _091320_, _091321_, _091322_, _091323_, _091324_, _091325_, _091326_, _091327_, _091328_, _091329_, _091330_, _091331_, _091332_, _091333_, _091334_, _091335_, _091336_, _091337_, _091338_, _091339_, _091340_, _091341_, _091342_, _091343_, _091344_, _091345_, _091346_, _091347_, _091348_, _091349_, _091350_, _091351_, _091352_, _091353_, _091354_, _091355_, _091356_, _091357_, _091358_, _091359_, _091360_, _091361_, _091362_, _091363_, _091364_, _091365_, _091366_, _091367_, _091368_, _091369_, _091370_, _091371_, _091372_, _091373_, _091374_, _091375_, _091376_, _091377_, _091378_, _091379_, _091380_, _091381_, _091382_, _091383_, _091384_, _091385_, _091386_, _091387_, _091388_, _091389_, _091390_, _091391_, _091392_, _091393_, _091394_, _091395_, _091396_, _091397_, _091398_, _091399_, _091400_, _091401_, _091402_, _091403_, _091404_, _091405_, _091406_, _091407_, _091408_, _091409_, _091410_, _091411_, _091412_, _091413_, _091414_, _091415_, _091416_, _091417_, _091418_, _091419_, _091420_, _091421_, _091422_, _091423_, _091424_, _091425_, _091426_, _091427_, _091428_, _091429_, _091430_, _091431_, _091432_, _091433_, _091434_, _091435_, _091436_, _091437_, _091438_, _091439_, _091440_, _091441_, _091442_, _091443_, _091444_, _091445_, _091446_, _091447_, _091448_, _091449_, _091450_, _091451_, _091452_, _091453_, _091454_, _091455_, _091456_, _091457_, _091458_, _091459_, _091460_, _091461_, _091462_, _091463_, _091464_, _091465_, _091466_, _091467_, _091468_, _091469_, _091470_, _091471_, _091472_, _091473_, _091474_, _091475_, _091476_, _091477_, _091478_, _091479_, _091480_, _091481_, _091482_, _091483_, _091484_, _091485_, _091486_, _091487_, _091488_, _091489_, _091490_, _091491_, _091492_, _091493_, _091494_, _091495_, _091496_, _091497_, _091498_, _091499_, _091500_, _091501_, _091502_, _091503_, _091504_, _091505_, _091506_, _091507_, _091508_, _091509_, _091510_, _091511_, _091512_, _091513_, _091514_, _091515_, _091516_, _091517_, _091518_, _091519_, _091520_, _091521_, _091522_, _091523_, _091524_, _091525_, _091526_, _091527_, _091528_, _091529_, _091530_, _091531_, _091532_, _091533_, _091534_, _091535_, _091536_, _091537_, _091538_, _091539_, _091540_, _091541_, _091542_, _091543_, _091544_, _091545_, _091546_, _091547_, _091548_, _091549_, _091550_, _091551_, _091552_, _091553_, _091554_, _091555_, _091556_, _091557_, _091558_, _091559_, _091560_, _091561_, _091562_, _091563_, _091564_, _091565_, _091566_, _091567_, _091568_, _091569_, _091570_, _091571_, _091572_, _091573_, _091574_, _091575_, _091576_, _091577_, _091578_, _091579_, _091580_, _091581_, _091582_, _091583_, _091584_, _091585_, _091586_, _091587_, _091588_, _091589_, _091590_, _091591_, _091592_, _091593_, _091594_, _091595_, _091596_, _091597_, _091598_, _091599_, _091600_, _091601_, _091602_, _091603_, _091604_, _091605_, _091606_, _091607_, _091608_, _091609_, _091610_, _091611_, _091612_, _091613_, _091614_, _091615_, _091616_, _091617_, _091618_, _091619_, _091620_, _091621_, _091622_, _091623_, _091624_, _091625_, _091626_, _091627_, _091628_, _091629_, _091630_, _091631_, _091632_, _091633_, _091634_, _091635_, _091636_, _091637_, _091638_, _091639_, _091640_, _091641_, _091642_, _091643_, _091644_, _091645_, _091646_, _091647_, _091648_, _091649_, _091650_, _091651_, _091652_, _091653_, _091654_, _091655_, _091656_, _091657_, _091658_, _091659_, _091660_, _091661_, _091662_, _091663_, _091664_, _091665_, _091666_, _091667_, _091668_, _091669_, _091670_, _091671_, _091672_, _091673_, _091674_, _091675_, _091676_, _091677_, _091678_, _091679_, _091680_, _091681_, _091682_, _091683_, _091684_, _091685_, _091686_, _091687_, _091688_, _091689_, _091690_, _091691_, _091692_, _091693_, _091694_, _091695_, _091696_, _091697_, _091698_, _091699_, _091700_, _091701_, _091702_, _091703_, _091704_, _091705_, _091706_, _091707_, _091708_, _091709_, _091710_, _091711_, _091712_, _091713_, _091714_, _091715_, _091716_, _091717_, _091718_, _091719_, _091720_, _091721_, _091722_, _091723_, _091724_, _091725_, _091726_, _091727_, _091728_, _091729_, _091730_, _091731_, _091732_, _091733_, _091734_, _091735_, _091736_, _091737_, _091738_, _091739_, _091740_, _091741_, _091742_, _091743_, _091744_, _091745_, _091746_, _091747_, _091748_, _091749_, _091750_, _091751_, _091752_, _091753_, _091754_, _091755_, _091756_, _091757_, _091758_, _091759_, _091760_, _091761_, _091762_, _091763_, _091764_, _091765_, _091766_, _091767_, _091768_, _091769_, _091770_, _091771_, _091772_, _091773_, _091774_, _091775_, _091776_, _091777_, _091778_, _091779_, _091780_, _091781_, _091782_, _091783_, _091784_, _091785_, _091786_, _091787_, _091788_, _091789_, _091790_, _091791_, _091792_, _091793_, _091794_, _091795_, _091796_, _091797_, _091798_, _091799_, _091800_, _091801_, _091802_, _091803_, _091804_, _091805_, _091806_, _091807_, _091808_, _091809_, _091810_, _091811_, _091812_, _091813_, _091814_, _091815_, _091816_, _091817_, _091818_, _091819_, _091820_, _091821_, _091822_, _091823_, _091824_, _091825_, _091826_, _091827_, _091828_, _091829_, _091830_, _091831_, _091832_, _091833_, _091834_, _091835_, _091836_, _091837_, _091838_, _091839_, _091840_, _091841_, _091842_, _091843_, _091844_, _091845_, _091846_, _091847_, _091848_, _091849_, _091850_, _091851_, _091852_, _091853_, _091854_, _091855_, _091856_, _091857_, _091858_, _091859_, _091860_, _091861_, _091862_, _091863_, _091864_, _091865_, _091866_, _091867_, _091868_, _091869_, _091870_, _091871_, _091872_, _091873_, _091874_, _091875_, _091876_, _091877_, _091878_, _091879_, _091880_, _091881_, _091882_, _091883_, _091884_, _091885_, _091886_, _091887_, _091888_, _091889_, _091890_, _091891_, _091892_, _091893_, _091894_, _091895_, _091896_, _091897_, _091898_, _091899_, _091900_, _091901_, _091902_, _091903_, _091904_, _091905_, _091906_, _091907_, _091908_, _091909_, _091910_, _091911_, _091912_, _091913_, _091914_, _091915_, _091916_, _091917_, _091918_, _091919_, _091920_, _091921_, _091922_, _091923_, _091924_, _091925_, _091926_, _091927_, _091928_, _091929_, _091930_, _091931_, _091932_, _091933_, _091934_, _091935_, _091936_, _091937_, _091938_, _091939_, _091940_, _091941_, _091942_, _091943_, _091944_, _091945_, _091946_, _091947_, _091948_, _091949_, _091950_, _091951_, _091952_, _091953_, _091954_, _091955_, _091956_, _091957_, _091958_, _091959_, _091960_, _091961_, _091962_, _091963_, _091964_, _091965_, _091966_, _091967_, _091968_, _091969_, _091970_, _091971_, _091972_, _091973_, _091974_, _091975_, _091976_, _091977_, _091978_, _091979_, _091980_, _091981_, _091982_, _091983_, _091984_, _091985_, _091986_, _091987_, _091988_, _091989_, _091990_, _091991_, _091992_, _091993_, _091994_, _091995_, _091996_, _091997_, _091998_, _091999_, _092000_, _092001_, _092002_, _092003_, _092004_, _092005_, _092006_, _092007_, _092008_, _092009_, _092010_, _092011_, _092012_, _092013_, _092014_, _092015_, _092016_, _092017_, _092018_, _092019_, _092020_, _092021_, _092022_, _092023_, _092024_, _092025_, _092026_, _092027_, _092028_, _092029_, _092030_, _092031_, _092032_, _092033_, _092034_, _092035_, _092036_, _092037_, _092038_, _092039_, _092040_, _092041_, _092042_, _092043_, _092044_, _092045_, _092046_, _092047_, _092048_, _092049_, _092050_, _092051_, _092052_, _092053_, _092054_, _092055_, _092056_, _092057_, _092058_, _092059_, _092060_, _092061_, _092062_, _092063_, _092064_, _092065_, _092066_, _092067_, _092068_, _092069_, _092070_, _092071_, _092072_, _092073_, _092074_, _092075_, _092076_, _092077_, _092078_, _092079_, _092080_, _092081_, _092082_, _092083_, _092084_, _092085_, _092086_, _092087_, _092088_, _092089_, _092090_, _092091_, _092092_, _092093_, _092094_, _092095_, _092096_, _092097_, _092098_, _092099_, _092100_, _092101_, _092102_, _092103_, _092104_, _092105_, _092106_, _092107_, _092108_, _092109_, _092110_, _092111_, _092112_, _092113_, _092114_, _092115_, _092116_, _092117_, _092118_, _092119_, _092120_, _092121_, _092122_, _092123_, _092124_, _092125_, _092126_, _092127_, _092128_, _092129_, _092130_, _092131_, _092132_, _092133_, _092134_, _092135_, _092136_, _092137_, _092138_, _092139_, _092140_, _092141_, _092142_, _092143_, _092144_, _092145_, _092146_, _092147_, _092148_, _092149_, _092150_, _092151_, _092152_, _092153_, _092154_, _092155_, _092156_, _092157_, _092158_, _092159_, _092160_, _092161_, _092162_, _092163_, _092164_, _092165_, _092166_, _092167_, _092168_, _092169_, _092170_, _092171_, _092172_, _092173_, _092174_, _092175_, _092176_, _092177_, _092178_, _092179_, _092180_, _092181_, _092182_, _092183_, _092184_, _092185_, _092186_, _092187_, _092188_, _092189_, _092190_, _092191_, _092192_, _092193_, _092194_, _092195_, _092196_, _092197_, _092198_, _092199_, _092200_, _092201_, _092202_, _092203_, _092204_, _092205_, _092206_, _092207_, _092208_, _092209_, _092210_, _092211_, _092212_, _092213_, _092214_, _092215_, _092216_, _092217_, _092218_, _092219_, _092220_, _092221_, _092222_, _092223_, _092224_, _092225_, _092226_, _092227_, _092228_, _092229_, _092230_, _092231_, _092232_, _092233_, _092234_, _092235_, _092236_, _092237_, _092238_, _092239_, _092240_, _092241_, _092242_, _092243_, _092244_, _092245_, _092246_, _092247_, _092248_, _092249_, _092250_, _092251_, _092252_, _092253_, _092254_, _092255_, _092256_, _092257_, _092258_, _092259_, _092260_, _092261_, _092262_, _092263_, _092264_, _092265_, _092266_, _092267_, _092268_, _092269_, _092270_, _092271_, _092272_, _092273_, _092274_, _092275_, _092276_, _092277_, _092278_, _092279_, _092280_, _092281_, _092282_, _092283_, _092284_, _092285_, _092286_, _092287_, _092288_, _092289_, _092290_, _092291_, _092292_, _092293_, _092294_, _092295_, _092296_, _092297_, _092298_, _092299_, _092300_, _092301_, _092302_, _092303_, _092304_, _092305_, _092306_, _092307_, _092308_, _092309_, _092310_, _092311_, _092312_, _092313_, _092314_, _092315_, _092316_, _092317_, _092318_, _092319_, _092320_, _092321_, _092322_, _092323_, _092324_, _092325_, _092326_, _092327_, _092328_, _092329_, _092330_, _092331_, _092332_, _092333_, _092334_, _092335_, _092336_, _092337_, _092338_, _092339_, _092340_, _092341_, _092342_, _092343_, _092344_, _092345_, _092346_, _092347_, _092348_, _092349_, _092350_, _092351_, _092352_, _092353_, _092354_, _092355_, _092356_, _092357_, _092358_, _092359_, _092360_, _092361_, _092362_, _092363_, _092364_, _092365_, _092366_, _092367_, _092368_, _092369_, _092370_, _092371_, _092372_, _092373_, _092374_, _092375_, _092376_, _092377_, _092378_, _092379_, _092380_, _092381_, _092382_, _092383_, _092384_, _092385_, _092386_, _092387_, _092388_, _092389_, _092390_, _092391_, _092392_, _092393_, _092394_, _092395_, _092396_, _092397_, _092398_, _092399_, _092400_, _092401_, _092402_, _092403_, _092404_, _092405_, _092406_, _092407_, _092408_, _092409_, _092410_, _092411_, _092412_, _092413_, _092414_, _092415_, _092416_, _092417_, _092418_, _092419_, _092420_, _092421_, _092422_, _092423_, _092424_, _092425_, _092426_, _092427_, _092428_, _092429_, _092430_, _092431_, _092432_, _092433_, _092434_, _092435_, _092436_, _092437_, _092438_, _092439_, _092440_, _092441_, _092442_, _092443_, _092444_, _092445_, _092446_, _092447_, _092448_, _092449_, _092450_, _092451_, _092452_, _092453_, _092454_, _092455_, _092456_, _092457_, _092458_, _092459_, _092460_, _092461_, _092462_, _092463_, _092464_, _092465_, _092466_, _092467_, _092468_, _092469_, _092470_, _092471_, _092472_, _092473_, _092474_, _092475_, _092476_, _092477_, _092478_, _092479_, _092480_, _092481_, _092482_, _092483_, _092484_, _092485_, _092486_, _092487_, _092488_, _092489_, _092490_, _092491_, _092492_, _092493_, _092494_, _092495_, _092496_, _092497_, _092498_, _092499_, _092500_, _092501_, _092502_, _092503_, _092504_, _092505_, _092506_, _092507_, _092508_, _092509_, _092510_, _092511_, _092512_, _092513_, _092514_, _092515_, _092516_, _092517_, _092518_, _092519_, _092520_, _092521_, _092522_, _092523_, _092524_, _092525_, _092526_, _092527_, _092528_, _092529_, _092530_, _092531_, _092532_, _092533_, _092534_, _092535_, _092536_, _092537_, _092538_, _092539_, _092540_, _092541_, _092542_, _092543_, _092544_, _092545_, _092546_, _092547_, _092548_, _092549_, _092550_, _092551_, _092552_, _092553_, _092554_, _092555_, _092556_, _092557_, _092558_, _092559_, _092560_, _092561_, _092562_, _092563_, _092564_, _092565_, _092566_, _092567_, _092568_, _092569_, _092570_, _092571_, _092572_, _092573_, _092574_, _092575_, _092576_, _092577_, _092578_, _092579_, _092580_, _092581_, _092582_, _092583_, _092584_, _092585_, _092586_, _092587_, _092588_, _092589_, _092590_, _092591_, _092592_, _092593_, _092594_, _092595_, _092596_, _092597_, _092598_, _092599_, _092600_, _092601_, _092602_, _092603_, _092604_, _092605_, _092606_, _092607_, _092608_, _092609_, _092610_, _092611_, _092612_, _092613_, _092614_, _092615_, _092616_, _092617_, _092618_, _092619_, _092620_, _092621_, _092622_, _092623_, _092624_, _092625_, _092626_, _092627_, _092628_, _092629_, _092630_, _092631_, _092632_, _092633_, _092634_, _092635_, _092636_, _092637_, _092638_, _092639_, _092640_, _092641_, _092642_, _092643_, _092644_, _092645_, _092646_, _092647_, _092648_, _092649_, _092650_, _092651_, _092652_, _092653_, _092654_, _092655_, _092656_, _092657_, _092658_, _092659_, _092660_, _092661_, _092662_, _092663_, _092664_, _092665_, _092666_, _092667_, _092668_, _092669_, _092670_, _092671_, _092672_, _092673_, _092674_, _092675_, _092676_, _092677_, _092678_, _092679_, _092680_, _092681_, _092682_, _092683_, _092684_, _092685_, _092686_, _092687_, _092688_, _092689_, _092690_, _092691_, _092692_, _092693_, _092694_, _092695_, _092696_, _092697_, _092698_, _092699_, _092700_, _092701_, _092702_, _092703_, _092704_, _092705_, _092706_, _092707_, _092708_, _092709_, _092710_, _092711_, _092712_, _092713_, _092714_, _092715_, _092716_, _092717_, _092718_, _092719_, _092720_, _092721_, _092722_, _092723_, _092724_, _092725_, _092726_, _092727_, _092728_, _092729_, _092730_, _092731_, _092732_, _092733_, _092734_, _092735_, _092736_, _092737_, _092738_, _092739_, _092740_, _092741_, _092742_, _092743_, _092744_, _092745_, _092746_, _092747_, _092748_, _092749_, _092750_, _092751_, _092752_, _092753_, _092754_, _092755_, _092756_, _092757_, _092758_, _092759_, _092760_, _092761_, _092762_, _092763_, _092764_, _092765_, _092766_, _092767_, _092768_, _092769_, _092770_, _092771_, _092772_, _092773_, _092774_, _092775_, _092776_, _092777_, _092778_, _092779_, _092780_, _092781_, _092782_, _092783_, _092784_, _092785_, _092786_, _092787_, _092788_, _092789_, _092790_, _092791_, _092792_, _092793_, _092794_, _092795_, _092796_, _092797_, _092798_, _092799_, _092800_, _092801_, _092802_, _092803_, _092804_, _092805_, _092806_, _092807_, _092808_, _092809_, _092810_, _092811_, _092812_, _092813_, _092814_, _092815_, _092816_, _092817_, _092818_, _092819_, _092820_, _092821_, _092822_, _092823_, _092824_, _092825_, _092826_, _092827_, _092828_, _092829_, _092830_, _092831_, _092832_, _092833_, _092834_, _092835_, _092836_, _092837_, _092838_, _092839_, _092840_, _092841_, _092842_, _092843_, _092844_, _092845_, _092846_, _092847_, _092848_, _092849_, _092850_, _092851_, _092852_, _092853_, _092854_, _092855_, _092856_, _092857_, _092858_, _092859_, _092860_, _092861_, _092862_, _092863_, _092864_, _092865_, _092866_, _092867_, _092868_, _092869_, _092870_, _092871_, _092872_, _092873_, _092874_, _092875_, _092876_, _092877_, _092878_, _092879_, _092880_, _092881_, _092882_, _092883_, _092884_, _092885_, _092886_, _092887_, _092888_, _092889_, _092890_, _092891_, _092892_, _092893_, _092894_, _092895_, _092896_, _092897_, _092898_, _092899_, _092900_, _092901_, _092902_, _092903_, _092904_, _092905_, _092906_, _092907_, _092908_, _092909_, _092910_, _092911_, _092912_, _092913_, _092914_, _092915_, _092916_, _092917_, _092918_, _092919_, _092920_, _092921_, _092922_, _092923_, _092924_, _092925_, _092926_, _092927_, _092928_, _092929_, _092930_, _092931_, _092932_, _092933_, _092934_, _092935_, _092936_, _092937_, _092938_, _092939_, _092940_, _092941_, _092942_, _092943_, _092944_, _092945_, _092946_, _092947_, _092948_, _092949_, _092950_, _092951_, _092952_, _092953_, _092954_, _092955_, _092956_, _092957_, _092958_, _092959_, _092960_, _092961_, _092962_, _092963_, _092964_, _092965_, _092966_, _092967_, _092968_, _092969_, _092970_, _092971_, _092972_, _092973_, _092974_, _092975_, _092976_, _092977_, _092978_, _092979_, _092980_, _092981_, _092982_, _092983_, _092984_, _092985_, _092986_, _092987_, _092988_, _092989_, _092990_, _092991_, _092992_, _092993_, _092994_, _092995_, _092996_, _092997_, _092998_, _092999_, _093000_, _093001_, _093002_, _093003_, _093004_, _093005_, _093006_, _093007_, _093008_, _093009_, _093010_, _093011_, _093012_, _093013_, _093014_, _093015_, _093016_, _093017_, _093018_, _093019_, _093020_, _093021_, _093022_, _093023_, _093024_, _093025_, _093026_, _093027_, _093028_, _093029_, _093030_, _093031_, _093032_, _093033_, _093034_, _093035_, _093036_, _093037_, _093038_, _093039_, _093040_, _093041_, _093042_, _093043_, _093044_, _093045_, _093046_, _093047_, _093048_, _093049_, _093050_, _093051_, _093052_, _093053_, _093054_, _093055_, _093056_, _093057_, _093058_, _093059_, _093060_, _093061_, _093062_, _093063_, _093064_, _093065_, _093066_, _093067_, _093068_, _093069_, _093070_, _093071_, _093072_, _093073_, _093074_, _093075_, _093076_, _093077_, _093078_, _093079_, _093080_, _093081_, _093082_, _093083_, _093084_, _093085_, _093086_, _093087_, _093088_, _093089_, _093090_, _093091_, _093092_, _093093_, _093094_, _093095_, _093096_, _093097_, _093098_, _093099_, _093100_, _093101_, _093102_, _093103_, _093104_, _093105_, _093106_, _093107_, _093108_, _093109_, _093110_, _093111_, _093112_, _093113_, _093114_, _093115_, _093116_, _093117_, _093118_, _093119_, _093120_, _093121_, _093122_, _093123_, _093124_, _093125_, _093126_, _093127_, _093128_, _093129_, _093130_, _093131_, _093132_, _093133_, _093134_, _093135_, _093136_, _093137_, _093138_, _093139_, _093140_, _093141_, _093142_, _093143_, _093144_, _093145_, _093146_, _093147_, _093148_, _093149_, _093150_, _093151_, _093152_, _093153_, _093154_, _093155_, _093156_, _093157_, _093158_, _093159_, _093160_, _093161_, _093162_, _093163_, _093164_, _093165_, _093166_, _093167_, _093168_, _093169_, _093170_, _093171_, _093172_, _093173_, _093174_, _093175_, _093176_, _093177_, _093178_, _093179_, _093180_, _093181_, _093182_, _093183_, _093184_, _093185_, _093186_, _093187_, _093188_, _093189_, _093190_, _093191_, _093192_, _093193_, _093194_, _093195_, _093196_, _093197_, _093198_, _093199_, _093200_, _093201_, _093202_, _093203_, _093204_, _093205_, _093206_, _093207_, _093208_, _093209_, _093210_, _093211_, _093212_, _093213_, _093214_, _093215_, _093216_, _093217_, _093218_, _093219_, _093220_, _093221_, _093222_, _093223_, _093224_, _093225_, _093226_, _093227_, _093228_, _093229_, _093230_, _093231_, _093232_, _093233_, _093234_, _093235_, _093236_, _093237_, _093238_, _093239_, _093240_, _093241_, _093242_, _093243_, _093244_, _093245_, _093246_, _093247_, _093248_, _093249_, _093250_, _093251_, _093252_, _093253_, _093254_, _093255_, _093256_, _093257_, _093258_, _093259_, _093260_, _093261_, _093262_, _093263_, _093264_, _093265_, _093266_, _093267_, _093268_, _093269_, _093270_, _093271_, _093272_, _093273_, _093274_, _093275_, _093276_, _093277_, _093278_, _093279_, _093280_, _093281_, _093282_, _093283_, _093284_, _093285_, _093286_, _093287_, _093288_, _093289_, _093290_, _093291_, _093292_, _093293_, _093294_, _093295_, _093296_, _093297_, _093298_, _093299_, _093300_, _093301_, _093302_, _093303_, _093304_, _093305_, _093306_, _093307_, _093308_, _093309_, _093310_, _093311_, _093312_, _093313_, _093314_, _093315_, _093316_, _093317_, _093318_, _093319_, _093320_, _093321_, _093322_, _093323_, _093324_, _093325_, _093326_, _093327_, _093328_, _093329_, _093330_, _093331_, _093332_, _093333_, _093334_, _093335_, _093336_, _093337_, _093338_, _093339_, _093340_, _093341_, _093342_, _093343_, _093344_, _093345_, _093346_, _093347_, _093348_, _093349_, _093350_, _093351_, _093352_, _093353_, _093354_, _093355_, _093356_, _093357_, _093358_, _093359_, _093360_, _093361_, _093362_, _093363_, _093364_, _093365_, _093366_, _093367_, _093368_, _093369_, _093370_, _093371_, _093372_, _093373_, _093374_, _093375_, _093376_, _093377_, _093378_, _093379_, _093380_, _093381_, _093382_, _093383_, _093384_, _093385_, _093386_, _093387_, _093388_, _093389_, _093390_, _093391_, _093392_, _093393_, _093394_, _093395_, _093396_, _093397_, _093398_, _093399_, _093400_, _093401_, _093402_, _093403_, _093404_, _093405_, _093406_, _093407_, _093408_, _093409_, _093410_, _093411_, _093412_, _093413_, _093414_, _093415_, _093416_, _093417_, _093418_, _093419_, _093420_, _093421_, _093422_, _093423_, _093424_, _093425_, _093426_, _093427_, _093428_, _093429_, _093430_, _093431_, _093432_, _093433_, _093434_, _093435_, _093436_, _093437_, _093438_, _093439_, _093440_, _093441_, _093442_, _093443_, _093444_, _093445_, _093446_, _093447_, _093448_, _093449_, _093450_, _093451_, _093452_, _093453_, _093454_, _093455_, _093456_, _093457_, _093458_, _093459_, _093460_, _093461_, _093462_, _093463_, _093464_, _093465_, _093466_, _093467_, _093468_, _093469_, _093470_, _093471_, _093472_, _093473_, _093474_, _093475_, _093476_, _093477_, _093478_, _093479_, _093480_, _093481_, _093482_, _093483_, _093484_, _093485_, _093486_, _093487_, _093488_, _093489_, _093490_, _093491_, _093492_, _093493_, _093494_, _093495_, _093496_, _093497_, _093498_, _093499_, _093500_, _093501_, _093502_, _093503_, _093504_, _093505_, _093506_, _093507_, _093508_, _093509_, _093510_, _093511_, _093512_, _093513_, _093514_, _093515_, _093516_, _093517_, _093518_, _093519_, _093520_, _093521_, _093522_, _093523_, _093524_, _093525_, _093526_, _093527_, _093528_, _093529_, _093530_, _093531_, _093532_, _093533_, _093534_, _093535_, _093536_, _093537_, _093538_, _093539_, _093540_, _093541_, _093542_, _093543_, _093544_, _093545_, _093546_, _093547_, _093548_, _093549_, _093550_, _093551_, _093552_, _093553_, _093554_, _093555_, _093556_, _093557_, _093558_, _093559_, _093560_, _093561_, _093562_, _093563_, _093564_, _093565_, _093566_, _093567_, _093568_, _093569_, _093570_, _093571_, _093572_, _093573_, _093574_, _093575_, _093576_, _093577_, _093578_, _093579_, _093580_, _093581_, _093582_, _093583_, _093584_, _093585_, _093586_, _093587_, _093588_, _093589_, _093590_, _093591_, _093592_, _093593_, _093594_, _093595_, _093596_, _093597_, _093598_, _093599_, _093600_, _093601_, _093602_, _093603_, _093604_, _093605_, _093606_, _093607_, _093608_, _093609_, _093610_, _093611_, _093612_, _093613_, _093614_, _093615_, _093616_, _093617_, _093618_, _093619_, _093620_, _093621_, _093622_, _093623_, _093624_, _093625_, _093626_, _093627_, _093628_, _093629_, _093630_, _093631_, _093632_, _093633_, _093634_, _093635_, _093636_, _093637_, _093638_, _093639_, _093640_, _093641_, _093642_, _093643_, _093644_, _093645_, _093646_, _093647_, _093648_, _093649_, _093650_, _093651_, _093652_, _093653_, _093654_, _093655_, _093656_, _093657_, _093658_, _093659_, _093660_, _093661_, _093662_, _093663_, _093664_, _093665_, _093666_, _093667_, _093668_, _093669_, _093670_, _093671_, _093672_, _093673_, _093674_, _093675_, _093676_, _093677_, _093678_, _093679_, _093680_, _093681_, _093682_, _093683_, _093684_, _093685_, _093686_, _093687_, _093688_, _093689_, _093690_, _093691_, _093692_, _093693_, _093694_, _093695_, _093696_, _093697_, _093698_, _093699_, _093700_, _093701_, _093702_, _093703_, _093704_, _093705_, _093706_, _093707_, _093708_, _093709_, _093710_, _093711_, _093712_, _093713_, _093714_, _093715_, _093716_, _093717_, _093718_, _093719_, _093720_, _093721_, _093722_, _093723_, _093724_, _093725_, _093726_, _093727_, _093728_, _093729_, _093730_, _093731_, _093732_, _093733_, _093734_, _093735_, _093736_, _093737_, _093738_, _093739_, _093740_, _093741_, _093742_, _093743_, _093744_, _093745_, _093746_, _093747_, _093748_, _093749_, _093750_, _093751_, _093752_, _093753_, _093754_, _093755_, _093756_, _093757_, _093758_, _093759_, _093760_, _093761_, _093762_, _093763_, _093764_, _093765_, _093766_, _093767_, _093768_, _093769_, _093770_, _093771_, _093772_, _093773_, _093774_, _093775_, _093776_, _093777_, _093778_, _093779_, _093780_, _093781_, _093782_, _093783_, _093784_, _093785_, _093786_, _093787_, _093788_, _093789_, _093790_, _093791_, _093792_, _093793_, _093794_, _093795_, _093796_, _093797_, _093798_, _093799_, _093800_, _093801_, _093802_, _093803_, _093804_, _093805_, _093806_, _093807_, _093808_, _093809_, _093810_, _093811_, _093812_, _093813_, _093814_, _093815_, _093816_, _093817_, _093818_, _093819_, _093820_, _093821_, _093822_, _093823_, _093824_, _093825_, _093826_, _093827_, _093828_, _093829_, _093830_, _093831_, _093832_, _093833_, _093834_, _093835_, _093836_, _093837_, _093838_, _093839_, _093840_, _093841_, _093842_, _093843_, _093844_, _093845_, _093846_, _093847_, _093848_, _093849_, _093850_, _093851_, _093852_, _093853_, _093854_, _093855_, _093856_, _093857_, _093858_, _093859_, _093860_, _093861_, _093862_, _093863_, _093864_, _093865_, _093866_, _093867_, _093868_, _093869_, _093870_, _093871_, _093872_, _093873_, _093874_, _093875_, _093876_, _093877_, _093878_, _093879_, _093880_, _093881_, _093882_, _093883_, _093884_, _093885_, _093886_, _093887_, _093888_, _093889_, _093890_, _093891_, _093892_, _093893_, _093894_, _093895_, _093896_, _093897_, _093898_, _093899_, _093900_, _093901_, _093902_, _093903_, _093904_, _093905_, _093906_, _093907_, _093908_, _093909_, _093910_, _093911_, _093912_, _093913_, _093914_, _093915_, _093916_, _093917_, _093918_, _093919_, _093920_, _093921_, _093922_, _093923_, _093924_, _093925_, _093926_, _093927_, _093928_, _093929_, _093930_, _093931_, _093932_, _093933_, _093934_, _093935_, _093936_, _093937_, _093938_, _093939_, _093940_, _093941_, _093942_, _093943_, _093944_, _093945_, _093946_, _093947_, _093948_, _093949_, _093950_, _093951_, _093952_, _093953_, _093954_, _093955_, _093956_, _093957_, _093958_, _093959_, _093960_, _093961_, _093962_, _093963_, _093964_, _093965_, _093966_, _093967_, _093968_, _093969_, _093970_, _093971_, _093972_, _093973_, _093974_, _093975_, _093976_, _093977_, _093978_, _093979_, _093980_, _093981_, _093982_, _093983_, _093984_, _093985_, _093986_, _093987_, _093988_, _093989_, _093990_, _093991_, _093992_, _093993_, _093994_, _093995_, _093996_, _093997_, _093998_, _093999_, _094000_, _094001_, _094002_, _094003_, _094004_, _094005_, _094006_, _094007_, _094008_, _094009_, _094010_, _094011_, _094012_, _094013_, _094014_, _094015_, _094016_, _094017_, _094018_, _094019_, _094020_, _094021_, _094022_, _094023_, _094024_, _094025_, _094026_, _094027_, _094028_, _094029_, _094030_, _094031_, _094032_, _094033_, _094034_, _094035_, _094036_, _094037_, _094038_, _094039_, _094040_, _094041_, _094042_, _094043_, _094044_, _094045_, _094046_, _094047_, _094048_, _094049_, _094050_, _094051_, _094052_, _094053_, _094054_, _094055_, _094056_, _094057_, _094058_, _094059_, _094060_, _094061_, _094062_, _094063_, _094064_, _094065_, _094066_, _094067_, _094068_, _094069_, _094070_, _094071_, _094072_, _094073_, _094074_, _094075_, _094076_, _094077_, _094078_, _094079_, _094080_, _094081_, _094082_, _094083_, _094084_, _094085_, _094086_, _094087_, _094088_, _094089_, _094090_, _094091_, _094092_, _094093_, _094094_, _094095_, _094096_, _094097_, _094098_, _094099_, _094100_, _094101_, _094102_, _094103_, _094104_, _094105_, _094106_, _094107_, _094108_, _094109_, _094110_, _094111_, _094112_, _094113_, _094114_, _094115_, _094116_, _094117_, _094118_, _094119_, _094120_, _094121_, _094122_, _094123_, _094124_, _094125_, _094126_, _094127_, _094128_, _094129_, _094130_, _094131_, _094132_, _094133_, _094134_, _094135_, _094136_, _094137_, _094138_, _094139_, _094140_, _094141_, _094142_, _094143_, _094144_, _094145_, _094146_, _094147_, _094148_, _094149_, _094150_, _094151_, _094152_, _094153_, _094154_, _094155_, _094156_, _094157_, _094158_, _094159_, _094160_, _094161_, _094162_, _094163_, _094164_, _094165_, _094166_, _094167_, _094168_, _094169_, _094170_, _094171_, _094172_, _094173_, _094174_, _094175_, _094176_, _094177_, _094178_, _094179_, _094180_, _094181_, _094182_, _094183_, _094184_, _094185_, _094186_, _094187_, _094188_, _094189_, _094190_, _094191_, _094192_, _094193_, _094194_, _094195_, _094196_, _094197_, _094198_, _094199_, _094200_, _094201_, _094202_, _094203_, _094204_, _094205_, _094206_, _094207_, _094208_, _094209_, _094210_, _094211_, _094212_, _094213_, _094214_, _094215_, _094216_, _094217_, _094218_, _094219_, _094220_, _094221_, _094222_, _094223_, _094224_, _094225_, _094226_, _094227_, _094228_, _094229_, _094230_, _094231_, _094232_, _094233_, _094234_, _094235_, _094236_, _094237_, _094238_, _094239_, _094240_, _094241_, _094242_, _094243_, _094244_, _094245_, _094246_, _094247_, _094248_, _094249_, _094250_, _094251_, _094252_, _094253_, _094254_, _094255_, _094256_, _094257_, _094258_, _094259_, _094260_, _094261_, _094262_, _094263_, _094264_, _094265_, _094266_, _094267_, _094268_, _094269_, _094270_, _094271_, _094272_, _094273_, _094274_, _094275_, _094276_, _094277_, _094278_, _094279_, _094280_, _094281_, _094282_, _094283_, _094284_, _094285_, _094286_, _094287_, _094288_, _094289_, _094290_, _094291_, _094292_, _094293_, _094294_, _094295_, _094296_, _094297_, _094298_, _094299_, _094300_, _094301_, _094302_, _094303_, _094304_, _094305_, _094306_, _094307_, _094308_, _094309_, _094310_, _094311_, _094312_, _094313_, _094314_, _094315_, _094316_, _094317_, _094318_, _094319_, _094320_, _094321_, _094322_, _094323_, _094324_, _094325_, _094326_, _094327_, _094328_, _094329_, _094330_, _094331_, _094332_, _094333_, _094334_, _094335_, _094336_, _094337_, _094338_, _094339_, _094340_, _094341_, _094342_, _094343_, _094344_, _094345_, _094346_, _094347_, _094348_, _094349_, _094350_, _094351_, _094352_, _094353_, _094354_, _094355_, _094356_, _094357_, _094358_, _094359_, _094360_, _094361_, _094362_, _094363_, _094364_, _094365_, _094366_, _094367_, _094368_, _094369_, _094370_, _094371_, _094372_, _094373_, _094374_, _094375_, _094376_, _094377_, _094378_, _094379_, _094380_, _094381_, _094382_, _094383_, _094384_, _094385_, _094386_, _094387_, _094388_, _094389_, _094390_, _094391_, _094392_, _094393_, _094394_, _094395_, _094396_, _094397_, _094398_, _094399_, _094400_, _094401_, _094402_, _094403_, _094404_, _094405_, _094406_, _094407_, _094408_, _094409_, _094410_, _094411_, _094412_, _094413_, _094414_, _094415_, _094416_, _094417_, _094418_, _094419_, _094420_, _094421_, _094422_, _094423_, _094424_, _094425_, _094426_, _094427_, _094428_, _094429_, _094430_, _094431_, _094432_, _094433_, _094434_, _094435_, _094436_, _094437_, _094438_, _094439_, _094440_, _094441_, _094442_, _094443_, _094444_, _094445_, _094446_, _094447_, _094448_, _094449_, _094450_, _094451_, _094452_, _094453_, _094454_, _094455_, _094456_, _094457_, _094458_, _094459_, _094460_, _094461_, _094462_, _094463_, _094464_, _094465_, _094466_, _094467_, _094468_, _094469_, _094470_, _094471_, _094472_, _094473_, _094474_, _094475_, _094476_, _094477_, _094478_, _094479_, _094480_, _094481_, _094482_, _094483_, _094484_, _094485_, _094486_, _094487_, _094488_, _094489_, _094490_, _094491_, _094492_, _094493_, _094494_, _094495_, _094496_, _094497_, _094498_, _094499_, _094500_, _094501_, _094502_, _094503_, _094504_, _094505_, _094506_, _094507_, _094508_, _094509_, _094510_, _094511_, _094512_, _094513_, _094514_, _094515_, _094516_, _094517_, _094518_, _094519_, _094520_, _094521_, _094522_, _094523_, _094524_, _094525_, _094526_, _094527_, _094528_, _094529_, _094530_, _094531_, _094532_, _094533_, _094534_, _094535_, _094536_, _094537_, _094538_, _094539_, _094540_, _094541_, _094542_, _094543_, _094544_, _094545_, _094546_, _094547_, _094548_, _094549_, _094550_, _094551_, _094552_, _094553_, _094554_, _094555_, _094556_, _094557_, _094558_, _094559_, _094560_, _094561_, _094562_, _094563_, _094564_, _094565_, _094566_, _094567_, _094568_, _094569_, _094570_, _094571_, _094572_, _094573_, _094574_, _094575_, _094576_, _094577_, _094578_, _094579_, _094580_, _094581_, _094582_, _094583_, _094584_, _094585_, _094586_, _094587_, _094588_, _094589_, _094590_, _094591_, _094592_, _094593_, _094594_, _094595_, _094596_, _094597_, _094598_, _094599_, _094600_, _094601_, _094602_, _094603_, _094604_, _094605_, _094606_, _094607_, _094608_, _094609_, _094610_, _094611_, _094612_, _094613_, _094614_, _094615_, _094616_, _094617_, _094618_, _094619_, _094620_, _094621_, _094622_, _094623_, _094624_, _094625_, _094626_, _094627_, _094628_, _094629_, _094630_, _094631_, _094632_, _094633_, _094634_, _094635_, _094636_, _094637_, _094638_, _094639_, _094640_, _094641_, _094642_, _094643_, _094644_, _094645_, _094646_, _094647_, _094648_, _094649_, _094650_, _094651_, _094652_, _094653_, _094654_, _094655_, _094656_, _094657_, _094658_, _094659_, _094660_, _094661_, _094662_, _094663_, _094664_, _094665_, _094666_, _094667_, _094668_, _094669_, _094670_, _094671_, _094672_, _094673_, _094674_, _094675_, _094676_, _094677_, _094678_, _094679_, _094680_, _094681_, _094682_, _094683_, _094684_, _094685_, _094686_, _094687_, _094688_, _094689_, _094690_, _094691_, _094692_, _094693_, _094694_, _094695_, _094696_, _094697_, _094698_, _094699_, _094700_, _094701_, _094702_, _094703_, _094704_, _094705_, _094706_, _094707_, _094708_, _094709_, _094710_, _094711_, _094712_, _094713_, _094714_, _094715_, _094716_, _094717_, _094718_, _094719_, _094720_, _094721_, _094722_, _094723_, _094724_, _094725_, _094726_, _094727_, _094728_, _094729_, _094730_, _094731_, _094732_, _094733_, _094734_, _094735_, _094736_, _094737_, _094738_, _094739_, _094740_, _094741_, _094742_, _094743_, _094744_, _094745_, _094746_, _094747_, _094748_, _094749_, _094750_, _094751_, _094752_, _094753_, _094754_, _094755_, _094756_, _094757_, _094758_, _094759_, _094760_, _094761_, _094762_, _094763_, _094764_, _094765_, _094766_, _094767_, _094768_, _094769_, _094770_, _094771_, _094772_, _094773_, _094774_, _094775_, _094776_, _094777_, _094778_, _094779_, _094780_, _094781_, _094782_, _094783_, _094784_, _094785_, _094786_, _094787_, _094788_, _094789_, _094790_, _094791_, _094792_, _094793_, _094794_, _094795_, _094796_, _094797_, _094798_, _094799_, _094800_, _094801_, _094802_, _094803_, _094804_, _094805_, _094806_, _094807_, _094808_, _094809_, _094810_, _094811_, _094812_, _094813_, _094814_, _094815_, _094816_, _094817_, _094818_, _094819_, _094820_, _094821_, _094822_, _094823_, _094824_, _094825_, _094826_, _094827_, _094828_, _094829_, _094830_, _094831_, _094832_, _094833_, _094834_, _094835_, _094836_, _094837_, _094838_, _094839_, _094840_, _094841_, _094842_, _094843_, _094844_, _094845_, _094846_, _094847_, _094848_, _094849_, _094850_, _094851_, _094852_, _094853_, _094854_, _094855_, _094856_, _094857_, _094858_, _094859_, _094860_, _094861_, _094862_, _094863_, _094864_, _094865_, _094866_, _094867_, _094868_, _094869_, _094870_, _094871_, _094872_, _094873_, _094874_, _094875_, _094876_, _094877_, _094878_, _094879_, _094880_, _094881_, _094882_, _094883_, _094884_, _094885_, _094886_, _094887_, _094888_, _094889_, _094890_, _094891_, _094892_, _094893_, _094894_, _094895_, _094896_, _094897_, _094898_, _094899_, _094900_, _094901_, _094902_, _094903_, _094904_, _094905_, _094906_, _094907_, _094908_, _094909_, _094910_, _094911_, _094912_, _094913_, _094914_, _094915_, _094916_, _094917_, _094918_, _094919_, _094920_, _094921_, _094922_, _094923_, _094924_, _094925_, _094926_, _094927_, _094928_, _094929_, _094930_, _094931_, _094932_, _094933_, _094934_, _094935_, _094936_, _094937_, _094938_, _094939_, _094940_, _094941_, _094942_, _094943_, _094944_, _094945_, _094946_, _094947_, _094948_, _094949_, _094950_, _094951_, _094952_, _094953_, _094954_, _094955_, _094956_, _094957_, _094958_, _094959_, _094960_, _094961_, _094962_, _094963_, _094964_, _094965_, _094966_, _094967_, _094968_, _094969_, _094970_, _094971_, _094972_, _094973_, _094974_, _094975_, _094976_, _094977_, _094978_, _094979_, _094980_, _094981_, _094982_, _094983_, _094984_, _094985_, _094986_, _094987_, _094988_, _094989_, _094990_, _094991_, _094992_, _094993_, _094994_, _094995_, _094996_, _094997_, _094998_, _094999_, _095000_, _095001_, _095002_, _095003_, _095004_, _095005_, _095006_, _095007_, _095008_, _095009_, _095010_, _095011_, _095012_, _095013_, _095014_, _095015_, _095016_, _095017_, _095018_, _095019_, _095020_, _095021_, _095022_, _095023_, _095024_, _095025_, _095026_, _095027_, _095028_, _095029_, _095030_, _095031_, _095032_, _095033_, _095034_, _095035_, _095036_, _095037_, _095038_, _095039_, _095040_, _095041_, _095042_, _095043_, _095044_, _095045_, _095046_, _095047_, _095048_, _095049_, _095050_, _095051_, _095052_, _095053_, _095054_, _095055_, _095056_, _095057_, _095058_, _095059_, _095060_, _095061_, _095062_, _095063_, _095064_, _095065_, _095066_, _095067_, _095068_, _095069_, _095070_, _095071_, _095072_, _095073_, _095074_, _095075_, _095076_, _095077_, _095078_, _095079_, _095080_, _095081_, _095082_, _095083_, _095084_, _095085_, _095086_, _095087_, _095088_, _095089_, _095090_, _095091_, _095092_, _095093_, _095094_, _095095_, _095096_, _095097_, _095098_, _095099_, _095100_, _095101_, _095102_, _095103_, _095104_, _095105_, _095106_, _095107_, _095108_, _095109_, _095110_, _095111_, _095112_, _095113_, _095114_, _095115_, _095116_, _095117_, _095118_, _095119_, _095120_, _095121_, _095122_, _095123_, _095124_, _095125_, _095126_, _095127_, _095128_, _095129_, _095130_, _095131_, _095132_, _095133_, _095134_, _095135_, _095136_, _095137_, _095138_, _095139_, _095140_, _095141_, _095142_, _095143_, _095144_, _095145_, _095146_, _095147_, _095148_, _095149_, _095150_, _095151_, _095152_, _095153_, _095154_, _095155_, _095156_, _095157_, _095158_, _095159_, _095160_, _095161_, _095162_, _095163_, _095164_, _095165_, _095166_, _095167_, _095168_, _095169_, _095170_, _095171_, _095172_, _095173_, _095174_, _095175_, _095176_, _095177_, _095178_, _095179_, _095180_, _095181_, _095182_, _095183_, _095184_, _095185_, _095186_, _095187_, _095188_, _095189_, _095190_, _095191_, _095192_, _095193_, _095194_, _095195_, _095196_, _095197_, _095198_, _095199_, _095200_, _095201_, _095202_, _095203_, _095204_, _095205_, _095206_, _095207_, _095208_, _095209_, _095210_, _095211_, _095212_, _095213_, _095214_, _095215_, _095216_, _095217_, _095218_, _095219_, _095220_, _095221_, _095222_, _095223_, _095224_, _095225_, _095226_, _095227_, _095228_, _095229_, _095230_, _095231_, _095232_, _095233_, _095234_, _095235_, _095236_, _095237_, _095238_, _095239_, _095240_, _095241_, _095242_, _095243_, _095244_, _095245_, _095246_, _095247_, _095248_, _095249_, _095250_, _095251_, _095252_, _095253_, _095254_, _095255_, _095256_, _095257_, _095258_, _095259_, _095260_, _095261_, _095262_, _095263_, _095264_, _095265_, _095266_, _095267_, _095268_, _095269_, _095270_, _095271_, _095272_, _095273_, _095274_, _095275_, _095276_, _095277_, _095278_, _095279_, _095280_, _095281_, _095282_, _095283_, _095284_, _095285_, _095286_, _095287_, _095288_, _095289_, _095290_, _095291_, _095292_, _095293_, _095294_, _095295_, _095296_, _095297_, _095298_, _095299_, _095300_, _095301_, _095302_, _095303_, _095304_, _095305_, _095306_, _095307_, _095308_, _095309_, _095310_, _095311_, _095312_, _095313_, _095314_, _095315_, _095316_, _095317_, _095318_, _095319_, _095320_, _095321_, _095322_, _095323_, _095324_, _095325_, _095326_, _095327_, _095328_, _095329_, _095330_, _095331_, _095332_, _095333_, _095334_, _095335_, _095336_, _095337_, _095338_, _095339_, _095340_, _095341_, _095342_, _095343_, _095344_, _095345_, _095346_, _095347_, _095348_, _095349_, _095350_, _095351_, _095352_, _095353_, _095354_, _095355_, _095356_, _095357_, _095358_, _095359_, _095360_, _095361_, _095362_, _095363_, _095364_, _095365_, _095366_, _095367_, _095368_, _095369_, _095370_, _095371_, _095372_, _095373_, _095374_, _095375_, _095376_, _095377_, _095378_, _095379_, _095380_, _095381_, _095382_, _095383_, _095384_, _095385_, _095386_, _095387_, _095388_, _095389_, _095390_, _095391_, _095392_, _095393_, _095394_, _095395_, _095396_, _095397_, _095398_, _095399_, _095400_, _095401_, _095402_, _095403_, _095404_, _095405_, _095406_, _095407_, _095408_, _095409_, _095410_, _095411_, _095412_, _095413_, _095414_, _095415_, _095416_, _095417_, _095418_, _095419_, _095420_, _095421_, _095422_, _095423_, _095424_, _095425_, _095426_, _095427_, _095428_, _095429_, _095430_, _095431_, _095432_, _095433_, _095434_, _095435_, _095436_, _095437_, _095438_, _095439_, _095440_, _095441_, _095442_, _095443_, _095444_, _095445_, _095446_, _095447_, _095448_, _095449_, _095450_, _095451_, _095452_, _095453_, _095454_, _095455_, _095456_, _095457_, _095458_, _095459_, _095460_, _095461_, _095462_, _095463_, _095464_, _095465_, _095466_, _095467_, _095468_, _095469_, _095470_, _095471_, _095472_, _095473_, _095474_, _095475_, _095476_, _095477_, _095478_, _095479_, _095480_, _095481_, _095482_, _095483_, _095484_, _095485_, _095486_, _095487_, _095488_, _095489_, _095490_, _095491_, _095492_, _095493_, _095494_, _095495_, _095496_, _095497_, _095498_, _095499_, _095500_, _095501_, _095502_, _095503_, _095504_, _095505_, _095506_, _095507_, _095508_, _095509_, _095510_, _095511_, _095512_, _095513_, _095514_, _095515_, _095516_, _095517_, _095518_, _095519_, _095520_, _095521_, _095522_, _095523_, _095524_, _095525_, _095526_, _095527_, _095528_, _095529_, _095530_, _095531_, _095532_, _095533_, _095534_, _095535_, _095536_, _095537_, _095538_, _095539_, _095540_, _095541_, _095542_, _095543_, _095544_, _095545_, _095546_, _095547_, _095548_, _095549_, _095550_, _095551_, _095552_, _095553_, _095554_, _095555_, _095556_, _095557_, _095558_, _095559_, _095560_, _095561_, _095562_, _095563_, _095564_, _095565_, _095566_, _095567_, _095568_, _095569_, _095570_, _095571_, _095572_, _095573_, _095574_, _095575_, _095576_, _095577_, _095578_, _095579_, _095580_, _095581_, _095582_, _095583_, _095584_, _095585_, _095586_, _095587_, _095588_, _095589_, _095590_, _095591_, _095592_, _095593_, _095594_, _095595_, _095596_, _095597_, _095598_, _095599_, _095600_, _095601_, _095602_, _095603_, _095604_, _095605_, _095606_, _095607_, _095608_, _095609_, _095610_, _095611_, _095612_, _095613_, _095614_, _095615_, _095616_, _095617_, _095618_, _095619_, _095620_, _095621_, _095622_, _095623_, _095624_, _095625_, _095626_, _095627_, _095628_, _095629_, _095630_, _095631_, _095632_, _095633_, _095634_, _095635_, _095636_, _095637_, _095638_, _095639_, _095640_, _095641_, _095642_, _095643_, _095644_, _095645_, _095646_, _095647_, _095648_, _095649_, _095650_, _095651_, _095652_, _095653_, _095654_, _095655_, _095656_, _095657_, _095658_, _095659_, _095660_, _095661_, _095662_, _095663_, _095664_, _095665_, _095666_, _095667_, _095668_, _095669_, _095670_, _095671_, _095672_, _095673_, _095674_, _095675_, _095676_, _095677_, _095678_, _095679_, _095680_, _095681_, _095682_, _095683_, _095684_, _095685_, _095686_, _095687_, _095688_, _095689_, _095690_, _095691_, _095692_, _095693_, _095694_, _095695_, _095696_, _095697_, _095698_, _095699_, _095700_, _095701_, _095702_, _095703_, _095704_, _095705_, _095706_, _095707_, _095708_, _095709_, _095710_, _095711_, _095712_, _095713_, _095714_, _095715_, _095716_, _095717_, _095718_, _095719_, _095720_, _095721_, _095722_, _095723_, _095724_, _095725_, _095726_, _095727_, _095728_, _095729_, _095730_, _095731_, _095732_, _095733_, _095734_, _095735_, _095736_, _095737_, _095738_, _095739_, _095740_, _095741_, _095742_, _095743_, _095744_, _095745_, _095746_, _095747_, _095748_, _095749_, _095750_, _095751_, _095752_, _095753_, _095754_, _095755_, _095756_, _095757_, _095758_, _095759_, _095760_, _095761_, _095762_, _095763_, _095764_, _095765_, _095766_, _095767_, _095768_, _095769_, _095770_, _095771_, _095772_, _095773_, _095774_, _095775_, _095776_, _095777_, _095778_, _095779_, _095780_, _095781_, _095782_, _095783_, _095784_, _095785_, _095786_, _095787_, _095788_, _095789_, _095790_, _095791_, _095792_, _095793_, _095794_, _095795_, _095796_, _095797_, _095798_, _095799_, _095800_, _095801_, _095802_, _095803_, _095804_, _095805_, _095806_, _095807_, _095808_, _095809_, _095810_, _095811_, _095812_, _095813_, _095814_, _095815_, _095816_, _095817_, _095818_, _095819_, _095820_, _095821_, _095822_, _095823_, _095824_, _095825_, _095826_, _095827_, _095828_, _095829_, _095830_, _095831_, _095832_, _095833_, _095834_, _095835_, _095836_, _095837_, _095838_, _095839_, _095840_, _095841_, _095842_, _095843_, _095844_, _095845_, _095846_, _095847_, _095848_, _095849_, _095850_, _095851_, _095852_, _095853_, _095854_, _095855_, _095856_, _095857_, _095858_, _095859_, _095860_, _095861_, _095862_, _095863_, _095864_, _095865_, _095866_, _095867_, _095868_, _095869_, _095870_, _095871_, _095872_, _095873_, _095874_, _095875_, _095876_, _095877_, _095878_, _095879_, _095880_, _095881_, _095882_, _095883_, _095884_, _095885_, _095886_, _095887_, _095888_, _095889_, _095890_, _095891_, _095892_, _095893_, _095894_, _095895_, _095896_, _095897_, _095898_, _095899_, _095900_, _095901_, _095902_, _095903_, _095904_, _095905_, _095906_, _095907_, _095908_, _095909_, _095910_, _095911_, _095912_, _095913_, _095914_, _095915_, _095916_, _095917_, _095918_, _095919_, _095920_, _095921_, _095922_, _095923_, _095924_, _095925_, _095926_, _095927_, _095928_, _095929_, _095930_, _095931_, _095932_, _095933_, _095934_, _095935_, _095936_, _095937_, _095938_, _095939_, _095940_, _095941_, _095942_, _095943_, _095944_, _095945_, _095946_, _095947_, _095948_, _095949_, _095950_, _095951_, _095952_, _095953_, _095954_, _095955_, _095956_, _095957_, _095958_, _095959_, _095960_, _095961_, _095962_, _095963_, _095964_, _095965_, _095966_, _095967_, _095968_, _095969_, _095970_, _095971_, _095972_, _095973_, _095974_, _095975_, _095976_, _095977_, _095978_, _095979_, _095980_, _095981_, _095982_, _095983_, _095984_, _095985_, _095986_, _095987_, _095988_, _095989_, _095990_, _095991_, _095992_, _095993_, _095994_, _095995_, _095996_, _095997_, _095998_, _095999_, _096000_, _096001_, _096002_, _096003_, _096004_, _096005_, _096006_, _096007_, _096008_, _096009_, _096010_, _096011_, _096012_, _096013_, _096014_, _096015_, _096016_, _096017_, _096018_, _096019_, _096020_, _096021_, _096022_, _096023_, _096024_, _096025_, _096026_, _096027_, _096028_, _096029_, _096030_, _096031_, _096032_, _096033_, _096034_, _096035_, _096036_, _096037_, _096038_, _096039_, _096040_, _096041_, _096042_, _096043_, _096044_, _096045_, _096046_, _096047_, _096048_, _096049_, _096050_, _096051_, _096052_, _096053_, _096054_, _096055_, _096056_, _096057_, _096058_, _096059_, _096060_, _096061_, _096062_, _096063_, _096064_, _096065_, _096066_, _096067_, _096068_, _096069_, _096070_, _096071_, _096072_, _096073_, _096074_, _096075_, _096076_, _096077_, _096078_, _096079_, _096080_, _096081_, _096082_, _096083_, _096084_, _096085_, _096086_, _096087_, _096088_, _096089_, _096090_, _096091_, _096092_, _096093_, _096094_, _096095_, _096096_, _096097_, _096098_, _096099_, _096100_, _096101_, _096102_, _096103_, _096104_, _096105_, _096106_, _096107_, _096108_, _096109_, _096110_, _096111_, _096112_, _096113_, _096114_, _096115_, _096116_, _096117_, _096118_, _096119_, _096120_, _096121_, _096122_, _096123_, _096124_, _096125_, _096126_, _096127_, _096128_, _096129_, _096130_, _096131_, _096132_, _096133_, _096134_, _096135_, _096136_, _096137_, _096138_, _096139_, _096140_, _096141_, _096142_, _096143_, _096144_, _096145_, _096146_, _096147_, _096148_, _096149_, _096150_, _096151_, _096152_, _096153_, _096154_, _096155_, _096156_, _096157_, _096158_, _096159_, _096160_, _096161_, _096162_, _096163_, _096164_, _096165_, _096166_, _096167_, _096168_, _096169_, _096170_, _096171_, _096172_, _096173_, _096174_, _096175_, _096176_, _096177_, _096178_, _096179_, _096180_, _096181_, _096182_, _096183_, _096184_, _096185_, _096186_, _096187_, _096188_, _096189_, _096190_, _096191_, _096192_, _096193_, _096194_, _096195_, _096196_, _096197_, _096198_, _096199_, _096200_, _096201_, _096202_, _096203_, _096204_, _096205_, _096206_, _096207_, _096208_, _096209_, _096210_, _096211_, _096212_, _096213_, _096214_, _096215_, _096216_, _096217_, _096218_, _096219_, _096220_, _096221_, _096222_, _096223_, _096224_, _096225_, _096226_, _096227_, _096228_, _096229_, _096230_, _096231_, _096232_, _096233_, _096234_, _096235_, _096236_, _096237_, _096238_, _096239_, _096240_, _096241_, _096242_, _096243_, _096244_, _096245_, _096246_, _096247_, _096248_, _096249_, _096250_, _096251_, _096252_, _096253_, _096254_, _096255_, _096256_, _096257_, _096258_, _096259_, _096260_, _096261_, _096262_, _096263_, _096264_, _096265_, _096266_, _096267_, _096268_, _096269_, _096270_, _096271_, _096272_, _096273_, _096274_, _096275_, _096276_, _096277_, _096278_, _096279_, _096280_, _096281_, _096282_, _096283_, _096284_, _096285_, _096286_, _096287_, _096288_, _096289_, _096290_, _096291_, _096292_, _096293_, _096294_, _096295_, _096296_, _096297_, _096298_, _096299_, _096300_, _096301_, _096302_, _096303_, _096304_, _096305_, _096306_, _096307_, _096308_, _096309_, _096310_, _096311_, _096312_, _096313_, _096314_, _096315_, _096316_, _096317_, _096318_, _096319_, _096320_, _096321_, _096322_, _096323_, _096324_, _096325_, _096326_, _096327_, _096328_, _096329_, _096330_, _096331_, _096332_, _096333_, _096334_, _096335_, _096336_, _096337_, _096338_, _096339_, _096340_, _096341_, _096342_, _096343_, _096344_, _096345_, _096346_, _096347_, _096348_, _096349_, _096350_, _096351_, _096352_, _096353_, _096354_, _096355_, _096356_, _096357_, _096358_, _096359_, _096360_, _096361_, _096362_, _096363_, _096364_, _096365_, _096366_, _096367_, _096368_, _096369_, _096370_, _096371_, _096372_, _096373_, _096374_, _096375_, _096376_, _096377_, _096378_, _096379_, _096380_, _096381_, _096382_, _096383_, _096384_, _096385_, _096386_, _096387_, _096388_, _096389_, _096390_, _096391_, _096392_, _096393_, _096394_, _096395_, _096396_, _096397_, _096398_, _096399_, _096400_, _096401_, _096402_, _096403_, _096404_, _096405_, _096406_, _096407_, _096408_, _096409_, _096410_, _096411_, _096412_, _096413_, _096414_, _096415_, _096416_, _096417_, _096418_, _096419_, _096420_, _096421_, _096422_, _096423_, _096424_, _096425_, _096426_, _096427_, _096428_, _096429_, _096430_, _096431_, _096432_, _096433_, _096434_, _096435_, _096436_, _096437_, _096438_, _096439_, _096440_, _096441_, _096442_, _096443_, _096444_, _096445_, _096446_, _096447_, _096448_, _096449_, _096450_, _096451_, _096452_, _096453_, _096454_, _096455_, _096456_, _096457_, _096458_, _096459_, _096460_, _096461_, _096462_, _096463_, _096464_, _096465_, _096466_, _096467_, _096468_, _096469_, _096470_, _096471_, _096472_, _096473_, _096474_, _096475_, _096476_, _096477_, _096478_, _096479_, _096480_, _096481_, _096482_, _096483_, _096484_, _096485_, _096486_, _096487_, _096488_, _096489_, _096490_, _096491_, _096492_, _096493_, _096494_, _096495_, _096496_, _096497_, _096498_, _096499_, _096500_, _096501_, _096502_, _096503_, _096504_, _096505_, _096506_, _096507_, _096508_, _096509_, _096510_, _096511_, _096512_, _096513_, _096514_, _096515_, _096516_, _096517_, _096518_, _096519_, _096520_, _096521_, _096522_, _096523_, _096524_, _096525_, _096526_, _096527_, _096528_, _096529_, _096530_, _096531_, _096532_, _096533_, _096534_, _096535_, _096536_, _096537_, _096538_, _096539_, _096540_, _096541_, _096542_, _096543_, _096544_, _096545_, _096546_, _096547_, _096548_, _096549_, _096550_, _096551_, _096552_, _096553_, _096554_, _096555_, _096556_, _096557_, _096558_, _096559_, _096560_, _096561_, _096562_, _096563_, _096564_, _096565_, _096566_, _096567_, _096568_, _096569_, _096570_, _096571_, _096572_, _096573_, _096574_, _096575_, _096576_, _096577_, _096578_, _096579_, _096580_, _096581_, _096582_, _096583_, _096584_, _096585_, _096586_, _096587_, _096588_, _096589_, _096590_, _096591_, _096592_, _096593_, _096594_, _096595_, _096596_, _096597_, _096598_, _096599_, _096600_, _096601_, _096602_, _096603_, _096604_, _096605_, _096606_, _096607_, _096608_, _096609_, _096610_, _096611_, _096612_, _096613_, _096614_, _096615_, _096616_, _096617_, _096618_, _096619_, _096620_, _096621_, _096622_, _096623_, _096624_, _096625_, _096626_, _096627_, _096628_, _096629_, _096630_, _096631_, _096632_, _096633_, _096634_, _096635_, _096636_, _096637_, _096638_, _096639_, _096640_, _096641_, _096642_, _096643_, _096644_, _096645_, _096646_, _096647_, _096648_, _096649_, _096650_, _096651_, _096652_, _096653_, _096654_, _096655_, _096656_, _096657_, _096658_, _096659_, _096660_, _096661_, _096662_, _096663_, _096664_, _096665_, _096666_, _096667_, _096668_, _096669_, _096670_, _096671_, _096672_, _096673_, _096674_, _096675_, _096676_, _096677_, _096678_, _096679_, _096680_, _096681_, _096682_, _096683_, _096684_, _096685_, _096686_, _096687_, _096688_, _096689_, _096690_, _096691_, _096692_, _096693_, _096694_, _096695_, _096696_, _096697_, _096698_, _096699_, _096700_, _096701_, _096702_, _096703_, _096704_, _096705_, _096706_, _096707_, _096708_, _096709_, _096710_, _096711_, _096712_, _096713_, _096714_, _096715_, _096716_, _096717_, _096718_, _096719_, _096720_, _096721_, _096722_, _096723_, _096724_, _096725_, _096726_, _096727_, _096728_, _096729_, _096730_, _096731_, _096732_, _096733_, _096734_, _096735_, _096736_, _096737_, _096738_, _096739_, _096740_, _096741_, _096742_, _096743_, _096744_, _096745_, _096746_, _096747_, _096748_, _096749_, _096750_, _096751_, _096752_, _096753_, _096754_, _096755_, _096756_, _096757_, _096758_, _096759_, _096760_, _096761_, _096762_, _096763_, _096764_, _096765_, _096766_, _096767_, _096768_, _096769_, _096770_, _096771_, _096772_, _096773_, _096774_, _096775_, _096776_, _096777_, _096778_, _096779_, _096780_, _096781_, _096782_, _096783_, _096784_, _096785_, _096786_, _096787_, _096788_, _096789_, _096790_, _096791_, _096792_, _096793_, _096794_, _096795_, _096796_, _096797_, _096798_, _096799_, _096800_, _096801_, _096802_, _096803_, _096804_, _096805_, _096806_, _096807_, _096808_, _096809_, _096810_, _096811_, _096812_, _096813_, _096814_, _096815_, _096816_, _096817_, _096818_, _096819_, _096820_, _096821_, _096822_, _096823_, _096824_, _096825_, _096826_, _096827_, _096828_, _096829_, _096830_, _096831_, _096832_, _096833_, _096834_, _096835_, _096836_, _096837_, _096838_, _096839_, _096840_, _096841_, _096842_, _096843_, _096844_, _096845_, _096846_, _096847_, _096848_, _096849_, _096850_, _096851_, _096852_, _096853_, _096854_, _096855_, _096856_, _096857_, _096858_, _096859_, _096860_, _096861_, _096862_, _096863_, _096864_, _096865_, _096866_, _096867_, _096868_, _096869_, _096870_, _096871_, _096872_, _096873_, _096874_, _096875_, _096876_, _096877_, _096878_, _096879_, _096880_, _096881_, _096882_, _096883_, _096884_, _096885_, _096886_, _096887_, _096888_, _096889_, _096890_, _096891_, _096892_, _096893_, _096894_, _096895_, _096896_, _096897_, _096898_, _096899_, _096900_, _096901_, _096902_, _096903_, _096904_, _096905_, _096906_, _096907_, _096908_, _096909_, _096910_, _096911_, _096912_, _096913_, _096914_, _096915_, _096916_, _096917_, _096918_, _096919_, _096920_, _096921_, _096922_, _096923_, _096924_, _096925_, _096926_, _096927_, _096928_, _096929_, _096930_, _096931_, _096932_, _096933_, _096934_, _096935_, _096936_, _096937_, _096938_, _096939_, _096940_, _096941_, _096942_, _096943_, _096944_, _096945_, _096946_, _096947_, _096948_, _096949_, _096950_, _096951_, _096952_, _096953_, _096954_, _096955_, _096956_, _096957_, _096958_, _096959_, _096960_, _096961_, _096962_, _096963_, _096964_, _096965_, _096966_, _096967_, _096968_, _096969_, _096970_, _096971_, _096972_, _096973_, _096974_, _096975_, _096976_, _096977_, _096978_, _096979_, _096980_, _096981_, _096982_, _096983_, _096984_, _096985_, _096986_, _096987_, _096988_, _096989_, _096990_, _096991_, _096992_, _096993_, _096994_, _096995_, _096996_, _096997_, _096998_, _096999_, _097000_, _097001_, _097002_, _097003_, _097004_, _097005_, _097006_, _097007_, _097008_, _097009_, _097010_, _097011_, _097012_, _097013_, _097014_, _097015_, _097016_, _097017_, _097018_, _097019_, _097020_, _097021_, _097022_, _097023_, _097024_, _097025_, _097026_, _097027_, _097028_, _097029_, _097030_, _097031_, _097032_, _097033_, _097034_, _097035_, _097036_, _097037_, _097038_, _097039_, _097040_, _097041_, _097042_, _097043_, _097044_, _097045_, _097046_, _097047_, _097048_, _097049_, _097050_, _097051_, _097052_, _097053_, _097054_, _097055_, _097056_, _097057_, _097058_, _097059_, _097060_, _097061_, _097062_, _097063_, _097064_, _097065_, _097066_, _097067_, _097068_, _097069_, _097070_, _097071_, _097072_, _097073_, _097074_, _097075_, _097076_, _097077_, _097078_, _097079_, _097080_, _097081_, _097082_, _097083_, _097084_, _097085_, _097086_, _097087_, _097088_, _097089_, _097090_, _097091_, _097092_, _097093_, _097094_, _097095_, _097096_, _097097_, _097098_, _097099_, _097100_, _097101_, _097102_, _097103_, _097104_, _097105_, _097106_, _097107_, _097108_, _097109_, _097110_, _097111_, _097112_, _097113_, _097114_, _097115_, _097116_, _097117_, _097118_, _097119_, _097120_, _097121_, _097122_, _097123_, _097124_, _097125_, _097126_, _097127_, _097128_, _097129_, _097130_, _097131_, _097132_, _097133_, _097134_, _097135_, _097136_, _097137_, _097138_, _097139_, _097140_, _097141_, _097142_, _097143_, _097144_, _097145_, _097146_, _097147_, _097148_, _097149_, _097150_, _097151_, _097152_, _097153_, _097154_, _097155_, _097156_, _097157_, _097158_, _097159_, _097160_, _097161_, _097162_, _097163_, _097164_, _097165_, _097166_, _097167_, _097168_, _097169_, _097170_, _097171_, _097172_, _097173_, _097174_, _097175_, _097176_, _097177_, _097178_, _097179_, _097180_, _097181_, _097182_, _097183_, _097184_, _097185_, _097186_, _097187_, _097188_, _097189_, _097190_, _097191_, _097192_, _097193_, _097194_, _097195_, _097196_, _097197_, _097198_, _097199_, _097200_, _097201_, _097202_, _097203_, _097204_, _097205_, _097206_, _097207_, _097208_, _097209_, _097210_, _097211_, _097212_, _097213_, _097214_, _097215_, _097216_, _097217_, _097218_, _097219_, _097220_, _097221_, _097222_, _097223_, _097224_, _097225_, _097226_, _097227_, _097228_, _097229_, _097230_, _097231_, _097232_, _097233_, _097234_, _097235_, _097236_, _097237_, _097238_, _097239_, _097240_, _097241_, _097242_, _097243_, _097244_, _097245_, _097246_, _097247_, _097248_, _097249_, _097250_, _097251_, _097252_, _097253_, _097254_, _097255_, _097256_, _097257_, _097258_, _097259_, _097260_, _097261_, _097262_, _097263_, _097264_, _097265_, _097266_, _097267_, _097268_, _097269_, _097270_, _097271_, _097272_, _097273_, _097274_, _097275_, _097276_, _097277_, _097278_, _097279_, _097280_, _097281_, _097282_, _097283_, _097284_, _097285_, _097286_, _097287_, _097288_, _097289_, _097290_, _097291_, _097292_, _097293_, _097294_, _097295_, _097296_, _097297_, _097298_, _097299_, _097300_, _097301_, _097302_, _097303_, _097304_, _097305_, _097306_, _097307_, _097308_, _097309_, _097310_, _097311_, _097312_, _097313_, _097314_, _097315_, _097316_, _097317_, _097318_, _097319_, _097320_, _097321_, _097322_, _097323_, _097324_, _097325_, _097326_, _097327_, _097328_, _097329_, _097330_, _097331_, _097332_, _097333_, _097334_, _097335_, _097336_, _097337_, _097338_, _097339_, _097340_, _097341_, _097342_, _097343_, _097344_, _097345_, _097346_, _097347_, _097348_, _097349_, _097350_, _097351_, _097352_, _097353_, _097354_, _097355_, _097356_, _097357_, _097358_, _097359_, _097360_, _097361_, _097362_, _097363_, _097364_, _097365_, _097366_, _097367_, _097368_, _097369_, _097370_, _097371_, _097372_, _097373_, _097374_, _097375_, _097376_, _097377_, _097378_, _097379_, _097380_, _097381_, _097382_, _097383_, _097384_, _097385_, _097386_, _097387_, _097388_, _097389_, _097390_, _097391_, _097392_, _097393_, _097394_, _097395_, _097396_, _097397_, _097398_, _097399_, _097400_, _097401_, _097402_, _097403_, _097404_, _097405_, _097406_, _097407_, _097408_, _097409_, _097410_, _097411_, _097412_, _097413_, _097414_, _097415_, _097416_, _097417_, _097418_, _097419_, _097420_, _097421_, _097422_, _097423_, _097424_, _097425_, _097426_, _097427_, _097428_, _097429_, _097430_, _097431_, _097432_, _097433_, _097434_, _097435_, _097436_, _097437_, _097438_, _097439_, _097440_, _097441_, _097442_, _097443_, _097444_, _097445_, _097446_, _097447_, _097448_, _097449_, _097450_, _097451_, _097452_, _097453_, _097454_, _097455_, _097456_, _097457_, _097458_, _097459_, _097460_, _097461_, _097462_, _097463_, _097464_, _097465_, _097466_, _097467_, _097468_, _097469_, _097470_, _097471_, _097472_, _097473_, _097474_, _097475_, _097476_, _097477_, _097478_, _097479_, _097480_, _097481_, _097482_, _097483_, _097484_, _097485_, _097486_, _097487_, _097488_, _097489_, _097490_, _097491_, _097492_, _097493_, _097494_, _097495_, _097496_, _097497_, _097498_, _097499_, _097500_, _097501_, _097502_, _097503_, _097504_, _097505_, _097506_, _097507_, _097508_, _097509_, _097510_, _097511_, _097512_, _097513_, _097514_, _097515_, _097516_, _097517_, _097518_, _097519_, _097520_, _097521_, _097522_, _097523_, _097524_, _097525_, _097526_, _097527_, _097528_, _097529_, _097530_, _097531_, _097532_, _097533_, _097534_, _097535_, _097536_, _097537_, _097538_, _097539_, _097540_, _097541_, _097542_, _097543_, _097544_, _097545_, _097546_, _097547_, _097548_, _097549_, _097550_, _097551_, _097552_, _097553_, _097554_, _097555_, _097556_, _097557_, _097558_, _097559_, _097560_, _097561_, _097562_, _097563_, _097564_, _097565_, _097566_, _097567_, _097568_, _097569_, _097570_, _097571_, _097572_, _097573_, _097574_, _097575_, _097576_, _097577_, _097578_, _097579_, _097580_, _097581_, _097582_, _097583_, _097584_, _097585_, _097586_, _097587_, _097588_, _097589_, _097590_, _097591_, _097592_, _097593_, _097594_, _097595_, _097596_, _097597_, _097598_, _097599_, _097600_, _097601_, _097602_, _097603_, _097604_, _097605_, _097606_, _097607_, _097608_, _097609_, _097610_, _097611_, _097612_, _097613_, _097614_, _097615_, _097616_, _097617_, _097618_, _097619_, _097620_, _097621_, _097622_, _097623_, _097624_, _097625_, _097626_, _097627_, _097628_, _097629_, _097630_, _097631_, _097632_, _097633_, _097634_, _097635_, _097636_, _097637_, _097638_, _097639_, _097640_, _097641_, _097642_, _097643_, _097644_, _097645_, _097646_, _097647_, _097648_, _097649_, _097650_, _097651_, _097652_, _097653_, _097654_, _097655_, _097656_, _097657_, _097658_, _097659_, _097660_, _097661_, _097662_, _097663_, _097664_, _097665_, _097666_, _097667_, _097668_, _097669_, _097670_, _097671_, _097672_, _097673_, _097674_, _097675_, _097676_, _097677_, _097678_, _097679_, _097680_, _097681_, _097682_, _097683_, _097684_, _097685_, _097686_, _097687_, _097688_, _097689_, _097690_, _097691_, _097692_, _097693_, _097694_, _097695_, _097696_, _097697_, _097698_, _097699_, _097700_, _097701_, _097702_, _097703_, _097704_, _097705_, _097706_, _097707_, _097708_, _097709_, _097710_, _097711_, _097712_, _097713_, _097714_, _097715_, _097716_, _097717_, _097718_, _097719_, _097720_, _097721_, _097722_, _097723_, _097724_, _097725_, _097726_, _097727_, _097728_, _097729_, _097730_, _097731_, _097732_, _097733_, _097734_, _097735_, _097736_, _097737_, _097738_, _097739_, _097740_, _097741_, _097742_, _097743_, _097744_, _097745_, _097746_, _097747_, _097748_, _097749_, _097750_, _097751_, _097752_, _097753_, _097754_, _097755_, _097756_, _097757_, _097758_, _097759_, _097760_, _097761_, _097762_, _097763_, _097764_, _097765_, _097766_, _097767_, _097768_, _097769_, _097770_, _097771_, _097772_, _097773_, _097774_, _097775_, _097776_, _097777_, _097778_, _097779_, _097780_, _097781_, _097782_, _097783_, _097784_, _097785_, _097786_, _097787_, _097788_, _097789_, _097790_, _097791_, _097792_, _097793_, _097794_, _097795_, _097796_, _097797_, _097798_, _097799_, _097800_, _097801_, _097802_, _097803_, _097804_, _097805_, _097806_, _097807_, _097808_, _097809_, _097810_, _097811_, _097812_, _097813_, _097814_, _097815_, _097816_, _097817_, _097818_, _097819_, _097820_, _097821_, _097822_, _097823_, _097824_, _097825_, _097826_, _097827_, _097828_, _097829_, _097830_, _097831_, _097832_, _097833_, _097834_, _097835_, _097836_, _097837_, _097838_, _097839_, _097840_, _097841_, _097842_, _097843_, _097844_, _097845_, _097846_, _097847_, _097848_, _097849_, _097850_, _097851_, _097852_, _097853_, _097854_, _097855_, _097856_, _097857_, _097858_, _097859_, _097860_, _097861_, _097862_, _097863_, _097864_, _097865_, _097866_, _097867_, _097868_, _097869_, _097870_, _097871_, _097872_, _097873_, _097874_, _097875_, _097876_, _097877_, _097878_, _097879_, _097880_, _097881_, _097882_, _097883_, _097884_, _097885_, _097886_, _097887_, _097888_, _097889_, _097890_, _097891_, _097892_, _097893_, _097894_, _097895_, _097896_, _097897_, _097898_, _097899_, _097900_, _097901_, _097902_, _097903_, _097904_, _097905_, _097906_, _097907_, _097908_, _097909_, _097910_, _097911_, _097912_, _097913_, _097914_, _097915_, _097916_, _097917_, _097918_, _097919_, _097920_, _097921_, _097922_, _097923_, _097924_, _097925_, _097926_, _097927_, _097928_, _097929_, _097930_, _097931_, _097932_, _097933_, _097934_, _097935_, _097936_, _097937_, _097938_, _097939_, _097940_, _097941_, _097942_, _097943_, _097944_, _097945_, _097946_, _097947_, _097948_, _097949_, _097950_, _097951_, _097952_, _097953_, _097954_, _097955_, _097956_, _097957_, _097958_, _097959_, _097960_, _097961_, _097962_, _097963_, _097964_, _097965_, _097966_, _097967_, _097968_, _097969_, _097970_, _097971_, _097972_, _097973_, _097974_, _097975_, _097976_, _097977_, _097978_, _097979_, _097980_, _097981_, _097982_, _097983_, _097984_, _097985_, _097986_, _097987_, _097988_, _097989_, _097990_, _097991_, _097992_, _097993_, _097994_, _097995_, _097996_, _097997_, _097998_, _097999_, _098000_, _098001_, _098002_, _098003_, _098004_, _098005_, _098006_, _098007_, _098008_, _098009_, _098010_, _098011_, _098012_, _098013_, _098014_, _098015_, _098016_, _098017_, _098018_, _098019_, _098020_, _098021_, _098022_, _098023_, _098024_, _098025_, _098026_, _098027_, _098028_, _098029_, _098030_, _098031_, _098032_, _098033_, _098034_, _098035_, _098036_, _098037_, _098038_, _098039_, _098040_, _098041_, _098042_, _098043_, _098044_, _098045_, _098046_, _098047_, _098048_, _098049_, _098050_, _098051_, _098052_, _098053_, _098054_, _098055_, _098056_, _098057_, _098058_, _098059_, _098060_, _098061_, _098062_, _098063_, _098064_, _098065_, _098066_, _098067_, _098068_, _098069_, _098070_, _098071_, _098072_, _098073_, _098074_, _098075_, _098076_, _098077_, _098078_, _098079_, _098080_, _098081_, _098082_, _098083_, _098084_, _098085_, _098086_, _098087_, _098088_, _098089_, _098090_, _098091_, _098092_, _098093_, _098094_, _098095_, _098096_, _098097_, _098098_, _098099_, _098100_, _098101_, _098102_, _098103_, _098104_, _098105_, _098106_, _098107_, _098108_, _098109_, _098110_, _098111_, _098112_, _098113_, _098114_, _098115_, _098116_, _098117_, _098118_, _098119_, _098120_, _098121_, _098122_, _098123_, _098124_, _098125_, _098126_, _098127_, _098128_, _098129_, _098130_, _098131_, _098132_, _098133_, _098134_, _098135_, _098136_, _098137_, _098138_, _098139_, _098140_, _098141_, _098142_, _098143_, _098144_, _098145_, _098146_, _098147_, _098148_, _098149_, _098150_, _098151_, _098152_, _098153_, _098154_, _098155_, _098156_, _098157_, _098158_, _098159_, _098160_, _098161_, _098162_, _098163_, _098164_, _098165_, _098166_, _098167_, _098168_, _098169_, _098170_, _098171_, _098172_, _098173_, _098174_, _098175_, _098176_, _098177_, _098178_, _098179_, _098180_, _098181_, _098182_, _098183_, _098184_, _098185_, _098186_, _098187_, _098188_, _098189_, _098190_, _098191_, _098192_, _098193_, _098194_, _098195_, _098196_, _098197_, _098198_, _098199_, _098200_, _098201_, _098202_, _098203_, _098204_, _098205_, _098206_, _098207_, _098208_, _098209_, _098210_, _098211_, _098212_, _098213_, _098214_, _098215_, _098216_, _098217_, _098218_, _098219_, _098220_, _098221_, _098222_, _098223_, _098224_, _098225_, _098226_, _098227_, _098228_, _098229_, _098230_, _098231_, _098232_, _098233_, _098234_, _098235_, _098236_, _098237_, _098238_, _098239_, _098240_, _098241_, _098242_, _098243_, _098244_, _098245_, _098246_, _098247_, _098248_, _098249_, _098250_, _098251_, _098252_, _098253_, _098254_, _098255_, _098256_, _098257_, _098258_, _098259_, _098260_, _098261_, _098262_, _098263_, _098264_, _098265_, _098266_, _098267_, _098268_, _098269_, _098270_, _098271_, _098272_, _098273_, _098274_, _098275_, _098276_, _098277_, _098278_, _098279_, _098280_, _098281_, _098282_, _098283_, _098284_, _098285_, _098286_, _098287_, _098288_, _098289_, _098290_, _098291_, _098292_, _098293_, _098294_, _098295_, _098296_, _098297_, _098298_, _098299_, _098300_, _098301_, _098302_, _098303_, _098304_, _098305_, _098306_, _098307_, _098308_, _098309_, _098310_, _098311_, _098312_, _098313_, _098314_, _098315_, _098316_, _098317_, _098318_, _098319_, _098320_, _098321_, _098322_, _098323_, _098324_, _098325_, _098326_, _098327_, _098328_, _098329_, _098330_, _098331_, _098332_, _098333_, _098334_, _098335_, _098336_, _098337_, _098338_, _098339_, _098340_, _098341_, _098342_, _098343_, _098344_, _098345_, _098346_, _098347_, _098348_, _098349_, _098350_, _098351_, _098352_, _098353_, _098354_, _098355_, _098356_, _098357_, _098358_, _098359_, _098360_, _098361_, _098362_, _098363_, _098364_, _098365_, _098366_, _098367_, _098368_, _098369_, _098370_, _098371_, _098372_, _098373_, _098374_, _098375_, _098376_, _098377_, _098378_, _098379_, _098380_, _098381_, _098382_, _098383_, _098384_, _098385_, _098386_, _098387_, _098388_, _098389_, _098390_, _098391_, _098392_, _098393_, _098394_, _098395_, _098396_, _098397_, _098398_, _098399_, _098400_, _098401_, _098402_, _098403_, _098404_, _098405_, _098406_, _098407_, _098408_, _098409_, _098410_, _098411_, _098412_, _098413_, _098414_, _098415_, _098416_, _098417_, _098418_, _098419_, _098420_, _098421_, _098422_, _098423_, _098424_, _098425_, _098426_, _098427_, _098428_, _098429_, _098430_, _098431_, _098432_, _098433_, _098434_, _098435_, _098436_, _098437_, _098438_, _098439_, _098440_, _098441_, _098442_, _098443_, _098444_, _098445_, _098446_, _098447_, _098448_, _098449_, _098450_, _098451_, _098452_, _098453_, _098454_, _098455_, _098456_, _098457_, _098458_, _098459_, _098460_, _098461_, _098462_, _098463_, _098464_, _098465_, _098466_, _098467_, _098468_, _098469_, _098470_, _098471_, _098472_, _098473_, _098474_, _098475_, _098476_, _098477_, _098478_, _098479_, _098480_, _098481_, _098482_, _098483_, _098484_, _098485_, _098486_, _098487_, _098488_, _098489_, _098490_, _098491_, _098492_, _098493_, _098494_, _098495_, _098496_, _098497_, _098498_, _098499_, _098500_, _098501_, _098502_, _098503_, _098504_, _098505_, _098506_, _098507_, _098508_, _098509_, _098510_, _098511_, _098512_, _098513_, _098514_, _098515_, _098516_, _098517_, _098518_, _098519_, _098520_, _098521_, _098522_, _098523_, _098524_, _098525_, _098526_, _098527_, _098528_, _098529_, _098530_, _098531_, _098532_, _098533_, _098534_, _098535_, _098536_, _098537_, _098538_, _098539_, _098540_, _098541_, _098542_, _098543_, _098544_, _098545_, _098546_, _098547_, _098548_, _098549_, _098550_, _098551_, _098552_, _098553_, _098554_, _098555_, _098556_, _098557_, _098558_, _098559_, _098560_, _098561_, _098562_, _098563_, _098564_, _098565_, _098566_, _098567_, _098568_, _098569_, _098570_, _098571_, _098572_, _098573_, _098574_, _098575_, _098576_, _098577_, _098578_, _098579_, _098580_, _098581_, _098582_, _098583_, _098584_, _098585_, _098586_, _098587_, _098588_, _098589_, _098590_, _098591_, _098592_, _098593_, _098594_, _098595_, _098596_, _098597_, _098598_, _098599_, _098600_, _098601_, _098602_, _098603_, _098604_, _098605_, _098606_, _098607_, _098608_, _098609_, _098610_, _098611_, _098612_, _098613_, _098614_, _098615_, _098616_, _098617_, _098618_, _098619_, _098620_, _098621_, _098622_, _098623_, _098624_, _098625_, _098626_, _098627_, _098628_, _098629_, _098630_, _098631_, _098632_, _098633_, _098634_, _098635_, _098636_, _098637_, _098638_, _098639_, _098640_, _098641_, _098642_, _098643_, _098644_, _098645_, _098646_, _098647_, _098648_, _098649_, _098650_, _098651_, _098652_, _098653_, _098654_, _098655_, _098656_, _098657_, _098658_, _098659_, _098660_, _098661_, _098662_, _098663_, _098664_, _098665_, _098666_, _098667_, _098668_, _098669_, _098670_, _098671_, _098672_, _098673_, _098674_, _098675_, _098676_, _098677_, _098678_, _098679_, _098680_, _098681_, _098682_, _098683_, _098684_, _098685_, _098686_, _098687_, _098688_, _098689_, _098690_, _098691_, _098692_, _098693_, _098694_, _098695_, _098696_, _098697_, _098698_, _098699_, _098700_, _098701_, _098702_, _098703_, _098704_, _098705_, _098706_, _098707_, _098708_, _098709_, _098710_, _098711_, _098712_, _098713_, _098714_, _098715_, _098716_, _098717_, _098718_, _098719_, _098720_, _098721_, _098722_, _098723_, _098724_, _098725_, _098726_, _098727_, _098728_, _098729_, _098730_, _098731_, _098732_, _098733_, _098734_, _098735_, _098736_, _098737_, _098738_, _098739_, _098740_, _098741_, _098742_, _098743_, _098744_, _098745_, _098746_, _098747_, _098748_, _098749_, _098750_, _098751_, _098752_, _098753_, _098754_, _098755_, _098756_, _098757_, _098758_, _098759_, _098760_, _098761_, _098762_, _098763_, _098764_, _098765_, _098766_, _098767_, _098768_, _098769_, _098770_, _098771_, _098772_, _098773_, _098774_, _098775_, _098776_, _098777_, _098778_, _098779_, _098780_, _098781_, _098782_, _098783_, _098784_, _098785_, _098786_, _098787_, _098788_, _098789_, _098790_, _098791_, _098792_, _098793_, _098794_, _098795_, _098796_, _098797_, _098798_, _098799_, _098800_, _098801_, _098802_, _098803_, _098804_, _098805_, _098806_, _098807_, _098808_, _098809_, _098810_, _098811_, _098812_, _098813_, _098814_, _098815_, _098816_, _098817_, _098818_, _098819_, _098820_, _098821_, _098822_, _098823_, _098824_, _098825_, _098826_, _098827_, _098828_, _098829_, _098830_, _098831_, _098832_, _098833_, _098834_, _098835_, _098836_, _098837_, _098838_, _098839_, _098840_, _098841_, _098842_, _098843_, _098844_, _098845_, _098846_, _098847_, _098848_, _098849_, _098850_, _098851_, _098852_, _098853_, _098854_, _098855_, _098856_, _098857_, _098858_, _098859_, _098860_, _098861_, _098862_, _098863_, _098864_, _098865_, _098866_, _098867_, _098868_, _098869_, _098870_, _098871_, _098872_, _098873_, _098874_, _098875_, _098876_, _098877_, _098878_, _098879_, _098880_, _098881_, _098882_, _098883_, _098884_, _098885_, _098886_, _098887_, _098888_, _098889_, _098890_, _098891_, _098892_, _098893_, _098894_, _098895_, _098896_, _098897_, _098898_, _098899_, _098900_, _098901_, _098902_, _098903_, _098904_, _098905_, _098906_, _098907_, _098908_, _098909_, _098910_, _098911_, _098912_, _098913_, _098914_, _098915_, _098916_, _098917_, _098918_, _098919_, _098920_, _098921_, _098922_, _098923_, _098924_, _098925_, _098926_, _098927_, _098928_, _098929_, _098930_, _098931_, _098932_, _098933_, _098934_, _098935_, _098936_, _098937_, _098938_, _098939_, _098940_, _098941_, _098942_, _098943_, _098944_, _098945_, _098946_, _098947_, _098948_, _098949_, _098950_, _098951_, _098952_, _098953_, _098954_, _098955_, _098956_, _098957_, _098958_, _098959_, _098960_, _098961_, _098962_, _098963_, _098964_, _098965_, _098966_, _098967_, _098968_, _098969_, _098970_, _098971_, _098972_, _098973_, _098974_, _098975_, _098976_, _098977_, _098978_, _098979_, _098980_, _098981_, _098982_, _098983_, _098984_, _098985_, _098986_, _098987_, _098988_, _098989_, _098990_, _098991_, _098992_, _098993_, _098994_, _098995_, _098996_, _098997_, _098998_, _098999_, _099000_, _099001_, _099002_, _099003_, _099004_, _099005_, _099006_, _099007_, _099008_, _099009_, _099010_, _099011_, _099012_, _099013_, _099014_, _099015_, _099016_, _099017_, _099018_, _099019_, _099020_, _099021_, _099022_, _099023_, _099024_, _099025_, _099026_, _099027_, _099028_, _099029_, _099030_, _099031_, _099032_, _099033_, _099034_, _099035_, _099036_, _099037_, _099038_, _099039_, _099040_, _099041_, _099042_, _099043_, _099044_, _099045_, _099046_, _099047_, _099048_, _099049_, _099050_, _099051_, _099052_, _099053_, _099054_, _099055_, _099056_, _099057_, _099058_, _099059_, _099060_, _099061_, _099062_, _099063_, _099064_, _099065_, _099066_, _099067_, _099068_, _099069_, _099070_, _099071_, _099072_, _099073_, _099074_, _099075_, _099076_, _099077_, _099078_, _099079_, _099080_, _099081_, _099082_, _099083_, _099084_, _099085_, _099086_, _099087_, _099088_, _099089_, _099090_, _099091_, _099092_, _099093_, _099094_, _099095_, _099096_, _099097_, _099098_, _099099_, _099100_, _099101_, _099102_, _099103_, _099104_, _099105_, _099106_, _099107_, _099108_, _099109_, _099110_, _099111_, _099112_, _099113_, _099114_, _099115_, _099116_, _099117_, _099118_, _099119_, _099120_, _099121_, _099122_, _099123_, _099124_, _099125_, _099126_, _099127_, _099128_, _099129_, _099130_, _099131_, _099132_, _099133_, _099134_, _099135_, _099136_, _099137_, _099138_, _099139_, _099140_, _099141_, _099142_, _099143_, _099144_, _099145_, _099146_, _099147_, _099148_, _099149_, _099150_, _099151_, _099152_, _099153_, _099154_, _099155_, _099156_, _099157_, _099158_, _099159_, _099160_, _099161_, _099162_, _099163_, _099164_, _099165_, _099166_, _099167_, _099168_, _099169_, _099170_, _099171_, _099172_, _099173_, _099174_, _099175_, _099176_, _099177_, _099178_, _099179_, _099180_, _099181_, _099182_, _099183_, _099184_, _099185_, _099186_, _099187_, _099188_, _099189_, _099190_, _099191_, _099192_, _099193_, _099194_, _099195_, _099196_, _099197_, _099198_, _099199_, _099200_, _099201_, _099202_, _099203_, _099204_, _099205_, _099206_, _099207_, _099208_, _099209_, _099210_, _099211_, _099212_, _099213_, _099214_, _099215_, _099216_, _099217_, _099218_, _099219_, _099220_, _099221_, _099222_, _099223_, _099224_, _099225_, _099226_, _099227_, _099228_, _099229_, _099230_, _099231_, _099232_, _099233_, _099234_, _099235_, _099236_, _099237_, _099238_, _099239_, _099240_, _099241_, _099242_, _099243_, _099244_, _099245_, _099246_, _099247_, _099248_, _099249_, _099250_, _099251_, _099252_, _099253_, _099254_, _099255_, _099256_, _099257_, _099258_, _099259_, _099260_, _099261_, _099262_, , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , , ;
  input [479:0] set1;
  input [479:0] set2;
  input set1[0], set1[1], set1[2], set1[3], set1[4], set1[5], set1[6], set1[7], set1[8], set1[9], set1[10], set1[11], set1[12], set1[13], set1[14], set1[15], set1[16], set1[17], set1[18], set1[19], set1[20], set1[21], set1[22], set1[23], set1[24], set1[25], set1[26], set1[27], set1[28], set1[29], set1[30], set1[31], set1[32], set1[33], set1[34], set1[35], set1[36], set1[37], set1[38], set1[39], set1[40], set1[41], set1[42], set1[43], set1[44], set1[45], set1[46], set1[47], set1[48], set1[49], set1[50], set1[51], set1[52], set1[53], set1[54], set1[55], set1[56], set1[57], set1[58], set1[59], set1[60], set1[61], set1[62], set1[63], set1[64], set1[65], set1[66], set1[67], set1[68], set1[69], set1[70], set1[71], set1[72], set1[73], set1[74], set1[75], set1[76], set1[77], set1[78], set1[79], set1[80], set1[81], set1[82], set1[83], set1[84], set1[85], set1[86], set1[87], set1[88], set1[89], set1[90], set1[91], set1[92], set1[93], set1[94], set1[95], set1[96], set1[97], set1[98], set1[99], set1[100], set1[101], set1[102], set1[103], set1[104], set1[105], set1[106], set1[107], set1[108], set1[109], set1[110], set1[111], set1[112], set1[113], set1[114], set1[115], set1[116], set1[117], set1[118], set1[119], set1[120], set1[121], set1[122], set1[123], set1[124], set1[125], set1[126], set1[127], set1[128], set1[129], set1[130], set1[131], set1[132], set1[133], set1[134], set1[135], set1[136], set1[137], set1[138], set1[139], set1[140], set1[141], set1[142], set1[143], set1[144], set1[145], set1[146], set1[147], set1[148], set1[149], set1[150], set1[151], set1[152], set1[153], set1[154], set1[155], set1[156], set1[157], set1[158], set1[159], set1[160], set1[161], set1[162], set1[163], set1[164], set1[165], set1[166], set1[167], set1[168], set1[169], set1[170], set1[171], set1[172], set1[173], set1[174], set1[175], set1[176], set1[177], set1[178], set1[179], set1[180], set1[181], set1[182], set1[183], set1[184], set1[185], set1[186], set1[187], set1[188], set1[189], set1[190], set1[191], set1[192], set1[193], set1[194], set1[195], set1[196], set1[197], set1[198], set1[199], set1[200], set1[201], set1[202], set1[203], set1[204], set1[205], set1[206], set1[207], set1[208], set1[209], set1[210], set1[211], set1[212], set1[213], set1[214], set1[215], set1[216], set1[217], set1[218], set1[219], set1[220], set1[221], set1[222], set1[223], set1[224], set1[225], set1[226], set1[227], set1[228], set1[229], set1[230], set1[231], set1[232], set1[233], set1[234], set1[235], set1[236], set1[237], set1[238], set1[239], set1[240], set1[241], set1[242], set1[243], set1[244], set1[245], set1[246], set1[247], set1[248], set1[249], set1[250], set1[251], set1[252], set1[253], set1[254], set1[255], set1[256], set1[257], set1[258], set1[259], set1[260], set1[261], set1[262], set1[263], set1[264], set1[265], set1[266], set1[267], set1[268], set1[269], set1[270], set1[271], set1[272], set1[273], set1[274], set1[275], set1[276], set1[277], set1[278], set1[279], set1[280], set1[281], set1[282], set1[283], set1[284], set1[285], set1[286], set1[287], set1[288], set1[289], set1[290], set1[291], set1[292], set1[293], set1[294], set1[295], set1[296], set1[297], set1[298], set1[299], set1[300], set1[301], set1[302], set1[303], set1[304], set1[305], set1[306], set1[307], set1[308], set1[309], set1[310], set1[311], set1[312], set1[313], set1[314], set1[315], set1[316], set1[317], set1[318], set1[319], set1[320], set1[321], set1[322], set1[323], set1[324], set1[325], set1[326], set1[327], set1[328], set1[329], set1[330], set1[331], set1[332], set1[333], set1[334], set1[335], set1[336], set1[337], set1[338], set1[339], set1[340], set1[341], set1[342], set1[343], set1[344], set1[345], set1[346], set1[347], set1[348], set1[349], set1[350], set1[351], set1[352], set1[353], set1[354], set1[355], set1[356], set1[357], set1[358], set1[359], set1[360], set1[361], set1[362], set1[363], set1[364], set1[365], set1[366], set1[367], set1[368], set1[369], set1[370], set1[371], set1[372], set1[373], set1[374], set1[375], set1[376], set1[377], set1[378], set1[379], set1[380], set1[381], set1[382], set1[383], set1[384], set1[385], set1[386], set1[387], set1[388], set1[389], set1[390], set1[391], set1[392], set1[393], set1[394], set1[395], set1[396], set1[397], set1[398], set1[399], set1[400], set1[401], set1[402], set1[403], set1[404], set1[405], set1[406], set1[407], set1[408], set1[409], set1[410], set1[411], set1[412], set1[413], set1[414], set1[415], set1[416], set1[417], set1[418], set1[419], set1[420], set1[421], set1[422], set1[423], set1[424], set1[425], set1[426], set1[427], set1[428], set1[429], set1[430], set1[431], set1[432], set1[433], set1[434], set1[435], set1[436], set1[437], set1[438], set1[439], set1[440], set1[441], set1[442], set1[443], set1[444], set1[445], set1[446], set1[447], set1[448], set1[449], set1[450], set1[451], set1[452], set1[453], set1[454], set1[455], set1[456], set1[457], set1[458], set1[459], set1[460], set1[461], set1[462], set1[463], set1[464], set1[465], set1[466], set1[467], set1[468], set1[469], set1[470], set1[471], set1[472], set1[473], set1[474], set1[475], set1[476], set1[477], set1[478], set1[479], set2[0], set2[1], set2[2], set2[3], set2[4], set2[5], set2[6], set2[7], set2[8], set2[9], set2[10], set2[11], set2[12], set2[13], set2[14], set2[15], set2[16], set2[17], set2[18], set2[19], set2[20], set2[21], set2[22], set2[23], set2[24], set2[25], set2[26], set2[27], set2[28], set2[29], set2[30], set2[31], set2[32], set2[33], set2[34], set2[35], set2[36], set2[37], set2[38], set2[39], set2[40], set2[41], set2[42], set2[43], set2[44], set2[45], set2[46], set2[47], set2[48], set2[49], set2[50], set2[51], set2[52], set2[53], set2[54], set2[55], set2[56], set2[57], set2[58], set2[59], set2[60], set2[61], set2[62], set2[63], set2[64], set2[65], set2[66], set2[67], set2[68], set2[69], set2[70], set2[71], set2[72], set2[73], set2[74], set2[75], set2[76], set2[77], set2[78], set2[79], set2[80], set2[81], set2[82], set2[83], set2[84], set2[85], set2[86], set2[87], set2[88], set2[89], set2[90], set2[91], set2[92], set2[93], set2[94], set2[95], set2[96], set2[97], set2[98], set2[99], set2[100], set2[101], set2[102], set2[103], set2[104], set2[105], set2[106], set2[107], set2[108], set2[109], set2[110], set2[111], set2[112], set2[113], set2[114], set2[115], set2[116], set2[117], set2[118], set2[119], set2[120], set2[121], set2[122], set2[123], set2[124], set2[125], set2[126], set2[127], set2[128], set2[129], set2[130], set2[131], set2[132], set2[133], set2[134], set2[135], set2[136], set2[137], set2[138], set2[139], set2[140], set2[141], set2[142], set2[143], set2[144], set2[145], set2[146], set2[147], set2[148], set2[149], set2[150], set2[151], set2[152], set2[153], set2[154], set2[155], set2[156], set2[157], set2[158], set2[159], set2[160], set2[161], set2[162], set2[163], set2[164], set2[165], set2[166], set2[167], set2[168], set2[169], set2[170], set2[171], set2[172], set2[173], set2[174], set2[175], set2[176], set2[177], set2[178], set2[179], set2[180], set2[181], set2[182], set2[183], set2[184], set2[185], set2[186], set2[187], set2[188], set2[189], set2[190], set2[191], set2[192], set2[193], set2[194], set2[195], set2[196], set2[197], set2[198], set2[199], set2[200], set2[201], set2[202], set2[203], set2[204], set2[205], set2[206], set2[207], set2[208], set2[209], set2[210], set2[211], set2[212], set2[213], set2[214], set2[215], set2[216], set2[217], set2[218], set2[219], set2[220], set2[221], set2[222], set2[223], set2[224], set2[225], set2[226], set2[227], set2[228], set2[229], set2[230], set2[231], set2[232], set2[233], set2[234], set2[235], set2[236], set2[237], set2[238], set2[239], set2[240], set2[241], set2[242], set2[243], set2[244], set2[245], set2[246], set2[247], set2[248], set2[249], set2[250], set2[251], set2[252], set2[253], set2[254], set2[255], set2[256], set2[257], set2[258], set2[259], set2[260], set2[261], set2[262], set2[263], set2[264], set2[265], set2[266], set2[267], set2[268], set2[269], set2[270], set2[271], set2[272], set2[273], set2[274], set2[275], set2[276], set2[277], set2[278], set2[279], set2[280], set2[281], set2[282], set2[283], set2[284], set2[285], set2[286], set2[287], set2[288], set2[289], set2[290], set2[291], set2[292], set2[293], set2[294], set2[295], set2[296], set2[297], set2[298], set2[299], set2[300], set2[301], set2[302], set2[303], set2[304], set2[305], set2[306], set2[307], set2[308], set2[309], set2[310], set2[311], set2[312], set2[313], set2[314], set2[315], set2[316], set2[317], set2[318], set2[319], set2[320], set2[321], set2[322], set2[323], set2[324], set2[325], set2[326], set2[327], set2[328], set2[329], set2[330], set2[331], set2[332], set2[333], set2[334], set2[335], set2[336], set2[337], set2[338], set2[339], set2[340], set2[341], set2[342], set2[343], set2[344], set2[345], set2[346], set2[347], set2[348], set2[349], set2[350], set2[351], set2[352], set2[353], set2[354], set2[355], set2[356], set2[357], set2[358], set2[359], set2[360], set2[361], set2[362], set2[363], set2[364], set2[365], set2[366], set2[367], set2[368], set2[369], set2[370], set2[371], set2[372], set2[373], set2[374], set2[375], set2[376], set2[377], set2[378], set2[379], set2[380], set2[381], set2[382], set2[383], set2[384], set2[385], set2[386], set2[387], set2[388], set2[389], set2[390], set2[391], set2[392], set2[393], set2[394], set2[395], set2[396], set2[397], set2[398], set2[399], set2[400], set2[401], set2[402], set2[403], set2[404], set2[405], set2[406], set2[407], set2[408], set2[409], set2[410], set2[411], set2[412], set2[413], set2[414], set2[415], set2[416], set2[417], set2[418], set2[419], set2[420], set2[421], set2[422], set2[423], set2[424], set2[425], set2[426], set2[427], set2[428], set2[429], set2[430], set2[431], set2[432], set2[433], set2[434], set2[435], set2[436], set2[437], set2[438], set2[439], set2[440], set2[441], set2[442], set2[443], set2[444], set2[445], set2[446], set2[447], set2[448], set2[449], set2[450], set2[451], set2[452], set2[453], set2[454], set2[455], set2[456], set2[457], set2[458], set2[459], set2[460], set2[461], set2[462], set2[463], set2[464], set2[465], set2[466], set2[467], set2[468], set2[469], set2[470], set2[471], set2[472], set2[473], set2[474], set2[475], set2[476], set2[477], set2[478], set2[479];
  output out[0], out[1], out[2], out[3], out[4], out[5], out[6], out[7], out[8], out[9], out[10], out[11], out[12], out[13], out[14], out[15], out[16], out[17], out[18], out[19], out[20], out[21], out[22], out[23], out[24], out[25], out[26], out[27], out[28], out[29], out[30], out[31], out[32], out[33], out[34], out[35], out[36], out[37], out[38], out[39], out[40], out[41], out[42], out[43], out[44], out[45], out[46], out[47], out[48], out[49], out[50], out[51], out[52], out[53], out[54], out[55], out[56], out[57], out[58], out[59], out[60], out[61], out[62], out[63], out[64], out[65], out[66], out[67], out[68], out[69], out[70], out[71], out[72], out[73], out[74], out[75], out[76], out[77], out[78], out[79], out[80], out[81], out[82], out[83], out[84], out[85], out[86], out[87], out[88], out[89], out[90], out[91], out[92], out[93], out[94], out[95], out[96], out[97], out[98], out[99], out[100], out[101], out[102], out[103], out[104], out[105], out[106], out[107], out[108], out[109], out[110], out[111], out[112], out[113], out[114], out[115], out[116], out[117], out[118], out[119], out[120], out[121], out[122], out[123], out[124], out[125], out[126], out[127], out[128], out[129], out[130], out[131], out[132], out[133], out[134], out[135], out[136], out[137], out[138], out[139], out[140], out[141], out[142], out[143], out[144], out[145], out[146], out[147], out[148], out[149], out[150], out[151], out[152], out[153], out[154], out[155], out[156], out[157], out[158], out[159], out[160], out[161], out[162], out[163], out[164], out[165], out[166], out[167], out[168], out[169], out[170], out[171], out[172], out[173], out[174], out[175], out[176], out[177], out[178], out[179], out[180], out[181], out[182], out[183], out[184], out[185], out[186], out[187], out[188], out[189], out[190], out[191], out[192], out[193], out[194], out[195], out[196], out[197], out[198], out[199], out[200], out[201], out[202], out[203], out[204], out[205], out[206], out[207], out[208], out[209], out[210], out[211], out[212], out[213], out[214], out[215], out[216], out[217], out[218], out[219], out[220], out[221], out[222], out[223], out[224], out[225], out[226], out[227], out[228], out[229], out[230], out[231], out[232], out[233], out[234], out[235], out[236], out[237], out[238], out[239], out[240], out[241], out[242], out[243], out[244], out[245], out[246], out[247], out[248], out[249], out[250], out[251], out[252], out[253], out[254], out[255], out[256], out[257], out[258], out[259], out[260], out[261], out[262], out[263], out[264], out[265], out[266], out[267], out[268], out[269], out[270], out[271], out[272], out[273], out[274], out[275], out[276], out[277], out[278], out[279], out[280], out[281], out[282], out[283], out[284], out[285], out[286], out[287], out[288], out[289], out[290], out[291], out[292], out[293], out[294], out[295], out[296], out[297], out[298], out[299], out[300], out[301], out[302], out[303], out[304], out[305], out[306], out[307], out[308], out[309], out[310], out[311], out[312], out[313], out[314], out[315], out[316], out[317], out[318], out[319], out[320], out[321], out[322], out[323], out[324], out[325], out[326], out[327], out[328], out[329], out[330], out[331], out[332], out[333], out[334], out[335], out[336], out[337], out[338], out[339], out[340], out[341], out[342], out[343], out[344], out[345], out[346], out[347], out[348], out[349], out[350], out[351], out[352], out[353], out[354], out[355], out[356], out[357], out[358], out[359], out[360], out[361], out[362], out[363], out[364], out[365], out[366], out[367], out[368], out[369], out[370], out[371], out[372], out[373], out[374], out[375], out[376], out[377], out[378], out[379], out[380], out[381], out[382], out[383], out[384], out[385], out[386], out[387], out[388], out[389], out[390], out[391], out[392], out[393], out[394], out[395], out[396], out[397], out[398], out[399], out[400], out[401], out[402], out[403], out[404], out[405], out[406], out[407], out[408], out[409], out[410], out[411], out[412], out[413], out[414], out[415], out[416], out[417], out[418], out[419], out[420], out[421], out[422], out[423], out[424], out[425], out[426], out[427], out[428], out[429], out[430], out[431], out[432], out[433], out[434], out[435], out[436], out[437], out[438], out[439], out[440], out[441], out[442], out[443], out[444], out[445], out[446], out[447], out[448], out[449], out[450], out[451], out[452], out[453], out[454], out[455], out[456], out[457], out[458], out[459], out[460], out[461], out[462], out[463], out[464], out[465], out[466], out[467], out[468], out[469], out[470], out[471], out[472], out[473], out[474], out[475], out[476], out[477], out[478], out[479], out[480], out[481], out[482], out[483], out[484], out[485], out[486], out[487], out[488], out[489], out[490], out[491], out[492], out[493], out[494], out[495], out[496], out[497], out[498], out[499], out[500], out[501], out[502], out[503], out[504], out[505], out[506], out[507], out[508], out[509], out[510], out[511], out[512], out[513], out[514], out[515], out[516], out[517], out[518], out[519], out[520], out[521], out[522], out[523], out[524], out[525], out[526], out[527], out[528], out[529], out[530], out[531], out[532], out[533], out[534], out[535], out[536], out[537], out[538], out[539], out[540], out[541], out[542], out[543], out[544], out[545], out[546], out[547], out[548], out[549], out[550], out[551], out[552], out[553], out[554], out[555], out[556], out[557], out[558], out[559], out[560], out[561], out[562], out[563], out[564], out[565], out[566], out[567], out[568], out[569], out[570], out[571], out[572], out[573], out[574], out[575], out[576], out[577], out[578], out[579], out[580], out[581], out[582], out[583], out[584], out[585], out[586], out[587], out[588], out[589], out[590], out[591], out[592], out[593], out[594], out[595], out[596], out[597], out[598], out[599], out[600], out[601], out[602], out[603], out[604], out[605], out[606], out[607], out[608], out[609], out[610], out[611], out[612], out[613], out[614], out[615], out[616], out[617], out[618], out[619], out[620], out[621], out[622], out[623], out[624], out[625], out[626], out[627], out[628], out[629], out[630], out[631], out[632], out[633], out[634], out[635], out[636], out[637], out[638], out[639], out[640], out[641], out[642], out[643], out[644], out[645], out[646], out[647], out[648], out[649], out[650], out[651], out[652], out[653], out[654], out[655], out[656], out[657], out[658], out[659], out[660], out[661], out[662], out[663], out[664], out[665], out[666], out[667], out[668], out[669], out[670], out[671], out[672], out[673], out[674], out[675], out[676], out[677], out[678], out[679], out[680], out[681], out[682], out[683], out[684], out[685], out[686], out[687], out[688], out[689], out[690], out[691], out[692], out[693], out[694], out[695], out[696], out[697], out[698], out[699], out[700], out[701], out[702], out[703], out[704], out[705], out[706], out[707], out[708], out[709], out[710], out[711], out[712], out[713], out[714], out[715], out[716], out[717], out[718], out[719], out[720], out[721], out[722], out[723], out[724], out[725], out[726], out[727], out[728], out[729], out[730], out[731], out[732], out[733], out[734], out[735], out[736], out[737], out[738], out[739], out[740], out[741], out[742], out[743], out[744], out[745], out[746], out[747], out[748], out[749], out[750], out[751], out[752], out[753], out[754], out[755], out[756], out[757], out[758], out[759], out[760], out[761], out[762], out[763], out[764], out[765], out[766], out[767], out[768], out[769], out[770], out[771], out[772], out[773], out[774], out[775], out[776], out[777], out[778], out[779], out[780], out[781], out[782], out[783], out[784], out[785], out[786], out[787], out[788], out[789], out[790], out[791], out[792], out[793], out[794], out[795], out[796], out[797], out[798], out[799], out[800], out[801], out[802], out[803], out[804], out[805], out[806], out[807], out[808], out[809], out[810], out[811], out[812], out[813], out[814], out[815], out[816], out[817], out[818], out[819], out[820], out[821], out[822], out[823], out[824], out[825], out[826], out[827], out[828], out[829], out[830], out[831], out[832], out[833], out[834], out[835], out[836], out[837], out[838], out[839], out[840], out[841], out[842], out[843], out[844], out[845], out[846], out[847], out[848], out[849], out[850], out[851], out[852], out[853], out[854], out[855], out[856], out[857], out[858], out[859], out[860], out[861], out[862], out[863], out[864], out[865], out[866], out[867], out[868], out[869], out[870], out[871], out[872], out[873], out[874], out[875], out[876], out[877], out[878], out[879], out[880], out[881], out[882], out[883], out[884], out[885], out[886], out[887], out[888], out[889], out[890], out[891], out[892], out[893], out[894], out[895], out[896], out[897], out[898], out[899], out[900], out[901], out[902], out[903], out[904], out[905], out[906], out[907], out[908], out[909], out[910], out[911], out[912], out[913], out[914], out[915], out[916], out[917], out[918], out[919], out[920], out[921], out[922], out[923], out[924], out[925], out[926], out[927], out[928], out[929], out[930], out[931], out[932], out[933], out[934], out[935], out[936], out[937], out[938], out[939], out[940], out[941], out[942], out[943], out[944], out[945], out[946], out[947], out[948], out[949], out[950], out[951], out[952], out[953], out[954], out[955], out[956], out[957], out[958], out[959], out[960], out[961], out[962], out[963], out[964], out[965], out[966], out[967];
  not g_099263_(out[481], _097964_);
  not g_099264_(out[482], _097975_);
  not g_099265_(out[487], _097986_);
  not g_099266_(out[7], _097997_);
  not g_099267_(out[488], _098008_);
  not g_099268_(out[489], _098019_);
  not g_099269_(out[491], _098030_);
  not g_099270_(out[11], _098041_);
  not g_099271_(out[492], _098052_);
  not g_099272_(out[27], _098063_);
  not g_099273_(out[28], _098074_);
  not g_099274_(out[39], _098085_);
  not g_099275_(out[43], _098096_);
  not g_099276_(out[59], _098107_);
  not g_099277_(out[75], _098118_);
  not g_099278_(out[91], _098129_);
  not g_099279_(out[107], _098140_);
  not g_099280_(out[123], _098151_);
  not g_099281_(out[139], _098162_);
  not g_099282_(out[155], _098173_);
  not g_099283_(out[171], _098184_);
  not g_099284_(out[187], _098195_);
  not g_099285_(out[203], _098206_);
  not g_099286_(out[219], _098217_);
  not g_099287_(out[235], _098228_);
  not g_099288_(out[251], _098239_);
  not g_099289_(out[267], _098250_);
  not g_099290_(out[283], _098261_);
  not g_099291_(out[299], _098272_);
  not g_099292_(out[315], _098283_);
  not g_099293_(out[331], _098294_);
  not g_099294_(out[347], _049400_);
  not g_099295_(out[363], _049411_);
  not g_099296_(out[379], _049422_);
  not g_099297_(out[395], _049433_);
  not g_099298_(out[411], _049444_);
  not g_099299_(out[427], _049455_);
  not g_099300_(out[443], _049466_);
  not g_099301_(out[459], _049477_);
  not g_099302_(out[471], _049488_);
  not g_099303_(out[475], _049499_);
  not g_099304_(out[507], _049510_);
  not g_099305_(out[523], _049521_);
  not g_099306_(out[539], _049532_);
  not g_099307_(out[555], _049543_);
  not g_099308_(out[571], _049554_);
  not g_099309_(out[587], _049565_);
  not g_099310_(out[603], _049576_);
  not g_099311_(out[619], _049587_);
  not g_099312_(out[635], _049598_);
  not g_099313_(out[651], _049609_);
  not g_099314_(out[667], _049620_);
  not g_099315_(out[683], _049631_);
  not g_099316_(out[699], _049642_);
  not g_099317_(out[715], _049653_);
  not g_099318_(out[731], _049664_);
  not g_099319_(out[747], _049675_);
  not g_099320_(out[763], _049686_);
  not g_099321_(out[779], _049697_);
  not g_099322_(out[795], _049708_);
  not g_099323_(out[811], _049719_);
  not g_099324_(out[827], _049730_);
  not g_099325_(out[843], _049741_);
  not g_099326_(out[859], _049752_);
  not g_099327_(out[875], _049763_);
  not g_099328_(out[891], _049774_);
  not g_099329_(out[907], _049785_);
  not g_099330_(out[923], _049796_);
  not g_099331_(out[939], _049807_);
  not g_099332_(out[951], _049818_);
  not g_099333_(out[955], _049829_);
  xor g_099334_(out[473], out[953], _049840_);
  and g_099335_(_049488_, out[951], _049851_);
  and g_099336_(out[471], _049818_, _049862_);
  xor g_099337_(out[467], out[947], _049873_);
  xor g_099338_(out[477], out[957], _049884_);
  xor g_099339_(out[470], out[950], _049895_);
  xor g_099340_(out[474], out[954], _049906_);
  or g_099341_(_049895_, _049906_, _049917_);
  xor g_099342_(out[469], out[949], _049928_);
  xor g_099343_(out[465], out[945], _049939_);
  xor g_099344_(out[475], out[955], _049950_);
  xor g_099345_(out[464], out[944], _049961_);
  xor g_099346_(out[472], out[952], _049972_);
  xor g_099347_(out[476], out[956], _049983_);
  xor g_099348_(out[468], out[948], _049994_);
  or g_099349_(_049873_, _049994_, _050005_);
  xor g_099350_(out[478], out[958], _050016_);
  or g_099351_(_049917_, _050005_, _050027_);
  or g_099352_(_049928_, _049950_, _050038_);
  or g_099353_(_049884_, _050038_, _050049_);
  or g_099354_(_050027_, _050049_, _050060_);
  or g_099355_(_049961_, _049983_, _050071_);
  or g_099356_(_050060_, _050071_, _050082_);
  xor g_099357_(out[466], out[946], _050093_);
  or g_099358_(_049851_, _050093_, _050104_);
  xor g_099359_(out[479], out[959], _050115_);
  or g_099360_(_050016_, _050115_, _050126_);
  or g_099361_(_050104_, _050126_, _050137_);
  or g_099362_(_049840_, _049862_, _050148_);
  or g_099363_(_049939_, _050148_, _050159_);
  or g_099364_(_050137_, _050159_, _050170_);
  or g_099365_(_049972_, _050170_, _050181_);
  or g_099366_(_050082_, _050181_, _050192_);
  xor g_099367_(out[455], out[951], _050203_);
  and g_099368_(_049477_, out[955], _050214_);
  xor g_099369_(out[462], out[958], _050225_);
  xor g_099370_(out[456], out[952], _050236_);
  xor g_099371_(out[449], out[945], _050247_);
  xor g_099372_(out[461], out[957], _050258_);
  xor g_099373_(out[457], out[953], _050269_);
  xor g_099374_(out[452], out[948], _050280_);
  xor g_099375_(out[450], out[946], _050291_);
  and g_099376_(out[459], _049829_, _050302_);
  xor g_099377_(out[451], out[947], _050313_);
  xor g_099378_(out[454], out[950], _050324_);
  xor g_099379_(out[463], out[959], _050335_);
  xor g_099380_(out[458], out[954], _050346_);
  xor g_099381_(out[453], out[949], _050357_);
  xor g_099382_(out[448], out[944], _050368_);
  or g_099383_(_050225_, _050280_, _050379_);
  or g_099384_(_050236_, _050258_, _050390_);
  or g_099385_(_050291_, _050346_, _050401_);
  or g_099386_(_050390_, _050401_, _050412_);
  or g_099387_(_050269_, _050313_, _050423_);
  or g_099388_(_050357_, _050368_, _050434_);
  or g_099389_(_050423_, _050434_, _050445_);
  or g_099390_(_050412_, _050445_, _050456_);
  xor g_099391_(out[460], out[956], _050467_);
  or g_099392_(_050214_, _050467_, _050478_);
  or g_099393_(_050203_, _050324_, _050489_);
  or g_099394_(_050478_, _050489_, _050500_);
  or g_099395_(_050247_, _050302_, _050511_);
  or g_099396_(_050335_, _050511_, _050522_);
  or g_099397_(_050500_, _050522_, _050533_);
  or g_099398_(_050456_, _050533_, _050544_);
  or g_099399_(_050379_, _050544_, _050555_);
  xor g_099400_(out[433], out[945], _050566_);
  and g_099401_(out[443], _049829_, _050577_);
  xor g_099402_(out[446], out[958], _050588_);
  xor g_099403_(out[435], out[947], _050599_);
  xor g_099404_(out[436], out[948], _050610_);
  xor g_099405_(out[434], out[946], _050621_);
  xor g_099406_(out[441], out[953], _050632_);
  xor g_099407_(out[432], out[944], _050643_);
  and g_099408_(_049466_, out[955], _050654_);
  xor g_099409_(out[438], out[950], _050665_);
  xor g_099410_(out[442], out[954], _050676_);
  xor g_099411_(out[437], out[949], _050687_);
  xor g_099412_(out[447], out[959], _050698_);
  xor g_099413_(out[445], out[957], _050709_);
  xor g_099414_(out[440], out[952], _050720_);
  or g_099415_(_050588_, _050610_, _050731_);
  or g_099416_(_050709_, _050720_, _050742_);
  or g_099417_(_050621_, _050676_, _050753_);
  or g_099418_(_050742_, _050753_, _050764_);
  or g_099419_(_050599_, _050632_, _050775_);
  or g_099420_(_050643_, _050687_, _050786_);
  or g_099421_(_050775_, _050786_, _050797_);
  or g_099422_(_050764_, _050797_, _050808_);
  xor g_099423_(out[444], out[956], _050819_);
  or g_099424_(_050654_, _050819_, _050830_);
  xor g_099425_(out[439], out[951], _050841_);
  or g_099426_(_050665_, _050841_, _050852_);
  or g_099427_(_050830_, _050852_, _050863_);
  or g_099428_(_050566_, _050577_, _050874_);
  or g_099429_(_050698_, _050874_, _050885_);
  or g_099430_(_050863_, _050885_, _050896_);
  or g_099431_(_050808_, _050896_, _050907_);
  or g_099432_(_050731_, _050907_, _050918_);
  xor g_099433_(out[423], out[951], _050929_);
  and g_099434_(_049455_, out[955], _050940_);
  xor g_099435_(out[430], out[958], _050951_);
  xor g_099436_(out[424], out[952], _050962_);
  xor g_099437_(out[417], out[945], _050973_);
  xor g_099438_(out[429], out[957], _050984_);
  xor g_099439_(out[425], out[953], _050995_);
  xor g_099440_(out[420], out[948], _051006_);
  xor g_099441_(out[418], out[946], _051017_);
  and g_099442_(out[427], _049829_, _051028_);
  xor g_099443_(out[419], out[947], _051039_);
  xor g_099444_(out[422], out[950], _051050_);
  xor g_099445_(out[431], out[959], _051061_);
  xor g_099446_(out[426], out[954], _051072_);
  xor g_099447_(out[421], out[949], _051083_);
  xor g_099448_(out[416], out[944], _051094_);
  or g_099449_(_050951_, _051006_, _051105_);
  or g_099450_(_050962_, _050984_, _051116_);
  or g_099451_(_051017_, _051072_, _051127_);
  or g_099452_(_051116_, _051127_, _051138_);
  or g_099453_(_050995_, _051039_, _051149_);
  or g_099454_(_051083_, _051094_, _051160_);
  or g_099455_(_051149_, _051160_, _051171_);
  or g_099456_(_051138_, _051171_, _051182_);
  xor g_099457_(out[428], out[956], _051193_);
  or g_099458_(_050940_, _051193_, _051204_);
  or g_099459_(_050929_, _051050_, _051215_);
  or g_099460_(_051204_, _051215_, _051226_);
  or g_099461_(_050973_, _051028_, _051237_);
  or g_099462_(_051061_, _051237_, _051248_);
  or g_099463_(_051226_, _051248_, _051259_);
  or g_099464_(_051182_, _051259_, _051270_);
  or g_099465_(_051105_, _051270_, _051281_);
  xor g_099466_(out[408], out[952], _051292_);
  xor g_099467_(out[405], out[949], _051303_);
  xor g_099468_(out[403], out[947], _051314_);
  xor g_099469_(out[414], out[958], _051325_);
  xor g_099470_(out[413], out[957], _051336_);
  xor g_099471_(out[402], out[946], _051347_);
  xor g_099472_(out[409], out[953], _051358_);
  xor g_099473_(out[406], out[950], _051369_);
  xor g_099474_(out[415], out[959], _051380_);
  xor g_099475_(out[410], out[954], _051391_);
  xor g_099476_(out[404], out[948], _051402_);
  xor g_099477_(out[400], out[944], _051413_);
  and g_099478_(_049444_, out[955], _051424_);
  and g_099479_(out[411], _049829_, _051435_);
  or g_099480_(_051292_, _051336_, _051446_);
  xor g_099481_(out[401], out[945], _051457_);
  or g_099482_(_051347_, _051391_, _051468_);
  or g_099483_(_051446_, _051468_, _051479_);
  or g_099484_(_051314_, _051358_, _051490_);
  or g_099485_(_051303_, _051490_, _051501_);
  or g_099486_(_051479_, _051501_, _051512_);
  or g_099487_(_051325_, _051402_, _051523_);
  or g_099488_(_051512_, _051523_, _051534_);
  xor g_099489_(out[412], out[956], _051545_);
  or g_099490_(_051424_, _051545_, _051556_);
  xor g_099491_(out[407], out[951], _051567_);
  or g_099492_(_051369_, _051567_, _051578_);
  or g_099493_(_051556_, _051578_, _051589_);
  or g_099494_(_051435_, _051457_, _051600_);
  or g_099495_(_051380_, _051600_, _051611_);
  or g_099496_(_051589_, _051611_, _051622_);
  or g_099497_(_051413_, _051622_, _051633_);
  or g_099498_(_051534_, _051633_, _051644_);
  xor g_099499_(out[391], out[951], _051655_);
  and g_099500_(_049433_, out[955], _051666_);
  xor g_099501_(out[398], out[958], _051677_);
  xor g_099502_(out[392], out[952], _051688_);
  xor g_099503_(out[385], out[945], _051699_);
  xor g_099504_(out[397], out[957], _051710_);
  xor g_099505_(out[393], out[953], _051721_);
  xor g_099506_(out[388], out[948], _051732_);
  xor g_099507_(out[386], out[946], _051743_);
  and g_099508_(out[395], _049829_, _051754_);
  xor g_099509_(out[387], out[947], _051765_);
  xor g_099510_(out[390], out[950], _051776_);
  xor g_099511_(out[399], out[959], _051787_);
  xor g_099512_(out[394], out[954], _051798_);
  xor g_099513_(out[389], out[949], _051809_);
  xor g_099514_(out[384], out[944], _051820_);
  or g_099515_(_051677_, _051732_, _051831_);
  or g_099516_(_051688_, _051710_, _051842_);
  or g_099517_(_051743_, _051798_, _051853_);
  or g_099518_(_051842_, _051853_, _051864_);
  or g_099519_(_051721_, _051765_, _051875_);
  or g_099520_(_051809_, _051820_, _051886_);
  or g_099521_(_051875_, _051886_, _051897_);
  or g_099522_(_051864_, _051897_, _051908_);
  xor g_099523_(out[396], out[956], _051919_);
  or g_099524_(_051666_, _051919_, _051930_);
  or g_099525_(_051655_, _051776_, _051941_);
  or g_099526_(_051930_, _051941_, _051952_);
  or g_099527_(_051699_, _051754_, _051963_);
  or g_099528_(_051787_, _051963_, _051974_);
  or g_099529_(_051952_, _051974_, _051985_);
  or g_099530_(_051908_, _051985_, _051996_);
  or g_099531_(_051831_, _051996_, _052007_);
  xor g_099532_(out[369], out[945], _052018_);
  and g_099533_(out[379], _049829_, _052029_);
  xor g_099534_(out[382], out[958], _052040_);
  xor g_099535_(out[371], out[947], _052051_);
  xor g_099536_(out[372], out[948], _052062_);
  xor g_099537_(out[370], out[946], _052073_);
  xor g_099538_(out[377], out[953], _052084_);
  xor g_099539_(out[368], out[944], _052095_);
  and g_099540_(_049422_, out[955], _052106_);
  xor g_099541_(out[374], out[950], _052117_);
  xor g_099542_(out[378], out[954], _052128_);
  xor g_099543_(out[373], out[949], _052139_);
  xor g_099544_(out[383], out[959], _052150_);
  xor g_099545_(out[381], out[957], _052161_);
  xor g_099546_(out[376], out[952], _052172_);
  or g_099547_(_052040_, _052062_, _052183_);
  or g_099548_(_052161_, _052172_, _052194_);
  or g_099549_(_052073_, _052128_, _052205_);
  or g_099550_(_052194_, _052205_, _052216_);
  or g_099551_(_052051_, _052084_, _052227_);
  or g_099552_(_052095_, _052139_, _052238_);
  or g_099553_(_052227_, _052238_, _052249_);
  or g_099554_(_052216_, _052249_, _052260_);
  xor g_099555_(out[380], out[956], _052271_);
  or g_099556_(_052106_, _052271_, _052282_);
  xor g_099557_(out[375], out[951], _052293_);
  or g_099558_(_052117_, _052293_, _052304_);
  or g_099559_(_052282_, _052304_, _052315_);
  or g_099560_(_052018_, _052029_, _052326_);
  or g_099561_(_052150_, _052326_, _052337_);
  or g_099562_(_052315_, _052337_, _052348_);
  or g_099563_(_052260_, _052348_, _052359_);
  or g_099564_(_052183_, _052359_, _052370_);
  xor g_099565_(out[359], out[951], _052381_);
  and g_099566_(_049411_, out[955], _052392_);
  xor g_099567_(out[366], out[958], _052403_);
  xor g_099568_(out[360], out[952], _052414_);
  xor g_099569_(out[353], out[945], _052425_);
  xor g_099570_(out[365], out[957], _052436_);
  xor g_099571_(out[361], out[953], _052447_);
  xor g_099572_(out[356], out[948], _052458_);
  xor g_099573_(out[354], out[946], _052469_);
  and g_099574_(out[363], _049829_, _052480_);
  xor g_099575_(out[355], out[947], _052491_);
  xor g_099576_(out[358], out[950], _052502_);
  xor g_099577_(out[367], out[959], _052513_);
  xor g_099578_(out[362], out[954], _052524_);
  xor g_099579_(out[357], out[949], _052535_);
  xor g_099580_(out[352], out[944], _052546_);
  or g_099581_(_052403_, _052458_, _052557_);
  or g_099582_(_052414_, _052436_, _052568_);
  or g_099583_(_052469_, _052524_, _052579_);
  or g_099584_(_052568_, _052579_, _052590_);
  or g_099585_(_052447_, _052491_, _052601_);
  or g_099586_(_052535_, _052546_, _052612_);
  or g_099587_(_052601_, _052612_, _052623_);
  or g_099588_(_052590_, _052623_, _052634_);
  xor g_099589_(out[364], out[956], _052645_);
  or g_099590_(_052392_, _052645_, _052656_);
  or g_099591_(_052381_, _052502_, _052667_);
  or g_099592_(_052656_, _052667_, _052678_);
  or g_099593_(_052425_, _052480_, _052689_);
  or g_099594_(_052513_, _052689_, _052700_);
  or g_099595_(_052678_, _052700_, _052711_);
  or g_099596_(_052634_, _052711_, _052722_);
  or g_099597_(_052557_, _052722_, _052733_);
  xor g_099598_(out[337], out[945], _052744_);
  and g_099599_(out[347], _049829_, _052755_);
  xor g_099600_(out[345], out[953], _052766_);
  xor g_099601_(out[336], out[944], _052777_);
  xor g_099602_(out[350], out[958], _052788_);
  xor g_099603_(out[340], out[948], _052799_);
  or g_099604_(_052788_, _052799_, _052810_);
  xor g_099605_(out[349], out[957], _052821_);
  xor g_099606_(out[339], out[947], _052832_);
  and g_099607_(_049400_, out[955], _052843_);
  xor g_099608_(out[342], out[950], _052854_);
  xor g_099609_(out[346], out[954], _052865_);
  xor g_099610_(out[341], out[949], _052876_);
  xor g_099611_(out[351], out[959], _052887_);
  xor g_099612_(out[344], out[952], _052898_);
  or g_099613_(_052821_, _052898_, _052909_);
  xor g_099614_(out[338], out[946], _052920_);
  or g_099615_(_052865_, _052920_, _052931_);
  or g_099616_(_052909_, _052931_, _052942_);
  or g_099617_(_052766_, _052832_, _052953_);
  or g_099618_(_052876_, _052953_, _052964_);
  or g_099619_(_052942_, _052964_, _052975_);
  or g_099620_(_052810_, _052975_, _052986_);
  xor g_099621_(out[348], out[956], _052997_);
  or g_099622_(_052843_, _052997_, _053008_);
  xor g_099623_(out[343], out[951], _053019_);
  or g_099624_(_052854_, _053019_, _053030_);
  or g_099625_(_053008_, _053030_, _053041_);
  or g_099626_(_052744_, _052755_, _053052_);
  or g_099627_(_052887_, _053052_, _053063_);
  or g_099628_(_053041_, _053063_, _053074_);
  or g_099629_(_052777_, _053074_, _053085_);
  or g_099630_(_052986_, _053085_, _053096_);
  xor g_099631_(out[327], out[951], _053107_);
  and g_099632_(_098294_, out[955], _053118_);
  xor g_099633_(out[334], out[958], _053129_);
  xor g_099634_(out[328], out[952], _053140_);
  xor g_099635_(out[321], out[945], _053151_);
  xor g_099636_(out[333], out[957], _053162_);
  xor g_099637_(out[329], out[953], _053173_);
  xor g_099638_(out[324], out[948], _053184_);
  xor g_099639_(out[322], out[946], _053195_);
  and g_099640_(out[331], _049829_, _053206_);
  xor g_099641_(out[323], out[947], _053217_);
  xor g_099642_(out[326], out[950], _053228_);
  xor g_099643_(out[335], out[959], _053239_);
  xor g_099644_(out[330], out[954], _053250_);
  xor g_099645_(out[325], out[949], _053261_);
  xor g_099646_(out[320], out[944], _053272_);
  or g_099647_(_053129_, _053184_, _053283_);
  or g_099648_(_053140_, _053162_, _053294_);
  or g_099649_(_053195_, _053250_, _053305_);
  or g_099650_(_053294_, _053305_, _053316_);
  or g_099651_(_053173_, _053217_, _053327_);
  or g_099652_(_053261_, _053272_, _053338_);
  or g_099653_(_053327_, _053338_, _053349_);
  or g_099654_(_053316_, _053349_, _053360_);
  xor g_099655_(out[332], out[956], _053371_);
  or g_099656_(_053118_, _053371_, _053382_);
  or g_099657_(_053107_, _053228_, _053393_);
  or g_099658_(_053382_, _053393_, _053404_);
  or g_099659_(_053151_, _053206_, _053415_);
  or g_099660_(_053239_, _053415_, _053426_);
  or g_099661_(_053404_, _053426_, _053437_);
  or g_099662_(_053360_, _053437_, _053448_);
  or g_099663_(_053283_, _053448_, _053459_);
  xor g_099664_(out[316], out[956], _053470_);
  and g_099665_(_098283_, out[955], _053481_);
  xor g_099666_(out[312], out[952], _053492_);
  xor g_099667_(out[310], out[950], _053503_);
  xor g_099668_(out[317], out[957], _053514_);
  xor g_099669_(out[318], out[958], _053525_);
  xor g_099670_(out[306], out[946], _053536_);
  xor g_099671_(out[313], out[953], _053547_);
  xor g_099672_(out[309], out[949], _053558_);
  xor g_099673_(out[305], out[945], _053569_);
  and g_099674_(out[315], _049829_, _053580_);
  or g_099675_(_053492_, _053514_, _053591_);
  xor g_099676_(out[319], out[959], _053602_);
  xor g_099677_(out[314], out[954], _053613_);
  xor g_099678_(out[308], out[948], _053624_);
  xor g_099679_(out[307], out[947], _053635_);
  xor g_099680_(out[304], out[944], _053646_);
  or g_099681_(_053536_, _053613_, _053657_);
  or g_099682_(_053591_, _053657_, _053668_);
  or g_099683_(_053547_, _053635_, _053679_);
  or g_099684_(_053558_, _053679_, _053690_);
  or g_099685_(_053668_, _053690_, _053701_);
  or g_099686_(_053525_, _053624_, _053712_);
  or g_099687_(_053701_, _053712_, _053723_);
  or g_099688_(_053470_, _053481_, _053734_);
  xor g_099689_(out[311], out[951], _053745_);
  or g_099690_(_053503_, _053745_, _053756_);
  or g_099691_(_053734_, _053756_, _053767_);
  or g_099692_(_053569_, _053580_, _053778_);
  or g_099693_(_053602_, _053778_, _053789_);
  or g_099694_(_053767_, _053789_, _053800_);
  or g_099695_(_053646_, _053800_, _053811_);
  or g_099696_(_053723_, _053811_, _053822_);
  xor g_099697_(out[295], out[951], _053833_);
  and g_099698_(_098272_, out[955], _053844_);
  xor g_099699_(out[302], out[958], _053855_);
  xor g_099700_(out[296], out[952], _053866_);
  xor g_099701_(out[289], out[945], _053877_);
  xor g_099702_(out[301], out[957], _053888_);
  xor g_099703_(out[297], out[953], _053899_);
  xor g_099704_(out[292], out[948], _053910_);
  xor g_099705_(out[290], out[946], _053921_);
  and g_099706_(out[299], _049829_, _053932_);
  xor g_099707_(out[291], out[947], _053943_);
  xor g_099708_(out[294], out[950], _053954_);
  xor g_099709_(out[303], out[959], _053965_);
  xor g_099710_(out[298], out[954], _053976_);
  xor g_099711_(out[293], out[949], _053987_);
  xor g_099712_(out[288], out[944], _053998_);
  or g_099713_(_053855_, _053910_, _054009_);
  or g_099714_(_053866_, _053888_, _054020_);
  or g_099715_(_053921_, _053976_, _054031_);
  or g_099716_(_054020_, _054031_, _054042_);
  or g_099717_(_053899_, _053943_, _054053_);
  or g_099718_(_053987_, _053998_, _054064_);
  or g_099719_(_054053_, _054064_, _054075_);
  or g_099720_(_054042_, _054075_, _054086_);
  xor g_099721_(out[300], out[956], _054097_);
  or g_099722_(_053844_, _054097_, _054108_);
  or g_099723_(_053833_, _053954_, _054119_);
  or g_099724_(_054108_, _054119_, _054130_);
  or g_099725_(_053877_, _053932_, _054141_);
  or g_099726_(_053965_, _054141_, _054152_);
  or g_099727_(_054130_, _054152_, _054163_);
  or g_099728_(_054086_, _054163_, _054174_);
  or g_099729_(_054009_, _054174_, _054185_);
  xor g_099730_(out[273], out[945], _054196_);
  and g_099731_(out[283], _049829_, _054207_);
  xor g_099732_(out[286], out[958], _054218_);
  xor g_099733_(out[275], out[947], _054229_);
  xor g_099734_(out[276], out[948], _054240_);
  xor g_099735_(out[274], out[946], _054251_);
  xor g_099736_(out[281], out[953], _054262_);
  xor g_099737_(out[272], out[944], _054273_);
  and g_099738_(_098261_, out[955], _054284_);
  xor g_099739_(out[278], out[950], _054295_);
  xor g_099740_(out[282], out[954], _054306_);
  xor g_099741_(out[277], out[949], _054317_);
  xor g_099742_(out[287], out[959], _054328_);
  xor g_099743_(out[285], out[957], _054339_);
  xor g_099744_(out[280], out[952], _054350_);
  or g_099745_(_054218_, _054240_, _054361_);
  or g_099746_(_054339_, _054350_, _054372_);
  or g_099747_(_054251_, _054306_, _054383_);
  or g_099748_(_054372_, _054383_, _054394_);
  or g_099749_(_054229_, _054262_, _054405_);
  or g_099750_(_054273_, _054317_, _054416_);
  or g_099751_(_054405_, _054416_, _054427_);
  or g_099752_(_054394_, _054427_, _054438_);
  xor g_099753_(out[284], out[956], _054449_);
  or g_099754_(_054284_, _054449_, _054460_);
  xor g_099755_(out[279], out[951], _054471_);
  or g_099756_(_054295_, _054471_, _054482_);
  or g_099757_(_054460_, _054482_, _054493_);
  or g_099758_(_054196_, _054207_, _054504_);
  or g_099759_(_054328_, _054504_, _054515_);
  or g_099760_(_054493_, _054515_, _054526_);
  or g_099761_(_054438_, _054526_, _054537_);
  or g_099762_(_054361_, _054537_, _054548_);
  xor g_099763_(out[263], out[951], _054559_);
  and g_099764_(_098250_, out[955], _054570_);
  xor g_099765_(out[270], out[958], _054581_);
  xor g_099766_(out[264], out[952], _054592_);
  xor g_099767_(out[257], out[945], _054603_);
  xor g_099768_(out[269], out[957], _054614_);
  xor g_099769_(out[265], out[953], _054625_);
  xor g_099770_(out[260], out[948], _054636_);
  xor g_099771_(out[258], out[946], _054647_);
  and g_099772_(out[267], _049829_, _054658_);
  xor g_099773_(out[259], out[947], _054669_);
  xor g_099774_(out[262], out[950], _054680_);
  xor g_099775_(out[271], out[959], _054691_);
  xor g_099776_(out[266], out[954], _054702_);
  xor g_099777_(out[261], out[949], _054713_);
  xor g_099778_(out[256], out[944], _054724_);
  or g_099779_(_054581_, _054636_, _054735_);
  or g_099780_(_054592_, _054614_, _054746_);
  or g_099781_(_054647_, _054702_, _054757_);
  or g_099782_(_054746_, _054757_, _054768_);
  or g_099783_(_054625_, _054669_, _054779_);
  or g_099784_(_054713_, _054724_, _054790_);
  or g_099785_(_054779_, _054790_, _054801_);
  or g_099786_(_054768_, _054801_, _054812_);
  xor g_099787_(out[268], out[956], _054823_);
  or g_099788_(_054570_, _054823_, _054834_);
  or g_099789_(_054559_, _054680_, _054845_);
  or g_099790_(_054834_, _054845_, _054856_);
  or g_099791_(_054603_, _054658_, _054867_);
  or g_099792_(_054691_, _054867_, _054878_);
  or g_099793_(_054856_, _054878_, _054889_);
  or g_099794_(_054812_, _054889_, _054900_);
  or g_099795_(_054735_, _054900_, _054911_);
  xor g_099796_(out[252], out[956], _054922_);
  and g_099797_(_098239_, out[955], _054933_);
  xor g_099798_(out[248], out[952], _054944_);
  xor g_099799_(out[246], out[950], _054955_);
  xor g_099800_(out[253], out[957], _054966_);
  xor g_099801_(out[254], out[958], _054977_);
  xor g_099802_(out[242], out[946], _054988_);
  xor g_099803_(out[249], out[953], _054999_);
  xor g_099804_(out[245], out[949], _055010_);
  xor g_099805_(out[241], out[945], _055021_);
  and g_099806_(out[251], _049829_, _055032_);
  or g_099807_(_054944_, _054966_, _055043_);
  xor g_099808_(out[255], out[959], _055054_);
  xor g_099809_(out[250], out[954], _055065_);
  xor g_099810_(out[244], out[948], _055076_);
  xor g_099811_(out[243], out[947], _055087_);
  xor g_099812_(out[240], out[944], _055098_);
  or g_099813_(_054988_, _055065_, _055109_);
  or g_099814_(_055043_, _055109_, _055120_);
  or g_099815_(_054999_, _055087_, _055131_);
  or g_099816_(_055010_, _055131_, _055142_);
  or g_099817_(_055120_, _055142_, _055153_);
  or g_099818_(_054977_, _055076_, _055164_);
  or g_099819_(_055153_, _055164_, _055175_);
  or g_099820_(_054922_, _054933_, _055186_);
  xor g_099821_(out[247], out[951], _055197_);
  or g_099822_(_054955_, _055197_, _055208_);
  or g_099823_(_055186_, _055208_, _055219_);
  or g_099824_(_055021_, _055032_, _055230_);
  or g_099825_(_055054_, _055230_, _055241_);
  or g_099826_(_055219_, _055241_, _055252_);
  or g_099827_(_055098_, _055252_, _055263_);
  or g_099828_(_055175_, _055263_, _055274_);
  xor g_099829_(out[231], out[951], _055285_);
  and g_099830_(_098228_, out[955], _055296_);
  xor g_099831_(out[238], out[958], _055307_);
  xor g_099832_(out[232], out[952], _055318_);
  xor g_099833_(out[225], out[945], _055329_);
  xor g_099834_(out[237], out[957], _055340_);
  xor g_099835_(out[233], out[953], _055351_);
  xor g_099836_(out[228], out[948], _055362_);
  xor g_099837_(out[226], out[946], _055373_);
  and g_099838_(out[235], _049829_, _055384_);
  xor g_099839_(out[227], out[947], _055395_);
  xor g_099840_(out[230], out[950], _055406_);
  xor g_099841_(out[239], out[959], _055417_);
  xor g_099842_(out[234], out[954], _055428_);
  xor g_099843_(out[229], out[949], _055439_);
  xor g_099844_(out[224], out[944], _055450_);
  or g_099845_(_055307_, _055362_, _055461_);
  or g_099846_(_055318_, _055340_, _055472_);
  or g_099847_(_055373_, _055428_, _055483_);
  or g_099848_(_055472_, _055483_, _055494_);
  or g_099849_(_055351_, _055395_, _055505_);
  or g_099850_(_055439_, _055450_, _055516_);
  or g_099851_(_055505_, _055516_, _055527_);
  or g_099852_(_055494_, _055527_, _055538_);
  xor g_099853_(out[236], out[956], _055549_);
  or g_099854_(_055296_, _055549_, _055560_);
  or g_099855_(_055285_, _055406_, _055571_);
  or g_099856_(_055560_, _055571_, _055582_);
  or g_099857_(_055329_, _055384_, _055593_);
  or g_099858_(_055417_, _055593_, _055604_);
  or g_099859_(_055582_, _055604_, _055615_);
  or g_099860_(_055538_, _055615_, _055626_);
  or g_099861_(_055461_, _055626_, _055637_);
  xor g_099862_(out[209], out[945], _055648_);
  and g_099863_(out[219], _049829_, _055659_);
  xor g_099864_(out[222], out[958], _055670_);
  xor g_099865_(out[211], out[947], _055681_);
  xor g_099866_(out[212], out[948], _055692_);
  xor g_099867_(out[210], out[946], _055703_);
  xor g_099868_(out[217], out[953], _055714_);
  xor g_099869_(out[208], out[944], _055725_);
  and g_099870_(_098217_, out[955], _055736_);
  xor g_099871_(out[214], out[950], _055747_);
  xor g_099872_(out[218], out[954], _055758_);
  xor g_099873_(out[213], out[949], _055769_);
  xor g_099874_(out[223], out[959], _055780_);
  xor g_099875_(out[221], out[957], _055791_);
  xor g_099876_(out[216], out[952], _055802_);
  or g_099877_(_055670_, _055692_, _055813_);
  or g_099878_(_055791_, _055802_, _055824_);
  or g_099879_(_055703_, _055758_, _055835_);
  or g_099880_(_055824_, _055835_, _055846_);
  or g_099881_(_055681_, _055714_, _055857_);
  or g_099882_(_055725_, _055769_, _055868_);
  or g_099883_(_055857_, _055868_, _055879_);
  or g_099884_(_055846_, _055879_, _055890_);
  xor g_099885_(out[220], out[956], _055901_);
  or g_099886_(_055736_, _055901_, _055912_);
  xor g_099887_(out[215], out[951], _055923_);
  or g_099888_(_055747_, _055923_, _055934_);
  or g_099889_(_055912_, _055934_, _055945_);
  or g_099890_(_055648_, _055659_, _055956_);
  or g_099891_(_055780_, _055956_, _055967_);
  or g_099892_(_055945_, _055967_, _055978_);
  or g_099893_(_055890_, _055978_, _055989_);
  or g_099894_(_055813_, _055989_, _056000_);
  xor g_099895_(out[199], out[951], _056011_);
  and g_099896_(_098206_, out[955], _056022_);
  xor g_099897_(out[206], out[958], _056033_);
  xor g_099898_(out[200], out[952], _056044_);
  xor g_099899_(out[193], out[945], _056055_);
  xor g_099900_(out[205], out[957], _056066_);
  xor g_099901_(out[201], out[953], _056077_);
  xor g_099902_(out[196], out[948], _056088_);
  xor g_099903_(out[194], out[946], _056099_);
  and g_099904_(out[203], _049829_, _056110_);
  xor g_099905_(out[195], out[947], _056121_);
  xor g_099906_(out[198], out[950], _056132_);
  xor g_099907_(out[207], out[959], _056143_);
  xor g_099908_(out[202], out[954], _056154_);
  xor g_099909_(out[197], out[949], _056165_);
  xor g_099910_(out[192], out[944], _056176_);
  or g_099911_(_056033_, _056088_, _056187_);
  or g_099912_(_056044_, _056066_, _056198_);
  or g_099913_(_056099_, _056154_, _056209_);
  or g_099914_(_056198_, _056209_, _056220_);
  or g_099915_(_056077_, _056121_, _056231_);
  or g_099916_(_056165_, _056176_, _056242_);
  or g_099917_(_056231_, _056242_, _056253_);
  or g_099918_(_056220_, _056253_, _056264_);
  xor g_099919_(out[204], out[956], _056275_);
  or g_099920_(_056022_, _056275_, _056286_);
  or g_099921_(_056011_, _056132_, _056297_);
  or g_099922_(_056286_, _056297_, _056308_);
  or g_099923_(_056055_, _056110_, _056319_);
  or g_099924_(_056143_, _056319_, _056330_);
  or g_099925_(_056308_, _056330_, _056341_);
  or g_099926_(_056264_, _056341_, _056352_);
  or g_099927_(_056187_, _056352_, _056363_);
  xor g_099928_(out[189], out[957], _056374_);
  xor g_099929_(out[178], out[946], _056385_);
  xor g_099930_(out[181], out[949], _056396_);
  xor g_099931_(out[185], out[953], _056407_);
  xor g_099932_(out[180], out[948], _056418_);
  xor g_099933_(out[184], out[952], _056429_);
  xor g_099934_(out[190], out[958], _056440_);
  xor g_099935_(out[182], out[950], _056451_);
  xor g_099936_(out[191], out[959], _056462_);
  xor g_099937_(out[186], out[954], _056473_);
  xor g_099938_(out[176], out[944], _056484_);
  xor g_099939_(out[179], out[947], _056495_);
  and g_099940_(_098195_, out[955], _056506_);
  and g_099941_(out[187], _049829_, _056517_);
  xor g_099942_(out[177], out[945], _056528_);
  or g_099943_(_056418_, _056440_, _056539_);
  or g_099944_(_056374_, _056429_, _056550_);
  or g_099945_(_056385_, _056473_, _056561_);
  or g_099946_(_056550_, _056561_, _056572_);
  or g_099947_(_056407_, _056495_, _056583_);
  or g_099948_(_056396_, _056484_, _056594_);
  or g_099949_(_056583_, _056594_, _056605_);
  or g_099950_(_056572_, _056605_, _056616_);
  xor g_099951_(out[188], out[956], _056627_);
  or g_099952_(_056506_, _056627_, _056638_);
  xor g_099953_(out[183], out[951], _056649_);
  or g_099954_(_056451_, _056649_, _056660_);
  or g_099955_(_056638_, _056660_, _056671_);
  or g_099956_(_056517_, _056528_, _056682_);
  or g_099957_(_056462_, _056682_, _056693_);
  or g_099958_(_056671_, _056693_, _056704_);
  or g_099959_(_056616_, _056704_, _056715_);
  or g_099960_(_056539_, _056715_, _056726_);
  xor g_099961_(out[167], out[951], _056737_);
  and g_099962_(_098184_, out[955], _056748_);
  xor g_099963_(out[174], out[958], _056759_);
  xor g_099964_(out[168], out[952], _056770_);
  xor g_099965_(out[161], out[945], _056781_);
  xor g_099966_(out[173], out[957], _056792_);
  xor g_099967_(out[169], out[953], _056803_);
  xor g_099968_(out[164], out[948], _056814_);
  xor g_099969_(out[162], out[946], _056825_);
  and g_099970_(out[171], _049829_, _056836_);
  xor g_099971_(out[163], out[947], _056847_);
  xor g_099972_(out[166], out[950], _056858_);
  xor g_099973_(out[175], out[959], _056869_);
  xor g_099974_(out[170], out[954], _056880_);
  xor g_099975_(out[165], out[949], _056891_);
  xor g_099976_(out[160], out[944], _056902_);
  or g_099977_(_056759_, _056814_, _056913_);
  or g_099978_(_056770_, _056792_, _056924_);
  or g_099979_(_056825_, _056880_, _056935_);
  or g_099980_(_056924_, _056935_, _056946_);
  or g_099981_(_056803_, _056847_, _056957_);
  or g_099982_(_056891_, _056902_, _056968_);
  or g_099983_(_056957_, _056968_, _056979_);
  or g_099984_(_056946_, _056979_, _056990_);
  xor g_099985_(out[172], out[956], _057001_);
  or g_099986_(_056748_, _057001_, _057012_);
  or g_099987_(_056737_, _056858_, _057023_);
  or g_099988_(_057012_, _057023_, _057034_);
  or g_099989_(_056781_, _056836_, _057045_);
  or g_099990_(_056869_, _057045_, _057056_);
  or g_099991_(_057034_, _057056_, _057067_);
  or g_099992_(_056990_, _057067_, _057078_);
  or g_099993_(_056913_, _057078_, _057089_);
  xor g_099994_(out[145], out[945], _057100_);
  and g_099995_(out[155], _049829_, _057111_);
  xor g_099996_(out[153], out[953], _057122_);
  xor g_099997_(out[144], out[944], _057133_);
  xor g_099998_(out[158], out[958], _057144_);
  xor g_099999_(out[148], out[948], _057155_);
  or g_100000_(_057144_, _057155_, _057166_);
  xor g_100001_(out[157], out[957], _057177_);
  xor g_100002_(out[147], out[947], _057188_);
  and g_100003_(_098173_, out[955], _057199_);
  xor g_100004_(out[150], out[950], _057210_);
  xor g_100005_(out[154], out[954], _057221_);
  xor g_100006_(out[149], out[949], _057232_);
  xor g_100007_(out[159], out[959], _057243_);
  xor g_100008_(out[152], out[952], _057254_);
  or g_100009_(_057177_, _057254_, _057265_);
  xor g_100010_(out[146], out[946], _057276_);
  or g_100011_(_057221_, _057276_, _057287_);
  or g_100012_(_057265_, _057287_, _057298_);
  or g_100013_(_057122_, _057188_, _057309_);
  or g_100014_(_057232_, _057309_, _057320_);
  or g_100015_(_057298_, _057320_, _057331_);
  or g_100016_(_057166_, _057331_, _057342_);
  xor g_100017_(out[156], out[956], _057353_);
  or g_100018_(_057199_, _057353_, _057364_);
  xor g_100019_(out[151], out[951], _057375_);
  or g_100020_(_057210_, _057375_, _057386_);
  or g_100021_(_057364_, _057386_, _057397_);
  or g_100022_(_057100_, _057111_, _057408_);
  or g_100023_(_057243_, _057408_, _057419_);
  or g_100024_(_057397_, _057419_, _057430_);
  or g_100025_(_057133_, _057430_, _057441_);
  or g_100026_(_057342_, _057441_, _057452_);
  xor g_100027_(out[135], out[951], _057463_);
  and g_100028_(_098162_, out[955], _057474_);
  xor g_100029_(out[142], out[958], _057485_);
  xor g_100030_(out[136], out[952], _057496_);
  xor g_100031_(out[129], out[945], _057507_);
  xor g_100032_(out[141], out[957], _057518_);
  xor g_100033_(out[137], out[953], _057529_);
  xor g_100034_(out[132], out[948], _057540_);
  xor g_100035_(out[130], out[946], _057551_);
  and g_100036_(out[139], _049829_, _057562_);
  xor g_100037_(out[131], out[947], _057573_);
  xor g_100038_(out[134], out[950], _057584_);
  xor g_100039_(out[143], out[959], _057595_);
  xor g_100040_(out[138], out[954], _057606_);
  xor g_100041_(out[133], out[949], _057617_);
  xor g_100042_(out[128], out[944], _057628_);
  or g_100043_(_057485_, _057540_, _057639_);
  or g_100044_(_057496_, _057518_, _057650_);
  or g_100045_(_057551_, _057606_, _057661_);
  or g_100046_(_057650_, _057661_, _057672_);
  or g_100047_(_057529_, _057573_, _057683_);
  or g_100048_(_057617_, _057628_, _057694_);
  or g_100049_(_057683_, _057694_, _057705_);
  or g_100050_(_057672_, _057705_, _057716_);
  xor g_100051_(out[140], out[956], _057727_);
  or g_100052_(_057474_, _057727_, _057738_);
  or g_100053_(_057463_, _057584_, _057749_);
  or g_100054_(_057738_, _057749_, _057760_);
  or g_100055_(_057507_, _057562_, _057771_);
  or g_100056_(_057595_, _057771_, _057782_);
  or g_100057_(_057760_, _057782_, _057793_);
  or g_100058_(_057716_, _057793_, _057804_);
  or g_100059_(_057639_, _057804_, _057815_);
  xor g_100060_(out[113], out[945], _057826_);
  and g_100061_(out[123], _049829_, _057837_);
  xor g_100062_(out[121], out[953], _057848_);
  xor g_100063_(out[112], out[944], _057859_);
  xor g_100064_(out[126], out[958], _057870_);
  xor g_100065_(out[116], out[948], _057881_);
  or g_100066_(_057870_, _057881_, _057892_);
  xor g_100067_(out[125], out[957], _057903_);
  xor g_100068_(out[115], out[947], _057914_);
  and g_100069_(_098151_, out[955], _057925_);
  xor g_100070_(out[118], out[950], _057936_);
  xor g_100071_(out[122], out[954], _057947_);
  xor g_100072_(out[117], out[949], _057958_);
  xor g_100073_(out[127], out[959], _057969_);
  xor g_100074_(out[120], out[952], _057980_);
  or g_100075_(_057903_, _057980_, _057991_);
  xor g_100076_(out[114], out[946], _058002_);
  or g_100077_(_057947_, _058002_, _058013_);
  or g_100078_(_057991_, _058013_, _058024_);
  or g_100079_(_057848_, _057914_, _058035_);
  or g_100080_(_057958_, _058035_, _058046_);
  or g_100081_(_058024_, _058046_, _058057_);
  or g_100082_(_057892_, _058057_, _058068_);
  xor g_100083_(out[124], out[956], _058079_);
  or g_100084_(_057925_, _058079_, _058090_);
  xor g_100085_(out[119], out[951], _058101_);
  or g_100086_(_057936_, _058101_, _058112_);
  or g_100087_(_058090_, _058112_, _058123_);
  or g_100088_(_057826_, _057837_, _058134_);
  or g_100089_(_057969_, _058134_, _058145_);
  or g_100090_(_058123_, _058145_, _058156_);
  or g_100091_(_057859_, _058156_, _058167_);
  or g_100092_(_058068_, _058167_, _058178_);
  xor g_100093_(out[103], out[951], _058189_);
  and g_100094_(_098140_, out[955], _058200_);
  xor g_100095_(out[110], out[958], _058211_);
  xor g_100096_(out[104], out[952], _058222_);
  xor g_100097_(out[97], out[945], _058233_);
  xor g_100098_(out[109], out[957], _058244_);
  xor g_100099_(out[105], out[953], _058255_);
  xor g_100100_(out[100], out[948], _058266_);
  xor g_100101_(out[98], out[946], _058277_);
  and g_100102_(out[107], _049829_, _058288_);
  xor g_100103_(out[99], out[947], _058299_);
  xor g_100104_(out[102], out[950], _058310_);
  xor g_100105_(out[111], out[959], _058321_);
  xor g_100106_(out[106], out[954], _058332_);
  xor g_100107_(out[101], out[949], _058343_);
  xor g_100108_(out[96], out[944], _058354_);
  or g_100109_(_058211_, _058266_, _058365_);
  or g_100110_(_058222_, _058244_, _058376_);
  or g_100111_(_058277_, _058332_, _058387_);
  or g_100112_(_058376_, _058387_, _058398_);
  or g_100113_(_058255_, _058299_, _058409_);
  or g_100114_(_058343_, _058354_, _058420_);
  or g_100115_(_058409_, _058420_, _058431_);
  or g_100116_(_058398_, _058431_, _058442_);
  xor g_100117_(out[108], out[956], _058453_);
  or g_100118_(_058200_, _058453_, _058464_);
  or g_100119_(_058189_, _058310_, _058475_);
  or g_100120_(_058464_, _058475_, _058486_);
  or g_100121_(_058233_, _058288_, _058497_);
  or g_100122_(_058321_, _058497_, _058508_);
  or g_100123_(_058486_, _058508_, _058519_);
  or g_100124_(_058442_, _058519_, _058530_);
  or g_100125_(_058365_, _058530_, _058541_);
  xor g_100126_(out[90], out[954], _058552_);
  xor g_100127_(out[82], out[946], _058563_);
  xor g_100128_(out[81], out[945], _058574_);
  and g_100129_(_098129_, out[955], _058585_);
  and g_100130_(out[91], _049829_, _058596_);
  xor g_100131_(out[93], out[957], _058607_);
  xor g_100132_(out[83], out[947], _058618_);
  xor g_100133_(out[94], out[958], _058629_);
  xor g_100134_(out[92], out[956], _058640_);
  xor g_100135_(out[88], out[952], _058651_);
  xor g_100136_(out[95], out[959], _058662_);
  xor g_100137_(out[85], out[949], _058673_);
  xor g_100138_(out[86], out[950], _058684_);
  xor g_100139_(out[80], out[944], _058695_);
  xor g_100140_(out[84], out[948], _058706_);
  or g_100141_(_058607_, _058651_, _058717_);
  xor g_100142_(out[89], out[953], _058728_);
  or g_100143_(_058552_, _058563_, _058739_);
  or g_100144_(_058717_, _058739_, _058750_);
  or g_100145_(_058618_, _058728_, _058761_);
  or g_100146_(_058673_, _058761_, _058772_);
  or g_100147_(_058750_, _058772_, _058783_);
  or g_100148_(_058629_, _058706_, _058794_);
  or g_100149_(_058783_, _058794_, _058805_);
  or g_100150_(_058585_, _058640_, _058816_);
  xor g_100151_(out[87], out[951], _058827_);
  or g_100152_(_058684_, _058827_, _058838_);
  or g_100153_(_058816_, _058838_, _058849_);
  or g_100154_(_058574_, _058596_, _058860_);
  or g_100155_(_058662_, _058860_, _058871_);
  or g_100156_(_058849_, _058871_, _058882_);
  or g_100157_(_058695_, _058882_, _058893_);
  or g_100158_(_058805_, _058893_, _058904_);
  xor g_100159_(out[71], out[951], _058915_);
  and g_100160_(_098118_, out[955], _058926_);
  xor g_100161_(out[78], out[958], _058937_);
  xor g_100162_(out[72], out[952], _058948_);
  xor g_100163_(out[65], out[945], _058959_);
  xor g_100164_(out[77], out[957], _058970_);
  xor g_100165_(out[73], out[953], _058981_);
  xor g_100166_(out[68], out[948], _058992_);
  xor g_100167_(out[66], out[946], _059003_);
  and g_100168_(out[75], _049829_, _059014_);
  xor g_100169_(out[67], out[947], _059025_);
  xor g_100170_(out[70], out[950], _059036_);
  xor g_100171_(out[79], out[959], _059047_);
  xor g_100172_(out[74], out[954], _059058_);
  xor g_100173_(out[69], out[949], _059069_);
  xor g_100174_(out[64], out[944], _059080_);
  or g_100175_(_058937_, _058992_, _059091_);
  or g_100176_(_058948_, _058970_, _059102_);
  or g_100177_(_059003_, _059058_, _059113_);
  or g_100178_(_059102_, _059113_, _059124_);
  or g_100179_(_058981_, _059025_, _059135_);
  or g_100180_(_059069_, _059080_, _059146_);
  or g_100181_(_059135_, _059146_, _059157_);
  or g_100182_(_059124_, _059157_, _059168_);
  xor g_100183_(out[76], out[956], _059179_);
  or g_100184_(_058926_, _059179_, _059190_);
  or g_100185_(_058915_, _059036_, _059201_);
  or g_100186_(_059190_, _059201_, _059212_);
  or g_100187_(_058959_, _059014_, _059223_);
  or g_100188_(_059047_, _059223_, _059234_);
  or g_100189_(_059212_, _059234_, _059245_);
  or g_100190_(_059168_, _059245_, _059256_);
  or g_100191_(_059091_, _059256_, _059267_);
  xor g_100192_(out[60], out[956], _059278_);
  and g_100193_(_098107_, out[955], _059289_);
  xor g_100194_(out[56], out[952], _059300_);
  xor g_100195_(out[54], out[950], _059311_);
  xor g_100196_(out[61], out[957], _059322_);
  xor g_100197_(out[62], out[958], _059333_);
  xor g_100198_(out[50], out[946], _059344_);
  xor g_100199_(out[57], out[953], _059355_);
  xor g_100200_(out[53], out[949], _059366_);
  xor g_100201_(out[49], out[945], _059377_);
  and g_100202_(out[59], _049829_, _059388_);
  or g_100203_(_059300_, _059322_, _059399_);
  xor g_100204_(out[63], out[959], _059410_);
  xor g_100205_(out[58], out[954], _059421_);
  xor g_100206_(out[52], out[948], _059432_);
  xor g_100207_(out[51], out[947], _059443_);
  xor g_100208_(out[48], out[944], _059454_);
  or g_100209_(_059344_, _059421_, _059465_);
  or g_100210_(_059399_, _059465_, _059476_);
  or g_100211_(_059355_, _059443_, _059487_);
  or g_100212_(_059366_, _059487_, _059498_);
  or g_100213_(_059476_, _059498_, _059509_);
  or g_100214_(_059333_, _059432_, _059520_);
  or g_100215_(_059509_, _059520_, _059531_);
  or g_100216_(_059278_, _059289_, _059542_);
  xor g_100217_(out[55], out[951], _059553_);
  or g_100218_(_059311_, _059553_, _059564_);
  or g_100219_(_059542_, _059564_, _059575_);
  or g_100220_(_059377_, _059388_, _059586_);
  or g_100221_(_059410_, _059586_, _059597_);
  or g_100222_(_059575_, _059597_, _059608_);
  or g_100223_(_059454_, _059608_, _059619_);
  or g_100224_(_059531_, _059619_, _059630_);
  xor g_100225_(out[39], out[951], _059641_);
  and g_100226_(_098096_, out[955], _059652_);
  xor g_100227_(out[46], out[958], _059663_);
  xor g_100228_(out[40], out[952], _059674_);
  xor g_100229_(out[33], out[945], _059685_);
  xor g_100230_(out[45], out[957], _059696_);
  xor g_100231_(out[41], out[953], _059707_);
  xor g_100232_(out[36], out[948], _059718_);
  xor g_100233_(out[34], out[946], _059729_);
  and g_100234_(out[43], _049829_, _059740_);
  xor g_100235_(out[35], out[947], _059751_);
  xor g_100236_(out[38], out[950], _059762_);
  xor g_100237_(out[47], out[959], _059773_);
  xor g_100238_(out[42], out[954], _059784_);
  xor g_100239_(out[37], out[949], _059795_);
  xor g_100240_(out[32], out[944], _059806_);
  or g_100241_(_059663_, _059718_, _059817_);
  or g_100242_(_059674_, _059696_, _059828_);
  or g_100243_(_059729_, _059784_, _059839_);
  or g_100244_(_059828_, _059839_, _059850_);
  or g_100245_(_059707_, _059751_, _059861_);
  or g_100246_(_059795_, _059806_, _059872_);
  or g_100247_(_059861_, _059872_, _059883_);
  or g_100248_(_059850_, _059883_, _059894_);
  xor g_100249_(out[44], out[956], _059905_);
  or g_100250_(_059652_, _059905_, _059916_);
  or g_100251_(_059641_, _059762_, _059927_);
  or g_100252_(_059916_, _059927_, _059938_);
  or g_100253_(_059685_, _059740_, _059949_);
  or g_100254_(_059773_, _059949_, _059960_);
  or g_100255_(_059938_, _059960_, _059971_);
  or g_100256_(_059894_, _059971_, _059982_);
  or g_100257_(_059817_, _059982_, _059993_);
  xor g_100258_(out[17], out[945], _060004_);
  and g_100259_(out[27], _049829_, _060015_);
  xor g_100260_(out[25], out[953], _060026_);
  xor g_100261_(out[16], out[944], _060037_);
  xor g_100262_(out[30], out[958], _060048_);
  xor g_100263_(out[20], out[948], _060059_);
  or g_100264_(_060048_, _060059_, _060070_);
  xor g_100265_(out[29], out[957], _060081_);
  xor g_100266_(out[19], out[947], _060092_);
  and g_100267_(_098063_, out[955], _060103_);
  xor g_100268_(out[22], out[950], _060114_);
  xor g_100269_(out[26], out[954], _060125_);
  xor g_100270_(out[21], out[949], _060136_);
  xor g_100271_(out[31], out[959], _060147_);
  xor g_100272_(out[24], out[952], _060158_);
  or g_100273_(_060081_, _060158_, _060169_);
  xor g_100274_(out[18], out[946], _060180_);
  or g_100275_(_060125_, _060180_, _060191_);
  or g_100276_(_060169_, _060191_, _060202_);
  or g_100277_(_060026_, _060092_, _060213_);
  or g_100278_(_060136_, _060213_, _060224_);
  or g_100279_(_060202_, _060224_, _060235_);
  or g_100280_(_060070_, _060235_, _060246_);
  xor g_100281_(out[28], out[956], _060257_);
  or g_100282_(_060103_, _060257_, _060268_);
  xor g_100283_(out[23], out[951], _060279_);
  or g_100284_(_060114_, _060279_, _060290_);
  or g_100285_(_060268_, _060290_, _060301_);
  or g_100286_(_060004_, _060015_, _060312_);
  or g_100287_(_060147_, _060312_, _060323_);
  or g_100288_(_060301_, _060323_, _060334_);
  or g_100289_(_060037_, _060334_, _060345_);
  or g_100290_(_060246_, _060345_, _060356_);
  xor g_100291_(out[1], out[945], _060367_);
  and g_100292_(_098041_, out[955], _060378_);
  and g_100293_(out[11], _049829_, _060389_);
  xor g_100294_(out[8], out[952], _060400_);
  xor g_100295_(out[10], out[954], _060411_);
  xor g_100296_(out[2], out[946], _060422_);
  xor g_100297_(out[4], out[948], _060433_);
  xor g_100298_(out[5], out[949], _060444_);
  xor g_100299_(out[9], out[953], _060455_);
  xor g_100300_(out[3], out[947], _060466_);
  xor g_100301_(out[14], out[958], _060477_);
  xor g_100302_(out[0], out[944], _060488_);
  xor g_100303_(out[15], out[959], _060499_);
  xor g_100304_(out[13], out[957], _060510_);
  or g_100305_(_060400_, _060510_, _060521_);
  xor g_100306_(out[6], out[950], _060532_);
  or g_100307_(_060411_, _060422_, _060543_);
  or g_100308_(_060521_, _060543_, _060554_);
  or g_100309_(_060455_, _060466_, _060565_);
  or g_100310_(_060444_, _060565_, _060576_);
  or g_100311_(_060554_, _060576_, _060587_);
  or g_100312_(_060433_, _060477_, _060598_);
  or g_100313_(_060587_, _060598_, _060609_);
  xor g_100314_(out[12], out[956], _060620_);
  or g_100315_(_060378_, _060620_, _060631_);
  xor g_100316_(out[7], out[951], _060642_);
  or g_100317_(_060532_, _060642_, _060653_);
  or g_100318_(_060631_, _060653_, _060664_);
  or g_100319_(_060367_, _060389_, _060675_);
  or g_100320_(_060499_, _060675_, _060686_);
  or g_100321_(_060664_, _060686_, _060697_);
  or g_100322_(_060488_, _060697_, _060708_);
  or g_100323_(_060609_, _060708_, _060719_);
  xor g_100324_(out[471], out[935], _060730_);
  and g_100325_(_049499_, out[939], _060741_);
  xor g_100326_(out[478], out[942], _060752_);
  xor g_100327_(out[472], out[936], _060763_);
  xor g_100328_(out[465], out[929], _060774_);
  xor g_100329_(out[477], out[941], _060785_);
  xor g_100330_(out[473], out[937], _060796_);
  xor g_100331_(out[468], out[932], _060807_);
  xor g_100332_(out[466], out[930], _060818_);
  and g_100333_(out[475], _049807_, _060829_);
  xor g_100334_(out[467], out[931], _060840_);
  xor g_100335_(out[470], out[934], _060851_);
  xor g_100336_(out[479], out[943], _060862_);
  xor g_100337_(out[474], out[938], _060873_);
  xor g_100338_(out[469], out[933], _060884_);
  xor g_100339_(out[464], out[928], _060895_);
  or g_100340_(_060752_, _060807_, _060906_);
  or g_100341_(_060763_, _060785_, _060917_);
  or g_100342_(_060818_, _060873_, _060928_);
  or g_100343_(_060917_, _060928_, _060939_);
  or g_100344_(_060796_, _060840_, _060950_);
  or g_100345_(_060884_, _060895_, _060961_);
  or g_100346_(_060950_, _060961_, _060972_);
  or g_100347_(_060939_, _060972_, _060983_);
  xor g_100348_(out[476], out[940], _060994_);
  or g_100349_(_060741_, _060994_, _061005_);
  or g_100350_(_060730_, _060851_, _061016_);
  or g_100351_(_061005_, _061016_, _061027_);
  or g_100352_(_060774_, _060829_, _061038_);
  or g_100353_(_060862_, _061038_, _061049_);
  or g_100354_(_061027_, _061049_, _061060_);
  or g_100355_(_060983_, _061060_, _061071_);
  or g_100356_(_060906_, _061071_, _061082_);
  xor g_100357_(out[449], out[929], _061093_);
  and g_100358_(out[459], _049807_, _061104_);
  xor g_100359_(out[457], out[937], _061115_);
  xor g_100360_(out[448], out[928], _061126_);
  xor g_100361_(out[462], out[942], _061137_);
  xor g_100362_(out[452], out[932], _061148_);
  or g_100363_(_061137_, _061148_, _061159_);
  xor g_100364_(out[461], out[941], _061170_);
  xor g_100365_(out[451], out[931], _061181_);
  and g_100366_(_049477_, out[939], _061192_);
  xor g_100367_(out[454], out[934], _061203_);
  xor g_100368_(out[458], out[938], _061214_);
  xor g_100369_(out[453], out[933], _061225_);
  xor g_100370_(out[463], out[943], _061236_);
  xor g_100371_(out[456], out[936], _061247_);
  or g_100372_(_061170_, _061247_, _061258_);
  xor g_100373_(out[450], out[930], _061269_);
  or g_100374_(_061214_, _061269_, _061280_);
  or g_100375_(_061258_, _061280_, _061291_);
  or g_100376_(_061115_, _061181_, _061302_);
  or g_100377_(_061225_, _061302_, _061313_);
  or g_100378_(_061291_, _061313_, _061324_);
  or g_100379_(_061159_, _061324_, _061335_);
  xor g_100380_(out[460], out[940], _061346_);
  or g_100381_(_061192_, _061346_, _061357_);
  xor g_100382_(out[455], out[935], _061368_);
  or g_100383_(_061203_, _061368_, _061379_);
  or g_100384_(_061357_, _061379_, _061390_);
  or g_100385_(_061093_, _061104_, _061401_);
  or g_100386_(_061236_, _061401_, _061412_);
  or g_100387_(_061390_, _061412_, _061423_);
  or g_100388_(_061126_, _061423_, _061434_);
  or g_100389_(_061335_, _061434_, _061445_);
  xor g_100390_(out[439], out[935], _061456_);
  and g_100391_(_049466_, out[939], _061467_);
  xor g_100392_(out[446], out[942], _061478_);
  xor g_100393_(out[440], out[936], _061489_);
  xor g_100394_(out[433], out[929], _061500_);
  xor g_100395_(out[445], out[941], _061511_);
  xor g_100396_(out[441], out[937], _061522_);
  xor g_100397_(out[436], out[932], _061533_);
  xor g_100398_(out[434], out[930], _061544_);
  and g_100399_(out[443], _049807_, _061555_);
  xor g_100400_(out[435], out[931], _061566_);
  xor g_100401_(out[438], out[934], _061577_);
  xor g_100402_(out[447], out[943], _061588_);
  xor g_100403_(out[442], out[938], _061599_);
  xor g_100404_(out[437], out[933], _061610_);
  xor g_100405_(out[432], out[928], _061621_);
  or g_100406_(_061478_, _061533_, _061632_);
  or g_100407_(_061489_, _061511_, _061643_);
  or g_100408_(_061544_, _061599_, _061654_);
  or g_100409_(_061643_, _061654_, _061665_);
  or g_100410_(_061522_, _061566_, _061676_);
  or g_100411_(_061610_, _061621_, _061687_);
  or g_100412_(_061676_, _061687_, _061698_);
  or g_100413_(_061665_, _061698_, _061709_);
  xor g_100414_(out[444], out[940], _061720_);
  or g_100415_(_061467_, _061720_, _061731_);
  or g_100416_(_061456_, _061577_, _061742_);
  or g_100417_(_061731_, _061742_, _061753_);
  or g_100418_(_061500_, _061555_, _061764_);
  or g_100419_(_061588_, _061764_, _061775_);
  or g_100420_(_061753_, _061775_, _061786_);
  or g_100421_(_061709_, _061786_, _061797_);
  or g_100422_(_061632_, _061797_, _061808_);
  not g_100423_(_061808_, _061819_);
  xor g_100424_(out[424], out[936], _061830_);
  xor g_100425_(out[421], out[933], _061841_);
  xor g_100426_(out[419], out[931], _061852_);
  xor g_100427_(out[430], out[942], _061863_);
  xor g_100428_(out[429], out[941], _061874_);
  xor g_100429_(out[418], out[930], _061885_);
  xor g_100430_(out[425], out[937], _061896_);
  xor g_100431_(out[422], out[934], _061907_);
  xor g_100432_(out[431], out[943], _061918_);
  xor g_100433_(out[426], out[938], _061929_);
  xor g_100434_(out[420], out[932], _061940_);
  xor g_100435_(out[416], out[928], _061951_);
  and g_100436_(_049455_, out[939], _061962_);
  and g_100437_(out[427], _049807_, _061973_);
  or g_100438_(_061830_, _061874_, _061984_);
  xor g_100439_(out[417], out[929], _061995_);
  or g_100440_(_061885_, _061929_, _062006_);
  or g_100441_(_061984_, _062006_, _062017_);
  or g_100442_(_061852_, _061896_, _062028_);
  or g_100443_(_061841_, _062028_, _062039_);
  or g_100444_(_062017_, _062039_, _062050_);
  or g_100445_(_061863_, _061940_, _062061_);
  or g_100446_(_062050_, _062061_, _062072_);
  xor g_100447_(out[428], out[940], _062083_);
  or g_100448_(_061962_, _062083_, _062094_);
  xor g_100449_(out[423], out[935], _062105_);
  or g_100450_(_061907_, _062105_, _062116_);
  or g_100451_(_062094_, _062116_, _062127_);
  or g_100452_(_061973_, _061995_, _062138_);
  or g_100453_(_061918_, _062138_, _062149_);
  or g_100454_(_062127_, _062149_, _062160_);
  or g_100455_(_061951_, _062160_, _062171_);
  or g_100456_(_062072_, _062171_, _062182_);
  xor g_100457_(out[407], out[935], _062193_);
  and g_100458_(_049444_, out[939], _062204_);
  xor g_100459_(out[414], out[942], _062215_);
  xor g_100460_(out[408], out[936], _062226_);
  xor g_100461_(out[401], out[929], _062237_);
  xor g_100462_(out[413], out[941], _062248_);
  xor g_100463_(out[409], out[937], _062259_);
  xor g_100464_(out[404], out[932], _062270_);
  xor g_100465_(out[402], out[930], _062281_);
  and g_100466_(out[411], _049807_, _062292_);
  xor g_100467_(out[403], out[931], _062303_);
  xor g_100468_(out[406], out[934], _062314_);
  xor g_100469_(out[415], out[943], _062325_);
  xor g_100470_(out[410], out[938], _062336_);
  xor g_100471_(out[405], out[933], _062347_);
  xor g_100472_(out[400], out[928], _062358_);
  or g_100473_(_062215_, _062270_, _062369_);
  or g_100474_(_062226_, _062248_, _062380_);
  or g_100475_(_062281_, _062336_, _062391_);
  or g_100476_(_062380_, _062391_, _062402_);
  or g_100477_(_062259_, _062303_, _062413_);
  or g_100478_(_062347_, _062358_, _062424_);
  or g_100479_(_062413_, _062424_, _062435_);
  or g_100480_(_062402_, _062435_, _062446_);
  xor g_100481_(out[412], out[940], _062457_);
  or g_100482_(_062204_, _062457_, _062468_);
  or g_100483_(_062193_, _062314_, _062479_);
  or g_100484_(_062468_, _062479_, _062490_);
  or g_100485_(_062237_, _062292_, _062501_);
  or g_100486_(_062325_, _062501_, _062512_);
  or g_100487_(_062490_, _062512_, _062523_);
  or g_100488_(_062446_, _062523_, _062534_);
  or g_100489_(_062369_, _062534_, _062545_);
  xor g_100490_(out[388], out[932], _062556_);
  xor g_100491_(out[396], out[940], _062567_);
  and g_100492_(_049433_, out[939], _062578_);
  xor g_100493_(out[394], out[938], _062589_);
  xor g_100494_(out[390], out[934], _062600_);
  xor g_100495_(out[389], out[933], _062611_);
  xor g_100496_(out[387], out[931], _062622_);
  xor g_100497_(out[397], out[941], _062633_);
  xor g_100498_(out[398], out[942], _062644_);
  xor g_100499_(out[385], out[929], _062655_);
  xor g_100500_(out[386], out[930], _062666_);
  and g_100501_(out[395], _049807_, _062677_);
  xor g_100502_(out[384], out[928], _062688_);
  xor g_100503_(out[399], out[943], _062699_);
  xor g_100504_(out[392], out[936], _062710_);
  or g_100505_(_062633_, _062710_, _062721_);
  xor g_100506_(out[393], out[937], _062732_);
  or g_100507_(_062589_, _062666_, _062743_);
  or g_100508_(_062721_, _062743_, _062754_);
  or g_100509_(_062622_, _062732_, _062765_);
  or g_100510_(_062611_, _062765_, _062776_);
  or g_100511_(_062754_, _062776_, _062787_);
  or g_100512_(_062556_, _062644_, _062798_);
  or g_100513_(_062787_, _062798_, _062809_);
  or g_100514_(_062567_, _062578_, _062820_);
  xor g_100515_(out[391], out[935], _062831_);
  or g_100516_(_062600_, _062831_, _062842_);
  or g_100517_(_062820_, _062842_, _062853_);
  or g_100518_(_062655_, _062677_, _062864_);
  or g_100519_(_062699_, _062864_, _062875_);
  or g_100520_(_062853_, _062875_, _062886_);
  or g_100521_(_062688_, _062886_, _062897_);
  or g_100522_(_062809_, _062897_, _062908_);
  not g_100523_(_062908_, _062919_);
  xor g_100524_(out[375], out[935], _062930_);
  and g_100525_(_049422_, out[939], _062941_);
  xor g_100526_(out[382], out[942], _062952_);
  xor g_100527_(out[376], out[936], _062963_);
  xor g_100528_(out[369], out[929], _062974_);
  xor g_100529_(out[381], out[941], _062985_);
  xor g_100530_(out[377], out[937], _062996_);
  xor g_100531_(out[372], out[932], _063007_);
  xor g_100532_(out[370], out[930], _063018_);
  and g_100533_(out[379], _049807_, _063029_);
  xor g_100534_(out[371], out[931], _063040_);
  xor g_100535_(out[374], out[934], _063051_);
  xor g_100536_(out[383], out[943], _063062_);
  xor g_100537_(out[378], out[938], _063073_);
  xor g_100538_(out[373], out[933], _063084_);
  xor g_100539_(out[368], out[928], _063095_);
  or g_100540_(_062952_, _063007_, _063106_);
  or g_100541_(_062963_, _062985_, _063117_);
  or g_100542_(_063018_, _063073_, _063128_);
  or g_100543_(_063117_, _063128_, _063139_);
  or g_100544_(_062996_, _063040_, _063150_);
  or g_100545_(_063084_, _063095_, _063161_);
  or g_100546_(_063150_, _063161_, _063172_);
  or g_100547_(_063139_, _063172_, _063183_);
  xor g_100548_(out[380], out[940], _063194_);
  or g_100549_(_062941_, _063194_, _063205_);
  or g_100550_(_062930_, _063051_, _063216_);
  or g_100551_(_063205_, _063216_, _063227_);
  or g_100552_(_062974_, _063029_, _063238_);
  or g_100553_(_063062_, _063238_, _063249_);
  or g_100554_(_063227_, _063249_, _063260_);
  or g_100555_(_063183_, _063260_, _063271_);
  or g_100556_(_063106_, _063271_, _063282_);
  not g_100557_(_063282_, _063293_);
  and g_100558_(out[363], _049807_, _063304_);
  xor g_100559_(out[356], out[932], _063315_);
  xor g_100560_(out[366], out[942], _063326_);
  or g_100561_(_063315_, _063326_, _063337_);
  xor g_100562_(out[365], out[941], _063348_);
  xor g_100563_(out[355], out[931], _063359_);
  xor g_100564_(out[352], out[928], _063370_);
  and g_100565_(_049411_, out[939], _063381_);
  xor g_100566_(out[362], out[938], _063392_);
  xor g_100567_(out[367], out[943], _063403_);
  xor g_100568_(out[358], out[934], _063414_);
  xor g_100569_(out[357], out[933], _063425_);
  xor g_100570_(out[360], out[936], _063436_);
  or g_100571_(_063348_, _063436_, _063447_);
  xor g_100572_(out[354], out[930], _063458_);
  xor g_100573_(out[361], out[937], _063469_);
  xor g_100574_(out[353], out[929], _063480_);
  or g_100575_(_063392_, _063458_, _063491_);
  or g_100576_(_063447_, _063491_, _063502_);
  or g_100577_(_063359_, _063469_, _063513_);
  or g_100578_(_063425_, _063513_, _063524_);
  or g_100579_(_063502_, _063524_, _063535_);
  or g_100580_(_063337_, _063535_, _063546_);
  xor g_100581_(out[364], out[940], _063557_);
  or g_100582_(_063381_, _063557_, _063568_);
  xor g_100583_(out[359], out[935], _063579_);
  or g_100584_(_063414_, _063579_, _063590_);
  or g_100585_(_063568_, _063590_, _063601_);
  or g_100586_(_063304_, _063480_, _063612_);
  or g_100587_(_063403_, _063612_, _063623_);
  or g_100588_(_063601_, _063623_, _063634_);
  or g_100589_(_063370_, _063634_, _063645_);
  or g_100590_(_063546_, _063645_, _063656_);
  xor g_100591_(out[343], out[935], _063667_);
  and g_100592_(_049400_, out[939], _063678_);
  xor g_100593_(out[350], out[942], _063689_);
  xor g_100594_(out[344], out[936], _063700_);
  xor g_100595_(out[337], out[929], _063711_);
  xor g_100596_(out[349], out[941], _063722_);
  xor g_100597_(out[345], out[937], _063733_);
  xor g_100598_(out[340], out[932], _063744_);
  xor g_100599_(out[338], out[930], _063755_);
  and g_100600_(out[347], _049807_, _063766_);
  xor g_100601_(out[339], out[931], _063777_);
  xor g_100602_(out[342], out[934], _063788_);
  xor g_100603_(out[351], out[943], _063799_);
  xor g_100604_(out[346], out[938], _063810_);
  xor g_100605_(out[341], out[933], _063821_);
  xor g_100606_(out[336], out[928], _063832_);
  or g_100607_(_063689_, _063744_, _063843_);
  or g_100608_(_063700_, _063722_, _063854_);
  or g_100609_(_063755_, _063810_, _063865_);
  or g_100610_(_063854_, _063865_, _063876_);
  or g_100611_(_063733_, _063777_, _063887_);
  or g_100612_(_063821_, _063832_, _063898_);
  or g_100613_(_063887_, _063898_, _063909_);
  or g_100614_(_063876_, _063909_, _063920_);
  xor g_100615_(out[348], out[940], _063931_);
  or g_100616_(_063678_, _063931_, _063942_);
  or g_100617_(_063667_, _063788_, _063953_);
  or g_100618_(_063942_, _063953_, _063964_);
  or g_100619_(_063711_, _063766_, _063975_);
  or g_100620_(_063799_, _063975_, _063986_);
  or g_100621_(_063964_, _063986_, _063997_);
  or g_100622_(_063920_, _063997_, _064008_);
  or g_100623_(_063843_, _064008_, _064019_);
  and g_100624_(out[331], _049807_, _064030_);
  xor g_100625_(out[324], out[932], _064041_);
  xor g_100626_(out[334], out[942], _064052_);
  or g_100627_(_064041_, _064052_, _064063_);
  xor g_100628_(out[333], out[941], _064074_);
  xor g_100629_(out[323], out[931], _064085_);
  xor g_100630_(out[320], out[928], _064096_);
  and g_100631_(_098294_, out[939], _064107_);
  xor g_100632_(out[330], out[938], _064118_);
  xor g_100633_(out[335], out[943], _064129_);
  xor g_100634_(out[326], out[934], _064140_);
  xor g_100635_(out[325], out[933], _064151_);
  xor g_100636_(out[328], out[936], _064162_);
  or g_100637_(_064074_, _064162_, _064173_);
  xor g_100638_(out[322], out[930], _064184_);
  xor g_100639_(out[329], out[937], _064195_);
  xor g_100640_(out[321], out[929], _064206_);
  or g_100641_(_064118_, _064184_, _064217_);
  or g_100642_(_064173_, _064217_, _064228_);
  or g_100643_(_064085_, _064195_, _064239_);
  or g_100644_(_064151_, _064239_, _064250_);
  or g_100645_(_064228_, _064250_, _064261_);
  or g_100646_(_064063_, _064261_, _064272_);
  xor g_100647_(out[332], out[940], _064283_);
  or g_100648_(_064107_, _064283_, _064294_);
  xor g_100649_(out[327], out[935], _064305_);
  or g_100650_(_064140_, _064305_, _064316_);
  or g_100651_(_064294_, _064316_, _064327_);
  or g_100652_(_064030_, _064206_, _064338_);
  or g_100653_(_064129_, _064338_, _064349_);
  or g_100654_(_064327_, _064349_, _064360_);
  or g_100655_(_064096_, _064360_, _064371_);
  or g_100656_(_064272_, _064371_, _064382_);
  xor g_100657_(out[311], out[935], _064393_);
  and g_100658_(_098283_, out[939], _064404_);
  xor g_100659_(out[318], out[942], _064415_);
  xor g_100660_(out[312], out[936], _064426_);
  xor g_100661_(out[305], out[929], _064437_);
  xor g_100662_(out[317], out[941], _064448_);
  xor g_100663_(out[313], out[937], _064459_);
  xor g_100664_(out[308], out[932], _064470_);
  xor g_100665_(out[306], out[930], _064481_);
  and g_100666_(out[315], _049807_, _064492_);
  xor g_100667_(out[307], out[931], _064503_);
  xor g_100668_(out[310], out[934], _064514_);
  xor g_100669_(out[319], out[943], _064525_);
  xor g_100670_(out[314], out[938], _064536_);
  xor g_100671_(out[309], out[933], _064547_);
  xor g_100672_(out[304], out[928], _064558_);
  or g_100673_(_064415_, _064470_, _064569_);
  or g_100674_(_064426_, _064448_, _064580_);
  or g_100675_(_064481_, _064536_, _064591_);
  or g_100676_(_064580_, _064591_, _064602_);
  or g_100677_(_064459_, _064503_, _064613_);
  or g_100678_(_064547_, _064558_, _064624_);
  or g_100679_(_064613_, _064624_, _064635_);
  or g_100680_(_064602_, _064635_, _064646_);
  xor g_100681_(out[316], out[940], _064657_);
  or g_100682_(_064404_, _064657_, _064668_);
  or g_100683_(_064393_, _064514_, _064679_);
  or g_100684_(_064668_, _064679_, _064690_);
  or g_100685_(_064437_, _064492_, _064701_);
  or g_100686_(_064525_, _064701_, _064712_);
  or g_100687_(_064690_, _064712_, _064723_);
  or g_100688_(_064646_, _064723_, _064734_);
  or g_100689_(_064569_, _064734_, _064745_);
  xor g_100690_(out[289], out[929], _064756_);
  and g_100691_(out[299], _049807_, _064767_);
  xor g_100692_(out[297], out[937], _064778_);
  xor g_100693_(out[288], out[928], _064789_);
  xor g_100694_(out[302], out[942], _064800_);
  xor g_100695_(out[292], out[932], _064811_);
  or g_100696_(_064800_, _064811_, _064822_);
  xor g_100697_(out[301], out[941], _064833_);
  xor g_100698_(out[291], out[931], _064844_);
  and g_100699_(_098272_, out[939], _064855_);
  xor g_100700_(out[294], out[934], _064866_);
  xor g_100701_(out[298], out[938], _064877_);
  xor g_100702_(out[293], out[933], _064888_);
  xor g_100703_(out[303], out[943], _064899_);
  xor g_100704_(out[296], out[936], _064910_);
  or g_100705_(_064833_, _064910_, _064921_);
  xor g_100706_(out[290], out[930], _064932_);
  or g_100707_(_064877_, _064932_, _064943_);
  or g_100708_(_064921_, _064943_, _064954_);
  or g_100709_(_064778_, _064844_, _064965_);
  or g_100710_(_064888_, _064965_, _064976_);
  or g_100711_(_064954_, _064976_, _064987_);
  or g_100712_(_064822_, _064987_, _064998_);
  xor g_100713_(out[300], out[940], _065009_);
  or g_100714_(_064855_, _065009_, _065020_);
  xor g_100715_(out[295], out[935], _065031_);
  or g_100716_(_064866_, _065031_, _065042_);
  or g_100717_(_065020_, _065042_, _065053_);
  or g_100718_(_064756_, _064767_, _065064_);
  or g_100719_(_064899_, _065064_, _065075_);
  or g_100720_(_065053_, _065075_, _065086_);
  or g_100721_(_064789_, _065086_, _065097_);
  or g_100722_(_064998_, _065097_, _065108_);
  xor g_100723_(out[279], out[935], _065119_);
  and g_100724_(_098261_, out[939], _065130_);
  xor g_100725_(out[286], out[942], _065141_);
  xor g_100726_(out[280], out[936], _065152_);
  xor g_100727_(out[273], out[929], _065163_);
  xor g_100728_(out[285], out[941], _065174_);
  xor g_100729_(out[281], out[937], _065185_);
  xor g_100730_(out[276], out[932], _065196_);
  xor g_100731_(out[274], out[930], _065207_);
  and g_100732_(out[283], _049807_, _065218_);
  xor g_100733_(out[275], out[931], _065229_);
  xor g_100734_(out[278], out[934], _065240_);
  xor g_100735_(out[287], out[943], _065251_);
  xor g_100736_(out[282], out[938], _065262_);
  xor g_100737_(out[277], out[933], _065273_);
  xor g_100738_(out[272], out[928], _065284_);
  or g_100739_(_065141_, _065196_, _065295_);
  or g_100740_(_065152_, _065174_, _065306_);
  or g_100741_(_065207_, _065262_, _065317_);
  or g_100742_(_065306_, _065317_, _065328_);
  or g_100743_(_065185_, _065229_, _065339_);
  or g_100744_(_065273_, _065284_, _065350_);
  or g_100745_(_065339_, _065350_, _065361_);
  or g_100746_(_065328_, _065361_, _065372_);
  xor g_100747_(out[284], out[940], _065383_);
  or g_100748_(_065130_, _065383_, _065394_);
  or g_100749_(_065119_, _065240_, _065405_);
  or g_100750_(_065394_, _065405_, _065416_);
  or g_100751_(_065163_, _065218_, _065427_);
  or g_100752_(_065251_, _065427_, _065438_);
  or g_100753_(_065416_, _065438_, _065449_);
  or g_100754_(_065372_, _065449_, _065460_);
  or g_100755_(_065295_, _065460_, _065471_);
  xor g_100756_(out[268], out[940], _065482_);
  and g_100757_(_098250_, out[939], _065493_);
  xor g_100758_(out[269], out[941], _065504_);
  xor g_100759_(out[262], out[934], _065515_);
  xor g_100760_(out[264], out[936], _065526_);
  xor g_100761_(out[265], out[937], _065537_);
  xor g_100762_(out[270], out[942], _065548_);
  xor g_100763_(out[260], out[932], _065559_);
  or g_100764_(_065548_, _065559_, _065570_);
  xor g_100765_(out[261], out[933], _065581_);
  xor g_100766_(out[257], out[929], _065592_);
  and g_100767_(out[267], _049807_, _065603_);
  xor g_100768_(out[271], out[943], _065614_);
  xor g_100769_(out[266], out[938], _065625_);
  xor g_100770_(out[256], out[928], _065636_);
  xor g_100771_(out[258], out[930], _065647_);
  xor g_100772_(out[259], out[931], _065658_);
  or g_100773_(_065504_, _065526_, _065669_);
  or g_100774_(_065625_, _065647_, _065680_);
  or g_100775_(_065669_, _065680_, _065691_);
  or g_100776_(_065537_, _065658_, _065702_);
  or g_100777_(_065581_, _065636_, _065713_);
  or g_100778_(_065702_, _065713_, _065724_);
  or g_100779_(_065691_, _065724_, _065735_);
  or g_100780_(_065482_, _065493_, _065746_);
  xor g_100781_(out[263], out[935], _065757_);
  or g_100782_(_065515_, _065757_, _065768_);
  or g_100783_(_065746_, _065768_, _065779_);
  or g_100784_(_065592_, _065603_, _065790_);
  or g_100785_(_065614_, _065790_, _065801_);
  or g_100786_(_065779_, _065801_, _065812_);
  or g_100787_(_065735_, _065812_, _065823_);
  or g_100788_(_065570_, _065823_, _065834_);
  not g_100789_(_065834_, _065845_);
  xor g_100790_(out[247], out[935], _065856_);
  and g_100791_(_098239_, out[939], _065867_);
  xor g_100792_(out[254], out[942], _065878_);
  xor g_100793_(out[248], out[936], _065889_);
  xor g_100794_(out[241], out[929], _065900_);
  xor g_100795_(out[253], out[941], _065911_);
  xor g_100796_(out[249], out[937], _065922_);
  xor g_100797_(out[244], out[932], _065933_);
  xor g_100798_(out[242], out[930], _065944_);
  and g_100799_(out[251], _049807_, _065955_);
  xor g_100800_(out[243], out[931], _065966_);
  xor g_100801_(out[246], out[934], _065977_);
  xor g_100802_(out[255], out[943], _065988_);
  xor g_100803_(out[250], out[938], _065999_);
  xor g_100804_(out[245], out[933], _066010_);
  xor g_100805_(out[240], out[928], _066021_);
  or g_100806_(_065878_, _065933_, _066032_);
  or g_100807_(_065889_, _065911_, _066043_);
  or g_100808_(_065944_, _065999_, _066054_);
  or g_100809_(_066043_, _066054_, _066065_);
  or g_100810_(_065922_, _065966_, _066076_);
  or g_100811_(_066010_, _066021_, _066087_);
  or g_100812_(_066076_, _066087_, _066098_);
  or g_100813_(_066065_, _066098_, _066109_);
  xor g_100814_(out[252], out[940], _066120_);
  or g_100815_(_065867_, _066120_, _066131_);
  or g_100816_(_065856_, _065977_, _066142_);
  or g_100817_(_066131_, _066142_, _066153_);
  or g_100818_(_065900_, _065955_, _066164_);
  or g_100819_(_065988_, _066164_, _066175_);
  or g_100820_(_066153_, _066175_, _066186_);
  or g_100821_(_066109_, _066186_, _066197_);
  or g_100822_(_066032_, _066197_, _066208_);
  xor g_100823_(out[236], out[940], _066219_);
  and g_100824_(_098228_, out[939], _066230_);
  xor g_100825_(out[232], out[936], _066241_);
  xor g_100826_(out[230], out[934], _066252_);
  xor g_100827_(out[237], out[941], _066263_);
  xor g_100828_(out[238], out[942], _066274_);
  xor g_100829_(out[226], out[930], _066285_);
  xor g_100830_(out[233], out[937], _066296_);
  xor g_100831_(out[229], out[933], _066307_);
  xor g_100832_(out[225], out[929], _066318_);
  and g_100833_(out[235], _049807_, _066329_);
  or g_100834_(_066241_, _066263_, _066340_);
  xor g_100835_(out[239], out[943], _066351_);
  xor g_100836_(out[234], out[938], _066362_);
  xor g_100837_(out[228], out[932], _066373_);
  xor g_100838_(out[227], out[931], _066384_);
  xor g_100839_(out[224], out[928], _066395_);
  or g_100840_(_066285_, _066362_, _066406_);
  or g_100841_(_066340_, _066406_, _066417_);
  or g_100842_(_066296_, _066384_, _066428_);
  or g_100843_(_066307_, _066428_, _066439_);
  or g_100844_(_066417_, _066439_, _066450_);
  or g_100845_(_066274_, _066373_, _066461_);
  or g_100846_(_066450_, _066461_, _066472_);
  or g_100847_(_066219_, _066230_, _066483_);
  xor g_100848_(out[231], out[935], _066494_);
  or g_100849_(_066252_, _066494_, _066505_);
  or g_100850_(_066483_, _066505_, _066516_);
  or g_100851_(_066318_, _066329_, _066527_);
  or g_100852_(_066351_, _066527_, _066538_);
  or g_100853_(_066516_, _066538_, _066549_);
  or g_100854_(_066395_, _066549_, _066560_);
  or g_100855_(_066472_, _066560_, _066571_);
  xor g_100856_(out[215], out[935], _066582_);
  and g_100857_(_098217_, out[939], _066593_);
  xor g_100858_(out[222], out[942], _066604_);
  xor g_100859_(out[216], out[936], _066615_);
  xor g_100860_(out[209], out[929], _066626_);
  xor g_100861_(out[221], out[941], _066637_);
  xor g_100862_(out[217], out[937], _066648_);
  xor g_100863_(out[212], out[932], _066659_);
  xor g_100864_(out[210], out[930], _066670_);
  and g_100865_(out[219], _049807_, _066681_);
  xor g_100866_(out[211], out[931], _066692_);
  xor g_100867_(out[214], out[934], _066703_);
  xor g_100868_(out[223], out[943], _066714_);
  xor g_100869_(out[218], out[938], _066725_);
  xor g_100870_(out[213], out[933], _066736_);
  xor g_100871_(out[208], out[928], _066747_);
  or g_100872_(_066604_, _066659_, _066758_);
  or g_100873_(_066615_, _066637_, _066769_);
  or g_100874_(_066670_, _066725_, _066780_);
  or g_100875_(_066769_, _066780_, _066791_);
  or g_100876_(_066648_, _066692_, _066802_);
  or g_100877_(_066736_, _066747_, _066813_);
  or g_100878_(_066802_, _066813_, _066824_);
  or g_100879_(_066791_, _066824_, _066835_);
  xor g_100880_(out[220], out[940], _066846_);
  or g_100881_(_066593_, _066846_, _066857_);
  or g_100882_(_066582_, _066703_, _066868_);
  or g_100883_(_066857_, _066868_, _066879_);
  or g_100884_(_066626_, _066681_, _066890_);
  or g_100885_(_066714_, _066890_, _066901_);
  or g_100886_(_066879_, _066901_, _066912_);
  or g_100887_(_066835_, _066912_, _066923_);
  or g_100888_(_066758_, _066923_, _066934_);
  xor g_100889_(out[193], out[929], _066945_);
  and g_100890_(out[203], _049807_, _066956_);
  xor g_100891_(out[201], out[937], _066967_);
  xor g_100892_(out[192], out[928], _066978_);
  xor g_100893_(out[206], out[942], _066989_);
  xor g_100894_(out[196], out[932], _067000_);
  or g_100895_(_066989_, _067000_, _067011_);
  xor g_100896_(out[205], out[941], _067022_);
  xor g_100897_(out[195], out[931], _067033_);
  and g_100898_(_098206_, out[939], _067044_);
  xor g_100899_(out[198], out[934], _067055_);
  xor g_100900_(out[202], out[938], _067066_);
  xor g_100901_(out[197], out[933], _067077_);
  xor g_100902_(out[207], out[943], _067088_);
  xor g_100903_(out[200], out[936], _067099_);
  or g_100904_(_067022_, _067099_, _067110_);
  xor g_100905_(out[194], out[930], _067121_);
  or g_100906_(_067066_, _067121_, _067132_);
  or g_100907_(_067110_, _067132_, _067143_);
  or g_100908_(_066967_, _067033_, _067154_);
  or g_100909_(_067077_, _067154_, _067165_);
  or g_100910_(_067143_, _067165_, _067176_);
  or g_100911_(_067011_, _067176_, _067187_);
  xor g_100912_(out[204], out[940], _067198_);
  or g_100913_(_067044_, _067198_, _067209_);
  xor g_100914_(out[199], out[935], _067220_);
  or g_100915_(_067055_, _067220_, _067231_);
  or g_100916_(_067209_, _067231_, _067242_);
  or g_100917_(_066945_, _066956_, _067253_);
  or g_100918_(_067088_, _067253_, _067264_);
  or g_100919_(_067242_, _067264_, _067275_);
  or g_100920_(_066978_, _067275_, _067286_);
  or g_100921_(_067187_, _067286_, _067297_);
  xor g_100922_(out[183], out[935], _067308_);
  and g_100923_(_098195_, out[939], _067319_);
  xor g_100924_(out[190], out[942], _067330_);
  xor g_100925_(out[184], out[936], _067341_);
  xor g_100926_(out[177], out[929], _067352_);
  xor g_100927_(out[189], out[941], _067363_);
  xor g_100928_(out[185], out[937], _067374_);
  xor g_100929_(out[180], out[932], _067385_);
  xor g_100930_(out[178], out[930], _067396_);
  and g_100931_(out[187], _049807_, _067407_);
  xor g_100932_(out[179], out[931], _067418_);
  xor g_100933_(out[182], out[934], _067429_);
  xor g_100934_(out[191], out[943], _067440_);
  xor g_100935_(out[186], out[938], _067451_);
  xor g_100936_(out[181], out[933], _067462_);
  xor g_100937_(out[176], out[928], _067473_);
  or g_100938_(_067330_, _067385_, _067484_);
  or g_100939_(_067341_, _067363_, _067495_);
  or g_100940_(_067396_, _067451_, _067506_);
  or g_100941_(_067495_, _067506_, _067517_);
  or g_100942_(_067374_, _067418_, _067528_);
  or g_100943_(_067462_, _067473_, _067539_);
  or g_100944_(_067528_, _067539_, _067550_);
  or g_100945_(_067517_, _067550_, _067561_);
  xor g_100946_(out[188], out[940], _067572_);
  or g_100947_(_067319_, _067572_, _067583_);
  or g_100948_(_067308_, _067429_, _067594_);
  or g_100949_(_067583_, _067594_, _067605_);
  or g_100950_(_067352_, _067407_, _067616_);
  or g_100951_(_067440_, _067616_, _067627_);
  or g_100952_(_067605_, _067627_, _067638_);
  or g_100953_(_067561_, _067638_, _067649_);
  or g_100954_(_067484_, _067649_, _067660_);
  xor g_100955_(out[161], out[929], _067671_);
  and g_100956_(_098184_, out[939], _067682_);
  and g_100957_(out[171], _049807_, _067693_);
  xor g_100958_(out[174], out[942], _067704_);
  xor g_100959_(out[163], out[931], _067715_);
  xor g_100960_(out[164], out[932], _067726_);
  xor g_100961_(out[162], out[930], _067737_);
  xor g_100962_(out[169], out[937], _067748_);
  xor g_100963_(out[160], out[928], _067759_);
  xor g_100964_(out[172], out[940], _067770_);
  xor g_100965_(out[166], out[934], _067781_);
  xor g_100966_(out[170], out[938], _067792_);
  xor g_100967_(out[165], out[933], _067803_);
  xor g_100968_(out[175], out[943], _067814_);
  xor g_100969_(out[173], out[941], _067825_);
  xor g_100970_(out[168], out[936], _067836_);
  or g_100971_(_067704_, _067726_, _067847_);
  or g_100972_(_067825_, _067836_, _067858_);
  or g_100973_(_067737_, _067792_, _067869_);
  or g_100974_(_067858_, _067869_, _067880_);
  or g_100975_(_067715_, _067748_, _067891_);
  or g_100976_(_067759_, _067803_, _067902_);
  or g_100977_(_067891_, _067902_, _067913_);
  or g_100978_(_067880_, _067913_, _067924_);
  or g_100979_(_067682_, _067770_, _067935_);
  xor g_100980_(out[167], out[935], _067946_);
  or g_100981_(_067781_, _067946_, _067957_);
  or g_100982_(_067935_, _067957_, _067968_);
  or g_100983_(_067671_, _067693_, _067979_);
  or g_100984_(_067814_, _067979_, _067990_);
  or g_100985_(_067968_, _067990_, _068001_);
  or g_100986_(_067924_, _068001_, _068012_);
  or g_100987_(_067847_, _068012_, _068023_);
  xor g_100988_(out[151], out[935], _068034_);
  and g_100989_(_098173_, out[939], _068045_);
  xor g_100990_(out[158], out[942], _068056_);
  xor g_100991_(out[152], out[936], _068067_);
  xor g_100992_(out[145], out[929], _068078_);
  xor g_100993_(out[157], out[941], _068089_);
  xor g_100994_(out[153], out[937], _068100_);
  xor g_100995_(out[148], out[932], _068111_);
  xor g_100996_(out[146], out[930], _068122_);
  and g_100997_(out[155], _049807_, _068133_);
  xor g_100998_(out[147], out[931], _068144_);
  xor g_100999_(out[150], out[934], _068155_);
  xor g_101000_(out[159], out[943], _068166_);
  xor g_101001_(out[154], out[938], _068177_);
  xor g_101002_(out[149], out[933], _068188_);
  xor g_101003_(out[144], out[928], _068199_);
  or g_101004_(_068056_, _068111_, _068210_);
  or g_101005_(_068067_, _068089_, _068221_);
  or g_101006_(_068122_, _068177_, _068232_);
  or g_101007_(_068221_, _068232_, _068243_);
  or g_101008_(_068100_, _068144_, _068254_);
  or g_101009_(_068188_, _068199_, _068265_);
  or g_101010_(_068254_, _068265_, _068276_);
  or g_101011_(_068243_, _068276_, _068287_);
  xor g_101012_(out[156], out[940], _068298_);
  or g_101013_(_068045_, _068298_, _068309_);
  or g_101014_(_068034_, _068155_, _068320_);
  or g_101015_(_068309_, _068320_, _068331_);
  or g_101016_(_068078_, _068133_, _068342_);
  or g_101017_(_068166_, _068342_, _068353_);
  or g_101018_(_068331_, _068353_, _068364_);
  or g_101019_(_068287_, _068364_, _068375_);
  or g_101020_(_068210_, _068375_, _068386_);
  xor g_101021_(out[129], out[929], _068397_);
  and g_101022_(out[139], _049807_, _068408_);
  xor g_101023_(out[137], out[937], _068419_);
  xor g_101024_(out[128], out[928], _068430_);
  xor g_101025_(out[142], out[942], _068441_);
  xor g_101026_(out[132], out[932], _068452_);
  or g_101027_(_068441_, _068452_, _068463_);
  xor g_101028_(out[141], out[941], _068474_);
  xor g_101029_(out[131], out[931], _068485_);
  and g_101030_(_098162_, out[939], _068496_);
  xor g_101031_(out[134], out[934], _068507_);
  xor g_101032_(out[138], out[938], _068518_);
  xor g_101033_(out[133], out[933], _068529_);
  xor g_101034_(out[143], out[943], _068540_);
  xor g_101035_(out[136], out[936], _068551_);
  or g_101036_(_068474_, _068551_, _068562_);
  xor g_101037_(out[130], out[930], _068573_);
  or g_101038_(_068518_, _068573_, _068584_);
  or g_101039_(_068562_, _068584_, _068595_);
  or g_101040_(_068419_, _068485_, _068606_);
  or g_101041_(_068529_, _068606_, _068617_);
  or g_101042_(_068595_, _068617_, _068628_);
  or g_101043_(_068463_, _068628_, _068639_);
  xor g_101044_(out[140], out[940], _068650_);
  or g_101045_(_068496_, _068650_, _068661_);
  xor g_101046_(out[135], out[935], _068672_);
  or g_101047_(_068507_, _068672_, _068683_);
  or g_101048_(_068661_, _068683_, _068694_);
  or g_101049_(_068397_, _068408_, _068705_);
  or g_101050_(_068540_, _068705_, _068716_);
  or g_101051_(_068694_, _068716_, _068727_);
  or g_101052_(_068430_, _068727_, _068738_);
  or g_101053_(_068639_, _068738_, _068749_);
  xor g_101054_(out[119], out[935], _068760_);
  and g_101055_(_098151_, out[939], _068771_);
  xor g_101056_(out[126], out[942], _068782_);
  xor g_101057_(out[120], out[936], _068793_);
  xor g_101058_(out[113], out[929], _068804_);
  xor g_101059_(out[125], out[941], _068815_);
  xor g_101060_(out[121], out[937], _068826_);
  xor g_101061_(out[116], out[932], _068837_);
  xor g_101062_(out[114], out[930], _068848_);
  and g_101063_(out[123], _049807_, _068859_);
  xor g_101064_(out[115], out[931], _068870_);
  xor g_101065_(out[118], out[934], _068881_);
  xor g_101066_(out[127], out[943], _068892_);
  xor g_101067_(out[122], out[938], _068903_);
  xor g_101068_(out[117], out[933], _068914_);
  xor g_101069_(out[112], out[928], _068925_);
  or g_101070_(_068782_, _068837_, _068936_);
  or g_101071_(_068793_, _068815_, _068947_);
  or g_101072_(_068848_, _068903_, _068958_);
  or g_101073_(_068947_, _068958_, _068969_);
  or g_101074_(_068826_, _068870_, _068980_);
  or g_101075_(_068914_, _068925_, _068991_);
  or g_101076_(_068980_, _068991_, _069002_);
  or g_101077_(_068969_, _069002_, _069013_);
  xor g_101078_(out[124], out[940], _069024_);
  or g_101079_(_068771_, _069024_, _069035_);
  or g_101080_(_068760_, _068881_, _069046_);
  or g_101081_(_069035_, _069046_, _069057_);
  or g_101082_(_068804_, _068859_, _069068_);
  or g_101083_(_068892_, _069068_, _069079_);
  or g_101084_(_069057_, _069079_, _069090_);
  or g_101085_(_069013_, _069090_, _069101_);
  or g_101086_(_068936_, _069101_, _069112_);
  xor g_101087_(out[104], out[936], _069123_);
  xor g_101088_(out[101], out[933], _069134_);
  xor g_101089_(out[99], out[931], _069145_);
  xor g_101090_(out[110], out[942], _069156_);
  xor g_101091_(out[109], out[941], _069167_);
  xor g_101092_(out[98], out[930], _069178_);
  xor g_101093_(out[105], out[937], _069189_);
  xor g_101094_(out[102], out[934], _069200_);
  xor g_101095_(out[111], out[943], _069211_);
  xor g_101096_(out[106], out[938], _069222_);
  xor g_101097_(out[100], out[932], _069233_);
  xor g_101098_(out[96], out[928], _069244_);
  and g_101099_(_098140_, out[939], _069255_);
  and g_101100_(out[107], _049807_, _069266_);
  or g_101101_(_069123_, _069167_, _069277_);
  xor g_101102_(out[97], out[929], _069288_);
  or g_101103_(_069178_, _069222_, _069299_);
  or g_101104_(_069277_, _069299_, _069310_);
  or g_101105_(_069145_, _069189_, _069321_);
  or g_101106_(_069134_, _069321_, _069332_);
  or g_101107_(_069310_, _069332_, _069343_);
  or g_101108_(_069156_, _069233_, _069354_);
  or g_101109_(_069343_, _069354_, _069365_);
  xor g_101110_(out[108], out[940], _069376_);
  or g_101111_(_069255_, _069376_, _069387_);
  xor g_101112_(out[103], out[935], _069398_);
  or g_101113_(_069200_, _069398_, _069409_);
  or g_101114_(_069387_, _069409_, _069420_);
  or g_101115_(_069266_, _069288_, _069431_);
  or g_101116_(_069211_, _069431_, _069442_);
  or g_101117_(_069420_, _069442_, _069453_);
  or g_101118_(_069244_, _069453_, _069464_);
  or g_101119_(_069365_, _069464_, _069475_);
  not g_101120_(_069475_, _069486_);
  xor g_101121_(out[87], out[935], _069497_);
  and g_101122_(_098129_, out[939], _069508_);
  xor g_101123_(out[94], out[942], _069519_);
  xor g_101124_(out[88], out[936], _069530_);
  xor g_101125_(out[81], out[929], _069541_);
  xor g_101126_(out[93], out[941], _069552_);
  xor g_101127_(out[89], out[937], _069563_);
  xor g_101128_(out[84], out[932], _069574_);
  xor g_101129_(out[82], out[930], _069585_);
  and g_101130_(out[91], _049807_, _069596_);
  xor g_101131_(out[83], out[931], _069607_);
  xor g_101132_(out[86], out[934], _069618_);
  xor g_101133_(out[95], out[943], _069629_);
  xor g_101134_(out[90], out[938], _069640_);
  xor g_101135_(out[85], out[933], _069651_);
  xor g_101136_(out[80], out[928], _069662_);
  or g_101137_(_069519_, _069574_, _069673_);
  or g_101138_(_069530_, _069552_, _069684_);
  or g_101139_(_069585_, _069640_, _069695_);
  or g_101140_(_069684_, _069695_, _069706_);
  or g_101141_(_069563_, _069607_, _069717_);
  or g_101142_(_069651_, _069662_, _069728_);
  or g_101143_(_069717_, _069728_, _069739_);
  or g_101144_(_069706_, _069739_, _069750_);
  xor g_101145_(out[92], out[940], _069761_);
  or g_101146_(_069508_, _069761_, _069772_);
  or g_101147_(_069497_, _069618_, _069783_);
  or g_101148_(_069772_, _069783_, _069794_);
  or g_101149_(_069541_, _069596_, _069805_);
  or g_101150_(_069629_, _069805_, _069816_);
  or g_101151_(_069794_, _069816_, _069827_);
  or g_101152_(_069750_, _069827_, _069838_);
  or g_101153_(_069673_, _069838_, _069849_);
  not g_101154_(_069849_, _069860_);
  and g_101155_(out[75], _049807_, _069871_);
  xor g_101156_(out[68], out[932], _069882_);
  xor g_101157_(out[66], out[930], _069893_);
  xor g_101158_(out[73], out[937], _069904_);
  xor g_101159_(out[64], out[928], _069915_);
  xor g_101160_(out[67], out[931], _069926_);
  and g_101161_(_098118_, out[939], _069937_);
  xor g_101162_(out[74], out[938], _069948_);
  xor g_101163_(out[79], out[943], _069959_);
  xor g_101164_(out[70], out[934], _069970_);
  xor g_101165_(out[69], out[933], _069981_);
  xor g_101166_(out[77], out[941], _069992_);
  xor g_101167_(out[78], out[942], _070003_);
  xor g_101168_(out[72], out[936], _070014_);
  xor g_101169_(out[65], out[929], _070025_);
  or g_101170_(_069882_, _070003_, _070036_);
  or g_101171_(_069992_, _070014_, _070047_);
  or g_101172_(_069893_, _069948_, _070058_);
  or g_101173_(_070047_, _070058_, _070069_);
  or g_101174_(_069904_, _069926_, _070080_);
  or g_101175_(_069915_, _069981_, _070091_);
  or g_101176_(_070080_, _070091_, _070102_);
  or g_101177_(_070069_, _070102_, _070113_);
  xor g_101178_(out[76], out[940], _070124_);
  or g_101179_(_069937_, _070124_, _070135_);
  xor g_101180_(out[71], out[935], _070146_);
  or g_101181_(_069970_, _070146_, _070157_);
  or g_101182_(_070135_, _070157_, _070168_);
  or g_101183_(_069871_, _070025_, _070179_);
  or g_101184_(_069959_, _070179_, _070190_);
  or g_101185_(_070168_, _070190_, _070201_);
  or g_101186_(_070113_, _070201_, _070212_);
  or g_101187_(_070036_, _070212_, _070223_);
  xor g_101188_(out[55], out[935], _070234_);
  and g_101189_(_098107_, out[939], _070245_);
  xor g_101190_(out[62], out[942], _070256_);
  xor g_101191_(out[56], out[936], _070267_);
  xor g_101192_(out[49], out[929], _070278_);
  xor g_101193_(out[61], out[941], _070289_);
  xor g_101194_(out[57], out[937], _070300_);
  xor g_101195_(out[52], out[932], _070311_);
  xor g_101196_(out[50], out[930], _070322_);
  and g_101197_(out[59], _049807_, _070333_);
  xor g_101198_(out[51], out[931], _070344_);
  xor g_101199_(out[54], out[934], _070355_);
  xor g_101200_(out[63], out[943], _070366_);
  xor g_101201_(out[58], out[938], _070377_);
  xor g_101202_(out[53], out[933], _070388_);
  xor g_101203_(out[48], out[928], _070399_);
  or g_101204_(_070256_, _070311_, _070410_);
  or g_101205_(_070267_, _070289_, _070421_);
  or g_101206_(_070322_, _070377_, _070432_);
  or g_101207_(_070421_, _070432_, _070443_);
  or g_101208_(_070300_, _070344_, _070454_);
  or g_101209_(_070388_, _070399_, _070465_);
  or g_101210_(_070454_, _070465_, _070476_);
  or g_101211_(_070443_, _070476_, _070487_);
  xor g_101212_(out[60], out[940], _070498_);
  or g_101213_(_070245_, _070498_, _070509_);
  or g_101214_(_070234_, _070355_, _070520_);
  or g_101215_(_070509_, _070520_, _070531_);
  or g_101216_(_070278_, _070333_, _070542_);
  or g_101217_(_070366_, _070542_, _070553_);
  or g_101218_(_070531_, _070553_, _070564_);
  or g_101219_(_070487_, _070564_, _070575_);
  or g_101220_(_070410_, _070575_, _070586_);
  xor g_101221_(out[33], out[929], _070597_);
  and g_101222_(out[43], _049807_, _070608_);
  xor g_101223_(out[41], out[937], _070619_);
  xor g_101224_(out[32], out[928], _070630_);
  xor g_101225_(out[46], out[942], _070641_);
  xor g_101226_(out[36], out[932], _070652_);
  or g_101227_(_070641_, _070652_, _070663_);
  xor g_101228_(out[45], out[941], _070674_);
  xor g_101229_(out[35], out[931], _070685_);
  and g_101230_(_098096_, out[939], _070696_);
  xor g_101231_(out[38], out[934], _070707_);
  xor g_101232_(out[42], out[938], _070718_);
  xor g_101233_(out[37], out[933], _070729_);
  xor g_101234_(out[47], out[943], _070740_);
  xor g_101235_(out[40], out[936], _070751_);
  or g_101236_(_070674_, _070751_, _070762_);
  xor g_101237_(out[34], out[930], _070773_);
  or g_101238_(_070718_, _070773_, _070784_);
  or g_101239_(_070762_, _070784_, _070795_);
  or g_101240_(_070619_, _070685_, _070806_);
  or g_101241_(_070729_, _070806_, _070817_);
  or g_101242_(_070795_, _070817_, _070828_);
  or g_101243_(_070663_, _070828_, _070839_);
  xor g_101244_(out[44], out[940], _070850_);
  or g_101245_(_070696_, _070850_, _070861_);
  xor g_101246_(out[39], out[935], _070872_);
  or g_101247_(_070707_, _070872_, _070883_);
  or g_101248_(_070861_, _070883_, _070894_);
  or g_101249_(_070597_, _070608_, _070905_);
  or g_101250_(_070740_, _070905_, _070916_);
  or g_101251_(_070894_, _070916_, _070927_);
  or g_101252_(_070630_, _070927_, _070938_);
  or g_101253_(_070839_, _070938_, _070949_);
  xor g_101254_(out[23], out[935], _070960_);
  and g_101255_(_098063_, out[939], _070971_);
  xor g_101256_(out[30], out[942], _070982_);
  xor g_101257_(out[24], out[936], _070993_);
  xor g_101258_(out[17], out[929], _071004_);
  xor g_101259_(out[29], out[941], _071015_);
  xor g_101260_(out[25], out[937], _071026_);
  xor g_101261_(out[20], out[932], _071037_);
  xor g_101262_(out[18], out[930], _071048_);
  and g_101263_(out[27], _049807_, _071059_);
  xor g_101264_(out[19], out[931], _071070_);
  xor g_101265_(out[22], out[934], _071081_);
  xor g_101266_(out[31], out[943], _071092_);
  xor g_101267_(out[26], out[938], _071103_);
  xor g_101268_(out[21], out[933], _071114_);
  xor g_101269_(out[16], out[928], _071125_);
  or g_101270_(_070982_, _071037_, _071136_);
  or g_101271_(_070993_, _071015_, _071147_);
  or g_101272_(_071048_, _071103_, _071158_);
  or g_101273_(_071147_, _071158_, _071169_);
  or g_101274_(_071026_, _071070_, _071180_);
  or g_101275_(_071114_, _071125_, _071191_);
  or g_101276_(_071180_, _071191_, _071202_);
  or g_101277_(_071169_, _071202_, _071213_);
  xor g_101278_(out[28], out[940], _071224_);
  or g_101279_(_070971_, _071224_, _071235_);
  or g_101280_(_070960_, _071081_, _071246_);
  or g_101281_(_071235_, _071246_, _071257_);
  or g_101282_(_071004_, _071059_, _071268_);
  or g_101283_(_071092_, _071268_, _071279_);
  or g_101284_(_071257_, _071279_, _071290_);
  or g_101285_(_071213_, _071290_, _071301_);
  or g_101286_(_071136_, _071301_, _071312_);
  xor g_101287_(out[1], out[929], _071323_);
  and g_101288_(_098041_, out[939], _071334_);
  and g_101289_(out[11], _049807_, _071345_);
  xor g_101290_(out[9], out[937], _071356_);
  xor g_101291_(out[0], out[928], _071367_);
  xor g_101292_(out[14], out[942], _071378_);
  xor g_101293_(out[4], out[932], _071389_);
  or g_101294_(_071378_, _071389_, _071400_);
  xor g_101295_(out[13], out[941], _071411_);
  xor g_101296_(out[3], out[931], _071422_);
  xor g_101297_(out[12], out[940], _071433_);
  xor g_101298_(out[6], out[934], _071444_);
  xor g_101299_(out[10], out[938], _071455_);
  xor g_101300_(out[5], out[933], _071466_);
  xor g_101301_(out[15], out[943], _071477_);
  xor g_101302_(out[8], out[936], _071488_);
  or g_101303_(_071411_, _071488_, _071499_);
  xor g_101304_(out[2], out[930], _071510_);
  or g_101305_(_071455_, _071510_, _071521_);
  or g_101306_(_071499_, _071521_, _071532_);
  or g_101307_(_071356_, _071422_, _071543_);
  or g_101308_(_071466_, _071543_, _071554_);
  or g_101309_(_071532_, _071554_, _071565_);
  or g_101310_(_071400_, _071565_, _071576_);
  or g_101311_(_071334_, _071433_, _071587_);
  xor g_101312_(out[7], out[935], _071598_);
  or g_101313_(_071444_, _071598_, _071609_);
  or g_101314_(_071587_, _071609_, _071620_);
  or g_101315_(_071323_, _071345_, _071631_);
  or g_101316_(_071477_, _071631_, _071642_);
  or g_101317_(_071620_, _071642_, _071653_);
  or g_101318_(_071367_, _071653_, _071664_);
  or g_101319_(_071576_, _071664_, _071675_);
  not g_101320_(_071675_, _071686_);
  xor g_101321_(out[467], out[915], _071697_);
  xor g_101322_(out[468], out[916], _071708_);
  xor g_101323_(out[478], out[926], _071719_);
  xor g_101324_(out[466], out[914], _071730_);
  xor g_101325_(out[469], out[917], _071741_);
  xor g_101326_(out[473], out[921], _071752_);
  xor g_101327_(out[472], out[920], _071763_);
  xor g_101328_(out[479], out[927], _071774_);
  xor g_101329_(out[474], out[922], _071785_);
  xor g_101330_(out[470], out[918], _071796_);
  xor g_101331_(out[464], out[912], _071807_);
  and g_101332_(_049499_, out[923], _071818_);
  and g_101333_(out[475], _049796_, _071829_);
  xor g_101334_(out[477], out[925], _071840_);
  or g_101335_(_071763_, _071840_, _071851_);
  xor g_101336_(out[465], out[913], _071862_);
  or g_101337_(_071730_, _071785_, _071873_);
  or g_101338_(_071851_, _071873_, _071884_);
  or g_101339_(_071697_, _071752_, _071895_);
  or g_101340_(_071741_, _071895_, _071906_);
  or g_101341_(_071884_, _071906_, _071917_);
  or g_101342_(_071708_, _071719_, _071928_);
  or g_101343_(_071917_, _071928_, _071939_);
  xor g_101344_(out[476], out[924], _071950_);
  or g_101345_(_071818_, _071950_, _071961_);
  xor g_101346_(out[471], out[919], _071972_);
  or g_101347_(_071796_, _071972_, _071983_);
  or g_101348_(_071961_, _071983_, _071994_);
  or g_101349_(_071829_, _071862_, _072005_);
  or g_101350_(_071774_, _072005_, _072016_);
  or g_101351_(_071994_, _072016_, _072027_);
  or g_101352_(_071807_, _072027_, _072038_);
  or g_101353_(_071939_, _072038_, _072049_);
  not g_101354_(_072049_, _072060_);
  xor g_101355_(out[455], out[919], _072071_);
  and g_101356_(_049477_, out[923], _072082_);
  xor g_101357_(out[462], out[926], _072093_);
  xor g_101358_(out[456], out[920], _072104_);
  xor g_101359_(out[449], out[913], _072115_);
  xor g_101360_(out[461], out[925], _072126_);
  xor g_101361_(out[457], out[921], _072137_);
  xor g_101362_(out[452], out[916], _072148_);
  xor g_101363_(out[450], out[914], _072159_);
  and g_101364_(out[459], _049796_, _072170_);
  xor g_101365_(out[451], out[915], _072181_);
  xor g_101366_(out[454], out[918], _072192_);
  xor g_101367_(out[463], out[927], _072203_);
  xor g_101368_(out[458], out[922], _072214_);
  xor g_101369_(out[453], out[917], _072225_);
  xor g_101370_(out[448], out[912], _072236_);
  or g_101371_(_072093_, _072148_, _072247_);
  or g_101372_(_072104_, _072126_, _072258_);
  or g_101373_(_072159_, _072214_, _072269_);
  or g_101374_(_072258_, _072269_, _072280_);
  or g_101375_(_072137_, _072181_, _072291_);
  or g_101376_(_072225_, _072236_, _072302_);
  or g_101377_(_072291_, _072302_, _072313_);
  or g_101378_(_072280_, _072313_, _072324_);
  xor g_101379_(out[460], out[924], _072335_);
  or g_101380_(_072082_, _072335_, _072346_);
  or g_101381_(_072071_, _072192_, _072357_);
  or g_101382_(_072346_, _072357_, _072368_);
  or g_101383_(_072115_, _072170_, _072379_);
  or g_101384_(_072203_, _072379_, _072390_);
  or g_101385_(_072368_, _072390_, _072401_);
  or g_101386_(_072324_, _072401_, _072412_);
  or g_101387_(_072247_, _072412_, _072423_);
  not g_101388_(_072423_, _072434_);
  xor g_101389_(out[433], out[913], _072445_);
  and g_101390_(out[443], _049796_, _072456_);
  xor g_101391_(out[441], out[921], _072467_);
  xor g_101392_(out[432], out[912], _072478_);
  xor g_101393_(out[446], out[926], _072489_);
  xor g_101394_(out[436], out[916], _072500_);
  or g_101395_(_072489_, _072500_, _072511_);
  xor g_101396_(out[445], out[925], _072522_);
  xor g_101397_(out[435], out[915], _072533_);
  and g_101398_(_049466_, out[923], _072544_);
  xor g_101399_(out[438], out[918], _072555_);
  xor g_101400_(out[442], out[922], _072566_);
  xor g_101401_(out[437], out[917], _072577_);
  xor g_101402_(out[447], out[927], _072588_);
  xor g_101403_(out[440], out[920], _072599_);
  or g_101404_(_072522_, _072599_, _072610_);
  xor g_101405_(out[434], out[914], _072621_);
  or g_101406_(_072566_, _072621_, _072632_);
  or g_101407_(_072610_, _072632_, _072643_);
  or g_101408_(_072467_, _072533_, _072654_);
  or g_101409_(_072577_, _072654_, _072665_);
  or g_101410_(_072643_, _072665_, _072676_);
  or g_101411_(_072511_, _072676_, _072687_);
  xor g_101412_(out[444], out[924], _072698_);
  or g_101413_(_072544_, _072698_, _072709_);
  xor g_101414_(out[439], out[919], _072720_);
  or g_101415_(_072555_, _072720_, _072731_);
  or g_101416_(_072709_, _072731_, _072742_);
  or g_101417_(_072445_, _072456_, _072753_);
  or g_101418_(_072588_, _072753_, _072764_);
  or g_101419_(_072742_, _072764_, _072775_);
  or g_101420_(_072478_, _072775_, _072786_);
  or g_101421_(_072687_, _072786_, _072797_);
  xor g_101422_(out[423], out[919], _072808_);
  and g_101423_(_049455_, out[923], _072819_);
  xor g_101424_(out[430], out[926], _072830_);
  xor g_101425_(out[424], out[920], _072841_);
  xor g_101426_(out[417], out[913], _072852_);
  xor g_101427_(out[429], out[925], _072863_);
  xor g_101428_(out[425], out[921], _072874_);
  xor g_101429_(out[420], out[916], _072885_);
  xor g_101430_(out[418], out[914], _072896_);
  and g_101431_(out[427], _049796_, _072907_);
  xor g_101432_(out[419], out[915], _072918_);
  xor g_101433_(out[422], out[918], _072929_);
  xor g_101434_(out[431], out[927], _072940_);
  xor g_101435_(out[426], out[922], _072951_);
  xor g_101436_(out[421], out[917], _072962_);
  xor g_101437_(out[416], out[912], _072973_);
  or g_101438_(_072830_, _072885_, _072984_);
  or g_101439_(_072841_, _072863_, _072995_);
  or g_101440_(_072896_, _072951_, _073006_);
  or g_101441_(_072995_, _073006_, _073017_);
  or g_101442_(_072874_, _072918_, _073028_);
  or g_101443_(_072962_, _072973_, _073039_);
  or g_101444_(_073028_, _073039_, _073050_);
  or g_101445_(_073017_, _073050_, _073061_);
  xor g_101446_(out[428], out[924], _073072_);
  or g_101447_(_072819_, _073072_, _073083_);
  or g_101448_(_072808_, _072929_, _073094_);
  or g_101449_(_073083_, _073094_, _073105_);
  or g_101450_(_072852_, _072907_, _073116_);
  or g_101451_(_072940_, _073116_, _073127_);
  or g_101452_(_073105_, _073127_, _073138_);
  or g_101453_(_073061_, _073138_, _073149_);
  or g_101454_(_072984_, _073149_, _073160_);
  xor g_101455_(out[408], out[920], _073171_);
  xor g_101456_(out[405], out[917], _073182_);
  xor g_101457_(out[403], out[915], _073193_);
  xor g_101458_(out[414], out[926], _073204_);
  xor g_101459_(out[413], out[925], _073215_);
  xor g_101460_(out[402], out[914], _073226_);
  xor g_101461_(out[409], out[921], _073237_);
  xor g_101462_(out[406], out[918], _073248_);
  xor g_101463_(out[415], out[927], _073259_);
  xor g_101464_(out[410], out[922], _073270_);
  xor g_101465_(out[404], out[916], _073281_);
  xor g_101466_(out[400], out[912], _073292_);
  and g_101467_(_049444_, out[923], _073303_);
  and g_101468_(out[411], _049796_, _073314_);
  or g_101469_(_073171_, _073215_, _073325_);
  xor g_101470_(out[401], out[913], _073336_);
  or g_101471_(_073226_, _073270_, _073347_);
  or g_101472_(_073325_, _073347_, _073358_);
  or g_101473_(_073193_, _073237_, _073369_);
  or g_101474_(_073182_, _073369_, _073380_);
  or g_101475_(_073358_, _073380_, _073391_);
  or g_101476_(_073204_, _073281_, _073402_);
  or g_101477_(_073391_, _073402_, _073413_);
  xor g_101478_(out[412], out[924], _073424_);
  or g_101479_(_073303_, _073424_, _073435_);
  xor g_101480_(out[407], out[919], _073446_);
  or g_101481_(_073248_, _073446_, _073457_);
  or g_101482_(_073435_, _073457_, _073468_);
  or g_101483_(_073314_, _073336_, _073479_);
  or g_101484_(_073259_, _073479_, _073490_);
  or g_101485_(_073468_, _073490_, _073501_);
  or g_101486_(_073292_, _073501_, _073512_);
  or g_101487_(_073413_, _073512_, _073523_);
  xor g_101488_(out[391], out[919], _073534_);
  and g_101489_(_049433_, out[923], _073545_);
  xor g_101490_(out[398], out[926], _073556_);
  xor g_101491_(out[392], out[920], _073567_);
  xor g_101492_(out[385], out[913], _073578_);
  xor g_101493_(out[397], out[925], _073589_);
  xor g_101494_(out[393], out[921], _073600_);
  xor g_101495_(out[388], out[916], _073611_);
  xor g_101496_(out[386], out[914], _073622_);
  and g_101497_(out[395], _049796_, _073633_);
  xor g_101498_(out[387], out[915], _073644_);
  xor g_101499_(out[390], out[918], _073655_);
  xor g_101500_(out[399], out[927], _073666_);
  xor g_101501_(out[394], out[922], _073677_);
  xor g_101502_(out[389], out[917], _073688_);
  xor g_101503_(out[384], out[912], _073699_);
  or g_101504_(_073556_, _073611_, _073710_);
  or g_101505_(_073567_, _073589_, _073721_);
  or g_101506_(_073622_, _073677_, _073732_);
  or g_101507_(_073721_, _073732_, _073743_);
  or g_101508_(_073600_, _073644_, _073754_);
  or g_101509_(_073688_, _073699_, _073765_);
  or g_101510_(_073754_, _073765_, _073776_);
  or g_101511_(_073743_, _073776_, _073787_);
  xor g_101512_(out[396], out[924], _073798_);
  or g_101513_(_073545_, _073798_, _073809_);
  or g_101514_(_073534_, _073655_, _073820_);
  or g_101515_(_073809_, _073820_, _073831_);
  or g_101516_(_073578_, _073633_, _073842_);
  or g_101517_(_073666_, _073842_, _073853_);
  or g_101518_(_073831_, _073853_, _073864_);
  or g_101519_(_073787_, _073864_, _073875_);
  or g_101520_(_073710_, _073875_, _073886_);
  not g_101521_(_073886_, _073897_);
  and g_101522_(out[379], _049796_, _073908_);
  and g_101523_(_049422_, out[923], _073919_);
  xor g_101524_(out[371], out[915], _073930_);
  xor g_101525_(out[369], out[913], _073941_);
  xor g_101526_(out[382], out[926], _073952_);
  xor g_101527_(out[373], out[917], _073963_);
  xor g_101528_(out[376], out[920], _073974_);
  xor g_101529_(out[378], out[922], _073985_);
  xor g_101530_(out[374], out[918], _073996_);
  xor g_101531_(out[372], out[916], _074007_);
  xor g_101532_(out[381], out[925], _074018_);
  xor g_101533_(out[383], out[927], _074029_);
  xor g_101534_(out[368], out[912], _074040_);
  xor g_101535_(out[370], out[914], _074051_);
  xor g_101536_(out[377], out[921], _074062_);
  or g_101537_(_073952_, _074007_, _074073_);
  or g_101538_(_073974_, _074018_, _074084_);
  or g_101539_(_073985_, _074051_, _074095_);
  or g_101540_(_074084_, _074095_, _074106_);
  or g_101541_(_073930_, _074062_, _074117_);
  or g_101542_(_073963_, _074040_, _074128_);
  or g_101543_(_074117_, _074128_, _074139_);
  or g_101544_(_074106_, _074139_, _074150_);
  xor g_101545_(out[380], out[924], _074161_);
  or g_101546_(_073919_, _074161_, _074172_);
  xor g_101547_(out[375], out[919], _074183_);
  or g_101548_(_073996_, _074183_, _074194_);
  or g_101549_(_074172_, _074194_, _074205_);
  or g_101550_(_073908_, _073941_, _074216_);
  or g_101551_(_074029_, _074216_, _074227_);
  or g_101552_(_074205_, _074227_, _074238_);
  or g_101553_(_074150_, _074238_, _074249_);
  or g_101554_(_074073_, _074249_, _074260_);
  xor g_101555_(out[359], out[919], _074271_);
  and g_101556_(_049411_, out[923], _074282_);
  xor g_101557_(out[366], out[926], _074293_);
  xor g_101558_(out[360], out[920], _074304_);
  xor g_101559_(out[353], out[913], _074315_);
  xor g_101560_(out[365], out[925], _074326_);
  xor g_101561_(out[361], out[921], _074337_);
  xor g_101562_(out[356], out[916], _074348_);
  xor g_101563_(out[354], out[914], _074359_);
  and g_101564_(out[363], _049796_, _074370_);
  xor g_101565_(out[355], out[915], _074381_);
  xor g_101566_(out[358], out[918], _074392_);
  xor g_101567_(out[367], out[927], _074403_);
  xor g_101568_(out[362], out[922], _074414_);
  xor g_101569_(out[357], out[917], _074425_);
  xor g_101570_(out[352], out[912], _074436_);
  or g_101571_(_074293_, _074348_, _074447_);
  or g_101572_(_074304_, _074326_, _074458_);
  or g_101573_(_074359_, _074414_, _074469_);
  or g_101574_(_074458_, _074469_, _074480_);
  or g_101575_(_074337_, _074381_, _074491_);
  or g_101576_(_074425_, _074436_, _074502_);
  or g_101577_(_074491_, _074502_, _074513_);
  or g_101578_(_074480_, _074513_, _074524_);
  xor g_101579_(out[364], out[924], _074535_);
  or g_101580_(_074282_, _074535_, _074546_);
  or g_101581_(_074271_, _074392_, _074557_);
  or g_101582_(_074546_, _074557_, _074568_);
  or g_101583_(_074315_, _074370_, _074579_);
  or g_101584_(_074403_, _074579_, _074590_);
  or g_101585_(_074568_, _074590_, _074601_);
  or g_101586_(_074524_, _074601_, _074612_);
  or g_101587_(_074447_, _074612_, _074623_);
  xor g_101588_(out[337], out[913], _074634_);
  and g_101589_(out[347], _049796_, _074645_);
  xor g_101590_(out[345], out[921], _074656_);
  xor g_101591_(out[336], out[912], _074667_);
  xor g_101592_(out[350], out[926], _074678_);
  xor g_101593_(out[340], out[916], _074689_);
  or g_101594_(_074678_, _074689_, _074700_);
  xor g_101595_(out[349], out[925], _074711_);
  xor g_101596_(out[339], out[915], _074722_);
  and g_101597_(_049400_, out[923], _074733_);
  xor g_101598_(out[342], out[918], _074744_);
  xor g_101599_(out[346], out[922], _074755_);
  xor g_101600_(out[341], out[917], _074766_);
  xor g_101601_(out[351], out[927], _074777_);
  xor g_101602_(out[344], out[920], _074788_);
  or g_101603_(_074711_, _074788_, _074799_);
  xor g_101604_(out[338], out[914], _074810_);
  or g_101605_(_074755_, _074810_, _074821_);
  or g_101606_(_074799_, _074821_, _074832_);
  or g_101607_(_074656_, _074722_, _074843_);
  or g_101608_(_074766_, _074843_, _074854_);
  or g_101609_(_074832_, _074854_, _074865_);
  or g_101610_(_074700_, _074865_, _074876_);
  xor g_101611_(out[348], out[924], _074887_);
  or g_101612_(_074733_, _074887_, _074898_);
  xor g_101613_(out[343], out[919], _074909_);
  or g_101614_(_074744_, _074909_, _074920_);
  or g_101615_(_074898_, _074920_, _074931_);
  or g_101616_(_074634_, _074645_, _074942_);
  or g_101617_(_074777_, _074942_, _074953_);
  or g_101618_(_074931_, _074953_, _074964_);
  or g_101619_(_074667_, _074964_, _074975_);
  or g_101620_(_074876_, _074975_, _074986_);
  xor g_101621_(out[327], out[919], _074997_);
  and g_101622_(_098294_, out[923], _075008_);
  xor g_101623_(out[334], out[926], _075019_);
  xor g_101624_(out[328], out[920], _075030_);
  xor g_101625_(out[321], out[913], _075041_);
  xor g_101626_(out[333], out[925], _075052_);
  xor g_101627_(out[329], out[921], _075063_);
  xor g_101628_(out[324], out[916], _075074_);
  xor g_101629_(out[322], out[914], _075085_);
  and g_101630_(out[331], _049796_, _075096_);
  xor g_101631_(out[323], out[915], _075107_);
  xor g_101632_(out[326], out[918], _075118_);
  xor g_101633_(out[335], out[927], _075129_);
  xor g_101634_(out[330], out[922], _075140_);
  xor g_101635_(out[325], out[917], _075151_);
  xor g_101636_(out[320], out[912], _075162_);
  or g_101637_(_075019_, _075074_, _075173_);
  or g_101638_(_075030_, _075052_, _075184_);
  or g_101639_(_075085_, _075140_, _075195_);
  or g_101640_(_075184_, _075195_, _075206_);
  or g_101641_(_075063_, _075107_, _075217_);
  or g_101642_(_075151_, _075162_, _075228_);
  or g_101643_(_075217_, _075228_, _075239_);
  or g_101644_(_075206_, _075239_, _075250_);
  xor g_101645_(out[332], out[924], _075261_);
  or g_101646_(_075008_, _075261_, _075272_);
  or g_101647_(_074997_, _075118_, _075283_);
  or g_101648_(_075272_, _075283_, _075294_);
  or g_101649_(_075041_, _075096_, _075305_);
  or g_101650_(_075129_, _075305_, _075316_);
  or g_101651_(_075294_, _075316_, _075327_);
  or g_101652_(_075250_, _075327_, _075338_);
  or g_101653_(_075173_, _075338_, _075349_);
  xor g_101654_(out[305], out[913], _075359_);
  and g_101655_(out[315], _049796_, _075370_);
  xor g_101656_(out[313], out[921], _075381_);
  xor g_101657_(out[304], out[912], _075392_);
  xor g_101658_(out[318], out[926], _075403_);
  xor g_101659_(out[308], out[916], _075414_);
  or g_101660_(_075403_, _075414_, _075425_);
  xor g_101661_(out[317], out[925], _075436_);
  xor g_101662_(out[307], out[915], _075447_);
  and g_101663_(_098283_, out[923], _075458_);
  xor g_101664_(out[310], out[918], _075469_);
  xor g_101665_(out[314], out[922], _075480_);
  xor g_101666_(out[309], out[917], _075491_);
  xor g_101667_(out[319], out[927], _075502_);
  xor g_101668_(out[312], out[920], _075513_);
  or g_101669_(_075436_, _075513_, _075524_);
  xor g_101670_(out[306], out[914], _075535_);
  or g_101671_(_075480_, _075535_, _075546_);
  or g_101672_(_075524_, _075546_, _075557_);
  or g_101673_(_075381_, _075447_, _075568_);
  or g_101674_(_075491_, _075568_, _075579_);
  or g_101675_(_075557_, _075579_, _075590_);
  or g_101676_(_075425_, _075590_, _075601_);
  xor g_101677_(out[316], out[924], _075612_);
  or g_101678_(_075458_, _075612_, _075623_);
  xor g_101679_(out[311], out[919], _075634_);
  or g_101680_(_075469_, _075634_, _075645_);
  or g_101681_(_075623_, _075645_, _075656_);
  or g_101682_(_075359_, _075370_, _075667_);
  or g_101683_(_075502_, _075667_, _075678_);
  or g_101684_(_075656_, _075678_, _075689_);
  or g_101685_(_075392_, _075689_, _075700_);
  or g_101686_(_075601_, _075700_, _075711_);
  xor g_101687_(out[295], out[919], _075722_);
  and g_101688_(_098272_, out[923], _075733_);
  xor g_101689_(out[302], out[926], _075744_);
  xor g_101690_(out[296], out[920], _075755_);
  xor g_101691_(out[289], out[913], _075766_);
  xor g_101692_(out[301], out[925], _075777_);
  xor g_101693_(out[297], out[921], _075788_);
  xor g_101694_(out[292], out[916], _075799_);
  xor g_101695_(out[290], out[914], _075810_);
  and g_101696_(out[299], _049796_, _075821_);
  xor g_101697_(out[291], out[915], _075832_);
  xor g_101698_(out[294], out[918], _075843_);
  xor g_101699_(out[303], out[927], _075854_);
  xor g_101700_(out[298], out[922], _075865_);
  xor g_101701_(out[293], out[917], _075876_);
  xor g_101702_(out[288], out[912], _075887_);
  or g_101703_(_075744_, _075799_, _075898_);
  or g_101704_(_075755_, _075777_, _075909_);
  or g_101705_(_075810_, _075865_, _075920_);
  or g_101706_(_075909_, _075920_, _075931_);
  or g_101707_(_075788_, _075832_, _075942_);
  or g_101708_(_075876_, _075887_, _075953_);
  or g_101709_(_075942_, _075953_, _075964_);
  or g_101710_(_075931_, _075964_, _075975_);
  xor g_101711_(out[300], out[924], _075986_);
  or g_101712_(_075733_, _075986_, _075997_);
  or g_101713_(_075722_, _075843_, _076008_);
  or g_101714_(_075997_, _076008_, _076019_);
  or g_101715_(_075766_, _075821_, _076030_);
  or g_101716_(_075854_, _076030_, _076041_);
  or g_101717_(_076019_, _076041_, _076052_);
  or g_101718_(_075975_, _076052_, _076063_);
  or g_101719_(_075898_, _076063_, _076074_);
  not g_101720_(_076074_, _076085_);
  xor g_101721_(out[273], out[913], _076096_);
  and g_101722_(out[283], _049796_, _076107_);
  xor g_101723_(out[281], out[921], _076118_);
  xor g_101724_(out[272], out[912], _076129_);
  xor g_101725_(out[286], out[926], _076140_);
  xor g_101726_(out[276], out[916], _076151_);
  or g_101727_(_076140_, _076151_, _076162_);
  xor g_101728_(out[285], out[925], _076173_);
  xor g_101729_(out[275], out[915], _076184_);
  and g_101730_(_098261_, out[923], _076195_);
  xor g_101731_(out[278], out[918], _076206_);
  xor g_101732_(out[282], out[922], _076217_);
  xor g_101733_(out[277], out[917], _076228_);
  xor g_101734_(out[287], out[927], _076239_);
  xor g_101735_(out[280], out[920], _076250_);
  or g_101736_(_076173_, _076250_, _076261_);
  xor g_101737_(out[274], out[914], _076272_);
  or g_101738_(_076217_, _076272_, _076283_);
  or g_101739_(_076261_, _076283_, _076294_);
  or g_101740_(_076118_, _076184_, _076305_);
  or g_101741_(_076228_, _076305_, _076316_);
  or g_101742_(_076294_, _076316_, _076327_);
  or g_101743_(_076162_, _076327_, _076338_);
  xor g_101744_(out[284], out[924], _076349_);
  or g_101745_(_076195_, _076349_, _076360_);
  xor g_101746_(out[279], out[919], _076371_);
  or g_101747_(_076206_, _076371_, _076382_);
  or g_101748_(_076360_, _076382_, _076393_);
  or g_101749_(_076096_, _076107_, _076404_);
  or g_101750_(_076239_, _076404_, _076415_);
  or g_101751_(_076393_, _076415_, _076426_);
  or g_101752_(_076129_, _076426_, _076437_);
  or g_101753_(_076338_, _076437_, _076448_);
  xor g_101754_(out[263], out[919], _076459_);
  and g_101755_(_098250_, out[923], _076470_);
  xor g_101756_(out[270], out[926], _076481_);
  xor g_101757_(out[264], out[920], _076492_);
  xor g_101758_(out[257], out[913], _076503_);
  xor g_101759_(out[269], out[925], _076514_);
  xor g_101760_(out[265], out[921], _076525_);
  xor g_101761_(out[260], out[916], _076536_);
  xor g_101762_(out[258], out[914], _076547_);
  and g_101763_(out[267], _049796_, _076558_);
  xor g_101764_(out[259], out[915], _076569_);
  xor g_101765_(out[262], out[918], _076580_);
  xor g_101766_(out[271], out[927], _076591_);
  xor g_101767_(out[266], out[922], _076602_);
  xor g_101768_(out[261], out[917], _076613_);
  xor g_101769_(out[256], out[912], _076624_);
  or g_101770_(_076481_, _076536_, _076635_);
  or g_101771_(_076492_, _076514_, _076646_);
  or g_101772_(_076547_, _076602_, _076657_);
  or g_101773_(_076646_, _076657_, _076668_);
  or g_101774_(_076525_, _076569_, _076679_);
  or g_101775_(_076613_, _076624_, _076690_);
  or g_101776_(_076679_, _076690_, _076701_);
  or g_101777_(_076668_, _076701_, _076712_);
  xor g_101778_(out[268], out[924], _076723_);
  or g_101779_(_076470_, _076723_, _076734_);
  or g_101780_(_076459_, _076580_, _076745_);
  or g_101781_(_076734_, _076745_, _076756_);
  or g_101782_(_076503_, _076558_, _076767_);
  or g_101783_(_076591_, _076767_, _076778_);
  or g_101784_(_076756_, _076778_, _076789_);
  or g_101785_(_076712_, _076789_, _076800_);
  or g_101786_(_076635_, _076800_, _076811_);
  xor g_101787_(out[252], out[924], _076822_);
  and g_101788_(_098239_, out[923], _076833_);
  xor g_101789_(out[248], out[920], _076844_);
  xor g_101790_(out[246], out[918], _076855_);
  xor g_101791_(out[253], out[925], _076866_);
  xor g_101792_(out[254], out[926], _076877_);
  xor g_101793_(out[242], out[914], _076888_);
  xor g_101794_(out[249], out[921], _076899_);
  xor g_101795_(out[245], out[917], _076910_);
  xor g_101796_(out[241], out[913], _076921_);
  and g_101797_(out[251], _049796_, _076932_);
  or g_101798_(_076844_, _076866_, _076943_);
  xor g_101799_(out[255], out[927], _076954_);
  xor g_101800_(out[250], out[922], _076965_);
  xor g_101801_(out[244], out[916], _076976_);
  xor g_101802_(out[243], out[915], _076987_);
  xor g_101803_(out[240], out[912], _076998_);
  or g_101804_(_076888_, _076965_, _077009_);
  or g_101805_(_076943_, _077009_, _077020_);
  or g_101806_(_076899_, _076987_, _077031_);
  or g_101807_(_076910_, _077031_, _077042_);
  or g_101808_(_077020_, _077042_, _077053_);
  or g_101809_(_076877_, _076976_, _077064_);
  or g_101810_(_077053_, _077064_, _077075_);
  or g_101811_(_076822_, _076833_, _077086_);
  xor g_101812_(out[247], out[919], _077097_);
  or g_101813_(_076855_, _077097_, _077108_);
  or g_101814_(_077086_, _077108_, _077119_);
  or g_101815_(_076921_, _076932_, _077130_);
  or g_101816_(_076954_, _077130_, _077141_);
  or g_101817_(_077119_, _077141_, _077152_);
  or g_101818_(_076998_, _077152_, _077163_);
  or g_101819_(_077075_, _077163_, _077174_);
  not g_101820_(_077174_, _077185_);
  xor g_101821_(out[231], out[919], _077196_);
  and g_101822_(_098228_, out[923], _077207_);
  xor g_101823_(out[238], out[926], _077218_);
  xor g_101824_(out[232], out[920], _077229_);
  xor g_101825_(out[225], out[913], _077240_);
  xor g_101826_(out[237], out[925], _077251_);
  xor g_101827_(out[233], out[921], _077262_);
  xor g_101828_(out[228], out[916], _077273_);
  xor g_101829_(out[226], out[914], _077284_);
  and g_101830_(out[235], _049796_, _077295_);
  xor g_101831_(out[227], out[915], _077306_);
  xor g_101832_(out[230], out[918], _077317_);
  xor g_101833_(out[239], out[927], _077328_);
  xor g_101834_(out[234], out[922], _077339_);
  xor g_101835_(out[229], out[917], _077350_);
  xor g_101836_(out[224], out[912], _077361_);
  or g_101837_(_077218_, _077273_, _077372_);
  or g_101838_(_077229_, _077251_, _077383_);
  or g_101839_(_077284_, _077339_, _077394_);
  or g_101840_(_077383_, _077394_, _077405_);
  or g_101841_(_077262_, _077306_, _077416_);
  or g_101842_(_077350_, _077361_, _077427_);
  or g_101843_(_077416_, _077427_, _077438_);
  or g_101844_(_077405_, _077438_, _077449_);
  xor g_101845_(out[236], out[924], _077460_);
  or g_101846_(_077207_, _077460_, _077471_);
  or g_101847_(_077196_, _077317_, _077482_);
  or g_101848_(_077471_, _077482_, _077493_);
  or g_101849_(_077240_, _077295_, _077504_);
  or g_101850_(_077328_, _077504_, _077515_);
  or g_101851_(_077493_, _077515_, _077526_);
  or g_101852_(_077449_, _077526_, _077537_);
  or g_101853_(_077372_, _077537_, _077548_);
  not g_101854_(_077548_, _077559_);
  xor g_101855_(out[209], out[913], _077570_);
  and g_101856_(out[219], _049796_, _077581_);
  xor g_101857_(out[217], out[921], _077592_);
  xor g_101858_(out[208], out[912], _077603_);
  xor g_101859_(out[222], out[926], _077614_);
  xor g_101860_(out[212], out[916], _077625_);
  or g_101861_(_077614_, _077625_, _077636_);
  xor g_101862_(out[221], out[925], _077647_);
  xor g_101863_(out[211], out[915], _077658_);
  and g_101864_(_098217_, out[923], _077669_);
  xor g_101865_(out[214], out[918], _077680_);
  xor g_101866_(out[218], out[922], _077691_);
  xor g_101867_(out[213], out[917], _077702_);
  xor g_101868_(out[223], out[927], _077713_);
  xor g_101869_(out[216], out[920], _077724_);
  or g_101870_(_077647_, _077724_, _077735_);
  xor g_101871_(out[210], out[914], _077746_);
  or g_101872_(_077691_, _077746_, _077757_);
  or g_101873_(_077735_, _077757_, _077768_);
  or g_101874_(_077592_, _077658_, _077779_);
  or g_101875_(_077702_, _077779_, _077790_);
  or g_101876_(_077768_, _077790_, _077801_);
  or g_101877_(_077636_, _077801_, _077812_);
  xor g_101878_(out[220], out[924], _077823_);
  or g_101879_(_077669_, _077823_, _077834_);
  xor g_101880_(out[215], out[919], _077845_);
  or g_101881_(_077680_, _077845_, _077856_);
  or g_101882_(_077834_, _077856_, _077867_);
  or g_101883_(_077570_, _077581_, _077878_);
  or g_101884_(_077713_, _077878_, _077889_);
  or g_101885_(_077867_, _077889_, _077900_);
  or g_101886_(_077603_, _077900_, _077911_);
  or g_101887_(_077812_, _077911_, _077922_);
  xor g_101888_(out[199], out[919], _077933_);
  and g_101889_(_098206_, out[923], _077944_);
  xor g_101890_(out[206], out[926], _077955_);
  xor g_101891_(out[200], out[920], _077966_);
  xor g_101892_(out[193], out[913], _077977_);
  xor g_101893_(out[205], out[925], _077988_);
  xor g_101894_(out[201], out[921], _077999_);
  xor g_101895_(out[196], out[916], _078010_);
  xor g_101896_(out[194], out[914], _078021_);
  and g_101897_(out[203], _049796_, _078032_);
  xor g_101898_(out[195], out[915], _078043_);
  xor g_101899_(out[198], out[918], _078054_);
  xor g_101900_(out[207], out[927], _078065_);
  xor g_101901_(out[202], out[922], _078076_);
  xor g_101902_(out[197], out[917], _078087_);
  xor g_101903_(out[192], out[912], _078098_);
  or g_101904_(_077955_, _078010_, _078109_);
  or g_101905_(_077966_, _077988_, _078120_);
  or g_101906_(_078021_, _078076_, _078131_);
  or g_101907_(_078120_, _078131_, _078142_);
  or g_101908_(_077999_, _078043_, _078152_);
  or g_101909_(_078087_, _078098_, _078163_);
  or g_101910_(_078152_, _078163_, _078174_);
  or g_101911_(_078142_, _078174_, _078185_);
  xor g_101912_(out[204], out[924], _078196_);
  or g_101913_(_077944_, _078196_, _078207_);
  or g_101914_(_077933_, _078054_, _078218_);
  or g_101915_(_078207_, _078218_, _078229_);
  or g_101916_(_077977_, _078032_, _078240_);
  or g_101917_(_078065_, _078240_, _078251_);
  or g_101918_(_078229_, _078251_, _078262_);
  or g_101919_(_078185_, _078262_, _078273_);
  or g_101920_(_078109_, _078273_, _078284_);
  xor g_101921_(out[179], out[915], _078295_);
  xor g_101922_(out[180], out[916], _078306_);
  xor g_101923_(out[190], out[926], _078317_);
  xor g_101924_(out[178], out[914], _078328_);
  xor g_101925_(out[181], out[917], _078339_);
  xor g_101926_(out[185], out[921], _078350_);
  xor g_101927_(out[184], out[920], _078361_);
  xor g_101928_(out[191], out[927], _078372_);
  xor g_101929_(out[186], out[922], _078383_);
  xor g_101930_(out[182], out[918], _078394_);
  xor g_101931_(out[176], out[912], _078405_);
  and g_101932_(_098195_, out[923], _078416_);
  and g_101933_(out[187], _049796_, _078427_);
  xor g_101934_(out[189], out[925], _078438_);
  or g_101935_(_078361_, _078438_, _078449_);
  xor g_101936_(out[177], out[913], _078460_);
  or g_101937_(_078328_, _078383_, _078471_);
  or g_101938_(_078449_, _078471_, _078482_);
  or g_101939_(_078295_, _078350_, _078493_);
  or g_101940_(_078339_, _078493_, _078504_);
  or g_101941_(_078482_, _078504_, _078515_);
  or g_101942_(_078306_, _078317_, _078526_);
  or g_101943_(_078515_, _078526_, _078537_);
  xor g_101944_(out[188], out[924], _078548_);
  or g_101945_(_078416_, _078548_, _078559_);
  xor g_101946_(out[183], out[919], _078570_);
  or g_101947_(_078394_, _078570_, _078581_);
  or g_101948_(_078559_, _078581_, _078592_);
  or g_101949_(_078427_, _078460_, _078603_);
  or g_101950_(_078372_, _078603_, _078614_);
  or g_101951_(_078592_, _078614_, _078625_);
  or g_101952_(_078405_, _078625_, _078636_);
  or g_101953_(_078537_, _078636_, _078647_);
  not g_101954_(_078647_, _078658_);
  xor g_101955_(out[167], out[919], _078669_);
  and g_101956_(_098184_, out[923], _078680_);
  xor g_101957_(out[174], out[926], _078691_);
  xor g_101958_(out[168], out[920], _078702_);
  xor g_101959_(out[161], out[913], _078713_);
  xor g_101960_(out[173], out[925], _078724_);
  xor g_101961_(out[169], out[921], _078735_);
  xor g_101962_(out[164], out[916], _078746_);
  xor g_101963_(out[162], out[914], _078757_);
  and g_101964_(out[171], _049796_, _078768_);
  xor g_101965_(out[163], out[915], _078779_);
  xor g_101966_(out[166], out[918], _078790_);
  xor g_101967_(out[175], out[927], _078801_);
  xor g_101968_(out[170], out[922], _078812_);
  xor g_101969_(out[165], out[917], _078823_);
  xor g_101970_(out[160], out[912], _078834_);
  or g_101971_(_078691_, _078746_, _078845_);
  or g_101972_(_078702_, _078724_, _078856_);
  or g_101973_(_078757_, _078812_, _078867_);
  or g_101974_(_078856_, _078867_, _078878_);
  or g_101975_(_078735_, _078779_, _078889_);
  or g_101976_(_078823_, _078834_, _078900_);
  or g_101977_(_078889_, _078900_, _078911_);
  or g_101978_(_078878_, _078911_, _078922_);
  xor g_101979_(out[172], out[924], _078933_);
  or g_101980_(_078680_, _078933_, _078944_);
  or g_101981_(_078669_, _078790_, _078955_);
  or g_101982_(_078944_, _078955_, _078966_);
  or g_101983_(_078713_, _078768_, _078977_);
  or g_101984_(_078801_, _078977_, _078988_);
  or g_101985_(_078966_, _078988_, _078999_);
  or g_101986_(_078922_, _078999_, _079010_);
  or g_101987_(_078845_, _079010_, _079021_);
  not g_101988_(_079021_, _079032_);
  xor g_101989_(out[145], out[913], _079043_);
  and g_101990_(out[155], _049796_, _079054_);
  xor g_101991_(out[158], out[926], _079065_);
  xor g_101992_(out[147], out[915], _079076_);
  xor g_101993_(out[148], out[916], _079087_);
  xor g_101994_(out[146], out[914], _079098_);
  xor g_101995_(out[153], out[921], _079109_);
  xor g_101996_(out[144], out[912], _079120_);
  and g_101997_(_098173_, out[923], _079131_);
  xor g_101998_(out[150], out[918], _079142_);
  xor g_101999_(out[154], out[922], _079153_);
  xor g_102000_(out[149], out[917], _079164_);
  xor g_102001_(out[159], out[927], _079175_);
  xor g_102002_(out[157], out[925], _079186_);
  xor g_102003_(out[152], out[920], _079197_);
  or g_102004_(_079065_, _079087_, _079208_);
  or g_102005_(_079186_, _079197_, _079219_);
  or g_102006_(_079098_, _079153_, _079230_);
  or g_102007_(_079219_, _079230_, _079241_);
  or g_102008_(_079076_, _079109_, _079252_);
  or g_102009_(_079120_, _079164_, _079263_);
  or g_102010_(_079252_, _079263_, _079274_);
  or g_102011_(_079241_, _079274_, _079285_);
  xor g_102012_(out[156], out[924], _079296_);
  or g_102013_(_079131_, _079296_, _079307_);
  xor g_102014_(out[151], out[919], _079318_);
  or g_102015_(_079142_, _079318_, _079329_);
  or g_102016_(_079307_, _079329_, _079340_);
  or g_102017_(_079043_, _079054_, _079351_);
  or g_102018_(_079175_, _079351_, _079362_);
  or g_102019_(_079340_, _079362_, _079373_);
  or g_102020_(_079285_, _079373_, _079384_);
  or g_102021_(_079208_, _079384_, _079395_);
  xor g_102022_(out[135], out[919], _079406_);
  and g_102023_(_098162_, out[923], _079417_);
  xor g_102024_(out[142], out[926], _079428_);
  xor g_102025_(out[136], out[920], _079439_);
  xor g_102026_(out[129], out[913], _079450_);
  xor g_102027_(out[141], out[925], _079461_);
  xor g_102028_(out[137], out[921], _079472_);
  xor g_102029_(out[132], out[916], _079483_);
  xor g_102030_(out[130], out[914], _079494_);
  and g_102031_(out[139], _049796_, _079505_);
  xor g_102032_(out[131], out[915], _079516_);
  xor g_102033_(out[134], out[918], _079527_);
  xor g_102034_(out[143], out[927], _079538_);
  xor g_102035_(out[138], out[922], _079549_);
  xor g_102036_(out[133], out[917], _079560_);
  xor g_102037_(out[128], out[912], _079571_);
  or g_102038_(_079428_, _079483_, _079582_);
  or g_102039_(_079439_, _079461_, _079593_);
  or g_102040_(_079494_, _079549_, _079604_);
  or g_102041_(_079593_, _079604_, _079615_);
  or g_102042_(_079472_, _079516_, _079626_);
  or g_102043_(_079560_, _079571_, _079637_);
  or g_102044_(_079626_, _079637_, _079648_);
  or g_102045_(_079615_, _079648_, _079659_);
  xor g_102046_(out[140], out[924], _079670_);
  or g_102047_(_079417_, _079670_, _079681_);
  or g_102048_(_079406_, _079527_, _079692_);
  or g_102049_(_079681_, _079692_, _079703_);
  or g_102050_(_079450_, _079505_, _079714_);
  or g_102051_(_079538_, _079714_, _079725_);
  or g_102052_(_079703_, _079725_, _079736_);
  or g_102053_(_079659_, _079736_, _079747_);
  or g_102054_(_079582_, _079747_, _079758_);
  xor g_102055_(out[114], out[914], _079769_);
  xor g_102056_(out[112], out[912], _079780_);
  xor g_102057_(out[121], out[921], _079791_);
  xor g_102058_(out[120], out[920], _079802_);
  xor g_102059_(out[117], out[917], _079813_);
  xor g_102060_(out[126], out[926], _079824_);
  xor g_102061_(out[125], out[925], _079835_);
  xor g_102062_(out[127], out[927], _079846_);
  xor g_102063_(out[122], out[922], _079857_);
  xor g_102064_(out[118], out[918], _079868_);
  xor g_102065_(out[115], out[915], _079879_);
  and g_102066_(_098151_, out[923], _079890_);
  and g_102067_(out[123], _049796_, _079901_);
  xor g_102068_(out[116], out[916], _079912_);
  xor g_102069_(out[113], out[913], _079923_);
  or g_102070_(_079824_, _079912_, _079934_);
  or g_102071_(_079802_, _079835_, _079945_);
  or g_102072_(_079769_, _079857_, _079956_);
  or g_102073_(_079945_, _079956_, _079967_);
  or g_102074_(_079791_, _079879_, _079978_);
  or g_102075_(_079780_, _079813_, _079989_);
  or g_102076_(_079978_, _079989_, _080000_);
  or g_102077_(_079967_, _080000_, _080011_);
  xor g_102078_(out[124], out[924], _080022_);
  or g_102079_(_079890_, _080022_, _080033_);
  xor g_102080_(out[119], out[919], _080044_);
  or g_102081_(_079868_, _080044_, _080055_);
  or g_102082_(_080033_, _080055_, _080066_);
  or g_102083_(_079901_, _079923_, _080077_);
  or g_102084_(_079846_, _080077_, _080088_);
  or g_102085_(_080066_, _080088_, _080099_);
  or g_102086_(_080011_, _080099_, _080110_);
  or g_102087_(_079934_, _080110_, _080121_);
  xor g_102088_(out[103], out[919], _080132_);
  and g_102089_(_098140_, out[923], _080143_);
  xor g_102090_(out[110], out[926], _080154_);
  xor g_102091_(out[104], out[920], _080165_);
  xor g_102092_(out[97], out[913], _080176_);
  xor g_102093_(out[109], out[925], _080187_);
  xor g_102094_(out[105], out[921], _080198_);
  xor g_102095_(out[100], out[916], _080209_);
  xor g_102096_(out[98], out[914], _080220_);
  and g_102097_(out[107], _049796_, _080231_);
  xor g_102098_(out[99], out[915], _080242_);
  xor g_102099_(out[102], out[918], _080253_);
  xor g_102100_(out[111], out[927], _080264_);
  xor g_102101_(out[106], out[922], _080275_);
  xor g_102102_(out[101], out[917], _080286_);
  xor g_102103_(out[96], out[912], _080297_);
  or g_102104_(_080154_, _080209_, _080308_);
  or g_102105_(_080165_, _080187_, _080319_);
  or g_102106_(_080220_, _080275_, _080330_);
  or g_102107_(_080319_, _080330_, _080341_);
  or g_102108_(_080198_, _080242_, _080352_);
  or g_102109_(_080286_, _080297_, _080363_);
  or g_102110_(_080352_, _080363_, _080374_);
  or g_102111_(_080341_, _080374_, _080385_);
  xor g_102112_(out[108], out[924], _080396_);
  or g_102113_(_080143_, _080396_, _080407_);
  or g_102114_(_080132_, _080253_, _080418_);
  or g_102115_(_080407_, _080418_, _080429_);
  or g_102116_(_080176_, _080231_, _080440_);
  or g_102117_(_080264_, _080440_, _080451_);
  or g_102118_(_080429_, _080451_, _080462_);
  or g_102119_(_080385_, _080462_, _080473_);
  or g_102120_(_080308_, _080473_, _080484_);
  xor g_102121_(out[92], out[924], _080495_);
  and g_102122_(_098129_, out[923], _080506_);
  xor g_102123_(out[88], out[920], _080517_);
  xor g_102124_(out[86], out[918], _080528_);
  xor g_102125_(out[93], out[925], _080539_);
  xor g_102126_(out[94], out[926], _080550_);
  xor g_102127_(out[82], out[914], _080561_);
  xor g_102128_(out[89], out[921], _080572_);
  xor g_102129_(out[85], out[917], _080583_);
  xor g_102130_(out[81], out[913], _080594_);
  and g_102131_(out[91], _049796_, _080605_);
  or g_102132_(_080517_, _080539_, _080616_);
  xor g_102133_(out[95], out[927], _080627_);
  xor g_102134_(out[90], out[922], _080638_);
  xor g_102135_(out[84], out[916], _080649_);
  xor g_102136_(out[83], out[915], _080660_);
  xor g_102137_(out[80], out[912], _080671_);
  or g_102138_(_080561_, _080638_, _080682_);
  or g_102139_(_080616_, _080682_, _080693_);
  or g_102140_(_080572_, _080660_, _080704_);
  or g_102141_(_080583_, _080704_, _080715_);
  or g_102142_(_080693_, _080715_, _080726_);
  or g_102143_(_080550_, _080649_, _080737_);
  or g_102144_(_080726_, _080737_, _080748_);
  or g_102145_(_080495_, _080506_, _080759_);
  xor g_102146_(out[87], out[919], _080770_);
  or g_102147_(_080528_, _080770_, _080781_);
  or g_102148_(_080759_, _080781_, _080792_);
  or g_102149_(_080594_, _080605_, _080803_);
  or g_102150_(_080627_, _080803_, _080814_);
  or g_102151_(_080792_, _080814_, _080825_);
  or g_102152_(_080671_, _080825_, _080836_);
  or g_102153_(_080748_, _080836_, _080847_);
  not g_102154_(_080847_, _080858_);
  xor g_102155_(out[71], out[919], _080869_);
  and g_102156_(_098118_, out[923], _080880_);
  xor g_102157_(out[78], out[926], _080891_);
  xor g_102158_(out[72], out[920], _080902_);
  xor g_102159_(out[65], out[913], _080913_);
  xor g_102160_(out[77], out[925], _080924_);
  xor g_102161_(out[73], out[921], _080935_);
  xor g_102162_(out[68], out[916], _080945_);
  xor g_102163_(out[66], out[914], _080956_);
  and g_102164_(out[75], _049796_, _080967_);
  xor g_102165_(out[67], out[915], _080978_);
  xor g_102166_(out[70], out[918], _080989_);
  xor g_102167_(out[79], out[927], _081000_);
  xor g_102168_(out[74], out[922], _081011_);
  xor g_102169_(out[69], out[917], _081022_);
  xor g_102170_(out[64], out[912], _081033_);
  or g_102171_(_080891_, _080945_, _081044_);
  or g_102172_(_080902_, _080924_, _081055_);
  or g_102173_(_080956_, _081011_, _081066_);
  or g_102174_(_081055_, _081066_, _081077_);
  or g_102175_(_080935_, _080978_, _081088_);
  or g_102176_(_081022_, _081033_, _081099_);
  or g_102177_(_081088_, _081099_, _081110_);
  or g_102178_(_081077_, _081110_, _081121_);
  xor g_102179_(out[76], out[924], _081132_);
  or g_102180_(_080880_, _081132_, _081143_);
  or g_102181_(_080869_, _080989_, _081154_);
  or g_102182_(_081143_, _081154_, _081165_);
  or g_102183_(_080913_, _080967_, _081176_);
  or g_102184_(_081000_, _081176_, _081187_);
  or g_102185_(_081165_, _081187_, _081198_);
  or g_102186_(_081121_, _081198_, _081209_);
  or g_102187_(_081044_, _081209_, _081220_);
  not g_102188_(_081220_, _081231_);
  xor g_102189_(out[49], out[913], _081242_);
  and g_102190_(out[59], _049796_, _081253_);
  xor g_102191_(out[57], out[921], _081264_);
  xor g_102192_(out[48], out[912], _081275_);
  xor g_102193_(out[62], out[926], _081286_);
  xor g_102194_(out[52], out[916], _081297_);
  or g_102195_(_081286_, _081297_, _081308_);
  xor g_102196_(out[61], out[925], _081319_);
  xor g_102197_(out[51], out[915], _081330_);
  and g_102198_(_098107_, out[923], _081341_);
  xor g_102199_(out[54], out[918], _081352_);
  xor g_102200_(out[58], out[922], _081363_);
  xor g_102201_(out[53], out[917], _081374_);
  xor g_102202_(out[63], out[927], _081385_);
  xor g_102203_(out[56], out[920], _081396_);
  or g_102204_(_081319_, _081396_, _081407_);
  xor g_102205_(out[50], out[914], _081418_);
  or g_102206_(_081363_, _081418_, _081429_);
  or g_102207_(_081407_, _081429_, _081440_);
  or g_102208_(_081264_, _081330_, _081451_);
  or g_102209_(_081374_, _081451_, _081462_);
  or g_102210_(_081440_, _081462_, _081473_);
  or g_102211_(_081308_, _081473_, _081484_);
  xor g_102212_(out[60], out[924], _081495_);
  or g_102213_(_081341_, _081495_, _081506_);
  xor g_102214_(out[55], out[919], _081517_);
  or g_102215_(_081352_, _081517_, _081528_);
  or g_102216_(_081506_, _081528_, _081539_);
  or g_102217_(_081242_, _081253_, _081550_);
  or g_102218_(_081385_, _081550_, _081561_);
  or g_102219_(_081539_, _081561_, _081572_);
  or g_102220_(_081275_, _081572_, _081583_);
  or g_102221_(_081484_, _081583_, _081594_);
  xor g_102222_(out[39], out[919], _081605_);
  and g_102223_(_098096_, out[923], _081616_);
  xor g_102224_(out[46], out[926], _081627_);
  xor g_102225_(out[40], out[920], _081638_);
  xor g_102226_(out[33], out[913], _081649_);
  xor g_102227_(out[45], out[925], _081660_);
  xor g_102228_(out[41], out[921], _081671_);
  xor g_102229_(out[36], out[916], _081682_);
  xor g_102230_(out[34], out[914], _081693_);
  and g_102231_(out[43], _049796_, _081704_);
  xor g_102232_(out[35], out[915], _081715_);
  xor g_102233_(out[38], out[918], _081726_);
  xor g_102234_(out[47], out[927], _081737_);
  xor g_102235_(out[42], out[922], _081748_);
  xor g_102236_(out[37], out[917], _081759_);
  xor g_102237_(out[32], out[912], _081770_);
  or g_102238_(_081627_, _081682_, _081781_);
  or g_102239_(_081638_, _081660_, _081792_);
  or g_102240_(_081693_, _081748_, _081803_);
  or g_102241_(_081792_, _081803_, _081814_);
  or g_102242_(_081671_, _081715_, _081825_);
  or g_102243_(_081759_, _081770_, _081836_);
  or g_102244_(_081825_, _081836_, _081847_);
  or g_102245_(_081814_, _081847_, _081858_);
  xor g_102246_(out[44], out[924], _081869_);
  or g_102247_(_081616_, _081869_, _081880_);
  or g_102248_(_081605_, _081726_, _081891_);
  or g_102249_(_081880_, _081891_, _081902_);
  or g_102250_(_081649_, _081704_, _081913_);
  or g_102251_(_081737_, _081913_, _081924_);
  or g_102252_(_081902_, _081924_, _081935_);
  or g_102253_(_081858_, _081935_, _081946_);
  or g_102254_(_081781_, _081946_, _081957_);
  xor g_102255_(out[17], out[913], _081968_);
  and g_102256_(out[27], _049796_, _081979_);
  xor g_102257_(out[25], out[921], _081990_);
  xor g_102258_(out[16], out[912], _082001_);
  xor g_102259_(out[30], out[926], _082012_);
  xor g_102260_(out[20], out[916], _082023_);
  or g_102261_(_082012_, _082023_, _082034_);
  xor g_102262_(out[29], out[925], _082045_);
  xor g_102263_(out[19], out[915], _082056_);
  and g_102264_(_098063_, out[923], _082067_);
  xor g_102265_(out[22], out[918], _082078_);
  xor g_102266_(out[26], out[922], _082089_);
  xor g_102267_(out[21], out[917], _082100_);
  xor g_102268_(out[31], out[927], _082111_);
  xor g_102269_(out[24], out[920], _082122_);
  or g_102270_(_082045_, _082122_, _082133_);
  xor g_102271_(out[18], out[914], _082144_);
  or g_102272_(_082089_, _082144_, _082155_);
  or g_102273_(_082133_, _082155_, _082166_);
  or g_102274_(_081990_, _082056_, _082177_);
  or g_102275_(_082100_, _082177_, _082188_);
  or g_102276_(_082166_, _082188_, _082199_);
  or g_102277_(_082034_, _082199_, _082210_);
  xor g_102278_(out[28], out[924], _082221_);
  or g_102279_(_082067_, _082221_, _082232_);
  xor g_102280_(out[23], out[919], _082243_);
  or g_102281_(_082078_, _082243_, _082254_);
  or g_102282_(_082232_, _082254_, _082265_);
  or g_102283_(_081968_, _081979_, _082276_);
  or g_102284_(_082111_, _082276_, _082287_);
  or g_102285_(_082265_, _082287_, _082298_);
  or g_102286_(_082001_, _082298_, _082309_);
  or g_102287_(_082210_, _082309_, _082320_);
  not g_102288_(_082320_, _082331_);
  xor g_102289_(out[6], out[918], _082342_);
  xor g_102290_(out[1], out[913], _082353_);
  xor g_102291_(out[0], out[912], _082364_);
  xor g_102292_(out[2], out[914], _082375_);
  xor g_102293_(out[3], out[915], _082386_);
  xor g_102294_(out[9], out[921], _082397_);
  xor g_102295_(out[14], out[926], _082408_);
  and g_102296_(_098041_, out[923], _082419_);
  xor g_102297_(out[7], out[919], _082430_);
  and g_102298_(out[11], _049796_, _082441_);
  xor g_102299_(out[13], out[925], _082452_);
  xor g_102300_(out[8], out[920], _082463_);
  or g_102301_(_082452_, _082463_, _082474_);
  xor g_102302_(out[15], out[927], _082485_);
  xor g_102303_(out[10], out[922], _082496_);
  xor g_102304_(out[5], out[917], _082507_);
  xor g_102305_(out[4], out[916], _082518_);
  or g_102306_(_082375_, _082496_, _082529_);
  or g_102307_(_082474_, _082529_, _082540_);
  or g_102308_(_082386_, _082397_, _082551_);
  or g_102309_(_082507_, _082551_, _082562_);
  or g_102310_(_082540_, _082562_, _082573_);
  or g_102311_(_082408_, _082518_, _082584_);
  or g_102312_(_082573_, _082584_, _082595_);
  xor g_102313_(out[12], out[924], _082606_);
  or g_102314_(_082419_, _082606_, _082617_);
  or g_102315_(_082342_, _082430_, _082628_);
  or g_102316_(_082617_, _082628_, _082639_);
  or g_102317_(_082353_, _082441_, _082650_);
  or g_102318_(_082485_, _082650_, _082661_);
  or g_102319_(_082639_, _082661_, _082672_);
  or g_102320_(_082364_, _082672_, _082683_);
  or g_102321_(_082595_, _082683_, _082694_);
  xor g_102322_(out[471], out[903], _082705_);
  and g_102323_(_049499_, out[907], _082716_);
  xor g_102324_(out[478], out[910], _082727_);
  xor g_102325_(out[472], out[904], _082738_);
  xor g_102326_(out[465], out[897], _082749_);
  xor g_102327_(out[477], out[909], _082760_);
  xor g_102328_(out[473], out[905], _082771_);
  xor g_102329_(out[468], out[900], _082782_);
  xor g_102330_(out[466], out[898], _082793_);
  and g_102331_(out[475], _049785_, _082804_);
  xor g_102332_(out[467], out[899], _082815_);
  xor g_102333_(out[470], out[902], _082826_);
  xor g_102334_(out[479], out[911], _082837_);
  xor g_102335_(out[474], out[906], _082848_);
  xor g_102336_(out[469], out[901], _082859_);
  xor g_102337_(out[464], out[896], _082870_);
  or g_102338_(_082727_, _082782_, _082881_);
  or g_102339_(_082738_, _082760_, _082892_);
  or g_102340_(_082793_, _082848_, _082903_);
  or g_102341_(_082892_, _082903_, _082914_);
  or g_102342_(_082771_, _082815_, _082925_);
  or g_102343_(_082859_, _082870_, _082936_);
  or g_102344_(_082925_, _082936_, _082947_);
  or g_102345_(_082914_, _082947_, _082958_);
  xor g_102346_(out[476], out[908], _082969_);
  or g_102347_(_082716_, _082969_, _082980_);
  or g_102348_(_082705_, _082826_, _082991_);
  or g_102349_(_082980_, _082991_, _083002_);
  or g_102350_(_082749_, _082804_, _083013_);
  or g_102351_(_082837_, _083013_, _083024_);
  or g_102352_(_083002_, _083024_, _083035_);
  or g_102353_(_082958_, _083035_, _083046_);
  or g_102354_(_082881_, _083046_, _083057_);
  xor g_102355_(out[458], out[906], _083068_);
  xor g_102356_(out[456], out[904], _083079_);
  xor g_102357_(out[449], out[897], _083090_);
  and g_102358_(_049477_, out[907], _083101_);
  and g_102359_(out[459], _049785_, _083112_);
  xor g_102360_(out[450], out[898], _083123_);
  xor g_102361_(out[453], out[901], _083134_);
  xor g_102362_(out[457], out[905], _083145_);
  xor g_102363_(out[460], out[908], _083156_);
  xor g_102364_(out[461], out[909], _083167_);
  xor g_102365_(out[463], out[911], _083178_);
  xor g_102366_(out[452], out[900], _083189_);
  xor g_102367_(out[454], out[902], _083200_);
  xor g_102368_(out[451], out[899], _083211_);
  xor g_102369_(out[448], out[896], _083222_);
  xor g_102370_(out[462], out[910], _083233_);
  or g_102371_(_083189_, _083233_, _083244_);
  or g_102372_(_083079_, _083167_, _083255_);
  or g_102373_(_083068_, _083123_, _083266_);
  or g_102374_(_083255_, _083266_, _083277_);
  or g_102375_(_083145_, _083211_, _083288_);
  or g_102376_(_083134_, _083222_, _083299_);
  or g_102377_(_083288_, _083299_, _083310_);
  or g_102378_(_083277_, _083310_, _083321_);
  or g_102379_(_083101_, _083156_, _083332_);
  xor g_102380_(out[455], out[903], _083343_);
  or g_102381_(_083200_, _083343_, _083354_);
  or g_102382_(_083332_, _083354_, _083365_);
  or g_102383_(_083090_, _083112_, _083376_);
  or g_102384_(_083178_, _083376_, _083387_);
  or g_102385_(_083365_, _083387_, _083398_);
  or g_102386_(_083321_, _083398_, _083409_);
  or g_102387_(_083244_, _083409_, _083420_);
  not g_102388_(_083420_, _083431_);
  xor g_102389_(out[439], out[903], _083442_);
  and g_102390_(_049466_, out[907], _083453_);
  xor g_102391_(out[446], out[910], _083464_);
  xor g_102392_(out[440], out[904], _083475_);
  xor g_102393_(out[433], out[897], _083486_);
  xor g_102394_(out[445], out[909], _083497_);
  xor g_102395_(out[441], out[905], _083508_);
  xor g_102396_(out[436], out[900], _083519_);
  xor g_102397_(out[434], out[898], _083530_);
  and g_102398_(out[443], _049785_, _083541_);
  xor g_102399_(out[435], out[899], _083552_);
  xor g_102400_(out[438], out[902], _083563_);
  xor g_102401_(out[447], out[911], _083574_);
  xor g_102402_(out[442], out[906], _083585_);
  xor g_102403_(out[437], out[901], _083596_);
  xor g_102404_(out[432], out[896], _083607_);
  or g_102405_(_083464_, _083519_, _083618_);
  or g_102406_(_083475_, _083497_, _083629_);
  or g_102407_(_083530_, _083585_, _083640_);
  or g_102408_(_083629_, _083640_, _083651_);
  or g_102409_(_083508_, _083552_, _083662_);
  or g_102410_(_083596_, _083607_, _083673_);
  or g_102411_(_083662_, _083673_, _083684_);
  or g_102412_(_083651_, _083684_, _083695_);
  xor g_102413_(out[444], out[908], _083706_);
  or g_102414_(_083453_, _083706_, _083717_);
  or g_102415_(_083442_, _083563_, _083728_);
  or g_102416_(_083717_, _083728_, _083739_);
  or g_102417_(_083486_, _083541_, _083750_);
  or g_102418_(_083574_, _083750_, _083761_);
  or g_102419_(_083739_, _083761_, _083772_);
  or g_102420_(_083695_, _083772_, _083783_);
  or g_102421_(_083618_, _083783_, _083794_);
  xor g_102422_(out[424], out[904], _083805_);
  xor g_102423_(out[421], out[901], _083816_);
  xor g_102424_(out[419], out[899], _083827_);
  xor g_102425_(out[430], out[910], _083838_);
  xor g_102426_(out[429], out[909], _083849_);
  xor g_102427_(out[418], out[898], _083860_);
  xor g_102428_(out[425], out[905], _083871_);
  xor g_102429_(out[422], out[902], _083882_);
  xor g_102430_(out[431], out[911], _083893_);
  xor g_102431_(out[426], out[906], _083904_);
  xor g_102432_(out[420], out[900], _083915_);
  xor g_102433_(out[416], out[896], _083926_);
  and g_102434_(_049455_, out[907], _083936_);
  and g_102435_(out[427], _049785_, _083947_);
  or g_102436_(_083805_, _083849_, _083958_);
  xor g_102437_(out[417], out[897], _083969_);
  or g_102438_(_083860_, _083904_, _083980_);
  or g_102439_(_083958_, _083980_, _083991_);
  or g_102440_(_083827_, _083871_, _084002_);
  or g_102441_(_083816_, _084002_, _084013_);
  or g_102442_(_083991_, _084013_, _084024_);
  or g_102443_(_083838_, _083915_, _084035_);
  or g_102444_(_084024_, _084035_, _084046_);
  xor g_102445_(out[428], out[908], _084057_);
  or g_102446_(_083936_, _084057_, _084068_);
  xor g_102447_(out[423], out[903], _084079_);
  or g_102448_(_083882_, _084079_, _084090_);
  or g_102449_(_084068_, _084090_, _084101_);
  or g_102450_(_083947_, _083969_, _084112_);
  or g_102451_(_083893_, _084112_, _084123_);
  or g_102452_(_084101_, _084123_, _084134_);
  or g_102453_(_083926_, _084134_, _084145_);
  or g_102454_(_084046_, _084145_, _084156_);
  xor g_102455_(out[407], out[903], _084167_);
  and g_102456_(_049444_, out[907], _084178_);
  xor g_102457_(out[414], out[910], _084189_);
  xor g_102458_(out[408], out[904], _084200_);
  xor g_102459_(out[401], out[897], _084211_);
  xor g_102460_(out[413], out[909], _084222_);
  xor g_102461_(out[409], out[905], _084233_);
  xor g_102462_(out[404], out[900], _084244_);
  xor g_102463_(out[402], out[898], _084255_);
  and g_102464_(out[411], _049785_, _084266_);
  xor g_102465_(out[403], out[899], _084277_);
  xor g_102466_(out[406], out[902], _084288_);
  xor g_102467_(out[415], out[911], _084299_);
  xor g_102468_(out[410], out[906], _084310_);
  xor g_102469_(out[405], out[901], _084321_);
  xor g_102470_(out[400], out[896], _084332_);
  or g_102471_(_084189_, _084244_, _084343_);
  or g_102472_(_084200_, _084222_, _084354_);
  or g_102473_(_084255_, _084310_, _084365_);
  or g_102474_(_084354_, _084365_, _084376_);
  or g_102475_(_084233_, _084277_, _084387_);
  or g_102476_(_084321_, _084332_, _084398_);
  or g_102477_(_084387_, _084398_, _084409_);
  or g_102478_(_084376_, _084409_, _084420_);
  xor g_102479_(out[412], out[908], _084431_);
  or g_102480_(_084178_, _084431_, _084442_);
  or g_102481_(_084167_, _084288_, _084453_);
  or g_102482_(_084442_, _084453_, _084464_);
  or g_102483_(_084211_, _084266_, _084475_);
  or g_102484_(_084299_, _084475_, _084486_);
  or g_102485_(_084464_, _084486_, _084497_);
  or g_102486_(_084420_, _084497_, _084508_);
  or g_102487_(_084343_, _084508_, _084519_);
  xor g_102488_(out[394], out[906], _084530_);
  xor g_102489_(out[386], out[898], _084541_);
  xor g_102490_(out[385], out[897], _084552_);
  and g_102491_(_049433_, out[907], _084563_);
  and g_102492_(out[395], _049785_, _084574_);
  xor g_102493_(out[397], out[909], _084585_);
  xor g_102494_(out[387], out[899], _084596_);
  xor g_102495_(out[398], out[910], _084607_);
  xor g_102496_(out[396], out[908], _084618_);
  xor g_102497_(out[392], out[904], _084629_);
  xor g_102498_(out[399], out[911], _084640_);
  xor g_102499_(out[389], out[901], _084651_);
  xor g_102500_(out[390], out[902], _084662_);
  xor g_102501_(out[384], out[896], _084673_);
  xor g_102502_(out[388], out[900], _084684_);
  or g_102503_(_084585_, _084629_, _084695_);
  xor g_102504_(out[393], out[905], _084706_);
  or g_102505_(_084530_, _084541_, _084717_);
  or g_102506_(_084695_, _084717_, _084728_);
  or g_102507_(_084596_, _084706_, _084739_);
  or g_102508_(_084651_, _084739_, _084750_);
  or g_102509_(_084728_, _084750_, _084761_);
  or g_102510_(_084607_, _084684_, _084772_);
  or g_102511_(_084761_, _084772_, _084783_);
  or g_102512_(_084563_, _084618_, _084794_);
  xor g_102513_(out[391], out[903], _084805_);
  or g_102514_(_084662_, _084805_, _084816_);
  or g_102515_(_084794_, _084816_, _084827_);
  or g_102516_(_084552_, _084574_, _084838_);
  or g_102517_(_084640_, _084838_, _084849_);
  or g_102518_(_084827_, _084849_, _084860_);
  or g_102519_(_084673_, _084860_, _084871_);
  or g_102520_(_084783_, _084871_, _084882_);
  xor g_102521_(out[375], out[903], _084893_);
  and g_102522_(_049422_, out[907], _084904_);
  xor g_102523_(out[382], out[910], _084915_);
  xor g_102524_(out[376], out[904], _084926_);
  xor g_102525_(out[369], out[897], _084937_);
  xor g_102526_(out[381], out[909], _084948_);
  xor g_102527_(out[377], out[905], _084959_);
  xor g_102528_(out[372], out[900], _084970_);
  xor g_102529_(out[370], out[898], _084981_);
  and g_102530_(out[379], _049785_, _084992_);
  xor g_102531_(out[371], out[899], _085003_);
  xor g_102532_(out[374], out[902], _085014_);
  xor g_102533_(out[383], out[911], _085025_);
  xor g_102534_(out[378], out[906], _085036_);
  xor g_102535_(out[373], out[901], _085047_);
  xor g_102536_(out[368], out[896], _085058_);
  or g_102537_(_084915_, _084970_, _085069_);
  or g_102538_(_084926_, _084948_, _085080_);
  or g_102539_(_084981_, _085036_, _085091_);
  or g_102540_(_085080_, _085091_, _085102_);
  or g_102541_(_084959_, _085003_, _085113_);
  or g_102542_(_085047_, _085058_, _085124_);
  or g_102543_(_085113_, _085124_, _085135_);
  or g_102544_(_085102_, _085135_, _085146_);
  xor g_102545_(out[380], out[908], _085157_);
  or g_102546_(_084904_, _085157_, _085168_);
  or g_102547_(_084893_, _085014_, _085179_);
  or g_102548_(_085168_, _085179_, _085190_);
  or g_102549_(_084937_, _084992_, _085201_);
  or g_102550_(_085025_, _085201_, _085212_);
  or g_102551_(_085190_, _085212_, _085223_);
  or g_102552_(_085146_, _085223_, _085234_);
  or g_102553_(_085069_, _085234_, _085245_);
  xor g_102554_(out[360], out[904], _085256_);
  xor g_102555_(out[357], out[901], _085267_);
  xor g_102556_(out[355], out[899], _085278_);
  xor g_102557_(out[366], out[910], _085289_);
  xor g_102558_(out[365], out[909], _085300_);
  xor g_102559_(out[354], out[898], _085311_);
  xor g_102560_(out[361], out[905], _085322_);
  xor g_102561_(out[358], out[902], _085333_);
  xor g_102562_(out[367], out[911], _085344_);
  xor g_102563_(out[362], out[906], _085355_);
  xor g_102564_(out[356], out[900], _085366_);
  xor g_102565_(out[352], out[896], _085377_);
  and g_102566_(_049411_, out[907], _085388_);
  and g_102567_(out[363], _049785_, _085399_);
  or g_102568_(_085256_, _085300_, _085410_);
  xor g_102569_(out[353], out[897], _085421_);
  or g_102570_(_085311_, _085355_, _085432_);
  or g_102571_(_085410_, _085432_, _085443_);
  or g_102572_(_085278_, _085322_, _085454_);
  or g_102573_(_085267_, _085454_, _085465_);
  or g_102574_(_085443_, _085465_, _085476_);
  or g_102575_(_085289_, _085366_, _085487_);
  or g_102576_(_085476_, _085487_, _085498_);
  xor g_102577_(out[364], out[908], _085509_);
  or g_102578_(_085388_, _085509_, _085520_);
  xor g_102579_(out[359], out[903], _085531_);
  or g_102580_(_085333_, _085531_, _085542_);
  or g_102581_(_085520_, _085542_, _085553_);
  or g_102582_(_085399_, _085421_, _085564_);
  or g_102583_(_085344_, _085564_, _085575_);
  or g_102584_(_085553_, _085575_, _085586_);
  or g_102585_(_085377_, _085586_, _085597_);
  or g_102586_(_085498_, _085597_, _085608_);
  xor g_102587_(out[343], out[903], _085619_);
  and g_102588_(_049400_, out[907], _085630_);
  xor g_102589_(out[350], out[910], _085641_);
  xor g_102590_(out[344], out[904], _085652_);
  xor g_102591_(out[337], out[897], _085663_);
  xor g_102592_(out[349], out[909], _085674_);
  xor g_102593_(out[345], out[905], _085685_);
  xor g_102594_(out[340], out[900], _085696_);
  xor g_102595_(out[338], out[898], _085707_);
  and g_102596_(out[347], _049785_, _085718_);
  xor g_102597_(out[339], out[899], _085729_);
  xor g_102598_(out[342], out[902], _085740_);
  xor g_102599_(out[351], out[911], _085751_);
  xor g_102600_(out[346], out[906], _085762_);
  xor g_102601_(out[341], out[901], _085773_);
  xor g_102602_(out[336], out[896], _085784_);
  or g_102603_(_085641_, _085696_, _085795_);
  or g_102604_(_085652_, _085674_, _085806_);
  or g_102605_(_085707_, _085762_, _085817_);
  or g_102606_(_085806_, _085817_, _085828_);
  or g_102607_(_085685_, _085729_, _085839_);
  or g_102608_(_085773_, _085784_, _085850_);
  or g_102609_(_085839_, _085850_, _085861_);
  or g_102610_(_085828_, _085861_, _085872_);
  xor g_102611_(out[348], out[908], _085883_);
  or g_102612_(_085630_, _085883_, _085894_);
  or g_102613_(_085619_, _085740_, _085905_);
  or g_102614_(_085894_, _085905_, _085916_);
  or g_102615_(_085663_, _085718_, _085927_);
  or g_102616_(_085751_, _085927_, _085938_);
  or g_102617_(_085916_, _085938_, _085949_);
  or g_102618_(_085872_, _085949_, _085960_);
  or g_102619_(_085795_, _085960_, _085971_);
  not g_102620_(_085971_, _085982_);
  xor g_102621_(out[321], out[897], _085993_);
  and g_102622_(out[331], _049785_, _086004_);
  xor g_102623_(out[329], out[905], _086015_);
  xor g_102624_(out[320], out[896], _086026_);
  xor g_102625_(out[334], out[910], _086037_);
  xor g_102626_(out[324], out[900], _086048_);
  or g_102627_(_086037_, _086048_, _086059_);
  xor g_102628_(out[333], out[909], _086070_);
  xor g_102629_(out[323], out[899], _086081_);
  and g_102630_(_098294_, out[907], _086092_);
  xor g_102631_(out[326], out[902], _086103_);
  xor g_102632_(out[330], out[906], _086114_);
  xor g_102633_(out[325], out[901], _086125_);
  xor g_102634_(out[335], out[911], _086136_);
  xor g_102635_(out[328], out[904], _086147_);
  or g_102636_(_086070_, _086147_, _086158_);
  xor g_102637_(out[322], out[898], _086169_);
  or g_102638_(_086114_, _086169_, _086180_);
  or g_102639_(_086158_, _086180_, _086191_);
  or g_102640_(_086015_, _086081_, _086202_);
  or g_102641_(_086125_, _086202_, _086213_);
  or g_102642_(_086191_, _086213_, _086224_);
  or g_102643_(_086059_, _086224_, _086235_);
  xor g_102644_(out[332], out[908], _086246_);
  or g_102645_(_086092_, _086246_, _086257_);
  xor g_102646_(out[327], out[903], _086268_);
  or g_102647_(_086103_, _086268_, _086279_);
  or g_102648_(_086257_, _086279_, _086290_);
  or g_102649_(_085993_, _086004_, _086301_);
  or g_102650_(_086136_, _086301_, _086312_);
  or g_102651_(_086290_, _086312_, _086323_);
  or g_102652_(_086026_, _086323_, _086334_);
  or g_102653_(_086235_, _086334_, _086345_);
  xor g_102654_(out[311], out[903], _086356_);
  and g_102655_(_098283_, out[907], _086367_);
  xor g_102656_(out[318], out[910], _086378_);
  xor g_102657_(out[312], out[904], _086389_);
  xor g_102658_(out[305], out[897], _086400_);
  xor g_102659_(out[317], out[909], _086411_);
  xor g_102660_(out[313], out[905], _086422_);
  xor g_102661_(out[308], out[900], _086433_);
  xor g_102662_(out[306], out[898], _086444_);
  and g_102663_(out[315], _049785_, _086455_);
  xor g_102664_(out[307], out[899], _086466_);
  xor g_102665_(out[310], out[902], _086477_);
  xor g_102666_(out[319], out[911], _086488_);
  xor g_102667_(out[314], out[906], _086499_);
  xor g_102668_(out[309], out[901], _086510_);
  xor g_102669_(out[304], out[896], _086521_);
  or g_102670_(_086378_, _086433_, _086532_);
  or g_102671_(_086389_, _086411_, _086543_);
  or g_102672_(_086444_, _086499_, _086554_);
  or g_102673_(_086543_, _086554_, _086565_);
  or g_102674_(_086422_, _086466_, _086576_);
  or g_102675_(_086510_, _086521_, _086587_);
  or g_102676_(_086576_, _086587_, _086598_);
  or g_102677_(_086565_, _086598_, _086609_);
  xor g_102678_(out[316], out[908], _086620_);
  or g_102679_(_086367_, _086620_, _086631_);
  or g_102680_(_086356_, _086477_, _086642_);
  or g_102681_(_086631_, _086642_, _086653_);
  or g_102682_(_086400_, _086455_, _086664_);
  or g_102683_(_086488_, _086664_, _086675_);
  or g_102684_(_086653_, _086675_, _086686_);
  or g_102685_(_086609_, _086686_, _086697_);
  or g_102686_(_086532_, _086697_, _086708_);
  xor g_102687_(out[296], out[904], _086719_);
  xor g_102688_(out[293], out[901], _086730_);
  xor g_102689_(out[291], out[899], _086741_);
  xor g_102690_(out[302], out[910], _086752_);
  xor g_102691_(out[301], out[909], _086763_);
  xor g_102692_(out[290], out[898], _086774_);
  xor g_102693_(out[297], out[905], _086785_);
  xor g_102694_(out[294], out[902], _086795_);
  xor g_102695_(out[303], out[911], _086806_);
  xor g_102696_(out[298], out[906], _086817_);
  xor g_102697_(out[292], out[900], _086828_);
  xor g_102698_(out[288], out[896], _086839_);
  and g_102699_(_098272_, out[907], _086850_);
  and g_102700_(out[299], _049785_, _086861_);
  or g_102701_(_086719_, _086763_, _086872_);
  xor g_102702_(out[289], out[897], _086883_);
  or g_102703_(_086774_, _086817_, _086894_);
  or g_102704_(_086872_, _086894_, _086905_);
  or g_102705_(_086741_, _086785_, _086916_);
  or g_102706_(_086730_, _086916_, _086927_);
  or g_102707_(_086905_, _086927_, _086938_);
  or g_102708_(_086752_, _086828_, _086949_);
  or g_102709_(_086938_, _086949_, _086960_);
  xor g_102710_(out[300], out[908], _086971_);
  or g_102711_(_086850_, _086971_, _086982_);
  xor g_102712_(out[295], out[903], _086993_);
  or g_102713_(_086795_, _086993_, _087004_);
  or g_102714_(_086982_, _087004_, _087015_);
  or g_102715_(_086861_, _086883_, _087026_);
  or g_102716_(_086806_, _087026_, _087037_);
  or g_102717_(_087015_, _087037_, _087048_);
  or g_102718_(_086839_, _087048_, _087059_);
  or g_102719_(_086960_, _087059_, _087070_);
  not g_102720_(_087070_, _087081_);
  xor g_102721_(out[279], out[903], _087092_);
  and g_102722_(_098261_, out[907], _087103_);
  xor g_102723_(out[286], out[910], _087114_);
  xor g_102724_(out[280], out[904], _087125_);
  xor g_102725_(out[273], out[897], _087136_);
  xor g_102726_(out[285], out[909], _087147_);
  xor g_102727_(out[281], out[905], _087158_);
  xor g_102728_(out[276], out[900], _087169_);
  xor g_102729_(out[274], out[898], _087180_);
  and g_102730_(out[283], _049785_, _087191_);
  xor g_102731_(out[275], out[899], _087202_);
  xor g_102732_(out[278], out[902], _087213_);
  xor g_102733_(out[287], out[911], _087224_);
  xor g_102734_(out[282], out[906], _087235_);
  xor g_102735_(out[277], out[901], _087246_);
  xor g_102736_(out[272], out[896], _087257_);
  or g_102737_(_087114_, _087169_, _087268_);
  or g_102738_(_087125_, _087147_, _087279_);
  or g_102739_(_087180_, _087235_, _087290_);
  or g_102740_(_087279_, _087290_, _087301_);
  or g_102741_(_087158_, _087202_, _087312_);
  or g_102742_(_087246_, _087257_, _087323_);
  or g_102743_(_087312_, _087323_, _087334_);
  or g_102744_(_087301_, _087334_, _087345_);
  xor g_102745_(out[284], out[908], _087356_);
  or g_102746_(_087103_, _087356_, _087367_);
  or g_102747_(_087092_, _087213_, _087378_);
  or g_102748_(_087367_, _087378_, _087389_);
  or g_102749_(_087136_, _087191_, _087400_);
  or g_102750_(_087224_, _087400_, _087411_);
  or g_102751_(_087389_, _087411_, _087422_);
  or g_102752_(_087345_, _087422_, _087433_);
  or g_102753_(_087268_, _087433_, _087444_);
  not g_102754_(_087444_, _087455_);
  xor g_102755_(out[268], out[908], _087466_);
  and g_102756_(_098250_, out[907], _087477_);
  xor g_102757_(out[264], out[904], _087488_);
  xor g_102758_(out[262], out[902], _087499_);
  xor g_102759_(out[269], out[909], _087510_);
  xor g_102760_(out[270], out[910], _087521_);
  xor g_102761_(out[258], out[898], _087532_);
  xor g_102762_(out[265], out[905], _087543_);
  xor g_102763_(out[261], out[901], _087554_);
  xor g_102764_(out[257], out[897], _087565_);
  and g_102765_(out[267], _049785_, _087576_);
  or g_102766_(_087488_, _087510_, _087587_);
  xor g_102767_(out[271], out[911], _087598_);
  xor g_102768_(out[266], out[906], _087609_);
  xor g_102769_(out[260], out[900], _087620_);
  xor g_102770_(out[259], out[899], _087631_);
  xor g_102771_(out[256], out[896], _087642_);
  or g_102772_(_087532_, _087609_, _087653_);
  or g_102773_(_087587_, _087653_, _087664_);
  or g_102774_(_087543_, _087631_, _087675_);
  or g_102775_(_087554_, _087675_, _087686_);
  or g_102776_(_087664_, _087686_, _087697_);
  or g_102777_(_087521_, _087620_, _087708_);
  or g_102778_(_087697_, _087708_, _087719_);
  or g_102779_(_087466_, _087477_, _087730_);
  xor g_102780_(out[263], out[903], _087741_);
  or g_102781_(_087499_, _087741_, _087752_);
  or g_102782_(_087730_, _087752_, _087763_);
  or g_102783_(_087565_, _087576_, _087774_);
  or g_102784_(_087598_, _087774_, _087785_);
  or g_102785_(_087763_, _087785_, _087796_);
  or g_102786_(_087642_, _087796_, _087807_);
  or g_102787_(_087719_, _087807_, _087818_);
  not g_102788_(_087818_, _087829_);
  xor g_102789_(out[247], out[903], _087840_);
  and g_102790_(_098239_, out[907], _087851_);
  xor g_102791_(out[254], out[910], _087862_);
  xor g_102792_(out[248], out[904], _087873_);
  xor g_102793_(out[241], out[897], _087884_);
  xor g_102794_(out[253], out[909], _087895_);
  xor g_102795_(out[249], out[905], _087906_);
  xor g_102796_(out[244], out[900], _087917_);
  xor g_102797_(out[242], out[898], _087928_);
  and g_102798_(out[251], _049785_, _087939_);
  xor g_102799_(out[243], out[899], _087950_);
  xor g_102800_(out[246], out[902], _087961_);
  xor g_102801_(out[255], out[911], _087972_);
  xor g_102802_(out[250], out[906], _087983_);
  xor g_102803_(out[245], out[901], _087994_);
  xor g_102804_(out[240], out[896], _088005_);
  or g_102805_(_087862_, _087917_, _088016_);
  or g_102806_(_087873_, _087895_, _088027_);
  or g_102807_(_087928_, _087983_, _088038_);
  or g_102808_(_088027_, _088038_, _088049_);
  or g_102809_(_087906_, _087950_, _088060_);
  or g_102810_(_087994_, _088005_, _088071_);
  or g_102811_(_088060_, _088071_, _088082_);
  or g_102812_(_088049_, _088082_, _088093_);
  xor g_102813_(out[252], out[908], _088104_);
  or g_102814_(_087851_, _088104_, _088115_);
  or g_102815_(_087840_, _087961_, _088126_);
  or g_102816_(_088115_, _088126_, _088137_);
  or g_102817_(_087884_, _087939_, _088148_);
  or g_102818_(_087972_, _088148_, _088159_);
  or g_102819_(_088137_, _088159_, _088170_);
  or g_102820_(_088093_, _088170_, _088181_);
  or g_102821_(_088016_, _088181_, _088192_);
  xor g_102822_(out[225], out[897], _088203_);
  and g_102823_(out[235], _049785_, _088214_);
  xor g_102824_(out[233], out[905], _088225_);
  xor g_102825_(out[224], out[896], _088236_);
  xor g_102826_(out[238], out[910], _088247_);
  xor g_102827_(out[228], out[900], _088258_);
  or g_102828_(_088247_, _088258_, _088269_);
  xor g_102829_(out[237], out[909], _088280_);
  xor g_102830_(out[227], out[899], _088291_);
  and g_102831_(_098228_, out[907], _088302_);
  xor g_102832_(out[230], out[902], _088313_);
  xor g_102833_(out[234], out[906], _088324_);
  xor g_102834_(out[229], out[901], _088335_);
  xor g_102835_(out[239], out[911], _088346_);
  xor g_102836_(out[232], out[904], _088357_);
  or g_102837_(_088280_, _088357_, _088368_);
  xor g_102838_(out[226], out[898], _088379_);
  or g_102839_(_088324_, _088379_, _088390_);
  or g_102840_(_088368_, _088390_, _088401_);
  or g_102841_(_088225_, _088291_, _088412_);
  or g_102842_(_088335_, _088412_, _088423_);
  or g_102843_(_088401_, _088423_, _088434_);
  or g_102844_(_088269_, _088434_, _088445_);
  xor g_102845_(out[236], out[908], _088456_);
  or g_102846_(_088302_, _088456_, _088467_);
  xor g_102847_(out[231], out[903], _088478_);
  or g_102848_(_088313_, _088478_, _088489_);
  or g_102849_(_088467_, _088489_, _088500_);
  or g_102850_(_088203_, _088214_, _088511_);
  or g_102851_(_088346_, _088511_, _088522_);
  or g_102852_(_088500_, _088522_, _088533_);
  or g_102853_(_088236_, _088533_, _088544_);
  or g_102854_(_088445_, _088544_, _088555_);
  not g_102855_(_088555_, _088566_);
  xor g_102856_(out[215], out[903], _088577_);
  and g_102857_(_098217_, out[907], _088588_);
  xor g_102858_(out[222], out[910], _088599_);
  xor g_102859_(out[216], out[904], _088610_);
  xor g_102860_(out[209], out[897], _088621_);
  xor g_102861_(out[221], out[909], _088632_);
  xor g_102862_(out[217], out[905], _088643_);
  xor g_102863_(out[212], out[900], _088654_);
  xor g_102864_(out[210], out[898], _088665_);
  and g_102865_(out[219], _049785_, _088676_);
  xor g_102866_(out[211], out[899], _088687_);
  xor g_102867_(out[214], out[902], _088698_);
  xor g_102868_(out[223], out[911], _088709_);
  xor g_102869_(out[218], out[906], _088720_);
  xor g_102870_(out[213], out[901], _088731_);
  xor g_102871_(out[208], out[896], _088742_);
  or g_102872_(_088599_, _088654_, _088753_);
  or g_102873_(_088610_, _088632_, _088764_);
  or g_102874_(_088665_, _088720_, _088775_);
  or g_102875_(_088764_, _088775_, _088786_);
  or g_102876_(_088643_, _088687_, _088797_);
  or g_102877_(_088731_, _088742_, _088808_);
  or g_102878_(_088797_, _088808_, _088819_);
  or g_102879_(_088786_, _088819_, _088830_);
  xor g_102880_(out[220], out[908], _088841_);
  or g_102881_(_088588_, _088841_, _088852_);
  or g_102882_(_088577_, _088698_, _088863_);
  or g_102883_(_088852_, _088863_, _088874_);
  or g_102884_(_088621_, _088676_, _088885_);
  or g_102885_(_088709_, _088885_, _088896_);
  or g_102886_(_088874_, _088896_, _088907_);
  or g_102887_(_088830_, _088907_, _088918_);
  or g_102888_(_088753_, _088918_, _088929_);
  xor g_102889_(out[202], out[906], _088940_);
  xor g_102890_(out[194], out[898], _088951_);
  xor g_102891_(out[193], out[897], _088962_);
  and g_102892_(_098206_, out[907], _088973_);
  and g_102893_(out[203], _049785_, _088984_);
  xor g_102894_(out[205], out[909], _088995_);
  xor g_102895_(out[195], out[899], _089006_);
  xor g_102896_(out[206], out[910], _089017_);
  xor g_102897_(out[204], out[908], _089028_);
  xor g_102898_(out[200], out[904], _089039_);
  xor g_102899_(out[207], out[911], _089050_);
  xor g_102900_(out[197], out[901], _089061_);
  xor g_102901_(out[198], out[902], _089072_);
  xor g_102902_(out[192], out[896], _089083_);
  xor g_102903_(out[196], out[900], _089094_);
  or g_102904_(_088995_, _089039_, _089105_);
  xor g_102905_(out[201], out[905], _089116_);
  or g_102906_(_088940_, _088951_, _089127_);
  or g_102907_(_089105_, _089127_, _089138_);
  or g_102908_(_089006_, _089116_, _089149_);
  or g_102909_(_089061_, _089149_, _089160_);
  or g_102910_(_089138_, _089160_, _089171_);
  or g_102911_(_089017_, _089094_, _089182_);
  or g_102912_(_089171_, _089182_, _089193_);
  or g_102913_(_088973_, _089028_, _089204_);
  xor g_102914_(out[199], out[903], _089215_);
  or g_102915_(_089072_, _089215_, _089226_);
  or g_102916_(_089204_, _089226_, _089237_);
  or g_102917_(_088962_, _088984_, _089248_);
  or g_102918_(_089050_, _089248_, _089259_);
  or g_102919_(_089237_, _089259_, _089270_);
  or g_102920_(_089083_, _089270_, _089281_);
  or g_102921_(_089193_, _089281_, _089292_);
  not g_102922_(_089292_, _089303_);
  xor g_102923_(out[183], out[903], _089314_);
  and g_102924_(_098195_, out[907], _089325_);
  xor g_102925_(out[190], out[910], _089336_);
  xor g_102926_(out[184], out[904], _089347_);
  xor g_102927_(out[177], out[897], _089358_);
  xor g_102928_(out[189], out[909], _089369_);
  xor g_102929_(out[185], out[905], _089380_);
  xor g_102930_(out[180], out[900], _089391_);
  xor g_102931_(out[178], out[898], _089402_);
  and g_102932_(out[187], _049785_, _089413_);
  xor g_102933_(out[179], out[899], _089424_);
  xor g_102934_(out[182], out[902], _089435_);
  xor g_102935_(out[191], out[911], _089446_);
  xor g_102936_(out[186], out[906], _089457_);
  xor g_102937_(out[181], out[901], _089468_);
  xor g_102938_(out[176], out[896], _089479_);
  or g_102939_(_089336_, _089391_, _089490_);
  or g_102940_(_089347_, _089369_, _089501_);
  or g_102941_(_089402_, _089457_, _089512_);
  or g_102942_(_089501_, _089512_, _089523_);
  or g_102943_(_089380_, _089424_, _089534_);
  or g_102944_(_089468_, _089479_, _089545_);
  or g_102945_(_089534_, _089545_, _089556_);
  or g_102946_(_089523_, _089556_, _089567_);
  xor g_102947_(out[188], out[908], _089578_);
  or g_102948_(_089325_, _089578_, _089589_);
  or g_102949_(_089314_, _089435_, _089600_);
  or g_102950_(_089589_, _089600_, _089611_);
  or g_102951_(_089358_, _089413_, _089621_);
  or g_102952_(_089446_, _089621_, _089632_);
  or g_102953_(_089611_, _089632_, _089643_);
  or g_102954_(_089567_, _089643_, _089654_);
  or g_102955_(_089490_, _089654_, _089665_);
  xor g_102956_(out[162], out[898], _089676_);
  xor g_102957_(out[160], out[896], _089687_);
  xor g_102958_(out[169], out[905], _089698_);
  xor g_102959_(out[168], out[904], _089709_);
  xor g_102960_(out[165], out[901], _089720_);
  xor g_102961_(out[174], out[910], _089731_);
  xor g_102962_(out[173], out[909], _089742_);
  xor g_102963_(out[175], out[911], _089753_);
  xor g_102964_(out[170], out[906], _089764_);
  xor g_102965_(out[166], out[902], _089775_);
  xor g_102966_(out[163], out[899], _089786_);
  and g_102967_(_098184_, out[907], _089797_);
  and g_102968_(out[171], _049785_, _089808_);
  xor g_102969_(out[164], out[900], _089819_);
  xor g_102970_(out[161], out[897], _089830_);
  or g_102971_(_089731_, _089819_, _089841_);
  or g_102972_(_089709_, _089742_, _089852_);
  or g_102973_(_089676_, _089764_, _089863_);
  or g_102974_(_089852_, _089863_, _089874_);
  or g_102975_(_089698_, _089786_, _089885_);
  or g_102976_(_089687_, _089720_, _089896_);
  or g_102977_(_089885_, _089896_, _089907_);
  or g_102978_(_089874_, _089907_, _089918_);
  xor g_102979_(out[172], out[908], _089929_);
  or g_102980_(_089797_, _089929_, _089940_);
  xor g_102981_(out[167], out[903], _089951_);
  or g_102982_(_089775_, _089951_, _089962_);
  or g_102983_(_089940_, _089962_, _089973_);
  or g_102984_(_089808_, _089830_, _089984_);
  or g_102985_(_089753_, _089984_, _089995_);
  or g_102986_(_089973_, _089995_, _090006_);
  or g_102987_(_089918_, _090006_, _090017_);
  or g_102988_(_089841_, _090017_, _090028_);
  xor g_102989_(out[151], out[903], _090039_);
  and g_102990_(_098173_, out[907], _090050_);
  xor g_102991_(out[158], out[910], _090061_);
  xor g_102992_(out[152], out[904], _090072_);
  xor g_102993_(out[145], out[897], _090083_);
  xor g_102994_(out[157], out[909], _090094_);
  xor g_102995_(out[153], out[905], _090105_);
  xor g_102996_(out[148], out[900], _090116_);
  xor g_102997_(out[146], out[898], _090127_);
  and g_102998_(out[155], _049785_, _090138_);
  xor g_102999_(out[147], out[899], _090149_);
  xor g_103000_(out[150], out[902], _090160_);
  xor g_103001_(out[159], out[911], _090171_);
  xor g_103002_(out[154], out[906], _090182_);
  xor g_103003_(out[149], out[901], _090193_);
  xor g_103004_(out[144], out[896], _090204_);
  or g_103005_(_090061_, _090116_, _090215_);
  or g_103006_(_090072_, _090094_, _090226_);
  or g_103007_(_090127_, _090182_, _090237_);
  or g_103008_(_090226_, _090237_, _090248_);
  or g_103009_(_090105_, _090149_, _090259_);
  or g_103010_(_090193_, _090204_, _090270_);
  or g_103011_(_090259_, _090270_, _090281_);
  or g_103012_(_090248_, _090281_, _090292_);
  xor g_103013_(out[156], out[908], _090303_);
  or g_103014_(_090050_, _090303_, _090314_);
  or g_103015_(_090039_, _090160_, _090325_);
  or g_103016_(_090314_, _090325_, _090336_);
  or g_103017_(_090083_, _090138_, _090347_);
  or g_103018_(_090171_, _090347_, _090358_);
  or g_103019_(_090336_, _090358_, _090369_);
  or g_103020_(_090292_, _090369_, _090380_);
  or g_103021_(_090215_, _090380_, _090391_);
  not g_103022_(_090391_, _090402_);
  xor g_103023_(out[129], out[897], _090413_);
  and g_103024_(out[139], _049785_, _090424_);
  xor g_103025_(out[137], out[905], _090435_);
  xor g_103026_(out[128], out[896], _090446_);
  xor g_103027_(out[142], out[910], _090457_);
  xor g_103028_(out[132], out[900], _090468_);
  or g_103029_(_090457_, _090468_, _090479_);
  xor g_103030_(out[141], out[909], _090490_);
  xor g_103031_(out[131], out[899], _090501_);
  and g_103032_(_098162_, out[907], _090512_);
  xor g_103033_(out[134], out[902], _090523_);
  xor g_103034_(out[138], out[906], _090534_);
  xor g_103035_(out[133], out[901], _090545_);
  xor g_103036_(out[143], out[911], _090556_);
  xor g_103037_(out[136], out[904], _090567_);
  or g_103038_(_090490_, _090567_, _090578_);
  xor g_103039_(out[130], out[898], _090589_);
  or g_103040_(_090534_, _090589_, _090600_);
  or g_103041_(_090578_, _090600_, _090611_);
  or g_103042_(_090435_, _090501_, _090622_);
  or g_103043_(_090545_, _090622_, _090633_);
  or g_103044_(_090611_, _090633_, _090644_);
  or g_103045_(_090479_, _090644_, _090655_);
  xor g_103046_(out[140], out[908], _090666_);
  or g_103047_(_090512_, _090666_, _090677_);
  xor g_103048_(out[135], out[903], _090688_);
  or g_103049_(_090523_, _090688_, _090699_);
  or g_103050_(_090677_, _090699_, _090710_);
  or g_103051_(_090413_, _090424_, _090721_);
  or g_103052_(_090556_, _090721_, _090732_);
  or g_103053_(_090710_, _090732_, _090743_);
  or g_103054_(_090446_, _090743_, _090754_);
  or g_103055_(_090655_, _090754_, _090765_);
  xor g_103056_(out[119], out[903], _090776_);
  and g_103057_(_098151_, out[907], _090787_);
  xor g_103058_(out[126], out[910], _090798_);
  xor g_103059_(out[120], out[904], _090809_);
  xor g_103060_(out[113], out[897], _090820_);
  xor g_103061_(out[125], out[909], _090831_);
  xor g_103062_(out[121], out[905], _090842_);
  xor g_103063_(out[116], out[900], _090853_);
  xor g_103064_(out[114], out[898], _090864_);
  and g_103065_(out[123], _049785_, _090875_);
  xor g_103066_(out[115], out[899], _090886_);
  xor g_103067_(out[118], out[902], _090897_);
  xor g_103068_(out[127], out[911], _090908_);
  xor g_103069_(out[122], out[906], _090919_);
  xor g_103070_(out[117], out[901], _090930_);
  xor g_103071_(out[112], out[896], _090941_);
  or g_103072_(_090798_, _090853_, _090952_);
  or g_103073_(_090809_, _090831_, _090963_);
  or g_103074_(_090864_, _090919_, _090974_);
  or g_103075_(_090963_, _090974_, _090985_);
  or g_103076_(_090842_, _090886_, _090996_);
  or g_103077_(_090930_, _090941_, _091007_);
  or g_103078_(_090996_, _091007_, _091018_);
  or g_103079_(_090985_, _091018_, _091029_);
  xor g_103080_(out[124], out[908], _091040_);
  or g_103081_(_090787_, _091040_, _091051_);
  or g_103082_(_090776_, _090897_, _091062_);
  or g_103083_(_091051_, _091062_, _091073_);
  or g_103084_(_090820_, _090875_, _091084_);
  or g_103085_(_090908_, _091084_, _091095_);
  or g_103086_(_091073_, _091095_, _091106_);
  or g_103087_(_091029_, _091106_, _091117_);
  or g_103088_(_090952_, _091117_, _091128_);
  xor g_103089_(out[97], out[897], _091139_);
  and g_103090_(out[107], _049785_, _091150_);
  xor g_103091_(out[105], out[905], _091161_);
  xor g_103092_(out[96], out[896], _091172_);
  xor g_103093_(out[110], out[910], _091183_);
  xor g_103094_(out[100], out[900], _091194_);
  or g_103095_(_091183_, _091194_, _091205_);
  xor g_103096_(out[109], out[909], _091216_);
  xor g_103097_(out[99], out[899], _091227_);
  and g_103098_(_098140_, out[907], _091238_);
  xor g_103099_(out[102], out[902], _091249_);
  xor g_103100_(out[106], out[906], _091260_);
  xor g_103101_(out[101], out[901], _091271_);
  xor g_103102_(out[111], out[911], _091282_);
  xor g_103103_(out[104], out[904], _091293_);
  or g_103104_(_091216_, _091293_, _091304_);
  xor g_103105_(out[98], out[898], _091315_);
  or g_103106_(_091260_, _091315_, _091326_);
  or g_103107_(_091304_, _091326_, _091337_);
  or g_103108_(_091161_, _091227_, _091348_);
  or g_103109_(_091271_, _091348_, _091359_);
  or g_103110_(_091337_, _091359_, _091370_);
  or g_103111_(_091205_, _091370_, _091381_);
  xor g_103112_(out[108], out[908], _091392_);
  or g_103113_(_091238_, _091392_, _091403_);
  xor g_103114_(out[103], out[903], _091414_);
  or g_103115_(_091249_, _091414_, _091425_);
  or g_103116_(_091403_, _091425_, _091436_);
  or g_103117_(_091139_, _091150_, _091447_);
  or g_103118_(_091282_, _091447_, _091458_);
  or g_103119_(_091436_, _091458_, _091469_);
  or g_103120_(_091172_, _091469_, _091480_);
  or g_103121_(_091381_, _091480_, _091491_);
  xor g_103122_(out[87], out[903], _091502_);
  and g_103123_(_098129_, out[907], _091513_);
  xor g_103124_(out[94], out[910], _091524_);
  xor g_103125_(out[88], out[904], _091535_);
  xor g_103126_(out[81], out[897], _091546_);
  xor g_103127_(out[93], out[909], _091557_);
  xor g_103128_(out[89], out[905], _091568_);
  xor g_103129_(out[84], out[900], _091579_);
  xor g_103130_(out[82], out[898], _091590_);
  and g_103131_(out[91], _049785_, _091601_);
  xor g_103132_(out[83], out[899], _091612_);
  xor g_103133_(out[86], out[902], _091623_);
  xor g_103134_(out[95], out[911], _091634_);
  xor g_103135_(out[90], out[906], _091645_);
  xor g_103136_(out[85], out[901], _091656_);
  xor g_103137_(out[80], out[896], _091667_);
  or g_103138_(_091524_, _091579_, _091678_);
  or g_103139_(_091535_, _091557_, _091689_);
  or g_103140_(_091590_, _091645_, _091700_);
  or g_103141_(_091689_, _091700_, _091711_);
  or g_103142_(_091568_, _091612_, _091722_);
  or g_103143_(_091656_, _091667_, _091733_);
  or g_103144_(_091722_, _091733_, _091744_);
  or g_103145_(_091711_, _091744_, _091755_);
  xor g_103146_(out[92], out[908], _091766_);
  or g_103147_(_091513_, _091766_, _091777_);
  or g_103148_(_091502_, _091623_, _091788_);
  or g_103149_(_091777_, _091788_, _091799_);
  or g_103150_(_091546_, _091601_, _091810_);
  or g_103151_(_091634_, _091810_, _091821_);
  or g_103152_(_091799_, _091821_, _091832_);
  or g_103153_(_091755_, _091832_, _091843_);
  or g_103154_(_091678_, _091843_, _091854_);
  xor g_103155_(out[65], out[897], _091865_);
  and g_103156_(out[75], _049785_, _091876_);
  xor g_103157_(out[73], out[905], _091887_);
  xor g_103158_(out[64], out[896], _091898_);
  xor g_103159_(out[78], out[910], _091909_);
  xor g_103160_(out[68], out[900], _091920_);
  or g_103161_(_091909_, _091920_, _091931_);
  xor g_103162_(out[77], out[909], _091942_);
  xor g_103163_(out[67], out[899], _091953_);
  and g_103164_(_098118_, out[907], _091964_);
  xor g_103165_(out[70], out[902], _091975_);
  xor g_103166_(out[74], out[906], _091986_);
  xor g_103167_(out[69], out[901], _091997_);
  xor g_103168_(out[79], out[911], _092008_);
  xor g_103169_(out[72], out[904], _092019_);
  or g_103170_(_091942_, _092019_, _092030_);
  xor g_103171_(out[66], out[898], _092041_);
  or g_103172_(_091986_, _092041_, _092052_);
  or g_103173_(_092030_, _092052_, _092063_);
  or g_103174_(_091887_, _091953_, _092074_);
  or g_103175_(_091997_, _092074_, _092085_);
  or g_103176_(_092063_, _092085_, _092096_);
  or g_103177_(_091931_, _092096_, _092107_);
  xor g_103178_(out[76], out[908], _092118_);
  or g_103179_(_091964_, _092118_, _092129_);
  xor g_103180_(out[71], out[903], _092140_);
  or g_103181_(_091975_, _092140_, _092151_);
  or g_103182_(_092129_, _092151_, _092162_);
  or g_103183_(_091865_, _091876_, _092173_);
  or g_103184_(_092008_, _092173_, _092184_);
  or g_103185_(_092162_, _092184_, _092195_);
  or g_103186_(_091898_, _092195_, _092206_);
  or g_103187_(_092107_, _092206_, _092216_);
  xor g_103188_(out[55], out[903], _092227_);
  and g_103189_(_098107_, out[907], _092238_);
  xor g_103190_(out[62], out[910], _092249_);
  xor g_103191_(out[56], out[904], _092260_);
  xor g_103192_(out[49], out[897], _092271_);
  xor g_103193_(out[61], out[909], _092282_);
  xor g_103194_(out[57], out[905], _092293_);
  xor g_103195_(out[52], out[900], _092304_);
  xor g_103196_(out[50], out[898], _092315_);
  and g_103197_(out[59], _049785_, _092326_);
  xor g_103198_(out[51], out[899], _092337_);
  xor g_103199_(out[54], out[902], _092348_);
  xor g_103200_(out[63], out[911], _092359_);
  xor g_103201_(out[58], out[906], _092370_);
  xor g_103202_(out[53], out[901], _092381_);
  xor g_103203_(out[48], out[896], _092392_);
  or g_103204_(_092249_, _092304_, _092403_);
  or g_103205_(_092260_, _092282_, _092414_);
  or g_103206_(_092315_, _092370_, _092425_);
  or g_103207_(_092414_, _092425_, _092436_);
  or g_103208_(_092293_, _092337_, _092447_);
  or g_103209_(_092381_, _092392_, _092458_);
  or g_103210_(_092447_, _092458_, _092469_);
  or g_103211_(_092436_, _092469_, _092480_);
  xor g_103212_(out[60], out[908], _092491_);
  or g_103213_(_092238_, _092491_, _092502_);
  or g_103214_(_092227_, _092348_, _092513_);
  or g_103215_(_092502_, _092513_, _092524_);
  or g_103216_(_092271_, _092326_, _092535_);
  or g_103217_(_092359_, _092535_, _092546_);
  or g_103218_(_092524_, _092546_, _092557_);
  or g_103219_(_092480_, _092557_, _092568_);
  or g_103220_(_092403_, _092568_, _092579_);
  xor g_103221_(out[33], out[897], _092590_);
  and g_103222_(out[43], _049785_, _092601_);
  xor g_103223_(out[46], out[910], _092612_);
  xor g_103224_(out[35], out[899], _092623_);
  xor g_103225_(out[36], out[900], _092634_);
  xor g_103226_(out[34], out[898], _092645_);
  xor g_103227_(out[41], out[905], _092656_);
  xor g_103228_(out[32], out[896], _092667_);
  and g_103229_(_098096_, out[907], _092678_);
  xor g_103230_(out[38], out[902], _092689_);
  xor g_103231_(out[42], out[906], _092700_);
  xor g_103232_(out[37], out[901], _092711_);
  xor g_103233_(out[47], out[911], _092722_);
  xor g_103234_(out[45], out[909], _092733_);
  xor g_103235_(out[40], out[904], _092744_);
  or g_103236_(_092612_, _092634_, _092755_);
  or g_103237_(_092733_, _092744_, _092766_);
  or g_103238_(_092645_, _092700_, _092777_);
  or g_103239_(_092766_, _092777_, _092788_);
  or g_103240_(_092623_, _092656_, _092799_);
  or g_103241_(_092667_, _092711_, _092810_);
  or g_103242_(_092799_, _092810_, _092821_);
  or g_103243_(_092788_, _092821_, _092832_);
  xor g_103244_(out[44], out[908], _092843_);
  or g_103245_(_092678_, _092843_, _092854_);
  xor g_103246_(out[39], out[903], _092865_);
  or g_103247_(_092689_, _092865_, _092876_);
  or g_103248_(_092854_, _092876_, _092887_);
  or g_103249_(_092590_, _092601_, _092898_);
  or g_103250_(_092722_, _092898_, _092909_);
  or g_103251_(_092887_, _092909_, _092920_);
  or g_103252_(_092832_, _092920_, _092931_);
  or g_103253_(_092755_, _092931_, _092942_);
  xor g_103254_(out[23], out[903], _092953_);
  and g_103255_(_098063_, out[907], _092964_);
  xor g_103256_(out[30], out[910], _092975_);
  xor g_103257_(out[24], out[904], _092986_);
  xor g_103258_(out[17], out[897], _092997_);
  xor g_103259_(out[29], out[909], _093008_);
  xor g_103260_(out[25], out[905], _093019_);
  xor g_103261_(out[20], out[900], _093030_);
  xor g_103262_(out[18], out[898], _093041_);
  and g_103263_(out[27], _049785_, _093052_);
  xor g_103264_(out[19], out[899], _093063_);
  xor g_103265_(out[22], out[902], _093074_);
  xor g_103266_(out[31], out[911], _093085_);
  xor g_103267_(out[26], out[906], _093096_);
  xor g_103268_(out[21], out[901], _093107_);
  xor g_103269_(out[16], out[896], _093118_);
  or g_103270_(_092975_, _093030_, _093129_);
  or g_103271_(_092986_, _093008_, _093140_);
  or g_103272_(_093041_, _093096_, _093151_);
  or g_103273_(_093140_, _093151_, _093162_);
  or g_103274_(_093019_, _093063_, _093173_);
  or g_103275_(_093107_, _093118_, _093184_);
  or g_103276_(_093173_, _093184_, _093195_);
  or g_103277_(_093162_, _093195_, _093206_);
  xor g_103278_(out[28], out[908], _093217_);
  or g_103279_(_092964_, _093217_, _093228_);
  or g_103280_(_092953_, _093074_, _093239_);
  or g_103281_(_093228_, _093239_, _093250_);
  or g_103282_(_092997_, _093052_, _093252_);
  or g_103283_(_093085_, _093252_, _093253_);
  or g_103284_(_093250_, _093253_, _093254_);
  or g_103285_(_093206_, _093254_, _093255_);
  or g_103286_(_093129_, _093255_, _093256_);
  xor g_103287_(out[12], out[908], _093257_);
  and g_103288_(_098041_, out[907], _093258_);
  xor g_103289_(out[8], out[904], _093259_);
  xor g_103290_(out[6], out[902], _093260_);
  xor g_103291_(out[13], out[909], _093261_);
  xor g_103292_(out[14], out[910], _093262_);
  xor g_103293_(out[2], out[898], _093263_);
  xor g_103294_(out[9], out[905], _093264_);
  xor g_103295_(out[5], out[901], _093265_);
  xor g_103296_(out[1], out[897], _093266_);
  and g_103297_(out[11], _049785_, _093267_);
  or g_103298_(_093259_, _093261_, _093268_);
  xor g_103299_(out[15], out[911], _093269_);
  xor g_103300_(out[10], out[906], _093270_);
  xor g_103301_(out[4], out[900], _093271_);
  xor g_103302_(out[3], out[899], _093272_);
  xor g_103303_(out[0], out[896], _093273_);
  or g_103304_(_093263_, _093270_, _093274_);
  or g_103305_(_093268_, _093274_, _093275_);
  or g_103306_(_093264_, _093272_, _093276_);
  or g_103307_(_093265_, _093276_, _093277_);
  or g_103308_(_093275_, _093277_, _093278_);
  or g_103309_(_093262_, _093271_, _093279_);
  or g_103310_(_093278_, _093279_, _093280_);
  or g_103311_(_093257_, _093258_, _093281_);
  xor g_103312_(out[7], out[903], _093282_);
  or g_103313_(_093260_, _093282_, _093283_);
  or g_103314_(_093281_, _093283_, _093284_);
  or g_103315_(_093266_, _093267_, _093285_);
  or g_103316_(_093269_, _093285_, _093286_);
  or g_103317_(_093284_, _093286_, _093287_);
  or g_103318_(_093273_, _093287_, _093288_);
  or g_103319_(_093280_, _093288_, _093289_);
  not g_103320_(_093289_, _093290_);
  xor g_103321_(out[472], out[888], _093291_);
  xor g_103322_(out[469], out[885], _093292_);
  xor g_103323_(out[467], out[883], _093293_);
  xor g_103324_(out[478], out[894], _093294_);
  xor g_103325_(out[477], out[893], _093295_);
  xor g_103326_(out[466], out[882], _093296_);
  xor g_103327_(out[473], out[889], _093297_);
  xor g_103328_(out[470], out[886], _093298_);
  xor g_103329_(out[479], out[895], _093299_);
  xor g_103330_(out[474], out[890], _093300_);
  xor g_103331_(out[468], out[884], _093301_);
  xor g_103332_(out[464], out[880], _093302_);
  and g_103333_(_049499_, out[891], _093303_);
  and g_103334_(out[475], _049774_, _093304_);
  or g_103335_(_093291_, _093295_, _093305_);
  xor g_103336_(out[465], out[881], _093306_);
  or g_103337_(_093296_, _093300_, _093307_);
  or g_103338_(_093305_, _093307_, _093308_);
  or g_103339_(_093293_, _093297_, _093309_);
  or g_103340_(_093292_, _093309_, _093310_);
  or g_103341_(_093308_, _093310_, _093311_);
  or g_103342_(_093294_, _093301_, _093312_);
  or g_103343_(_093311_, _093312_, _093313_);
  xor g_103344_(out[476], out[892], _093314_);
  or g_103345_(_093303_, _093314_, _093315_);
  xor g_103346_(out[471], out[887], _093316_);
  or g_103347_(_093298_, _093316_, _093317_);
  or g_103348_(_093315_, _093317_, _093318_);
  or g_103349_(_093304_, _093306_, _093319_);
  or g_103350_(_093299_, _093319_, _093320_);
  or g_103351_(_093318_, _093320_, _093321_);
  or g_103352_(_093302_, _093321_, _093322_);
  or g_103353_(_093313_, _093322_, _093323_);
  not g_103354_(_093323_, _093324_);
  xor g_103355_(out[455], out[887], _093325_);
  and g_103356_(_049477_, out[891], _093326_);
  xor g_103357_(out[462], out[894], _093327_);
  xor g_103358_(out[456], out[888], _093328_);
  xor g_103359_(out[449], out[881], _093329_);
  xor g_103360_(out[461], out[893], _093330_);
  xor g_103361_(out[457], out[889], _093331_);
  xor g_103362_(out[452], out[884], _093332_);
  xor g_103363_(out[450], out[882], _093333_);
  and g_103364_(out[459], _049774_, _093334_);
  xor g_103365_(out[451], out[883], _093335_);
  xor g_103366_(out[454], out[886], _093336_);
  xor g_103367_(out[463], out[895], _093337_);
  xor g_103368_(out[458], out[890], _093338_);
  xor g_103369_(out[453], out[885], _093339_);
  xor g_103370_(out[448], out[880], _093340_);
  or g_103371_(_093327_, _093332_, _093341_);
  or g_103372_(_093328_, _093330_, _093342_);
  or g_103373_(_093333_, _093338_, _093343_);
  or g_103374_(_093342_, _093343_, _093344_);
  or g_103375_(_093331_, _093335_, _093345_);
  or g_103376_(_093339_, _093340_, _093346_);
  or g_103377_(_093345_, _093346_, _093347_);
  or g_103378_(_093344_, _093347_, _093348_);
  xor g_103379_(out[460], out[892], _093349_);
  or g_103380_(_093326_, _093349_, _093350_);
  or g_103381_(_093325_, _093336_, _093351_);
  or g_103382_(_093350_, _093351_, _093352_);
  or g_103383_(_093329_, _093334_, _093353_);
  or g_103384_(_093337_, _093353_, _093354_);
  or g_103385_(_093352_, _093354_, _093355_);
  or g_103386_(_093348_, _093355_, _093356_);
  or g_103387_(_093341_, _093356_, _093357_);
  not g_103388_(_093357_, _093358_);
  xor g_103389_(out[444], out[892], _093359_);
  and g_103390_(_049466_, out[891], _093360_);
  xor g_103391_(out[440], out[888], _093361_);
  xor g_103392_(out[438], out[886], _093362_);
  xor g_103393_(out[445], out[893], _093363_);
  xor g_103394_(out[446], out[894], _093364_);
  xor g_103395_(out[434], out[882], _093365_);
  xor g_103396_(out[441], out[889], _093366_);
  xor g_103397_(out[437], out[885], _093367_);
  xor g_103398_(out[433], out[881], _093368_);
  and g_103399_(out[443], _049774_, _093369_);
  or g_103400_(_093361_, _093363_, _093370_);
  xor g_103401_(out[447], out[895], _093371_);
  xor g_103402_(out[442], out[890], _093372_);
  xor g_103403_(out[436], out[884], _093373_);
  xor g_103404_(out[435], out[883], _093374_);
  xor g_103405_(out[432], out[880], _093375_);
  or g_103406_(_093365_, _093372_, _093376_);
  or g_103407_(_093370_, _093376_, _093377_);
  or g_103408_(_093366_, _093374_, _093378_);
  or g_103409_(_093367_, _093378_, _093379_);
  or g_103410_(_093377_, _093379_, _093380_);
  or g_103411_(_093364_, _093373_, _093381_);
  or g_103412_(_093380_, _093381_, _093382_);
  or g_103413_(_093359_, _093360_, _093383_);
  xor g_103414_(out[439], out[887], _093384_);
  or g_103415_(_093362_, _093384_, _093385_);
  or g_103416_(_093383_, _093385_, _093386_);
  or g_103417_(_093368_, _093369_, _093387_);
  or g_103418_(_093371_, _093387_, _093388_);
  or g_103419_(_093386_, _093388_, _093389_);
  or g_103420_(_093375_, _093389_, _093390_);
  or g_103421_(_093382_, _093390_, _093391_);
  not g_103422_(_093391_, _093392_);
  xor g_103423_(out[423], out[887], _093393_);
  and g_103424_(_049455_, out[891], _093394_);
  xor g_103425_(out[430], out[894], _093395_);
  xor g_103426_(out[424], out[888], _093396_);
  xor g_103427_(out[417], out[881], _093397_);
  xor g_103428_(out[429], out[893], _093398_);
  xor g_103429_(out[425], out[889], _093399_);
  xor g_103430_(out[420], out[884], _093400_);
  xor g_103431_(out[418], out[882], _093401_);
  and g_103432_(out[427], _049774_, _093402_);
  xor g_103433_(out[419], out[883], _093403_);
  xor g_103434_(out[422], out[886], _093404_);
  xor g_103435_(out[431], out[895], _093405_);
  xor g_103436_(out[426], out[890], _093406_);
  xor g_103437_(out[421], out[885], _093407_);
  xor g_103438_(out[416], out[880], _093408_);
  or g_103439_(_093395_, _093400_, _093409_);
  or g_103440_(_093396_, _093398_, _093410_);
  or g_103441_(_093401_, _093406_, _093411_);
  or g_103442_(_093410_, _093411_, _093412_);
  or g_103443_(_093399_, _093403_, _093413_);
  or g_103444_(_093407_, _093408_, _093414_);
  or g_103445_(_093413_, _093414_, _093415_);
  or g_103446_(_093412_, _093415_, _093416_);
  xor g_103447_(out[428], out[892], _093417_);
  or g_103448_(_093394_, _093417_, _093418_);
  or g_103449_(_093393_, _093404_, _093419_);
  or g_103450_(_093418_, _093419_, _093420_);
  or g_103451_(_093397_, _093402_, _093421_);
  or g_103452_(_093405_, _093421_, _093422_);
  or g_103453_(_093420_, _093422_, _093423_);
  or g_103454_(_093416_, _093423_, _093424_);
  or g_103455_(_093409_, _093424_, _093425_);
  xor g_103456_(out[403], out[883], _093426_);
  xor g_103457_(out[404], out[884], _093427_);
  xor g_103458_(out[414], out[894], _093428_);
  xor g_103459_(out[402], out[882], _093429_);
  xor g_103460_(out[405], out[885], _093430_);
  xor g_103461_(out[409], out[889], _093431_);
  xor g_103462_(out[408], out[888], _093432_);
  xor g_103463_(out[415], out[895], _093433_);
  xor g_103464_(out[410], out[890], _093434_);
  xor g_103465_(out[406], out[886], _093435_);
  xor g_103466_(out[400], out[880], _093436_);
  and g_103467_(_049444_, out[891], _093437_);
  and g_103468_(out[411], _049774_, _093438_);
  xor g_103469_(out[413], out[893], _093439_);
  or g_103470_(_093432_, _093439_, _093440_);
  xor g_103471_(out[401], out[881], _093441_);
  or g_103472_(_093429_, _093434_, _093442_);
  or g_103473_(_093440_, _093442_, _093443_);
  or g_103474_(_093426_, _093431_, _093444_);
  or g_103475_(_093430_, _093444_, _093445_);
  or g_103476_(_093443_, _093445_, _093446_);
  or g_103477_(_093427_, _093428_, _093447_);
  or g_103478_(_093446_, _093447_, _093448_);
  xor g_103479_(out[412], out[892], _093449_);
  or g_103480_(_093437_, _093449_, _093450_);
  xor g_103481_(out[407], out[887], _093451_);
  or g_103482_(_093435_, _093451_, _093452_);
  or g_103483_(_093450_, _093452_, _093453_);
  or g_103484_(_093438_, _093441_, _093454_);
  or g_103485_(_093433_, _093454_, _093455_);
  or g_103486_(_093453_, _093455_, _093456_);
  or g_103487_(_093436_, _093456_, _093457_);
  or g_103488_(_093448_, _093457_, _093458_);
  xor g_103489_(out[391], out[887], _093459_);
  and g_103490_(_049433_, out[891], _093460_);
  xor g_103491_(out[398], out[894], _093461_);
  xor g_103492_(out[392], out[888], _093462_);
  xor g_103493_(out[385], out[881], _093463_);
  xor g_103494_(out[397], out[893], _093464_);
  xor g_103495_(out[393], out[889], _093465_);
  xor g_103496_(out[388], out[884], _093466_);
  xor g_103497_(out[386], out[882], _093467_);
  and g_103498_(out[395], _049774_, _093468_);
  xor g_103499_(out[387], out[883], _093469_);
  xor g_103500_(out[390], out[886], _093470_);
  xor g_103501_(out[399], out[895], _093471_);
  xor g_103502_(out[394], out[890], _093472_);
  xor g_103503_(out[389], out[885], _093473_);
  xor g_103504_(out[384], out[880], _093474_);
  or g_103505_(_093461_, _093466_, _093475_);
  or g_103506_(_093462_, _093464_, _093476_);
  or g_103507_(_093467_, _093472_, _093477_);
  or g_103508_(_093476_, _093477_, _093478_);
  or g_103509_(_093465_, _093469_, _093479_);
  or g_103510_(_093473_, _093474_, _093480_);
  or g_103511_(_093479_, _093480_, _093481_);
  or g_103512_(_093478_, _093481_, _093482_);
  xor g_103513_(out[396], out[892], _093483_);
  or g_103514_(_093460_, _093483_, _093484_);
  or g_103515_(_093459_, _093470_, _093485_);
  or g_103516_(_093484_, _093485_, _093486_);
  or g_103517_(_093463_, _093468_, _093487_);
  or g_103518_(_093471_, _093487_, _093488_);
  or g_103519_(_093486_, _093488_, _093489_);
  or g_103520_(_093482_, _093489_, _093490_);
  or g_103521_(_093475_, _093490_, _093491_);
  not g_103522_(_093491_, _093492_);
  xor g_103523_(out[369], out[881], _093493_);
  and g_103524_(out[379], _049774_, _093494_);
  xor g_103525_(out[377], out[889], _093495_);
  xor g_103526_(out[368], out[880], _093496_);
  xor g_103527_(out[382], out[894], _093497_);
  xor g_103528_(out[372], out[884], _093498_);
  or g_103529_(_093497_, _093498_, _093499_);
  xor g_103530_(out[381], out[893], _093500_);
  xor g_103531_(out[371], out[883], _093501_);
  and g_103532_(_049422_, out[891], _093502_);
  xor g_103533_(out[374], out[886], _093503_);
  xor g_103534_(out[378], out[890], _093504_);
  xor g_103535_(out[373], out[885], _093505_);
  xor g_103536_(out[383], out[895], _093506_);
  xor g_103537_(out[376], out[888], _093507_);
  or g_103538_(_093500_, _093507_, _093508_);
  xor g_103539_(out[370], out[882], _093509_);
  or g_103540_(_093504_, _093509_, _093510_);
  or g_103541_(_093508_, _093510_, _093511_);
  or g_103542_(_093495_, _093501_, _093512_);
  or g_103543_(_093505_, _093512_, _093513_);
  or g_103544_(_093511_, _093513_, _093514_);
  or g_103545_(_093499_, _093514_, _093515_);
  xor g_103546_(out[380], out[892], _093516_);
  or g_103547_(_093502_, _093516_, _093517_);
  xor g_103548_(out[375], out[887], _093518_);
  or g_103549_(_093503_, _093518_, _093519_);
  or g_103550_(_093517_, _093519_, _093520_);
  or g_103551_(_093493_, _093494_, _093521_);
  or g_103552_(_093506_, _093521_, _093522_);
  or g_103553_(_093520_, _093522_, _093523_);
  or g_103554_(_093496_, _093523_, _093524_);
  or g_103555_(_093515_, _093524_, _093525_);
  xor g_103556_(out[359], out[887], _093526_);
  and g_103557_(_049411_, out[891], _093527_);
  xor g_103558_(out[366], out[894], _093528_);
  xor g_103559_(out[360], out[888], _093529_);
  xor g_103560_(out[353], out[881], _093530_);
  xor g_103561_(out[365], out[893], _093531_);
  xor g_103562_(out[361], out[889], _093532_);
  xor g_103563_(out[356], out[884], _093533_);
  xor g_103564_(out[354], out[882], _093534_);
  and g_103565_(out[363], _049774_, _093535_);
  xor g_103566_(out[355], out[883], _093536_);
  xor g_103567_(out[358], out[886], _093537_);
  xor g_103568_(out[367], out[895], _093538_);
  xor g_103569_(out[362], out[890], _093539_);
  xor g_103570_(out[357], out[885], _093540_);
  xor g_103571_(out[352], out[880], _093541_);
  or g_103572_(_093528_, _093533_, _093542_);
  or g_103573_(_093529_, _093531_, _093543_);
  or g_103574_(_093534_, _093539_, _093544_);
  or g_103575_(_093543_, _093544_, _093545_);
  or g_103576_(_093532_, _093536_, _093546_);
  or g_103577_(_093540_, _093541_, _093547_);
  or g_103578_(_093546_, _093547_, _093548_);
  or g_103579_(_093545_, _093548_, _093549_);
  xor g_103580_(out[364], out[892], _093550_);
  or g_103581_(_093527_, _093550_, _093551_);
  or g_103582_(_093526_, _093537_, _093552_);
  or g_103583_(_093551_, _093552_, _093553_);
  or g_103584_(_093530_, _093535_, _093554_);
  or g_103585_(_093538_, _093554_, _093555_);
  or g_103586_(_093553_, _093555_, _093556_);
  or g_103587_(_093549_, _093556_, _093557_);
  or g_103588_(_093542_, _093557_, _093558_);
  xor g_103589_(out[337], out[881], _093559_);
  and g_103590_(out[347], _049774_, _093560_);
  xor g_103591_(out[345], out[889], _093561_);
  xor g_103592_(out[336], out[880], _093562_);
  xor g_103593_(out[350], out[894], _093563_);
  xor g_103594_(out[340], out[884], _093564_);
  or g_103595_(_093563_, _093564_, _093565_);
  xor g_103596_(out[349], out[893], _093566_);
  xor g_103597_(out[339], out[883], _093567_);
  and g_103598_(_049400_, out[891], _093568_);
  xor g_103599_(out[342], out[886], _093569_);
  xor g_103600_(out[346], out[890], _093570_);
  xor g_103601_(out[341], out[885], _093571_);
  xor g_103602_(out[351], out[895], _093572_);
  xor g_103603_(out[344], out[888], _093573_);
  or g_103604_(_093566_, _093573_, _093574_);
  xor g_103605_(out[338], out[882], _093575_);
  or g_103606_(_093570_, _093575_, _093576_);
  or g_103607_(_093574_, _093576_, _093577_);
  or g_103608_(_093561_, _093567_, _093578_);
  or g_103609_(_093571_, _093578_, _093579_);
  or g_103610_(_093577_, _093579_, _093580_);
  or g_103611_(_093565_, _093580_, _093581_);
  xor g_103612_(out[348], out[892], _093582_);
  or g_103613_(_093568_, _093582_, _093583_);
  xor g_103614_(out[343], out[887], _093584_);
  or g_103615_(_093569_, _093584_, _093585_);
  or g_103616_(_093583_, _093585_, _093586_);
  or g_103617_(_093559_, _093560_, _093587_);
  or g_103618_(_093572_, _093587_, _093588_);
  or g_103619_(_093586_, _093588_, _093589_);
  or g_103620_(_093562_, _093589_, _093590_);
  or g_103621_(_093581_, _093590_, _093591_);
  xor g_103622_(out[327], out[887], _093592_);
  and g_103623_(_098294_, out[891], _093593_);
  xor g_103624_(out[334], out[894], _093594_);
  xor g_103625_(out[328], out[888], _093595_);
  xor g_103626_(out[321], out[881], _093596_);
  xor g_103627_(out[333], out[893], _093597_);
  xor g_103628_(out[329], out[889], _093598_);
  xor g_103629_(out[324], out[884], _093599_);
  xor g_103630_(out[322], out[882], _093600_);
  and g_103631_(out[331], _049774_, _093601_);
  xor g_103632_(out[323], out[883], _093602_);
  xor g_103633_(out[326], out[886], _093603_);
  xor g_103634_(out[335], out[895], _093604_);
  xor g_103635_(out[330], out[890], _093605_);
  xor g_103636_(out[325], out[885], _093606_);
  xor g_103637_(out[320], out[880], _093607_);
  or g_103638_(_093594_, _093599_, _093608_);
  or g_103639_(_093595_, _093597_, _093609_);
  or g_103640_(_093600_, _093605_, _093610_);
  or g_103641_(_093609_, _093610_, _093611_);
  or g_103642_(_093598_, _093602_, _093612_);
  or g_103643_(_093606_, _093607_, _093613_);
  or g_103644_(_093612_, _093613_, _093614_);
  or g_103645_(_093611_, _093614_, _093615_);
  xor g_103646_(out[332], out[892], _093616_);
  or g_103647_(_093593_, _093616_, _093617_);
  or g_103648_(_093592_, _093603_, _093618_);
  or g_103649_(_093617_, _093618_, _093619_);
  or g_103650_(_093596_, _093601_, _093620_);
  or g_103651_(_093604_, _093620_, _093621_);
  or g_103652_(_093619_, _093621_, _093622_);
  or g_103653_(_093615_, _093622_, _093623_);
  or g_103654_(_093608_, _093623_, _093624_);
  xor g_103655_(out[316], out[892], _093625_);
  and g_103656_(_098283_, out[891], _093626_);
  xor g_103657_(out[317], out[893], _093627_);
  xor g_103658_(out[310], out[886], _093628_);
  xor g_103659_(out[312], out[888], _093629_);
  xor g_103660_(out[313], out[889], _093630_);
  xor g_103661_(out[318], out[894], _093631_);
  xor g_103662_(out[308], out[884], _093632_);
  or g_103663_(_093631_, _093632_, _093633_);
  xor g_103664_(out[309], out[885], _093634_);
  xor g_103665_(out[305], out[881], _093635_);
  and g_103666_(out[315], _049774_, _093636_);
  xor g_103667_(out[319], out[895], _093637_);
  xor g_103668_(out[314], out[890], _093638_);
  xor g_103669_(out[304], out[880], _093639_);
  xor g_103670_(out[306], out[882], _093640_);
  xor g_103671_(out[307], out[883], _093641_);
  or g_103672_(_093627_, _093629_, _093642_);
  or g_103673_(_093638_, _093640_, _093643_);
  or g_103674_(_093642_, _093643_, _093644_);
  or g_103675_(_093630_, _093641_, _093645_);
  or g_103676_(_093634_, _093639_, _093646_);
  or g_103677_(_093645_, _093646_, _093647_);
  or g_103678_(_093644_, _093647_, _093648_);
  or g_103679_(_093625_, _093626_, _093649_);
  xor g_103680_(out[311], out[887], _093650_);
  or g_103681_(_093628_, _093650_, _093651_);
  or g_103682_(_093649_, _093651_, _093652_);
  or g_103683_(_093635_, _093636_, _093653_);
  or g_103684_(_093637_, _093653_, _093654_);
  or g_103685_(_093652_, _093654_, _093655_);
  or g_103686_(_093648_, _093655_, _093656_);
  or g_103687_(_093633_, _093656_, _093657_);
  not g_103688_(_093657_, _093658_);
  xor g_103689_(out[295], out[887], _093659_);
  and g_103690_(_098272_, out[891], _093660_);
  xor g_103691_(out[302], out[894], _093661_);
  xor g_103692_(out[296], out[888], _093662_);
  xor g_103693_(out[289], out[881], _093663_);
  xor g_103694_(out[301], out[893], _093664_);
  xor g_103695_(out[297], out[889], _093665_);
  xor g_103696_(out[292], out[884], _093666_);
  xor g_103697_(out[290], out[882], _093667_);
  and g_103698_(out[299], _049774_, _093668_);
  xor g_103699_(out[291], out[883], _093669_);
  xor g_103700_(out[294], out[886], _093670_);
  xor g_103701_(out[303], out[895], _093671_);
  xor g_103702_(out[298], out[890], _093672_);
  xor g_103703_(out[293], out[885], _093673_);
  xor g_103704_(out[288], out[880], _093674_);
  or g_103705_(_093661_, _093666_, _093675_);
  or g_103706_(_093662_, _093664_, _093676_);
  or g_103707_(_093667_, _093672_, _093677_);
  or g_103708_(_093676_, _093677_, _093678_);
  or g_103709_(_093665_, _093669_, _093679_);
  or g_103710_(_093673_, _093674_, _093680_);
  or g_103711_(_093679_, _093680_, _093681_);
  or g_103712_(_093678_, _093681_, _093682_);
  xor g_103713_(out[300], out[892], _093683_);
  or g_103714_(_093660_, _093683_, _093684_);
  or g_103715_(_093659_, _093670_, _093685_);
  or g_103716_(_093684_, _093685_, _093686_);
  or g_103717_(_093663_, _093668_, _093687_);
  or g_103718_(_093671_, _093687_, _093688_);
  or g_103719_(_093686_, _093688_, _093689_);
  or g_103720_(_093682_, _093689_, _093690_);
  or g_103721_(_093675_, _093690_, _093691_);
  xor g_103722_(out[273], out[881], _093692_);
  and g_103723_(out[283], _049774_, _093693_);
  xor g_103724_(out[281], out[889], _093694_);
  xor g_103725_(out[272], out[880], _093695_);
  xor g_103726_(out[286], out[894], _093696_);
  xor g_103727_(out[276], out[884], _093697_);
  or g_103728_(_093696_, _093697_, _093698_);
  xor g_103729_(out[285], out[893], _093699_);
  xor g_103730_(out[275], out[883], _093700_);
  and g_103731_(_098261_, out[891], _093701_);
  xor g_103732_(out[278], out[886], _093702_);
  xor g_103733_(out[282], out[890], _093703_);
  xor g_103734_(out[277], out[885], _093704_);
  xor g_103735_(out[287], out[895], _093705_);
  xor g_103736_(out[280], out[888], _093706_);
  or g_103737_(_093699_, _093706_, _093707_);
  xor g_103738_(out[274], out[882], _093708_);
  or g_103739_(_093703_, _093708_, _093709_);
  or g_103740_(_093707_, _093709_, _093710_);
  or g_103741_(_093694_, _093700_, _093711_);
  or g_103742_(_093704_, _093711_, _093712_);
  or g_103743_(_093710_, _093712_, _093713_);
  or g_103744_(_093698_, _093713_, _093714_);
  xor g_103745_(out[284], out[892], _093715_);
  or g_103746_(_093701_, _093715_, _093716_);
  xor g_103747_(out[279], out[887], _093717_);
  or g_103748_(_093702_, _093717_, _093718_);
  or g_103749_(_093716_, _093718_, _093719_);
  or g_103750_(_093692_, _093693_, _093720_);
  or g_103751_(_093705_, _093720_, _093721_);
  or g_103752_(_093719_, _093721_, _093722_);
  or g_103753_(_093695_, _093722_, _093723_);
  or g_103754_(_093714_, _093723_, _093724_);
  xor g_103755_(out[263], out[887], _093725_);
  and g_103756_(_098250_, out[891], _093726_);
  xor g_103757_(out[270], out[894], _093727_);
  xor g_103758_(out[264], out[888], _093728_);
  xor g_103759_(out[257], out[881], _093729_);
  xor g_103760_(out[269], out[893], _093730_);
  xor g_103761_(out[265], out[889], _093731_);
  xor g_103762_(out[260], out[884], _093732_);
  xor g_103763_(out[258], out[882], _093733_);
  and g_103764_(out[267], _049774_, _093734_);
  xor g_103765_(out[259], out[883], _093735_);
  xor g_103766_(out[262], out[886], _093736_);
  xor g_103767_(out[271], out[895], _093737_);
  xor g_103768_(out[266], out[890], _093738_);
  xor g_103769_(out[261], out[885], _093739_);
  xor g_103770_(out[256], out[880], _093740_);
  or g_103771_(_093727_, _093732_, _093741_);
  or g_103772_(_093728_, _093730_, _093742_);
  or g_103773_(_093733_, _093738_, _093743_);
  or g_103774_(_093742_, _093743_, _093744_);
  or g_103775_(_093731_, _093735_, _093745_);
  or g_103776_(_093739_, _093740_, _093746_);
  or g_103777_(_093745_, _093746_, _093747_);
  or g_103778_(_093744_, _093747_, _093748_);
  xor g_103779_(out[268], out[892], _093749_);
  or g_103780_(_093726_, _093749_, _093750_);
  or g_103781_(_093725_, _093736_, _093751_);
  or g_103782_(_093750_, _093751_, _093752_);
  or g_103783_(_093729_, _093734_, _093753_);
  or g_103784_(_093737_, _093753_, _093754_);
  or g_103785_(_093752_, _093754_, _093755_);
  or g_103786_(_093748_, _093755_, _093756_);
  or g_103787_(_093741_, _093756_, _093757_);
  and g_103788_(out[251], _049774_, _093758_);
  xor g_103789_(out[244], out[884], _093759_);
  xor g_103790_(out[254], out[894], _093760_);
  or g_103791_(_093759_, _093760_, _093761_);
  xor g_103792_(out[253], out[893], _093762_);
  xor g_103793_(out[243], out[883], _093763_);
  xor g_103794_(out[240], out[880], _093764_);
  and g_103795_(_098239_, out[891], _093765_);
  xor g_103796_(out[250], out[890], _093766_);
  xor g_103797_(out[255], out[895], _093767_);
  xor g_103798_(out[246], out[886], _093768_);
  xor g_103799_(out[245], out[885], _093769_);
  xor g_103800_(out[248], out[888], _093770_);
  or g_103801_(_093762_, _093770_, _093771_);
  xor g_103802_(out[242], out[882], _093772_);
  xor g_103803_(out[249], out[889], _093773_);
  xor g_103804_(out[241], out[881], _093774_);
  or g_103805_(_093766_, _093772_, _093775_);
  or g_103806_(_093771_, _093775_, _093776_);
  or g_103807_(_093763_, _093773_, _093777_);
  or g_103808_(_093769_, _093777_, _093778_);
  or g_103809_(_093776_, _093778_, _093779_);
  or g_103810_(_093761_, _093779_, _093780_);
  xor g_103811_(out[252], out[892], _093781_);
  or g_103812_(_093765_, _093781_, _093782_);
  xor g_103813_(out[247], out[887], _093783_);
  or g_103814_(_093768_, _093783_, _093784_);
  or g_103815_(_093782_, _093784_, _093785_);
  or g_103816_(_093758_, _093774_, _093786_);
  or g_103817_(_093767_, _093786_, _093787_);
  or g_103818_(_093785_, _093787_, _093788_);
  or g_103819_(_093764_, _093788_, _093789_);
  or g_103820_(_093780_, _093789_, _093790_);
  xor g_103821_(out[231], out[887], _093791_);
  and g_103822_(_098228_, out[891], _093792_);
  xor g_103823_(out[238], out[894], _093793_);
  xor g_103824_(out[232], out[888], _093794_);
  xor g_103825_(out[225], out[881], _093795_);
  xor g_103826_(out[237], out[893], _093796_);
  xor g_103827_(out[233], out[889], _093797_);
  xor g_103828_(out[228], out[884], _093798_);
  xor g_103829_(out[226], out[882], _093799_);
  and g_103830_(out[235], _049774_, _093800_);
  xor g_103831_(out[227], out[883], _093801_);
  xor g_103832_(out[230], out[886], _093802_);
  xor g_103833_(out[239], out[895], _093803_);
  xor g_103834_(out[234], out[890], _093804_);
  xor g_103835_(out[229], out[885], _093805_);
  xor g_103836_(out[224], out[880], _093806_);
  or g_103837_(_093793_, _093798_, _093807_);
  or g_103838_(_093794_, _093796_, _093808_);
  or g_103839_(_093799_, _093804_, _093809_);
  or g_103840_(_093808_, _093809_, _093810_);
  or g_103841_(_093797_, _093801_, _093811_);
  or g_103842_(_093805_, _093806_, _093812_);
  or g_103843_(_093811_, _093812_, _093813_);
  or g_103844_(_093810_, _093813_, _093814_);
  xor g_103845_(out[236], out[892], _093815_);
  or g_103846_(_093792_, _093815_, _093816_);
  or g_103847_(_093791_, _093802_, _093817_);
  or g_103848_(_093816_, _093817_, _093818_);
  or g_103849_(_093795_, _093800_, _093819_);
  or g_103850_(_093803_, _093819_, _093820_);
  or g_103851_(_093818_, _093820_, _093821_);
  or g_103852_(_093814_, _093821_, _093822_);
  or g_103853_(_093807_, _093822_, _093823_);
  and g_103854_(out[219], _049774_, _093824_);
  xor g_103855_(out[212], out[884], _093825_);
  xor g_103856_(out[222], out[894], _093826_);
  or g_103857_(_093825_, _093826_, _093827_);
  xor g_103858_(out[221], out[893], _093828_);
  xor g_103859_(out[211], out[883], _093829_);
  xor g_103860_(out[208], out[880], _093830_);
  and g_103861_(_098217_, out[891], _093831_);
  xor g_103862_(out[218], out[890], _093832_);
  xor g_103863_(out[223], out[895], _093833_);
  xor g_103864_(out[214], out[886], _093834_);
  xor g_103865_(out[213], out[885], _093835_);
  xor g_103866_(out[216], out[888], _093836_);
  or g_103867_(_093828_, _093836_, _093837_);
  xor g_103868_(out[210], out[882], _093838_);
  xor g_103869_(out[217], out[889], _093839_);
  xor g_103870_(out[209], out[881], _093840_);
  or g_103871_(_093832_, _093838_, _093841_);
  or g_103872_(_093837_, _093841_, _093842_);
  or g_103873_(_093829_, _093839_, _093843_);
  or g_103874_(_093835_, _093843_, _093844_);
  or g_103875_(_093842_, _093844_, _093845_);
  or g_103876_(_093827_, _093845_, _093846_);
  xor g_103877_(out[220], out[892], _093847_);
  or g_103878_(_093831_, _093847_, _093848_);
  xor g_103879_(out[215], out[887], _093849_);
  or g_103880_(_093834_, _093849_, _093850_);
  or g_103881_(_093848_, _093850_, _093851_);
  or g_103882_(_093824_, _093840_, _093852_);
  or g_103883_(_093833_, _093852_, _093853_);
  or g_103884_(_093851_, _093853_, _093854_);
  or g_103885_(_093830_, _093854_, _093855_);
  or g_103886_(_093846_, _093855_, _093856_);
  xor g_103887_(out[199], out[887], _093857_);
  and g_103888_(_098206_, out[891], _093858_);
  xor g_103889_(out[206], out[894], _093859_);
  xor g_103890_(out[200], out[888], _093860_);
  xor g_103891_(out[193], out[881], _093861_);
  xor g_103892_(out[205], out[893], _093862_);
  xor g_103893_(out[201], out[889], _093863_);
  xor g_103894_(out[196], out[884], _093864_);
  xor g_103895_(out[194], out[882], _093865_);
  and g_103896_(out[203], _049774_, _093866_);
  xor g_103897_(out[195], out[883], _093867_);
  xor g_103898_(out[198], out[886], _093868_);
  xor g_103899_(out[207], out[895], _093869_);
  xor g_103900_(out[202], out[890], _093870_);
  xor g_103901_(out[197], out[885], _093871_);
  xor g_103902_(out[192], out[880], _093872_);
  or g_103903_(_093859_, _093864_, _093873_);
  or g_103904_(_093860_, _093862_, _093874_);
  or g_103905_(_093865_, _093870_, _093875_);
  or g_103906_(_093874_, _093875_, _093876_);
  or g_103907_(_093863_, _093867_, _093877_);
  or g_103908_(_093871_, _093872_, _093878_);
  or g_103909_(_093877_, _093878_, _093879_);
  or g_103910_(_093876_, _093879_, _093880_);
  xor g_103911_(out[204], out[892], _093881_);
  or g_103912_(_093858_, _093881_, _093882_);
  or g_103913_(_093857_, _093868_, _093883_);
  or g_103914_(_093882_, _093883_, _093884_);
  or g_103915_(_093861_, _093866_, _093885_);
  or g_103916_(_093869_, _093885_, _093886_);
  or g_103917_(_093884_, _093886_, _093887_);
  or g_103918_(_093880_, _093887_, _093888_);
  or g_103919_(_093873_, _093888_, _093889_);
  xor g_103920_(out[188], out[892], _093890_);
  and g_103921_(_098195_, out[891], _093891_);
  xor g_103922_(out[184], out[888], _093892_);
  xor g_103923_(out[182], out[886], _093893_);
  xor g_103924_(out[189], out[893], _093894_);
  xor g_103925_(out[190], out[894], _093895_);
  xor g_103926_(out[178], out[882], _093896_);
  xor g_103927_(out[185], out[889], _093897_);
  xor g_103928_(out[181], out[885], _093898_);
  xor g_103929_(out[177], out[881], _093899_);
  and g_103930_(out[187], _049774_, _093900_);
  or g_103931_(_093892_, _093894_, _093901_);
  xor g_103932_(out[191], out[895], _093902_);
  xor g_103933_(out[186], out[890], _093903_);
  xor g_103934_(out[180], out[884], _093904_);
  xor g_103935_(out[179], out[883], _093905_);
  xor g_103936_(out[176], out[880], _093906_);
  or g_103937_(_093896_, _093903_, _093907_);
  or g_103938_(_093901_, _093907_, _093908_);
  or g_103939_(_093897_, _093905_, _093909_);
  or g_103940_(_093898_, _093909_, _093910_);
  or g_103941_(_093908_, _093910_, _093911_);
  or g_103942_(_093895_, _093904_, _093912_);
  or g_103943_(_093911_, _093912_, _093913_);
  or g_103944_(_093890_, _093891_, _093914_);
  xor g_103945_(out[183], out[887], _093915_);
  or g_103946_(_093893_, _093915_, _093916_);
  or g_103947_(_093914_, _093916_, _093917_);
  or g_103948_(_093899_, _093900_, _093918_);
  or g_103949_(_093902_, _093918_, _093919_);
  or g_103950_(_093917_, _093919_, _093920_);
  or g_103951_(_093906_, _093920_, _093921_);
  or g_103952_(_093913_, _093921_, _093922_);
  not g_103953_(_093922_, _093923_);
  xor g_103954_(out[167], out[887], _093924_);
  and g_103955_(_098184_, out[891], _093925_);
  xor g_103956_(out[174], out[894], _093926_);
  xor g_103957_(out[168], out[888], _093927_);
  xor g_103958_(out[161], out[881], _093928_);
  xor g_103959_(out[173], out[893], _093929_);
  xor g_103960_(out[169], out[889], _093930_);
  xor g_103961_(out[164], out[884], _093931_);
  xor g_103962_(out[162], out[882], _093932_);
  and g_103963_(out[171], _049774_, _093933_);
  xor g_103964_(out[163], out[883], _093934_);
  xor g_103965_(out[166], out[886], _093935_);
  xor g_103966_(out[175], out[895], _093936_);
  xor g_103967_(out[170], out[890], _093937_);
  xor g_103968_(out[165], out[885], _093938_);
  xor g_103969_(out[160], out[880], _093939_);
  or g_103970_(_093926_, _093931_, _093940_);
  or g_103971_(_093927_, _093929_, _093941_);
  or g_103972_(_093932_, _093937_, _093942_);
  or g_103973_(_093941_, _093942_, _093943_);
  or g_103974_(_093930_, _093934_, _093944_);
  or g_103975_(_093938_, _093939_, _093945_);
  or g_103976_(_093944_, _093945_, _093946_);
  or g_103977_(_093943_, _093946_, _093947_);
  xor g_103978_(out[172], out[892], _093948_);
  or g_103979_(_093925_, _093948_, _093949_);
  or g_103980_(_093924_, _093935_, _093950_);
  or g_103981_(_093949_, _093950_, _093951_);
  or g_103982_(_093928_, _093933_, _093952_);
  or g_103983_(_093936_, _093952_, _093953_);
  or g_103984_(_093951_, _093953_, _093954_);
  or g_103985_(_093947_, _093954_, _093955_);
  or g_103986_(_093940_, _093955_, _093956_);
  not g_103987_(_093956_, _093957_);
  xor g_103988_(out[145], out[881], _093958_);
  and g_103989_(out[155], _049774_, _093959_);
  xor g_103990_(out[153], out[889], _093960_);
  xor g_103991_(out[144], out[880], _093961_);
  xor g_103992_(out[158], out[894], _093962_);
  xor g_103993_(out[148], out[884], _093963_);
  or g_103994_(_093962_, _093963_, _093964_);
  xor g_103995_(out[157], out[893], _093965_);
  xor g_103996_(out[147], out[883], _093966_);
  and g_103997_(_098173_, out[891], _093967_);
  xor g_103998_(out[150], out[886], _093968_);
  xor g_103999_(out[154], out[890], _093969_);
  xor g_104000_(out[149], out[885], _093970_);
  xor g_104001_(out[159], out[895], _093971_);
  xor g_104002_(out[152], out[888], _093972_);
  or g_104003_(_093965_, _093972_, _093973_);
  xor g_104004_(out[146], out[882], _093974_);
  or g_104005_(_093969_, _093974_, _093975_);
  or g_104006_(_093973_, _093975_, _093976_);
  or g_104007_(_093960_, _093966_, _093977_);
  or g_104008_(_093970_, _093977_, _093978_);
  or g_104009_(_093976_, _093978_, _093979_);
  or g_104010_(_093964_, _093979_, _093980_);
  xor g_104011_(out[156], out[892], _093981_);
  or g_104012_(_093967_, _093981_, _093982_);
  xor g_104013_(out[151], out[887], _093983_);
  or g_104014_(_093968_, _093983_, _093984_);
  or g_104015_(_093982_, _093984_, _093985_);
  or g_104016_(_093958_, _093959_, _093986_);
  or g_104017_(_093971_, _093986_, _093987_);
  or g_104018_(_093985_, _093987_, _093988_);
  or g_104019_(_093961_, _093988_, _093989_);
  or g_104020_(_093980_, _093989_, _093990_);
  not g_104021_(_093990_, _093991_);
  xor g_104022_(out[135], out[887], _093992_);
  and g_104023_(_098162_, out[891], _093993_);
  xor g_104024_(out[142], out[894], _093994_);
  xor g_104025_(out[136], out[888], _093995_);
  xor g_104026_(out[129], out[881], _093996_);
  xor g_104027_(out[141], out[893], _093997_);
  xor g_104028_(out[137], out[889], _093998_);
  xor g_104029_(out[132], out[884], _093999_);
  xor g_104030_(out[130], out[882], _094000_);
  and g_104031_(out[139], _049774_, _094001_);
  xor g_104032_(out[131], out[883], _094002_);
  xor g_104033_(out[134], out[886], _094003_);
  xor g_104034_(out[143], out[895], _094004_);
  xor g_104035_(out[138], out[890], _094005_);
  xor g_104036_(out[133], out[885], _094006_);
  xor g_104037_(out[128], out[880], _094007_);
  or g_104038_(_093994_, _093999_, _094008_);
  or g_104039_(_093995_, _093997_, _094009_);
  or g_104040_(_094000_, _094005_, _094010_);
  or g_104041_(_094009_, _094010_, _094011_);
  or g_104042_(_093998_, _094002_, _094012_);
  or g_104043_(_094006_, _094007_, _094013_);
  or g_104044_(_094012_, _094013_, _094014_);
  or g_104045_(_094011_, _094014_, _094015_);
  xor g_104046_(out[140], out[892], _094016_);
  or g_104047_(_093993_, _094016_, _094017_);
  or g_104048_(_093992_, _094003_, _094018_);
  or g_104049_(_094017_, _094018_, _094019_);
  or g_104050_(_093996_, _094001_, _094020_);
  or g_104051_(_094004_, _094020_, _094021_);
  or g_104052_(_094019_, _094021_, _094022_);
  or g_104053_(_094015_, _094022_, _094023_);
  or g_104054_(_094008_, _094023_, _094024_);
  xor g_104055_(out[113], out[881], _094025_);
  and g_104056_(out[123], _049774_, _094026_);
  xor g_104057_(out[126], out[894], _094027_);
  xor g_104058_(out[115], out[883], _094028_);
  xor g_104059_(out[116], out[884], _094029_);
  xor g_104060_(out[114], out[882], _094030_);
  xor g_104061_(out[121], out[889], _094031_);
  xor g_104062_(out[112], out[880], _094032_);
  and g_104063_(_098151_, out[891], _094033_);
  xor g_104064_(out[118], out[886], _094034_);
  xor g_104065_(out[122], out[890], _094035_);
  xor g_104066_(out[117], out[885], _094036_);
  xor g_104067_(out[127], out[895], _094037_);
  xor g_104068_(out[125], out[893], _094038_);
  xor g_104069_(out[120], out[888], _094039_);
  or g_104070_(_094027_, _094029_, _094040_);
  or g_104071_(_094038_, _094039_, _094041_);
  or g_104072_(_094030_, _094035_, _094042_);
  or g_104073_(_094041_, _094042_, _094043_);
  or g_104074_(_094028_, _094031_, _094044_);
  or g_104075_(_094032_, _094036_, _094045_);
  or g_104076_(_094044_, _094045_, _094046_);
  or g_104077_(_094043_, _094046_, _094047_);
  xor g_104078_(out[124], out[892], _094048_);
  or g_104079_(_094033_, _094048_, _094049_);
  xor g_104080_(out[119], out[887], _094050_);
  or g_104081_(_094034_, _094050_, _094051_);
  or g_104082_(_094049_, _094051_, _094052_);
  or g_104083_(_094025_, _094026_, _094053_);
  or g_104084_(_094037_, _094053_, _094054_);
  or g_104085_(_094052_, _094054_, _094055_);
  or g_104086_(_094047_, _094055_, _094056_);
  or g_104087_(_094040_, _094056_, _094057_);
  not g_104088_(_094057_, _094058_);
  xor g_104089_(out[103], out[887], _094059_);
  and g_104090_(_098140_, out[891], _094060_);
  xor g_104091_(out[110], out[894], _094061_);
  xor g_104092_(out[104], out[888], _094062_);
  xor g_104093_(out[97], out[881], _094063_);
  xor g_104094_(out[109], out[893], _094064_);
  xor g_104095_(out[105], out[889], _094065_);
  xor g_104096_(out[100], out[884], _094066_);
  xor g_104097_(out[98], out[882], _094067_);
  and g_104098_(out[107], _049774_, _094068_);
  xor g_104099_(out[99], out[883], _094069_);
  xor g_104100_(out[102], out[886], _094070_);
  xor g_104101_(out[111], out[895], _094071_);
  xor g_104102_(out[106], out[890], _094072_);
  xor g_104103_(out[101], out[885], _094073_);
  xor g_104104_(out[96], out[880], _094074_);
  or g_104105_(_094061_, _094066_, _094075_);
  or g_104106_(_094062_, _094064_, _094076_);
  or g_104107_(_094067_, _094072_, _094077_);
  or g_104108_(_094076_, _094077_, _094078_);
  or g_104109_(_094065_, _094069_, _094079_);
  or g_104110_(_094073_, _094074_, _094080_);
  or g_104111_(_094079_, _094080_, _094081_);
  or g_104112_(_094078_, _094081_, _094082_);
  xor g_104113_(out[108], out[892], _094083_);
  or g_104114_(_094060_, _094083_, _094084_);
  or g_104115_(_094059_, _094070_, _094085_);
  or g_104116_(_094084_, _094085_, _094086_);
  or g_104117_(_094063_, _094068_, _094087_);
  or g_104118_(_094071_, _094087_, _094088_);
  or g_104119_(_094086_, _094088_, _094089_);
  or g_104120_(_094082_, _094089_, _094090_);
  or g_104121_(_094075_, _094090_, _094091_);
  not g_104122_(_094091_, _094092_);
  and g_104123_(out[91], _049774_, _094093_);
  and g_104124_(_098129_, out[891], _094094_);
  xor g_104125_(out[84], out[884], _094095_);
  xor g_104126_(out[90], out[890], _094096_);
  xor g_104127_(out[85], out[885], _094097_);
  xor g_104128_(out[92], out[892], _094098_);
  xor g_104129_(out[83], out[883], _094099_);
  xor g_104130_(out[88], out[888], _094100_);
  xor g_104131_(out[82], out[882], _094101_);
  xor g_104132_(out[94], out[894], _094102_);
  xor g_104133_(out[89], out[889], _094103_);
  xor g_104134_(out[95], out[895], _094104_);
  xor g_104135_(out[81], out[881], _094105_);
  xor g_104136_(out[86], out[886], _094106_);
  xor g_104137_(out[80], out[880], _094107_);
  xor g_104138_(out[93], out[893], _094108_);
  or g_104139_(_094095_, _094102_, _094109_);
  or g_104140_(_094100_, _094108_, _094110_);
  or g_104141_(_094096_, _094101_, _094111_);
  or g_104142_(_094110_, _094111_, _094112_);
  or g_104143_(_094099_, _094103_, _094113_);
  or g_104144_(_094097_, _094107_, _094114_);
  or g_104145_(_094113_, _094114_, _094115_);
  or g_104146_(_094112_, _094115_, _094116_);
  or g_104147_(_094094_, _094098_, _094117_);
  xor g_104148_(out[87], out[887], _094118_);
  or g_104149_(_094106_, _094118_, _094119_);
  or g_104150_(_094117_, _094119_, _094120_);
  or g_104151_(_094093_, _094105_, _094121_);
  or g_104152_(_094104_, _094121_, _094122_);
  or g_104153_(_094120_, _094122_, _094123_);
  or g_104154_(_094116_, _094123_, _094124_);
  or g_104155_(_094109_, _094124_, _094125_);
  xor g_104156_(out[71], out[887], _094126_);
  and g_104157_(_098118_, out[891], _094127_);
  xor g_104158_(out[78], out[894], _094128_);
  xor g_104159_(out[72], out[888], _094129_);
  xor g_104160_(out[65], out[881], _094130_);
  xor g_104161_(out[77], out[893], _094131_);
  xor g_104162_(out[73], out[889], _094132_);
  xor g_104163_(out[68], out[884], _094133_);
  xor g_104164_(out[66], out[882], _094134_);
  and g_104165_(out[75], _049774_, _094135_);
  xor g_104166_(out[67], out[883], _094136_);
  xor g_104167_(out[70], out[886], _094137_);
  xor g_104168_(out[79], out[895], _094138_);
  xor g_104169_(out[74], out[890], _094139_);
  xor g_104170_(out[69], out[885], _094140_);
  xor g_104171_(out[64], out[880], _094141_);
  or g_104172_(_094128_, _094133_, _094142_);
  or g_104173_(_094129_, _094131_, _094143_);
  or g_104174_(_094134_, _094139_, _094144_);
  or g_104175_(_094143_, _094144_, _094145_);
  or g_104176_(_094132_, _094136_, _094146_);
  or g_104177_(_094140_, _094141_, _094147_);
  or g_104178_(_094146_, _094147_, _094148_);
  or g_104179_(_094145_, _094148_, _094149_);
  xor g_104180_(out[76], out[892], _094150_);
  or g_104181_(_094127_, _094150_, _094151_);
  or g_104182_(_094126_, _094137_, _094152_);
  or g_104183_(_094151_, _094152_, _094153_);
  or g_104184_(_094130_, _094135_, _094154_);
  or g_104185_(_094138_, _094154_, _094155_);
  or g_104186_(_094153_, _094155_, _094156_);
  or g_104187_(_094149_, _094156_, _094157_);
  or g_104188_(_094142_, _094157_, _094158_);
  xor g_104189_(out[50], out[882], _094159_);
  xor g_104190_(out[48], out[880], _094160_);
  xor g_104191_(out[57], out[889], _094161_);
  xor g_104192_(out[56], out[888], _094162_);
  xor g_104193_(out[53], out[885], _094163_);
  xor g_104194_(out[62], out[894], _094164_);
  xor g_104195_(out[61], out[893], _094165_);
  xor g_104196_(out[63], out[895], _094166_);
  xor g_104197_(out[58], out[890], _094167_);
  xor g_104198_(out[54], out[886], _094168_);
  xor g_104199_(out[51], out[883], _094169_);
  and g_104200_(_098107_, out[891], _094170_);
  and g_104201_(out[59], _049774_, _094171_);
  xor g_104202_(out[52], out[884], _094172_);
  xor g_104203_(out[49], out[881], _094173_);
  or g_104204_(_094164_, _094172_, _094174_);
  or g_104205_(_094162_, _094165_, _094175_);
  or g_104206_(_094159_, _094167_, _094176_);
  or g_104207_(_094175_, _094176_, _094177_);
  or g_104208_(_094161_, _094169_, _094178_);
  or g_104209_(_094160_, _094163_, _094179_);
  or g_104210_(_094178_, _094179_, _094180_);
  or g_104211_(_094177_, _094180_, _094181_);
  xor g_104212_(out[60], out[892], _094182_);
  or g_104213_(_094170_, _094182_, _094183_);
  xor g_104214_(out[55], out[887], _094184_);
  or g_104215_(_094168_, _094184_, _094185_);
  or g_104216_(_094183_, _094185_, _094186_);
  or g_104217_(_094171_, _094173_, _094187_);
  or g_104218_(_094166_, _094187_, _094188_);
  or g_104219_(_094186_, _094188_, _094189_);
  or g_104220_(_094181_, _094189_, _094190_);
  or g_104221_(_094174_, _094190_, _094191_);
  not g_104222_(_094191_, _094192_);
  xor g_104223_(out[39], out[887], _094193_);
  and g_104224_(_098096_, out[891], _094194_);
  xor g_104225_(out[46], out[894], _094195_);
  xor g_104226_(out[40], out[888], _094196_);
  xor g_104227_(out[33], out[881], _094197_);
  xor g_104228_(out[45], out[893], _094198_);
  xor g_104229_(out[41], out[889], _094199_);
  xor g_104230_(out[36], out[884], _094200_);
  xor g_104231_(out[34], out[882], _094201_);
  and g_104232_(out[43], _049774_, _094202_);
  xor g_104233_(out[35], out[883], _094203_);
  xor g_104234_(out[38], out[886], _094204_);
  xor g_104235_(out[47], out[895], _094205_);
  xor g_104236_(out[42], out[890], _094206_);
  xor g_104237_(out[37], out[885], _094207_);
  xor g_104238_(out[32], out[880], _094208_);
  or g_104239_(_094195_, _094200_, _094209_);
  or g_104240_(_094196_, _094198_, _094210_);
  or g_104241_(_094201_, _094206_, _094211_);
  or g_104242_(_094210_, _094211_, _094212_);
  or g_104243_(_094199_, _094203_, _094213_);
  or g_104244_(_094207_, _094208_, _094214_);
  or g_104245_(_094213_, _094214_, _094215_);
  or g_104246_(_094212_, _094215_, _094216_);
  xor g_104247_(out[44], out[892], _094217_);
  or g_104248_(_094194_, _094217_, _094218_);
  or g_104249_(_094193_, _094204_, _094219_);
  or g_104250_(_094218_, _094219_, _094220_);
  or g_104251_(_094197_, _094202_, _094221_);
  or g_104252_(_094205_, _094221_, _094222_);
  or g_104253_(_094220_, _094222_, _094223_);
  or g_104254_(_094216_, _094223_, _094224_);
  or g_104255_(_094209_, _094224_, _094225_);
  not g_104256_(_094225_, _094226_);
  and g_104257_(out[27], _049774_, _094227_);
  and g_104258_(_098063_, out[891], _094228_);
  xor g_104259_(out[29], out[893], _094229_);
  xor g_104260_(out[26], out[890], _094230_);
  xor g_104261_(out[21], out[885], _094231_);
  xor g_104262_(out[28], out[892], _094232_);
  xor g_104263_(out[16], out[880], _094233_);
  xor g_104264_(out[18], out[882], _094234_);
  xor g_104265_(out[19], out[883], _094235_);
  xor g_104266_(out[25], out[889], _094236_);
  xor g_104267_(out[30], out[894], _094237_);
  xor g_104268_(out[31], out[895], _094238_);
  xor g_104269_(out[17], out[881], _094239_);
  xor g_104270_(out[22], out[886], _094240_);
  xor g_104271_(out[20], out[884], _094241_);
  xor g_104272_(out[24], out[888], _094242_);
  or g_104273_(_094229_, _094242_, _094243_);
  or g_104274_(_094230_, _094234_, _094244_);
  or g_104275_(_094243_, _094244_, _094245_);
  or g_104276_(_094235_, _094236_, _094246_);
  or g_104277_(_094231_, _094246_, _094247_);
  or g_104278_(_094245_, _094247_, _094248_);
  or g_104279_(_094237_, _094241_, _094249_);
  or g_104280_(_094248_, _094249_, _094250_);
  or g_104281_(_094228_, _094232_, _094251_);
  xor g_104282_(out[23], out[887], _094252_);
  or g_104283_(_094240_, _094252_, _094253_);
  or g_104284_(_094251_, _094253_, _094254_);
  or g_104285_(_094227_, _094239_, _094255_);
  or g_104286_(_094238_, _094255_, _094256_);
  or g_104287_(_094254_, _094256_, _094257_);
  or g_104288_(_094233_, _094257_, _094258_);
  or g_104289_(_094250_, _094258_, _094259_);
  not g_104290_(_094259_, _094260_);
  xor g_104291_(out[0], out[880], _094261_);
  xor g_104292_(out[8], out[888], _094262_);
  xor g_104293_(out[6], out[886], _094263_);
  xor g_104294_(out[2], out[882], _094264_);
  and g_104295_(_098041_, out[891], _094265_);
  and g_104296_(out[11], _049774_, _094266_);
  xor g_104297_(out[4], out[884], _094267_);
  xor g_104298_(out[1], out[881], _094268_);
  xor g_104299_(out[13], out[893], _094269_);
  xor g_104300_(out[3], out[883], _094270_);
  xor g_104301_(out[5], out[885], _094271_);
  xor g_104302_(out[15], out[895], _094272_);
  xor g_104303_(out[10], out[890], _094273_);
  xor g_104304_(out[14], out[894], _094274_);
  or g_104305_(_094262_, _094269_, _094275_);
  xor g_104306_(out[9], out[889], _094276_);
  or g_104307_(_094264_, _094273_, _094277_);
  or g_104308_(_094275_, _094277_, _094278_);
  or g_104309_(_094270_, _094276_, _094279_);
  or g_104310_(_094271_, _094279_, _094280_);
  or g_104311_(_094278_, _094280_, _094281_);
  or g_104312_(_094267_, _094274_, _094282_);
  or g_104313_(_094281_, _094282_, _094283_);
  xor g_104314_(out[12], out[892], _094284_);
  or g_104315_(_094265_, _094284_, _094285_);
  xor g_104316_(out[7], out[887], _094286_);
  or g_104317_(_094263_, _094286_, _094287_);
  or g_104318_(_094285_, _094287_, _094288_);
  or g_104319_(_094266_, _094268_, _094289_);
  or g_104320_(_094272_, _094289_, _094290_);
  or g_104321_(_094288_, _094290_, _094291_);
  or g_104322_(_094261_, _094291_, _094292_);
  or g_104323_(_094283_, _094292_, _094293_);
  not g_104324_(_094293_, _094294_);
  xor g_104325_(out[471], out[871], _094295_);
  and g_104326_(_049499_, out[875], _094296_);
  xor g_104327_(out[478], out[878], _094297_);
  xor g_104328_(out[472], out[872], _094298_);
  xor g_104329_(out[465], out[865], _094299_);
  xor g_104330_(out[477], out[877], _094300_);
  xor g_104331_(out[473], out[873], _094301_);
  xor g_104332_(out[468], out[868], _094302_);
  xor g_104333_(out[466], out[866], _094303_);
  and g_104334_(out[475], _049763_, _094304_);
  xor g_104335_(out[467], out[867], _094305_);
  xor g_104336_(out[470], out[870], _094306_);
  xor g_104337_(out[479], out[879], _094307_);
  xor g_104338_(out[474], out[874], _094308_);
  xor g_104339_(out[469], out[869], _094309_);
  xor g_104340_(out[464], out[864], _094310_);
  or g_104341_(_094297_, _094302_, _094311_);
  or g_104342_(_094298_, _094300_, _094312_);
  or g_104343_(_094303_, _094308_, _094313_);
  or g_104344_(_094312_, _094313_, _094314_);
  or g_104345_(_094301_, _094305_, _094315_);
  or g_104346_(_094309_, _094310_, _094316_);
  or g_104347_(_094315_, _094316_, _094317_);
  or g_104348_(_094314_, _094317_, _094318_);
  xor g_104349_(out[476], out[876], _094319_);
  or g_104350_(_094296_, _094319_, _094320_);
  or g_104351_(_094295_, _094306_, _094321_);
  or g_104352_(_094320_, _094321_, _094322_);
  or g_104353_(_094299_, _094304_, _094323_);
  or g_104354_(_094307_, _094323_, _094324_);
  or g_104355_(_094322_, _094324_, _094325_);
  or g_104356_(_094318_, _094325_, _094326_);
  or g_104357_(_094311_, _094326_, _094327_);
  not g_104358_(_094327_, _094328_);
  and g_104359_(out[459], _049763_, _094329_);
  xor g_104360_(out[452], out[868], _094330_);
  xor g_104361_(out[462], out[878], _094331_);
  or g_104362_(_094330_, _094331_, _094332_);
  xor g_104363_(out[461], out[877], _094333_);
  xor g_104364_(out[451], out[867], _094334_);
  xor g_104365_(out[448], out[864], _094335_);
  and g_104366_(_049477_, out[875], _094336_);
  xor g_104367_(out[458], out[874], _094337_);
  xor g_104368_(out[463], out[879], _094338_);
  xor g_104369_(out[454], out[870], _094339_);
  xor g_104370_(out[453], out[869], _094340_);
  xor g_104371_(out[456], out[872], _094341_);
  or g_104372_(_094333_, _094341_, _094342_);
  xor g_104373_(out[450], out[866], _094343_);
  xor g_104374_(out[457], out[873], _094344_);
  xor g_104375_(out[449], out[865], _094345_);
  or g_104376_(_094337_, _094343_, _094346_);
  or g_104377_(_094342_, _094346_, _094347_);
  or g_104378_(_094334_, _094344_, _094348_);
  or g_104379_(_094340_, _094348_, _094349_);
  or g_104380_(_094347_, _094349_, _094350_);
  or g_104381_(_094332_, _094350_, _094351_);
  xor g_104382_(out[460], out[876], _094352_);
  or g_104383_(_094336_, _094352_, _094353_);
  xor g_104384_(out[455], out[871], _094354_);
  or g_104385_(_094339_, _094354_, _094355_);
  or g_104386_(_094353_, _094355_, _094356_);
  or g_104387_(_094329_, _094345_, _094357_);
  or g_104388_(_094338_, _094357_, _094358_);
  or g_104389_(_094356_, _094358_, _094359_);
  or g_104390_(_094335_, _094359_, _094360_);
  or g_104391_(_094351_, _094360_, _094361_);
  xor g_104392_(out[439], out[871], _094362_);
  and g_104393_(_049466_, out[875], _094363_);
  xor g_104394_(out[446], out[878], _094364_);
  xor g_104395_(out[440], out[872], _094365_);
  xor g_104396_(out[433], out[865], _094366_);
  xor g_104397_(out[445], out[877], _094367_);
  xor g_104398_(out[441], out[873], _094368_);
  xor g_104399_(out[436], out[868], _094369_);
  xor g_104400_(out[434], out[866], _094370_);
  and g_104401_(out[443], _049763_, _094371_);
  xor g_104402_(out[435], out[867], _094372_);
  xor g_104403_(out[438], out[870], _094373_);
  xor g_104404_(out[447], out[879], _094374_);
  xor g_104405_(out[442], out[874], _094375_);
  xor g_104406_(out[437], out[869], _094376_);
  xor g_104407_(out[432], out[864], _094377_);
  or g_104408_(_094364_, _094369_, _094378_);
  or g_104409_(_094365_, _094367_, _094379_);
  or g_104410_(_094370_, _094375_, _094380_);
  or g_104411_(_094379_, _094380_, _094381_);
  or g_104412_(_094368_, _094372_, _094382_);
  or g_104413_(_094376_, _094377_, _094383_);
  or g_104414_(_094382_, _094383_, _094384_);
  or g_104415_(_094381_, _094384_, _094385_);
  xor g_104416_(out[444], out[876], _094386_);
  or g_104417_(_094363_, _094386_, _094387_);
  or g_104418_(_094362_, _094373_, _094388_);
  or g_104419_(_094387_, _094388_, _094389_);
  or g_104420_(_094366_, _094371_, _094390_);
  or g_104421_(_094374_, _094390_, _094391_);
  or g_104422_(_094389_, _094391_, _094392_);
  or g_104423_(_094385_, _094392_, _094393_);
  or g_104424_(_094378_, _094393_, _094394_);
  xor g_104425_(out[424], out[872], _094395_);
  xor g_104426_(out[421], out[869], _094396_);
  xor g_104427_(out[419], out[867], _094397_);
  xor g_104428_(out[430], out[878], _094398_);
  xor g_104429_(out[429], out[877], _094399_);
  xor g_104430_(out[418], out[866], _094400_);
  xor g_104431_(out[425], out[873], _094401_);
  xor g_104432_(out[422], out[870], _094402_);
  xor g_104433_(out[431], out[879], _094403_);
  xor g_104434_(out[426], out[874], _094404_);
  xor g_104435_(out[420], out[868], _094405_);
  xor g_104436_(out[416], out[864], _094406_);
  and g_104437_(_049455_, out[875], _094407_);
  and g_104438_(out[427], _049763_, _094408_);
  or g_104439_(_094395_, _094399_, _094409_);
  xor g_104440_(out[417], out[865], _094410_);
  or g_104441_(_094400_, _094404_, _094411_);
  or g_104442_(_094409_, _094411_, _094412_);
  or g_104443_(_094397_, _094401_, _094413_);
  or g_104444_(_094396_, _094413_, _094414_);
  or g_104445_(_094412_, _094414_, _094415_);
  or g_104446_(_094398_, _094405_, _094416_);
  or g_104447_(_094415_, _094416_, _094417_);
  xor g_104448_(out[428], out[876], _094418_);
  or g_104449_(_094407_, _094418_, _094419_);
  xor g_104450_(out[423], out[871], _094420_);
  or g_104451_(_094402_, _094420_, _094421_);
  or g_104452_(_094419_, _094421_, _094422_);
  or g_104453_(_094408_, _094410_, _094423_);
  or g_104454_(_094403_, _094423_, _094424_);
  or g_104455_(_094422_, _094424_, _094425_);
  or g_104456_(_094406_, _094425_, _094426_);
  or g_104457_(_094417_, _094426_, _094427_);
  xor g_104458_(out[407], out[871], _094428_);
  and g_104459_(_049444_, out[875], _094429_);
  xor g_104460_(out[414], out[878], _094430_);
  xor g_104461_(out[408], out[872], _094431_);
  xor g_104462_(out[401], out[865], _094432_);
  xor g_104463_(out[413], out[877], _094433_);
  xor g_104464_(out[409], out[873], _094434_);
  xor g_104465_(out[404], out[868], _094435_);
  xor g_104466_(out[402], out[866], _094436_);
  and g_104467_(out[411], _049763_, _094437_);
  xor g_104468_(out[403], out[867], _094438_);
  xor g_104469_(out[406], out[870], _094439_);
  xor g_104470_(out[415], out[879], _094440_);
  xor g_104471_(out[410], out[874], _094441_);
  xor g_104472_(out[405], out[869], _094442_);
  xor g_104473_(out[400], out[864], _094443_);
  or g_104474_(_094430_, _094435_, _094444_);
  or g_104475_(_094431_, _094433_, _094445_);
  or g_104476_(_094436_, _094441_, _094446_);
  or g_104477_(_094445_, _094446_, _094447_);
  or g_104478_(_094434_, _094438_, _094448_);
  or g_104479_(_094442_, _094443_, _094449_);
  or g_104480_(_094448_, _094449_, _094450_);
  or g_104481_(_094447_, _094450_, _094451_);
  xor g_104482_(out[412], out[876], _094452_);
  or g_104483_(_094429_, _094452_, _094453_);
  or g_104484_(_094428_, _094439_, _094454_);
  or g_104485_(_094453_, _094454_, _094455_);
  or g_104486_(_094432_, _094437_, _094456_);
  or g_104487_(_094440_, _094456_, _094457_);
  or g_104488_(_094455_, _094457_, _094458_);
  or g_104489_(_094451_, _094458_, _094459_);
  or g_104490_(_094444_, _094459_, _094460_);
  xor g_104491_(out[394], out[874], _094461_);
  xor g_104492_(out[386], out[866], _094462_);
  xor g_104493_(out[385], out[865], _094463_);
  and g_104494_(_049433_, out[875], _094464_);
  and g_104495_(out[395], _049763_, _094465_);
  xor g_104496_(out[397], out[877], _094466_);
  xor g_104497_(out[387], out[867], _094467_);
  xor g_104498_(out[398], out[878], _094468_);
  xor g_104499_(out[396], out[876], _094469_);
  xor g_104500_(out[392], out[872], _094470_);
  xor g_104501_(out[399], out[879], _094471_);
  xor g_104502_(out[389], out[869], _094472_);
  xor g_104503_(out[390], out[870], _094473_);
  xor g_104504_(out[384], out[864], _094474_);
  xor g_104505_(out[388], out[868], _094475_);
  or g_104506_(_094466_, _094470_, _094476_);
  xor g_104507_(out[393], out[873], _094477_);
  or g_104508_(_094461_, _094462_, _094478_);
  or g_104509_(_094476_, _094478_, _094479_);
  or g_104510_(_094467_, _094477_, _094480_);
  or g_104511_(_094472_, _094480_, _094481_);
  or g_104512_(_094479_, _094481_, _094482_);
  or g_104513_(_094468_, _094475_, _094483_);
  or g_104514_(_094482_, _094483_, _094484_);
  or g_104515_(_094464_, _094469_, _094485_);
  xor g_104516_(out[391], out[871], _094486_);
  or g_104517_(_094473_, _094486_, _094487_);
  or g_104518_(_094485_, _094487_, _094488_);
  or g_104519_(_094463_, _094465_, _094489_);
  or g_104520_(_094471_, _094489_, _094490_);
  or g_104521_(_094488_, _094490_, _094491_);
  or g_104522_(_094474_, _094491_, _094492_);
  or g_104523_(_094484_, _094492_, _094493_);
  xor g_104524_(out[375], out[871], _094494_);
  and g_104525_(_049422_, out[875], _094495_);
  xor g_104526_(out[382], out[878], _094496_);
  xor g_104527_(out[376], out[872], _094497_);
  xor g_104528_(out[369], out[865], _094498_);
  xor g_104529_(out[381], out[877], _094499_);
  xor g_104530_(out[377], out[873], _094500_);
  xor g_104531_(out[372], out[868], _094501_);
  xor g_104532_(out[370], out[866], _094502_);
  and g_104533_(out[379], _049763_, _094503_);
  xor g_104534_(out[371], out[867], _094504_);
  xor g_104535_(out[374], out[870], _094505_);
  xor g_104536_(out[383], out[879], _094506_);
  xor g_104537_(out[378], out[874], _094507_);
  xor g_104538_(out[373], out[869], _094508_);
  xor g_104539_(out[368], out[864], _094509_);
  or g_104540_(_094496_, _094501_, _094510_);
  or g_104541_(_094497_, _094499_, _094511_);
  or g_104542_(_094502_, _094507_, _094512_);
  or g_104543_(_094511_, _094512_, _094513_);
  or g_104544_(_094500_, _094504_, _094514_);
  or g_104545_(_094508_, _094509_, _094515_);
  or g_104546_(_094514_, _094515_, _094516_);
  or g_104547_(_094513_, _094516_, _094517_);
  xor g_104548_(out[380], out[876], _094518_);
  or g_104549_(_094495_, _094518_, _094519_);
  or g_104550_(_094494_, _094505_, _094520_);
  or g_104551_(_094519_, _094520_, _094521_);
  or g_104552_(_094498_, _094503_, _094522_);
  or g_104553_(_094506_, _094522_, _094523_);
  or g_104554_(_094521_, _094523_, _094524_);
  or g_104555_(_094517_, _094524_, _094525_);
  or g_104556_(_094510_, _094525_, _094526_);
  xor g_104557_(out[360], out[872], _094527_);
  xor g_104558_(out[357], out[869], _094528_);
  xor g_104559_(out[355], out[867], _094529_);
  xor g_104560_(out[366], out[878], _094530_);
  xor g_104561_(out[365], out[877], _094531_);
  xor g_104562_(out[354], out[866], _094532_);
  xor g_104563_(out[361], out[873], _094533_);
  xor g_104564_(out[358], out[870], _094534_);
  xor g_104565_(out[367], out[879], _094535_);
  xor g_104566_(out[362], out[874], _094536_);
  xor g_104567_(out[356], out[868], _094537_);
  xor g_104568_(out[352], out[864], _094538_);
  and g_104569_(_049411_, out[875], _094539_);
  and g_104570_(out[363], _049763_, _094540_);
  or g_104571_(_094527_, _094531_, _094541_);
  xor g_104572_(out[353], out[865], _094542_);
  or g_104573_(_094532_, _094536_, _094543_);
  or g_104574_(_094541_, _094543_, _094544_);
  or g_104575_(_094529_, _094533_, _094545_);
  or g_104576_(_094528_, _094545_, _094546_);
  or g_104577_(_094544_, _094546_, _094547_);
  or g_104578_(_094530_, _094537_, _094548_);
  or g_104579_(_094547_, _094548_, _094549_);
  xor g_104580_(out[364], out[876], _094550_);
  or g_104581_(_094539_, _094550_, _094551_);
  xor g_104582_(out[359], out[871], _094552_);
  or g_104583_(_094534_, _094552_, _094553_);
  or g_104584_(_094551_, _094553_, _094554_);
  or g_104585_(_094540_, _094542_, _094555_);
  or g_104586_(_094535_, _094555_, _094556_);
  or g_104587_(_094554_, _094556_, _094557_);
  or g_104588_(_094538_, _094557_, _094558_);
  or g_104589_(_094549_, _094558_, _094559_);
  xor g_104590_(out[343], out[871], _094560_);
  and g_104591_(_049400_, out[875], _094561_);
  xor g_104592_(out[350], out[878], _094562_);
  xor g_104593_(out[344], out[872], _094563_);
  xor g_104594_(out[337], out[865], _094564_);
  xor g_104595_(out[349], out[877], _094565_);
  xor g_104596_(out[345], out[873], _094566_);
  xor g_104597_(out[340], out[868], _094567_);
  xor g_104598_(out[338], out[866], _094568_);
  and g_104599_(out[347], _049763_, _094569_);
  xor g_104600_(out[339], out[867], _094570_);
  xor g_104601_(out[342], out[870], _094571_);
  xor g_104602_(out[351], out[879], _094572_);
  xor g_104603_(out[346], out[874], _094573_);
  xor g_104604_(out[341], out[869], _094574_);
  xor g_104605_(out[336], out[864], _094575_);
  or g_104606_(_094562_, _094567_, _094576_);
  not g_104607_(_094576_, _094577_);
  or g_104608_(_094563_, _094565_, _094578_);
  or g_104609_(_094568_, _094573_, _094579_);
  or g_104610_(_094578_, _094579_, _094580_);
  or g_104611_(_094566_, _094570_, _094581_);
  or g_104612_(_094574_, _094575_, _094582_);
  or g_104613_(_094581_, _094582_, _094583_);
  or g_104614_(_094580_, _094583_, _094584_);
  xor g_104615_(out[348], out[876], _094585_);
  or g_104616_(_094561_, _094585_, _094586_);
  or g_104617_(_094560_, _094571_, _094587_);
  or g_104618_(_094586_, _094587_, _094588_);
  or g_104619_(_094564_, _094569_, _094589_);
  or g_104620_(_094572_, _094589_, _094590_);
  or g_104621_(_094588_, _094590_, _094591_);
  or g_104622_(_094584_, _094591_, _094592_);
  not g_104623_(_094592_, _094593_);
  and g_104624_(_094577_, _094593_, _094594_);
  not g_104625_(_094594_, _094595_);
  xor g_104626_(out[321], out[865], _094596_);
  and g_104627_(out[331], _049763_, _094597_);
  xor g_104628_(out[329], out[873], _094598_);
  xor g_104629_(out[320], out[864], _094599_);
  xor g_104630_(out[334], out[878], _094600_);
  xor g_104631_(out[324], out[868], _094601_);
  or g_104632_(_094600_, _094601_, _094602_);
  xor g_104633_(out[333], out[877], _094603_);
  xor g_104634_(out[323], out[867], _094604_);
  and g_104635_(_098294_, out[875], _094605_);
  xor g_104636_(out[326], out[870], _094606_);
  xor g_104637_(out[330], out[874], _094607_);
  xor g_104638_(out[325], out[869], _094608_);
  xor g_104639_(out[335], out[879], _094609_);
  xor g_104640_(out[328], out[872], _094610_);
  or g_104641_(_094603_, _094610_, _094611_);
  xor g_104642_(out[322], out[866], _094612_);
  or g_104643_(_094607_, _094612_, _094613_);
  or g_104644_(_094611_, _094613_, _094614_);
  or g_104645_(_094598_, _094604_, _094615_);
  or g_104646_(_094608_, _094615_, _094616_);
  or g_104647_(_094614_, _094616_, _094617_);
  or g_104648_(_094602_, _094617_, _094618_);
  xor g_104649_(out[332], out[876], _094619_);
  or g_104650_(_094605_, _094619_, _094620_);
  xor g_104651_(out[327], out[871], _094621_);
  or g_104652_(_094606_, _094621_, _094622_);
  or g_104653_(_094620_, _094622_, _094623_);
  or g_104654_(_094596_, _094597_, _094624_);
  or g_104655_(_094609_, _094624_, _094625_);
  or g_104656_(_094623_, _094625_, _094626_);
  or g_104657_(_094599_, _094626_, _094627_);
  or g_104658_(_094618_, _094627_, _094628_);
  not g_104659_(_094628_, _094629_);
  xor g_104660_(out[311], out[871], _094630_);
  and g_104661_(_098283_, out[875], _094631_);
  xor g_104662_(out[318], out[878], _094632_);
  xor g_104663_(out[312], out[872], _094633_);
  xor g_104664_(out[305], out[865], _094634_);
  xor g_104665_(out[317], out[877], _094635_);
  xor g_104666_(out[313], out[873], _094636_);
  xor g_104667_(out[308], out[868], _094637_);
  xor g_104668_(out[306], out[866], _094638_);
  and g_104669_(out[315], _049763_, _094639_);
  xor g_104670_(out[307], out[867], _094640_);
  xor g_104671_(out[310], out[870], _094641_);
  xor g_104672_(out[319], out[879], _094642_);
  xor g_104673_(out[314], out[874], _094643_);
  xor g_104674_(out[309], out[869], _094644_);
  xor g_104675_(out[304], out[864], _094645_);
  or g_104676_(_094632_, _094637_, _094646_);
  or g_104677_(_094633_, _094635_, _094647_);
  or g_104678_(_094638_, _094643_, _094648_);
  or g_104679_(_094647_, _094648_, _094649_);
  or g_104680_(_094636_, _094640_, _094650_);
  or g_104681_(_094644_, _094645_, _094651_);
  or g_104682_(_094650_, _094651_, _094652_);
  or g_104683_(_094649_, _094652_, _094653_);
  xor g_104684_(out[316], out[876], _094654_);
  or g_104685_(_094631_, _094654_, _094655_);
  or g_104686_(_094630_, _094641_, _094656_);
  or g_104687_(_094655_, _094656_, _094657_);
  or g_104688_(_094634_, _094639_, _094658_);
  or g_104689_(_094642_, _094658_, _094659_);
  or g_104690_(_094657_, _094659_, _094660_);
  or g_104691_(_094653_, _094660_, _094661_);
  or g_104692_(_094646_, _094661_, _094662_);
  and g_104693_(out[299], _049763_, _094663_);
  xor g_104694_(out[292], out[868], _094664_);
  xor g_104695_(out[291], out[867], _094665_);
  xor g_104696_(out[295], out[871], _094666_);
  xor g_104697_(out[302], out[878], _094667_);
  and g_104698_(_098272_, out[875], _094668_);
  xor g_104699_(out[301], out[877], _094669_);
  xor g_104700_(out[290], out[866], _094670_);
  xor g_104701_(out[297], out[873], _094671_);
  xor g_104702_(out[288], out[864], _094672_);
  xor g_104703_(out[296], out[872], _094673_);
  xor g_104704_(out[294], out[870], _094674_);
  xor g_104705_(out[293], out[869], _094675_);
  xor g_104706_(out[303], out[879], _094676_);
  xor g_104707_(out[298], out[874], _094677_);
  or g_104708_(_094669_, _094673_, _094678_);
  xor g_104709_(out[289], out[865], _094679_);
  or g_104710_(_094670_, _094677_, _094680_);
  or g_104711_(_094678_, _094680_, _094681_);
  or g_104712_(_094665_, _094671_, _094682_);
  or g_104713_(_094675_, _094682_, _094683_);
  or g_104714_(_094681_, _094683_, _094684_);
  or g_104715_(_094664_, _094667_, _094685_);
  or g_104716_(_094684_, _094685_, _094686_);
  xor g_104717_(out[300], out[876], _094687_);
  or g_104718_(_094668_, _094687_, _094688_);
  or g_104719_(_094666_, _094674_, _094689_);
  or g_104720_(_094688_, _094689_, _094690_);
  or g_104721_(_094663_, _094679_, _094691_);
  or g_104722_(_094676_, _094691_, _094692_);
  or g_104723_(_094690_, _094692_, _094693_);
  or g_104724_(_094672_, _094693_, _094694_);
  or g_104725_(_094686_, _094694_, _094695_);
  not g_104726_(_094695_, _094696_);
  xor g_104727_(out[279], out[871], _094697_);
  and g_104728_(_098261_, out[875], _094698_);
  xor g_104729_(out[286], out[878], _094699_);
  xor g_104730_(out[280], out[872], _094700_);
  xor g_104731_(out[273], out[865], _094701_);
  xor g_104732_(out[285], out[877], _094702_);
  xor g_104733_(out[281], out[873], _094703_);
  xor g_104734_(out[276], out[868], _094704_);
  xor g_104735_(out[274], out[866], _094705_);
  and g_104736_(out[283], _049763_, _094706_);
  xor g_104737_(out[275], out[867], _094707_);
  xor g_104738_(out[278], out[870], _094708_);
  xor g_104739_(out[287], out[879], _094709_);
  xor g_104740_(out[282], out[874], _094710_);
  xor g_104741_(out[277], out[869], _094711_);
  xor g_104742_(out[272], out[864], _094712_);
  or g_104743_(_094699_, _094704_, _094713_);
  or g_104744_(_094700_, _094702_, _094714_);
  or g_104745_(_094705_, _094710_, _094715_);
  or g_104746_(_094714_, _094715_, _094716_);
  or g_104747_(_094703_, _094707_, _094717_);
  or g_104748_(_094711_, _094712_, _094718_);
  or g_104749_(_094717_, _094718_, _094719_);
  or g_104750_(_094716_, _094719_, _094720_);
  xor g_104751_(out[284], out[876], _094721_);
  or g_104752_(_094698_, _094721_, _094722_);
  or g_104753_(_094697_, _094708_, _094723_);
  or g_104754_(_094722_, _094723_, _094724_);
  or g_104755_(_094701_, _094706_, _094725_);
  or g_104756_(_094709_, _094725_, _094726_);
  or g_104757_(_094724_, _094726_, _094727_);
  or g_104758_(_094720_, _094727_, _094728_);
  or g_104759_(_094713_, _094728_, _094729_);
  not g_104760_(_094729_, _094730_);
  xor g_104761_(out[257], out[865], _094731_);
  and g_104762_(out[267], _049763_, _094732_);
  xor g_104763_(out[265], out[873], _094733_);
  xor g_104764_(out[256], out[864], _094734_);
  xor g_104765_(out[270], out[878], _094735_);
  xor g_104766_(out[260], out[868], _094736_);
  or g_104767_(_094735_, _094736_, _094737_);
  xor g_104768_(out[269], out[877], _094738_);
  xor g_104769_(out[259], out[867], _094739_);
  and g_104770_(_098250_, out[875], _094740_);
  xor g_104771_(out[262], out[870], _094741_);
  xor g_104772_(out[266], out[874], _094742_);
  xor g_104773_(out[261], out[869], _094743_);
  xor g_104774_(out[271], out[879], _094744_);
  xor g_104775_(out[264], out[872], _094745_);
  or g_104776_(_094738_, _094745_, _094746_);
  xor g_104777_(out[258], out[866], _094747_);
  or g_104778_(_094742_, _094747_, _094748_);
  or g_104779_(_094746_, _094748_, _094749_);
  or g_104780_(_094733_, _094739_, _094750_);
  or g_104781_(_094743_, _094750_, _094751_);
  or g_104782_(_094749_, _094751_, _094752_);
  or g_104783_(_094737_, _094752_, _094753_);
  xor g_104784_(out[268], out[876], _094754_);
  or g_104785_(_094740_, _094754_, _094755_);
  xor g_104786_(out[263], out[871], _094756_);
  or g_104787_(_094741_, _094756_, _094757_);
  or g_104788_(_094755_, _094757_, _094758_);
  or g_104789_(_094731_, _094732_, _094759_);
  or g_104790_(_094744_, _094759_, _094760_);
  or g_104791_(_094758_, _094760_, _094761_);
  or g_104792_(_094734_, _094761_, _094762_);
  or g_104793_(_094753_, _094762_, _094763_);
  xor g_104794_(out[247], out[871], _094764_);
  and g_104795_(_098239_, out[875], _094765_);
  xor g_104796_(out[254], out[878], _094766_);
  xor g_104797_(out[248], out[872], _094767_);
  xor g_104798_(out[241], out[865], _094768_);
  xor g_104799_(out[253], out[877], _094769_);
  xor g_104800_(out[249], out[873], _094770_);
  xor g_104801_(out[244], out[868], _094771_);
  xor g_104802_(out[242], out[866], _094772_);
  and g_104803_(out[251], _049763_, _094773_);
  xor g_104804_(out[243], out[867], _094774_);
  xor g_104805_(out[246], out[870], _094775_);
  xor g_104806_(out[255], out[879], _094776_);
  xor g_104807_(out[250], out[874], _094777_);
  xor g_104808_(out[245], out[869], _094778_);
  xor g_104809_(out[240], out[864], _094779_);
  or g_104810_(_094766_, _094771_, _094780_);
  or g_104811_(_094767_, _094769_, _094781_);
  or g_104812_(_094772_, _094777_, _094782_);
  or g_104813_(_094781_, _094782_, _094783_);
  or g_104814_(_094770_, _094774_, _094784_);
  or g_104815_(_094778_, _094779_, _094785_);
  or g_104816_(_094784_, _094785_, _094786_);
  or g_104817_(_094783_, _094786_, _094787_);
  xor g_104818_(out[252], out[876], _094788_);
  or g_104819_(_094765_, _094788_, _094789_);
  or g_104820_(_094764_, _094775_, _094790_);
  or g_104821_(_094789_, _094790_, _094791_);
  or g_104822_(_094768_, _094773_, _094792_);
  or g_104823_(_094776_, _094792_, _094793_);
  or g_104824_(_094791_, _094793_, _094794_);
  or g_104825_(_094787_, _094794_, _094795_);
  or g_104826_(_094780_, _094795_, _094796_);
  xor g_104827_(out[232], out[872], _094797_);
  xor g_104828_(out[229], out[869], _094798_);
  xor g_104829_(out[227], out[867], _094799_);
  xor g_104830_(out[238], out[878], _094800_);
  xor g_104831_(out[237], out[877], _094801_);
  xor g_104832_(out[226], out[866], _094802_);
  xor g_104833_(out[233], out[873], _094803_);
  xor g_104834_(out[230], out[870], _094804_);
  xor g_104835_(out[239], out[879], _094805_);
  xor g_104836_(out[234], out[874], _094806_);
  xor g_104837_(out[228], out[868], _094807_);
  xor g_104838_(out[224], out[864], _094808_);
  and g_104839_(_098228_, out[875], _094809_);
  and g_104840_(out[235], _049763_, _094810_);
  or g_104841_(_094797_, _094801_, _094811_);
  xor g_104842_(out[225], out[865], _094812_);
  or g_104843_(_094802_, _094806_, _094813_);
  or g_104844_(_094811_, _094813_, _094814_);
  or g_104845_(_094799_, _094803_, _094815_);
  or g_104846_(_094798_, _094815_, _094816_);
  or g_104847_(_094814_, _094816_, _094817_);
  or g_104848_(_094800_, _094807_, _094818_);
  or g_104849_(_094817_, _094818_, _094819_);
  xor g_104850_(out[236], out[876], _094820_);
  or g_104851_(_094809_, _094820_, _094821_);
  xor g_104852_(out[231], out[871], _094822_);
  or g_104853_(_094804_, _094822_, _094823_);
  or g_104854_(_094821_, _094823_, _094824_);
  or g_104855_(_094810_, _094812_, _094825_);
  or g_104856_(_094805_, _094825_, _094826_);
  or g_104857_(_094824_, _094826_, _094827_);
  or g_104858_(_094808_, _094827_, _094828_);
  or g_104859_(_094819_, _094828_, _094829_);
  not g_104860_(_094829_, _094830_);
  xor g_104861_(out[215], out[871], _094831_);
  and g_104862_(_098217_, out[875], _094832_);
  xor g_104863_(out[222], out[878], _094833_);
  xor g_104864_(out[216], out[872], _094834_);
  xor g_104865_(out[209], out[865], _094835_);
  xor g_104866_(out[221], out[877], _094836_);
  xor g_104867_(out[217], out[873], _094837_);
  xor g_104868_(out[212], out[868], _094838_);
  xor g_104869_(out[210], out[866], _094839_);
  and g_104870_(out[219], _049763_, _094840_);
  xor g_104871_(out[211], out[867], _094841_);
  xor g_104872_(out[214], out[870], _094842_);
  xor g_104873_(out[223], out[879], _094843_);
  xor g_104874_(out[218], out[874], _094844_);
  xor g_104875_(out[213], out[869], _094845_);
  xor g_104876_(out[208], out[864], _094846_);
  or g_104877_(_094833_, _094838_, _094847_);
  or g_104878_(_094834_, _094836_, _094848_);
  or g_104879_(_094839_, _094844_, _094849_);
  or g_104880_(_094848_, _094849_, _094850_);
  or g_104881_(_094837_, _094841_, _094851_);
  or g_104882_(_094845_, _094846_, _094852_);
  or g_104883_(_094851_, _094852_, _094853_);
  or g_104884_(_094850_, _094853_, _094854_);
  xor g_104885_(out[220], out[876], _094855_);
  or g_104886_(_094832_, _094855_, _094856_);
  or g_104887_(_094831_, _094842_, _094857_);
  or g_104888_(_094856_, _094857_, _094858_);
  or g_104889_(_094835_, _094840_, _094859_);
  or g_104890_(_094843_, _094859_, _094860_);
  or g_104891_(_094858_, _094860_, _094861_);
  or g_104892_(_094854_, _094861_, _094862_);
  or g_104893_(_094847_, _094862_, _094863_);
  xor g_104894_(out[204], out[876], _094864_);
  and g_104895_(_098206_, out[875], _094865_);
  xor g_104896_(out[200], out[872], _094866_);
  xor g_104897_(out[198], out[870], _094867_);
  xor g_104898_(out[205], out[877], _094868_);
  xor g_104899_(out[206], out[878], _094869_);
  xor g_104900_(out[194], out[866], _094870_);
  xor g_104901_(out[201], out[873], _094871_);
  xor g_104902_(out[197], out[869], _094872_);
  xor g_104903_(out[193], out[865], _094873_);
  and g_104904_(out[203], _049763_, _094874_);
  or g_104905_(_094866_, _094868_, _094875_);
  xor g_104906_(out[207], out[879], _094876_);
  xor g_104907_(out[202], out[874], _094877_);
  xor g_104908_(out[196], out[868], _094878_);
  xor g_104909_(out[195], out[867], _094879_);
  xor g_104910_(out[192], out[864], _094880_);
  or g_104911_(_094870_, _094877_, _094881_);
  or g_104912_(_094875_, _094881_, _094882_);
  or g_104913_(_094871_, _094879_, _094883_);
  or g_104914_(_094872_, _094883_, _094884_);
  or g_104915_(_094882_, _094884_, _094885_);
  or g_104916_(_094869_, _094878_, _094886_);
  or g_104917_(_094885_, _094886_, _094887_);
  or g_104918_(_094864_, _094865_, _094888_);
  xor g_104919_(out[199], out[871], _094889_);
  or g_104920_(_094867_, _094889_, _094890_);
  or g_104921_(_094888_, _094890_, _094891_);
  or g_104922_(_094873_, _094874_, _094892_);
  or g_104923_(_094876_, _094892_, _094893_);
  or g_104924_(_094891_, _094893_, _094894_);
  or g_104925_(_094880_, _094894_, _094895_);
  or g_104926_(_094887_, _094895_, _094896_);
  xor g_104927_(out[183], out[871], _094897_);
  and g_104928_(_098195_, out[875], _094898_);
  xor g_104929_(out[190], out[878], _094899_);
  xor g_104930_(out[184], out[872], _094900_);
  xor g_104931_(out[177], out[865], _094901_);
  xor g_104932_(out[189], out[877], _094902_);
  xor g_104933_(out[185], out[873], _094903_);
  xor g_104934_(out[180], out[868], _094904_);
  xor g_104935_(out[178], out[866], _094905_);
  and g_104936_(out[187], _049763_, _094906_);
  xor g_104937_(out[179], out[867], _094907_);
  xor g_104938_(out[182], out[870], _094908_);
  xor g_104939_(out[191], out[879], _094909_);
  xor g_104940_(out[186], out[874], _094910_);
  xor g_104941_(out[181], out[869], _094911_);
  xor g_104942_(out[176], out[864], _094912_);
  or g_104943_(_094899_, _094904_, _094913_);
  or g_104944_(_094900_, _094902_, _094914_);
  or g_104945_(_094905_, _094910_, _094915_);
  or g_104946_(_094914_, _094915_, _094916_);
  or g_104947_(_094903_, _094907_, _094917_);
  or g_104948_(_094911_, _094912_, _094918_);
  or g_104949_(_094917_, _094918_, _094919_);
  or g_104950_(_094916_, _094919_, _094920_);
  xor g_104951_(out[188], out[876], _094921_);
  or g_104952_(_094898_, _094921_, _094922_);
  or g_104953_(_094897_, _094908_, _094923_);
  or g_104954_(_094922_, _094923_, _094924_);
  or g_104955_(_094901_, _094906_, _094925_);
  or g_104956_(_094909_, _094925_, _094926_);
  or g_104957_(_094924_, _094926_, _094927_);
  or g_104958_(_094920_, _094927_, _094928_);
  or g_104959_(_094913_, _094928_, _094929_);
  not g_104960_(_094929_, _094930_);
  and g_104961_(out[171], _049763_, _094931_);
  and g_104962_(_098184_, out[875], _094932_);
  xor g_104963_(out[168], out[872], _094933_);
  xor g_104964_(out[175], out[879], _094934_);
  xor g_104965_(out[161], out[865], _094935_);
  xor g_104966_(out[162], out[866], _094936_);
  xor g_104967_(out[164], out[868], _094937_);
  xor g_104968_(out[173], out[877], _094938_);
  xor g_104969_(out[169], out[873], _094939_);
  xor g_104970_(out[163], out[867], _094940_);
  xor g_104971_(out[165], out[869], _094941_);
  xor g_104972_(out[174], out[878], _094942_);
  xor g_104973_(out[160], out[864], _094943_);
  xor g_104974_(out[170], out[874], _094944_);
  or g_104975_(_094933_, _094938_, _094945_);
  xor g_104976_(out[166], out[870], _094946_);
  or g_104977_(_094936_, _094944_, _094947_);
  or g_104978_(_094945_, _094947_, _094948_);
  or g_104979_(_094939_, _094940_, _094949_);
  or g_104980_(_094941_, _094949_, _094950_);
  or g_104981_(_094948_, _094950_, _094951_);
  or g_104982_(_094937_, _094942_, _094952_);
  or g_104983_(_094951_, _094952_, _094953_);
  xor g_104984_(out[172], out[876], _094954_);
  or g_104985_(_094932_, _094954_, _094955_);
  xor g_104986_(out[167], out[871], _094956_);
  or g_104987_(_094946_, _094956_, _094957_);
  or g_104988_(_094955_, _094957_, _094958_);
  or g_104989_(_094931_, _094935_, _094959_);
  or g_104990_(_094934_, _094959_, _094960_);
  or g_104991_(_094958_, _094960_, _094961_);
  or g_104992_(_094943_, _094961_, _094962_);
  or g_104993_(_094953_, _094962_, _094963_);
  not g_104994_(_094963_, _094964_);
  xor g_104995_(out[151], out[871], _094965_);
  and g_104996_(_098173_, out[875], _094966_);
  xor g_104997_(out[158], out[878], _094967_);
  xor g_104998_(out[152], out[872], _094968_);
  xor g_104999_(out[145], out[865], _094969_);
  xor g_105000_(out[157], out[877], _094970_);
  xor g_105001_(out[153], out[873], _094971_);
  xor g_105002_(out[148], out[868], _094972_);
  xor g_105003_(out[146], out[866], _094973_);
  and g_105004_(out[155], _049763_, _094974_);
  xor g_105005_(out[147], out[867], _094975_);
  xor g_105006_(out[150], out[870], _094976_);
  xor g_105007_(out[159], out[879], _094977_);
  xor g_105008_(out[154], out[874], _094978_);
  xor g_105009_(out[149], out[869], _094979_);
  xor g_105010_(out[144], out[864], _094980_);
  or g_105011_(_094967_, _094972_, _094981_);
  or g_105012_(_094968_, _094970_, _094982_);
  or g_105013_(_094973_, _094978_, _094983_);
  or g_105014_(_094982_, _094983_, _094984_);
  or g_105015_(_094971_, _094975_, _094985_);
  or g_105016_(_094979_, _094980_, _094986_);
  or g_105017_(_094985_, _094986_, _094987_);
  or g_105018_(_094984_, _094987_, _094988_);
  xor g_105019_(out[156], out[876], _094989_);
  or g_105020_(_094966_, _094989_, _094990_);
  or g_105021_(_094965_, _094976_, _094991_);
  or g_105022_(_094990_, _094991_, _094992_);
  or g_105023_(_094969_, _094974_, _094993_);
  or g_105024_(_094977_, _094993_, _094994_);
  or g_105025_(_094992_, _094994_, _094995_);
  or g_105026_(_094988_, _094995_, _094996_);
  or g_105027_(_094981_, _094996_, _094997_);
  xor g_105028_(out[138], out[874], _094998_);
  xor g_105029_(out[130], out[866], _094999_);
  xor g_105030_(out[129], out[865], _095000_);
  and g_105031_(_098162_, out[875], _095001_);
  and g_105032_(out[139], _049763_, _095002_);
  xor g_105033_(out[141], out[877], _095003_);
  xor g_105034_(out[131], out[867], _095004_);
  xor g_105035_(out[142], out[878], _095005_);
  xor g_105036_(out[140], out[876], _095006_);
  xor g_105037_(out[136], out[872], _095007_);
  xor g_105038_(out[143], out[879], _095008_);
  xor g_105039_(out[133], out[869], _095009_);
  xor g_105040_(out[134], out[870], _095010_);
  xor g_105041_(out[128], out[864], _095011_);
  xor g_105042_(out[132], out[868], _095012_);
  or g_105043_(_095003_, _095007_, _095013_);
  xor g_105044_(out[137], out[873], _095014_);
  or g_105045_(_094998_, _094999_, _095015_);
  or g_105046_(_095013_, _095015_, _095016_);
  or g_105047_(_095004_, _095014_, _095017_);
  or g_105048_(_095009_, _095017_, _095018_);
  or g_105049_(_095016_, _095018_, _095019_);
  or g_105050_(_095005_, _095012_, _095020_);
  or g_105051_(_095019_, _095020_, _095021_);
  or g_105052_(_095001_, _095006_, _095022_);
  xor g_105053_(out[135], out[871], _095023_);
  or g_105054_(_095010_, _095023_, _095024_);
  or g_105055_(_095022_, _095024_, _095025_);
  or g_105056_(_095000_, _095002_, _095026_);
  or g_105057_(_095008_, _095026_, _095027_);
  or g_105058_(_095025_, _095027_, _095028_);
  or g_105059_(_095011_, _095028_, _095029_);
  or g_105060_(_095021_, _095029_, _095030_);
  xor g_105061_(out[119], out[871], _095031_);
  and g_105062_(_098151_, out[875], _095032_);
  xor g_105063_(out[126], out[878], _095033_);
  xor g_105064_(out[120], out[872], _095034_);
  xor g_105065_(out[113], out[865], _095035_);
  xor g_105066_(out[125], out[877], _095036_);
  xor g_105067_(out[121], out[873], _095037_);
  xor g_105068_(out[116], out[868], _095038_);
  xor g_105069_(out[114], out[866], _095039_);
  and g_105070_(out[123], _049763_, _095040_);
  xor g_105071_(out[115], out[867], _095041_);
  xor g_105072_(out[118], out[870], _095042_);
  xor g_105073_(out[127], out[879], _095043_);
  xor g_105074_(out[122], out[874], _095044_);
  xor g_105075_(out[117], out[869], _095045_);
  xor g_105076_(out[112], out[864], _095046_);
  or g_105077_(_095033_, _095038_, _095047_);
  or g_105078_(_095034_, _095036_, _095048_);
  or g_105079_(_095039_, _095044_, _095049_);
  or g_105080_(_095048_, _095049_, _095050_);
  or g_105081_(_095037_, _095041_, _095051_);
  or g_105082_(_095045_, _095046_, _095052_);
  or g_105083_(_095051_, _095052_, _095053_);
  or g_105084_(_095050_, _095053_, _095054_);
  xor g_105085_(out[124], out[876], _095055_);
  or g_105086_(_095032_, _095055_, _095056_);
  or g_105087_(_095031_, _095042_, _095057_);
  or g_105088_(_095056_, _095057_, _095058_);
  or g_105089_(_095035_, _095040_, _095059_);
  or g_105090_(_095043_, _095059_, _095060_);
  or g_105091_(_095058_, _095060_, _095061_);
  or g_105092_(_095054_, _095061_, _095062_);
  or g_105093_(_095047_, _095062_, _095063_);
  xor g_105094_(out[98], out[866], _095064_);
  xor g_105095_(out[96], out[864], _095065_);
  xor g_105096_(out[105], out[873], _095066_);
  xor g_105097_(out[104], out[872], _095067_);
  xor g_105098_(out[101], out[869], _095068_);
  xor g_105099_(out[110], out[878], _095069_);
  xor g_105100_(out[109], out[877], _095070_);
  xor g_105101_(out[111], out[879], _095071_);
  xor g_105102_(out[106], out[874], _095072_);
  xor g_105103_(out[102], out[870], _095073_);
  xor g_105104_(out[99], out[867], _095074_);
  and g_105105_(_098140_, out[875], _095075_);
  and g_105106_(out[107], _049763_, _095076_);
  xor g_105107_(out[100], out[868], _095077_);
  xor g_105108_(out[97], out[865], _095078_);
  or g_105109_(_095069_, _095077_, _095079_);
  or g_105110_(_095067_, _095070_, _095080_);
  or g_105111_(_095064_, _095072_, _095081_);
  or g_105112_(_095080_, _095081_, _095082_);
  or g_105113_(_095066_, _095074_, _095083_);
  or g_105114_(_095065_, _095068_, _095084_);
  or g_105115_(_095083_, _095084_, _095085_);
  or g_105116_(_095082_, _095085_, _095086_);
  xor g_105117_(out[108], out[876], _095087_);
  or g_105118_(_095075_, _095087_, _095088_);
  xor g_105119_(out[103], out[871], _095089_);
  or g_105120_(_095073_, _095089_, _095090_);
  or g_105121_(_095088_, _095090_, _095091_);
  or g_105122_(_095076_, _095078_, _095092_);
  or g_105123_(_095071_, _095092_, _095093_);
  or g_105124_(_095091_, _095093_, _095094_);
  or g_105125_(_095086_, _095094_, _095095_);
  or g_105126_(_095079_, _095095_, _095096_);
  xor g_105127_(out[87], out[871], _095097_);
  and g_105128_(_098129_, out[875], _095098_);
  xor g_105129_(out[94], out[878], _095099_);
  xor g_105130_(out[88], out[872], _095100_);
  xor g_105131_(out[81], out[865], _095101_);
  xor g_105132_(out[93], out[877], _095102_);
  xor g_105133_(out[89], out[873], _095103_);
  xor g_105134_(out[84], out[868], _095104_);
  xor g_105135_(out[82], out[866], _095105_);
  and g_105136_(out[91], _049763_, _095106_);
  xor g_105137_(out[83], out[867], _095107_);
  xor g_105138_(out[86], out[870], _095108_);
  xor g_105139_(out[95], out[879], _095109_);
  xor g_105140_(out[90], out[874], _095110_);
  xor g_105141_(out[85], out[869], _095111_);
  xor g_105142_(out[80], out[864], _095112_);
  or g_105143_(_095099_, _095104_, _095113_);
  or g_105144_(_095100_, _095102_, _095114_);
  or g_105145_(_095105_, _095110_, _095115_);
  or g_105146_(_095114_, _095115_, _095116_);
  or g_105147_(_095103_, _095107_, _095117_);
  or g_105148_(_095111_, _095112_, _095118_);
  or g_105149_(_095117_, _095118_, _095119_);
  or g_105150_(_095116_, _095119_, _095120_);
  xor g_105151_(out[92], out[876], _095121_);
  or g_105152_(_095098_, _095121_, _095122_);
  or g_105153_(_095097_, _095108_, _095123_);
  or g_105154_(_095122_, _095123_, _095124_);
  or g_105155_(_095101_, _095106_, _095125_);
  or g_105156_(_095109_, _095125_, _095126_);
  or g_105157_(_095124_, _095126_, _095127_);
  or g_105158_(_095120_, _095127_, _095128_);
  or g_105159_(_095113_, _095128_, _095129_);
  not g_105160_(_095129_, _095130_);
  xor g_105161_(out[72], out[872], _095131_);
  xor g_105162_(out[69], out[869], _095132_);
  xor g_105163_(out[67], out[867], _095133_);
  xor g_105164_(out[78], out[878], _095134_);
  xor g_105165_(out[77], out[877], _095135_);
  xor g_105166_(out[66], out[866], _095136_);
  xor g_105167_(out[73], out[873], _095137_);
  xor g_105168_(out[70], out[870], _095138_);
  xor g_105169_(out[79], out[879], _095139_);
  xor g_105170_(out[74], out[874], _095140_);
  xor g_105171_(out[68], out[868], _095141_);
  xor g_105172_(out[64], out[864], _095142_);
  and g_105173_(_098118_, out[875], _095143_);
  and g_105174_(out[75], _049763_, _095144_);
  or g_105175_(_095131_, _095135_, _095145_);
  xor g_105176_(out[65], out[865], _095146_);
  or g_105177_(_095136_, _095140_, _095147_);
  or g_105178_(_095145_, _095147_, _095148_);
  or g_105179_(_095133_, _095137_, _095149_);
  or g_105180_(_095132_, _095149_, _095150_);
  or g_105181_(_095148_, _095150_, _095151_);
  or g_105182_(_095134_, _095141_, _095152_);
  or g_105183_(_095151_, _095152_, _095153_);
  xor g_105184_(out[76], out[876], _095154_);
  or g_105185_(_095143_, _095154_, _095155_);
  xor g_105186_(out[71], out[871], _095156_);
  or g_105187_(_095138_, _095156_, _095157_);
  or g_105188_(_095155_, _095157_, _095158_);
  or g_105189_(_095144_, _095146_, _095159_);
  or g_105190_(_095139_, _095159_, _095160_);
  or g_105191_(_095158_, _095160_, _095161_);
  or g_105192_(_095142_, _095161_, _095162_);
  or g_105193_(_095153_, _095162_, _095163_);
  not g_105194_(_095163_, _095164_);
  xor g_105195_(out[55], out[871], _095165_);
  and g_105196_(_098107_, out[875], _095166_);
  xor g_105197_(out[62], out[878], _095167_);
  xor g_105198_(out[56], out[872], _095168_);
  xor g_105199_(out[49], out[865], _095169_);
  xor g_105200_(out[61], out[877], _095170_);
  xor g_105201_(out[57], out[873], _095171_);
  xor g_105202_(out[52], out[868], _095172_);
  xor g_105203_(out[50], out[866], _095173_);
  and g_105204_(out[59], _049763_, _095174_);
  xor g_105205_(out[51], out[867], _095175_);
  xor g_105206_(out[54], out[870], _095176_);
  xor g_105207_(out[63], out[879], _095177_);
  xor g_105208_(out[58], out[874], _095178_);
  xor g_105209_(out[53], out[869], _095179_);
  xor g_105210_(out[48], out[864], _095180_);
  or g_105211_(_095167_, _095172_, _095181_);
  or g_105212_(_095168_, _095170_, _095182_);
  or g_105213_(_095173_, _095178_, _095183_);
  or g_105214_(_095182_, _095183_, _095184_);
  or g_105215_(_095171_, _095175_, _095185_);
  or g_105216_(_095179_, _095180_, _095186_);
  or g_105217_(_095185_, _095186_, _095187_);
  or g_105218_(_095184_, _095187_, _095188_);
  xor g_105219_(out[60], out[876], _095189_);
  or g_105220_(_095166_, _095189_, _095190_);
  or g_105221_(_095165_, _095176_, _095191_);
  or g_105222_(_095190_, _095191_, _095192_);
  or g_105223_(_095169_, _095174_, _095193_);
  or g_105224_(_095177_, _095193_, _095194_);
  or g_105225_(_095192_, _095194_, _095195_);
  or g_105226_(_095188_, _095195_, _095196_);
  or g_105227_(_095181_, _095196_, _095197_);
  not g_105228_(_095197_, _095198_);
  and g_105229_(_098096_, out[875], _095199_);
  and g_105230_(out[43], _049763_, _095200_);
  xor g_105231_(out[36], out[868], _095201_);
  xor g_105232_(out[46], out[878], _095202_);
  or g_105233_(_095201_, _095202_, _095203_);
  xor g_105234_(out[45], out[877], _095204_);
  xor g_105235_(out[35], out[867], _095205_);
  xor g_105236_(out[32], out[864], _095206_);
  xor g_105237_(out[42], out[874], _095207_);
  xor g_105238_(out[47], out[879], _095208_);
  xor g_105239_(out[38], out[870], _095209_);
  xor g_105240_(out[37], out[869], _095210_);
  xor g_105241_(out[40], out[872], _095211_);
  or g_105242_(_095204_, _095211_, _095212_);
  xor g_105243_(out[34], out[866], _095213_);
  xor g_105244_(out[41], out[873], _095214_);
  xor g_105245_(out[33], out[865], _095215_);
  or g_105246_(_095207_, _095213_, _095216_);
  or g_105247_(_095212_, _095216_, _095217_);
  or g_105248_(_095205_, _095214_, _095218_);
  or g_105249_(_095210_, _095218_, _095219_);
  or g_105250_(_095217_, _095219_, _095220_);
  or g_105251_(_095203_, _095220_, _095221_);
  xor g_105252_(out[44], out[876], _095222_);
  or g_105253_(_095199_, _095222_, _095223_);
  xor g_105254_(out[39], out[871], _095224_);
  or g_105255_(_095209_, _095224_, _095225_);
  or g_105256_(_095223_, _095225_, _095226_);
  or g_105257_(_095200_, _095215_, _095227_);
  or g_105258_(_095208_, _095227_, _095228_);
  or g_105259_(_095226_, _095228_, _095229_);
  or g_105260_(_095206_, _095229_, _095230_);
  or g_105261_(_095221_, _095230_, _095231_);
  xor g_105262_(out[23], out[871], _095232_);
  and g_105263_(_098063_, out[875], _095233_);
  xor g_105264_(out[30], out[878], _095234_);
  xor g_105265_(out[24], out[872], _095235_);
  xor g_105266_(out[17], out[865], _095236_);
  xor g_105267_(out[29], out[877], _095237_);
  xor g_105268_(out[25], out[873], _095238_);
  xor g_105269_(out[20], out[868], _095239_);
  xor g_105270_(out[18], out[866], _095240_);
  and g_105271_(out[27], _049763_, _095241_);
  xor g_105272_(out[19], out[867], _095242_);
  xor g_105273_(out[22], out[870], _095243_);
  xor g_105274_(out[31], out[879], _095244_);
  xor g_105275_(out[26], out[874], _095245_);
  xor g_105276_(out[21], out[869], _095246_);
  xor g_105277_(out[16], out[864], _095247_);
  or g_105278_(_095234_, _095239_, _095248_);
  or g_105279_(_095235_, _095237_, _095249_);
  or g_105280_(_095240_, _095245_, _095250_);
  or g_105281_(_095249_, _095250_, _095251_);
  or g_105282_(_095238_, _095242_, _095252_);
  or g_105283_(_095246_, _095247_, _095253_);
  or g_105284_(_095252_, _095253_, _095254_);
  or g_105285_(_095251_, _095254_, _095255_);
  xor g_105286_(out[28], out[876], _095256_);
  or g_105287_(_095233_, _095256_, _095257_);
  or g_105288_(_095232_, _095243_, _095258_);
  or g_105289_(_095257_, _095258_, _095259_);
  or g_105290_(_095236_, _095241_, _095260_);
  or g_105291_(_095244_, _095260_, _095261_);
  or g_105292_(_095259_, _095261_, _095262_);
  or g_105293_(_095255_, _095262_, _095263_);
  or g_105294_(_095248_, _095263_, _095264_);
  xor g_105295_(out[10], out[874], _095265_);
  xor g_105296_(out[8], out[872], _095266_);
  xor g_105297_(out[1], out[865], _095267_);
  and g_105298_(_098041_, out[875], _095268_);
  and g_105299_(out[11], _049763_, _095269_);
  xor g_105300_(out[2], out[866], _095270_);
  xor g_105301_(out[5], out[869], _095271_);
  xor g_105302_(out[9], out[873], _095272_);
  xor g_105303_(out[12], out[876], _095273_);
  xor g_105304_(out[13], out[877], _095274_);
  xor g_105305_(out[15], out[879], _095275_);
  xor g_105306_(out[4], out[868], _095276_);
  xor g_105307_(out[6], out[870], _095277_);
  xor g_105308_(out[3], out[867], _095278_);
  xor g_105309_(out[0], out[864], _095279_);
  xor g_105310_(out[14], out[878], _095280_);
  or g_105311_(_095276_, _095280_, _095281_);
  or g_105312_(_095266_, _095274_, _095282_);
  or g_105313_(_095265_, _095270_, _095283_);
  or g_105314_(_095282_, _095283_, _095284_);
  or g_105315_(_095272_, _095278_, _095285_);
  or g_105316_(_095271_, _095279_, _095286_);
  or g_105317_(_095285_, _095286_, _095287_);
  or g_105318_(_095284_, _095287_, _095288_);
  or g_105319_(_095268_, _095273_, _095289_);
  xor g_105320_(out[7], out[871], _095290_);
  or g_105321_(_095277_, _095290_, _095291_);
  or g_105322_(_095289_, _095291_, _095292_);
  or g_105323_(_095267_, _095269_, _095293_);
  or g_105324_(_095275_, _095293_, _095294_);
  or g_105325_(_095292_, _095294_, _095295_);
  or g_105326_(_095288_, _095295_, _095296_);
  or g_105327_(_095281_, _095296_, _095297_);
  not g_105328_(_095297_, _095298_);
  xor g_105329_(out[472], out[856], _095299_);
  xor g_105330_(out[469], out[853], _095300_);
  xor g_105331_(out[467], out[851], _095301_);
  xor g_105332_(out[478], out[862], _095302_);
  xor g_105333_(out[477], out[861], _095303_);
  xor g_105334_(out[466], out[850], _095304_);
  xor g_105335_(out[473], out[857], _095305_);
  xor g_105336_(out[470], out[854], _095306_);
  xor g_105337_(out[479], out[863], _095307_);
  xor g_105338_(out[474], out[858], _095308_);
  xor g_105339_(out[468], out[852], _095309_);
  xor g_105340_(out[464], out[848], _095310_);
  and g_105341_(_049499_, out[859], _095311_);
  and g_105342_(out[475], _049752_, _095312_);
  or g_105343_(_095299_, _095303_, _095313_);
  xor g_105344_(out[465], out[849], _095314_);
  or g_105345_(_095304_, _095308_, _095315_);
  or g_105346_(_095313_, _095315_, _095316_);
  or g_105347_(_095301_, _095305_, _095317_);
  or g_105348_(_095300_, _095317_, _095318_);
  or g_105349_(_095316_, _095318_, _095319_);
  or g_105350_(_095302_, _095309_, _095320_);
  or g_105351_(_095319_, _095320_, _095321_);
  xor g_105352_(out[476], out[860], _095322_);
  or g_105353_(_095311_, _095322_, _095323_);
  xor g_105354_(out[471], out[855], _095324_);
  or g_105355_(_095306_, _095324_, _095325_);
  or g_105356_(_095323_, _095325_, _095326_);
  or g_105357_(_095312_, _095314_, _095327_);
  or g_105358_(_095307_, _095327_, _095328_);
  or g_105359_(_095326_, _095328_, _095329_);
  or g_105360_(_095310_, _095329_, _095330_);
  or g_105361_(_095321_, _095330_, _095331_);
  not g_105362_(_095331_, _095332_);
  xor g_105363_(out[455], out[855], _095333_);
  and g_105364_(_049477_, out[859], _095334_);
  xor g_105365_(out[462], out[862], _095335_);
  xor g_105366_(out[456], out[856], _095336_);
  xor g_105367_(out[449], out[849], _095337_);
  xor g_105368_(out[461], out[861], _095338_);
  xor g_105369_(out[457], out[857], _095339_);
  xor g_105370_(out[452], out[852], _095340_);
  xor g_105371_(out[450], out[850], _095341_);
  and g_105372_(out[459], _049752_, _095342_);
  xor g_105373_(out[451], out[851], _095343_);
  xor g_105374_(out[454], out[854], _095344_);
  xor g_105375_(out[463], out[863], _095345_);
  xor g_105376_(out[458], out[858], _095346_);
  xor g_105377_(out[453], out[853], _095347_);
  xor g_105378_(out[448], out[848], _095348_);
  or g_105379_(_095335_, _095340_, _095349_);
  or g_105380_(_095336_, _095338_, _095350_);
  or g_105381_(_095341_, _095346_, _095351_);
  or g_105382_(_095350_, _095351_, _095352_);
  or g_105383_(_095339_, _095343_, _095353_);
  or g_105384_(_095347_, _095348_, _095354_);
  or g_105385_(_095353_, _095354_, _095355_);
  or g_105386_(_095352_, _095355_, _095356_);
  xor g_105387_(out[460], out[860], _095357_);
  or g_105388_(_095334_, _095357_, _095358_);
  or g_105389_(_095333_, _095344_, _095359_);
  or g_105390_(_095358_, _095359_, _095360_);
  or g_105391_(_095337_, _095342_, _095361_);
  or g_105392_(_095345_, _095361_, _095362_);
  or g_105393_(_095360_, _095362_, _095363_);
  or g_105394_(_095356_, _095363_, _095364_);
  or g_105395_(_095349_, _095364_, _095365_);
  not g_105396_(_095365_, _095366_);
  xor g_105397_(out[433], out[849], _095367_);
  and g_105398_(out[443], _049752_, _095368_);
  xor g_105399_(out[441], out[857], _095369_);
  xor g_105400_(out[432], out[848], _095370_);
  xor g_105401_(out[446], out[862], _095371_);
  xor g_105402_(out[436], out[852], _095372_);
  or g_105403_(_095371_, _095372_, _095373_);
  xor g_105404_(out[445], out[861], _095374_);
  xor g_105405_(out[435], out[851], _095375_);
  and g_105406_(_049466_, out[859], _095376_);
  xor g_105407_(out[438], out[854], _095377_);
  xor g_105408_(out[442], out[858], _095378_);
  xor g_105409_(out[437], out[853], _095379_);
  xor g_105410_(out[447], out[863], _095380_);
  xor g_105411_(out[440], out[856], _095381_);
  or g_105412_(_095374_, _095381_, _095382_);
  xor g_105413_(out[434], out[850], _095383_);
  or g_105414_(_095378_, _095383_, _095384_);
  or g_105415_(_095382_, _095384_, _095385_);
  or g_105416_(_095369_, _095375_, _095386_);
  or g_105417_(_095379_, _095386_, _095387_);
  or g_105418_(_095385_, _095387_, _095388_);
  or g_105419_(_095373_, _095388_, _095389_);
  xor g_105420_(out[444], out[860], _095390_);
  or g_105421_(_095376_, _095390_, _095391_);
  xor g_105422_(out[439], out[855], _095392_);
  or g_105423_(_095377_, _095392_, _095393_);
  or g_105424_(_095391_, _095393_, _095394_);
  or g_105425_(_095367_, _095368_, _095395_);
  or g_105426_(_095380_, _095395_, _095396_);
  or g_105427_(_095394_, _095396_, _095397_);
  or g_105428_(_095370_, _095397_, _095398_);
  or g_105429_(_095389_, _095398_, _095399_);
  xor g_105430_(out[423], out[855], _095400_);
  and g_105431_(_049455_, out[859], _095401_);
  xor g_105432_(out[430], out[862], _095402_);
  xor g_105433_(out[424], out[856], _095403_);
  xor g_105434_(out[417], out[849], _095404_);
  xor g_105435_(out[429], out[861], _095405_);
  xor g_105436_(out[425], out[857], _095406_);
  xor g_105437_(out[420], out[852], _095407_);
  xor g_105438_(out[418], out[850], _095408_);
  and g_105439_(out[427], _049752_, _095409_);
  xor g_105440_(out[419], out[851], _095410_);
  xor g_105441_(out[422], out[854], _095411_);
  xor g_105442_(out[431], out[863], _095412_);
  xor g_105443_(out[426], out[858], _095413_);
  xor g_105444_(out[421], out[853], _095414_);
  xor g_105445_(out[416], out[848], _095415_);
  or g_105446_(_095402_, _095407_, _095416_);
  or g_105447_(_095403_, _095405_, _095417_);
  or g_105448_(_095408_, _095413_, _095418_);
  or g_105449_(_095417_, _095418_, _095419_);
  or g_105450_(_095406_, _095410_, _095420_);
  or g_105451_(_095414_, _095415_, _095421_);
  or g_105452_(_095420_, _095421_, _095422_);
  or g_105453_(_095419_, _095422_, _095423_);
  xor g_105454_(out[428], out[860], _095424_);
  or g_105455_(_095401_, _095424_, _095425_);
  or g_105456_(_095400_, _095411_, _095426_);
  or g_105457_(_095425_, _095426_, _095427_);
  or g_105458_(_095404_, _095409_, _095428_);
  or g_105459_(_095412_, _095428_, _095429_);
  or g_105460_(_095427_, _095429_, _095430_);
  or g_105461_(_095423_, _095430_, _095431_);
  or g_105462_(_095416_, _095431_, _095432_);
  xor g_105463_(out[401], out[849], _095433_);
  and g_105464_(out[411], _049752_, _095434_);
  xor g_105465_(out[409], out[857], _095435_);
  xor g_105466_(out[400], out[848], _095436_);
  xor g_105467_(out[414], out[862], _095437_);
  xor g_105468_(out[404], out[852], _095438_);
  or g_105469_(_095437_, _095438_, _095439_);
  xor g_105470_(out[413], out[861], _095440_);
  xor g_105471_(out[403], out[851], _095441_);
  and g_105472_(_049444_, out[859], _095442_);
  xor g_105473_(out[406], out[854], _095443_);
  xor g_105474_(out[410], out[858], _095444_);
  xor g_105475_(out[405], out[853], _095445_);
  xor g_105476_(out[415], out[863], _095446_);
  xor g_105477_(out[408], out[856], _095447_);
  or g_105478_(_095440_, _095447_, _095448_);
  xor g_105479_(out[402], out[850], _095449_);
  or g_105480_(_095444_, _095449_, _095450_);
  or g_105481_(_095448_, _095450_, _095451_);
  or g_105482_(_095435_, _095441_, _095452_);
  or g_105483_(_095445_, _095452_, _095453_);
  or g_105484_(_095451_, _095453_, _095454_);
  or g_105485_(_095439_, _095454_, _095455_);
  xor g_105486_(out[412], out[860], _095456_);
  or g_105487_(_095442_, _095456_, _095457_);
  xor g_105488_(out[407], out[855], _095458_);
  or g_105489_(_095443_, _095458_, _095459_);
  or g_105490_(_095457_, _095459_, _095460_);
  or g_105491_(_095433_, _095434_, _095461_);
  or g_105492_(_095446_, _095461_, _095462_);
  or g_105493_(_095460_, _095462_, _095463_);
  or g_105494_(_095436_, _095463_, _095464_);
  or g_105495_(_095455_, _095464_, _095465_);
  xor g_105496_(out[391], out[855], _095466_);
  and g_105497_(_049433_, out[859], _095467_);
  xor g_105498_(out[398], out[862], _095468_);
  xor g_105499_(out[392], out[856], _095469_);
  xor g_105500_(out[385], out[849], _095470_);
  xor g_105501_(out[397], out[861], _095471_);
  xor g_105502_(out[393], out[857], _095472_);
  xor g_105503_(out[388], out[852], _095473_);
  xor g_105504_(out[386], out[850], _095474_);
  and g_105505_(out[395], _049752_, _095475_);
  xor g_105506_(out[387], out[851], _095476_);
  xor g_105507_(out[390], out[854], _095477_);
  xor g_105508_(out[399], out[863], _095478_);
  xor g_105509_(out[394], out[858], _095479_);
  xor g_105510_(out[389], out[853], _095480_);
  xor g_105511_(out[384], out[848], _095481_);
  or g_105512_(_095468_, _095473_, _095482_);
  or g_105513_(_095469_, _095471_, _095483_);
  or g_105514_(_095474_, _095479_, _095484_);
  or g_105515_(_095483_, _095484_, _095485_);
  or g_105516_(_095472_, _095476_, _095486_);
  or g_105517_(_095480_, _095481_, _095487_);
  or g_105518_(_095486_, _095487_, _095488_);
  or g_105519_(_095485_, _095488_, _095489_);
  xor g_105520_(out[396], out[860], _095490_);
  or g_105521_(_095467_, _095490_, _095491_);
  or g_105522_(_095466_, _095477_, _095492_);
  or g_105523_(_095491_, _095492_, _095493_);
  or g_105524_(_095470_, _095475_, _095494_);
  or g_105525_(_095478_, _095494_, _095495_);
  or g_105526_(_095493_, _095495_, _095496_);
  or g_105527_(_095489_, _095496_, _095497_);
  or g_105528_(_095482_, _095497_, _095498_);
  xor g_105529_(out[380], out[860], _095499_);
  and g_105530_(_049422_, out[859], _095500_);
  xor g_105531_(out[376], out[856], _095501_);
  xor g_105532_(out[374], out[854], _095502_);
  xor g_105533_(out[381], out[861], _095503_);
  xor g_105534_(out[382], out[862], _095504_);
  xor g_105535_(out[370], out[850], _095505_);
  xor g_105536_(out[377], out[857], _095506_);
  xor g_105537_(out[373], out[853], _095507_);
  xor g_105538_(out[369], out[849], _095508_);
  and g_105539_(out[379], _049752_, _095509_);
  or g_105540_(_095501_, _095503_, _095510_);
  xor g_105541_(out[383], out[863], _095511_);
  xor g_105542_(out[378], out[858], _095512_);
  xor g_105543_(out[372], out[852], _095513_);
  xor g_105544_(out[371], out[851], _095514_);
  xor g_105545_(out[368], out[848], _095515_);
  or g_105546_(_095505_, _095512_, _095516_);
  or g_105547_(_095510_, _095516_, _095517_);
  or g_105548_(_095506_, _095514_, _095518_);
  or g_105549_(_095507_, _095518_, _095519_);
  or g_105550_(_095517_, _095519_, _095520_);
  or g_105551_(_095504_, _095513_, _095521_);
  or g_105552_(_095520_, _095521_, _095522_);
  or g_105553_(_095499_, _095500_, _095523_);
  xor g_105554_(out[375], out[855], _095524_);
  or g_105555_(_095502_, _095524_, _095525_);
  or g_105556_(_095523_, _095525_, _095526_);
  or g_105557_(_095508_, _095509_, _095527_);
  or g_105558_(_095511_, _095527_, _095528_);
  or g_105559_(_095526_, _095528_, _095529_);
  or g_105560_(_095515_, _095529_, _095530_);
  or g_105561_(_095522_, _095530_, _095531_);
  not g_105562_(_095531_, _095532_);
  xor g_105563_(out[359], out[855], _095533_);
  and g_105564_(_049411_, out[859], _095534_);
  xor g_105565_(out[366], out[862], _095535_);
  xor g_105566_(out[360], out[856], _095536_);
  xor g_105567_(out[353], out[849], _095537_);
  xor g_105568_(out[365], out[861], _095538_);
  xor g_105569_(out[361], out[857], _095539_);
  xor g_105570_(out[356], out[852], _095540_);
  xor g_105571_(out[354], out[850], _095541_);
  and g_105572_(out[363], _049752_, _095542_);
  xor g_105573_(out[355], out[851], _095543_);
  xor g_105574_(out[358], out[854], _095544_);
  xor g_105575_(out[367], out[863], _095545_);
  xor g_105576_(out[362], out[858], _095546_);
  xor g_105577_(out[357], out[853], _095547_);
  xor g_105578_(out[352], out[848], _095548_);
  or g_105579_(_095535_, _095540_, _095549_);
  or g_105580_(_095536_, _095538_, _095550_);
  or g_105581_(_095541_, _095546_, _095551_);
  or g_105582_(_095550_, _095551_, _095552_);
  or g_105583_(_095539_, _095543_, _095553_);
  or g_105584_(_095547_, _095548_, _095554_);
  or g_105585_(_095553_, _095554_, _095555_);
  or g_105586_(_095552_, _095555_, _095556_);
  xor g_105587_(out[364], out[860], _095557_);
  or g_105588_(_095534_, _095557_, _095558_);
  or g_105589_(_095533_, _095544_, _095559_);
  or g_105590_(_095558_, _095559_, _095560_);
  or g_105591_(_095537_, _095542_, _095561_);
  or g_105592_(_095545_, _095561_, _095562_);
  or g_105593_(_095560_, _095562_, _095563_);
  or g_105594_(_095556_, _095563_, _095564_);
  or g_105595_(_095549_, _095564_, _095565_);
  not g_105596_(_095565_, _095566_);
  xor g_105597_(out[337], out[849], _095567_);
  and g_105598_(out[347], _049752_, _095568_);
  xor g_105599_(out[345], out[857], _095569_);
  xor g_105600_(out[336], out[848], _095570_);
  xor g_105601_(out[350], out[862], _095571_);
  xor g_105602_(out[340], out[852], _095572_);
  or g_105603_(_095571_, _095572_, _095573_);
  xor g_105604_(out[349], out[861], _095574_);
  xor g_105605_(out[339], out[851], _095575_);
  and g_105606_(_049400_, out[859], _095576_);
  xor g_105607_(out[342], out[854], _095577_);
  xor g_105608_(out[346], out[858], _095578_);
  xor g_105609_(out[341], out[853], _095579_);
  xor g_105610_(out[351], out[863], _095580_);
  xor g_105611_(out[344], out[856], _095581_);
  or g_105612_(_095574_, _095581_, _095582_);
  xor g_105613_(out[338], out[850], _095583_);
  or g_105614_(_095578_, _095583_, _095584_);
  or g_105615_(_095582_, _095584_, _095585_);
  or g_105616_(_095569_, _095575_, _095586_);
  or g_105617_(_095579_, _095586_, _095587_);
  or g_105618_(_095585_, _095587_, _095588_);
  or g_105619_(_095573_, _095588_, _095589_);
  xor g_105620_(out[348], out[860], _095590_);
  or g_105621_(_095576_, _095590_, _095591_);
  xor g_105622_(out[343], out[855], _095592_);
  or g_105623_(_095577_, _095592_, _095593_);
  or g_105624_(_095591_, _095593_, _095594_);
  or g_105625_(_095567_, _095568_, _095595_);
  or g_105626_(_095580_, _095595_, _095596_);
  or g_105627_(_095594_, _095596_, _095597_);
  or g_105628_(_095570_, _095597_, _095598_);
  or g_105629_(_095589_, _095598_, _095599_);
  xor g_105630_(out[327], out[855], _095600_);
  and g_105631_(_098294_, out[859], _095601_);
  xor g_105632_(out[334], out[862], _095602_);
  xor g_105633_(out[328], out[856], _095603_);
  xor g_105634_(out[321], out[849], _095604_);
  xor g_105635_(out[333], out[861], _095605_);
  xor g_105636_(out[329], out[857], _095606_);
  xor g_105637_(out[324], out[852], _095607_);
  xor g_105638_(out[322], out[850], _095608_);
  and g_105639_(out[331], _049752_, _095609_);
  xor g_105640_(out[323], out[851], _095610_);
  xor g_105641_(out[326], out[854], _095611_);
  xor g_105642_(out[335], out[863], _095612_);
  xor g_105643_(out[330], out[858], _095613_);
  xor g_105644_(out[325], out[853], _095614_);
  xor g_105645_(out[320], out[848], _095615_);
  or g_105646_(_095602_, _095607_, _095616_);
  or g_105647_(_095603_, _095605_, _095617_);
  or g_105648_(_095608_, _095613_, _095618_);
  or g_105649_(_095617_, _095618_, _095619_);
  or g_105650_(_095606_, _095610_, _095620_);
  or g_105651_(_095614_, _095615_, _095621_);
  or g_105652_(_095620_, _095621_, _095622_);
  or g_105653_(_095619_, _095622_, _095623_);
  xor g_105654_(out[332], out[860], _095624_);
  or g_105655_(_095601_, _095624_, _095625_);
  or g_105656_(_095600_, _095611_, _095626_);
  or g_105657_(_095625_, _095626_, _095627_);
  or g_105658_(_095604_, _095609_, _095628_);
  or g_105659_(_095612_, _095628_, _095629_);
  or g_105660_(_095627_, _095629_, _095630_);
  or g_105661_(_095623_, _095630_, _095631_);
  or g_105662_(_095616_, _095631_, _095632_);
  xor g_105663_(out[316], out[860], _095633_);
  and g_105664_(_098283_, out[859], _095634_);
  xor g_105665_(out[312], out[856], _095635_);
  xor g_105666_(out[310], out[854], _095636_);
  xor g_105667_(out[317], out[861], _095637_);
  xor g_105668_(out[318], out[862], _095638_);
  xor g_105669_(out[306], out[850], _095639_);
  xor g_105670_(out[313], out[857], _095640_);
  xor g_105671_(out[309], out[853], _095641_);
  xor g_105672_(out[305], out[849], _095642_);
  and g_105673_(out[315], _049752_, _095643_);
  or g_105674_(_095635_, _095637_, _095644_);
  xor g_105675_(out[319], out[863], _095645_);
  xor g_105676_(out[314], out[858], _095646_);
  xor g_105677_(out[308], out[852], _095647_);
  xor g_105678_(out[307], out[851], _095648_);
  xor g_105679_(out[304], out[848], _095649_);
  or g_105680_(_095639_, _095646_, _095650_);
  or g_105681_(_095644_, _095650_, _095651_);
  or g_105682_(_095640_, _095648_, _095652_);
  or g_105683_(_095641_, _095652_, _095653_);
  or g_105684_(_095651_, _095653_, _095654_);
  or g_105685_(_095638_, _095647_, _095655_);
  or g_105686_(_095654_, _095655_, _095656_);
  or g_105687_(_095633_, _095634_, _095657_);
  xor g_105688_(out[311], out[855], _095658_);
  or g_105689_(_095636_, _095658_, _095659_);
  or g_105690_(_095657_, _095659_, _095660_);
  or g_105691_(_095642_, _095643_, _095661_);
  or g_105692_(_095645_, _095661_, _095662_);
  or g_105693_(_095660_, _095662_, _095663_);
  or g_105694_(_095649_, _095663_, _095664_);
  or g_105695_(_095656_, _095664_, _095665_);
  not g_105696_(_095665_, _095666_);
  xor g_105697_(out[295], out[855], _095667_);
  and g_105698_(_098272_, out[859], _095668_);
  xor g_105699_(out[302], out[862], _095669_);
  xor g_105700_(out[296], out[856], _095670_);
  xor g_105701_(out[289], out[849], _095671_);
  xor g_105702_(out[301], out[861], _095672_);
  xor g_105703_(out[297], out[857], _095673_);
  xor g_105704_(out[292], out[852], _095674_);
  xor g_105705_(out[290], out[850], _095675_);
  and g_105706_(out[299], _049752_, _095676_);
  xor g_105707_(out[291], out[851], _095677_);
  xor g_105708_(out[294], out[854], _095678_);
  xor g_105709_(out[303], out[863], _095679_);
  xor g_105710_(out[298], out[858], _095680_);
  xor g_105711_(out[293], out[853], _095681_);
  xor g_105712_(out[288], out[848], _095682_);
  or g_105713_(_095669_, _095674_, _095683_);
  or g_105714_(_095670_, _095672_, _095684_);
  or g_105715_(_095675_, _095680_, _095685_);
  or g_105716_(_095684_, _095685_, _095686_);
  or g_105717_(_095673_, _095677_, _095687_);
  or g_105718_(_095681_, _095682_, _095688_);
  or g_105719_(_095687_, _095688_, _095689_);
  or g_105720_(_095686_, _095689_, _095690_);
  xor g_105721_(out[300], out[860], _095691_);
  or g_105722_(_095668_, _095691_, _095692_);
  or g_105723_(_095667_, _095678_, _095693_);
  or g_105724_(_095692_, _095693_, _095694_);
  or g_105725_(_095671_, _095676_, _095695_);
  or g_105726_(_095679_, _095695_, _095696_);
  or g_105727_(_095694_, _095696_, _095697_);
  or g_105728_(_095690_, _095697_, _095698_);
  or g_105729_(_095683_, _095698_, _095699_);
  xor g_105730_(out[273], out[849], _095700_);
  and g_105731_(_098261_, out[859], _095701_);
  and g_105732_(out[283], _049752_, _095702_);
  xor g_105733_(out[280], out[856], _095703_);
  xor g_105734_(out[282], out[858], _095704_);
  xor g_105735_(out[274], out[850], _095705_);
  xor g_105736_(out[276], out[852], _095706_);
  xor g_105737_(out[285], out[861], _095707_);
  xor g_105738_(out[281], out[857], _095708_);
  xor g_105739_(out[275], out[851], _095709_);
  xor g_105740_(out[277], out[853], _095710_);
  xor g_105741_(out[286], out[862], _095711_);
  xor g_105742_(out[272], out[848], _095712_);
  xor g_105743_(out[287], out[863], _095713_);
  or g_105744_(_095703_, _095707_, _095714_);
  xor g_105745_(out[278], out[854], _095715_);
  or g_105746_(_095704_, _095705_, _095716_);
  or g_105747_(_095714_, _095716_, _095717_);
  or g_105748_(_095708_, _095709_, _095718_);
  or g_105749_(_095710_, _095718_, _095719_);
  or g_105750_(_095717_, _095719_, _095720_);
  or g_105751_(_095706_, _095711_, _095721_);
  or g_105752_(_095720_, _095721_, _095722_);
  xor g_105753_(out[284], out[860], _095723_);
  or g_105754_(_095701_, _095723_, _095724_);
  xor g_105755_(out[279], out[855], _095725_);
  or g_105756_(_095715_, _095725_, _095726_);
  or g_105757_(_095724_, _095726_, _095727_);
  or g_105758_(_095700_, _095702_, _095728_);
  or g_105759_(_095713_, _095728_, _095729_);
  or g_105760_(_095727_, _095729_, _095730_);
  or g_105761_(_095712_, _095730_, _095731_);
  or g_105762_(_095722_, _095731_, _095732_);
  xor g_105763_(out[263], out[855], _095733_);
  and g_105764_(_098250_, out[859], _095734_);
  xor g_105765_(out[270], out[862], _095735_);
  xor g_105766_(out[264], out[856], _095736_);
  xor g_105767_(out[257], out[849], _095737_);
  xor g_105768_(out[269], out[861], _095738_);
  xor g_105769_(out[265], out[857], _095739_);
  xor g_105770_(out[260], out[852], _095740_);
  xor g_105771_(out[258], out[850], _095741_);
  and g_105772_(out[267], _049752_, _095742_);
  xor g_105773_(out[259], out[851], _095743_);
  xor g_105774_(out[262], out[854], _095744_);
  xor g_105775_(out[271], out[863], _095745_);
  xor g_105776_(out[266], out[858], _095746_);
  xor g_105777_(out[261], out[853], _095747_);
  xor g_105778_(out[256], out[848], _095748_);
  or g_105779_(_095735_, _095740_, _095749_);
  or g_105780_(_095736_, _095738_, _095750_);
  or g_105781_(_095741_, _095746_, _095751_);
  or g_105782_(_095750_, _095751_, _095752_);
  or g_105783_(_095739_, _095743_, _095753_);
  or g_105784_(_095747_, _095748_, _095754_);
  or g_105785_(_095753_, _095754_, _095755_);
  or g_105786_(_095752_, _095755_, _095756_);
  xor g_105787_(out[268], out[860], _095757_);
  or g_105788_(_095734_, _095757_, _095758_);
  or g_105789_(_095733_, _095744_, _095759_);
  or g_105790_(_095758_, _095759_, _095760_);
  or g_105791_(_095737_, _095742_, _095761_);
  or g_105792_(_095745_, _095761_, _095762_);
  or g_105793_(_095760_, _095762_, _095763_);
  or g_105794_(_095756_, _095763_, _095764_);
  or g_105795_(_095749_, _095764_, _095765_);
  xor g_105796_(out[252], out[860], _095766_);
  and g_105797_(_098239_, out[859], _095767_);
  xor g_105798_(out[253], out[861], _095768_);
  xor g_105799_(out[246], out[854], _095769_);
  xor g_105800_(out[248], out[856], _095770_);
  xor g_105801_(out[249], out[857], _095771_);
  xor g_105802_(out[254], out[862], _095772_);
  xor g_105803_(out[244], out[852], _095773_);
  or g_105804_(_095772_, _095773_, _095774_);
  xor g_105805_(out[245], out[853], _095775_);
  xor g_105806_(out[241], out[849], _095776_);
  and g_105807_(out[251], _049752_, _095777_);
  xor g_105808_(out[255], out[863], _095778_);
  xor g_105809_(out[250], out[858], _095779_);
  xor g_105810_(out[240], out[848], _095780_);
  xor g_105811_(out[242], out[850], _095781_);
  xor g_105812_(out[243], out[851], _095782_);
  or g_105813_(_095768_, _095770_, _095783_);
  or g_105814_(_095779_, _095781_, _095784_);
  or g_105815_(_095783_, _095784_, _095785_);
  or g_105816_(_095771_, _095782_, _095786_);
  or g_105817_(_095775_, _095780_, _095787_);
  or g_105818_(_095786_, _095787_, _095788_);
  or g_105819_(_095785_, _095788_, _095789_);
  or g_105820_(_095766_, _095767_, _095790_);
  xor g_105821_(out[247], out[855], _095791_);
  or g_105822_(_095769_, _095791_, _095792_);
  or g_105823_(_095790_, _095792_, _095793_);
  or g_105824_(_095776_, _095777_, _095794_);
  or g_105825_(_095778_, _095794_, _095795_);
  or g_105826_(_095793_, _095795_, _095796_);
  or g_105827_(_095789_, _095796_, _095797_);
  or g_105828_(_095774_, _095797_, _095798_);
  xor g_105829_(out[231], out[855], _095799_);
  and g_105830_(_098228_, out[859], _095800_);
  xor g_105831_(out[238], out[862], _095801_);
  xor g_105832_(out[232], out[856], _095802_);
  xor g_105833_(out[225], out[849], _095803_);
  xor g_105834_(out[237], out[861], _095804_);
  xor g_105835_(out[233], out[857], _095805_);
  xor g_105836_(out[228], out[852], _095806_);
  xor g_105837_(out[226], out[850], _095807_);
  and g_105838_(out[235], _049752_, _095808_);
  xor g_105839_(out[227], out[851], _095809_);
  xor g_105840_(out[230], out[854], _095810_);
  xor g_105841_(out[239], out[863], _095811_);
  xor g_105842_(out[234], out[858], _095812_);
  xor g_105843_(out[229], out[853], _095813_);
  xor g_105844_(out[224], out[848], _095814_);
  or g_105845_(_095801_, _095806_, _095815_);
  or g_105846_(_095802_, _095804_, _095816_);
  or g_105847_(_095807_, _095812_, _095817_);
  or g_105848_(_095816_, _095817_, _095818_);
  or g_105849_(_095805_, _095809_, _095819_);
  or g_105850_(_095813_, _095814_, _095820_);
  or g_105851_(_095819_, _095820_, _095821_);
  or g_105852_(_095818_, _095821_, _095822_);
  xor g_105853_(out[236], out[860], _095823_);
  or g_105854_(_095800_, _095823_, _095824_);
  or g_105855_(_095799_, _095810_, _095825_);
  or g_105856_(_095824_, _095825_, _095826_);
  or g_105857_(_095803_, _095808_, _095827_);
  or g_105858_(_095811_, _095827_, _095828_);
  or g_105859_(_095826_, _095828_, _095829_);
  or g_105860_(_095822_, _095829_, _095830_);
  or g_105861_(_095815_, _095830_, _095831_);
  not g_105862_(_095831_, _095832_);
  xor g_105863_(out[209], out[849], _095833_);
  and g_105864_(out[219], _049752_, _095834_);
  xor g_105865_(out[217], out[857], _095835_);
  xor g_105866_(out[208], out[848], _095836_);
  xor g_105867_(out[222], out[862], _095837_);
  xor g_105868_(out[212], out[852], _095838_);
  or g_105869_(_095837_, _095838_, _095839_);
  xor g_105870_(out[221], out[861], _095840_);
  xor g_105871_(out[211], out[851], _095841_);
  and g_105872_(_098217_, out[859], _095842_);
  xor g_105873_(out[214], out[854], _095843_);
  xor g_105874_(out[218], out[858], _095844_);
  xor g_105875_(out[213], out[853], _095845_);
  xor g_105876_(out[223], out[863], _095846_);
  xor g_105877_(out[216], out[856], _095847_);
  or g_105878_(_095840_, _095847_, _095848_);
  xor g_105879_(out[210], out[850], _095849_);
  or g_105880_(_095844_, _095849_, _095850_);
  or g_105881_(_095848_, _095850_, _095851_);
  or g_105882_(_095835_, _095841_, _095852_);
  or g_105883_(_095845_, _095852_, _095853_);
  or g_105884_(_095851_, _095853_, _095854_);
  or g_105885_(_095839_, _095854_, _095855_);
  xor g_105886_(out[220], out[860], _095856_);
  or g_105887_(_095842_, _095856_, _095857_);
  xor g_105888_(out[215], out[855], _095858_);
  or g_105889_(_095843_, _095858_, _095859_);
  or g_105890_(_095857_, _095859_, _095860_);
  or g_105891_(_095833_, _095834_, _095861_);
  or g_105892_(_095846_, _095861_, _095862_);
  or g_105893_(_095860_, _095862_, _095863_);
  or g_105894_(_095836_, _095863_, _095864_);
  or g_105895_(_095855_, _095864_, _095865_);
  xor g_105896_(out[199], out[855], _095866_);
  and g_105897_(_098206_, out[859], _095867_);
  xor g_105898_(out[206], out[862], _095868_);
  xor g_105899_(out[200], out[856], _095869_);
  xor g_105900_(out[193], out[849], _095870_);
  xor g_105901_(out[205], out[861], _095871_);
  xor g_105902_(out[201], out[857], _095872_);
  xor g_105903_(out[196], out[852], _095873_);
  xor g_105904_(out[194], out[850], _095874_);
  and g_105905_(out[203], _049752_, _095875_);
  xor g_105906_(out[195], out[851], _095876_);
  xor g_105907_(out[198], out[854], _095877_);
  xor g_105908_(out[207], out[863], _095878_);
  xor g_105909_(out[202], out[858], _095879_);
  xor g_105910_(out[197], out[853], _095880_);
  xor g_105911_(out[192], out[848], _095881_);
  or g_105912_(_095868_, _095873_, _095882_);
  or g_105913_(_095869_, _095871_, _095883_);
  or g_105914_(_095874_, _095879_, _095884_);
  or g_105915_(_095883_, _095884_, _095885_);
  or g_105916_(_095872_, _095876_, _095886_);
  or g_105917_(_095880_, _095881_, _095887_);
  or g_105918_(_095886_, _095887_, _095888_);
  or g_105919_(_095885_, _095888_, _095889_);
  xor g_105920_(out[204], out[860], _095890_);
  or g_105921_(_095867_, _095890_, _095891_);
  or g_105922_(_095866_, _095877_, _095892_);
  or g_105923_(_095891_, _095892_, _095893_);
  or g_105924_(_095870_, _095875_, _095894_);
  or g_105925_(_095878_, _095894_, _095895_);
  or g_105926_(_095893_, _095895_, _095896_);
  or g_105927_(_095889_, _095896_, _095897_);
  or g_105928_(_095882_, _095897_, _095898_);
  xor g_105929_(out[177], out[849], _095899_);
  and g_105930_(out[187], _049752_, _095900_);
  xor g_105931_(out[185], out[857], _095901_);
  xor g_105932_(out[176], out[848], _095902_);
  xor g_105933_(out[190], out[862], _095903_);
  xor g_105934_(out[180], out[852], _095904_);
  or g_105935_(_095903_, _095904_, _095905_);
  xor g_105936_(out[189], out[861], _095906_);
  xor g_105937_(out[179], out[851], _095907_);
  and g_105938_(_098195_, out[859], _095908_);
  xor g_105939_(out[182], out[854], _095909_);
  xor g_105940_(out[186], out[858], _095910_);
  xor g_105941_(out[181], out[853], _095911_);
  xor g_105942_(out[191], out[863], _095912_);
  xor g_105943_(out[184], out[856], _095913_);
  or g_105944_(_095906_, _095913_, _095914_);
  xor g_105945_(out[178], out[850], _095915_);
  or g_105946_(_095910_, _095915_, _095916_);
  or g_105947_(_095914_, _095916_, _095917_);
  or g_105948_(_095901_, _095907_, _095918_);
  or g_105949_(_095911_, _095918_, _095919_);
  or g_105950_(_095917_, _095919_, _095920_);
  or g_105951_(_095905_, _095920_, _095921_);
  xor g_105952_(out[188], out[860], _095922_);
  or g_105953_(_095908_, _095922_, _095923_);
  xor g_105954_(out[183], out[855], _095924_);
  or g_105955_(_095909_, _095924_, _095925_);
  or g_105956_(_095923_, _095925_, _095926_);
  or g_105957_(_095899_, _095900_, _095927_);
  or g_105958_(_095912_, _095927_, _095928_);
  or g_105959_(_095926_, _095928_, _095929_);
  or g_105960_(_095902_, _095929_, _095930_);
  or g_105961_(_095921_, _095930_, _095931_);
  xor g_105962_(out[167], out[855], _095932_);
  and g_105963_(_098184_, out[859], _095933_);
  xor g_105964_(out[174], out[862], _095934_);
  xor g_105965_(out[168], out[856], _095935_);
  xor g_105966_(out[161], out[849], _095936_);
  xor g_105967_(out[173], out[861], _095937_);
  xor g_105968_(out[169], out[857], _095938_);
  xor g_105969_(out[164], out[852], _095939_);
  xor g_105970_(out[162], out[850], _095940_);
  and g_105971_(out[171], _049752_, _095941_);
  xor g_105972_(out[163], out[851], _095942_);
  xor g_105973_(out[166], out[854], _095943_);
  xor g_105974_(out[175], out[863], _095944_);
  xor g_105975_(out[170], out[858], _095945_);
  xor g_105976_(out[165], out[853], _095946_);
  xor g_105977_(out[160], out[848], _095947_);
  or g_105978_(_095934_, _095939_, _095948_);
  or g_105979_(_095935_, _095937_, _095949_);
  or g_105980_(_095940_, _095945_, _095950_);
  or g_105981_(_095949_, _095950_, _095951_);
  or g_105982_(_095938_, _095942_, _095952_);
  or g_105983_(_095946_, _095947_, _095953_);
  or g_105984_(_095952_, _095953_, _095954_);
  or g_105985_(_095951_, _095954_, _095955_);
  xor g_105986_(out[172], out[860], _095956_);
  or g_105987_(_095933_, _095956_, _095957_);
  or g_105988_(_095932_, _095943_, _095958_);
  or g_105989_(_095957_, _095958_, _095959_);
  or g_105990_(_095936_, _095941_, _095960_);
  or g_105991_(_095944_, _095960_, _095961_);
  or g_105992_(_095959_, _095961_, _095962_);
  or g_105993_(_095955_, _095962_, _095963_);
  or g_105994_(_095948_, _095963_, _095964_);
  xor g_105995_(out[145], out[849], _095965_);
  and g_105996_(out[155], _049752_, _095966_);
  xor g_105997_(out[153], out[857], _095967_);
  xor g_105998_(out[144], out[848], _095968_);
  xor g_105999_(out[158], out[862], _095969_);
  xor g_106000_(out[148], out[852], _095970_);
  or g_106001_(_095969_, _095970_, _095971_);
  xor g_106002_(out[157], out[861], _095972_);
  xor g_106003_(out[147], out[851], _095973_);
  and g_106004_(_098173_, out[859], _095974_);
  xor g_106005_(out[150], out[854], _095975_);
  xor g_106006_(out[154], out[858], _095976_);
  xor g_106007_(out[149], out[853], _095977_);
  xor g_106008_(out[159], out[863], _095978_);
  xor g_106009_(out[152], out[856], _095979_);
  or g_106010_(_095972_, _095979_, _095980_);
  xor g_106011_(out[146], out[850], _095981_);
  or g_106012_(_095976_, _095981_, _095982_);
  or g_106013_(_095980_, _095982_, _095983_);
  or g_106014_(_095967_, _095973_, _095984_);
  or g_106015_(_095977_, _095984_, _095985_);
  or g_106016_(_095983_, _095985_, _095986_);
  or g_106017_(_095971_, _095986_, _095987_);
  xor g_106018_(out[156], out[860], _095988_);
  or g_106019_(_095974_, _095988_, _095989_);
  xor g_106020_(out[151], out[855], _095990_);
  or g_106021_(_095975_, _095990_, _095991_);
  or g_106022_(_095989_, _095991_, _095992_);
  or g_106023_(_095965_, _095966_, _095993_);
  or g_106024_(_095978_, _095993_, _095994_);
  or g_106025_(_095992_, _095994_, _095995_);
  or g_106026_(_095968_, _095995_, _095996_);
  or g_106027_(_095987_, _095996_, _095997_);
  xor g_106028_(out[135], out[855], _095998_);
  and g_106029_(_098162_, out[859], _095999_);
  xor g_106030_(out[142], out[862], _096000_);
  xor g_106031_(out[136], out[856], _096001_);
  xor g_106032_(out[129], out[849], _096002_);
  xor g_106033_(out[141], out[861], _096003_);
  xor g_106034_(out[137], out[857], _096004_);
  xor g_106035_(out[132], out[852], _096005_);
  xor g_106036_(out[130], out[850], _096006_);
  and g_106037_(out[139], _049752_, _096007_);
  xor g_106038_(out[131], out[851], _096008_);
  xor g_106039_(out[134], out[854], _096009_);
  xor g_106040_(out[143], out[863], _096010_);
  xor g_106041_(out[138], out[858], _096011_);
  xor g_106042_(out[133], out[853], _096012_);
  xor g_106043_(out[128], out[848], _096013_);
  or g_106044_(_096000_, _096005_, _096014_);
  or g_106045_(_096001_, _096003_, _096015_);
  or g_106046_(_096006_, _096011_, _096016_);
  or g_106047_(_096015_, _096016_, _096017_);
  or g_106048_(_096004_, _096008_, _096018_);
  or g_106049_(_096012_, _096013_, _096019_);
  or g_106050_(_096018_, _096019_, _096020_);
  or g_106051_(_096017_, _096020_, _096021_);
  xor g_106052_(out[140], out[860], _096022_);
  or g_106053_(_095999_, _096022_, _096023_);
  or g_106054_(_095998_, _096009_, _096024_);
  or g_106055_(_096023_, _096024_, _096025_);
  or g_106056_(_096002_, _096007_, _096026_);
  or g_106057_(_096010_, _096026_, _096027_);
  or g_106058_(_096025_, _096027_, _096028_);
  or g_106059_(_096021_, _096028_, _096029_);
  or g_106060_(_096014_, _096029_, _096030_);
  xor g_106061_(out[124], out[860], _096031_);
  and g_106062_(_098151_, out[859], _096032_);
  xor g_106063_(out[120], out[856], _096033_);
  xor g_106064_(out[118], out[854], _096034_);
  xor g_106065_(out[125], out[861], _096035_);
  xor g_106066_(out[126], out[862], _096036_);
  xor g_106067_(out[114], out[850], _096037_);
  xor g_106068_(out[121], out[857], _096038_);
  xor g_106069_(out[117], out[853], _096039_);
  xor g_106070_(out[113], out[849], _096040_);
  and g_106071_(out[123], _049752_, _096041_);
  or g_106072_(_096033_, _096035_, _096042_);
  xor g_106073_(out[127], out[863], _096043_);
  xor g_106074_(out[122], out[858], _096044_);
  xor g_106075_(out[116], out[852], _096045_);
  xor g_106076_(out[115], out[851], _096046_);
  xor g_106077_(out[112], out[848], _096047_);
  or g_106078_(_096037_, _096044_, _096048_);
  or g_106079_(_096042_, _096048_, _096049_);
  or g_106080_(_096038_, _096046_, _096050_);
  or g_106081_(_096039_, _096050_, _096051_);
  or g_106082_(_096049_, _096051_, _096052_);
  or g_106083_(_096036_, _096045_, _096053_);
  or g_106084_(_096052_, _096053_, _096054_);
  or g_106085_(_096031_, _096032_, _096055_);
  xor g_106086_(out[119], out[855], _096056_);
  or g_106087_(_096034_, _096056_, _096057_);
  or g_106088_(_096055_, _096057_, _096058_);
  or g_106089_(_096040_, _096041_, _096059_);
  or g_106090_(_096043_, _096059_, _096060_);
  or g_106091_(_096058_, _096060_, _096061_);
  or g_106092_(_096047_, _096061_, _096062_);
  or g_106093_(_096054_, _096062_, _096063_);
  xor g_106094_(out[103], out[855], _096064_);
  and g_106095_(_098140_, out[859], _096065_);
  xor g_106096_(out[110], out[862], _096066_);
  xor g_106097_(out[104], out[856], _096067_);
  xor g_106098_(out[97], out[849], _096068_);
  xor g_106099_(out[109], out[861], _096069_);
  xor g_106100_(out[105], out[857], _096070_);
  xor g_106101_(out[100], out[852], _096071_);
  xor g_106102_(out[98], out[850], _096072_);
  and g_106103_(out[107], _049752_, _096073_);
  xor g_106104_(out[99], out[851], _096074_);
  xor g_106105_(out[102], out[854], _096075_);
  xor g_106106_(out[111], out[863], _096076_);
  xor g_106107_(out[106], out[858], _096077_);
  xor g_106108_(out[101], out[853], _096078_);
  xor g_106109_(out[96], out[848], _096079_);
  or g_106110_(_096066_, _096071_, _096080_);
  or g_106111_(_096067_, _096069_, _096081_);
  or g_106112_(_096072_, _096077_, _096082_);
  or g_106113_(_096081_, _096082_, _096083_);
  or g_106114_(_096070_, _096074_, _096084_);
  or g_106115_(_096078_, _096079_, _096085_);
  or g_106116_(_096084_, _096085_, _096086_);
  or g_106117_(_096083_, _096086_, _096087_);
  xor g_106118_(out[108], out[860], _096088_);
  or g_106119_(_096065_, _096088_, _096089_);
  or g_106120_(_096064_, _096075_, _096090_);
  or g_106121_(_096089_, _096090_, _096091_);
  or g_106122_(_096068_, _096073_, _096092_);
  or g_106123_(_096076_, _096092_, _096093_);
  or g_106124_(_096091_, _096093_, _096094_);
  or g_106125_(_096087_, _096094_, _096095_);
  or g_106126_(_096080_, _096095_, _096096_);
  not g_106127_(_096096_, _096097_);
  and g_106128_(_098129_, out[859], _096098_);
  and g_106129_(out[91], _049752_, _096099_);
  xor g_106130_(out[84], out[852], _096100_);
  xor g_106131_(out[82], out[850], _096101_);
  xor g_106132_(out[89], out[857], _096102_);
  xor g_106133_(out[80], out[848], _096103_);
  xor g_106134_(out[83], out[851], _096104_);
  xor g_106135_(out[90], out[858], _096105_);
  xor g_106136_(out[95], out[863], _096106_);
  xor g_106137_(out[86], out[854], _096107_);
  xor g_106138_(out[85], out[853], _096108_);
  xor g_106139_(out[93], out[861], _096109_);
  xor g_106140_(out[94], out[862], _096110_);
  xor g_106141_(out[88], out[856], _096111_);
  xor g_106142_(out[81], out[849], _096112_);
  or g_106143_(_096100_, _096110_, _096113_);
  or g_106144_(_096109_, _096111_, _096114_);
  or g_106145_(_096101_, _096105_, _096115_);
  or g_106146_(_096114_, _096115_, _096116_);
  or g_106147_(_096102_, _096104_, _096117_);
  or g_106148_(_096103_, _096108_, _096118_);
  or g_106149_(_096117_, _096118_, _096119_);
  or g_106150_(_096116_, _096119_, _096120_);
  xor g_106151_(out[92], out[860], _096121_);
  or g_106152_(_096098_, _096121_, _096122_);
  xor g_106153_(out[87], out[855], _096123_);
  or g_106154_(_096107_, _096123_, _096124_);
  or g_106155_(_096122_, _096124_, _096125_);
  or g_106156_(_096099_, _096112_, _096126_);
  or g_106157_(_096106_, _096126_, _096127_);
  or g_106158_(_096125_, _096127_, _096128_);
  or g_106159_(_096120_, _096128_, _096129_);
  or g_106160_(_096113_, _096129_, _096130_);
  xor g_106161_(out[71], out[855], _096131_);
  and g_106162_(_098118_, out[859], _096132_);
  xor g_106163_(out[78], out[862], _096133_);
  xor g_106164_(out[72], out[856], _096134_);
  xor g_106165_(out[65], out[849], _096135_);
  xor g_106166_(out[77], out[861], _096136_);
  xor g_106167_(out[73], out[857], _096137_);
  xor g_106168_(out[68], out[852], _096138_);
  xor g_106169_(out[66], out[850], _096139_);
  and g_106170_(out[75], _049752_, _096140_);
  xor g_106171_(out[67], out[851], _096141_);
  xor g_106172_(out[70], out[854], _096142_);
  xor g_106173_(out[79], out[863], _096143_);
  xor g_106174_(out[74], out[858], _096144_);
  xor g_106175_(out[69], out[853], _096145_);
  xor g_106176_(out[64], out[848], _096146_);
  or g_106177_(_096133_, _096138_, _096147_);
  or g_106178_(_096134_, _096136_, _096148_);
  or g_106179_(_096139_, _096144_, _096149_);
  or g_106180_(_096148_, _096149_, _096150_);
  or g_106181_(_096137_, _096141_, _096151_);
  or g_106182_(_096145_, _096146_, _096152_);
  or g_106183_(_096151_, _096152_, _096153_);
  or g_106184_(_096150_, _096153_, _096154_);
  xor g_106185_(out[76], out[860], _096155_);
  or g_106186_(_096132_, _096155_, _096156_);
  or g_106187_(_096131_, _096142_, _096157_);
  or g_106188_(_096156_, _096157_, _096158_);
  or g_106189_(_096135_, _096140_, _096159_);
  or g_106190_(_096143_, _096159_, _096160_);
  or g_106191_(_096158_, _096160_, _096161_);
  or g_106192_(_096154_, _096161_, _096162_);
  or g_106193_(_096147_, _096162_, _096163_);
  xor g_106194_(out[56], out[856], _096164_);
  xor g_106195_(out[53], out[853], _096165_);
  xor g_106196_(out[51], out[851], _096166_);
  xor g_106197_(out[62], out[862], _096167_);
  xor g_106198_(out[61], out[861], _096168_);
  xor g_106199_(out[50], out[850], _096169_);
  xor g_106200_(out[57], out[857], _096170_);
  xor g_106201_(out[54], out[854], _096171_);
  xor g_106202_(out[63], out[863], _096172_);
  xor g_106203_(out[58], out[858], _096173_);
  xor g_106204_(out[52], out[852], _096174_);
  xor g_106205_(out[48], out[848], _096175_);
  and g_106206_(_098107_, out[859], _096176_);
  and g_106207_(out[59], _049752_, _096177_);
  or g_106208_(_096164_, _096168_, _096178_);
  xor g_106209_(out[49], out[849], _096179_);
  or g_106210_(_096169_, _096173_, _096180_);
  or g_106211_(_096178_, _096180_, _096181_);
  or g_106212_(_096166_, _096170_, _096182_);
  or g_106213_(_096165_, _096182_, _096183_);
  or g_106214_(_096181_, _096183_, _096184_);
  or g_106215_(_096167_, _096174_, _096185_);
  or g_106216_(_096184_, _096185_, _096186_);
  xor g_106217_(out[60], out[860], _096187_);
  or g_106218_(_096176_, _096187_, _096188_);
  xor g_106219_(out[55], out[855], _096189_);
  or g_106220_(_096171_, _096189_, _096190_);
  or g_106221_(_096188_, _096190_, _096191_);
  or g_106222_(_096177_, _096179_, _096192_);
  or g_106223_(_096172_, _096192_, _096193_);
  or g_106224_(_096191_, _096193_, _096194_);
  or g_106225_(_096175_, _096194_, _096195_);
  or g_106226_(_096186_, _096195_, _096196_);
  not g_106227_(_096196_, _096197_);
  xor g_106228_(out[39], out[855], _096198_);
  and g_106229_(_098096_, out[859], _096199_);
  xor g_106230_(out[46], out[862], _096200_);
  xor g_106231_(out[40], out[856], _096201_);
  xor g_106232_(out[33], out[849], _096202_);
  xor g_106233_(out[45], out[861], _096203_);
  xor g_106234_(out[41], out[857], _096204_);
  xor g_106235_(out[36], out[852], _096205_);
  xor g_106236_(out[34], out[850], _096206_);
  and g_106237_(out[43], _049752_, _096207_);
  xor g_106238_(out[35], out[851], _096208_);
  xor g_106239_(out[38], out[854], _096209_);
  xor g_106240_(out[47], out[863], _096210_);
  xor g_106241_(out[42], out[858], _096211_);
  xor g_106242_(out[37], out[853], _096212_);
  xor g_106243_(out[32], out[848], _096213_);
  or g_106244_(_096200_, _096205_, _096214_);
  or g_106245_(_096201_, _096203_, _096215_);
  or g_106246_(_096206_, _096211_, _096216_);
  or g_106247_(_096215_, _096216_, _096217_);
  or g_106248_(_096204_, _096208_, _096218_);
  or g_106249_(_096212_, _096213_, _096219_);
  or g_106250_(_096218_, _096219_, _096220_);
  or g_106251_(_096217_, _096220_, _096221_);
  xor g_106252_(out[44], out[860], _096222_);
  or g_106253_(_096199_, _096222_, _096223_);
  or g_106254_(_096198_, _096209_, _096224_);
  or g_106255_(_096223_, _096224_, _096225_);
  or g_106256_(_096202_, _096207_, _096226_);
  or g_106257_(_096210_, _096226_, _096227_);
  or g_106258_(_096225_, _096227_, _096228_);
  or g_106259_(_096221_, _096228_, _096229_);
  or g_106260_(_096214_, _096229_, _096230_);
  xor g_106261_(out[17], out[849], _096231_);
  and g_106262_(out[27], _049752_, _096232_);
  xor g_106263_(out[25], out[857], _096233_);
  xor g_106264_(out[16], out[848], _096234_);
  xor g_106265_(out[30], out[862], _096235_);
  xor g_106266_(out[20], out[852], _096236_);
  or g_106267_(_096235_, _096236_, _096237_);
  xor g_106268_(out[29], out[861], _096238_);
  xor g_106269_(out[19], out[851], _096239_);
  and g_106270_(_098063_, out[859], _096240_);
  xor g_106271_(out[22], out[854], _096241_);
  xor g_106272_(out[26], out[858], _096242_);
  xor g_106273_(out[21], out[853], _096243_);
  xor g_106274_(out[31], out[863], _096244_);
  xor g_106275_(out[24], out[856], _096245_);
  or g_106276_(_096238_, _096245_, _096246_);
  xor g_106277_(out[18], out[850], _096247_);
  or g_106278_(_096242_, _096247_, _096248_);
  or g_106279_(_096246_, _096248_, _096249_);
  or g_106280_(_096233_, _096239_, _096250_);
  or g_106281_(_096243_, _096250_, _096251_);
  or g_106282_(_096249_, _096251_, _096252_);
  or g_106283_(_096237_, _096252_, _096253_);
  xor g_106284_(out[28], out[860], _096254_);
  or g_106285_(_096240_, _096254_, _096255_);
  xor g_106286_(out[23], out[855], _096256_);
  or g_106287_(_096241_, _096256_, _096257_);
  or g_106288_(_096255_, _096257_, _096258_);
  or g_106289_(_096231_, _096232_, _096259_);
  or g_106290_(_096244_, _096259_, _096260_);
  or g_106291_(_096258_, _096260_, _096261_);
  or g_106292_(_096234_, _096261_, _096262_);
  or g_106293_(_096253_, _096262_, _096263_);
  xor g_106294_(out[1], out[849], _096264_);
  and g_106295_(out[11], _049752_, _096265_);
  xor g_106296_(out[9], out[857], _096266_);
  xor g_106297_(out[0], out[848], _096267_);
  xor g_106298_(out[14], out[862], _096268_);
  xor g_106299_(out[4], out[852], _096269_);
  or g_106300_(_096268_, _096269_, _096270_);
  xor g_106301_(out[13], out[861], _096271_);
  xor g_106302_(out[3], out[851], _096272_);
  and g_106303_(_098041_, out[859], _096273_);
  xor g_106304_(out[6], out[854], _096274_);
  xor g_106305_(out[10], out[858], _096275_);
  xor g_106306_(out[5], out[853], _096276_);
  xor g_106307_(out[15], out[863], _096277_);
  xor g_106308_(out[8], out[856], _096278_);
  or g_106309_(_096271_, _096278_, _096279_);
  xor g_106310_(out[2], out[850], _096280_);
  or g_106311_(_096275_, _096280_, _096281_);
  or g_106312_(_096279_, _096281_, _096282_);
  or g_106313_(_096266_, _096272_, _096283_);
  or g_106314_(_096276_, _096283_, _096284_);
  or g_106315_(_096282_, _096284_, _096285_);
  or g_106316_(_096270_, _096285_, _096286_);
  xor g_106317_(out[12], out[860], _096287_);
  or g_106318_(_096273_, _096287_, _096288_);
  xor g_106319_(out[7], out[855], _096289_);
  or g_106320_(_096274_, _096289_, _096290_);
  or g_106321_(_096288_, _096290_, _096291_);
  or g_106322_(_096264_, _096265_, _096292_);
  or g_106323_(_096277_, _096292_, _096293_);
  or g_106324_(_096291_, _096293_, _096294_);
  or g_106325_(_096267_, _096294_, _096295_);
  or g_106326_(_096286_, _096295_, _096296_);
  not g_106327_(_096296_, _096297_);
  xor g_106328_(out[471], out[839], _096298_);
  and g_106329_(_049499_, out[843], _096299_);
  xor g_106330_(out[478], out[846], _096300_);
  xor g_106331_(out[472], out[840], _096301_);
  xor g_106332_(out[465], out[833], _096302_);
  xor g_106333_(out[477], out[845], _096303_);
  xor g_106334_(out[473], out[841], _096304_);
  xor g_106335_(out[468], out[836], _096305_);
  xor g_106336_(out[466], out[834], _096306_);
  and g_106337_(out[475], _049741_, _096307_);
  xor g_106338_(out[467], out[835], _096308_);
  xor g_106339_(out[470], out[838], _096309_);
  xor g_106340_(out[479], out[847], _096310_);
  xor g_106341_(out[474], out[842], _096311_);
  xor g_106342_(out[469], out[837], _096312_);
  xor g_106343_(out[464], out[832], _096313_);
  or g_106344_(_096300_, _096305_, _096314_);
  or g_106345_(_096301_, _096303_, _096315_);
  or g_106346_(_096306_, _096311_, _096316_);
  or g_106347_(_096315_, _096316_, _096317_);
  or g_106348_(_096304_, _096308_, _096318_);
  or g_106349_(_096312_, _096313_, _096319_);
  or g_106350_(_096318_, _096319_, _096320_);
  or g_106351_(_096317_, _096320_, _096321_);
  xor g_106352_(out[476], out[844], _096322_);
  or g_106353_(_096299_, _096322_, _096323_);
  or g_106354_(_096298_, _096309_, _096324_);
  or g_106355_(_096323_, _096324_, _096325_);
  or g_106356_(_096302_, _096307_, _096326_);
  or g_106357_(_096310_, _096326_, _096327_);
  or g_106358_(_096325_, _096327_, _096328_);
  or g_106359_(_096321_, _096328_, _096329_);
  or g_106360_(_096314_, _096329_, _096330_);
  not g_106361_(_096330_, _096331_);
  xor g_106362_(out[452], out[836], _096332_);
  xor g_106363_(out[460], out[844], _096333_);
  and g_106364_(_049477_, out[843], _096334_);
  xor g_106365_(out[458], out[842], _096335_);
  xor g_106366_(out[454], out[838], _096336_);
  xor g_106367_(out[453], out[837], _096337_);
  xor g_106368_(out[451], out[835], _096338_);
  xor g_106369_(out[461], out[845], _096339_);
  xor g_106370_(out[462], out[846], _096340_);
  xor g_106371_(out[449], out[833], _096341_);
  xor g_106372_(out[450], out[834], _096342_);
  and g_106373_(out[459], _049741_, _096343_);
  xor g_106374_(out[448], out[832], _096344_);
  xor g_106375_(out[463], out[847], _096345_);
  xor g_106376_(out[456], out[840], _096346_);
  or g_106377_(_096339_, _096346_, _096347_);
  xor g_106378_(out[457], out[841], _096348_);
  or g_106379_(_096335_, _096342_, _096349_);
  or g_106380_(_096347_, _096349_, _096350_);
  or g_106381_(_096338_, _096348_, _096351_);
  or g_106382_(_096337_, _096351_, _096352_);
  or g_106383_(_096350_, _096352_, _096353_);
  or g_106384_(_096332_, _096340_, _096354_);
  or g_106385_(_096353_, _096354_, _096355_);
  or g_106386_(_096333_, _096334_, _096356_);
  xor g_106387_(out[455], out[839], _096357_);
  or g_106388_(_096336_, _096357_, _096358_);
  or g_106389_(_096356_, _096358_, _096359_);
  or g_106390_(_096341_, _096343_, _096360_);
  or g_106391_(_096345_, _096360_, _096361_);
  or g_106392_(_096359_, _096361_, _096362_);
  or g_106393_(_096344_, _096362_, _096363_);
  or g_106394_(_096355_, _096363_, _096364_);
  not g_106395_(_096364_, _096365_);
  xor g_106396_(out[439], out[839], _096366_);
  and g_106397_(_049466_, out[843], _096367_);
  xor g_106398_(out[446], out[846], _096368_);
  xor g_106399_(out[440], out[840], _096369_);
  xor g_106400_(out[433], out[833], _096370_);
  xor g_106401_(out[445], out[845], _096371_);
  xor g_106402_(out[441], out[841], _096372_);
  xor g_106403_(out[436], out[836], _096373_);
  xor g_106404_(out[434], out[834], _096374_);
  and g_106405_(out[443], _049741_, _096375_);
  xor g_106406_(out[435], out[835], _096376_);
  xor g_106407_(out[438], out[838], _096377_);
  xor g_106408_(out[447], out[847], _096378_);
  xor g_106409_(out[442], out[842], _096379_);
  xor g_106410_(out[437], out[837], _096380_);
  xor g_106411_(out[432], out[832], _096381_);
  or g_106412_(_096368_, _096373_, _096382_);
  or g_106413_(_096369_, _096371_, _096383_);
  or g_106414_(_096374_, _096379_, _096384_);
  or g_106415_(_096383_, _096384_, _096385_);
  or g_106416_(_096372_, _096376_, _096386_);
  or g_106417_(_096380_, _096381_, _096387_);
  or g_106418_(_096386_, _096387_, _096388_);
  or g_106419_(_096385_, _096388_, _096389_);
  xor g_106420_(out[444], out[844], _096390_);
  or g_106421_(_096367_, _096390_, _096391_);
  or g_106422_(_096366_, _096377_, _096392_);
  or g_106423_(_096391_, _096392_, _096393_);
  or g_106424_(_096370_, _096375_, _096394_);
  or g_106425_(_096378_, _096394_, _096395_);
  or g_106426_(_096393_, _096395_, _096396_);
  or g_106427_(_096389_, _096396_, _096397_);
  or g_106428_(_096382_, _096397_, _096398_);
  not g_106429_(_096398_, _096399_);
  xor g_106430_(out[417], out[833], _096400_);
  and g_106431_(out[427], _049741_, _096401_);
  xor g_106432_(out[425], out[841], _096402_);
  xor g_106433_(out[416], out[832], _096403_);
  xor g_106434_(out[430], out[846], _096404_);
  xor g_106435_(out[420], out[836], _096405_);
  or g_106436_(_096404_, _096405_, _096406_);
  xor g_106437_(out[429], out[845], _096407_);
  xor g_106438_(out[419], out[835], _096408_);
  and g_106439_(_049455_, out[843], _096409_);
  xor g_106440_(out[422], out[838], _096410_);
  xor g_106441_(out[426], out[842], _096411_);
  xor g_106442_(out[421], out[837], _096412_);
  xor g_106443_(out[431], out[847], _096413_);
  xor g_106444_(out[424], out[840], _096414_);
  or g_106445_(_096407_, _096414_, _096415_);
  xor g_106446_(out[418], out[834], _096416_);
  or g_106447_(_096411_, _096416_, _096417_);
  or g_106448_(_096415_, _096417_, _096418_);
  or g_106449_(_096402_, _096408_, _096419_);
  or g_106450_(_096412_, _096419_, _096420_);
  or g_106451_(_096418_, _096420_, _096421_);
  or g_106452_(_096406_, _096421_, _096422_);
  xor g_106453_(out[428], out[844], _096423_);
  or g_106454_(_096409_, _096423_, _096424_);
  xor g_106455_(out[423], out[839], _096425_);
  or g_106456_(_096410_, _096425_, _096426_);
  or g_106457_(_096424_, _096426_, _096427_);
  or g_106458_(_096400_, _096401_, _096428_);
  or g_106459_(_096413_, _096428_, _096429_);
  or g_106460_(_096427_, _096429_, _096430_);
  or g_106461_(_096403_, _096430_, _096431_);
  or g_106462_(_096422_, _096431_, _096432_);
  xor g_106463_(out[407], out[839], _096433_);
  and g_106464_(_049444_, out[843], _096434_);
  xor g_106465_(out[414], out[846], _096435_);
  xor g_106466_(out[408], out[840], _096436_);
  xor g_106467_(out[401], out[833], _096437_);
  xor g_106468_(out[413], out[845], _096438_);
  xor g_106469_(out[409], out[841], _096439_);
  xor g_106470_(out[404], out[836], _096440_);
  xor g_106471_(out[402], out[834], _096441_);
  and g_106472_(out[411], _049741_, _096442_);
  xor g_106473_(out[403], out[835], _096443_);
  xor g_106474_(out[406], out[838], _096444_);
  xor g_106475_(out[415], out[847], _096445_);
  xor g_106476_(out[410], out[842], _096446_);
  xor g_106477_(out[405], out[837], _096447_);
  xor g_106478_(out[400], out[832], _096448_);
  or g_106479_(_096435_, _096440_, _096449_);
  or g_106480_(_096436_, _096438_, _096450_);
  or g_106481_(_096441_, _096446_, _096451_);
  or g_106482_(_096450_, _096451_, _096452_);
  or g_106483_(_096439_, _096443_, _096453_);
  or g_106484_(_096447_, _096448_, _096454_);
  or g_106485_(_096453_, _096454_, _096455_);
  or g_106486_(_096452_, _096455_, _096456_);
  xor g_106487_(out[412], out[844], _096457_);
  or g_106488_(_096434_, _096457_, _096458_);
  or g_106489_(_096433_, _096444_, _096459_);
  or g_106490_(_096458_, _096459_, _096460_);
  or g_106491_(_096437_, _096442_, _096461_);
  or g_106492_(_096445_, _096461_, _096462_);
  or g_106493_(_096460_, _096462_, _096463_);
  or g_106494_(_096456_, _096463_, _096464_);
  or g_106495_(_096449_, _096464_, _096465_);
  and g_106496_(out[395], _049741_, _096466_);
  and g_106497_(_049433_, out[843], _096467_);
  xor g_106498_(out[392], out[840], _096468_);
  xor g_106499_(out[399], out[847], _096469_);
  xor g_106500_(out[385], out[833], _096470_);
  xor g_106501_(out[386], out[834], _096471_);
  xor g_106502_(out[388], out[836], _096472_);
  xor g_106503_(out[389], out[837], _096473_);
  xor g_106504_(out[393], out[841], _096474_);
  xor g_106505_(out[387], out[835], _096475_);
  xor g_106506_(out[398], out[846], _096476_);
  xor g_106507_(out[384], out[832], _096477_);
  xor g_106508_(out[394], out[842], _096478_);
  xor g_106509_(out[397], out[845], _096479_);
  or g_106510_(_096468_, _096479_, _096480_);
  xor g_106511_(out[390], out[838], _096481_);
  or g_106512_(_096471_, _096478_, _096482_);
  or g_106513_(_096480_, _096482_, _096483_);
  or g_106514_(_096474_, _096475_, _096484_);
  or g_106515_(_096473_, _096484_, _096485_);
  or g_106516_(_096483_, _096485_, _096486_);
  or g_106517_(_096472_, _096476_, _096487_);
  or g_106518_(_096486_, _096487_, _096488_);
  xor g_106519_(out[396], out[844], _096489_);
  or g_106520_(_096467_, _096489_, _096490_);
  xor g_106521_(out[391], out[839], _096491_);
  or g_106522_(_096481_, _096491_, _096492_);
  or g_106523_(_096490_, _096492_, _096493_);
  or g_106524_(_096466_, _096470_, _096494_);
  or g_106525_(_096469_, _096494_, _096495_);
  or g_106526_(_096493_, _096495_, _096496_);
  or g_106527_(_096477_, _096496_, _096497_);
  or g_106528_(_096488_, _096497_, _096498_);
  xor g_106529_(out[375], out[839], _096499_);
  and g_106530_(_049422_, out[843], _096500_);
  xor g_106531_(out[382], out[846], _096501_);
  xor g_106532_(out[376], out[840], _096502_);
  xor g_106533_(out[369], out[833], _096503_);
  xor g_106534_(out[381], out[845], _096504_);
  xor g_106535_(out[377], out[841], _096505_);
  xor g_106536_(out[372], out[836], _096506_);
  xor g_106537_(out[370], out[834], _096507_);
  and g_106538_(out[379], _049741_, _096508_);
  xor g_106539_(out[371], out[835], _096509_);
  xor g_106540_(out[374], out[838], _096510_);
  xor g_106541_(out[383], out[847], _096511_);
  xor g_106542_(out[378], out[842], _096512_);
  xor g_106543_(out[373], out[837], _096513_);
  xor g_106544_(out[368], out[832], _096514_);
  or g_106545_(_096501_, _096506_, _096515_);
  or g_106546_(_096502_, _096504_, _096516_);
  or g_106547_(_096507_, _096512_, _096517_);
  or g_106548_(_096516_, _096517_, _096518_);
  or g_106549_(_096505_, _096509_, _096519_);
  or g_106550_(_096513_, _096514_, _096520_);
  or g_106551_(_096519_, _096520_, _096521_);
  or g_106552_(_096518_, _096521_, _096522_);
  xor g_106553_(out[380], out[844], _096523_);
  or g_106554_(_096500_, _096523_, _096524_);
  or g_106555_(_096499_, _096510_, _096525_);
  or g_106556_(_096524_, _096525_, _096526_);
  or g_106557_(_096503_, _096508_, _096527_);
  or g_106558_(_096511_, _096527_, _096528_);
  or g_106559_(_096526_, _096528_, _096529_);
  or g_106560_(_096522_, _096529_, _096530_);
  or g_106561_(_096515_, _096530_, _096531_);
  xor g_106562_(out[362], out[842], _096532_);
  xor g_106563_(out[354], out[834], _096533_);
  xor g_106564_(out[353], out[833], _096534_);
  and g_106565_(_049411_, out[843], _096535_);
  and g_106566_(out[363], _049741_, _096536_);
  xor g_106567_(out[365], out[845], _096537_);
  xor g_106568_(out[355], out[835], _096538_);
  xor g_106569_(out[366], out[846], _096539_);
  xor g_106570_(out[364], out[844], _096540_);
  xor g_106571_(out[360], out[840], _096541_);
  xor g_106572_(out[367], out[847], _096542_);
  xor g_106573_(out[357], out[837], _096543_);
  xor g_106574_(out[358], out[838], _096544_);
  xor g_106575_(out[352], out[832], _096545_);
  xor g_106576_(out[356], out[836], _096546_);
  or g_106577_(_096537_, _096541_, _096547_);
  xor g_106578_(out[361], out[841], _096548_);
  or g_106579_(_096532_, _096533_, _096549_);
  or g_106580_(_096547_, _096549_, _096550_);
  or g_106581_(_096538_, _096548_, _096551_);
  or g_106582_(_096543_, _096551_, _096552_);
  or g_106583_(_096550_, _096552_, _096553_);
  or g_106584_(_096539_, _096546_, _096554_);
  or g_106585_(_096553_, _096554_, _096555_);
  or g_106586_(_096535_, _096540_, _096556_);
  xor g_106587_(out[359], out[839], _096557_);
  or g_106588_(_096544_, _096557_, _096558_);
  or g_106589_(_096556_, _096558_, _096559_);
  or g_106590_(_096534_, _096536_, _096560_);
  or g_106591_(_096542_, _096560_, _096561_);
  or g_106592_(_096559_, _096561_, _096562_);
  or g_106593_(_096545_, _096562_, _096563_);
  or g_106594_(_096555_, _096563_, _096564_);
  not g_106595_(_096564_, _096565_);
  xor g_106596_(out[343], out[839], _096566_);
  and g_106597_(_049400_, out[843], _096567_);
  xor g_106598_(out[350], out[846], _096568_);
  xor g_106599_(out[344], out[840], _096569_);
  xor g_106600_(out[337], out[833], _096570_);
  xor g_106601_(out[349], out[845], _096571_);
  xor g_106602_(out[345], out[841], _096572_);
  xor g_106603_(out[340], out[836], _096573_);
  xor g_106604_(out[338], out[834], _096574_);
  and g_106605_(out[347], _049741_, _096575_);
  xor g_106606_(out[339], out[835], _096576_);
  xor g_106607_(out[342], out[838], _096577_);
  xor g_106608_(out[351], out[847], _096578_);
  xor g_106609_(out[346], out[842], _096579_);
  xor g_106610_(out[341], out[837], _096580_);
  xor g_106611_(out[336], out[832], _096581_);
  or g_106612_(_096568_, _096573_, _096582_);
  or g_106613_(_096569_, _096571_, _096583_);
  or g_106614_(_096574_, _096579_, _096584_);
  or g_106615_(_096583_, _096584_, _096585_);
  or g_106616_(_096572_, _096576_, _096586_);
  or g_106617_(_096580_, _096581_, _096587_);
  or g_106618_(_096586_, _096587_, _096588_);
  or g_106619_(_096585_, _096588_, _096589_);
  xor g_106620_(out[348], out[844], _096590_);
  or g_106621_(_096567_, _096590_, _096591_);
  or g_106622_(_096566_, _096577_, _096592_);
  or g_106623_(_096591_, _096592_, _096593_);
  or g_106624_(_096570_, _096575_, _096594_);
  or g_106625_(_096578_, _096594_, _096595_);
  or g_106626_(_096593_, _096595_, _096596_);
  or g_106627_(_096589_, _096596_, _096597_);
  or g_106628_(_096582_, _096597_, _096598_);
  xor g_106629_(out[328], out[840], _096599_);
  xor g_106630_(out[325], out[837], _096600_);
  xor g_106631_(out[323], out[835], _096601_);
  xor g_106632_(out[334], out[846], _096602_);
  xor g_106633_(out[333], out[845], _096603_);
  xor g_106634_(out[322], out[834], _096604_);
  xor g_106635_(out[329], out[841], _096605_);
  xor g_106636_(out[326], out[838], _096606_);
  xor g_106637_(out[335], out[847], _096607_);
  xor g_106638_(out[330], out[842], _096608_);
  xor g_106639_(out[324], out[836], _096609_);
  xor g_106640_(out[320], out[832], _096610_);
  and g_106641_(_098294_, out[843], _096611_);
  and g_106642_(out[331], _049741_, _096612_);
  or g_106643_(_096599_, _096603_, _096613_);
  xor g_106644_(out[321], out[833], _096614_);
  or g_106645_(_096604_, _096608_, _096615_);
  or g_106646_(_096613_, _096615_, _096616_);
  or g_106647_(_096601_, _096605_, _096617_);
  or g_106648_(_096600_, _096617_, _096618_);
  or g_106649_(_096616_, _096618_, _096619_);
  or g_106650_(_096602_, _096609_, _096620_);
  or g_106651_(_096619_, _096620_, _096621_);
  xor g_106652_(out[332], out[844], _096622_);
  or g_106653_(_096611_, _096622_, _096623_);
  xor g_106654_(out[327], out[839], _096624_);
  or g_106655_(_096606_, _096624_, _096625_);
  or g_106656_(_096623_, _096625_, _096626_);
  or g_106657_(_096612_, _096614_, _096627_);
  or g_106658_(_096607_, _096627_, _096628_);
  or g_106659_(_096626_, _096628_, _096629_);
  or g_106660_(_096610_, _096629_, _096630_);
  or g_106661_(_096621_, _096630_, _096631_);
  xor g_106662_(out[311], out[839], _096632_);
  and g_106663_(_098283_, out[843], _096633_);
  xor g_106664_(out[318], out[846], _096634_);
  xor g_106665_(out[312], out[840], _096635_);
  xor g_106666_(out[305], out[833], _096636_);
  xor g_106667_(out[317], out[845], _096637_);
  xor g_106668_(out[313], out[841], _096638_);
  xor g_106669_(out[308], out[836], _096639_);
  xor g_106670_(out[306], out[834], _096640_);
  and g_106671_(out[315], _049741_, _096641_);
  xor g_106672_(out[307], out[835], _096642_);
  xor g_106673_(out[310], out[838], _096643_);
  xor g_106674_(out[319], out[847], _096644_);
  xor g_106675_(out[314], out[842], _096645_);
  xor g_106676_(out[309], out[837], _096646_);
  xor g_106677_(out[304], out[832], _096647_);
  or g_106678_(_096634_, _096639_, _096648_);
  or g_106679_(_096635_, _096637_, _096649_);
  or g_106680_(_096640_, _096645_, _096650_);
  or g_106681_(_096649_, _096650_, _096651_);
  or g_106682_(_096638_, _096642_, _096652_);
  or g_106683_(_096646_, _096647_, _096653_);
  or g_106684_(_096652_, _096653_, _096654_);
  or g_106685_(_096651_, _096654_, _096655_);
  xor g_106686_(out[316], out[844], _096656_);
  or g_106687_(_096633_, _096656_, _096657_);
  or g_106688_(_096632_, _096643_, _096658_);
  or g_106689_(_096657_, _096658_, _096659_);
  or g_106690_(_096636_, _096641_, _096660_);
  or g_106691_(_096644_, _096660_, _096661_);
  or g_106692_(_096659_, _096661_, _096662_);
  or g_106693_(_096655_, _096662_, _096663_);
  or g_106694_(_096648_, _096663_, _096664_);
  not g_106695_(_096664_, _096665_);
  xor g_106696_(out[289], out[833], _096666_);
  and g_106697_(out[299], _049741_, _096667_);
  xor g_106698_(out[297], out[841], _096668_);
  xor g_106699_(out[288], out[832], _096669_);
  xor g_106700_(out[302], out[846], _096670_);
  xor g_106701_(out[292], out[836], _096671_);
  or g_106702_(_096670_, _096671_, _096672_);
  xor g_106703_(out[301], out[845], _096673_);
  xor g_106704_(out[291], out[835], _096674_);
  and g_106705_(_098272_, out[843], _096675_);
  xor g_106706_(out[294], out[838], _096676_);
  xor g_106707_(out[298], out[842], _096677_);
  xor g_106708_(out[293], out[837], _096678_);
  xor g_106709_(out[303], out[847], _096679_);
  xor g_106710_(out[296], out[840], _096680_);
  or g_106711_(_096673_, _096680_, _096681_);
  xor g_106712_(out[290], out[834], _096682_);
  or g_106713_(_096677_, _096682_, _096683_);
  or g_106714_(_096681_, _096683_, _096684_);
  or g_106715_(_096668_, _096674_, _096685_);
  or g_106716_(_096678_, _096685_, _096686_);
  or g_106717_(_096684_, _096686_, _096687_);
  or g_106718_(_096672_, _096687_, _096688_);
  xor g_106719_(out[300], out[844], _096689_);
  or g_106720_(_096675_, _096689_, _096690_);
  xor g_106721_(out[295], out[839], _096691_);
  or g_106722_(_096676_, _096691_, _096692_);
  or g_106723_(_096690_, _096692_, _096693_);
  or g_106724_(_096666_, _096667_, _096694_);
  or g_106725_(_096679_, _096694_, _096695_);
  or g_106726_(_096693_, _096695_, _096696_);
  or g_106727_(_096669_, _096696_, _096697_);
  or g_106728_(_096688_, _096697_, _096698_);
  xor g_106729_(out[279], out[839], _096699_);
  and g_106730_(_098261_, out[843], _096700_);
  xor g_106731_(out[286], out[846], _096701_);
  xor g_106732_(out[280], out[840], _096702_);
  xor g_106733_(out[273], out[833], _096703_);
  xor g_106734_(out[285], out[845], _096704_);
  xor g_106735_(out[281], out[841], _096705_);
  xor g_106736_(out[276], out[836], _096706_);
  xor g_106737_(out[274], out[834], _096707_);
  and g_106738_(out[283], _049741_, _096708_);
  xor g_106739_(out[275], out[835], _096709_);
  xor g_106740_(out[278], out[838], _096710_);
  xor g_106741_(out[287], out[847], _096711_);
  xor g_106742_(out[282], out[842], _096712_);
  xor g_106743_(out[277], out[837], _096713_);
  xor g_106744_(out[272], out[832], _096714_);
  or g_106745_(_096701_, _096706_, _096715_);
  or g_106746_(_096702_, _096704_, _096716_);
  or g_106747_(_096707_, _096712_, _096717_);
  or g_106748_(_096716_, _096717_, _096718_);
  or g_106749_(_096705_, _096709_, _096719_);
  or g_106750_(_096713_, _096714_, _096720_);
  or g_106751_(_096719_, _096720_, _096721_);
  or g_106752_(_096718_, _096721_, _096722_);
  xor g_106753_(out[284], out[844], _096723_);
  or g_106754_(_096700_, _096723_, _096724_);
  or g_106755_(_096699_, _096710_, _096725_);
  or g_106756_(_096724_, _096725_, _096726_);
  or g_106757_(_096703_, _096708_, _096727_);
  or g_106758_(_096711_, _096727_, _096728_);
  or g_106759_(_096726_, _096728_, _096729_);
  or g_106760_(_096722_, _096729_, _096730_);
  or g_106761_(_096715_, _096730_, _096731_);
  xor g_106762_(out[269], out[845], _096732_);
  xor g_106763_(out[258], out[834], _096733_);
  xor g_106764_(out[261], out[837], _096734_);
  xor g_106765_(out[265], out[841], _096735_);
  xor g_106766_(out[260], out[836], _096736_);
  xor g_106767_(out[264], out[840], _096737_);
  xor g_106768_(out[270], out[846], _096738_);
  xor g_106769_(out[262], out[838], _096739_);
  xor g_106770_(out[271], out[847], _096740_);
  xor g_106771_(out[266], out[842], _096741_);
  xor g_106772_(out[256], out[832], _096742_);
  xor g_106773_(out[259], out[835], _096743_);
  and g_106774_(_098250_, out[843], _096744_);
  and g_106775_(out[267], _049741_, _096745_);
  xor g_106776_(out[257], out[833], _096746_);
  or g_106777_(_096736_, _096738_, _096747_);
  or g_106778_(_096732_, _096737_, _096748_);
  or g_106779_(_096733_, _096741_, _096749_);
  or g_106780_(_096748_, _096749_, _096750_);
  or g_106781_(_096735_, _096743_, _096751_);
  or g_106782_(_096734_, _096742_, _096752_);
  or g_106783_(_096751_, _096752_, _096753_);
  or g_106784_(_096750_, _096753_, _096754_);
  xor g_106785_(out[268], out[844], _096755_);
  or g_106786_(_096744_, _096755_, _096756_);
  xor g_106787_(out[263], out[839], _096757_);
  or g_106788_(_096739_, _096757_, _096758_);
  or g_106789_(_096756_, _096758_, _096759_);
  or g_106790_(_096745_, _096746_, _096760_);
  or g_106791_(_096740_, _096760_, _096761_);
  or g_106792_(_096759_, _096761_, _096762_);
  or g_106793_(_096754_, _096762_, _096763_);
  or g_106794_(_096747_, _096763_, _096764_);
  not g_106795_(_096764_, _096765_);
  xor g_106796_(out[247], out[839], _096766_);
  and g_106797_(_098239_, out[843], _096767_);
  xor g_106798_(out[254], out[846], _096768_);
  xor g_106799_(out[248], out[840], _096769_);
  xor g_106800_(out[241], out[833], _096770_);
  xor g_106801_(out[253], out[845], _096771_);
  xor g_106802_(out[249], out[841], _096772_);
  xor g_106803_(out[244], out[836], _096773_);
  xor g_106804_(out[242], out[834], _096774_);
  and g_106805_(out[251], _049741_, _096775_);
  xor g_106806_(out[243], out[835], _096776_);
  xor g_106807_(out[246], out[838], _096777_);
  xor g_106808_(out[255], out[847], _096778_);
  xor g_106809_(out[250], out[842], _096779_);
  xor g_106810_(out[245], out[837], _096780_);
  xor g_106811_(out[240], out[832], _096781_);
  or g_106812_(_096768_, _096773_, _096782_);
  or g_106813_(_096769_, _096771_, _096783_);
  or g_106814_(_096774_, _096779_, _096784_);
  or g_106815_(_096783_, _096784_, _096785_);
  or g_106816_(_096772_, _096776_, _096786_);
  or g_106817_(_096780_, _096781_, _096787_);
  or g_106818_(_096786_, _096787_, _096788_);
  or g_106819_(_096785_, _096788_, _096789_);
  xor g_106820_(out[252], out[844], _096790_);
  or g_106821_(_096767_, _096790_, _096791_);
  or g_106822_(_096766_, _096777_, _096792_);
  or g_106823_(_096791_, _096792_, _096793_);
  or g_106824_(_096770_, _096775_, _096794_);
  or g_106825_(_096778_, _096794_, _096795_);
  or g_106826_(_096793_, _096795_, _096796_);
  or g_106827_(_096789_, _096796_, _096797_);
  or g_106828_(_096782_, _096797_, _096798_);
  xor g_106829_(out[236], out[844], _096799_);
  and g_106830_(_098228_, out[843], _096800_);
  xor g_106831_(out[232], out[840], _096801_);
  xor g_106832_(out[230], out[838], _096802_);
  xor g_106833_(out[237], out[845], _096803_);
  xor g_106834_(out[238], out[846], _096804_);
  xor g_106835_(out[226], out[834], _096805_);
  xor g_106836_(out[233], out[841], _096806_);
  xor g_106837_(out[229], out[837], _096807_);
  xor g_106838_(out[225], out[833], _096808_);
  and g_106839_(out[235], _049741_, _096809_);
  or g_106840_(_096801_, _096803_, _096810_);
  xor g_106841_(out[239], out[847], _096811_);
  xor g_106842_(out[234], out[842], _096812_);
  xor g_106843_(out[228], out[836], _096813_);
  xor g_106844_(out[227], out[835], _096814_);
  xor g_106845_(out[224], out[832], _096815_);
  or g_106846_(_096805_, _096812_, _096816_);
  or g_106847_(_096810_, _096816_, _096817_);
  or g_106848_(_096806_, _096814_, _096818_);
  or g_106849_(_096807_, _096818_, _096819_);
  or g_106850_(_096817_, _096819_, _096820_);
  or g_106851_(_096804_, _096813_, _096821_);
  or g_106852_(_096820_, _096821_, _096822_);
  or g_106853_(_096799_, _096800_, _096823_);
  xor g_106854_(out[231], out[839], _096824_);
  or g_106855_(_096802_, _096824_, _096825_);
  or g_106856_(_096823_, _096825_, _096826_);
  or g_106857_(_096808_, _096809_, _096827_);
  or g_106858_(_096811_, _096827_, _096828_);
  or g_106859_(_096826_, _096828_, _096829_);
  or g_106860_(_096815_, _096829_, _096830_);
  or g_106861_(_096822_, _096830_, _096831_);
  xor g_106862_(out[215], out[839], _096832_);
  and g_106863_(_098217_, out[843], _096833_);
  xor g_106864_(out[222], out[846], _096834_);
  xor g_106865_(out[216], out[840], _096835_);
  xor g_106866_(out[209], out[833], _096836_);
  xor g_106867_(out[221], out[845], _096837_);
  xor g_106868_(out[217], out[841], _096838_);
  xor g_106869_(out[212], out[836], _096839_);
  xor g_106870_(out[210], out[834], _096840_);
  and g_106871_(out[219], _049741_, _096841_);
  xor g_106872_(out[211], out[835], _096842_);
  xor g_106873_(out[214], out[838], _096843_);
  xor g_106874_(out[223], out[847], _096844_);
  xor g_106875_(out[218], out[842], _096845_);
  xor g_106876_(out[213], out[837], _096846_);
  xor g_106877_(out[208], out[832], _096847_);
  or g_106878_(_096834_, _096839_, _096848_);
  or g_106879_(_096835_, _096837_, _096849_);
  or g_106880_(_096840_, _096845_, _096850_);
  or g_106881_(_096849_, _096850_, _096851_);
  or g_106882_(_096838_, _096842_, _096852_);
  or g_106883_(_096846_, _096847_, _096853_);
  or g_106884_(_096852_, _096853_, _096854_);
  or g_106885_(_096851_, _096854_, _096855_);
  xor g_106886_(out[220], out[844], _096856_);
  or g_106887_(_096833_, _096856_, _096857_);
  or g_106888_(_096832_, _096843_, _096858_);
  or g_106889_(_096857_, _096858_, _096859_);
  or g_106890_(_096836_, _096841_, _096860_);
  or g_106891_(_096844_, _096860_, _096861_);
  or g_106892_(_096859_, _096861_, _096862_);
  or g_106893_(_096855_, _096862_, _096863_);
  or g_106894_(_096848_, _096863_, _096864_);
  not g_106895_(_096864_, _096865_);
  xor g_106896_(out[193], out[833], _096866_);
  and g_106897_(out[203], _049741_, _096867_);
  xor g_106898_(out[201], out[841], _096868_);
  xor g_106899_(out[192], out[832], _096869_);
  xor g_106900_(out[206], out[846], _096870_);
  xor g_106901_(out[196], out[836], _096871_);
  or g_106902_(_096870_, _096871_, _096872_);
  xor g_106903_(out[205], out[845], _096873_);
  xor g_106904_(out[195], out[835], _096874_);
  and g_106905_(_098206_, out[843], _096875_);
  xor g_106906_(out[198], out[838], _096876_);
  xor g_106907_(out[202], out[842], _096877_);
  xor g_106908_(out[197], out[837], _096878_);
  xor g_106909_(out[207], out[847], _096879_);
  xor g_106910_(out[200], out[840], _096880_);
  or g_106911_(_096873_, _096880_, _096881_);
  xor g_106912_(out[194], out[834], _096882_);
  or g_106913_(_096877_, _096882_, _096883_);
  or g_106914_(_096881_, _096883_, _096884_);
  or g_106915_(_096868_, _096874_, _096885_);
  or g_106916_(_096878_, _096885_, _096886_);
  or g_106917_(_096884_, _096886_, _096887_);
  or g_106918_(_096872_, _096887_, _096888_);
  xor g_106919_(out[204], out[844], _096889_);
  or g_106920_(_096875_, _096889_, _096890_);
  xor g_106921_(out[199], out[839], _096891_);
  or g_106922_(_096876_, _096891_, _096892_);
  or g_106923_(_096890_, _096892_, _096893_);
  or g_106924_(_096866_, _096867_, _096894_);
  or g_106925_(_096879_, _096894_, _096895_);
  or g_106926_(_096893_, _096895_, _096896_);
  or g_106927_(_096869_, _096896_, _096897_);
  or g_106928_(_096888_, _096897_, _096898_);
  xor g_106929_(out[183], out[839], _096899_);
  and g_106930_(_098195_, out[843], _096900_);
  xor g_106931_(out[190], out[846], _096901_);
  xor g_106932_(out[184], out[840], _096902_);
  xor g_106933_(out[177], out[833], _096903_);
  xor g_106934_(out[189], out[845], _096904_);
  xor g_106935_(out[185], out[841], _096905_);
  xor g_106936_(out[180], out[836], _096906_);
  xor g_106937_(out[178], out[834], _096907_);
  and g_106938_(out[187], _049741_, _096908_);
  xor g_106939_(out[179], out[835], _096909_);
  xor g_106940_(out[182], out[838], _096910_);
  xor g_106941_(out[191], out[847], _096911_);
  xor g_106942_(out[186], out[842], _096912_);
  xor g_106943_(out[181], out[837], _096913_);
  xor g_106944_(out[176], out[832], _096914_);
  or g_106945_(_096901_, _096906_, _096915_);
  or g_106946_(_096902_, _096904_, _096916_);
  or g_106947_(_096907_, _096912_, _096917_);
  or g_106948_(_096916_, _096917_, _096918_);
  or g_106949_(_096905_, _096909_, _096919_);
  or g_106950_(_096913_, _096914_, _096920_);
  or g_106951_(_096919_, _096920_, _096921_);
  or g_106952_(_096918_, _096921_, _096922_);
  xor g_106953_(out[188], out[844], _096923_);
  or g_106954_(_096900_, _096923_, _096924_);
  or g_106955_(_096899_, _096910_, _096925_);
  or g_106956_(_096924_, _096925_, _096926_);
  or g_106957_(_096903_, _096908_, _096927_);
  or g_106958_(_096911_, _096927_, _096928_);
  or g_106959_(_096926_, _096928_, _096929_);
  or g_106960_(_096922_, _096929_, _096930_);
  or g_106961_(_096915_, _096930_, _096931_);
  xor g_106962_(out[161], out[833], _096932_);
  and g_106963_(out[171], _049741_, _096933_);
  xor g_106964_(out[174], out[846], _096934_);
  xor g_106965_(out[163], out[835], _096935_);
  xor g_106966_(out[164], out[836], _096936_);
  xor g_106967_(out[162], out[834], _096937_);
  xor g_106968_(out[169], out[841], _096938_);
  xor g_106969_(out[160], out[832], _096939_);
  and g_106970_(_098184_, out[843], _096940_);
  xor g_106971_(out[166], out[838], _096941_);
  xor g_106972_(out[170], out[842], _096942_);
  xor g_106973_(out[165], out[837], _096943_);
  xor g_106974_(out[175], out[847], _096944_);
  xor g_106975_(out[173], out[845], _096945_);
  xor g_106976_(out[168], out[840], _096946_);
  or g_106977_(_096934_, _096936_, _096947_);
  or g_106978_(_096945_, _096946_, _096948_);
  or g_106979_(_096937_, _096942_, _096949_);
  or g_106980_(_096948_, _096949_, _096950_);
  or g_106981_(_096935_, _096938_, _096951_);
  or g_106982_(_096939_, _096943_, _096952_);
  or g_106983_(_096951_, _096952_, _096953_);
  or g_106984_(_096950_, _096953_, _096954_);
  xor g_106985_(out[172], out[844], _096955_);
  or g_106986_(_096940_, _096955_, _096956_);
  xor g_106987_(out[167], out[839], _096957_);
  or g_106988_(_096941_, _096957_, _096958_);
  or g_106989_(_096956_, _096958_, _096959_);
  or g_106990_(_096932_, _096933_, _096960_);
  or g_106991_(_096944_, _096960_, _096961_);
  or g_106992_(_096959_, _096961_, _096962_);
  or g_106993_(_096954_, _096962_, _096963_);
  or g_106994_(_096947_, _096963_, _096964_);
  xor g_106995_(out[151], out[839], _096965_);
  and g_106996_(_098173_, out[843], _096966_);
  xor g_106997_(out[158], out[846], _096967_);
  xor g_106998_(out[152], out[840], _096968_);
  xor g_106999_(out[145], out[833], _096969_);
  xor g_107000_(out[157], out[845], _096970_);
  xor g_107001_(out[153], out[841], _096971_);
  xor g_107002_(out[148], out[836], _096972_);
  xor g_107003_(out[146], out[834], _096973_);
  and g_107004_(out[155], _049741_, _096974_);
  xor g_107005_(out[147], out[835], _096975_);
  xor g_107006_(out[150], out[838], _096976_);
  xor g_107007_(out[159], out[847], _096977_);
  xor g_107008_(out[154], out[842], _096978_);
  xor g_107009_(out[149], out[837], _096979_);
  xor g_107010_(out[144], out[832], _096980_);
  or g_107011_(_096967_, _096972_, _096981_);
  or g_107012_(_096968_, _096970_, _096982_);
  or g_107013_(_096973_, _096978_, _096983_);
  or g_107014_(_096982_, _096983_, _096984_);
  or g_107015_(_096971_, _096975_, _096985_);
  or g_107016_(_096979_, _096980_, _096986_);
  or g_107017_(_096985_, _096986_, _096987_);
  or g_107018_(_096984_, _096987_, _096988_);
  xor g_107019_(out[156], out[844], _096989_);
  or g_107020_(_096966_, _096989_, _096990_);
  or g_107021_(_096965_, _096976_, _096991_);
  or g_107022_(_096990_, _096991_, _096992_);
  or g_107023_(_096969_, _096974_, _096993_);
  or g_107024_(_096977_, _096993_, _096994_);
  or g_107025_(_096992_, _096994_, _096995_);
  or g_107026_(_096988_, _096995_, _096996_);
  or g_107027_(_096981_, _096996_, _096997_);
  xor g_107028_(out[129], out[833], _096998_);
  and g_107029_(out[139], _049741_, _096999_);
  xor g_107030_(out[137], out[841], _097000_);
  xor g_107031_(out[128], out[832], _097001_);
  xor g_107032_(out[142], out[846], _097002_);
  xor g_107033_(out[132], out[836], _097003_);
  or g_107034_(_097002_, _097003_, _097004_);
  xor g_107035_(out[141], out[845], _097005_);
  xor g_107036_(out[131], out[835], _097006_);
  and g_107037_(_098162_, out[843], _097007_);
  xor g_107038_(out[134], out[838], _097008_);
  xor g_107039_(out[138], out[842], _097009_);
  xor g_107040_(out[133], out[837], _097010_);
  xor g_107041_(out[143], out[847], _097011_);
  xor g_107042_(out[136], out[840], _097012_);
  or g_107043_(_097005_, _097012_, _097013_);
  xor g_107044_(out[130], out[834], _097014_);
  or g_107045_(_097009_, _097014_, _097015_);
  or g_107046_(_097013_, _097015_, _097016_);
  or g_107047_(_097000_, _097006_, _097017_);
  or g_107048_(_097010_, _097017_, _097018_);
  or g_107049_(_097016_, _097018_, _097019_);
  or g_107050_(_097004_, _097019_, _097020_);
  xor g_107051_(out[140], out[844], _097021_);
  or g_107052_(_097007_, _097021_, _097022_);
  xor g_107053_(out[135], out[839], _097023_);
  or g_107054_(_097008_, _097023_, _097024_);
  or g_107055_(_097022_, _097024_, _097025_);
  or g_107056_(_096998_, _096999_, _097026_);
  or g_107057_(_097011_, _097026_, _097027_);
  or g_107058_(_097025_, _097027_, _097028_);
  or g_107059_(_097001_, _097028_, _097029_);
  or g_107060_(_097020_, _097029_, _097030_);
  xor g_107061_(out[119], out[839], _097031_);
  and g_107062_(_098151_, out[843], _097032_);
  xor g_107063_(out[126], out[846], _097033_);
  xor g_107064_(out[120], out[840], _097034_);
  xor g_107065_(out[113], out[833], _097035_);
  xor g_107066_(out[125], out[845], _097036_);
  xor g_107067_(out[121], out[841], _097037_);
  xor g_107068_(out[116], out[836], _097038_);
  xor g_107069_(out[114], out[834], _097039_);
  and g_107070_(out[123], _049741_, _097040_);
  xor g_107071_(out[115], out[835], _097041_);
  xor g_107072_(out[118], out[838], _097042_);
  xor g_107073_(out[127], out[847], _097043_);
  xor g_107074_(out[122], out[842], _097044_);
  xor g_107075_(out[117], out[837], _097045_);
  xor g_107076_(out[112], out[832], _097046_);
  or g_107077_(_097033_, _097038_, _097047_);
  or g_107078_(_097034_, _097036_, _097048_);
  or g_107079_(_097039_, _097044_, _097049_);
  or g_107080_(_097048_, _097049_, _097050_);
  or g_107081_(_097037_, _097041_, _097051_);
  or g_107082_(_097045_, _097046_, _097052_);
  or g_107083_(_097051_, _097052_, _097053_);
  or g_107084_(_097050_, _097053_, _097054_);
  xor g_107085_(out[124], out[844], _097055_);
  or g_107086_(_097032_, _097055_, _097056_);
  or g_107087_(_097031_, _097042_, _097057_);
  or g_107088_(_097056_, _097057_, _097058_);
  or g_107089_(_097035_, _097040_, _097059_);
  or g_107090_(_097043_, _097059_, _097060_);
  or g_107091_(_097058_, _097060_, _097061_);
  or g_107092_(_097054_, _097061_, _097062_);
  or g_107093_(_097047_, _097062_, _097063_);
  xor g_107094_(out[97], out[833], _097064_);
  and g_107095_(_098140_, out[843], _097065_);
  and g_107096_(out[107], _049741_, _097066_);
  xor g_107097_(out[104], out[840], _097067_);
  xor g_107098_(out[106], out[842], _097068_);
  xor g_107099_(out[98], out[834], _097069_);
  xor g_107100_(out[100], out[836], _097070_);
  xor g_107101_(out[109], out[845], _097071_);
  xor g_107102_(out[105], out[841], _097072_);
  xor g_107103_(out[99], out[835], _097073_);
  xor g_107104_(out[101], out[837], _097074_);
  xor g_107105_(out[110], out[846], _097075_);
  xor g_107106_(out[96], out[832], _097076_);
  xor g_107107_(out[111], out[847], _097077_);
  or g_107108_(_097067_, _097071_, _097078_);
  xor g_107109_(out[102], out[838], _097079_);
  or g_107110_(_097068_, _097069_, _097080_);
  or g_107111_(_097078_, _097080_, _097081_);
  or g_107112_(_097072_, _097073_, _097082_);
  or g_107113_(_097074_, _097082_, _097083_);
  or g_107114_(_097081_, _097083_, _097084_);
  or g_107115_(_097070_, _097075_, _097085_);
  or g_107116_(_097084_, _097085_, _097086_);
  xor g_107117_(out[108], out[844], _097087_);
  or g_107118_(_097065_, _097087_, _097088_);
  xor g_107119_(out[103], out[839], _097089_);
  or g_107120_(_097079_, _097089_, _097090_);
  or g_107121_(_097088_, _097090_, _097091_);
  or g_107122_(_097064_, _097066_, _097092_);
  or g_107123_(_097077_, _097092_, _097093_);
  or g_107124_(_097091_, _097093_, _097094_);
  or g_107125_(_097076_, _097094_, _097095_);
  or g_107126_(_097086_, _097095_, _097096_);
  not g_107127_(_097096_, _097097_);
  xor g_107128_(out[87], out[839], _097098_);
  and g_107129_(_098129_, out[843], _097099_);
  xor g_107130_(out[94], out[846], _097100_);
  xor g_107131_(out[88], out[840], _097101_);
  xor g_107132_(out[81], out[833], _097102_);
  xor g_107133_(out[93], out[845], _097103_);
  xor g_107134_(out[89], out[841], _097104_);
  xor g_107135_(out[84], out[836], _097105_);
  xor g_107136_(out[82], out[834], _097106_);
  and g_107137_(out[91], _049741_, _097107_);
  xor g_107138_(out[83], out[835], _097108_);
  xor g_107139_(out[86], out[838], _097109_);
  xor g_107140_(out[95], out[847], _097110_);
  xor g_107141_(out[90], out[842], _097111_);
  xor g_107142_(out[85], out[837], _097112_);
  xor g_107143_(out[80], out[832], _097113_);
  or g_107144_(_097100_, _097105_, _097114_);
  or g_107145_(_097101_, _097103_, _097115_);
  or g_107146_(_097106_, _097111_, _097116_);
  or g_107147_(_097115_, _097116_, _097117_);
  or g_107148_(_097104_, _097108_, _097118_);
  or g_107149_(_097112_, _097113_, _097119_);
  or g_107150_(_097118_, _097119_, _097120_);
  or g_107151_(_097117_, _097120_, _097121_);
  xor g_107152_(out[92], out[844], _097122_);
  or g_107153_(_097099_, _097122_, _097123_);
  or g_107154_(_097098_, _097109_, _097124_);
  or g_107155_(_097123_, _097124_, _097125_);
  or g_107156_(_097102_, _097107_, _097126_);
  or g_107157_(_097110_, _097126_, _097127_);
  or g_107158_(_097125_, _097127_, _097128_);
  or g_107159_(_097121_, _097128_, _097129_);
  or g_107160_(_097114_, _097129_, _097130_);
  xor g_107161_(out[74], out[842], _097131_);
  xor g_107162_(out[72], out[840], _097132_);
  xor g_107163_(out[65], out[833], _097133_);
  and g_107164_(_098118_, out[843], _097134_);
  and g_107165_(out[75], _049741_, _097135_);
  xor g_107166_(out[66], out[834], _097136_);
  xor g_107167_(out[69], out[837], _097137_);
  xor g_107168_(out[73], out[841], _097138_);
  xor g_107169_(out[76], out[844], _097139_);
  xor g_107170_(out[77], out[845], _097140_);
  xor g_107171_(out[79], out[847], _097141_);
  xor g_107172_(out[68], out[836], _097142_);
  xor g_107173_(out[70], out[838], _097143_);
  xor g_107174_(out[67], out[835], _097144_);
  xor g_107175_(out[64], out[832], _097145_);
  xor g_107176_(out[78], out[846], _097146_);
  or g_107177_(_097142_, _097146_, _097147_);
  or g_107178_(_097132_, _097140_, _097148_);
  or g_107179_(_097131_, _097136_, _097149_);
  or g_107180_(_097148_, _097149_, _097150_);
  or g_107181_(_097138_, _097144_, _097151_);
  or g_107182_(_097137_, _097145_, _097152_);
  or g_107183_(_097151_, _097152_, _097153_);
  or g_107184_(_097150_, _097153_, _097154_);
  or g_107185_(_097134_, _097139_, _097155_);
  xor g_107186_(out[71], out[839], _097156_);
  or g_107187_(_097143_, _097156_, _097157_);
  or g_107188_(_097155_, _097157_, _097158_);
  or g_107189_(_097133_, _097135_, _097159_);
  or g_107190_(_097141_, _097159_, _097160_);
  or g_107191_(_097158_, _097160_, _097161_);
  or g_107192_(_097154_, _097161_, _097162_);
  or g_107193_(_097147_, _097162_, _097163_);
  xor g_107194_(out[55], out[839], _097164_);
  and g_107195_(_098107_, out[843], _097165_);
  xor g_107196_(out[62], out[846], _097166_);
  xor g_107197_(out[56], out[840], _097167_);
  xor g_107198_(out[49], out[833], _097168_);
  xor g_107199_(out[61], out[845], _097169_);
  xor g_107200_(out[57], out[841], _097170_);
  xor g_107201_(out[52], out[836], _097171_);
  xor g_107202_(out[50], out[834], _097172_);
  and g_107203_(out[59], _049741_, _097173_);
  xor g_107204_(out[51], out[835], _097174_);
  xor g_107205_(out[54], out[838], _097175_);
  xor g_107206_(out[63], out[847], _097176_);
  xor g_107207_(out[58], out[842], _097177_);
  xor g_107208_(out[53], out[837], _097178_);
  xor g_107209_(out[48], out[832], _097179_);
  or g_107210_(_097166_, _097171_, _097180_);
  or g_107211_(_097167_, _097169_, _097181_);
  or g_107212_(_097172_, _097177_, _097182_);
  or g_107213_(_097181_, _097182_, _097183_);
  or g_107214_(_097170_, _097174_, _097184_);
  or g_107215_(_097178_, _097179_, _097185_);
  or g_107216_(_097184_, _097185_, _097186_);
  or g_107217_(_097183_, _097186_, _097187_);
  xor g_107218_(out[60], out[844], _097188_);
  or g_107219_(_097165_, _097188_, _097189_);
  or g_107220_(_097164_, _097175_, _097190_);
  or g_107221_(_097189_, _097190_, _097191_);
  or g_107222_(_097168_, _097173_, _097192_);
  or g_107223_(_097176_, _097192_, _097193_);
  or g_107224_(_097191_, _097193_, _097194_);
  or g_107225_(_097187_, _097194_, _097195_);
  or g_107226_(_097180_, _097195_, _097196_);
  not g_107227_(_097196_, _097197_);
  xor g_107228_(out[33], out[833], _097198_);
  and g_107229_(out[43], _049741_, _097199_);
  xor g_107230_(out[41], out[841], _097200_);
  xor g_107231_(out[32], out[832], _097201_);
  xor g_107232_(out[46], out[846], _097202_);
  xor g_107233_(out[36], out[836], _097203_);
  or g_107234_(_097202_, _097203_, _097204_);
  xor g_107235_(out[45], out[845], _097205_);
  xor g_107236_(out[35], out[835], _097206_);
  and g_107237_(_098096_, out[843], _097207_);
  xor g_107238_(out[38], out[838], _097208_);
  xor g_107239_(out[42], out[842], _097209_);
  xor g_107240_(out[37], out[837], _097210_);
  xor g_107241_(out[47], out[847], _097211_);
  xor g_107242_(out[40], out[840], _097212_);
  or g_107243_(_097205_, _097212_, _097213_);
  xor g_107244_(out[34], out[834], _097214_);
  or g_107245_(_097209_, _097214_, _097215_);
  or g_107246_(_097213_, _097215_, _097216_);
  or g_107247_(_097200_, _097206_, _097217_);
  or g_107248_(_097210_, _097217_, _097218_);
  or g_107249_(_097216_, _097218_, _097219_);
  or g_107250_(_097204_, _097219_, _097220_);
  xor g_107251_(out[44], out[844], _097221_);
  or g_107252_(_097207_, _097221_, _097222_);
  xor g_107253_(out[39], out[839], _097223_);
  or g_107254_(_097208_, _097223_, _097224_);
  or g_107255_(_097222_, _097224_, _097225_);
  or g_107256_(_097198_, _097199_, _097226_);
  or g_107257_(_097211_, _097226_, _097227_);
  or g_107258_(_097225_, _097227_, _097228_);
  or g_107259_(_097201_, _097228_, _097229_);
  or g_107260_(_097220_, _097229_, _097230_);
  xor g_107261_(out[23], out[839], _097231_);
  and g_107262_(_098063_, out[843], _097232_);
  xor g_107263_(out[30], out[846], _097233_);
  xor g_107264_(out[24], out[840], _097234_);
  xor g_107265_(out[17], out[833], _097235_);
  xor g_107266_(out[29], out[845], _097236_);
  xor g_107267_(out[25], out[841], _097237_);
  xor g_107268_(out[20], out[836], _097238_);
  xor g_107269_(out[18], out[834], _097239_);
  and g_107270_(out[27], _049741_, _097240_);
  xor g_107271_(out[19], out[835], _097241_);
  xor g_107272_(out[22], out[838], _097242_);
  xor g_107273_(out[31], out[847], _097243_);
  xor g_107274_(out[26], out[842], _097244_);
  xor g_107275_(out[21], out[837], _097245_);
  xor g_107276_(out[16], out[832], _097246_);
  or g_107277_(_097233_, _097238_, _097247_);
  or g_107278_(_097234_, _097236_, _097248_);
  or g_107279_(_097239_, _097244_, _097249_);
  or g_107280_(_097248_, _097249_, _097250_);
  or g_107281_(_097237_, _097241_, _097251_);
  or g_107282_(_097245_, _097246_, _097252_);
  or g_107283_(_097251_, _097252_, _097253_);
  or g_107284_(_097250_, _097253_, _097254_);
  xor g_107285_(out[28], out[844], _097255_);
  or g_107286_(_097232_, _097255_, _097256_);
  or g_107287_(_097231_, _097242_, _097257_);
  or g_107288_(_097256_, _097257_, _097258_);
  or g_107289_(_097235_, _097240_, _097259_);
  or g_107290_(_097243_, _097259_, _097260_);
  or g_107291_(_097258_, _097260_, _097261_);
  or g_107292_(_097254_, _097261_, _097262_);
  or g_107293_(_097247_, _097262_, _097263_);
  xor g_107294_(out[10], out[842], _097264_);
  xor g_107295_(out[2], out[834], _097265_);
  xor g_107296_(out[1], out[833], _097266_);
  and g_107297_(_098041_, out[843], _097267_);
  and g_107298_(out[11], _049741_, _097268_);
  xor g_107299_(out[13], out[845], _097269_);
  xor g_107300_(out[3], out[835], _097270_);
  xor g_107301_(out[14], out[846], _097271_);
  xor g_107302_(out[12], out[844], _097272_);
  xor g_107303_(out[8], out[840], _097273_);
  xor g_107304_(out[15], out[847], _097274_);
  xor g_107305_(out[5], out[837], _097275_);
  xor g_107306_(out[6], out[838], _097276_);
  xor g_107307_(out[0], out[832], _097277_);
  xor g_107308_(out[4], out[836], _097278_);
  or g_107309_(_097269_, _097273_, _097279_);
  xor g_107310_(out[9], out[841], _097280_);
  or g_107311_(_097264_, _097265_, _097281_);
  or g_107312_(_097279_, _097281_, _097282_);
  or g_107313_(_097270_, _097280_, _097283_);
  or g_107314_(_097275_, _097283_, _097284_);
  or g_107315_(_097282_, _097284_, _097285_);
  or g_107316_(_097271_, _097278_, _097286_);
  or g_107317_(_097285_, _097286_, _097287_);
  or g_107318_(_097267_, _097272_, _097288_);
  xor g_107319_(out[7], out[839], _097289_);
  or g_107320_(_097276_, _097289_, _097290_);
  or g_107321_(_097288_, _097290_, _097291_);
  or g_107322_(_097266_, _097268_, _097292_);
  or g_107323_(_097274_, _097292_, _097293_);
  or g_107324_(_097291_, _097293_, _097294_);
  or g_107325_(_097277_, _097294_, _097295_);
  or g_107326_(_097287_, _097295_, _097296_);
  not g_107327_(_097296_, _097297_);
  and g_107328_(out[475], _049730_, _097298_);
  xor g_107329_(out[468], out[820], _097299_);
  xor g_107330_(out[478], out[830], _097300_);
  or g_107331_(_097299_, _097300_, _097301_);
  xor g_107332_(out[477], out[829], _097302_);
  xor g_107333_(out[467], out[819], _097303_);
  xor g_107334_(out[464], out[816], _097304_);
  and g_107335_(_049499_, out[827], _097305_);
  xor g_107336_(out[474], out[826], _097306_);
  xor g_107337_(out[479], out[831], _097307_);
  xor g_107338_(out[470], out[822], _097308_);
  xor g_107339_(out[469], out[821], _097309_);
  xor g_107340_(out[472], out[824], _097310_);
  or g_107341_(_097302_, _097310_, _097311_);
  xor g_107342_(out[466], out[818], _097312_);
  xor g_107343_(out[473], out[825], _097313_);
  xor g_107344_(out[465], out[817], _097314_);
  or g_107345_(_097306_, _097312_, _097315_);
  or g_107346_(_097311_, _097315_, _097316_);
  or g_107347_(_097303_, _097313_, _097317_);
  or g_107348_(_097309_, _097317_, _097318_);
  or g_107349_(_097316_, _097318_, _097319_);
  or g_107350_(_097301_, _097319_, _097320_);
  xor g_107351_(out[476], out[828], _097321_);
  or g_107352_(_097305_, _097321_, _097322_);
  xor g_107353_(out[471], out[823], _097323_);
  or g_107354_(_097308_, _097323_, _097324_);
  or g_107355_(_097322_, _097324_, _097325_);
  or g_107356_(_097298_, _097314_, _097326_);
  or g_107357_(_097307_, _097326_, _097327_);
  or g_107358_(_097325_, _097327_, _097328_);
  or g_107359_(_097304_, _097328_, _097329_);
  or g_107360_(_097320_, _097329_, _097330_);
  xor g_107361_(out[455], out[823], _097331_);
  and g_107362_(_049477_, out[827], _097332_);
  xor g_107363_(out[462], out[830], _097333_);
  xor g_107364_(out[456], out[824], _097334_);
  xor g_107365_(out[449], out[817], _097335_);
  xor g_107366_(out[461], out[829], _097336_);
  xor g_107367_(out[457], out[825], _097337_);
  xor g_107368_(out[452], out[820], _097338_);
  xor g_107369_(out[450], out[818], _097339_);
  and g_107370_(out[459], _049730_, _097340_);
  xor g_107371_(out[451], out[819], _097341_);
  xor g_107372_(out[454], out[822], _097342_);
  xor g_107373_(out[463], out[831], _097343_);
  xor g_107374_(out[458], out[826], _097344_);
  xor g_107375_(out[453], out[821], _097345_);
  xor g_107376_(out[448], out[816], _097346_);
  or g_107377_(_097333_, _097338_, _097347_);
  or g_107378_(_097334_, _097336_, _097348_);
  or g_107379_(_097339_, _097344_, _097349_);
  or g_107380_(_097348_, _097349_, _097350_);
  or g_107381_(_097337_, _097341_, _097351_);
  or g_107382_(_097345_, _097346_, _097352_);
  or g_107383_(_097351_, _097352_, _097353_);
  or g_107384_(_097350_, _097353_, _097354_);
  xor g_107385_(out[460], out[828], _097355_);
  or g_107386_(_097332_, _097355_, _097356_);
  or g_107387_(_097331_, _097342_, _097357_);
  or g_107388_(_097356_, _097357_, _097358_);
  or g_107389_(_097335_, _097340_, _097359_);
  or g_107390_(_097343_, _097359_, _097360_);
  or g_107391_(_097358_, _097360_, _097361_);
  or g_107392_(_097354_, _097361_, _097362_);
  or g_107393_(_097347_, _097362_, _097363_);
  xor g_107394_(out[434], out[818], _097364_);
  xor g_107395_(out[432], out[816], _097365_);
  xor g_107396_(out[441], out[825], _097366_);
  xor g_107397_(out[440], out[824], _097367_);
  xor g_107398_(out[437], out[821], _097368_);
  xor g_107399_(out[446], out[830], _097369_);
  xor g_107400_(out[445], out[829], _097370_);
  xor g_107401_(out[447], out[831], _097371_);
  xor g_107402_(out[442], out[826], _097372_);
  xor g_107403_(out[438], out[822], _097373_);
  xor g_107404_(out[435], out[819], _097374_);
  and g_107405_(_049466_, out[827], _097375_);
  and g_107406_(out[443], _049730_, _097376_);
  xor g_107407_(out[436], out[820], _097377_);
  xor g_107408_(out[433], out[817], _097378_);
  or g_107409_(_097369_, _097377_, _097379_);
  or g_107410_(_097367_, _097370_, _097380_);
  or g_107411_(_097364_, _097372_, _097381_);
  or g_107412_(_097380_, _097381_, _097382_);
  or g_107413_(_097366_, _097374_, _097383_);
  or g_107414_(_097365_, _097368_, _097384_);
  or g_107415_(_097383_, _097384_, _097385_);
  or g_107416_(_097382_, _097385_, _097386_);
  xor g_107417_(out[444], out[828], _097387_);
  or g_107418_(_097375_, _097387_, _097388_);
  xor g_107419_(out[439], out[823], _097389_);
  or g_107420_(_097373_, _097389_, _097390_);
  or g_107421_(_097388_, _097390_, _097391_);
  or g_107422_(_097376_, _097378_, _097392_);
  or g_107423_(_097371_, _097392_, _097393_);
  or g_107424_(_097391_, _097393_, _097394_);
  or g_107425_(_097386_, _097394_, _097395_);
  or g_107426_(_097379_, _097395_, _097396_);
  not g_107427_(_097396_, _097397_);
  xor g_107428_(out[423], out[823], _097398_);
  and g_107429_(_049455_, out[827], _097399_);
  xor g_107430_(out[430], out[830], _097400_);
  xor g_107431_(out[424], out[824], _097401_);
  xor g_107432_(out[417], out[817], _097402_);
  xor g_107433_(out[429], out[829], _097403_);
  xor g_107434_(out[425], out[825], _097404_);
  xor g_107435_(out[420], out[820], _097405_);
  xor g_107436_(out[418], out[818], _097406_);
  and g_107437_(out[427], _049730_, _097407_);
  xor g_107438_(out[419], out[819], _097408_);
  xor g_107439_(out[422], out[822], _097409_);
  xor g_107440_(out[431], out[831], _097410_);
  xor g_107441_(out[426], out[826], _097411_);
  xor g_107442_(out[421], out[821], _097412_);
  xor g_107443_(out[416], out[816], _097413_);
  or g_107444_(_097400_, _097405_, _097414_);
  or g_107445_(_097401_, _097403_, _097415_);
  or g_107446_(_097406_, _097411_, _097416_);
  or g_107447_(_097415_, _097416_, _097417_);
  or g_107448_(_097404_, _097408_, _097418_);
  or g_107449_(_097412_, _097413_, _097419_);
  or g_107450_(_097418_, _097419_, _097420_);
  or g_107451_(_097417_, _097420_, _097421_);
  xor g_107452_(out[428], out[828], _097422_);
  or g_107453_(_097399_, _097422_, _097423_);
  or g_107454_(_097398_, _097409_, _097424_);
  or g_107455_(_097423_, _097424_, _097425_);
  or g_107456_(_097402_, _097407_, _097426_);
  or g_107457_(_097410_, _097426_, _097427_);
  or g_107458_(_097425_, _097427_, _097428_);
  or g_107459_(_097421_, _097428_, _097429_);
  or g_107460_(_097414_, _097429_, _097430_);
  not g_107461_(_097430_, _097431_);
  xor g_107462_(out[412], out[828], _097432_);
  and g_107463_(_049444_, out[827], _097433_);
  xor g_107464_(out[408], out[824], _097434_);
  xor g_107465_(out[406], out[822], _097435_);
  xor g_107466_(out[413], out[829], _097436_);
  xor g_107467_(out[414], out[830], _097437_);
  xor g_107468_(out[402], out[818], _097438_);
  xor g_107469_(out[409], out[825], _097439_);
  xor g_107470_(out[405], out[821], _097440_);
  xor g_107471_(out[401], out[817], _097441_);
  and g_107472_(out[411], _049730_, _097442_);
  or g_107473_(_097434_, _097436_, _097443_);
  xor g_107474_(out[415], out[831], _097444_);
  xor g_107475_(out[410], out[826], _097445_);
  xor g_107476_(out[404], out[820], _097446_);
  xor g_107477_(out[403], out[819], _097447_);
  xor g_107478_(out[400], out[816], _097448_);
  or g_107479_(_097438_, _097445_, _097449_);
  or g_107480_(_097443_, _097449_, _097450_);
  or g_107481_(_097439_, _097447_, _097451_);
  or g_107482_(_097440_, _097451_, _097452_);
  or g_107483_(_097450_, _097452_, _097453_);
  or g_107484_(_097437_, _097446_, _097454_);
  or g_107485_(_097453_, _097454_, _097455_);
  or g_107486_(_097432_, _097433_, _097456_);
  xor g_107487_(out[407], out[823], _097457_);
  or g_107488_(_097435_, _097457_, _097458_);
  or g_107489_(_097456_, _097458_, _097459_);
  or g_107490_(_097441_, _097442_, _097460_);
  or g_107491_(_097444_, _097460_, _097461_);
  or g_107492_(_097459_, _097461_, _097462_);
  or g_107493_(_097448_, _097462_, _097463_);
  or g_107494_(_097455_, _097463_, _097464_);
  xor g_107495_(out[391], out[823], _097465_);
  and g_107496_(_049433_, out[827], _097466_);
  xor g_107497_(out[398], out[830], _097467_);
  xor g_107498_(out[392], out[824], _097468_);
  xor g_107499_(out[385], out[817], _097469_);
  xor g_107500_(out[397], out[829], _097470_);
  xor g_107501_(out[393], out[825], _097471_);
  xor g_107502_(out[388], out[820], _097472_);
  xor g_107503_(out[386], out[818], _097473_);
  and g_107504_(out[395], _049730_, _097474_);
  xor g_107505_(out[387], out[819], _097475_);
  xor g_107506_(out[390], out[822], _097476_);
  xor g_107507_(out[399], out[831], _097477_);
  xor g_107508_(out[394], out[826], _097478_);
  xor g_107509_(out[389], out[821], _097479_);
  xor g_107510_(out[384], out[816], _097480_);
  or g_107511_(_097467_, _097472_, _097481_);
  or g_107512_(_097468_, _097470_, _097482_);
  or g_107513_(_097473_, _097478_, _097483_);
  or g_107514_(_097482_, _097483_, _097484_);
  or g_107515_(_097471_, _097475_, _097485_);
  or g_107516_(_097479_, _097480_, _097486_);
  or g_107517_(_097485_, _097486_, _097487_);
  or g_107518_(_097484_, _097487_, _097488_);
  xor g_107519_(out[396], out[828], _097489_);
  or g_107520_(_097466_, _097489_, _097490_);
  or g_107521_(_097465_, _097476_, _097491_);
  or g_107522_(_097490_, _097491_, _097492_);
  or g_107523_(_097469_, _097474_, _097493_);
  or g_107524_(_097477_, _097493_, _097494_);
  or g_107525_(_097492_, _097494_, _097495_);
  or g_107526_(_097488_, _097495_, _097496_);
  or g_107527_(_097481_, _097496_, _097497_);
  xor g_107528_(out[369], out[817], _097498_);
  and g_107529_(out[379], _049730_, _097499_);
  xor g_107530_(out[377], out[825], _097500_);
  xor g_107531_(out[368], out[816], _097501_);
  xor g_107532_(out[382], out[830], _097502_);
  xor g_107533_(out[372], out[820], _097503_);
  or g_107534_(_097502_, _097503_, _097504_);
  xor g_107535_(out[381], out[829], _097505_);
  xor g_107536_(out[371], out[819], _097506_);
  and g_107537_(_049422_, out[827], _097507_);
  xor g_107538_(out[374], out[822], _097508_);
  xor g_107539_(out[378], out[826], _097509_);
  xor g_107540_(out[373], out[821], _097510_);
  xor g_107541_(out[383], out[831], _097511_);
  xor g_107542_(out[376], out[824], _097512_);
  or g_107543_(_097505_, _097512_, _097513_);
  xor g_107544_(out[370], out[818], _097514_);
  or g_107545_(_097509_, _097514_, _097515_);
  or g_107546_(_097513_, _097515_, _097516_);
  or g_107547_(_097500_, _097506_, _097517_);
  or g_107548_(_097510_, _097517_, _097518_);
  or g_107549_(_097516_, _097518_, _097519_);
  or g_107550_(_097504_, _097519_, _097520_);
  xor g_107551_(out[380], out[828], _097521_);
  or g_107552_(_097507_, _097521_, _097522_);
  xor g_107553_(out[375], out[823], _097523_);
  or g_107554_(_097508_, _097523_, _097524_);
  or g_107555_(_097522_, _097524_, _097525_);
  or g_107556_(_097498_, _097499_, _097526_);
  or g_107557_(_097511_, _097526_, _097527_);
  or g_107558_(_097525_, _097527_, _097528_);
  or g_107559_(_097501_, _097528_, _097529_);
  or g_107560_(_097520_, _097529_, _097530_);
  xor g_107561_(out[359], out[823], _097531_);
  and g_107562_(_049411_, out[827], _097532_);
  xor g_107563_(out[366], out[830], _097533_);
  xor g_107564_(out[360], out[824], _097534_);
  xor g_107565_(out[353], out[817], _097535_);
  xor g_107566_(out[365], out[829], _097536_);
  xor g_107567_(out[361], out[825], _097537_);
  xor g_107568_(out[356], out[820], _097538_);
  xor g_107569_(out[354], out[818], _097539_);
  and g_107570_(out[363], _049730_, _097540_);
  xor g_107571_(out[355], out[819], _097541_);
  xor g_107572_(out[358], out[822], _097542_);
  xor g_107573_(out[367], out[831], _097543_);
  xor g_107574_(out[362], out[826], _097544_);
  xor g_107575_(out[357], out[821], _097545_);
  xor g_107576_(out[352], out[816], _097546_);
  or g_107577_(_097533_, _097538_, _097547_);
  or g_107578_(_097534_, _097536_, _097548_);
  or g_107579_(_097539_, _097544_, _097549_);
  or g_107580_(_097548_, _097549_, _097550_);
  or g_107581_(_097537_, _097541_, _097551_);
  or g_107582_(_097545_, _097546_, _097552_);
  or g_107583_(_097551_, _097552_, _097553_);
  or g_107584_(_097550_, _097553_, _097554_);
  xor g_107585_(out[364], out[828], _097555_);
  or g_107586_(_097532_, _097555_, _097556_);
  or g_107587_(_097531_, _097542_, _097557_);
  or g_107588_(_097556_, _097557_, _097558_);
  or g_107589_(_097535_, _097540_, _097559_);
  or g_107590_(_097543_, _097559_, _097560_);
  or g_107591_(_097558_, _097560_, _097561_);
  or g_107592_(_097554_, _097561_, _097562_);
  or g_107593_(_097547_, _097562_, _097563_);
  and g_107594_(out[347], _049730_, _097564_);
  xor g_107595_(out[340], out[820], _097565_);
  xor g_107596_(out[350], out[830], _097566_);
  or g_107597_(_097565_, _097566_, _097567_);
  xor g_107598_(out[349], out[829], _097568_);
  xor g_107599_(out[339], out[819], _097569_);
  xor g_107600_(out[336], out[816], _097570_);
  and g_107601_(_049400_, out[827], _097571_);
  xor g_107602_(out[346], out[826], _097572_);
  xor g_107603_(out[351], out[831], _097573_);
  xor g_107604_(out[342], out[822], _097574_);
  xor g_107605_(out[341], out[821], _097575_);
  xor g_107606_(out[344], out[824], _097576_);
  or g_107607_(_097568_, _097576_, _097577_);
  xor g_107608_(out[338], out[818], _097578_);
  xor g_107609_(out[345], out[825], _097579_);
  xor g_107610_(out[337], out[817], _097580_);
  or g_107611_(_097572_, _097578_, _097581_);
  or g_107612_(_097577_, _097581_, _097582_);
  or g_107613_(_097569_, _097579_, _097583_);
  or g_107614_(_097575_, _097583_, _097584_);
  or g_107615_(_097582_, _097584_, _097585_);
  or g_107616_(_097567_, _097585_, _097586_);
  xor g_107617_(out[348], out[828], _097587_);
  or g_107618_(_097571_, _097587_, _097588_);
  xor g_107619_(out[343], out[823], _097589_);
  or g_107620_(_097574_, _097589_, _097590_);
  or g_107621_(_097588_, _097590_, _097591_);
  or g_107622_(_097564_, _097580_, _097592_);
  or g_107623_(_097573_, _097592_, _097593_);
  or g_107624_(_097591_, _097593_, _097594_);
  or g_107625_(_097570_, _097594_, _097595_);
  or g_107626_(_097586_, _097595_, _097596_);
  xor g_107627_(out[327], out[823], _097597_);
  and g_107628_(_098294_, out[827], _097598_);
  xor g_107629_(out[334], out[830], _097599_);
  xor g_107630_(out[328], out[824], _097600_);
  xor g_107631_(out[321], out[817], _097601_);
  xor g_107632_(out[333], out[829], _097602_);
  xor g_107633_(out[329], out[825], _097603_);
  xor g_107634_(out[324], out[820], _097604_);
  xor g_107635_(out[322], out[818], _097605_);
  and g_107636_(out[331], _049730_, _097606_);
  xor g_107637_(out[323], out[819], _097607_);
  xor g_107638_(out[326], out[822], _097608_);
  xor g_107639_(out[335], out[831], _097609_);
  xor g_107640_(out[330], out[826], _097610_);
  xor g_107641_(out[325], out[821], _097611_);
  xor g_107642_(out[320], out[816], _097612_);
  or g_107643_(_097599_, _097604_, _097613_);
  or g_107644_(_097600_, _097602_, _097614_);
  or g_107645_(_097605_, _097610_, _097615_);
  or g_107646_(_097614_, _097615_, _097616_);
  or g_107647_(_097603_, _097607_, _097617_);
  or g_107648_(_097611_, _097612_, _097618_);
  or g_107649_(_097617_, _097618_, _097619_);
  or g_107650_(_097616_, _097619_, _097620_);
  xor g_107651_(out[332], out[828], _097621_);
  or g_107652_(_097598_, _097621_, _097622_);
  or g_107653_(_097597_, _097608_, _097623_);
  or g_107654_(_097622_, _097623_, _097624_);
  or g_107655_(_097601_, _097606_, _097625_);
  or g_107656_(_097609_, _097625_, _097626_);
  or g_107657_(_097624_, _097626_, _097627_);
  or g_107658_(_097620_, _097627_, _097628_);
  or g_107659_(_097613_, _097628_, _097629_);
  xor g_107660_(out[316], out[828], _097630_);
  and g_107661_(_098283_, out[827], _097631_);
  xor g_107662_(out[312], out[824], _097632_);
  xor g_107663_(out[310], out[822], _097633_);
  xor g_107664_(out[317], out[829], _097634_);
  xor g_107665_(out[318], out[830], _097635_);
  xor g_107666_(out[306], out[818], _097636_);
  xor g_107667_(out[313], out[825], _097637_);
  xor g_107668_(out[309], out[821], _097638_);
  xor g_107669_(out[305], out[817], _097639_);
  and g_107670_(out[315], _049730_, _097640_);
  or g_107671_(_097632_, _097634_, _097641_);
  xor g_107672_(out[319], out[831], _097642_);
  xor g_107673_(out[314], out[826], _097643_);
  xor g_107674_(out[308], out[820], _097644_);
  xor g_107675_(out[307], out[819], _097645_);
  xor g_107676_(out[304], out[816], _097646_);
  or g_107677_(_097636_, _097643_, _097647_);
  or g_107678_(_097641_, _097647_, _097648_);
  or g_107679_(_097637_, _097645_, _097649_);
  or g_107680_(_097638_, _097649_, _097650_);
  or g_107681_(_097648_, _097650_, _097651_);
  or g_107682_(_097635_, _097644_, _097652_);
  or g_107683_(_097651_, _097652_, _097653_);
  or g_107684_(_097630_, _097631_, _097654_);
  xor g_107685_(out[311], out[823], _097655_);
  or g_107686_(_097633_, _097655_, _097656_);
  or g_107687_(_097654_, _097656_, _097657_);
  or g_107688_(_097639_, _097640_, _097658_);
  or g_107689_(_097642_, _097658_, _097659_);
  or g_107690_(_097657_, _097659_, _097660_);
  or g_107691_(_097646_, _097660_, _097661_);
  or g_107692_(_097653_, _097661_, _097662_);
  not g_107693_(_097662_, _097663_);
  xor g_107694_(out[295], out[823], _097664_);
  and g_107695_(_098272_, out[827], _097665_);
  xor g_107696_(out[302], out[830], _097666_);
  xor g_107697_(out[296], out[824], _097667_);
  xor g_107698_(out[289], out[817], _097668_);
  xor g_107699_(out[301], out[829], _097669_);
  xor g_107700_(out[297], out[825], _097670_);
  xor g_107701_(out[292], out[820], _097671_);
  xor g_107702_(out[290], out[818], _097672_);
  and g_107703_(out[299], _049730_, _097673_);
  xor g_107704_(out[291], out[819], _097674_);
  xor g_107705_(out[294], out[822], _097675_);
  xor g_107706_(out[303], out[831], _097676_);
  xor g_107707_(out[298], out[826], _097677_);
  xor g_107708_(out[293], out[821], _097678_);
  xor g_107709_(out[288], out[816], _097679_);
  or g_107710_(_097666_, _097671_, _097680_);
  or g_107711_(_097667_, _097669_, _097681_);
  or g_107712_(_097672_, _097677_, _097682_);
  or g_107713_(_097681_, _097682_, _097683_);
  or g_107714_(_097670_, _097674_, _097684_);
  or g_107715_(_097678_, _097679_, _097685_);
  or g_107716_(_097684_, _097685_, _097686_);
  or g_107717_(_097683_, _097686_, _097687_);
  xor g_107718_(out[300], out[828], _097688_);
  or g_107719_(_097665_, _097688_, _097689_);
  or g_107720_(_097664_, _097675_, _097690_);
  or g_107721_(_097689_, _097690_, _097691_);
  or g_107722_(_097668_, _097673_, _097692_);
  or g_107723_(_097676_, _097692_, _097693_);
  or g_107724_(_097691_, _097693_, _097694_);
  or g_107725_(_097687_, _097694_, _097695_);
  or g_107726_(_097680_, _097695_, _097696_);
  not g_107727_(_097696_, _097697_);
  xor g_107728_(out[282], out[826], _097698_);
  xor g_107729_(out[274], out[818], _097699_);
  xor g_107730_(out[273], out[817], _097700_);
  and g_107731_(_098261_, out[827], _097701_);
  and g_107732_(out[283], _049730_, _097702_);
  xor g_107733_(out[285], out[829], _097703_);
  xor g_107734_(out[275], out[819], _097704_);
  xor g_107735_(out[286], out[830], _097705_);
  xor g_107736_(out[284], out[828], _097706_);
  xor g_107737_(out[280], out[824], _097707_);
  xor g_107738_(out[287], out[831], _097708_);
  xor g_107739_(out[277], out[821], _097709_);
  xor g_107740_(out[278], out[822], _097710_);
  xor g_107741_(out[272], out[816], _097711_);
  xor g_107742_(out[276], out[820], _097712_);
  or g_107743_(_097703_, _097707_, _097713_);
  xor g_107744_(out[281], out[825], _097714_);
  or g_107745_(_097698_, _097699_, _097715_);
  or g_107746_(_097713_, _097715_, _097716_);
  or g_107747_(_097704_, _097714_, _097717_);
  or g_107748_(_097709_, _097717_, _097718_);
  or g_107749_(_097716_, _097718_, _097719_);
  or g_107750_(_097705_, _097712_, _097720_);
  or g_107751_(_097719_, _097720_, _097721_);
  or g_107752_(_097701_, _097706_, _097722_);
  xor g_107753_(out[279], out[823], _097723_);
  or g_107754_(_097710_, _097723_, _097724_);
  or g_107755_(_097722_, _097724_, _097725_);
  or g_107756_(_097700_, _097702_, _097726_);
  or g_107757_(_097708_, _097726_, _097727_);
  or g_107758_(_097725_, _097727_, _097728_);
  or g_107759_(_097711_, _097728_, _097729_);
  or g_107760_(_097721_, _097729_, _097730_);
  not g_107761_(_097730_, _097731_);
  xor g_107762_(out[263], out[823], _097732_);
  and g_107763_(_098250_, out[827], _097733_);
  xor g_107764_(out[270], out[830], _097734_);
  xor g_107765_(out[264], out[824], _097735_);
  xor g_107766_(out[257], out[817], _097736_);
  xor g_107767_(out[269], out[829], _097737_);
  xor g_107768_(out[265], out[825], _097738_);
  xor g_107769_(out[260], out[820], _097739_);
  xor g_107770_(out[258], out[818], _097740_);
  and g_107771_(out[267], _049730_, _097741_);
  xor g_107772_(out[259], out[819], _097742_);
  xor g_107773_(out[262], out[822], _097743_);
  xor g_107774_(out[271], out[831], _097744_);
  xor g_107775_(out[266], out[826], _097745_);
  xor g_107776_(out[261], out[821], _097746_);
  xor g_107777_(out[256], out[816], _097747_);
  or g_107778_(_097734_, _097739_, _097748_);
  or g_107779_(_097735_, _097737_, _097749_);
  or g_107780_(_097740_, _097745_, _097750_);
  or g_107781_(_097749_, _097750_, _097751_);
  or g_107782_(_097738_, _097742_, _097752_);
  or g_107783_(_097746_, _097747_, _097753_);
  or g_107784_(_097752_, _097753_, _097754_);
  or g_107785_(_097751_, _097754_, _097755_);
  xor g_107786_(out[268], out[828], _097756_);
  or g_107787_(_097733_, _097756_, _097757_);
  or g_107788_(_097732_, _097743_, _097758_);
  or g_107789_(_097757_, _097758_, _097759_);
  or g_107790_(_097736_, _097741_, _097760_);
  or g_107791_(_097744_, _097760_, _097761_);
  or g_107792_(_097759_, _097761_, _097762_);
  or g_107793_(_097755_, _097762_, _097763_);
  or g_107794_(_097748_, _097763_, _097764_);
  xor g_107795_(out[248], out[824], _097765_);
  xor g_107796_(out[245], out[821], _097766_);
  xor g_107797_(out[243], out[819], _097767_);
  xor g_107798_(out[254], out[830], _097768_);
  xor g_107799_(out[253], out[829], _097769_);
  xor g_107800_(out[242], out[818], _097770_);
  xor g_107801_(out[249], out[825], _097771_);
  xor g_107802_(out[246], out[822], _097772_);
  xor g_107803_(out[255], out[831], _097773_);
  xor g_107804_(out[250], out[826], _097774_);
  xor g_107805_(out[244], out[820], _097775_);
  xor g_107806_(out[240], out[816], _097776_);
  and g_107807_(_098239_, out[827], _097777_);
  and g_107808_(out[251], _049730_, _097778_);
  or g_107809_(_097765_, _097769_, _097779_);
  xor g_107810_(out[241], out[817], _097780_);
  or g_107811_(_097770_, _097774_, _097781_);
  or g_107812_(_097779_, _097781_, _097782_);
  or g_107813_(_097767_, _097771_, _097783_);
  or g_107814_(_097766_, _097783_, _097784_);
  or g_107815_(_097782_, _097784_, _097785_);
  or g_107816_(_097768_, _097775_, _097786_);
  or g_107817_(_097785_, _097786_, _097787_);
  xor g_107818_(out[252], out[828], _097788_);
  or g_107819_(_097777_, _097788_, _097789_);
  xor g_107820_(out[247], out[823], _097790_);
  or g_107821_(_097772_, _097790_, _097791_);
  or g_107822_(_097789_, _097791_, _097792_);
  or g_107823_(_097778_, _097780_, _097793_);
  or g_107824_(_097773_, _097793_, _097794_);
  or g_107825_(_097792_, _097794_, _097795_);
  or g_107826_(_097776_, _097795_, _097796_);
  or g_107827_(_097787_, _097796_, _097797_);
  xor g_107828_(out[231], out[823], _097798_);
  and g_107829_(_098228_, out[827], _097799_);
  xor g_107830_(out[238], out[830], _097800_);
  xor g_107831_(out[232], out[824], _097801_);
  xor g_107832_(out[225], out[817], _097802_);
  xor g_107833_(out[237], out[829], _097803_);
  xor g_107834_(out[233], out[825], _097804_);
  xor g_107835_(out[228], out[820], _097805_);
  xor g_107836_(out[226], out[818], _097806_);
  and g_107837_(out[235], _049730_, _097807_);
  xor g_107838_(out[227], out[819], _097808_);
  xor g_107839_(out[230], out[822], _097809_);
  xor g_107840_(out[239], out[831], _097810_);
  xor g_107841_(out[234], out[826], _097811_);
  xor g_107842_(out[229], out[821], _097812_);
  xor g_107843_(out[224], out[816], _097813_);
  or g_107844_(_097800_, _097805_, _097814_);
  or g_107845_(_097801_, _097803_, _097815_);
  or g_107846_(_097806_, _097811_, _097816_);
  or g_107847_(_097815_, _097816_, _097817_);
  or g_107848_(_097804_, _097808_, _097818_);
  or g_107849_(_097812_, _097813_, _097819_);
  or g_107850_(_097818_, _097819_, _097820_);
  or g_107851_(_097817_, _097820_, _097821_);
  xor g_107852_(out[236], out[828], _097822_);
  or g_107853_(_097799_, _097822_, _097823_);
  or g_107854_(_097798_, _097809_, _097824_);
  or g_107855_(_097823_, _097824_, _097825_);
  or g_107856_(_097802_, _097807_, _097826_);
  or g_107857_(_097810_, _097826_, _097827_);
  or g_107858_(_097825_, _097827_, _097828_);
  or g_107859_(_097821_, _097828_, _097829_);
  or g_107860_(_097814_, _097829_, _097830_);
  xor g_107861_(out[209], out[817], _097831_);
  and g_107862_(out[219], _049730_, _097832_);
  xor g_107863_(out[217], out[825], _097833_);
  xor g_107864_(out[208], out[816], _097834_);
  xor g_107865_(out[222], out[830], _097835_);
  xor g_107866_(out[212], out[820], _097836_);
  or g_107867_(_097835_, _097836_, _097837_);
  xor g_107868_(out[221], out[829], _097838_);
  xor g_107869_(out[211], out[819], _097839_);
  and g_107870_(_098217_, out[827], _097840_);
  xor g_107871_(out[214], out[822], _097841_);
  xor g_107872_(out[218], out[826], _097842_);
  xor g_107873_(out[213], out[821], _097843_);
  xor g_107874_(out[223], out[831], _097844_);
  xor g_107875_(out[216], out[824], _097845_);
  or g_107876_(_097838_, _097845_, _097846_);
  xor g_107877_(out[210], out[818], _097847_);
  or g_107878_(_097842_, _097847_, _097848_);
  or g_107879_(_097846_, _097848_, _097849_);
  or g_107880_(_097833_, _097839_, _097850_);
  or g_107881_(_097843_, _097850_, _097851_);
  or g_107882_(_097849_, _097851_, _097852_);
  or g_107883_(_097837_, _097852_, _097853_);
  xor g_107884_(out[220], out[828], _097854_);
  or g_107885_(_097840_, _097854_, _097855_);
  xor g_107886_(out[215], out[823], _097856_);
  or g_107887_(_097841_, _097856_, _097857_);
  or g_107888_(_097855_, _097857_, _097858_);
  or g_107889_(_097831_, _097832_, _097859_);
  or g_107890_(_097844_, _097859_, _097860_);
  or g_107891_(_097858_, _097860_, _097861_);
  or g_107892_(_097834_, _097861_, _097862_);
  or g_107893_(_097853_, _097862_, _097863_);
  xor g_107894_(out[199], out[823], _097864_);
  and g_107895_(_098206_, out[827], _097865_);
  xor g_107896_(out[206], out[830], _097866_);
  xor g_107897_(out[200], out[824], _097867_);
  xor g_107898_(out[193], out[817], _097868_);
  xor g_107899_(out[205], out[829], _097869_);
  xor g_107900_(out[201], out[825], _097870_);
  xor g_107901_(out[196], out[820], _097871_);
  xor g_107902_(out[194], out[818], _097872_);
  and g_107903_(out[203], _049730_, _097873_);
  xor g_107904_(out[195], out[819], _097874_);
  xor g_107905_(out[198], out[822], _097875_);
  xor g_107906_(out[207], out[831], _097876_);
  xor g_107907_(out[202], out[826], _097877_);
  xor g_107908_(out[197], out[821], _097878_);
  xor g_107909_(out[192], out[816], _097879_);
  or g_107910_(_097866_, _097871_, _097880_);
  or g_107911_(_097867_, _097869_, _097881_);
  or g_107912_(_097872_, _097877_, _097882_);
  or g_107913_(_097881_, _097882_, _097883_);
  or g_107914_(_097870_, _097874_, _097884_);
  or g_107915_(_097878_, _097879_, _097885_);
  or g_107916_(_097884_, _097885_, _097886_);
  or g_107917_(_097883_, _097886_, _097887_);
  xor g_107918_(out[204], out[828], _097888_);
  or g_107919_(_097865_, _097888_, _097889_);
  or g_107920_(_097864_, _097875_, _097890_);
  or g_107921_(_097889_, _097890_, _097891_);
  or g_107922_(_097868_, _097873_, _097892_);
  or g_107923_(_097876_, _097892_, _097893_);
  or g_107924_(_097891_, _097893_, _097894_);
  or g_107925_(_097887_, _097894_, _097895_);
  or g_107926_(_097880_, _097895_, _097896_);
  not g_107927_(_097896_, _097897_);
  xor g_107928_(out[177], out[817], _097898_);
  and g_107929_(out[187], _049730_, _097899_);
  xor g_107930_(out[190], out[830], _097900_);
  xor g_107931_(out[179], out[819], _097901_);
  xor g_107932_(out[180], out[820], _097902_);
  xor g_107933_(out[178], out[818], _097903_);
  xor g_107934_(out[185], out[825], _097904_);
  xor g_107935_(out[176], out[816], _097905_);
  and g_107936_(_098195_, out[827], _097906_);
  xor g_107937_(out[182], out[822], _097907_);
  xor g_107938_(out[186], out[826], _097908_);
  xor g_107939_(out[181], out[821], _097909_);
  xor g_107940_(out[191], out[831], _097910_);
  xor g_107941_(out[189], out[829], _097911_);
  xor g_107942_(out[184], out[824], _097912_);
  or g_107943_(_097900_, _097902_, _097913_);
  or g_107944_(_097911_, _097912_, _097914_);
  or g_107945_(_097903_, _097908_, _097915_);
  or g_107946_(_097914_, _097915_, _097916_);
  or g_107947_(_097901_, _097904_, _097917_);
  or g_107948_(_097905_, _097909_, _097918_);
  or g_107949_(_097917_, _097918_, _097919_);
  or g_107950_(_097916_, _097919_, _097920_);
  xor g_107951_(out[188], out[828], _097921_);
  or g_107952_(_097906_, _097921_, _097922_);
  xor g_107953_(out[183], out[823], _097923_);
  or g_107954_(_097907_, _097923_, _097924_);
  or g_107955_(_097922_, _097924_, _097925_);
  or g_107956_(_097898_, _097899_, _097926_);
  or g_107957_(_097910_, _097926_, _097927_);
  or g_107958_(_097925_, _097927_, _097928_);
  or g_107959_(_097920_, _097928_, _097929_);
  or g_107960_(_097913_, _097929_, _097930_);
  xor g_107961_(out[167], out[823], _097931_);
  and g_107962_(_098184_, out[827], _097932_);
  xor g_107963_(out[174], out[830], _097933_);
  xor g_107964_(out[168], out[824], _097934_);
  xor g_107965_(out[161], out[817], _097935_);
  xor g_107966_(out[173], out[829], _097936_);
  xor g_107967_(out[169], out[825], _097937_);
  xor g_107968_(out[164], out[820], _097938_);
  xor g_107969_(out[162], out[818], _097939_);
  and g_107970_(out[171], _049730_, _097940_);
  xor g_107971_(out[163], out[819], _097941_);
  xor g_107972_(out[166], out[822], _097942_);
  xor g_107973_(out[175], out[831], _097943_);
  xor g_107974_(out[170], out[826], _097944_);
  xor g_107975_(out[165], out[821], _097945_);
  xor g_107976_(out[160], out[816], _097946_);
  or g_107977_(_097933_, _097938_, _097947_);
  or g_107978_(_097934_, _097936_, _097948_);
  or g_107979_(_097939_, _097944_, _097949_);
  or g_107980_(_097948_, _097949_, _097950_);
  or g_107981_(_097937_, _097941_, _097951_);
  or g_107982_(_097945_, _097946_, _097952_);
  or g_107983_(_097951_, _097952_, _097953_);
  or g_107984_(_097950_, _097953_, _097954_);
  xor g_107985_(out[172], out[828], _097955_);
  or g_107986_(_097932_, _097955_, _097956_);
  or g_107987_(_097931_, _097942_, _097957_);
  or g_107988_(_097956_, _097957_, _097958_);
  or g_107989_(_097935_, _097940_, _097959_);
  or g_107990_(_097943_, _097959_, _097960_);
  or g_107991_(_097958_, _097960_, _097961_);
  or g_107992_(_097954_, _097961_, _097962_);
  or g_107993_(_097947_, _097962_, _097963_);
  and g_107994_(_098173_, out[827], _097965_);
  and g_107995_(out[155], _049730_, _097966_);
  xor g_107996_(out[154], out[826], _097967_);
  xor g_107997_(out[159], out[831], _097968_);
  xor g_107998_(out[158], out[830], _097969_);
  xor g_107999_(out[144], out[816], _097970_);
  xor g_108000_(out[146], out[818], _097971_);
  xor g_108001_(out[147], out[819], _097972_);
  xor g_108002_(out[153], out[825], _097973_);
  xor g_108003_(out[145], out[817], _097974_);
  xor g_108004_(out[149], out[821], _097976_);
  xor g_108005_(out[150], out[822], _097977_);
  xor g_108006_(out[148], out[820], _097978_);
  xor g_108007_(out[157], out[829], _097979_);
  xor g_108008_(out[152], out[824], _097980_);
  or g_108009_(_097979_, _097980_, _097981_);
  or g_108010_(_097967_, _097971_, _097982_);
  or g_108011_(_097981_, _097982_, _097983_);
  or g_108012_(_097972_, _097973_, _097984_);
  or g_108013_(_097976_, _097984_, _097985_);
  or g_108014_(_097983_, _097985_, _097987_);
  or g_108015_(_097969_, _097978_, _097988_);
  or g_108016_(_097987_, _097988_, _097989_);
  xor g_108017_(out[156], out[828], _097990_);
  or g_108018_(_097965_, _097990_, _097991_);
  xor g_108019_(out[151], out[823], _097992_);
  or g_108020_(_097977_, _097992_, _097993_);
  or g_108021_(_097991_, _097993_, _097994_);
  or g_108022_(_097966_, _097974_, _097995_);
  or g_108023_(_097968_, _097995_, _097996_);
  or g_108024_(_097994_, _097996_, _097998_);
  or g_108025_(_097970_, _097998_, _097999_);
  or g_108026_(_097989_, _097999_, _098000_);
  not g_108027_(_098000_, _098001_);
  xor g_108028_(out[135], out[823], _098002_);
  and g_108029_(_098162_, out[827], _098003_);
  xor g_108030_(out[142], out[830], _098004_);
  xor g_108031_(out[136], out[824], _098005_);
  xor g_108032_(out[129], out[817], _098006_);
  xor g_108033_(out[141], out[829], _098007_);
  xor g_108034_(out[137], out[825], _098009_);
  xor g_108035_(out[132], out[820], _098010_);
  xor g_108036_(out[130], out[818], _098011_);
  and g_108037_(out[139], _049730_, _098012_);
  xor g_108038_(out[131], out[819], _098013_);
  xor g_108039_(out[134], out[822], _098014_);
  xor g_108040_(out[143], out[831], _098015_);
  xor g_108041_(out[138], out[826], _098016_);
  xor g_108042_(out[133], out[821], _098017_);
  xor g_108043_(out[128], out[816], _098018_);
  or g_108044_(_098004_, _098010_, _098020_);
  or g_108045_(_098005_, _098007_, _098021_);
  or g_108046_(_098011_, _098016_, _098022_);
  or g_108047_(_098021_, _098022_, _098023_);
  or g_108048_(_098009_, _098013_, _098024_);
  or g_108049_(_098017_, _098018_, _098025_);
  or g_108050_(_098024_, _098025_, _098026_);
  or g_108051_(_098023_, _098026_, _098027_);
  xor g_108052_(out[140], out[828], _098028_);
  or g_108053_(_098003_, _098028_, _098029_);
  or g_108054_(_098002_, _098014_, _098031_);
  or g_108055_(_098029_, _098031_, _098032_);
  or g_108056_(_098006_, _098012_, _098033_);
  or g_108057_(_098015_, _098033_, _098034_);
  or g_108058_(_098032_, _098034_, _098035_);
  or g_108059_(_098027_, _098035_, _098036_);
  or g_108060_(_098020_, _098036_, _098037_);
  not g_108061_(_098037_, _098038_);
  xor g_108062_(out[113], out[817], _098039_);
  and g_108063_(out[123], _049730_, _098040_);
  xor g_108064_(out[121], out[825], _098042_);
  xor g_108065_(out[112], out[816], _098043_);
  xor g_108066_(out[126], out[830], _098044_);
  xor g_108067_(out[116], out[820], _098045_);
  or g_108068_(_098044_, _098045_, _098046_);
  xor g_108069_(out[125], out[829], _098047_);
  xor g_108070_(out[115], out[819], _098048_);
  and g_108071_(_098151_, out[827], _098049_);
  xor g_108072_(out[118], out[822], _098050_);
  xor g_108073_(out[122], out[826], _098051_);
  xor g_108074_(out[117], out[821], _098053_);
  xor g_108075_(out[127], out[831], _098054_);
  xor g_108076_(out[120], out[824], _098055_);
  or g_108077_(_098047_, _098055_, _098056_);
  xor g_108078_(out[114], out[818], _098057_);
  or g_108079_(_098051_, _098057_, _098058_);
  or g_108080_(_098056_, _098058_, _098059_);
  or g_108081_(_098042_, _098048_, _098060_);
  or g_108082_(_098053_, _098060_, _098061_);
  or g_108083_(_098059_, _098061_, _098062_);
  or g_108084_(_098046_, _098062_, _098064_);
  xor g_108085_(out[124], out[828], _098065_);
  or g_108086_(_098049_, _098065_, _098066_);
  xor g_108087_(out[119], out[823], _098067_);
  or g_108088_(_098050_, _098067_, _098068_);
  or g_108089_(_098066_, _098068_, _098069_);
  or g_108090_(_098039_, _098040_, _098070_);
  or g_108091_(_098054_, _098070_, _098071_);
  or g_108092_(_098069_, _098071_, _098072_);
  or g_108093_(_098043_, _098072_, _098073_);
  or g_108094_(_098064_, _098073_, _098075_);
  xor g_108095_(out[103], out[823], _098076_);
  and g_108096_(_098140_, out[827], _098077_);
  xor g_108097_(out[110], out[830], _098078_);
  xor g_108098_(out[104], out[824], _098079_);
  xor g_108099_(out[97], out[817], _098080_);
  xor g_108100_(out[109], out[829], _098081_);
  xor g_108101_(out[105], out[825], _098082_);
  xor g_108102_(out[100], out[820], _098083_);
  xor g_108103_(out[98], out[818], _098084_);
  and g_108104_(out[107], _049730_, _098086_);
  xor g_108105_(out[99], out[819], _098087_);
  xor g_108106_(out[102], out[822], _098088_);
  xor g_108107_(out[111], out[831], _098089_);
  xor g_108108_(out[106], out[826], _098090_);
  xor g_108109_(out[101], out[821], _098091_);
  xor g_108110_(out[96], out[816], _098092_);
  or g_108111_(_098078_, _098083_, _098093_);
  or g_108112_(_098079_, _098081_, _098094_);
  or g_108113_(_098084_, _098090_, _098095_);
  or g_108114_(_098094_, _098095_, _098097_);
  or g_108115_(_098082_, _098087_, _098098_);
  or g_108116_(_098091_, _098092_, _098099_);
  or g_108117_(_098098_, _098099_, _098100_);
  or g_108118_(_098097_, _098100_, _098101_);
  xor g_108119_(out[108], out[828], _098102_);
  or g_108120_(_098077_, _098102_, _098103_);
  or g_108121_(_098076_, _098088_, _098104_);
  or g_108122_(_098103_, _098104_, _098105_);
  or g_108123_(_098080_, _098086_, _098106_);
  or g_108124_(_098089_, _098106_, _098108_);
  or g_108125_(_098105_, _098108_, _098109_);
  or g_108126_(_098101_, _098109_, _098110_);
  or g_108127_(_098093_, _098110_, _098111_);
  xor g_108128_(out[84], out[820], _098112_);
  xor g_108129_(out[92], out[828], _098113_);
  and g_108130_(_098129_, out[827], _098114_);
  xor g_108131_(out[90], out[826], _098115_);
  xor g_108132_(out[86], out[822], _098116_);
  xor g_108133_(out[85], out[821], _098117_);
  xor g_108134_(out[83], out[819], _098119_);
  xor g_108135_(out[93], out[829], _098120_);
  xor g_108136_(out[94], out[830], _098121_);
  xor g_108137_(out[81], out[817], _098122_);
  xor g_108138_(out[82], out[818], _098123_);
  and g_108139_(out[91], _049730_, _098124_);
  xor g_108140_(out[80], out[816], _098125_);
  xor g_108141_(out[95], out[831], _098126_);
  xor g_108142_(out[88], out[824], _098127_);
  or g_108143_(_098120_, _098127_, _098128_);
  xor g_108144_(out[89], out[825], _098130_);
  or g_108145_(_098115_, _098123_, _098131_);
  or g_108146_(_098128_, _098131_, _098132_);
  or g_108147_(_098119_, _098130_, _098133_);
  or g_108148_(_098117_, _098133_, _098134_);
  or g_108149_(_098132_, _098134_, _098135_);
  or g_108150_(_098112_, _098121_, _098136_);
  or g_108151_(_098135_, _098136_, _098137_);
  or g_108152_(_098113_, _098114_, _098138_);
  xor g_108153_(out[87], out[823], _098139_);
  or g_108154_(_098116_, _098139_, _098141_);
  or g_108155_(_098138_, _098141_, _098142_);
  or g_108156_(_098122_, _098124_, _098143_);
  or g_108157_(_098126_, _098143_, _098144_);
  or g_108158_(_098142_, _098144_, _098145_);
  or g_108159_(_098125_, _098145_, _098146_);
  or g_108160_(_098137_, _098146_, _098147_);
  not g_108161_(_098147_, _098148_);
  xor g_108162_(out[71], out[823], _098149_);
  and g_108163_(_098118_, out[827], _098150_);
  xor g_108164_(out[78], out[830], _098152_);
  xor g_108165_(out[72], out[824], _098153_);
  xor g_108166_(out[65], out[817], _098154_);
  xor g_108167_(out[77], out[829], _098155_);
  xor g_108168_(out[73], out[825], _098156_);
  xor g_108169_(out[68], out[820], _098157_);
  xor g_108170_(out[66], out[818], _098158_);
  and g_108171_(out[75], _049730_, _098159_);
  xor g_108172_(out[67], out[819], _098160_);
  xor g_108173_(out[70], out[822], _098161_);
  xor g_108174_(out[79], out[831], _098163_);
  xor g_108175_(out[74], out[826], _098164_);
  xor g_108176_(out[69], out[821], _098165_);
  xor g_108177_(out[64], out[816], _098166_);
  or g_108178_(_098152_, _098157_, _098167_);
  or g_108179_(_098153_, _098155_, _098168_);
  or g_108180_(_098158_, _098164_, _098169_);
  or g_108181_(_098168_, _098169_, _098170_);
  or g_108182_(_098156_, _098160_, _098171_);
  or g_108183_(_098165_, _098166_, _098172_);
  or g_108184_(_098171_, _098172_, _098174_);
  or g_108185_(_098170_, _098174_, _098175_);
  xor g_108186_(out[76], out[828], _098176_);
  or g_108187_(_098150_, _098176_, _098177_);
  or g_108188_(_098149_, _098161_, _098178_);
  or g_108189_(_098177_, _098178_, _098179_);
  or g_108190_(_098154_, _098159_, _098180_);
  or g_108191_(_098163_, _098180_, _098181_);
  or g_108192_(_098179_, _098181_, _098182_);
  or g_108193_(_098175_, _098182_, _098183_);
  or g_108194_(_098167_, _098183_, _098185_);
  not g_108195_(_098185_, _098186_);
  xor g_108196_(out[49], out[817], _098187_);
  and g_108197_(out[59], _049730_, _098188_);
  xor g_108198_(out[62], out[830], _098189_);
  xor g_108199_(out[51], out[819], _098190_);
  xor g_108200_(out[52], out[820], _098191_);
  xor g_108201_(out[50], out[818], _098192_);
  xor g_108202_(out[57], out[825], _098193_);
  xor g_108203_(out[48], out[816], _098194_);
  and g_108204_(_098107_, out[827], _098196_);
  xor g_108205_(out[54], out[822], _098197_);
  xor g_108206_(out[58], out[826], _098198_);
  xor g_108207_(out[53], out[821], _098199_);
  xor g_108208_(out[63], out[831], _098200_);
  xor g_108209_(out[61], out[829], _098201_);
  xor g_108210_(out[56], out[824], _098202_);
  or g_108211_(_098189_, _098191_, _098203_);
  or g_108212_(_098201_, _098202_, _098204_);
  or g_108213_(_098192_, _098198_, _098205_);
  or g_108214_(_098204_, _098205_, _098207_);
  or g_108215_(_098190_, _098193_, _098208_);
  or g_108216_(_098194_, _098199_, _098209_);
  or g_108217_(_098208_, _098209_, _098210_);
  or g_108218_(_098207_, _098210_, _098211_);
  xor g_108219_(out[60], out[828], _098212_);
  or g_108220_(_098196_, _098212_, _098213_);
  xor g_108221_(out[55], out[823], _098214_);
  or g_108222_(_098197_, _098214_, _098215_);
  or g_108223_(_098213_, _098215_, _098216_);
  or g_108224_(_098187_, _098188_, _098218_);
  or g_108225_(_098200_, _098218_, _098219_);
  or g_108226_(_098216_, _098219_, _098220_);
  or g_108227_(_098211_, _098220_, _098221_);
  or g_108228_(_098203_, _098221_, _098222_);
  not g_108229_(_098222_, _098223_);
  xor g_108230_(out[39], out[823], _098224_);
  and g_108231_(_098096_, out[827], _098225_);
  xor g_108232_(out[46], out[830], _098226_);
  xor g_108233_(out[40], out[824], _098227_);
  xor g_108234_(out[33], out[817], _098229_);
  xor g_108235_(out[45], out[829], _098230_);
  xor g_108236_(out[41], out[825], _098231_);
  xor g_108237_(out[36], out[820], _098232_);
  xor g_108238_(out[34], out[818], _098233_);
  and g_108239_(out[43], _049730_, _098234_);
  xor g_108240_(out[35], out[819], _098235_);
  xor g_108241_(out[38], out[822], _098236_);
  xor g_108242_(out[47], out[831], _098237_);
  xor g_108243_(out[42], out[826], _098238_);
  xor g_108244_(out[37], out[821], _098240_);
  xor g_108245_(out[32], out[816], _098241_);
  or g_108246_(_098226_, _098232_, _098242_);
  or g_108247_(_098227_, _098230_, _098243_);
  or g_108248_(_098233_, _098238_, _098244_);
  or g_108249_(_098243_, _098244_, _098245_);
  or g_108250_(_098231_, _098235_, _098246_);
  or g_108251_(_098240_, _098241_, _098247_);
  or g_108252_(_098246_, _098247_, _098248_);
  or g_108253_(_098245_, _098248_, _098249_);
  xor g_108254_(out[44], out[828], _098251_);
  or g_108255_(_098225_, _098251_, _098252_);
  or g_108256_(_098224_, _098236_, _098253_);
  or g_108257_(_098252_, _098253_, _098254_);
  or g_108258_(_098229_, _098234_, _098255_);
  or g_108259_(_098237_, _098255_, _098256_);
  or g_108260_(_098254_, _098256_, _098257_);
  or g_108261_(_098249_, _098257_, _098258_);
  or g_108262_(_098242_, _098258_, _098259_);
  xor g_108263_(out[17], out[817], _098260_);
  and g_108264_(_098063_, out[827], _098262_);
  and g_108265_(out[27], _049730_, _098263_);
  xor g_108266_(out[30], out[830], _098264_);
  xor g_108267_(out[19], out[819], _098265_);
  xor g_108268_(out[20], out[820], _098266_);
  xor g_108269_(out[18], out[818], _098267_);
  xor g_108270_(out[25], out[825], _098268_);
  xor g_108271_(out[16], out[816], _098269_);
  xor g_108272_(out[28], out[828], _098270_);
  xor g_108273_(out[22], out[822], _098271_);
  xor g_108274_(out[26], out[826], _098273_);
  xor g_108275_(out[21], out[821], _098274_);
  xor g_108276_(out[31], out[831], _098275_);
  xor g_108277_(out[29], out[829], _098276_);
  xor g_108278_(out[24], out[824], _098277_);
  or g_108279_(_098264_, _098266_, _098278_);
  or g_108280_(_098276_, _098277_, _098279_);
  or g_108281_(_098267_, _098273_, _098280_);
  or g_108282_(_098279_, _098280_, _098281_);
  or g_108283_(_098265_, _098268_, _098282_);
  or g_108284_(_098269_, _098274_, _098284_);
  or g_108285_(_098282_, _098284_, _098285_);
  or g_108286_(_098281_, _098285_, _098286_);
  or g_108287_(_098262_, _098270_, _098287_);
  xor g_108288_(out[23], out[823], _098288_);
  or g_108289_(_098271_, _098288_, _098289_);
  or g_108290_(_098287_, _098289_, _098290_);
  or g_108291_(_098260_, _098263_, _098291_);
  or g_108292_(_098275_, _098291_, _098292_);
  or g_108293_(_098290_, _098292_, _098293_);
  or g_108294_(_098286_, _098293_, _049390_);
  or g_108295_(_098278_, _049390_, _049391_);
  not g_108296_(_049391_, _049392_);
  xor g_108297_(out[1], out[817], _049393_);
  and g_108298_(out[11], _049730_, _049394_);
  xor g_108299_(out[9], out[825], _049395_);
  xor g_108300_(out[0], out[816], _049396_);
  xor g_108301_(out[14], out[830], _049397_);
  xor g_108302_(out[4], out[820], _049398_);
  or g_108303_(_049397_, _049398_, _049399_);
  xor g_108304_(out[13], out[829], _049401_);
  xor g_108305_(out[3], out[819], _049402_);
  and g_108306_(_098041_, out[827], _049403_);
  xor g_108307_(out[6], out[822], _049404_);
  xor g_108308_(out[10], out[826], _049405_);
  xor g_108309_(out[5], out[821], _049406_);
  xor g_108310_(out[15], out[831], _049407_);
  xor g_108311_(out[8], out[824], _049408_);
  or g_108312_(_049401_, _049408_, _049409_);
  xor g_108313_(out[2], out[818], _049410_);
  or g_108314_(_049405_, _049410_, _049412_);
  or g_108315_(_049409_, _049412_, _049413_);
  or g_108316_(_049395_, _049402_, _049414_);
  or g_108317_(_049406_, _049414_, _049415_);
  or g_108318_(_049413_, _049415_, _049416_);
  or g_108319_(_049399_, _049416_, _049417_);
  xor g_108320_(out[12], out[828], _049418_);
  or g_108321_(_049403_, _049418_, _049419_);
  xor g_108322_(out[7], out[823], _049420_);
  or g_108323_(_049404_, _049420_, _049421_);
  or g_108324_(_049419_, _049421_, _049423_);
  or g_108325_(_049393_, _049394_, _049424_);
  or g_108326_(_049407_, _049424_, _049425_);
  or g_108327_(_049423_, _049425_, _049426_);
  or g_108328_(_049396_, _049426_, _049427_);
  or g_108329_(_049417_, _049427_, _049428_);
  xor g_108330_(out[471], out[807], _049429_);
  and g_108331_(_049499_, out[811], _049430_);
  xor g_108332_(out[478], out[814], _049431_);
  xor g_108333_(out[472], out[808], _049432_);
  xor g_108334_(out[465], out[801], _049434_);
  xor g_108335_(out[477], out[813], _049435_);
  xor g_108336_(out[473], out[809], _049436_);
  xor g_108337_(out[468], out[804], _049437_);
  xor g_108338_(out[466], out[802], _049438_);
  and g_108339_(out[475], _049719_, _049439_);
  xor g_108340_(out[467], out[803], _049440_);
  xor g_108341_(out[470], out[806], _049441_);
  xor g_108342_(out[479], out[815], _049442_);
  xor g_108343_(out[474], out[810], _049443_);
  xor g_108344_(out[469], out[805], _049445_);
  xor g_108345_(out[464], out[800], _049446_);
  or g_108346_(_049431_, _049437_, _049447_);
  or g_108347_(_049432_, _049435_, _049448_);
  or g_108348_(_049438_, _049443_, _049449_);
  or g_108349_(_049448_, _049449_, _049450_);
  or g_108350_(_049436_, _049440_, _049451_);
  or g_108351_(_049445_, _049446_, _049452_);
  or g_108352_(_049451_, _049452_, _049453_);
  or g_108353_(_049450_, _049453_, _049454_);
  xor g_108354_(out[476], out[812], _049456_);
  or g_108355_(_049430_, _049456_, _049457_);
  or g_108356_(_049429_, _049441_, _049458_);
  or g_108357_(_049457_, _049458_, _049459_);
  or g_108358_(_049434_, _049439_, _049460_);
  or g_108359_(_049442_, _049460_, _049461_);
  or g_108360_(_049459_, _049461_, _049462_);
  or g_108361_(_049454_, _049462_, _049463_);
  or g_108362_(_049447_, _049463_, _049464_);
  xor g_108363_(out[458], out[810], _049465_);
  xor g_108364_(out[450], out[802], _049467_);
  xor g_108365_(out[449], out[801], _049468_);
  and g_108366_(_049477_, out[811], _049469_);
  and g_108367_(out[459], _049719_, _049470_);
  xor g_108368_(out[461], out[813], _049471_);
  xor g_108369_(out[451], out[803], _049472_);
  xor g_108370_(out[462], out[814], _049473_);
  xor g_108371_(out[460], out[812], _049474_);
  xor g_108372_(out[456], out[808], _049475_);
  xor g_108373_(out[463], out[815], _049476_);
  xor g_108374_(out[453], out[805], _049478_);
  xor g_108375_(out[454], out[806], _049479_);
  xor g_108376_(out[448], out[800], _049480_);
  xor g_108377_(out[452], out[804], _049481_);
  or g_108378_(_049471_, _049475_, _049482_);
  xor g_108379_(out[457], out[809], _049483_);
  or g_108380_(_049465_, _049467_, _049484_);
  or g_108381_(_049482_, _049484_, _049485_);
  or g_108382_(_049472_, _049483_, _049486_);
  or g_108383_(_049478_, _049486_, _049487_);
  or g_108384_(_049485_, _049487_, _049489_);
  or g_108385_(_049473_, _049481_, _049490_);
  or g_108386_(_049489_, _049490_, _049491_);
  or g_108387_(_049469_, _049474_, _049492_);
  xor g_108388_(out[455], out[807], _049493_);
  or g_108389_(_049479_, _049493_, _049494_);
  or g_108390_(_049492_, _049494_, _049495_);
  or g_108391_(_049468_, _049470_, _049496_);
  or g_108392_(_049476_, _049496_, _049497_);
  or g_108393_(_049495_, _049497_, _049498_);
  or g_108394_(_049480_, _049498_, _049500_);
  or g_108395_(_049491_, _049500_, _049501_);
  not g_108396_(_049501_, _049502_);
  xor g_108397_(out[439], out[807], _049503_);
  and g_108398_(_049466_, out[811], _049504_);
  xor g_108399_(out[446], out[814], _049505_);
  xor g_108400_(out[440], out[808], _049506_);
  xor g_108401_(out[433], out[801], _049507_);
  xor g_108402_(out[445], out[813], _049508_);
  xor g_108403_(out[441], out[809], _049509_);
  xor g_108404_(out[436], out[804], _049511_);
  xor g_108405_(out[434], out[802], _049512_);
  and g_108406_(out[443], _049719_, _049513_);
  xor g_108407_(out[435], out[803], _049514_);
  xor g_108408_(out[438], out[806], _049515_);
  xor g_108409_(out[447], out[815], _049516_);
  xor g_108410_(out[442], out[810], _049517_);
  xor g_108411_(out[437], out[805], _049518_);
  xor g_108412_(out[432], out[800], _049519_);
  or g_108413_(_049505_, _049511_, _049520_);
  or g_108414_(_049506_, _049508_, _049522_);
  or g_108415_(_049512_, _049517_, _049523_);
  or g_108416_(_049522_, _049523_, _049524_);
  or g_108417_(_049509_, _049514_, _049525_);
  or g_108418_(_049518_, _049519_, _049526_);
  or g_108419_(_049525_, _049526_, _049527_);
  or g_108420_(_049524_, _049527_, _049528_);
  xor g_108421_(out[444], out[812], _049529_);
  or g_108422_(_049504_, _049529_, _049530_);
  or g_108423_(_049503_, _049515_, _049531_);
  or g_108424_(_049530_, _049531_, _049533_);
  or g_108425_(_049507_, _049513_, _049534_);
  or g_108426_(_049516_, _049534_, _049535_);
  or g_108427_(_049533_, _049535_, _049536_);
  or g_108428_(_049528_, _049536_, _049537_);
  or g_108429_(_049520_, _049537_, _049538_);
  xor g_108430_(out[417], out[801], _049539_);
  and g_108431_(_049455_, out[811], _049540_);
  and g_108432_(out[427], _049719_, _049541_);
  xor g_108433_(out[424], out[808], _049542_);
  xor g_108434_(out[426], out[810], _049544_);
  xor g_108435_(out[418], out[802], _049545_);
  xor g_108436_(out[420], out[804], _049546_);
  xor g_108437_(out[429], out[813], _049547_);
  xor g_108438_(out[425], out[809], _049548_);
  xor g_108439_(out[419], out[803], _049549_);
  xor g_108440_(out[421], out[805], _049550_);
  xor g_108441_(out[430], out[814], _049551_);
  xor g_108442_(out[416], out[800], _049552_);
  xor g_108443_(out[431], out[815], _049553_);
  or g_108444_(_049542_, _049547_, _049555_);
  xor g_108445_(out[422], out[806], _049556_);
  or g_108446_(_049544_, _049545_, _049557_);
  or g_108447_(_049555_, _049557_, _049558_);
  or g_108448_(_049548_, _049549_, _049559_);
  or g_108449_(_049550_, _049559_, _049560_);
  or g_108450_(_049558_, _049560_, _049561_);
  or g_108451_(_049546_, _049551_, _049562_);
  or g_108452_(_049561_, _049562_, _049563_);
  xor g_108453_(out[428], out[812], _049564_);
  or g_108454_(_049540_, _049564_, _049566_);
  xor g_108455_(out[423], out[807], _049567_);
  or g_108456_(_049556_, _049567_, _049568_);
  or g_108457_(_049566_, _049568_, _049569_);
  or g_108458_(_049539_, _049541_, _049570_);
  or g_108459_(_049553_, _049570_, _049571_);
  or g_108460_(_049569_, _049571_, _049572_);
  or g_108461_(_049552_, _049572_, _049573_);
  or g_108462_(_049563_, _049573_, _049574_);
  xor g_108463_(out[407], out[807], _049575_);
  and g_108464_(_049444_, out[811], _049577_);
  xor g_108465_(out[414], out[814], _049578_);
  xor g_108466_(out[408], out[808], _049579_);
  xor g_108467_(out[401], out[801], _049580_);
  xor g_108468_(out[413], out[813], _049581_);
  xor g_108469_(out[409], out[809], _049582_);
  xor g_108470_(out[404], out[804], _049583_);
  xor g_108471_(out[402], out[802], _049584_);
  and g_108472_(out[411], _049719_, _049585_);
  xor g_108473_(out[403], out[803], _049586_);
  xor g_108474_(out[406], out[806], _049588_);
  xor g_108475_(out[415], out[815], _049589_);
  xor g_108476_(out[410], out[810], _049590_);
  xor g_108477_(out[405], out[805], _049591_);
  xor g_108478_(out[400], out[800], _049592_);
  or g_108479_(_049578_, _049583_, _049593_);
  or g_108480_(_049579_, _049581_, _049594_);
  or g_108481_(_049584_, _049590_, _049595_);
  or g_108482_(_049594_, _049595_, _049596_);
  or g_108483_(_049582_, _049586_, _049597_);
  or g_108484_(_049591_, _049592_, _049599_);
  or g_108485_(_049597_, _049599_, _049600_);
  or g_108486_(_049596_, _049600_, _049601_);
  xor g_108487_(out[412], out[812], _049602_);
  or g_108488_(_049577_, _049602_, _049603_);
  or g_108489_(_049575_, _049588_, _049604_);
  or g_108490_(_049603_, _049604_, _049605_);
  or g_108491_(_049580_, _049585_, _049606_);
  or g_108492_(_049589_, _049606_, _049607_);
  or g_108493_(_049605_, _049607_, _049608_);
  or g_108494_(_049601_, _049608_, _049610_);
  or g_108495_(_049593_, _049610_, _049611_);
  xor g_108496_(out[385], out[801], _049612_);
  and g_108497_(out[395], _049719_, _049613_);
  xor g_108498_(out[393], out[809], _049614_);
  xor g_108499_(out[384], out[800], _049615_);
  xor g_108500_(out[398], out[814], _049616_);
  xor g_108501_(out[388], out[804], _049617_);
  or g_108502_(_049616_, _049617_, _049618_);
  xor g_108503_(out[397], out[813], _049619_);
  xor g_108504_(out[387], out[803], _049621_);
  and g_108505_(_049433_, out[811], _049622_);
  xor g_108506_(out[390], out[806], _049623_);
  xor g_108507_(out[394], out[810], _049624_);
  xor g_108508_(out[389], out[805], _049625_);
  xor g_108509_(out[399], out[815], _049626_);
  xor g_108510_(out[392], out[808], _049627_);
  or g_108511_(_049619_, _049627_, _049628_);
  xor g_108512_(out[386], out[802], _049629_);
  or g_108513_(_049624_, _049629_, _049630_);
  or g_108514_(_049628_, _049630_, _049632_);
  or g_108515_(_049614_, _049621_, _049633_);
  or g_108516_(_049625_, _049633_, _049634_);
  or g_108517_(_049632_, _049634_, _049635_);
  or g_108518_(_049618_, _049635_, _049636_);
  xor g_108519_(out[396], out[812], _049637_);
  or g_108520_(_049622_, _049637_, _049638_);
  xor g_108521_(out[391], out[807], _049639_);
  or g_108522_(_049623_, _049639_, _049640_);
  or g_108523_(_049638_, _049640_, _049641_);
  or g_108524_(_049612_, _049613_, _049643_);
  or g_108525_(_049626_, _049643_, _049644_);
  or g_108526_(_049641_, _049644_, _049645_);
  or g_108527_(_049615_, _049645_, _049646_);
  or g_108528_(_049636_, _049646_, _049647_);
  not g_108529_(_049647_, _049648_);
  xor g_108530_(out[375], out[807], _049649_);
  and g_108531_(_049422_, out[811], _049650_);
  xor g_108532_(out[382], out[814], _049651_);
  xor g_108533_(out[376], out[808], _049652_);
  xor g_108534_(out[369], out[801], _049654_);
  xor g_108535_(out[381], out[813], _049655_);
  xor g_108536_(out[377], out[809], _049656_);
  xor g_108537_(out[372], out[804], _049657_);
  xor g_108538_(out[370], out[802], _049658_);
  and g_108539_(out[379], _049719_, _049659_);
  xor g_108540_(out[371], out[803], _049660_);
  xor g_108541_(out[374], out[806], _049661_);
  xor g_108542_(out[383], out[815], _049662_);
  xor g_108543_(out[378], out[810], _049663_);
  xor g_108544_(out[373], out[805], _049665_);
  xor g_108545_(out[368], out[800], _049666_);
  or g_108546_(_049651_, _049657_, _049667_);
  or g_108547_(_049652_, _049655_, _049668_);
  or g_108548_(_049658_, _049663_, _049669_);
  or g_108549_(_049668_, _049669_, _049670_);
  or g_108550_(_049656_, _049660_, _049671_);
  or g_108551_(_049665_, _049666_, _049672_);
  or g_108552_(_049671_, _049672_, _049673_);
  or g_108553_(_049670_, _049673_, _049674_);
  xor g_108554_(out[380], out[812], _049676_);
  or g_108555_(_049650_, _049676_, _049677_);
  or g_108556_(_049649_, _049661_, _049678_);
  or g_108557_(_049677_, _049678_, _049679_);
  or g_108558_(_049654_, _049659_, _049680_);
  or g_108559_(_049662_, _049680_, _049681_);
  or g_108560_(_049679_, _049681_, _049682_);
  or g_108561_(_049674_, _049682_, _049683_);
  or g_108562_(_049667_, _049683_, _049684_);
  not g_108563_(_049684_, _049685_);
  xor g_108564_(out[355], out[803], _049687_);
  xor g_108565_(out[356], out[804], _049688_);
  xor g_108566_(out[366], out[814], _049689_);
  xor g_108567_(out[354], out[802], _049690_);
  xor g_108568_(out[357], out[805], _049691_);
  xor g_108569_(out[361], out[809], _049692_);
  xor g_108570_(out[360], out[808], _049693_);
  xor g_108571_(out[367], out[815], _049694_);
  xor g_108572_(out[362], out[810], _049695_);
  xor g_108573_(out[358], out[806], _049696_);
  xor g_108574_(out[352], out[800], _049698_);
  and g_108575_(_049411_, out[811], _049699_);
  and g_108576_(out[363], _049719_, _049700_);
  xor g_108577_(out[365], out[813], _049701_);
  or g_108578_(_049693_, _049701_, _049702_);
  xor g_108579_(out[353], out[801], _049703_);
  or g_108580_(_049690_, _049695_, _049704_);
  or g_108581_(_049702_, _049704_, _049705_);
  or g_108582_(_049687_, _049692_, _049706_);
  or g_108583_(_049691_, _049706_, _049707_);
  or g_108584_(_049705_, _049707_, _049709_);
  or g_108585_(_049688_, _049689_, _049710_);
  or g_108586_(_049709_, _049710_, _049711_);
  xor g_108587_(out[364], out[812], _049712_);
  or g_108588_(_049699_, _049712_, _049713_);
  xor g_108589_(out[359], out[807], _049714_);
  or g_108590_(_049696_, _049714_, _049715_);
  or g_108591_(_049713_, _049715_, _049716_);
  or g_108592_(_049700_, _049703_, _049717_);
  or g_108593_(_049694_, _049717_, _049718_);
  or g_108594_(_049716_, _049718_, _049720_);
  or g_108595_(_049698_, _049720_, _049721_);
  or g_108596_(_049711_, _049721_, _049722_);
  xor g_108597_(out[343], out[807], _049723_);
  and g_108598_(_049400_, out[811], _049724_);
  xor g_108599_(out[350], out[814], _049725_);
  xor g_108600_(out[344], out[808], _049726_);
  xor g_108601_(out[337], out[801], _049727_);
  xor g_108602_(out[349], out[813], _049728_);
  xor g_108603_(out[345], out[809], _049729_);
  xor g_108604_(out[340], out[804], _049731_);
  xor g_108605_(out[338], out[802], _049732_);
  and g_108606_(out[347], _049719_, _049733_);
  xor g_108607_(out[339], out[803], _049734_);
  xor g_108608_(out[342], out[806], _049735_);
  xor g_108609_(out[351], out[815], _049736_);
  xor g_108610_(out[346], out[810], _049737_);
  xor g_108611_(out[341], out[805], _049738_);
  xor g_108612_(out[336], out[800], _049739_);
  or g_108613_(_049725_, _049731_, _049740_);
  or g_108614_(_049726_, _049728_, _049742_);
  or g_108615_(_049732_, _049737_, _049743_);
  or g_108616_(_049742_, _049743_, _049744_);
  or g_108617_(_049729_, _049734_, _049745_);
  or g_108618_(_049738_, _049739_, _049746_);
  or g_108619_(_049745_, _049746_, _049747_);
  or g_108620_(_049744_, _049747_, _049748_);
  xor g_108621_(out[348], out[812], _049749_);
  or g_108622_(_049724_, _049749_, _049750_);
  or g_108623_(_049723_, _049735_, _049751_);
  or g_108624_(_049750_, _049751_, _049753_);
  or g_108625_(_049727_, _049733_, _049754_);
  or g_108626_(_049736_, _049754_, _049755_);
  or g_108627_(_049753_, _049755_, _049756_);
  or g_108628_(_049748_, _049756_, _049757_);
  or g_108629_(_049740_, _049757_, _049758_);
  not g_108630_(_049758_, _049759_);
  xor g_108631_(out[321], out[801], _049760_);
  and g_108632_(out[331], _049719_, _049761_);
  xor g_108633_(out[329], out[809], _049762_);
  xor g_108634_(out[320], out[800], _049764_);
  xor g_108635_(out[334], out[814], _049765_);
  xor g_108636_(out[324], out[804], _049766_);
  or g_108637_(_049765_, _049766_, _049767_);
  xor g_108638_(out[333], out[813], _049768_);
  xor g_108639_(out[323], out[803], _049769_);
  and g_108640_(_098294_, out[811], _049770_);
  xor g_108641_(out[326], out[806], _049771_);
  xor g_108642_(out[330], out[810], _049772_);
  xor g_108643_(out[325], out[805], _049773_);
  xor g_108644_(out[335], out[815], _049775_);
  xor g_108645_(out[328], out[808], _049776_);
  or g_108646_(_049768_, _049776_, _049777_);
  xor g_108647_(out[322], out[802], _049778_);
  or g_108648_(_049772_, _049778_, _049779_);
  or g_108649_(_049777_, _049779_, _049780_);
  or g_108650_(_049762_, _049769_, _049781_);
  or g_108651_(_049773_, _049781_, _049782_);
  or g_108652_(_049780_, _049782_, _049783_);
  or g_108653_(_049767_, _049783_, _049784_);
  xor g_108654_(out[332], out[812], _049786_);
  or g_108655_(_049770_, _049786_, _049787_);
  xor g_108656_(out[327], out[807], _049788_);
  or g_108657_(_049771_, _049788_, _049789_);
  or g_108658_(_049787_, _049789_, _049790_);
  or g_108659_(_049760_, _049761_, _049791_);
  or g_108660_(_049775_, _049791_, _049792_);
  or g_108661_(_049790_, _049792_, _049793_);
  or g_108662_(_049764_, _049793_, _049794_);
  or g_108663_(_049784_, _049794_, _049795_);
  xor g_108664_(out[311], out[807], _049797_);
  and g_108665_(_098283_, out[811], _049798_);
  xor g_108666_(out[318], out[814], _049799_);
  xor g_108667_(out[312], out[808], _049800_);
  xor g_108668_(out[305], out[801], _049801_);
  xor g_108669_(out[317], out[813], _049802_);
  xor g_108670_(out[313], out[809], _049803_);
  xor g_108671_(out[308], out[804], _049804_);
  xor g_108672_(out[306], out[802], _049805_);
  and g_108673_(out[315], _049719_, _049806_);
  xor g_108674_(out[307], out[803], _049808_);
  xor g_108675_(out[310], out[806], _049809_);
  xor g_108676_(out[319], out[815], _049810_);
  xor g_108677_(out[314], out[810], _049811_);
  xor g_108678_(out[309], out[805], _049812_);
  xor g_108679_(out[304], out[800], _049813_);
  or g_108680_(_049799_, _049804_, _049814_);
  or g_108681_(_049800_, _049802_, _049815_);
  or g_108682_(_049805_, _049811_, _049816_);
  or g_108683_(_049815_, _049816_, _049817_);
  or g_108684_(_049803_, _049808_, _049819_);
  or g_108685_(_049812_, _049813_, _049820_);
  or g_108686_(_049819_, _049820_, _049821_);
  or g_108687_(_049817_, _049821_, _049822_);
  xor g_108688_(out[316], out[812], _049823_);
  or g_108689_(_049798_, _049823_, _049824_);
  or g_108690_(_049797_, _049809_, _049825_);
  or g_108691_(_049824_, _049825_, _049826_);
  or g_108692_(_049801_, _049806_, _049827_);
  or g_108693_(_049810_, _049827_, _049828_);
  or g_108694_(_049826_, _049828_, _049830_);
  or g_108695_(_049822_, _049830_, _049831_);
  or g_108696_(_049814_, _049831_, _049832_);
  and g_108697_(out[299], _049719_, _049833_);
  xor g_108698_(out[292], out[804], _049834_);
  xor g_108699_(out[290], out[802], _049835_);
  xor g_108700_(out[297], out[809], _049836_);
  xor g_108701_(out[288], out[800], _049837_);
  xor g_108702_(out[291], out[803], _049838_);
  and g_108703_(_098272_, out[811], _049839_);
  xor g_108704_(out[298], out[810], _049841_);
  xor g_108705_(out[303], out[815], _049842_);
  xor g_108706_(out[294], out[806], _049843_);
  xor g_108707_(out[293], out[805], _049844_);
  xor g_108708_(out[301], out[813], _049845_);
  xor g_108709_(out[302], out[814], _049846_);
  xor g_108710_(out[296], out[808], _049847_);
  xor g_108711_(out[289], out[801], _049848_);
  or g_108712_(_049834_, _049846_, _049849_);
  or g_108713_(_049845_, _049847_, _049850_);
  or g_108714_(_049835_, _049841_, _049852_);
  or g_108715_(_049850_, _049852_, _049853_);
  or g_108716_(_049836_, _049838_, _049854_);
  or g_108717_(_049837_, _049844_, _049855_);
  or g_108718_(_049854_, _049855_, _049856_);
  or g_108719_(_049853_, _049856_, _049857_);
  xor g_108720_(out[300], out[812], _049858_);
  or g_108721_(_049839_, _049858_, _049859_);
  xor g_108722_(out[295], out[807], _049860_);
  or g_108723_(_049843_, _049860_, _049861_);
  or g_108724_(_049859_, _049861_, _049863_);
  or g_108725_(_049833_, _049848_, _049864_);
  or g_108726_(_049842_, _049864_, _049865_);
  or g_108727_(_049863_, _049865_, _049866_);
  or g_108728_(_049857_, _049866_, _049867_);
  or g_108729_(_049849_, _049867_, _049868_);
  xor g_108730_(out[279], out[807], _049869_);
  and g_108731_(_098261_, out[811], _049870_);
  xor g_108732_(out[286], out[814], _049871_);
  xor g_108733_(out[280], out[808], _049872_);
  xor g_108734_(out[273], out[801], _049874_);
  xor g_108735_(out[285], out[813], _049875_);
  xor g_108736_(out[281], out[809], _049876_);
  xor g_108737_(out[276], out[804], _049877_);
  xor g_108738_(out[274], out[802], _049878_);
  and g_108739_(out[283], _049719_, _049879_);
  xor g_108740_(out[275], out[803], _049880_);
  xor g_108741_(out[278], out[806], _049881_);
  xor g_108742_(out[287], out[815], _049882_);
  xor g_108743_(out[282], out[810], _049883_);
  xor g_108744_(out[277], out[805], _049885_);
  xor g_108745_(out[272], out[800], _049886_);
  or g_108746_(_049871_, _049877_, _049887_);
  or g_108747_(_049872_, _049875_, _049888_);
  or g_108748_(_049878_, _049883_, _049889_);
  or g_108749_(_049888_, _049889_, _049890_);
  or g_108750_(_049876_, _049880_, _049891_);
  or g_108751_(_049885_, _049886_, _049892_);
  or g_108752_(_049891_, _049892_, _049893_);
  or g_108753_(_049890_, _049893_, _049894_);
  xor g_108754_(out[284], out[812], _049896_);
  or g_108755_(_049870_, _049896_, _049897_);
  or g_108756_(_049869_, _049881_, _049898_);
  or g_108757_(_049897_, _049898_, _049899_);
  or g_108758_(_049874_, _049879_, _049900_);
  or g_108759_(_049882_, _049900_, _049901_);
  or g_108760_(_049899_, _049901_, _049902_);
  or g_108761_(_049894_, _049902_, _049903_);
  or g_108762_(_049887_, _049903_, _049904_);
  xor g_108763_(out[266], out[810], _049905_);
  xor g_108764_(out[264], out[808], _049907_);
  xor g_108765_(out[257], out[801], _049908_);
  and g_108766_(_098250_, out[811], _049909_);
  and g_108767_(out[267], _049719_, _049910_);
  xor g_108768_(out[258], out[802], _049911_);
  xor g_108769_(out[261], out[805], _049912_);
  xor g_108770_(out[265], out[809], _049913_);
  xor g_108771_(out[268], out[812], _049914_);
  xor g_108772_(out[269], out[813], _049915_);
  xor g_108773_(out[271], out[815], _049916_);
  xor g_108774_(out[260], out[804], _049918_);
  xor g_108775_(out[262], out[806], _049919_);
  xor g_108776_(out[259], out[803], _049920_);
  xor g_108777_(out[256], out[800], _049921_);
  xor g_108778_(out[270], out[814], _049922_);
  or g_108779_(_049918_, _049922_, _049923_);
  or g_108780_(_049907_, _049915_, _049924_);
  or g_108781_(_049905_, _049911_, _049925_);
  or g_108782_(_049924_, _049925_, _049926_);
  or g_108783_(_049913_, _049920_, _049927_);
  or g_108784_(_049912_, _049921_, _049929_);
  or g_108785_(_049927_, _049929_, _049930_);
  or g_108786_(_049926_, _049930_, _049931_);
  or g_108787_(_049909_, _049914_, _049932_);
  xor g_108788_(out[263], out[807], _049933_);
  or g_108789_(_049919_, _049933_, _049934_);
  or g_108790_(_049932_, _049934_, _049935_);
  or g_108791_(_049908_, _049910_, _049936_);
  or g_108792_(_049916_, _049936_, _049937_);
  or g_108793_(_049935_, _049937_, _049938_);
  or g_108794_(_049931_, _049938_, _049940_);
  or g_108795_(_049923_, _049940_, _049941_);
  xor g_108796_(out[247], out[807], _049942_);
  and g_108797_(_098239_, out[811], _049943_);
  xor g_108798_(out[254], out[814], _049944_);
  xor g_108799_(out[248], out[808], _049945_);
  xor g_108800_(out[241], out[801], _049946_);
  xor g_108801_(out[253], out[813], _049947_);
  xor g_108802_(out[249], out[809], _049948_);
  xor g_108803_(out[244], out[804], _049949_);
  xor g_108804_(out[242], out[802], _049951_);
  and g_108805_(out[251], _049719_, _049952_);
  xor g_108806_(out[243], out[803], _049953_);
  xor g_108807_(out[246], out[806], _049954_);
  xor g_108808_(out[255], out[815], _049955_);
  xor g_108809_(out[250], out[810], _049956_);
  xor g_108810_(out[245], out[805], _049957_);
  xor g_108811_(out[240], out[800], _049958_);
  or g_108812_(_049944_, _049949_, _049959_);
  or g_108813_(_049945_, _049947_, _049960_);
  or g_108814_(_049951_, _049956_, _049962_);
  or g_108815_(_049960_, _049962_, _049963_);
  or g_108816_(_049948_, _049953_, _049964_);
  or g_108817_(_049957_, _049958_, _049965_);
  or g_108818_(_049964_, _049965_, _049966_);
  or g_108819_(_049963_, _049966_, _049967_);
  xor g_108820_(out[252], out[812], _049968_);
  or g_108821_(_049943_, _049968_, _049969_);
  or g_108822_(_049942_, _049954_, _049970_);
  or g_108823_(_049969_, _049970_, _049971_);
  or g_108824_(_049946_, _049952_, _049973_);
  or g_108825_(_049955_, _049973_, _049974_);
  or g_108826_(_049971_, _049974_, _049975_);
  or g_108827_(_049967_, _049975_, _049976_);
  or g_108828_(_049959_, _049976_, _049977_);
  xor g_108829_(out[225], out[801], _049978_);
  and g_108830_(out[235], _049719_, _049979_);
  xor g_108831_(out[233], out[809], _049980_);
  xor g_108832_(out[224], out[800], _049981_);
  xor g_108833_(out[238], out[814], _049982_);
  xor g_108834_(out[228], out[804], _049984_);
  or g_108835_(_049982_, _049984_, _049985_);
  xor g_108836_(out[237], out[813], _049986_);
  xor g_108837_(out[227], out[803], _049987_);
  and g_108838_(_098228_, out[811], _049988_);
  xor g_108839_(out[230], out[806], _049989_);
  xor g_108840_(out[234], out[810], _049990_);
  xor g_108841_(out[229], out[805], _049991_);
  xor g_108842_(out[239], out[815], _049992_);
  xor g_108843_(out[232], out[808], _049993_);
  or g_108844_(_049986_, _049993_, _049995_);
  xor g_108845_(out[226], out[802], _049996_);
  or g_108846_(_049990_, _049996_, _049997_);
  or g_108847_(_049995_, _049997_, _049998_);
  or g_108848_(_049980_, _049987_, _049999_);
  or g_108849_(_049991_, _049999_, _050000_);
  or g_108850_(_049998_, _050000_, _050001_);
  or g_108851_(_049985_, _050001_, _050002_);
  xor g_108852_(out[236], out[812], _050003_);
  or g_108853_(_049988_, _050003_, _050004_);
  xor g_108854_(out[231], out[807], _050006_);
  or g_108855_(_049989_, _050006_, _050007_);
  or g_108856_(_050004_, _050007_, _050008_);
  or g_108857_(_049978_, _049979_, _050009_);
  or g_108858_(_049992_, _050009_, _050010_);
  or g_108859_(_050008_, _050010_, _050011_);
  or g_108860_(_049981_, _050011_, _050012_);
  or g_108861_(_050002_, _050012_, _050013_);
  xor g_108862_(out[215], out[807], _050014_);
  and g_108863_(_098217_, out[811], _050015_);
  xor g_108864_(out[222], out[814], _050017_);
  xor g_108865_(out[216], out[808], _050018_);
  xor g_108866_(out[209], out[801], _050019_);
  xor g_108867_(out[221], out[813], _050020_);
  xor g_108868_(out[217], out[809], _050021_);
  xor g_108869_(out[212], out[804], _050022_);
  xor g_108870_(out[210], out[802], _050023_);
  and g_108871_(out[219], _049719_, _050024_);
  xor g_108872_(out[211], out[803], _050025_);
  xor g_108873_(out[214], out[806], _050026_);
  xor g_108874_(out[223], out[815], _050028_);
  xor g_108875_(out[218], out[810], _050029_);
  xor g_108876_(out[213], out[805], _050030_);
  xor g_108877_(out[208], out[800], _050031_);
  or g_108878_(_050017_, _050022_, _050032_);
  or g_108879_(_050018_, _050020_, _050033_);
  or g_108880_(_050023_, _050029_, _050034_);
  or g_108881_(_050033_, _050034_, _050035_);
  or g_108882_(_050021_, _050025_, _050036_);
  or g_108883_(_050030_, _050031_, _050037_);
  or g_108884_(_050036_, _050037_, _050039_);
  or g_108885_(_050035_, _050039_, _050040_);
  xor g_108886_(out[220], out[812], _050041_);
  or g_108887_(_050015_, _050041_, _050042_);
  or g_108888_(_050014_, _050026_, _050043_);
  or g_108889_(_050042_, _050043_, _050044_);
  or g_108890_(_050019_, _050024_, _050045_);
  or g_108891_(_050028_, _050045_, _050046_);
  or g_108892_(_050044_, _050046_, _050047_);
  or g_108893_(_050040_, _050047_, _050048_);
  or g_108894_(_050032_, _050048_, _050050_);
  xor g_108895_(out[204], out[812], _050051_);
  and g_108896_(_098206_, out[811], _050052_);
  xor g_108897_(out[200], out[808], _050053_);
  xor g_108898_(out[198], out[806], _050054_);
  xor g_108899_(out[205], out[813], _050055_);
  xor g_108900_(out[206], out[814], _050056_);
  xor g_108901_(out[194], out[802], _050057_);
  xor g_108902_(out[201], out[809], _050058_);
  xor g_108903_(out[197], out[805], _050059_);
  xor g_108904_(out[193], out[801], _050061_);
  and g_108905_(out[203], _049719_, _050062_);
  or g_108906_(_050053_, _050055_, _050063_);
  xor g_108907_(out[207], out[815], _050064_);
  xor g_108908_(out[202], out[810], _050065_);
  xor g_108909_(out[196], out[804], _050066_);
  xor g_108910_(out[195], out[803], _050067_);
  xor g_108911_(out[192], out[800], _050068_);
  or g_108912_(_050057_, _050065_, _050069_);
  or g_108913_(_050063_, _050069_, _050070_);
  or g_108914_(_050058_, _050067_, _050072_);
  or g_108915_(_050059_, _050072_, _050073_);
  or g_108916_(_050070_, _050073_, _050074_);
  or g_108917_(_050056_, _050066_, _050075_);
  or g_108918_(_050074_, _050075_, _050076_);
  or g_108919_(_050051_, _050052_, _050077_);
  xor g_108920_(out[199], out[807], _050078_);
  or g_108921_(_050054_, _050078_, _050079_);
  or g_108922_(_050077_, _050079_, _050080_);
  or g_108923_(_050061_, _050062_, _050081_);
  or g_108924_(_050064_, _050081_, _050083_);
  or g_108925_(_050080_, _050083_, _050084_);
  or g_108926_(_050068_, _050084_, _050085_);
  or g_108927_(_050076_, _050085_, _050086_);
  xor g_108928_(out[183], out[807], _050087_);
  and g_108929_(_098195_, out[811], _050088_);
  xor g_108930_(out[190], out[814], _050089_);
  xor g_108931_(out[184], out[808], _050090_);
  xor g_108932_(out[177], out[801], _050091_);
  xor g_108933_(out[189], out[813], _050092_);
  xor g_108934_(out[185], out[809], _050094_);
  xor g_108935_(out[180], out[804], _050095_);
  xor g_108936_(out[178], out[802], _050096_);
  and g_108937_(out[187], _049719_, _050097_);
  xor g_108938_(out[179], out[803], _050098_);
  xor g_108939_(out[182], out[806], _050099_);
  xor g_108940_(out[191], out[815], _050100_);
  xor g_108941_(out[186], out[810], _050101_);
  xor g_108942_(out[181], out[805], _050102_);
  xor g_108943_(out[176], out[800], _050103_);
  or g_108944_(_050089_, _050095_, _050105_);
  or g_108945_(_050090_, _050092_, _050106_);
  or g_108946_(_050096_, _050101_, _050107_);
  or g_108947_(_050106_, _050107_, _050108_);
  or g_108948_(_050094_, _050098_, _050109_);
  or g_108949_(_050102_, _050103_, _050110_);
  or g_108950_(_050109_, _050110_, _050111_);
  or g_108951_(_050108_, _050111_, _050112_);
  xor g_108952_(out[188], out[812], _050113_);
  or g_108953_(_050088_, _050113_, _050114_);
  or g_108954_(_050087_, _050099_, _050116_);
  or g_108955_(_050114_, _050116_, _050117_);
  or g_108956_(_050091_, _050097_, _050118_);
  or g_108957_(_050100_, _050118_, _050119_);
  or g_108958_(_050117_, _050119_, _050120_);
  or g_108959_(_050112_, _050120_, _050121_);
  or g_108960_(_050105_, _050121_, _050122_);
  xor g_108961_(out[161], out[801], _050123_);
  and g_108962_(out[171], _049719_, _050124_);
  xor g_108963_(out[169], out[809], _050125_);
  xor g_108964_(out[160], out[800], _050127_);
  xor g_108965_(out[174], out[814], _050128_);
  xor g_108966_(out[164], out[804], _050129_);
  or g_108967_(_050128_, _050129_, _050130_);
  xor g_108968_(out[173], out[813], _050131_);
  xor g_108969_(out[163], out[803], _050132_);
  and g_108970_(_098184_, out[811], _050133_);
  xor g_108971_(out[166], out[806], _050134_);
  xor g_108972_(out[170], out[810], _050135_);
  xor g_108973_(out[165], out[805], _050136_);
  xor g_108974_(out[175], out[815], _050138_);
  xor g_108975_(out[168], out[808], _050139_);
  or g_108976_(_050131_, _050139_, _050140_);
  xor g_108977_(out[162], out[802], _050141_);
  or g_108978_(_050135_, _050141_, _050142_);
  or g_108979_(_050140_, _050142_, _050143_);
  or g_108980_(_050125_, _050132_, _050144_);
  or g_108981_(_050136_, _050144_, _050145_);
  or g_108982_(_050143_, _050145_, _050146_);
  or g_108983_(_050130_, _050146_, _050147_);
  xor g_108984_(out[172], out[812], _050149_);
  or g_108985_(_050133_, _050149_, _050150_);
  xor g_108986_(out[167], out[807], _050151_);
  or g_108987_(_050134_, _050151_, _050152_);
  or g_108988_(_050150_, _050152_, _050153_);
  or g_108989_(_050123_, _050124_, _050154_);
  or g_108990_(_050138_, _050154_, _050155_);
  or g_108991_(_050153_, _050155_, _050156_);
  or g_108992_(_050127_, _050156_, _050157_);
  or g_108993_(_050147_, _050157_, _050158_);
  xor g_108994_(out[151], out[807], _050160_);
  and g_108995_(_098173_, out[811], _050161_);
  xor g_108996_(out[158], out[814], _050162_);
  xor g_108997_(out[152], out[808], _050163_);
  xor g_108998_(out[145], out[801], _050164_);
  xor g_108999_(out[157], out[813], _050165_);
  xor g_109000_(out[153], out[809], _050166_);
  xor g_109001_(out[148], out[804], _050167_);
  xor g_109002_(out[146], out[802], _050168_);
  and g_109003_(out[155], _049719_, _050169_);
  xor g_109004_(out[147], out[803], _050171_);
  xor g_109005_(out[150], out[806], _050172_);
  xor g_109006_(out[159], out[815], _050173_);
  xor g_109007_(out[154], out[810], _050174_);
  xor g_109008_(out[149], out[805], _050175_);
  xor g_109009_(out[144], out[800], _050176_);
  or g_109010_(_050162_, _050167_, _050177_);
  or g_109011_(_050163_, _050165_, _050178_);
  or g_109012_(_050168_, _050174_, _050179_);
  or g_109013_(_050178_, _050179_, _050180_);
  or g_109014_(_050166_, _050171_, _050182_);
  or g_109015_(_050175_, _050176_, _050183_);
  or g_109016_(_050182_, _050183_, _050184_);
  or g_109017_(_050180_, _050184_, _050185_);
  xor g_109018_(out[156], out[812], _050186_);
  or g_109019_(_050161_, _050186_, _050187_);
  or g_109020_(_050160_, _050172_, _050188_);
  or g_109021_(_050187_, _050188_, _050189_);
  or g_109022_(_050164_, _050169_, _050190_);
  or g_109023_(_050173_, _050190_, _050191_);
  or g_109024_(_050189_, _050191_, _050193_);
  or g_109025_(_050185_, _050193_, _050194_);
  or g_109026_(_050177_, _050194_, _050195_);
  xor g_109027_(out[129], out[801], _050196_);
  and g_109028_(out[139], _049719_, _050197_);
  xor g_109029_(out[137], out[809], _050198_);
  xor g_109030_(out[128], out[800], _050199_);
  xor g_109031_(out[142], out[814], _050200_);
  xor g_109032_(out[132], out[804], _050201_);
  or g_109033_(_050200_, _050201_, _050202_);
  xor g_109034_(out[141], out[813], _050204_);
  xor g_109035_(out[131], out[803], _050205_);
  and g_109036_(_098162_, out[811], _050206_);
  xor g_109037_(out[134], out[806], _050207_);
  xor g_109038_(out[138], out[810], _050208_);
  xor g_109039_(out[133], out[805], _050209_);
  xor g_109040_(out[143], out[815], _050210_);
  xor g_109041_(out[136], out[808], _050211_);
  or g_109042_(_050204_, _050211_, _050212_);
  xor g_109043_(out[130], out[802], _050213_);
  or g_109044_(_050208_, _050213_, _050215_);
  or g_109045_(_050212_, _050215_, _050216_);
  or g_109046_(_050198_, _050205_, _050217_);
  or g_109047_(_050209_, _050217_, _050218_);
  or g_109048_(_050216_, _050218_, _050219_);
  or g_109049_(_050202_, _050219_, _050220_);
  xor g_109050_(out[140], out[812], _050221_);
  or g_109051_(_050206_, _050221_, _050222_);
  xor g_109052_(out[135], out[807], _050223_);
  or g_109053_(_050207_, _050223_, _050224_);
  or g_109054_(_050222_, _050224_, _050226_);
  or g_109055_(_050196_, _050197_, _050227_);
  or g_109056_(_050210_, _050227_, _050228_);
  or g_109057_(_050226_, _050228_, _050229_);
  or g_109058_(_050199_, _050229_, _050230_);
  or g_109059_(_050220_, _050230_, _050231_);
  xor g_109060_(out[119], out[807], _050232_);
  and g_109061_(_098151_, out[811], _050233_);
  xor g_109062_(out[126], out[814], _050234_);
  xor g_109063_(out[120], out[808], _050235_);
  xor g_109064_(out[113], out[801], _050237_);
  xor g_109065_(out[125], out[813], _050238_);
  xor g_109066_(out[121], out[809], _050239_);
  xor g_109067_(out[116], out[804], _050240_);
  xor g_109068_(out[114], out[802], _050241_);
  and g_109069_(out[123], _049719_, _050242_);
  xor g_109070_(out[115], out[803], _050243_);
  xor g_109071_(out[118], out[806], _050244_);
  xor g_109072_(out[127], out[815], _050245_);
  xor g_109073_(out[122], out[810], _050246_);
  xor g_109074_(out[117], out[805], _050248_);
  xor g_109075_(out[112], out[800], _050249_);
  or g_109076_(_050234_, _050240_, _050250_);
  or g_109077_(_050235_, _050238_, _050251_);
  or g_109078_(_050241_, _050246_, _050252_);
  or g_109079_(_050251_, _050252_, _050253_);
  or g_109080_(_050239_, _050243_, _050254_);
  or g_109081_(_050248_, _050249_, _050255_);
  or g_109082_(_050254_, _050255_, _050256_);
  or g_109083_(_050253_, _050256_, _050257_);
  xor g_109084_(out[124], out[812], _050259_);
  or g_109085_(_050233_, _050259_, _050260_);
  or g_109086_(_050232_, _050244_, _050261_);
  or g_109087_(_050260_, _050261_, _050262_);
  or g_109088_(_050237_, _050242_, _050263_);
  or g_109089_(_050245_, _050263_, _050264_);
  or g_109090_(_050262_, _050264_, _050265_);
  or g_109091_(_050257_, _050265_, _050266_);
  or g_109092_(_050250_, _050266_, _050267_);
  xor g_109093_(out[108], out[812], _050268_);
  and g_109094_(_098140_, out[811], _050270_);
  xor g_109095_(out[104], out[808], _050271_);
  xor g_109096_(out[102], out[806], _050272_);
  xor g_109097_(out[109], out[813], _050273_);
  xor g_109098_(out[110], out[814], _050274_);
  xor g_109099_(out[98], out[802], _050275_);
  xor g_109100_(out[105], out[809], _050276_);
  xor g_109101_(out[101], out[805], _050277_);
  xor g_109102_(out[97], out[801], _050278_);
  and g_109103_(out[107], _049719_, _050279_);
  or g_109104_(_050271_, _050273_, _050281_);
  xor g_109105_(out[111], out[815], _050282_);
  xor g_109106_(out[106], out[810], _050283_);
  xor g_109107_(out[100], out[804], _050284_);
  xor g_109108_(out[99], out[803], _050285_);
  xor g_109109_(out[96], out[800], _050286_);
  or g_109110_(_050275_, _050283_, _050287_);
  or g_109111_(_050281_, _050287_, _050288_);
  or g_109112_(_050276_, _050285_, _050289_);
  or g_109113_(_050277_, _050289_, _050290_);
  or g_109114_(_050288_, _050290_, _050292_);
  or g_109115_(_050274_, _050284_, _050293_);
  or g_109116_(_050292_, _050293_, _050294_);
  or g_109117_(_050268_, _050270_, _050295_);
  xor g_109118_(out[103], out[807], _050296_);
  or g_109119_(_050272_, _050296_, _050297_);
  or g_109120_(_050295_, _050297_, _050298_);
  or g_109121_(_050278_, _050279_, _050299_);
  or g_109122_(_050282_, _050299_, _050300_);
  or g_109123_(_050298_, _050300_, _050301_);
  or g_109124_(_050286_, _050301_, _050303_);
  or g_109125_(_050294_, _050303_, _050304_);
  not g_109126_(_050304_, _050305_);
  xor g_109127_(out[87], out[807], _050306_);
  and g_109128_(_098129_, out[811], _050307_);
  xor g_109129_(out[94], out[814], _050308_);
  xor g_109130_(out[88], out[808], _050309_);
  xor g_109131_(out[81], out[801], _050310_);
  xor g_109132_(out[93], out[813], _050311_);
  xor g_109133_(out[89], out[809], _050312_);
  xor g_109134_(out[84], out[804], _050314_);
  xor g_109135_(out[82], out[802], _050315_);
  and g_109136_(out[91], _049719_, _050316_);
  xor g_109137_(out[83], out[803], _050317_);
  xor g_109138_(out[86], out[806], _050318_);
  xor g_109139_(out[95], out[815], _050319_);
  xor g_109140_(out[90], out[810], _050320_);
  xor g_109141_(out[85], out[805], _050321_);
  xor g_109142_(out[80], out[800], _050322_);
  or g_109143_(_050308_, _050314_, _050323_);
  or g_109144_(_050309_, _050311_, _050325_);
  or g_109145_(_050315_, _050320_, _050326_);
  or g_109146_(_050325_, _050326_, _050327_);
  or g_109147_(_050312_, _050317_, _050328_);
  or g_109148_(_050321_, _050322_, _050329_);
  or g_109149_(_050328_, _050329_, _050330_);
  or g_109150_(_050327_, _050330_, _050331_);
  xor g_109151_(out[92], out[812], _050332_);
  or g_109152_(_050307_, _050332_, _050333_);
  or g_109153_(_050306_, _050318_, _050334_);
  or g_109154_(_050333_, _050334_, _050336_);
  or g_109155_(_050310_, _050316_, _050337_);
  or g_109156_(_050319_, _050337_, _050338_);
  or g_109157_(_050336_, _050338_, _050339_);
  or g_109158_(_050331_, _050339_, _050340_);
  or g_109159_(_050323_, _050340_, _050341_);
  xor g_109160_(out[65], out[801], _050342_);
  and g_109161_(out[75], _049719_, _050343_);
  xor g_109162_(out[73], out[809], _050344_);
  xor g_109163_(out[64], out[800], _050345_);
  xor g_109164_(out[78], out[814], _050347_);
  xor g_109165_(out[68], out[804], _050348_);
  or g_109166_(_050347_, _050348_, _050349_);
  xor g_109167_(out[77], out[813], _050350_);
  xor g_109168_(out[67], out[803], _050351_);
  and g_109169_(_098118_, out[811], _050352_);
  xor g_109170_(out[70], out[806], _050353_);
  xor g_109171_(out[74], out[810], _050354_);
  xor g_109172_(out[69], out[805], _050355_);
  xor g_109173_(out[79], out[815], _050356_);
  xor g_109174_(out[72], out[808], _050358_);
  or g_109175_(_050350_, _050358_, _050359_);
  xor g_109176_(out[66], out[802], _050360_);
  or g_109177_(_050354_, _050360_, _050361_);
  or g_109178_(_050359_, _050361_, _050362_);
  or g_109179_(_050344_, _050351_, _050363_);
  or g_109180_(_050355_, _050363_, _050364_);
  or g_109181_(_050362_, _050364_, _050365_);
  or g_109182_(_050349_, _050365_, _050366_);
  xor g_109183_(out[76], out[812], _050367_);
  or g_109184_(_050352_, _050367_, _050369_);
  xor g_109185_(out[71], out[807], _050370_);
  or g_109186_(_050353_, _050370_, _050371_);
  or g_109187_(_050369_, _050371_, _050372_);
  or g_109188_(_050342_, _050343_, _050373_);
  or g_109189_(_050356_, _050373_, _050374_);
  or g_109190_(_050372_, _050374_, _050375_);
  or g_109191_(_050345_, _050375_, _050376_);
  or g_109192_(_050366_, _050376_, _050377_);
  xor g_109193_(out[55], out[807], _050378_);
  and g_109194_(_098107_, out[811], _050380_);
  xor g_109195_(out[62], out[814], _050381_);
  xor g_109196_(out[56], out[808], _050382_);
  xor g_109197_(out[49], out[801], _050383_);
  xor g_109198_(out[61], out[813], _050384_);
  xor g_109199_(out[57], out[809], _050385_);
  xor g_109200_(out[52], out[804], _050386_);
  xor g_109201_(out[50], out[802], _050387_);
  and g_109202_(out[59], _049719_, _050388_);
  xor g_109203_(out[51], out[803], _050389_);
  xor g_109204_(out[54], out[806], _050391_);
  xor g_109205_(out[63], out[815], _050392_);
  xor g_109206_(out[58], out[810], _050393_);
  xor g_109207_(out[53], out[805], _050394_);
  xor g_109208_(out[48], out[800], _050395_);
  or g_109209_(_050381_, _050386_, _050396_);
  or g_109210_(_050382_, _050384_, _050397_);
  or g_109211_(_050387_, _050393_, _050398_);
  or g_109212_(_050397_, _050398_, _050399_);
  or g_109213_(_050385_, _050389_, _050400_);
  or g_109214_(_050394_, _050395_, _050402_);
  or g_109215_(_050400_, _050402_, _050403_);
  or g_109216_(_050399_, _050403_, _050404_);
  xor g_109217_(out[60], out[812], _050405_);
  or g_109218_(_050380_, _050405_, _050406_);
  or g_109219_(_050378_, _050391_, _050407_);
  or g_109220_(_050406_, _050407_, _050408_);
  or g_109221_(_050383_, _050388_, _050409_);
  or g_109222_(_050392_, _050409_, _050410_);
  or g_109223_(_050408_, _050410_, _050411_);
  or g_109224_(_050404_, _050411_, _050413_);
  or g_109225_(_050396_, _050413_, _050414_);
  xor g_109226_(out[33], out[801], _050415_);
  and g_109227_(out[43], _049719_, _050416_);
  xor g_109228_(out[41], out[809], _050417_);
  xor g_109229_(out[32], out[800], _050418_);
  xor g_109230_(out[46], out[814], _050419_);
  xor g_109231_(out[36], out[804], _050420_);
  or g_109232_(_050419_, _050420_, _050421_);
  xor g_109233_(out[45], out[813], _050422_);
  xor g_109234_(out[35], out[803], _050424_);
  and g_109235_(_098096_, out[811], _050425_);
  xor g_109236_(out[38], out[806], _050426_);
  xor g_109237_(out[42], out[810], _050427_);
  xor g_109238_(out[37], out[805], _050428_);
  xor g_109239_(out[47], out[815], _050429_);
  xor g_109240_(out[40], out[808], _050430_);
  or g_109241_(_050422_, _050430_, _050431_);
  xor g_109242_(out[34], out[802], _050432_);
  or g_109243_(_050427_, _050432_, _050433_);
  or g_109244_(_050431_, _050433_, _050435_);
  or g_109245_(_050417_, _050424_, _050436_);
  or g_109246_(_050428_, _050436_, _050437_);
  or g_109247_(_050435_, _050437_, _050438_);
  or g_109248_(_050421_, _050438_, _050439_);
  xor g_109249_(out[44], out[812], _050440_);
  or g_109250_(_050425_, _050440_, _050441_);
  xor g_109251_(out[39], out[807], _050442_);
  or g_109252_(_050426_, _050442_, _050443_);
  or g_109253_(_050441_, _050443_, _050444_);
  or g_109254_(_050415_, _050416_, _050446_);
  or g_109255_(_050429_, _050446_, _050447_);
  or g_109256_(_050444_, _050447_, _050448_);
  or g_109257_(_050418_, _050448_, _050449_);
  or g_109258_(_050439_, _050449_, _050450_);
  xor g_109259_(out[23], out[807], _050451_);
  and g_109260_(_098063_, out[811], _050452_);
  xor g_109261_(out[30], out[814], _050453_);
  xor g_109262_(out[24], out[808], _050454_);
  xor g_109263_(out[17], out[801], _050455_);
  xor g_109264_(out[29], out[813], _050457_);
  xor g_109265_(out[25], out[809], _050458_);
  xor g_109266_(out[20], out[804], _050459_);
  xor g_109267_(out[18], out[802], _050460_);
  and g_109268_(out[27], _049719_, _050461_);
  xor g_109269_(out[19], out[803], _050462_);
  xor g_109270_(out[22], out[806], _050463_);
  xor g_109271_(out[31], out[815], _050464_);
  xor g_109272_(out[26], out[810], _050465_);
  xor g_109273_(out[21], out[805], _050466_);
  xor g_109274_(out[16], out[800], _050468_);
  or g_109275_(_050453_, _050459_, _050469_);
  or g_109276_(_050454_, _050457_, _050470_);
  or g_109277_(_050460_, _050465_, _050471_);
  or g_109278_(_050470_, _050471_, _050472_);
  or g_109279_(_050458_, _050462_, _050473_);
  or g_109280_(_050466_, _050468_, _050474_);
  or g_109281_(_050473_, _050474_, _050475_);
  or g_109282_(_050472_, _050475_, _050476_);
  xor g_109283_(out[28], out[812], _050477_);
  or g_109284_(_050452_, _050477_, _050479_);
  or g_109285_(_050451_, _050463_, _050480_);
  or g_109286_(_050479_, _050480_, _050481_);
  or g_109287_(_050455_, _050461_, _050482_);
  or g_109288_(_050464_, _050482_, _050483_);
  or g_109289_(_050481_, _050483_, _050484_);
  or g_109290_(_050476_, _050484_, _050485_);
  or g_109291_(_050469_, _050485_, _050486_);
  and g_109292_(out[11], _049719_, _050487_);
  xor g_109293_(out[4], out[804], _050488_);
  xor g_109294_(out[14], out[814], _050490_);
  or g_109295_(_050488_, _050490_, _050491_);
  xor g_109296_(out[13], out[813], _050492_);
  xor g_109297_(out[3], out[803], _050493_);
  xor g_109298_(out[0], out[800], _050494_);
  and g_109299_(_098041_, out[811], _050495_);
  xor g_109300_(out[10], out[810], _050496_);
  xor g_109301_(out[15], out[815], _050497_);
  xor g_109302_(out[6], out[806], _050498_);
  xor g_109303_(out[5], out[805], _050499_);
  xor g_109304_(out[8], out[808], _050501_);
  or g_109305_(_050492_, _050501_, _050502_);
  xor g_109306_(out[2], out[802], _050503_);
  xor g_109307_(out[9], out[809], _050504_);
  xor g_109308_(out[1], out[801], _050505_);
  or g_109309_(_050496_, _050503_, _050506_);
  or g_109310_(_050502_, _050506_, _050507_);
  or g_109311_(_050493_, _050504_, _050508_);
  or g_109312_(_050499_, _050508_, _050509_);
  or g_109313_(_050507_, _050509_, _050510_);
  or g_109314_(_050491_, _050510_, _050512_);
  xor g_109315_(out[12], out[812], _050513_);
  or g_109316_(_050495_, _050513_, _050514_);
  xor g_109317_(out[7], out[807], _050515_);
  or g_109318_(_050498_, _050515_, _050516_);
  or g_109319_(_050514_, _050516_, _050517_);
  or g_109320_(_050487_, _050505_, _050518_);
  or g_109321_(_050497_, _050518_, _050519_);
  or g_109322_(_050517_, _050519_, _050520_);
  or g_109323_(_050494_, _050520_, _050521_);
  or g_109324_(_050512_, _050521_, _050523_);
  and g_109325_(out[475], _049708_, _050524_);
  xor g_109326_(out[476], out[796], _050525_);
  and g_109327_(_049499_, out[795], _050526_);
  xor g_109328_(out[473], out[793], _050527_);
  xor g_109329_(out[468], out[788], _050528_);
  xor g_109330_(out[469], out[789], _050529_);
  xor g_109331_(out[465], out[785], _050530_);
  xor g_109332_(out[477], out[797], _050531_);
  xor g_109333_(out[474], out[794], _050532_);
  xor g_109334_(out[470], out[790], _050534_);
  xor g_109335_(out[472], out[792], _050535_);
  or g_109336_(_050531_, _050535_, _050536_);
  xor g_109337_(out[466], out[786], _050537_);
  xor g_109338_(out[479], out[799], _050538_);
  xor g_109339_(out[467], out[787], _050539_);
  xor g_109340_(out[478], out[798], _050540_);
  xor g_109341_(out[464], out[784], _050541_);
  or g_109342_(_050532_, _050537_, _050542_);
  or g_109343_(_050536_, _050542_, _050543_);
  or g_109344_(_050527_, _050539_, _050545_);
  or g_109345_(_050529_, _050545_, _050546_);
  or g_109346_(_050543_, _050546_, _050547_);
  or g_109347_(_050528_, _050540_, _050548_);
  or g_109348_(_050547_, _050548_, _050549_);
  or g_109349_(_050525_, _050526_, _050550_);
  xor g_109350_(out[471], out[791], _050551_);
  or g_109351_(_050534_, _050551_, _050552_);
  or g_109352_(_050550_, _050552_, _050553_);
  or g_109353_(_050524_, _050530_, _050554_);
  or g_109354_(_050538_, _050554_, _050556_);
  or g_109355_(_050553_, _050556_, _050557_);
  or g_109356_(_050541_, _050557_, _050558_);
  or g_109357_(_050549_, _050558_, _050559_);
  xor g_109358_(out[455], out[791], _050560_);
  and g_109359_(_049477_, out[795], _050561_);
  xor g_109360_(out[462], out[798], _050562_);
  xor g_109361_(out[456], out[792], _050563_);
  xor g_109362_(out[449], out[785], _050564_);
  xor g_109363_(out[461], out[797], _050565_);
  xor g_109364_(out[457], out[793], _050567_);
  xor g_109365_(out[452], out[788], _050568_);
  xor g_109366_(out[450], out[786], _050569_);
  and g_109367_(out[459], _049708_, _050570_);
  xor g_109368_(out[451], out[787], _050571_);
  xor g_109369_(out[454], out[790], _050572_);
  xor g_109370_(out[463], out[799], _050573_);
  xor g_109371_(out[458], out[794], _050574_);
  xor g_109372_(out[453], out[789], _050575_);
  xor g_109373_(out[448], out[784], _050576_);
  or g_109374_(_050562_, _050568_, _050578_);
  or g_109375_(_050563_, _050565_, _050579_);
  or g_109376_(_050569_, _050574_, _050580_);
  or g_109377_(_050579_, _050580_, _050581_);
  or g_109378_(_050567_, _050571_, _050582_);
  or g_109379_(_050575_, _050576_, _050583_);
  or g_109380_(_050582_, _050583_, _050584_);
  or g_109381_(_050581_, _050584_, _050585_);
  xor g_109382_(out[460], out[796], _050586_);
  or g_109383_(_050561_, _050586_, _050587_);
  or g_109384_(_050560_, _050572_, _050589_);
  or g_109385_(_050587_, _050589_, _050590_);
  or g_109386_(_050564_, _050570_, _050591_);
  or g_109387_(_050573_, _050591_, _050592_);
  or g_109388_(_050590_, _050592_, _050593_);
  or g_109389_(_050585_, _050593_, _050594_);
  or g_109390_(_050578_, _050594_, _050595_);
  xor g_109391_(out[433], out[785], _050596_);
  and g_109392_(out[443], _049708_, _050597_);
  xor g_109393_(out[441], out[793], _050598_);
  xor g_109394_(out[432], out[784], _050600_);
  xor g_109395_(out[446], out[798], _050601_);
  xor g_109396_(out[436], out[788], _050602_);
  or g_109397_(_050601_, _050602_, _050603_);
  xor g_109398_(out[445], out[797], _050604_);
  xor g_109399_(out[435], out[787], _050605_);
  and g_109400_(_049466_, out[795], _050606_);
  xor g_109401_(out[438], out[790], _050607_);
  xor g_109402_(out[442], out[794], _050608_);
  xor g_109403_(out[437], out[789], _050609_);
  xor g_109404_(out[447], out[799], _050611_);
  xor g_109405_(out[440], out[792], _050612_);
  or g_109406_(_050604_, _050612_, _050613_);
  xor g_109407_(out[434], out[786], _050614_);
  or g_109408_(_050608_, _050614_, _050615_);
  or g_109409_(_050613_, _050615_, _050616_);
  or g_109410_(_050598_, _050605_, _050617_);
  or g_109411_(_050609_, _050617_, _050618_);
  or g_109412_(_050616_, _050618_, _050619_);
  or g_109413_(_050603_, _050619_, _050620_);
  xor g_109414_(out[444], out[796], _050622_);
  or g_109415_(_050606_, _050622_, _050623_);
  xor g_109416_(out[439], out[791], _050624_);
  or g_109417_(_050607_, _050624_, _050625_);
  or g_109418_(_050623_, _050625_, _050626_);
  or g_109419_(_050596_, _050597_, _050627_);
  or g_109420_(_050611_, _050627_, _050628_);
  or g_109421_(_050626_, _050628_, _050629_);
  or g_109422_(_050600_, _050629_, _050630_);
  or g_109423_(_050620_, _050630_, _050631_);
  not g_109424_(_050631_, _050633_);
  xor g_109425_(out[423], out[791], _050634_);
  and g_109426_(_049455_, out[795], _050635_);
  xor g_109427_(out[430], out[798], _050636_);
  xor g_109428_(out[424], out[792], _050637_);
  xor g_109429_(out[417], out[785], _050638_);
  xor g_109430_(out[429], out[797], _050639_);
  xor g_109431_(out[425], out[793], _050640_);
  xor g_109432_(out[420], out[788], _050641_);
  xor g_109433_(out[418], out[786], _050642_);
  and g_109434_(out[427], _049708_, _050644_);
  xor g_109435_(out[419], out[787], _050645_);
  xor g_109436_(out[422], out[790], _050646_);
  xor g_109437_(out[431], out[799], _050647_);
  xor g_109438_(out[426], out[794], _050648_);
  xor g_109439_(out[421], out[789], _050649_);
  xor g_109440_(out[416], out[784], _050650_);
  or g_109441_(_050636_, _050641_, _050651_);
  or g_109442_(_050637_, _050639_, _050652_);
  or g_109443_(_050642_, _050648_, _050653_);
  or g_109444_(_050652_, _050653_, _050655_);
  or g_109445_(_050640_, _050645_, _050656_);
  or g_109446_(_050649_, _050650_, _050657_);
  or g_109447_(_050656_, _050657_, _050658_);
  or g_109448_(_050655_, _050658_, _050659_);
  xor g_109449_(out[428], out[796], _050660_);
  or g_109450_(_050635_, _050660_, _050661_);
  or g_109451_(_050634_, _050646_, _050662_);
  or g_109452_(_050661_, _050662_, _050663_);
  or g_109453_(_050638_, _050644_, _050664_);
  or g_109454_(_050647_, _050664_, _050666_);
  or g_109455_(_050663_, _050666_, _050667_);
  or g_109456_(_050659_, _050667_, _050668_);
  or g_109457_(_050651_, _050668_, _050669_);
  xor g_109458_(out[401], out[785], _050670_);
  and g_109459_(out[411], _049708_, _050671_);
  xor g_109460_(out[409], out[793], _050672_);
  xor g_109461_(out[400], out[784], _050673_);
  xor g_109462_(out[414], out[798], _050674_);
  xor g_109463_(out[404], out[788], _050675_);
  or g_109464_(_050674_, _050675_, _050677_);
  xor g_109465_(out[413], out[797], _050678_);
  xor g_109466_(out[403], out[787], _050679_);
  and g_109467_(_049444_, out[795], _050680_);
  xor g_109468_(out[406], out[790], _050681_);
  xor g_109469_(out[410], out[794], _050682_);
  xor g_109470_(out[405], out[789], _050683_);
  xor g_109471_(out[415], out[799], _050684_);
  xor g_109472_(out[408], out[792], _050685_);
  or g_109473_(_050678_, _050685_, _050686_);
  xor g_109474_(out[402], out[786], _050688_);
  or g_109475_(_050682_, _050688_, _050689_);
  or g_109476_(_050686_, _050689_, _050690_);
  or g_109477_(_050672_, _050679_, _050691_);
  or g_109478_(_050683_, _050691_, _050692_);
  or g_109479_(_050690_, _050692_, _050693_);
  or g_109480_(_050677_, _050693_, _050694_);
  xor g_109481_(out[412], out[796], _050695_);
  or g_109482_(_050680_, _050695_, _050696_);
  xor g_109483_(out[407], out[791], _050697_);
  or g_109484_(_050681_, _050697_, _050699_);
  or g_109485_(_050696_, _050699_, _050700_);
  or g_109486_(_050670_, _050671_, _050701_);
  or g_109487_(_050684_, _050701_, _050702_);
  or g_109488_(_050700_, _050702_, _050703_);
  or g_109489_(_050673_, _050703_, _050704_);
  or g_109490_(_050694_, _050704_, _050705_);
  xor g_109491_(out[391], out[791], _050706_);
  and g_109492_(_049433_, out[795], _050707_);
  xor g_109493_(out[398], out[798], _050708_);
  xor g_109494_(out[392], out[792], _050710_);
  xor g_109495_(out[385], out[785], _050711_);
  xor g_109496_(out[397], out[797], _050712_);
  xor g_109497_(out[393], out[793], _050713_);
  xor g_109498_(out[388], out[788], _050714_);
  xor g_109499_(out[386], out[786], _050715_);
  and g_109500_(out[395], _049708_, _050716_);
  xor g_109501_(out[387], out[787], _050717_);
  xor g_109502_(out[390], out[790], _050718_);
  xor g_109503_(out[399], out[799], _050719_);
  xor g_109504_(out[394], out[794], _050721_);
  xor g_109505_(out[389], out[789], _050722_);
  xor g_109506_(out[384], out[784], _050723_);
  or g_109507_(_050708_, _050714_, _050724_);
  or g_109508_(_050710_, _050712_, _050725_);
  or g_109509_(_050715_, _050721_, _050726_);
  or g_109510_(_050725_, _050726_, _050727_);
  or g_109511_(_050713_, _050717_, _050728_);
  or g_109512_(_050722_, _050723_, _050729_);
  or g_109513_(_050728_, _050729_, _050730_);
  or g_109514_(_050727_, _050730_, _050732_);
  xor g_109515_(out[396], out[796], _050733_);
  or g_109516_(_050707_, _050733_, _050734_);
  or g_109517_(_050706_, _050718_, _050735_);
  or g_109518_(_050734_, _050735_, _050736_);
  or g_109519_(_050711_, _050716_, _050737_);
  or g_109520_(_050719_, _050737_, _050738_);
  or g_109521_(_050736_, _050738_, _050739_);
  or g_109522_(_050732_, _050739_, _050740_);
  or g_109523_(_050724_, _050740_, _050741_);
  not g_109524_(_050741_, _050743_);
  xor g_109525_(out[369], out[785], _050744_);
  and g_109526_(_049422_, out[795], _050745_);
  and g_109527_(out[379], _049708_, _050746_);
  xor g_109528_(out[382], out[798], _050747_);
  xor g_109529_(out[371], out[787], _050748_);
  xor g_109530_(out[372], out[788], _050749_);
  xor g_109531_(out[370], out[786], _050750_);
  xor g_109532_(out[377], out[793], _050751_);
  xor g_109533_(out[368], out[784], _050752_);
  xor g_109534_(out[380], out[796], _050754_);
  xor g_109535_(out[374], out[790], _050755_);
  xor g_109536_(out[378], out[794], _050756_);
  xor g_109537_(out[373], out[789], _050757_);
  xor g_109538_(out[383], out[799], _050758_);
  xor g_109539_(out[381], out[797], _050759_);
  xor g_109540_(out[376], out[792], _050760_);
  or g_109541_(_050747_, _050749_, _050761_);
  or g_109542_(_050759_, _050760_, _050762_);
  or g_109543_(_050750_, _050756_, _050763_);
  or g_109544_(_050762_, _050763_, _050765_);
  or g_109545_(_050748_, _050751_, _050766_);
  or g_109546_(_050752_, _050757_, _050767_);
  or g_109547_(_050766_, _050767_, _050768_);
  or g_109548_(_050765_, _050768_, _050769_);
  or g_109549_(_050745_, _050754_, _050770_);
  xor g_109550_(out[375], out[791], _050771_);
  or g_109551_(_050755_, _050771_, _050772_);
  or g_109552_(_050770_, _050772_, _050773_);
  or g_109553_(_050744_, _050746_, _050774_);
  or g_109554_(_050758_, _050774_, _050776_);
  or g_109555_(_050773_, _050776_, _050777_);
  or g_109556_(_050769_, _050777_, _050778_);
  or g_109557_(_050761_, _050778_, _050779_);
  not g_109558_(_050779_, _050780_);
  xor g_109559_(out[359], out[791], _050781_);
  and g_109560_(_049411_, out[795], _050782_);
  xor g_109561_(out[366], out[798], _050783_);
  xor g_109562_(out[360], out[792], _050784_);
  xor g_109563_(out[353], out[785], _050785_);
  xor g_109564_(out[365], out[797], _050787_);
  xor g_109565_(out[361], out[793], _050788_);
  xor g_109566_(out[356], out[788], _050789_);
  xor g_109567_(out[354], out[786], _050790_);
  and g_109568_(out[363], _049708_, _050791_);
  xor g_109569_(out[355], out[787], _050792_);
  xor g_109570_(out[358], out[790], _050793_);
  xor g_109571_(out[367], out[799], _050794_);
  xor g_109572_(out[362], out[794], _050795_);
  xor g_109573_(out[357], out[789], _050796_);
  xor g_109574_(out[352], out[784], _050798_);
  or g_109575_(_050783_, _050789_, _050799_);
  or g_109576_(_050784_, _050787_, _050800_);
  or g_109577_(_050790_, _050795_, _050801_);
  or g_109578_(_050800_, _050801_, _050802_);
  or g_109579_(_050788_, _050792_, _050803_);
  or g_109580_(_050796_, _050798_, _050804_);
  or g_109581_(_050803_, _050804_, _050805_);
  or g_109582_(_050802_, _050805_, _050806_);
  xor g_109583_(out[364], out[796], _050807_);
  or g_109584_(_050782_, _050807_, _050809_);
  or g_109585_(_050781_, _050793_, _050810_);
  or g_109586_(_050809_, _050810_, _050811_);
  or g_109587_(_050785_, _050791_, _050812_);
  or g_109588_(_050794_, _050812_, _050813_);
  or g_109589_(_050811_, _050813_, _050814_);
  or g_109590_(_050806_, _050814_, _050815_);
  or g_109591_(_050799_, _050815_, _050816_);
  not g_109592_(_050816_, _050817_);
  xor g_109593_(out[339], out[787], _050818_);
  xor g_109594_(out[340], out[788], _050820_);
  xor g_109595_(out[350], out[798], _050821_);
  xor g_109596_(out[338], out[786], _050822_);
  xor g_109597_(out[341], out[789], _050823_);
  xor g_109598_(out[345], out[793], _050824_);
  xor g_109599_(out[344], out[792], _050825_);
  xor g_109600_(out[351], out[799], _050826_);
  xor g_109601_(out[346], out[794], _050827_);
  xor g_109602_(out[342], out[790], _050828_);
  xor g_109603_(out[336], out[784], _050829_);
  and g_109604_(_049400_, out[795], _050831_);
  and g_109605_(out[347], _049708_, _050832_);
  xor g_109606_(out[349], out[797], _050833_);
  or g_109607_(_050825_, _050833_, _050834_);
  xor g_109608_(out[337], out[785], _050835_);
  or g_109609_(_050822_, _050827_, _050836_);
  or g_109610_(_050834_, _050836_, _050837_);
  or g_109611_(_050818_, _050824_, _050838_);
  or g_109612_(_050823_, _050838_, _050839_);
  or g_109613_(_050837_, _050839_, _050840_);
  or g_109614_(_050820_, _050821_, _050842_);
  or g_109615_(_050840_, _050842_, _050843_);
  xor g_109616_(out[348], out[796], _050844_);
  or g_109617_(_050831_, _050844_, _050845_);
  xor g_109618_(out[343], out[791], _050846_);
  or g_109619_(_050828_, _050846_, _050847_);
  or g_109620_(_050845_, _050847_, _050848_);
  or g_109621_(_050832_, _050835_, _050849_);
  or g_109622_(_050826_, _050849_, _050850_);
  or g_109623_(_050848_, _050850_, _050851_);
  or g_109624_(_050829_, _050851_, _050853_);
  or g_109625_(_050843_, _050853_, _050854_);
  not g_109626_(_050854_, _050855_);
  xor g_109627_(out[327], out[791], _050856_);
  and g_109628_(_098294_, out[795], _050857_);
  xor g_109629_(out[334], out[798], _050858_);
  xor g_109630_(out[328], out[792], _050859_);
  xor g_109631_(out[321], out[785], _050860_);
  xor g_109632_(out[333], out[797], _050861_);
  xor g_109633_(out[329], out[793], _050862_);
  xor g_109634_(out[324], out[788], _050864_);
  xor g_109635_(out[322], out[786], _050865_);
  and g_109636_(out[331], _049708_, _050866_);
  xor g_109637_(out[323], out[787], _050867_);
  xor g_109638_(out[326], out[790], _050868_);
  xor g_109639_(out[335], out[799], _050869_);
  xor g_109640_(out[330], out[794], _050870_);
  xor g_109641_(out[325], out[789], _050871_);
  xor g_109642_(out[320], out[784], _050872_);
  or g_109643_(_050858_, _050864_, _050873_);
  or g_109644_(_050859_, _050861_, _050875_);
  or g_109645_(_050865_, _050870_, _050876_);
  or g_109646_(_050875_, _050876_, _050877_);
  or g_109647_(_050862_, _050867_, _050878_);
  or g_109648_(_050871_, _050872_, _050879_);
  or g_109649_(_050878_, _050879_, _050880_);
  or g_109650_(_050877_, _050880_, _050881_);
  xor g_109651_(out[332], out[796], _050882_);
  or g_109652_(_050857_, _050882_, _050883_);
  or g_109653_(_050856_, _050868_, _050884_);
  or g_109654_(_050883_, _050884_, _050886_);
  or g_109655_(_050860_, _050866_, _050887_);
  or g_109656_(_050869_, _050887_, _050888_);
  or g_109657_(_050886_, _050888_, _050889_);
  or g_109658_(_050881_, _050889_, _050890_);
  or g_109659_(_050873_, _050890_, _050891_);
  xor g_109660_(out[316], out[796], _050892_);
  and g_109661_(_098283_, out[795], _050893_);
  xor g_109662_(out[312], out[792], _050894_);
  xor g_109663_(out[310], out[790], _050895_);
  xor g_109664_(out[317], out[797], _050897_);
  xor g_109665_(out[318], out[798], _050898_);
  xor g_109666_(out[306], out[786], _050899_);
  xor g_109667_(out[313], out[793], _050900_);
  xor g_109668_(out[309], out[789], _050901_);
  xor g_109669_(out[305], out[785], _050902_);
  and g_109670_(out[315], _049708_, _050903_);
  or g_109671_(_050894_, _050897_, _050904_);
  xor g_109672_(out[319], out[799], _050905_);
  xor g_109673_(out[314], out[794], _050906_);
  xor g_109674_(out[308], out[788], _050908_);
  xor g_109675_(out[307], out[787], _050909_);
  xor g_109676_(out[304], out[784], _050910_);
  or g_109677_(_050899_, _050906_, _050911_);
  or g_109678_(_050904_, _050911_, _050912_);
  or g_109679_(_050900_, _050909_, _050913_);
  or g_109680_(_050901_, _050913_, _050914_);
  or g_109681_(_050912_, _050914_, _050915_);
  or g_109682_(_050898_, _050908_, _050916_);
  or g_109683_(_050915_, _050916_, _050917_);
  or g_109684_(_050892_, _050893_, _050919_);
  xor g_109685_(out[311], out[791], _050920_);
  or g_109686_(_050895_, _050920_, _050921_);
  or g_109687_(_050919_, _050921_, _050922_);
  or g_109688_(_050902_, _050903_, _050923_);
  or g_109689_(_050905_, _050923_, _050924_);
  or g_109690_(_050922_, _050924_, _050925_);
  or g_109691_(_050910_, _050925_, _050926_);
  or g_109692_(_050917_, _050926_, _050927_);
  not g_109693_(_050927_, _050928_);
  xor g_109694_(out[295], out[791], _050930_);
  and g_109695_(_098272_, out[795], _050931_);
  xor g_109696_(out[302], out[798], _050932_);
  xor g_109697_(out[296], out[792], _050933_);
  xor g_109698_(out[289], out[785], _050934_);
  xor g_109699_(out[301], out[797], _050935_);
  xor g_109700_(out[297], out[793], _050936_);
  xor g_109701_(out[292], out[788], _050937_);
  xor g_109702_(out[290], out[786], _050938_);
  and g_109703_(out[299], _049708_, _050939_);
  xor g_109704_(out[291], out[787], _050941_);
  xor g_109705_(out[294], out[790], _050942_);
  xor g_109706_(out[303], out[799], _050943_);
  xor g_109707_(out[298], out[794], _050944_);
  xor g_109708_(out[293], out[789], _050945_);
  xor g_109709_(out[288], out[784], _050946_);
  or g_109710_(_050932_, _050937_, _050947_);
  or g_109711_(_050933_, _050935_, _050948_);
  or g_109712_(_050938_, _050944_, _050949_);
  or g_109713_(_050948_, _050949_, _050950_);
  or g_109714_(_050936_, _050941_, _050952_);
  or g_109715_(_050945_, _050946_, _050953_);
  or g_109716_(_050952_, _050953_, _050954_);
  or g_109717_(_050950_, _050954_, _050955_);
  xor g_109718_(out[300], out[796], _050956_);
  or g_109719_(_050931_, _050956_, _050957_);
  or g_109720_(_050930_, _050942_, _050958_);
  or g_109721_(_050957_, _050958_, _050959_);
  or g_109722_(_050934_, _050939_, _050960_);
  or g_109723_(_050943_, _050960_, _050961_);
  or g_109724_(_050959_, _050961_, _050963_);
  or g_109725_(_050955_, _050963_, _050964_);
  or g_109726_(_050947_, _050964_, _050965_);
  not g_109727_(_050965_, _050966_);
  xor g_109728_(out[280], out[792], _050967_);
  xor g_109729_(out[277], out[789], _050968_);
  xor g_109730_(out[275], out[787], _050969_);
  xor g_109731_(out[286], out[798], _050970_);
  xor g_109732_(out[285], out[797], _050971_);
  xor g_109733_(out[274], out[786], _050972_);
  xor g_109734_(out[281], out[793], _050974_);
  xor g_109735_(out[278], out[790], _050975_);
  xor g_109736_(out[287], out[799], _050976_);
  xor g_109737_(out[282], out[794], _050977_);
  xor g_109738_(out[276], out[788], _050978_);
  xor g_109739_(out[272], out[784], _050979_);
  and g_109740_(_098261_, out[795], _050980_);
  and g_109741_(out[283], _049708_, _050981_);
  or g_109742_(_050967_, _050971_, _050982_);
  xor g_109743_(out[273], out[785], _050983_);
  or g_109744_(_050972_, _050977_, _050985_);
  or g_109745_(_050982_, _050985_, _050986_);
  or g_109746_(_050969_, _050974_, _050987_);
  or g_109747_(_050968_, _050987_, _050988_);
  or g_109748_(_050986_, _050988_, _050989_);
  or g_109749_(_050970_, _050978_, _050990_);
  or g_109750_(_050989_, _050990_, _050991_);
  xor g_109751_(out[284], out[796], _050992_);
  or g_109752_(_050980_, _050992_, _050993_);
  xor g_109753_(out[279], out[791], _050994_);
  or g_109754_(_050975_, _050994_, _050996_);
  or g_109755_(_050993_, _050996_, _050997_);
  or g_109756_(_050981_, _050983_, _050998_);
  or g_109757_(_050976_, _050998_, _050999_);
  or g_109758_(_050997_, _050999_, _051000_);
  or g_109759_(_050979_, _051000_, _051001_);
  or g_109760_(_050991_, _051001_, _051002_);
  xor g_109761_(out[263], out[791], _051003_);
  and g_109762_(_098250_, out[795], _051004_);
  xor g_109763_(out[270], out[798], _051005_);
  xor g_109764_(out[264], out[792], _051007_);
  xor g_109765_(out[257], out[785], _051008_);
  xor g_109766_(out[269], out[797], _051009_);
  xor g_109767_(out[265], out[793], _051010_);
  xor g_109768_(out[260], out[788], _051011_);
  xor g_109769_(out[258], out[786], _051012_);
  and g_109770_(out[267], _049708_, _051013_);
  xor g_109771_(out[259], out[787], _051014_);
  xor g_109772_(out[262], out[790], _051015_);
  xor g_109773_(out[271], out[799], _051016_);
  xor g_109774_(out[266], out[794], _051018_);
  xor g_109775_(out[261], out[789], _051019_);
  xor g_109776_(out[256], out[784], _051020_);
  or g_109777_(_051005_, _051011_, _051021_);
  or g_109778_(_051007_, _051009_, _051022_);
  or g_109779_(_051012_, _051018_, _051023_);
  or g_109780_(_051022_, _051023_, _051024_);
  or g_109781_(_051010_, _051014_, _051025_);
  or g_109782_(_051019_, _051020_, _051026_);
  or g_109783_(_051025_, _051026_, _051027_);
  or g_109784_(_051024_, _051027_, _051029_);
  xor g_109785_(out[268], out[796], _051030_);
  or g_109786_(_051004_, _051030_, _051031_);
  or g_109787_(_051003_, _051015_, _051032_);
  or g_109788_(_051031_, _051032_, _051033_);
  or g_109789_(_051008_, _051013_, _051034_);
  or g_109790_(_051016_, _051034_, _051035_);
  or g_109791_(_051033_, _051035_, _051036_);
  or g_109792_(_051029_, _051036_, _051037_);
  or g_109793_(_051021_, _051037_, _051038_);
  xor g_109794_(out[252], out[796], _051040_);
  and g_109795_(_098239_, out[795], _051041_);
  xor g_109796_(out[248], out[792], _051042_);
  xor g_109797_(out[246], out[790], _051043_);
  xor g_109798_(out[253], out[797], _051044_);
  xor g_109799_(out[254], out[798], _051045_);
  xor g_109800_(out[242], out[786], _051046_);
  xor g_109801_(out[249], out[793], _051047_);
  xor g_109802_(out[245], out[789], _051048_);
  xor g_109803_(out[241], out[785], _051049_);
  and g_109804_(out[251], _049708_, _051051_);
  or g_109805_(_051042_, _051044_, _051052_);
  xor g_109806_(out[255], out[799], _051053_);
  xor g_109807_(out[250], out[794], _051054_);
  xor g_109808_(out[244], out[788], _051055_);
  xor g_109809_(out[243], out[787], _051056_);
  xor g_109810_(out[240], out[784], _051057_);
  or g_109811_(_051046_, _051054_, _051058_);
  or g_109812_(_051052_, _051058_, _051059_);
  or g_109813_(_051047_, _051056_, _051060_);
  or g_109814_(_051048_, _051060_, _051062_);
  or g_109815_(_051059_, _051062_, _051063_);
  or g_109816_(_051045_, _051055_, _051064_);
  or g_109817_(_051063_, _051064_, _051065_);
  or g_109818_(_051040_, _051041_, _051066_);
  xor g_109819_(out[247], out[791], _051067_);
  or g_109820_(_051043_, _051067_, _051068_);
  or g_109821_(_051066_, _051068_, _051069_);
  or g_109822_(_051049_, _051051_, _051070_);
  or g_109823_(_051053_, _051070_, _051071_);
  or g_109824_(_051069_, _051071_, _051073_);
  or g_109825_(_051057_, _051073_, _051074_);
  or g_109826_(_051065_, _051074_, _051075_);
  xor g_109827_(out[231], out[791], _051076_);
  and g_109828_(_098228_, out[795], _051077_);
  xor g_109829_(out[238], out[798], _051078_);
  xor g_109830_(out[232], out[792], _051079_);
  xor g_109831_(out[225], out[785], _051080_);
  xor g_109832_(out[237], out[797], _051081_);
  xor g_109833_(out[233], out[793], _051082_);
  xor g_109834_(out[228], out[788], _051084_);
  xor g_109835_(out[226], out[786], _051085_);
  and g_109836_(out[235], _049708_, _051086_);
  xor g_109837_(out[227], out[787], _051087_);
  xor g_109838_(out[230], out[790], _051088_);
  xor g_109839_(out[239], out[799], _051089_);
  xor g_109840_(out[234], out[794], _051090_);
  xor g_109841_(out[229], out[789], _051091_);
  xor g_109842_(out[224], out[784], _051092_);
  or g_109843_(_051078_, _051084_, _051093_);
  or g_109844_(_051079_, _051081_, _051095_);
  or g_109845_(_051085_, _051090_, _051096_);
  or g_109846_(_051095_, _051096_, _051097_);
  or g_109847_(_051082_, _051087_, _051098_);
  or g_109848_(_051091_, _051092_, _051099_);
  or g_109849_(_051098_, _051099_, _051100_);
  or g_109850_(_051097_, _051100_, _051101_);
  xor g_109851_(out[236], out[796], _051102_);
  or g_109852_(_051077_, _051102_, _051103_);
  or g_109853_(_051076_, _051088_, _051104_);
  or g_109854_(_051103_, _051104_, _051106_);
  or g_109855_(_051080_, _051086_, _051107_);
  or g_109856_(_051089_, _051107_, _051108_);
  or g_109857_(_051106_, _051108_, _051109_);
  or g_109858_(_051101_, _051109_, _051110_);
  or g_109859_(_051093_, _051110_, _051111_);
  not g_109860_(_051111_, _051112_);
  xor g_109861_(out[209], out[785], _051113_);
  and g_109862_(_098217_, out[795], _051114_);
  and g_109863_(out[219], _049708_, _051115_);
  xor g_109864_(out[217], out[793], _051117_);
  xor g_109865_(out[208], out[784], _051118_);
  xor g_109866_(out[222], out[798], _051119_);
  xor g_109867_(out[212], out[788], _051120_);
  or g_109868_(_051119_, _051120_, _051121_);
  xor g_109869_(out[221], out[797], _051122_);
  xor g_109870_(out[211], out[787], _051123_);
  xor g_109871_(out[220], out[796], _051124_);
  xor g_109872_(out[214], out[790], _051125_);
  xor g_109873_(out[218], out[794], _051126_);
  xor g_109874_(out[213], out[789], _051128_);
  xor g_109875_(out[223], out[799], _051129_);
  xor g_109876_(out[216], out[792], _051130_);
  or g_109877_(_051122_, _051130_, _051131_);
  xor g_109878_(out[210], out[786], _051132_);
  or g_109879_(_051126_, _051132_, _051133_);
  or g_109880_(_051131_, _051133_, _051134_);
  or g_109881_(_051117_, _051123_, _051135_);
  or g_109882_(_051128_, _051135_, _051136_);
  or g_109883_(_051134_, _051136_, _051137_);
  or g_109884_(_051121_, _051137_, _051139_);
  or g_109885_(_051114_, _051124_, _051140_);
  xor g_109886_(out[215], out[791], _051141_);
  or g_109887_(_051125_, _051141_, _051142_);
  or g_109888_(_051140_, _051142_, _051143_);
  or g_109889_(_051113_, _051115_, _051144_);
  or g_109890_(_051129_, _051144_, _051145_);
  or g_109891_(_051143_, _051145_, _051146_);
  or g_109892_(_051118_, _051146_, _051147_);
  or g_109893_(_051139_, _051147_, _051148_);
  not g_109894_(_051148_, _051150_);
  xor g_109895_(out[199], out[791], _051151_);
  and g_109896_(_098206_, out[795], _051152_);
  xor g_109897_(out[206], out[798], _051153_);
  xor g_109898_(out[200], out[792], _051154_);
  xor g_109899_(out[193], out[785], _051155_);
  xor g_109900_(out[205], out[797], _051156_);
  xor g_109901_(out[201], out[793], _051157_);
  xor g_109902_(out[196], out[788], _051158_);
  xor g_109903_(out[194], out[786], _051159_);
  and g_109904_(out[203], _049708_, _051161_);
  xor g_109905_(out[195], out[787], _051162_);
  xor g_109906_(out[198], out[790], _051163_);
  xor g_109907_(out[207], out[799], _051164_);
  xor g_109908_(out[202], out[794], _051165_);
  xor g_109909_(out[197], out[789], _051166_);
  xor g_109910_(out[192], out[784], _051167_);
  or g_109911_(_051153_, _051158_, _051168_);
  or g_109912_(_051154_, _051156_, _051169_);
  or g_109913_(_051159_, _051165_, _051170_);
  or g_109914_(_051169_, _051170_, _051172_);
  or g_109915_(_051157_, _051162_, _051173_);
  or g_109916_(_051166_, _051167_, _051174_);
  or g_109917_(_051173_, _051174_, _051175_);
  or g_109918_(_051172_, _051175_, _051176_);
  xor g_109919_(out[204], out[796], _051177_);
  or g_109920_(_051152_, _051177_, _051178_);
  or g_109921_(_051151_, _051163_, _051179_);
  or g_109922_(_051178_, _051179_, _051180_);
  or g_109923_(_051155_, _051161_, _051181_);
  or g_109924_(_051164_, _051181_, _051183_);
  or g_109925_(_051180_, _051183_, _051184_);
  or g_109926_(_051176_, _051184_, _051185_);
  or g_109927_(_051168_, _051185_, _051186_);
  xor g_109928_(out[186], out[794], _051187_);
  xor g_109929_(out[178], out[786], _051188_);
  xor g_109930_(out[177], out[785], _051189_);
  and g_109931_(_098195_, out[795], _051190_);
  and g_109932_(out[187], _049708_, _051191_);
  xor g_109933_(out[189], out[797], _051192_);
  xor g_109934_(out[179], out[787], _051194_);
  xor g_109935_(out[190], out[798], _051195_);
  xor g_109936_(out[188], out[796], _051196_);
  xor g_109937_(out[184], out[792], _051197_);
  xor g_109938_(out[191], out[799], _051198_);
  xor g_109939_(out[181], out[789], _051199_);
  xor g_109940_(out[182], out[790], _051200_);
  xor g_109941_(out[176], out[784], _051201_);
  xor g_109942_(out[180], out[788], _051202_);
  or g_109943_(_051192_, _051197_, _051203_);
  xor g_109944_(out[185], out[793], _051205_);
  or g_109945_(_051187_, _051188_, _051206_);
  or g_109946_(_051203_, _051206_, _051207_);
  or g_109947_(_051194_, _051205_, _051208_);
  or g_109948_(_051199_, _051208_, _051209_);
  or g_109949_(_051207_, _051209_, _051210_);
  or g_109950_(_051195_, _051202_, _051211_);
  or g_109951_(_051210_, _051211_, _051212_);
  or g_109952_(_051190_, _051196_, _051213_);
  xor g_109953_(out[183], out[791], _051214_);
  or g_109954_(_051200_, _051214_, _051216_);
  or g_109955_(_051213_, _051216_, _051217_);
  or g_109956_(_051189_, _051191_, _051218_);
  or g_109957_(_051198_, _051218_, _051219_);
  or g_109958_(_051217_, _051219_, _051220_);
  or g_109959_(_051201_, _051220_, _051221_);
  or g_109960_(_051212_, _051221_, _051222_);
  xor g_109961_(out[167], out[791], _051223_);
  and g_109962_(_098184_, out[795], _051224_);
  xor g_109963_(out[174], out[798], _051225_);
  xor g_109964_(out[168], out[792], _051227_);
  xor g_109965_(out[161], out[785], _051228_);
  xor g_109966_(out[173], out[797], _051229_);
  xor g_109967_(out[169], out[793], _051230_);
  xor g_109968_(out[164], out[788], _051231_);
  xor g_109969_(out[162], out[786], _051232_);
  and g_109970_(out[171], _049708_, _051233_);
  xor g_109971_(out[163], out[787], _051234_);
  xor g_109972_(out[166], out[790], _051235_);
  xor g_109973_(out[175], out[799], _051236_);
  xor g_109974_(out[170], out[794], _051238_);
  xor g_109975_(out[165], out[789], _051239_);
  xor g_109976_(out[160], out[784], _051240_);
  or g_109977_(_051225_, _051231_, _051241_);
  or g_109978_(_051227_, _051229_, _051242_);
  or g_109979_(_051232_, _051238_, _051243_);
  or g_109980_(_051242_, _051243_, _051244_);
  or g_109981_(_051230_, _051234_, _051245_);
  or g_109982_(_051239_, _051240_, _051246_);
  or g_109983_(_051245_, _051246_, _051247_);
  or g_109984_(_051244_, _051247_, _051249_);
  xor g_109985_(out[172], out[796], _051250_);
  or g_109986_(_051224_, _051250_, _051251_);
  or g_109987_(_051223_, _051235_, _051252_);
  or g_109988_(_051251_, _051252_, _051253_);
  or g_109989_(_051228_, _051233_, _051254_);
  or g_109990_(_051236_, _051254_, _051255_);
  or g_109991_(_051253_, _051255_, _051256_);
  or g_109992_(_051249_, _051256_, _051257_);
  or g_109993_(_051241_, _051257_, _051258_);
  not g_109994_(_051258_, _051260_);
  xor g_109995_(out[157], out[797], _051261_);
  xor g_109996_(out[146], out[786], _051262_);
  xor g_109997_(out[149], out[789], _051263_);
  xor g_109998_(out[153], out[793], _051264_);
  xor g_109999_(out[148], out[788], _051265_);
  xor g_110000_(out[152], out[792], _051266_);
  xor g_110001_(out[158], out[798], _051267_);
  xor g_110002_(out[150], out[790], _051268_);
  xor g_110003_(out[159], out[799], _051269_);
  xor g_110004_(out[154], out[794], _051271_);
  xor g_110005_(out[144], out[784], _051272_);
  xor g_110006_(out[147], out[787], _051273_);
  and g_110007_(_098173_, out[795], _051274_);
  and g_110008_(out[155], _049708_, _051275_);
  xor g_110009_(out[145], out[785], _051276_);
  or g_110010_(_051265_, _051267_, _051277_);
  or g_110011_(_051261_, _051266_, _051278_);
  or g_110012_(_051262_, _051271_, _051279_);
  or g_110013_(_051278_, _051279_, _051280_);
  or g_110014_(_051264_, _051273_, _051282_);
  or g_110015_(_051263_, _051272_, _051283_);
  or g_110016_(_051282_, _051283_, _051284_);
  or g_110017_(_051280_, _051284_, _051285_);
  xor g_110018_(out[156], out[796], _051286_);
  or g_110019_(_051274_, _051286_, _051287_);
  xor g_110020_(out[151], out[791], _051288_);
  or g_110021_(_051268_, _051288_, _051289_);
  or g_110022_(_051287_, _051289_, _051290_);
  or g_110023_(_051275_, _051276_, _051291_);
  or g_110024_(_051269_, _051291_, _051293_);
  or g_110025_(_051290_, _051293_, _051294_);
  or g_110026_(_051285_, _051294_, _051295_);
  or g_110027_(_051277_, _051295_, _051296_);
  xor g_110028_(out[135], out[791], _051297_);
  and g_110029_(_098162_, out[795], _051298_);
  xor g_110030_(out[142], out[798], _051299_);
  xor g_110031_(out[136], out[792], _051300_);
  xor g_110032_(out[129], out[785], _051301_);
  xor g_110033_(out[141], out[797], _051302_);
  xor g_110034_(out[137], out[793], _051304_);
  xor g_110035_(out[132], out[788], _051305_);
  xor g_110036_(out[130], out[786], _051306_);
  and g_110037_(out[139], _049708_, _051307_);
  xor g_110038_(out[131], out[787], _051308_);
  xor g_110039_(out[134], out[790], _051309_);
  xor g_110040_(out[143], out[799], _051310_);
  xor g_110041_(out[138], out[794], _051311_);
  xor g_110042_(out[133], out[789], _051312_);
  xor g_110043_(out[128], out[784], _051313_);
  or g_110044_(_051299_, _051305_, _051315_);
  or g_110045_(_051300_, _051302_, _051316_);
  or g_110046_(_051306_, _051311_, _051317_);
  or g_110047_(_051316_, _051317_, _051318_);
  or g_110048_(_051304_, _051308_, _051319_);
  or g_110049_(_051312_, _051313_, _051320_);
  or g_110050_(_051319_, _051320_, _051321_);
  or g_110051_(_051318_, _051321_, _051322_);
  xor g_110052_(out[140], out[796], _051323_);
  or g_110053_(_051298_, _051323_, _051324_);
  or g_110054_(_051297_, _051309_, _051326_);
  or g_110055_(_051324_, _051326_, _051327_);
  or g_110056_(_051301_, _051307_, _051328_);
  or g_110057_(_051310_, _051328_, _051329_);
  or g_110058_(_051327_, _051329_, _051330_);
  or g_110059_(_051322_, _051330_, _051331_);
  or g_110060_(_051315_, _051331_, _051332_);
  not g_110061_(_051332_, _051333_);
  xor g_110062_(out[113], out[785], _051334_);
  and g_110063_(out[123], _049708_, _051335_);
  xor g_110064_(out[126], out[798], _051337_);
  xor g_110065_(out[115], out[787], _051338_);
  xor g_110066_(out[116], out[788], _051339_);
  xor g_110067_(out[114], out[786], _051340_);
  xor g_110068_(out[121], out[793], _051341_);
  xor g_110069_(out[112], out[784], _051342_);
  and g_110070_(_098151_, out[795], _051343_);
  xor g_110071_(out[118], out[790], _051344_);
  xor g_110072_(out[122], out[794], _051345_);
  xor g_110073_(out[117], out[789], _051346_);
  xor g_110074_(out[127], out[799], _051348_);
  xor g_110075_(out[125], out[797], _051349_);
  xor g_110076_(out[120], out[792], _051350_);
  or g_110077_(_051337_, _051339_, _051351_);
  or g_110078_(_051349_, _051350_, _051352_);
  or g_110079_(_051340_, _051345_, _051353_);
  or g_110080_(_051352_, _051353_, _051354_);
  or g_110081_(_051338_, _051341_, _051355_);
  or g_110082_(_051342_, _051346_, _051356_);
  or g_110083_(_051355_, _051356_, _051357_);
  or g_110084_(_051354_, _051357_, _051359_);
  xor g_110085_(out[124], out[796], _051360_);
  or g_110086_(_051343_, _051360_, _051361_);
  xor g_110087_(out[119], out[791], _051362_);
  or g_110088_(_051344_, _051362_, _051363_);
  or g_110089_(_051361_, _051363_, _051364_);
  or g_110090_(_051334_, _051335_, _051365_);
  or g_110091_(_051348_, _051365_, _051366_);
  or g_110092_(_051364_, _051366_, _051367_);
  or g_110093_(_051359_, _051367_, _051368_);
  or g_110094_(_051351_, _051368_, _051370_);
  xor g_110095_(out[103], out[791], _051371_);
  and g_110096_(_098140_, out[795], _051372_);
  xor g_110097_(out[110], out[798], _051373_);
  xor g_110098_(out[104], out[792], _051374_);
  xor g_110099_(out[97], out[785], _051375_);
  xor g_110100_(out[109], out[797], _051376_);
  xor g_110101_(out[105], out[793], _051377_);
  xor g_110102_(out[100], out[788], _051378_);
  xor g_110103_(out[98], out[786], _051379_);
  and g_110104_(out[107], _049708_, _051381_);
  xor g_110105_(out[99], out[787], _051382_);
  xor g_110106_(out[102], out[790], _051383_);
  xor g_110107_(out[111], out[799], _051384_);
  xor g_110108_(out[106], out[794], _051385_);
  xor g_110109_(out[101], out[789], _051386_);
  xor g_110110_(out[96], out[784], _051387_);
  or g_110111_(_051373_, _051378_, _051388_);
  or g_110112_(_051374_, _051376_, _051389_);
  or g_110113_(_051379_, _051385_, _051390_);
  or g_110114_(_051389_, _051390_, _051392_);
  or g_110115_(_051377_, _051382_, _051393_);
  or g_110116_(_051386_, _051387_, _051394_);
  or g_110117_(_051393_, _051394_, _051395_);
  or g_110118_(_051392_, _051395_, _051396_);
  xor g_110119_(out[108], out[796], _051397_);
  or g_110120_(_051372_, _051397_, _051398_);
  or g_110121_(_051371_, _051383_, _051399_);
  or g_110122_(_051398_, _051399_, _051400_);
  or g_110123_(_051375_, _051381_, _051401_);
  or g_110124_(_051384_, _051401_, _051403_);
  or g_110125_(_051400_, _051403_, _051404_);
  or g_110126_(_051396_, _051404_, _051405_);
  or g_110127_(_051388_, _051405_, _051406_);
  xor g_110128_(out[81], out[785], _051407_);
  and g_110129_(out[91], _049708_, _051408_);
  xor g_110130_(out[89], out[793], _051409_);
  xor g_110131_(out[80], out[784], _051410_);
  xor g_110132_(out[94], out[798], _051411_);
  xor g_110133_(out[84], out[788], _051412_);
  or g_110134_(_051411_, _051412_, _051414_);
  xor g_110135_(out[93], out[797], _051415_);
  xor g_110136_(out[83], out[787], _051416_);
  and g_110137_(_098129_, out[795], _051417_);
  xor g_110138_(out[86], out[790], _051418_);
  xor g_110139_(out[90], out[794], _051419_);
  xor g_110140_(out[85], out[789], _051420_);
  xor g_110141_(out[95], out[799], _051421_);
  xor g_110142_(out[88], out[792], _051422_);
  or g_110143_(_051415_, _051422_, _051423_);
  xor g_110144_(out[82], out[786], _051425_);
  or g_110145_(_051419_, _051425_, _051426_);
  or g_110146_(_051423_, _051426_, _051427_);
  or g_110147_(_051409_, _051416_, _051428_);
  or g_110148_(_051420_, _051428_, _051429_);
  or g_110149_(_051427_, _051429_, _051430_);
  or g_110150_(_051414_, _051430_, _051431_);
  xor g_110151_(out[92], out[796], _051432_);
  or g_110152_(_051417_, _051432_, _051433_);
  xor g_110153_(out[87], out[791], _051434_);
  or g_110154_(_051418_, _051434_, _051436_);
  or g_110155_(_051433_, _051436_, _051437_);
  or g_110156_(_051407_, _051408_, _051438_);
  or g_110157_(_051421_, _051438_, _051439_);
  or g_110158_(_051437_, _051439_, _051440_);
  or g_110159_(_051410_, _051440_, _051441_);
  or g_110160_(_051431_, _051441_, _051442_);
  xor g_110161_(out[71], out[791], _051443_);
  and g_110162_(_098118_, out[795], _051444_);
  xor g_110163_(out[78], out[798], _051445_);
  xor g_110164_(out[72], out[792], _051447_);
  xor g_110165_(out[65], out[785], _051448_);
  xor g_110166_(out[77], out[797], _051449_);
  xor g_110167_(out[73], out[793], _051450_);
  xor g_110168_(out[68], out[788], _051451_);
  xor g_110169_(out[66], out[786], _051452_);
  and g_110170_(out[75], _049708_, _051453_);
  xor g_110171_(out[67], out[787], _051454_);
  xor g_110172_(out[70], out[790], _051455_);
  xor g_110173_(out[79], out[799], _051456_);
  xor g_110174_(out[74], out[794], _051458_);
  xor g_110175_(out[69], out[789], _051459_);
  xor g_110176_(out[64], out[784], _051460_);
  or g_110177_(_051445_, _051451_, _051461_);
  or g_110178_(_051447_, _051449_, _051462_);
  or g_110179_(_051452_, _051458_, _051463_);
  or g_110180_(_051462_, _051463_, _051464_);
  or g_110181_(_051450_, _051454_, _051465_);
  or g_110182_(_051459_, _051460_, _051466_);
  or g_110183_(_051465_, _051466_, _051467_);
  or g_110184_(_051464_, _051467_, _051469_);
  xor g_110185_(out[76], out[796], _051470_);
  or g_110186_(_051444_, _051470_, _051471_);
  or g_110187_(_051443_, _051455_, _051472_);
  or g_110188_(_051471_, _051472_, _051473_);
  or g_110189_(_051448_, _051453_, _051474_);
  or g_110190_(_051456_, _051474_, _051475_);
  or g_110191_(_051473_, _051475_, _051476_);
  or g_110192_(_051469_, _051476_, _051477_);
  or g_110193_(_051461_, _051477_, _051478_);
  xor g_110194_(out[56], out[792], _051480_);
  xor g_110195_(out[53], out[789], _051481_);
  xor g_110196_(out[51], out[787], _051482_);
  xor g_110197_(out[62], out[798], _051483_);
  xor g_110198_(out[61], out[797], _051484_);
  xor g_110199_(out[50], out[786], _051485_);
  xor g_110200_(out[57], out[793], _051486_);
  xor g_110201_(out[54], out[790], _051487_);
  xor g_110202_(out[63], out[799], _051488_);
  xor g_110203_(out[58], out[794], _051489_);
  xor g_110204_(out[52], out[788], _051491_);
  xor g_110205_(out[48], out[784], _051492_);
  and g_110206_(_098107_, out[795], _051493_);
  and g_110207_(out[59], _049708_, _051494_);
  or g_110208_(_051480_, _051484_, _051495_);
  xor g_110209_(out[49], out[785], _051496_);
  or g_110210_(_051485_, _051489_, _051497_);
  or g_110211_(_051495_, _051497_, _051498_);
  or g_110212_(_051482_, _051486_, _051499_);
  or g_110213_(_051481_, _051499_, _051500_);
  or g_110214_(_051498_, _051500_, _051502_);
  or g_110215_(_051483_, _051491_, _051503_);
  or g_110216_(_051502_, _051503_, _051504_);
  xor g_110217_(out[60], out[796], _051505_);
  or g_110218_(_051493_, _051505_, _051506_);
  xor g_110219_(out[55], out[791], _051507_);
  or g_110220_(_051487_, _051507_, _051508_);
  or g_110221_(_051506_, _051508_, _051509_);
  or g_110222_(_051494_, _051496_, _051510_);
  or g_110223_(_051488_, _051510_, _051511_);
  or g_110224_(_051509_, _051511_, _051513_);
  or g_110225_(_051492_, _051513_, _051514_);
  or g_110226_(_051504_, _051514_, _051515_);
  not g_110227_(_051515_, _051516_);
  xor g_110228_(out[39], out[791], _051517_);
  and g_110229_(_098096_, out[795], _051518_);
  xor g_110230_(out[46], out[798], _051519_);
  xor g_110231_(out[40], out[792], _051520_);
  xor g_110232_(out[33], out[785], _051521_);
  xor g_110233_(out[45], out[797], _051522_);
  xor g_110234_(out[41], out[793], _051524_);
  xor g_110235_(out[36], out[788], _051525_);
  xor g_110236_(out[34], out[786], _051526_);
  and g_110237_(out[43], _049708_, _051527_);
  xor g_110238_(out[35], out[787], _051528_);
  xor g_110239_(out[38], out[790], _051529_);
  xor g_110240_(out[47], out[799], _051530_);
  xor g_110241_(out[42], out[794], _051531_);
  xor g_110242_(out[37], out[789], _051532_);
  xor g_110243_(out[32], out[784], _051533_);
  or g_110244_(_051519_, _051525_, _051535_);
  or g_110245_(_051520_, _051522_, _051536_);
  or g_110246_(_051526_, _051531_, _051537_);
  or g_110247_(_051536_, _051537_, _051538_);
  or g_110248_(_051524_, _051528_, _051539_);
  or g_110249_(_051532_, _051533_, _051540_);
  or g_110250_(_051539_, _051540_, _051541_);
  or g_110251_(_051538_, _051541_, _051542_);
  xor g_110252_(out[44], out[796], _051543_);
  or g_110253_(_051518_, _051543_, _051544_);
  or g_110254_(_051517_, _051529_, _051546_);
  or g_110255_(_051544_, _051546_, _051547_);
  or g_110256_(_051521_, _051527_, _051548_);
  or g_110257_(_051530_, _051548_, _051549_);
  or g_110258_(_051547_, _051549_, _051550_);
  or g_110259_(_051542_, _051550_, _051551_);
  or g_110260_(_051535_, _051551_, _051552_);
  not g_110261_(_051552_, _051553_);
  and g_110262_(out[27], _049708_, _051554_);
  xor g_110263_(out[20], out[788], _051555_);
  xor g_110264_(out[30], out[798], _051557_);
  or g_110265_(_051555_, _051557_, _051558_);
  xor g_110266_(out[29], out[797], _051559_);
  xor g_110267_(out[19], out[787], _051560_);
  xor g_110268_(out[16], out[784], _051561_);
  and g_110269_(_098063_, out[795], _051562_);
  xor g_110270_(out[26], out[794], _051563_);
  xor g_110271_(out[31], out[799], _051564_);
  xor g_110272_(out[22], out[790], _051565_);
  xor g_110273_(out[21], out[789], _051566_);
  xor g_110274_(out[24], out[792], _051568_);
  or g_110275_(_051559_, _051568_, _051569_);
  xor g_110276_(out[18], out[786], _051570_);
  xor g_110277_(out[25], out[793], _051571_);
  xor g_110278_(out[17], out[785], _051572_);
  or g_110279_(_051563_, _051570_, _051573_);
  or g_110280_(_051569_, _051573_, _051574_);
  or g_110281_(_051560_, _051571_, _051575_);
  or g_110282_(_051566_, _051575_, _051576_);
  or g_110283_(_051574_, _051576_, _051577_);
  or g_110284_(_051558_, _051577_, _051579_);
  xor g_110285_(out[28], out[796], _051580_);
  or g_110286_(_051562_, _051580_, _051581_);
  xor g_110287_(out[23], out[791], _051582_);
  or g_110288_(_051565_, _051582_, _051583_);
  or g_110289_(_051581_, _051583_, _051584_);
  or g_110290_(_051554_, _051572_, _051585_);
  or g_110291_(_051564_, _051585_, _051586_);
  or g_110292_(_051584_, _051586_, _051587_);
  or g_110293_(_051561_, _051587_, _051588_);
  or g_110294_(_051579_, _051588_, _051590_);
  not g_110295_(_051590_, _051591_);
  xor g_110296_(out[1], out[785], _051592_);
  and g_110297_(out[11], _049708_, _051593_);
  xor g_110298_(out[14], out[798], _051594_);
  xor g_110299_(out[3], out[787], _051595_);
  xor g_110300_(out[4], out[788], _051596_);
  xor g_110301_(out[2], out[786], _051597_);
  xor g_110302_(out[9], out[793], _051598_);
  xor g_110303_(out[0], out[784], _051599_);
  and g_110304_(_098041_, out[795], _051601_);
  xor g_110305_(out[6], out[790], _051602_);
  xor g_110306_(out[10], out[794], _051603_);
  xor g_110307_(out[5], out[789], _051604_);
  xor g_110308_(out[15], out[799], _051605_);
  xor g_110309_(out[13], out[797], _051606_);
  xor g_110310_(out[8], out[792], _051607_);
  or g_110311_(_051594_, _051596_, _051608_);
  or g_110312_(_051606_, _051607_, _051609_);
  or g_110313_(_051597_, _051603_, _051610_);
  or g_110314_(_051609_, _051610_, _051612_);
  or g_110315_(_051595_, _051598_, _051613_);
  or g_110316_(_051599_, _051604_, _051614_);
  or g_110317_(_051613_, _051614_, _051615_);
  or g_110318_(_051612_, _051615_, _051616_);
  xor g_110319_(out[12], out[796], _051617_);
  or g_110320_(_051601_, _051617_, _051618_);
  xor g_110321_(out[7], out[791], _051619_);
  or g_110322_(_051602_, _051619_, _051620_);
  or g_110323_(_051618_, _051620_, _051621_);
  or g_110324_(_051592_, _051593_, _051623_);
  or g_110325_(_051605_, _051623_, _051624_);
  or g_110326_(_051621_, _051624_, _051625_);
  or g_110327_(_051616_, _051625_, _051626_);
  or g_110328_(_051608_, _051626_, _051627_);
  xor g_110329_(out[471], out[775], _051628_);
  and g_110330_(_049499_, out[779], _051629_);
  xor g_110331_(out[478], out[782], _051630_);
  xor g_110332_(out[472], out[776], _051631_);
  xor g_110333_(out[465], out[769], _051632_);
  xor g_110334_(out[477], out[781], _051634_);
  xor g_110335_(out[473], out[777], _051635_);
  xor g_110336_(out[468], out[772], _051636_);
  xor g_110337_(out[466], out[770], _051637_);
  and g_110338_(out[475], _049697_, _051638_);
  xor g_110339_(out[467], out[771], _051639_);
  xor g_110340_(out[470], out[774], _051640_);
  xor g_110341_(out[479], out[783], _051641_);
  xor g_110342_(out[474], out[778], _051642_);
  xor g_110343_(out[469], out[773], _051643_);
  xor g_110344_(out[464], out[768], _051645_);
  or g_110345_(_051630_, _051636_, _051646_);
  or g_110346_(_051631_, _051634_, _051647_);
  or g_110347_(_051637_, _051642_, _051648_);
  or g_110348_(_051647_, _051648_, _051649_);
  or g_110349_(_051635_, _051639_, _051650_);
  or g_110350_(_051643_, _051645_, _051651_);
  or g_110351_(_051650_, _051651_, _051652_);
  or g_110352_(_051649_, _051652_, _051653_);
  xor g_110353_(out[476], out[780], _051654_);
  or g_110354_(_051629_, _051654_, _051656_);
  or g_110355_(_051628_, _051640_, _051657_);
  or g_110356_(_051656_, _051657_, _051658_);
  or g_110357_(_051632_, _051638_, _051659_);
  or g_110358_(_051641_, _051659_, _051660_);
  or g_110359_(_051658_, _051660_, _051661_);
  or g_110360_(_051653_, _051661_, _051662_);
  or g_110361_(_051646_, _051662_, _051663_);
  xor g_110362_(out[449], out[769], _051664_);
  and g_110363_(out[459], _049697_, _051665_);
  xor g_110364_(out[457], out[777], _051667_);
  xor g_110365_(out[448], out[768], _051668_);
  xor g_110366_(out[462], out[782], _051669_);
  xor g_110367_(out[452], out[772], _051670_);
  or g_110368_(_051669_, _051670_, _051671_);
  xor g_110369_(out[461], out[781], _051672_);
  xor g_110370_(out[451], out[771], _051673_);
  and g_110371_(_049477_, out[779], _051674_);
  xor g_110372_(out[454], out[774], _051675_);
  xor g_110373_(out[458], out[778], _051676_);
  xor g_110374_(out[453], out[773], _051678_);
  xor g_110375_(out[463], out[783], _051679_);
  xor g_110376_(out[456], out[776], _051680_);
  or g_110377_(_051672_, _051680_, _051681_);
  xor g_110378_(out[450], out[770], _051682_);
  or g_110379_(_051676_, _051682_, _051683_);
  or g_110380_(_051681_, _051683_, _051684_);
  or g_110381_(_051667_, _051673_, _051685_);
  or g_110382_(_051678_, _051685_, _051686_);
  or g_110383_(_051684_, _051686_, _051687_);
  or g_110384_(_051671_, _051687_, _051689_);
  xor g_110385_(out[460], out[780], _051690_);
  or g_110386_(_051674_, _051690_, _051691_);
  xor g_110387_(out[455], out[775], _051692_);
  or g_110388_(_051675_, _051692_, _051693_);
  or g_110389_(_051691_, _051693_, _051694_);
  or g_110390_(_051664_, _051665_, _051695_);
  or g_110391_(_051679_, _051695_, _051696_);
  or g_110392_(_051694_, _051696_, _051697_);
  or g_110393_(_051668_, _051697_, _051698_);
  or g_110394_(_051689_, _051698_, _051700_);
  xor g_110395_(out[439], out[775], _051701_);
  and g_110396_(_049466_, out[779], _051702_);
  xor g_110397_(out[446], out[782], _051703_);
  xor g_110398_(out[440], out[776], _051704_);
  xor g_110399_(out[433], out[769], _051705_);
  xor g_110400_(out[445], out[781], _051706_);
  xor g_110401_(out[441], out[777], _051707_);
  xor g_110402_(out[436], out[772], _051708_);
  xor g_110403_(out[434], out[770], _051709_);
  and g_110404_(out[443], _049697_, _051711_);
  xor g_110405_(out[435], out[771], _051712_);
  xor g_110406_(out[438], out[774], _051713_);
  xor g_110407_(out[447], out[783], _051714_);
  xor g_110408_(out[442], out[778], _051715_);
  xor g_110409_(out[437], out[773], _051716_);
  xor g_110410_(out[432], out[768], _051717_);
  or g_110411_(_051703_, _051708_, _051718_);
  or g_110412_(_051704_, _051706_, _051719_);
  or g_110413_(_051709_, _051715_, _051720_);
  or g_110414_(_051719_, _051720_, _051722_);
  or g_110415_(_051707_, _051712_, _051723_);
  or g_110416_(_051716_, _051717_, _051724_);
  or g_110417_(_051723_, _051724_, _051725_);
  or g_110418_(_051722_, _051725_, _051726_);
  xor g_110419_(out[444], out[780], _051727_);
  or g_110420_(_051702_, _051727_, _051728_);
  or g_110421_(_051701_, _051713_, _051729_);
  or g_110422_(_051728_, _051729_, _051730_);
  or g_110423_(_051705_, _051711_, _051731_);
  or g_110424_(_051714_, _051731_, _051733_);
  or g_110425_(_051730_, _051733_, _051734_);
  or g_110426_(_051726_, _051734_, _051735_);
  or g_110427_(_051718_, _051735_, _051736_);
  xor g_110428_(out[428], out[780], _051737_);
  and g_110429_(_049455_, out[779], _051738_);
  xor g_110430_(out[424], out[776], _051739_);
  xor g_110431_(out[422], out[774], _051740_);
  xor g_110432_(out[429], out[781], _051741_);
  xor g_110433_(out[430], out[782], _051742_);
  xor g_110434_(out[418], out[770], _051744_);
  xor g_110435_(out[425], out[777], _051745_);
  xor g_110436_(out[421], out[773], _051746_);
  xor g_110437_(out[417], out[769], _051747_);
  and g_110438_(out[427], _049697_, _051748_);
  or g_110439_(_051739_, _051741_, _051749_);
  xor g_110440_(out[431], out[783], _051750_);
  xor g_110441_(out[426], out[778], _051751_);
  xor g_110442_(out[420], out[772], _051752_);
  xor g_110443_(out[419], out[771], _051753_);
  xor g_110444_(out[416], out[768], _051755_);
  or g_110445_(_051744_, _051751_, _051756_);
  or g_110446_(_051749_, _051756_, _051757_);
  or g_110447_(_051745_, _051753_, _051758_);
  or g_110448_(_051746_, _051758_, _051759_);
  or g_110449_(_051757_, _051759_, _051760_);
  or g_110450_(_051742_, _051752_, _051761_);
  or g_110451_(_051760_, _051761_, _051762_);
  or g_110452_(_051737_, _051738_, _051763_);
  xor g_110453_(out[423], out[775], _051764_);
  or g_110454_(_051740_, _051764_, _051766_);
  or g_110455_(_051763_, _051766_, _051767_);
  or g_110456_(_051747_, _051748_, _051768_);
  or g_110457_(_051750_, _051768_, _051769_);
  or g_110458_(_051767_, _051769_, _051770_);
  or g_110459_(_051755_, _051770_, _051771_);
  or g_110460_(_051762_, _051771_, _051772_);
  xor g_110461_(out[407], out[775], _051773_);
  and g_110462_(_049444_, out[779], _051774_);
  xor g_110463_(out[414], out[782], _051775_);
  xor g_110464_(out[408], out[776], _051777_);
  xor g_110465_(out[401], out[769], _051778_);
  xor g_110466_(out[413], out[781], _051779_);
  xor g_110467_(out[409], out[777], _051780_);
  xor g_110468_(out[404], out[772], _051781_);
  xor g_110469_(out[402], out[770], _051782_);
  and g_110470_(out[411], _049697_, _051783_);
  xor g_110471_(out[403], out[771], _051784_);
  xor g_110472_(out[406], out[774], _051785_);
  xor g_110473_(out[415], out[783], _051786_);
  xor g_110474_(out[410], out[778], _051788_);
  xor g_110475_(out[405], out[773], _051789_);
  xor g_110476_(out[400], out[768], _051790_);
  or g_110477_(_051775_, _051781_, _051791_);
  or g_110478_(_051777_, _051779_, _051792_);
  or g_110479_(_051782_, _051788_, _051793_);
  or g_110480_(_051792_, _051793_, _051794_);
  or g_110481_(_051780_, _051784_, _051795_);
  or g_110482_(_051789_, _051790_, _051796_);
  or g_110483_(_051795_, _051796_, _051797_);
  or g_110484_(_051794_, _051797_, _051799_);
  xor g_110485_(out[412], out[780], _051800_);
  or g_110486_(_051774_, _051800_, _051801_);
  or g_110487_(_051773_, _051785_, _051802_);
  or g_110488_(_051801_, _051802_, _051803_);
  or g_110489_(_051778_, _051783_, _051804_);
  or g_110490_(_051786_, _051804_, _051805_);
  or g_110491_(_051803_, _051805_, _051806_);
  or g_110492_(_051799_, _051806_, _051807_);
  or g_110493_(_051791_, _051807_, _051808_);
  xor g_110494_(out[385], out[769], _051810_);
  and g_110495_(out[395], _049697_, _051811_);
  xor g_110496_(out[393], out[777], _051812_);
  xor g_110497_(out[384], out[768], _051813_);
  xor g_110498_(out[398], out[782], _051814_);
  xor g_110499_(out[388], out[772], _051815_);
  or g_110500_(_051814_, _051815_, _051816_);
  xor g_110501_(out[397], out[781], _051817_);
  xor g_110502_(out[387], out[771], _051818_);
  and g_110503_(_049433_, out[779], _051819_);
  xor g_110504_(out[390], out[774], _051821_);
  xor g_110505_(out[394], out[778], _051822_);
  xor g_110506_(out[389], out[773], _051823_);
  xor g_110507_(out[399], out[783], _051824_);
  xor g_110508_(out[392], out[776], _051825_);
  or g_110509_(_051817_, _051825_, _051826_);
  xor g_110510_(out[386], out[770], _051827_);
  or g_110511_(_051822_, _051827_, _051828_);
  or g_110512_(_051826_, _051828_, _051829_);
  or g_110513_(_051812_, _051818_, _051830_);
  or g_110514_(_051823_, _051830_, _051832_);
  or g_110515_(_051829_, _051832_, _051833_);
  or g_110516_(_051816_, _051833_, _051834_);
  xor g_110517_(out[396], out[780], _051835_);
  or g_110518_(_051819_, _051835_, _051836_);
  xor g_110519_(out[391], out[775], _051837_);
  or g_110520_(_051821_, _051837_, _051838_);
  or g_110521_(_051836_, _051838_, _051839_);
  or g_110522_(_051810_, _051811_, _051840_);
  or g_110523_(_051824_, _051840_, _051841_);
  or g_110524_(_051839_, _051841_, _051843_);
  or g_110525_(_051813_, _051843_, _051844_);
  or g_110526_(_051834_, _051844_, _051845_);
  xor g_110527_(out[375], out[775], _051846_);
  and g_110528_(_049422_, out[779], _051847_);
  xor g_110529_(out[382], out[782], _051848_);
  xor g_110530_(out[376], out[776], _051849_);
  xor g_110531_(out[369], out[769], _051850_);
  xor g_110532_(out[381], out[781], _051851_);
  xor g_110533_(out[377], out[777], _051852_);
  xor g_110534_(out[372], out[772], _051854_);
  xor g_110535_(out[370], out[770], _051855_);
  and g_110536_(out[379], _049697_, _051856_);
  xor g_110537_(out[371], out[771], _051857_);
  xor g_110538_(out[374], out[774], _051858_);
  xor g_110539_(out[383], out[783], _051859_);
  xor g_110540_(out[378], out[778], _051860_);
  xor g_110541_(out[373], out[773], _051861_);
  xor g_110542_(out[368], out[768], _051862_);
  or g_110543_(_051848_, _051854_, _051863_);
  or g_110544_(_051849_, _051851_, _051865_);
  or g_110545_(_051855_, _051860_, _051866_);
  or g_110546_(_051865_, _051866_, _051867_);
  or g_110547_(_051852_, _051857_, _051868_);
  or g_110548_(_051861_, _051862_, _051869_);
  or g_110549_(_051868_, _051869_, _051870_);
  or g_110550_(_051867_, _051870_, _051871_);
  xor g_110551_(out[380], out[780], _051872_);
  or g_110552_(_051847_, _051872_, _051873_);
  or g_110553_(_051846_, _051858_, _051874_);
  or g_110554_(_051873_, _051874_, _051876_);
  or g_110555_(_051850_, _051856_, _051877_);
  or g_110556_(_051859_, _051877_, _051878_);
  or g_110557_(_051876_, _051878_, _051879_);
  or g_110558_(_051871_, _051879_, _051880_);
  or g_110559_(_051863_, _051880_, _051881_);
  not g_110560_(_051881_, _051882_);
  xor g_110561_(out[360], out[776], _051883_);
  xor g_110562_(out[357], out[773], _051884_);
  xor g_110563_(out[355], out[771], _051885_);
  xor g_110564_(out[366], out[782], _051887_);
  xor g_110565_(out[365], out[781], _051888_);
  xor g_110566_(out[354], out[770], _051889_);
  xor g_110567_(out[361], out[777], _051890_);
  xor g_110568_(out[358], out[774], _051891_);
  xor g_110569_(out[367], out[783], _051892_);
  xor g_110570_(out[362], out[778], _051893_);
  xor g_110571_(out[356], out[772], _051894_);
  xor g_110572_(out[352], out[768], _051895_);
  and g_110573_(_049411_, out[779], _051896_);
  and g_110574_(out[363], _049697_, _051898_);
  or g_110575_(_051883_, _051888_, _051899_);
  xor g_110576_(out[353], out[769], _051900_);
  or g_110577_(_051889_, _051893_, _051901_);
  or g_110578_(_051899_, _051901_, _051902_);
  or g_110579_(_051885_, _051890_, _051903_);
  or g_110580_(_051884_, _051903_, _051904_);
  or g_110581_(_051902_, _051904_, _051905_);
  or g_110582_(_051887_, _051894_, _051906_);
  or g_110583_(_051905_, _051906_, _051907_);
  xor g_110584_(out[364], out[780], _051909_);
  or g_110585_(_051896_, _051909_, _051910_);
  xor g_110586_(out[359], out[775], _051911_);
  or g_110587_(_051891_, _051911_, _051912_);
  or g_110588_(_051910_, _051912_, _051913_);
  or g_110589_(_051898_, _051900_, _051914_);
  or g_110590_(_051892_, _051914_, _051915_);
  or g_110591_(_051913_, _051915_, _051916_);
  or g_110592_(_051895_, _051916_, _051917_);
  or g_110593_(_051907_, _051917_, _051918_);
  not g_110594_(_051918_, _051920_);
  xor g_110595_(out[343], out[775], _051921_);
  and g_110596_(_049400_, out[779], _051922_);
  xor g_110597_(out[350], out[782], _051923_);
  xor g_110598_(out[344], out[776], _051924_);
  xor g_110599_(out[337], out[769], _051925_);
  xor g_110600_(out[349], out[781], _051926_);
  xor g_110601_(out[345], out[777], _051927_);
  xor g_110602_(out[340], out[772], _051928_);
  xor g_110603_(out[338], out[770], _051929_);
  and g_110604_(out[347], _049697_, _051931_);
  xor g_110605_(out[339], out[771], _051932_);
  xor g_110606_(out[342], out[774], _051933_);
  xor g_110607_(out[351], out[783], _051934_);
  xor g_110608_(out[346], out[778], _051935_);
  xor g_110609_(out[341], out[773], _051936_);
  xor g_110610_(out[336], out[768], _051937_);
  or g_110611_(_051923_, _051928_, _051938_);
  or g_110612_(_051924_, _051926_, _051939_);
  or g_110613_(_051929_, _051935_, _051940_);
  or g_110614_(_051939_, _051940_, _051942_);
  or g_110615_(_051927_, _051932_, _051943_);
  or g_110616_(_051936_, _051937_, _051944_);
  or g_110617_(_051943_, _051944_, _051945_);
  or g_110618_(_051942_, _051945_, _051946_);
  xor g_110619_(out[348], out[780], _051947_);
  or g_110620_(_051922_, _051947_, _051948_);
  or g_110621_(_051921_, _051933_, _051949_);
  or g_110622_(_051948_, _051949_, _051950_);
  or g_110623_(_051925_, _051931_, _051951_);
  or g_110624_(_051934_, _051951_, _051953_);
  or g_110625_(_051950_, _051953_, _051954_);
  or g_110626_(_051946_, _051954_, _051955_);
  or g_110627_(_051938_, _051955_, _051956_);
  not g_110628_(_051956_, _051957_);
  xor g_110629_(out[321], out[769], _051958_);
  and g_110630_(out[331], _049697_, _051959_);
  xor g_110631_(out[329], out[777], _051960_);
  xor g_110632_(out[320], out[768], _051961_);
  xor g_110633_(out[334], out[782], _051962_);
  xor g_110634_(out[324], out[772], _051964_);
  or g_110635_(_051962_, _051964_, _051965_);
  xor g_110636_(out[333], out[781], _051966_);
  xor g_110637_(out[323], out[771], _051967_);
  and g_110638_(_098294_, out[779], _051968_);
  xor g_110639_(out[326], out[774], _051969_);
  xor g_110640_(out[330], out[778], _051970_);
  xor g_110641_(out[325], out[773], _051971_);
  xor g_110642_(out[335], out[783], _051972_);
  xor g_110643_(out[328], out[776], _051973_);
  or g_110644_(_051966_, _051973_, _051975_);
  xor g_110645_(out[322], out[770], _051976_);
  or g_110646_(_051970_, _051976_, _051977_);
  or g_110647_(_051975_, _051977_, _051978_);
  or g_110648_(_051960_, _051967_, _051979_);
  or g_110649_(_051971_, _051979_, _051980_);
  or g_110650_(_051978_, _051980_, _051981_);
  or g_110651_(_051965_, _051981_, _051982_);
  xor g_110652_(out[332], out[780], _051983_);
  or g_110653_(_051968_, _051983_, _051984_);
  xor g_110654_(out[327], out[775], _051986_);
  or g_110655_(_051969_, _051986_, _051987_);
  or g_110656_(_051984_, _051987_, _051988_);
  or g_110657_(_051958_, _051959_, _051989_);
  or g_110658_(_051972_, _051989_, _051990_);
  or g_110659_(_051988_, _051990_, _051991_);
  or g_110660_(_051961_, _051991_, _051992_);
  or g_110661_(_051982_, _051992_, _051993_);
  xor g_110662_(out[311], out[775], _051994_);
  and g_110663_(_098283_, out[779], _051995_);
  xor g_110664_(out[318], out[782], _051997_);
  xor g_110665_(out[312], out[776], _051998_);
  xor g_110666_(out[305], out[769], _051999_);
  xor g_110667_(out[317], out[781], _052000_);
  xor g_110668_(out[313], out[777], _052001_);
  xor g_110669_(out[308], out[772], _052002_);
  xor g_110670_(out[306], out[770], _052003_);
  and g_110671_(out[315], _049697_, _052004_);
  xor g_110672_(out[307], out[771], _052005_);
  xor g_110673_(out[310], out[774], _052006_);
  xor g_110674_(out[319], out[783], _052008_);
  xor g_110675_(out[314], out[778], _052009_);
  xor g_110676_(out[309], out[773], _052010_);
  xor g_110677_(out[304], out[768], _052011_);
  or g_110678_(_051997_, _052002_, _052012_);
  or g_110679_(_051998_, _052000_, _052013_);
  or g_110680_(_052003_, _052009_, _052014_);
  or g_110681_(_052013_, _052014_, _052015_);
  or g_110682_(_052001_, _052005_, _052016_);
  or g_110683_(_052010_, _052011_, _052017_);
  or g_110684_(_052016_, _052017_, _052019_);
  or g_110685_(_052015_, _052019_, _052020_);
  xor g_110686_(out[316], out[780], _052021_);
  or g_110687_(_051995_, _052021_, _052022_);
  or g_110688_(_051994_, _052006_, _052023_);
  or g_110689_(_052022_, _052023_, _052024_);
  or g_110690_(_051999_, _052004_, _052025_);
  or g_110691_(_052008_, _052025_, _052026_);
  or g_110692_(_052024_, _052026_, _052027_);
  or g_110693_(_052020_, _052027_, _052028_);
  or g_110694_(_052012_, _052028_, _052030_);
  xor g_110695_(out[291], out[771], _052031_);
  xor g_110696_(out[292], out[772], _052032_);
  xor g_110697_(out[302], out[782], _052033_);
  xor g_110698_(out[290], out[770], _052034_);
  xor g_110699_(out[293], out[773], _052035_);
  xor g_110700_(out[297], out[777], _052036_);
  xor g_110701_(out[296], out[776], _052037_);
  xor g_110702_(out[303], out[783], _052038_);
  xor g_110703_(out[298], out[778], _052039_);
  xor g_110704_(out[294], out[774], _052041_);
  xor g_110705_(out[288], out[768], _052042_);
  and g_110706_(_098272_, out[779], _052043_);
  and g_110707_(out[299], _049697_, _052044_);
  xor g_110708_(out[301], out[781], _052045_);
  or g_110709_(_052037_, _052045_, _052046_);
  xor g_110710_(out[289], out[769], _052047_);
  or g_110711_(_052034_, _052039_, _052048_);
  or g_110712_(_052046_, _052048_, _052049_);
  or g_110713_(_052031_, _052036_, _052050_);
  or g_110714_(_052035_, _052050_, _052052_);
  or g_110715_(_052049_, _052052_, _052053_);
  or g_110716_(_052032_, _052033_, _052054_);
  or g_110717_(_052053_, _052054_, _052055_);
  xor g_110718_(out[300], out[780], _052056_);
  or g_110719_(_052043_, _052056_, _052057_);
  xor g_110720_(out[295], out[775], _052058_);
  or g_110721_(_052041_, _052058_, _052059_);
  or g_110722_(_052057_, _052059_, _052060_);
  or g_110723_(_052044_, _052047_, _052061_);
  or g_110724_(_052038_, _052061_, _052063_);
  or g_110725_(_052060_, _052063_, _052064_);
  or g_110726_(_052042_, _052064_, _052065_);
  or g_110727_(_052055_, _052065_, _052066_);
  not g_110728_(_052066_, _052067_);
  xor g_110729_(out[279], out[775], _052068_);
  and g_110730_(_098261_, out[779], _052069_);
  xor g_110731_(out[286], out[782], _052070_);
  xor g_110732_(out[280], out[776], _052071_);
  xor g_110733_(out[273], out[769], _052072_);
  xor g_110734_(out[285], out[781], _052074_);
  xor g_110735_(out[281], out[777], _052075_);
  xor g_110736_(out[276], out[772], _052076_);
  xor g_110737_(out[274], out[770], _052077_);
  and g_110738_(out[283], _049697_, _052078_);
  xor g_110739_(out[275], out[771], _052079_);
  xor g_110740_(out[278], out[774], _052080_);
  xor g_110741_(out[287], out[783], _052081_);
  xor g_110742_(out[282], out[778], _052082_);
  xor g_110743_(out[277], out[773], _052083_);
  xor g_110744_(out[272], out[768], _052085_);
  or g_110745_(_052070_, _052076_, _052086_);
  or g_110746_(_052071_, _052074_, _052087_);
  or g_110747_(_052077_, _052082_, _052088_);
  or g_110748_(_052087_, _052088_, _052089_);
  or g_110749_(_052075_, _052079_, _052090_);
  or g_110750_(_052083_, _052085_, _052091_);
  or g_110751_(_052090_, _052091_, _052092_);
  or g_110752_(_052089_, _052092_, _052093_);
  xor g_110753_(out[284], out[780], _052094_);
  or g_110754_(_052069_, _052094_, _052096_);
  or g_110755_(_052068_, _052080_, _052097_);
  or g_110756_(_052096_, _052097_, _052098_);
  or g_110757_(_052072_, _052078_, _052099_);
  or g_110758_(_052081_, _052099_, _052100_);
  or g_110759_(_052098_, _052100_, _052101_);
  or g_110760_(_052093_, _052101_, _052102_);
  or g_110761_(_052086_, _052102_, _052103_);
  not g_110762_(_052103_, _052104_);
  xor g_110763_(out[257], out[769], _052105_);
  and g_110764_(out[267], _049697_, _052107_);
  xor g_110765_(out[265], out[777], _052108_);
  xor g_110766_(out[256], out[768], _052109_);
  xor g_110767_(out[270], out[782], _052110_);
  xor g_110768_(out[260], out[772], _052111_);
  or g_110769_(_052110_, _052111_, _052112_);
  xor g_110770_(out[269], out[781], _052113_);
  xor g_110771_(out[259], out[771], _052114_);
  and g_110772_(_098250_, out[779], _052115_);
  xor g_110773_(out[262], out[774], _052116_);
  xor g_110774_(out[266], out[778], _052118_);
  xor g_110775_(out[261], out[773], _052119_);
  xor g_110776_(out[271], out[783], _052120_);
  xor g_110777_(out[264], out[776], _052121_);
  or g_110778_(_052113_, _052121_, _052122_);
  xor g_110779_(out[258], out[770], _052123_);
  or g_110780_(_052118_, _052123_, _052124_);
  or g_110781_(_052122_, _052124_, _052125_);
  or g_110782_(_052108_, _052114_, _052126_);
  or g_110783_(_052119_, _052126_, _052127_);
  or g_110784_(_052125_, _052127_, _052129_);
  or g_110785_(_052112_, _052129_, _052130_);
  xor g_110786_(out[268], out[780], _052131_);
  or g_110787_(_052115_, _052131_, _052132_);
  xor g_110788_(out[263], out[775], _052133_);
  or g_110789_(_052116_, _052133_, _052134_);
  or g_110790_(_052132_, _052134_, _052135_);
  or g_110791_(_052105_, _052107_, _052136_);
  or g_110792_(_052120_, _052136_, _052137_);
  or g_110793_(_052135_, _052137_, _052138_);
  or g_110794_(_052109_, _052138_, _052140_);
  or g_110795_(_052130_, _052140_, _052141_);
  xor g_110796_(out[247], out[775], _052142_);
  and g_110797_(_098239_, out[779], _052143_);
  xor g_110798_(out[254], out[782], _052144_);
  xor g_110799_(out[248], out[776], _052145_);
  xor g_110800_(out[241], out[769], _052146_);
  xor g_110801_(out[253], out[781], _052147_);
  xor g_110802_(out[249], out[777], _052148_);
  xor g_110803_(out[244], out[772], _052149_);
  xor g_110804_(out[242], out[770], _052151_);
  and g_110805_(out[251], _049697_, _052152_);
  xor g_110806_(out[243], out[771], _052153_);
  xor g_110807_(out[246], out[774], _052154_);
  xor g_110808_(out[255], out[783], _052155_);
  xor g_110809_(out[250], out[778], _052156_);
  xor g_110810_(out[245], out[773], _052157_);
  xor g_110811_(out[240], out[768], _052158_);
  or g_110812_(_052144_, _052149_, _052159_);
  or g_110813_(_052145_, _052147_, _052160_);
  or g_110814_(_052151_, _052156_, _052162_);
  or g_110815_(_052160_, _052162_, _052163_);
  or g_110816_(_052148_, _052153_, _052164_);
  or g_110817_(_052157_, _052158_, _052165_);
  or g_110818_(_052164_, _052165_, _052166_);
  or g_110819_(_052163_, _052166_, _052167_);
  xor g_110820_(out[252], out[780], _052168_);
  or g_110821_(_052143_, _052168_, _052169_);
  or g_110822_(_052142_, _052154_, _052170_);
  or g_110823_(_052169_, _052170_, _052171_);
  or g_110824_(_052146_, _052152_, _052173_);
  or g_110825_(_052155_, _052173_, _052174_);
  or g_110826_(_052171_, _052174_, _052175_);
  or g_110827_(_052167_, _052175_, _052176_);
  or g_110828_(_052159_, _052176_, _052177_);
  xor g_110829_(out[232], out[776], _052178_);
  xor g_110830_(out[229], out[773], _052179_);
  xor g_110831_(out[227], out[771], _052180_);
  xor g_110832_(out[238], out[782], _052181_);
  xor g_110833_(out[237], out[781], _052182_);
  xor g_110834_(out[226], out[770], _052184_);
  xor g_110835_(out[233], out[777], _052185_);
  xor g_110836_(out[230], out[774], _052186_);
  xor g_110837_(out[239], out[783], _052187_);
  xor g_110838_(out[234], out[778], _052188_);
  xor g_110839_(out[228], out[772], _052189_);
  xor g_110840_(out[224], out[768], _052190_);
  and g_110841_(_098228_, out[779], _052191_);
  and g_110842_(out[235], _049697_, _052192_);
  or g_110843_(_052178_, _052182_, _052193_);
  xor g_110844_(out[225], out[769], _052195_);
  or g_110845_(_052184_, _052188_, _052196_);
  or g_110846_(_052193_, _052196_, _052197_);
  or g_110847_(_052180_, _052185_, _052198_);
  or g_110848_(_052179_, _052198_, _052199_);
  or g_110849_(_052197_, _052199_, _052200_);
  or g_110850_(_052181_, _052189_, _052201_);
  or g_110851_(_052200_, _052201_, _052202_);
  xor g_110852_(out[236], out[780], _052203_);
  or g_110853_(_052191_, _052203_, _052204_);
  xor g_110854_(out[231], out[775], _052206_);
  or g_110855_(_052186_, _052206_, _052207_);
  or g_110856_(_052204_, _052207_, _052208_);
  or g_110857_(_052192_, _052195_, _052209_);
  or g_110858_(_052187_, _052209_, _052210_);
  or g_110859_(_052208_, _052210_, _052211_);
  or g_110860_(_052190_, _052211_, _052212_);
  or g_110861_(_052202_, _052212_, _052213_);
  not g_110862_(_052213_, _052214_);
  xor g_110863_(out[215], out[775], _052215_);
  and g_110864_(_098217_, out[779], _052217_);
  xor g_110865_(out[222], out[782], _052218_);
  xor g_110866_(out[216], out[776], _052219_);
  xor g_110867_(out[209], out[769], _052220_);
  xor g_110868_(out[221], out[781], _052221_);
  xor g_110869_(out[217], out[777], _052222_);
  xor g_110870_(out[212], out[772], _052223_);
  xor g_110871_(out[210], out[770], _052224_);
  and g_110872_(out[219], _049697_, _052225_);
  xor g_110873_(out[211], out[771], _052226_);
  xor g_110874_(out[214], out[774], _052228_);
  xor g_110875_(out[223], out[783], _052229_);
  xor g_110876_(out[218], out[778], _052230_);
  xor g_110877_(out[213], out[773], _052231_);
  xor g_110878_(out[208], out[768], _052232_);
  or g_110879_(_052218_, _052223_, _052233_);
  or g_110880_(_052219_, _052221_, _052234_);
  or g_110881_(_052224_, _052230_, _052235_);
  or g_110882_(_052234_, _052235_, _052236_);
  or g_110883_(_052222_, _052226_, _052237_);
  or g_110884_(_052231_, _052232_, _052239_);
  or g_110885_(_052237_, _052239_, _052240_);
  or g_110886_(_052236_, _052240_, _052241_);
  xor g_110887_(out[220], out[780], _052242_);
  or g_110888_(_052217_, _052242_, _052243_);
  or g_110889_(_052215_, _052228_, _052244_);
  or g_110890_(_052243_, _052244_, _052245_);
  or g_110891_(_052220_, _052225_, _052246_);
  or g_110892_(_052229_, _052246_, _052247_);
  or g_110893_(_052245_, _052247_, _052248_);
  or g_110894_(_052241_, _052248_, _052250_);
  or g_110895_(_052233_, _052250_, _052251_);
  xor g_110896_(out[204], out[780], _052252_);
  and g_110897_(_098206_, out[779], _052253_);
  xor g_110898_(out[205], out[781], _052254_);
  xor g_110899_(out[198], out[774], _052255_);
  xor g_110900_(out[200], out[776], _052256_);
  xor g_110901_(out[201], out[777], _052257_);
  xor g_110902_(out[206], out[782], _052258_);
  xor g_110903_(out[196], out[772], _052259_);
  or g_110904_(_052258_, _052259_, _052261_);
  xor g_110905_(out[197], out[773], _052262_);
  xor g_110906_(out[193], out[769], _052263_);
  and g_110907_(out[203], _049697_, _052264_);
  xor g_110908_(out[207], out[783], _052265_);
  xor g_110909_(out[202], out[778], _052266_);
  xor g_110910_(out[192], out[768], _052267_);
  xor g_110911_(out[194], out[770], _052268_);
  xor g_110912_(out[195], out[771], _052269_);
  or g_110913_(_052254_, _052256_, _052270_);
  or g_110914_(_052266_, _052268_, _052272_);
  or g_110915_(_052270_, _052272_, _052273_);
  or g_110916_(_052257_, _052269_, _052274_);
  or g_110917_(_052262_, _052267_, _052275_);
  or g_110918_(_052274_, _052275_, _052276_);
  or g_110919_(_052273_, _052276_, _052277_);
  or g_110920_(_052252_, _052253_, _052278_);
  xor g_110921_(out[199], out[775], _052279_);
  or g_110922_(_052255_, _052279_, _052280_);
  or g_110923_(_052278_, _052280_, _052281_);
  or g_110924_(_052263_, _052264_, _052283_);
  or g_110925_(_052265_, _052283_, _052284_);
  or g_110926_(_052281_, _052284_, _052285_);
  or g_110927_(_052277_, _052285_, _052286_);
  or g_110928_(_052261_, _052286_, _052287_);
  xor g_110929_(out[183], out[775], _052288_);
  and g_110930_(_098195_, out[779], _052289_);
  xor g_110931_(out[190], out[782], _052290_);
  xor g_110932_(out[184], out[776], _052291_);
  xor g_110933_(out[177], out[769], _052292_);
  xor g_110934_(out[189], out[781], _052294_);
  xor g_110935_(out[185], out[777], _052295_);
  xor g_110936_(out[180], out[772], _052296_);
  xor g_110937_(out[178], out[770], _052297_);
  and g_110938_(out[187], _049697_, _052298_);
  xor g_110939_(out[179], out[771], _052299_);
  xor g_110940_(out[182], out[774], _052300_);
  xor g_110941_(out[191], out[783], _052301_);
  xor g_110942_(out[186], out[778], _052302_);
  xor g_110943_(out[181], out[773], _052303_);
  xor g_110944_(out[176], out[768], _052305_);
  or g_110945_(_052290_, _052296_, _052306_);
  or g_110946_(_052291_, _052294_, _052307_);
  or g_110947_(_052297_, _052302_, _052308_);
  or g_110948_(_052307_, _052308_, _052309_);
  or g_110949_(_052295_, _052299_, _052310_);
  or g_110950_(_052303_, _052305_, _052311_);
  or g_110951_(_052310_, _052311_, _052312_);
  or g_110952_(_052309_, _052312_, _052313_);
  xor g_110953_(out[188], out[780], _052314_);
  or g_110954_(_052289_, _052314_, _052316_);
  or g_110955_(_052288_, _052300_, _052317_);
  or g_110956_(_052316_, _052317_, _052318_);
  or g_110957_(_052292_, _052298_, _052319_);
  or g_110958_(_052301_, _052319_, _052320_);
  or g_110959_(_052318_, _052320_, _052321_);
  or g_110960_(_052313_, _052321_, _052322_);
  or g_110961_(_052306_, _052322_, _052323_);
  not g_110962_(_052323_, _052324_);
  xor g_110963_(out[161], out[769], _052325_);
  and g_110964_(out[171], _049697_, _052327_);
  xor g_110965_(out[169], out[777], _052328_);
  xor g_110966_(out[160], out[768], _052329_);
  xor g_110967_(out[174], out[782], _052330_);
  xor g_110968_(out[164], out[772], _052331_);
  or g_110969_(_052330_, _052331_, _052332_);
  xor g_110970_(out[173], out[781], _052333_);
  xor g_110971_(out[163], out[771], _052334_);
  and g_110972_(_098184_, out[779], _052335_);
  xor g_110973_(out[166], out[774], _052336_);
  xor g_110974_(out[170], out[778], _052338_);
  xor g_110975_(out[165], out[773], _052339_);
  xor g_110976_(out[175], out[783], _052340_);
  xor g_110977_(out[168], out[776], _052341_);
  or g_110978_(_052333_, _052341_, _052342_);
  xor g_110979_(out[162], out[770], _052343_);
  or g_110980_(_052338_, _052343_, _052344_);
  or g_110981_(_052342_, _052344_, _052345_);
  or g_110982_(_052328_, _052334_, _052346_);
  or g_110983_(_052339_, _052346_, _052347_);
  or g_110984_(_052345_, _052347_, _052349_);
  or g_110985_(_052332_, _052349_, _052350_);
  xor g_110986_(out[172], out[780], _052351_);
  or g_110987_(_052335_, _052351_, _052352_);
  xor g_110988_(out[167], out[775], _052353_);
  or g_110989_(_052336_, _052353_, _052354_);
  or g_110990_(_052352_, _052354_, _052355_);
  or g_110991_(_052325_, _052327_, _052356_);
  or g_110992_(_052340_, _052356_, _052357_);
  or g_110993_(_052355_, _052357_, _052358_);
  or g_110994_(_052329_, _052358_, _052360_);
  or g_110995_(_052350_, _052360_, _052361_);
  xor g_110996_(out[151], out[775], _052362_);
  and g_110997_(_098173_, out[779], _052363_);
  xor g_110998_(out[158], out[782], _052364_);
  xor g_110999_(out[152], out[776], _052365_);
  xor g_111000_(out[145], out[769], _052366_);
  xor g_111001_(out[157], out[781], _052367_);
  xor g_111002_(out[153], out[777], _052368_);
  xor g_111003_(out[148], out[772], _052369_);
  xor g_111004_(out[146], out[770], _052371_);
  and g_111005_(out[155], _049697_, _052372_);
  xor g_111006_(out[147], out[771], _052373_);
  xor g_111007_(out[150], out[774], _052374_);
  xor g_111008_(out[159], out[783], _052375_);
  xor g_111009_(out[154], out[778], _052376_);
  xor g_111010_(out[149], out[773], _052377_);
  xor g_111011_(out[144], out[768], _052378_);
  or g_111012_(_052364_, _052369_, _052379_);
  or g_111013_(_052365_, _052367_, _052380_);
  or g_111014_(_052371_, _052376_, _052382_);
  or g_111015_(_052380_, _052382_, _052383_);
  or g_111016_(_052368_, _052373_, _052384_);
  or g_111017_(_052377_, _052378_, _052385_);
  or g_111018_(_052384_, _052385_, _052386_);
  or g_111019_(_052383_, _052386_, _052387_);
  xor g_111020_(out[156], out[780], _052388_);
  or g_111021_(_052363_, _052388_, _052389_);
  or g_111022_(_052362_, _052374_, _052390_);
  or g_111023_(_052389_, _052390_, _052391_);
  or g_111024_(_052366_, _052372_, _052393_);
  or g_111025_(_052375_, _052393_, _052394_);
  or g_111026_(_052391_, _052394_, _052395_);
  or g_111027_(_052387_, _052395_, _052396_);
  or g_111028_(_052379_, _052396_, _052397_);
  and g_111029_(out[139], _049697_, _052398_);
  xor g_111030_(out[132], out[772], _052399_);
  xor g_111031_(out[142], out[782], _052400_);
  or g_111032_(_052399_, _052400_, _052401_);
  xor g_111033_(out[141], out[781], _052402_);
  xor g_111034_(out[131], out[771], _052404_);
  xor g_111035_(out[128], out[768], _052405_);
  and g_111036_(_098162_, out[779], _052406_);
  xor g_111037_(out[138], out[778], _052407_);
  xor g_111038_(out[143], out[783], _052408_);
  xor g_111039_(out[134], out[774], _052409_);
  xor g_111040_(out[133], out[773], _052410_);
  xor g_111041_(out[136], out[776], _052411_);
  or g_111042_(_052402_, _052411_, _052412_);
  xor g_111043_(out[130], out[770], _052413_);
  xor g_111044_(out[137], out[777], _052415_);
  xor g_111045_(out[129], out[769], _052416_);
  or g_111046_(_052407_, _052413_, _052417_);
  or g_111047_(_052412_, _052417_, _052418_);
  or g_111048_(_052404_, _052415_, _052419_);
  or g_111049_(_052410_, _052419_, _052420_);
  or g_111050_(_052418_, _052420_, _052421_);
  or g_111051_(_052401_, _052421_, _052422_);
  xor g_111052_(out[140], out[780], _052423_);
  or g_111053_(_052406_, _052423_, _052424_);
  xor g_111054_(out[135], out[775], _052426_);
  or g_111055_(_052409_, _052426_, _052427_);
  or g_111056_(_052424_, _052427_, _052428_);
  or g_111057_(_052398_, _052416_, _052429_);
  or g_111058_(_052408_, _052429_, _052430_);
  or g_111059_(_052428_, _052430_, _052431_);
  or g_111060_(_052405_, _052431_, _052432_);
  or g_111061_(_052422_, _052432_, _052433_);
  xor g_111062_(out[119], out[775], _052434_);
  and g_111063_(_098151_, out[779], _052435_);
  xor g_111064_(out[126], out[782], _052437_);
  xor g_111065_(out[120], out[776], _052438_);
  xor g_111066_(out[113], out[769], _052439_);
  xor g_111067_(out[125], out[781], _052440_);
  xor g_111068_(out[121], out[777], _052441_);
  xor g_111069_(out[116], out[772], _052442_);
  xor g_111070_(out[114], out[770], _052443_);
  and g_111071_(out[123], _049697_, _052444_);
  xor g_111072_(out[115], out[771], _052445_);
  xor g_111073_(out[118], out[774], _052446_);
  xor g_111074_(out[127], out[783], _052448_);
  xor g_111075_(out[122], out[778], _052449_);
  xor g_111076_(out[117], out[773], _052450_);
  xor g_111077_(out[112], out[768], _052451_);
  or g_111078_(_052437_, _052442_, _052452_);
  or g_111079_(_052438_, _052440_, _052453_);
  or g_111080_(_052443_, _052449_, _052454_);
  or g_111081_(_052453_, _052454_, _052455_);
  or g_111082_(_052441_, _052445_, _052456_);
  or g_111083_(_052450_, _052451_, _052457_);
  or g_111084_(_052456_, _052457_, _052459_);
  or g_111085_(_052455_, _052459_, _052460_);
  xor g_111086_(out[124], out[780], _052461_);
  or g_111087_(_052435_, _052461_, _052462_);
  or g_111088_(_052434_, _052446_, _052463_);
  or g_111089_(_052462_, _052463_, _052464_);
  or g_111090_(_052439_, _052444_, _052465_);
  or g_111091_(_052448_, _052465_, _052466_);
  or g_111092_(_052464_, _052466_, _052467_);
  or g_111093_(_052460_, _052467_, _052468_);
  or g_111094_(_052452_, _052468_, _052470_);
  xor g_111095_(out[100], out[772], _052471_);
  xor g_111096_(out[108], out[780], _052472_);
  and g_111097_(_098140_, out[779], _052473_);
  xor g_111098_(out[106], out[778], _052474_);
  xor g_111099_(out[102], out[774], _052475_);
  xor g_111100_(out[101], out[773], _052476_);
  xor g_111101_(out[99], out[771], _052477_);
  xor g_111102_(out[109], out[781], _052478_);
  xor g_111103_(out[110], out[782], _052479_);
  xor g_111104_(out[97], out[769], _052481_);
  xor g_111105_(out[98], out[770], _052482_);
  and g_111106_(out[107], _049697_, _052483_);
  xor g_111107_(out[96], out[768], _052484_);
  xor g_111108_(out[111], out[783], _052485_);
  xor g_111109_(out[104], out[776], _052486_);
  or g_111110_(_052478_, _052486_, _052487_);
  xor g_111111_(out[105], out[777], _052488_);
  or g_111112_(_052474_, _052482_, _052489_);
  or g_111113_(_052487_, _052489_, _052490_);
  or g_111114_(_052477_, _052488_, _052492_);
  or g_111115_(_052476_, _052492_, _052493_);
  or g_111116_(_052490_, _052493_, _052494_);
  or g_111117_(_052471_, _052479_, _052495_);
  or g_111118_(_052494_, _052495_, _052496_);
  or g_111119_(_052472_, _052473_, _052497_);
  xor g_111120_(out[103], out[775], _052498_);
  or g_111121_(_052475_, _052498_, _052499_);
  or g_111122_(_052497_, _052499_, _052500_);
  or g_111123_(_052481_, _052483_, _052501_);
  or g_111124_(_052485_, _052501_, _052503_);
  or g_111125_(_052500_, _052503_, _052504_);
  or g_111126_(_052484_, _052504_, _052505_);
  or g_111127_(_052496_, _052505_, _052506_);
  not g_111128_(_052506_, _052507_);
  xor g_111129_(out[87], out[775], _052508_);
  and g_111130_(_098129_, out[779], _052509_);
  xor g_111131_(out[94], out[782], _052510_);
  xor g_111132_(out[88], out[776], _052511_);
  xor g_111133_(out[81], out[769], _052512_);
  xor g_111134_(out[93], out[781], _052514_);
  xor g_111135_(out[89], out[777], _052515_);
  xor g_111136_(out[84], out[772], _052516_);
  xor g_111137_(out[82], out[770], _052517_);
  and g_111138_(out[91], _049697_, _052518_);
  xor g_111139_(out[83], out[771], _052519_);
  xor g_111140_(out[86], out[774], _052520_);
  xor g_111141_(out[95], out[783], _052521_);
  xor g_111142_(out[90], out[778], _052522_);
  xor g_111143_(out[85], out[773], _052523_);
  xor g_111144_(out[80], out[768], _052525_);
  or g_111145_(_052510_, _052516_, _052526_);
  or g_111146_(_052511_, _052514_, _052527_);
  or g_111147_(_052517_, _052522_, _052528_);
  or g_111148_(_052527_, _052528_, _052529_);
  or g_111149_(_052515_, _052519_, _052530_);
  or g_111150_(_052523_, _052525_, _052531_);
  or g_111151_(_052530_, _052531_, _052532_);
  or g_111152_(_052529_, _052532_, _052533_);
  xor g_111153_(out[92], out[780], _052534_);
  or g_111154_(_052509_, _052534_, _052536_);
  or g_111155_(_052508_, _052520_, _052537_);
  or g_111156_(_052536_, _052537_, _052538_);
  or g_111157_(_052512_, _052518_, _052539_);
  or g_111158_(_052521_, _052539_, _052540_);
  or g_111159_(_052538_, _052540_, _052541_);
  or g_111160_(_052533_, _052541_, _052542_);
  or g_111161_(_052526_, _052542_, _052543_);
  xor g_111162_(out[74], out[778], _052544_);
  xor g_111163_(out[66], out[770], _052545_);
  xor g_111164_(out[65], out[769], _052547_);
  and g_111165_(_098118_, out[779], _052548_);
  and g_111166_(out[75], _049697_, _052549_);
  xor g_111167_(out[77], out[781], _052550_);
  xor g_111168_(out[67], out[771], _052551_);
  xor g_111169_(out[78], out[782], _052552_);
  xor g_111170_(out[76], out[780], _052553_);
  xor g_111171_(out[72], out[776], _052554_);
  xor g_111172_(out[79], out[783], _052555_);
  xor g_111173_(out[69], out[773], _052556_);
  xor g_111174_(out[70], out[774], _052558_);
  xor g_111175_(out[64], out[768], _052559_);
  xor g_111176_(out[68], out[772], _052560_);
  or g_111177_(_052550_, _052554_, _052561_);
  xor g_111178_(out[73], out[777], _052562_);
  or g_111179_(_052544_, _052545_, _052563_);
  or g_111180_(_052561_, _052563_, _052564_);
  or g_111181_(_052551_, _052562_, _052565_);
  or g_111182_(_052556_, _052565_, _052566_);
  or g_111183_(_052564_, _052566_, _052567_);
  or g_111184_(_052552_, _052560_, _052569_);
  or g_111185_(_052567_, _052569_, _052570_);
  or g_111186_(_052548_, _052553_, _052571_);
  xor g_111187_(out[71], out[775], _052572_);
  or g_111188_(_052558_, _052572_, _052573_);
  or g_111189_(_052571_, _052573_, _052574_);
  or g_111190_(_052547_, _052549_, _052575_);
  or g_111191_(_052555_, _052575_, _052576_);
  or g_111192_(_052574_, _052576_, _052577_);
  or g_111193_(_052559_, _052577_, _052578_);
  or g_111194_(_052570_, _052578_, _052580_);
  xor g_111195_(out[55], out[775], _052581_);
  and g_111196_(_098107_, out[779], _052582_);
  xor g_111197_(out[62], out[782], _052583_);
  xor g_111198_(out[56], out[776], _052584_);
  xor g_111199_(out[49], out[769], _052585_);
  xor g_111200_(out[61], out[781], _052586_);
  xor g_111201_(out[57], out[777], _052587_);
  xor g_111202_(out[52], out[772], _052588_);
  xor g_111203_(out[50], out[770], _052589_);
  and g_111204_(out[59], _049697_, _052591_);
  xor g_111205_(out[51], out[771], _052592_);
  xor g_111206_(out[54], out[774], _052593_);
  xor g_111207_(out[63], out[783], _052594_);
  xor g_111208_(out[58], out[778], _052595_);
  xor g_111209_(out[53], out[773], _052596_);
  xor g_111210_(out[48], out[768], _052597_);
  or g_111211_(_052583_, _052588_, _052598_);
  or g_111212_(_052584_, _052586_, _052599_);
  or g_111213_(_052589_, _052595_, _052600_);
  or g_111214_(_052599_, _052600_, _052602_);
  or g_111215_(_052587_, _052592_, _052603_);
  or g_111216_(_052596_, _052597_, _052604_);
  or g_111217_(_052603_, _052604_, _052605_);
  or g_111218_(_052602_, _052605_, _052606_);
  xor g_111219_(out[60], out[780], _052607_);
  or g_111220_(_052582_, _052607_, _052608_);
  or g_111221_(_052581_, _052593_, _052609_);
  or g_111222_(_052608_, _052609_, _052610_);
  or g_111223_(_052585_, _052591_, _052611_);
  or g_111224_(_052594_, _052611_, _052613_);
  or g_111225_(_052610_, _052613_, _052614_);
  or g_111226_(_052606_, _052614_, _052615_);
  or g_111227_(_052598_, _052615_, _052616_);
  xor g_111228_(out[33], out[769], _052617_);
  and g_111229_(_098096_, out[779], _052618_);
  and g_111230_(out[43], _049697_, _052619_);
  xor g_111231_(out[40], out[776], _052620_);
  xor g_111232_(out[42], out[778], _052621_);
  xor g_111233_(out[34], out[770], _052622_);
  xor g_111234_(out[36], out[772], _052624_);
  xor g_111235_(out[45], out[781], _052625_);
  xor g_111236_(out[41], out[777], _052626_);
  xor g_111237_(out[35], out[771], _052627_);
  xor g_111238_(out[37], out[773], _052628_);
  xor g_111239_(out[46], out[782], _052629_);
  xor g_111240_(out[32], out[768], _052630_);
  xor g_111241_(out[47], out[783], _052631_);
  or g_111242_(_052620_, _052625_, _052632_);
  xor g_111243_(out[38], out[774], _052633_);
  or g_111244_(_052621_, _052622_, _052635_);
  or g_111245_(_052632_, _052635_, _052636_);
  or g_111246_(_052626_, _052627_, _052637_);
  or g_111247_(_052628_, _052637_, _052638_);
  or g_111248_(_052636_, _052638_, _052639_);
  or g_111249_(_052624_, _052629_, _052640_);
  or g_111250_(_052639_, _052640_, _052641_);
  xor g_111251_(out[44], out[780], _052642_);
  or g_111252_(_052618_, _052642_, _052643_);
  xor g_111253_(out[39], out[775], _052644_);
  or g_111254_(_052633_, _052644_, _052646_);
  or g_111255_(_052643_, _052646_, _052647_);
  or g_111256_(_052617_, _052619_, _052648_);
  or g_111257_(_052631_, _052648_, _052649_);
  or g_111258_(_052647_, _052649_, _052650_);
  or g_111259_(_052630_, _052650_, _052651_);
  or g_111260_(_052641_, _052651_, _052652_);
  xor g_111261_(out[23], out[775], _052653_);
  and g_111262_(_098063_, out[779], _052654_);
  xor g_111263_(out[30], out[782], _052655_);
  xor g_111264_(out[24], out[776], _052657_);
  xor g_111265_(out[17], out[769], _052658_);
  xor g_111266_(out[29], out[781], _052659_);
  xor g_111267_(out[25], out[777], _052660_);
  xor g_111268_(out[20], out[772], _052661_);
  xor g_111269_(out[18], out[770], _052662_);
  and g_111270_(out[27], _049697_, _052663_);
  xor g_111271_(out[19], out[771], _052664_);
  xor g_111272_(out[22], out[774], _052665_);
  xor g_111273_(out[31], out[783], _052666_);
  xor g_111274_(out[26], out[778], _052668_);
  xor g_111275_(out[21], out[773], _052669_);
  xor g_111276_(out[16], out[768], _052670_);
  or g_111277_(_052655_, _052661_, _052671_);
  or g_111278_(_052657_, _052659_, _052672_);
  or g_111279_(_052662_, _052668_, _052673_);
  or g_111280_(_052672_, _052673_, _052674_);
  or g_111281_(_052660_, _052664_, _052675_);
  or g_111282_(_052669_, _052670_, _052676_);
  or g_111283_(_052675_, _052676_, _052677_);
  or g_111284_(_052674_, _052677_, _052679_);
  xor g_111285_(out[28], out[780], _052680_);
  or g_111286_(_052654_, _052680_, _052681_);
  or g_111287_(_052653_, _052665_, _052682_);
  or g_111288_(_052681_, _052682_, _052683_);
  or g_111289_(_052658_, _052663_, _052684_);
  or g_111290_(_052666_, _052684_, _052685_);
  or g_111291_(_052683_, _052685_, _052686_);
  or g_111292_(_052679_, _052686_, _052687_);
  or g_111293_(_052671_, _052687_, _052688_);
  not g_111294_(_052688_, _052690_);
  xor g_111295_(out[1], out[769], _052691_);
  and g_111296_(out[11], _049697_, _052692_);
  xor g_111297_(out[9], out[777], _052693_);
  xor g_111298_(out[0], out[768], _052694_);
  xor g_111299_(out[14], out[782], _052695_);
  xor g_111300_(out[4], out[772], _052696_);
  or g_111301_(_052695_, _052696_, _052697_);
  xor g_111302_(out[13], out[781], _052698_);
  xor g_111303_(out[3], out[771], _052699_);
  and g_111304_(_098041_, out[779], _052701_);
  xor g_111305_(out[6], out[774], _052702_);
  xor g_111306_(out[10], out[778], _052703_);
  xor g_111307_(out[5], out[773], _052704_);
  xor g_111308_(out[15], out[783], _052705_);
  xor g_111309_(out[8], out[776], _052706_);
  or g_111310_(_052698_, _052706_, _052707_);
  xor g_111311_(out[2], out[770], _052708_);
  or g_111312_(_052703_, _052708_, _052709_);
  or g_111313_(_052707_, _052709_, _052710_);
  or g_111314_(_052693_, _052699_, _052712_);
  or g_111315_(_052704_, _052712_, _052713_);
  or g_111316_(_052710_, _052713_, _052714_);
  or g_111317_(_052697_, _052714_, _052715_);
  xor g_111318_(out[12], out[780], _052716_);
  or g_111319_(_052701_, _052716_, _052717_);
  xor g_111320_(out[7], out[775], _052718_);
  or g_111321_(_052702_, _052718_, _052719_);
  or g_111322_(_052717_, _052719_, _052720_);
  or g_111323_(_052691_, _052692_, _052721_);
  or g_111324_(_052705_, _052721_, _052723_);
  or g_111325_(_052720_, _052723_, _052724_);
  or g_111326_(_052694_, _052724_, _052725_);
  or g_111327_(_052715_, _052725_, _052726_);
  xor g_111328_(out[476], out[764], _052727_);
  and g_111329_(_049499_, out[763], _052728_);
  xor g_111330_(out[477], out[765], _052729_);
  xor g_111331_(out[470], out[758], _052730_);
  xor g_111332_(out[472], out[760], _052731_);
  xor g_111333_(out[473], out[761], _052732_);
  xor g_111334_(out[478], out[766], _052734_);
  xor g_111335_(out[468], out[756], _052735_);
  or g_111336_(_052734_, _052735_, _052736_);
  xor g_111337_(out[469], out[757], _052737_);
  xor g_111338_(out[465], out[753], _052738_);
  and g_111339_(out[475], _049686_, _052739_);
  xor g_111340_(out[479], out[767], _052740_);
  xor g_111341_(out[474], out[762], _052741_);
  xor g_111342_(out[464], out[752], _052742_);
  xor g_111343_(out[466], out[754], _052743_);
  xor g_111344_(out[467], out[755], _052745_);
  or g_111345_(_052729_, _052731_, _052746_);
  or g_111346_(_052741_, _052743_, _052747_);
  or g_111347_(_052746_, _052747_, _052748_);
  or g_111348_(_052732_, _052745_, _052749_);
  or g_111349_(_052737_, _052742_, _052750_);
  or g_111350_(_052749_, _052750_, _052751_);
  or g_111351_(_052748_, _052751_, _052752_);
  or g_111352_(_052727_, _052728_, _052753_);
  xor g_111353_(out[471], out[759], _052754_);
  or g_111354_(_052730_, _052754_, _052756_);
  or g_111355_(_052753_, _052756_, _052757_);
  or g_111356_(_052738_, _052739_, _052758_);
  or g_111357_(_052740_, _052758_, _052759_);
  or g_111358_(_052757_, _052759_, _052760_);
  or g_111359_(_052752_, _052760_, _052761_);
  or g_111360_(_052736_, _052761_, _052762_);
  xor g_111361_(out[455], out[759], _052763_);
  and g_111362_(_049477_, out[763], _052764_);
  xor g_111363_(out[462], out[766], _052765_);
  xor g_111364_(out[456], out[760], _052767_);
  xor g_111365_(out[449], out[753], _052768_);
  xor g_111366_(out[461], out[765], _052769_);
  xor g_111367_(out[457], out[761], _052770_);
  xor g_111368_(out[452], out[756], _052771_);
  xor g_111369_(out[450], out[754], _052772_);
  and g_111370_(out[459], _049686_, _052773_);
  xor g_111371_(out[451], out[755], _052774_);
  xor g_111372_(out[454], out[758], _052775_);
  xor g_111373_(out[463], out[767], _052776_);
  xor g_111374_(out[458], out[762], _052778_);
  xor g_111375_(out[453], out[757], _052779_);
  xor g_111376_(out[448], out[752], _052780_);
  or g_111377_(_052765_, _052771_, _052781_);
  or g_111378_(_052767_, _052769_, _052782_);
  or g_111379_(_052772_, _052778_, _052783_);
  or g_111380_(_052782_, _052783_, _052784_);
  or g_111381_(_052770_, _052774_, _052785_);
  or g_111382_(_052779_, _052780_, _052786_);
  or g_111383_(_052785_, _052786_, _052787_);
  or g_111384_(_052784_, _052787_, _052789_);
  xor g_111385_(out[460], out[764], _052790_);
  or g_111386_(_052764_, _052790_, _052791_);
  or g_111387_(_052763_, _052775_, _052792_);
  or g_111388_(_052791_, _052792_, _052793_);
  or g_111389_(_052768_, _052773_, _052794_);
  or g_111390_(_052776_, _052794_, _052795_);
  or g_111391_(_052793_, _052795_, _052796_);
  or g_111392_(_052789_, _052796_, _052797_);
  or g_111393_(_052781_, _052797_, _052798_);
  xor g_111394_(out[444], out[764], _052800_);
  and g_111395_(_049466_, out[763], _052801_);
  xor g_111396_(out[440], out[760], _052802_);
  xor g_111397_(out[438], out[758], _052803_);
  xor g_111398_(out[445], out[765], _052804_);
  xor g_111399_(out[446], out[766], _052805_);
  xor g_111400_(out[434], out[754], _052806_);
  xor g_111401_(out[441], out[761], _052807_);
  xor g_111402_(out[437], out[757], _052808_);
  xor g_111403_(out[433], out[753], _052809_);
  and g_111404_(out[443], _049686_, _052811_);
  or g_111405_(_052802_, _052804_, _052812_);
  xor g_111406_(out[447], out[767], _052813_);
  xor g_111407_(out[442], out[762], _052814_);
  xor g_111408_(out[436], out[756], _052815_);
  xor g_111409_(out[435], out[755], _052816_);
  xor g_111410_(out[432], out[752], _052817_);
  or g_111411_(_052806_, _052814_, _052818_);
  or g_111412_(_052812_, _052818_, _052819_);
  or g_111413_(_052807_, _052816_, _052820_);
  or g_111414_(_052808_, _052820_, _052822_);
  or g_111415_(_052819_, _052822_, _052823_);
  or g_111416_(_052805_, _052815_, _052824_);
  or g_111417_(_052823_, _052824_, _052825_);
  or g_111418_(_052800_, _052801_, _052826_);
  xor g_111419_(out[439], out[759], _052827_);
  or g_111420_(_052803_, _052827_, _052828_);
  or g_111421_(_052826_, _052828_, _052829_);
  or g_111422_(_052809_, _052811_, _052830_);
  or g_111423_(_052813_, _052830_, _052831_);
  or g_111424_(_052829_, _052831_, _052833_);
  or g_111425_(_052817_, _052833_, _052834_);
  or g_111426_(_052825_, _052834_, _052835_);
  xor g_111427_(out[423], out[759], _052836_);
  and g_111428_(_049455_, out[763], _052837_);
  xor g_111429_(out[430], out[766], _052838_);
  xor g_111430_(out[424], out[760], _052839_);
  xor g_111431_(out[417], out[753], _052840_);
  xor g_111432_(out[429], out[765], _052841_);
  xor g_111433_(out[425], out[761], _052842_);
  xor g_111434_(out[420], out[756], _052844_);
  xor g_111435_(out[418], out[754], _052845_);
  and g_111436_(out[427], _049686_, _052846_);
  xor g_111437_(out[419], out[755], _052847_);
  xor g_111438_(out[422], out[758], _052848_);
  xor g_111439_(out[431], out[767], _052849_);
  xor g_111440_(out[426], out[762], _052850_);
  xor g_111441_(out[421], out[757], _052851_);
  xor g_111442_(out[416], out[752], _052852_);
  or g_111443_(_052838_, _052844_, _052853_);
  or g_111444_(_052839_, _052841_, _052855_);
  or g_111445_(_052845_, _052850_, _052856_);
  or g_111446_(_052855_, _052856_, _052857_);
  or g_111447_(_052842_, _052847_, _052858_);
  or g_111448_(_052851_, _052852_, _052859_);
  or g_111449_(_052858_, _052859_, _052860_);
  or g_111450_(_052857_, _052860_, _052861_);
  xor g_111451_(out[428], out[764], _052862_);
  or g_111452_(_052837_, _052862_, _052863_);
  or g_111453_(_052836_, _052848_, _052864_);
  or g_111454_(_052863_, _052864_, _052866_);
  or g_111455_(_052840_, _052846_, _052867_);
  or g_111456_(_052849_, _052867_, _052868_);
  or g_111457_(_052866_, _052868_, _052869_);
  or g_111458_(_052861_, _052869_, _052870_);
  or g_111459_(_052853_, _052870_, _052871_);
  xor g_111460_(out[404], out[756], _052872_);
  xor g_111461_(out[412], out[764], _052873_);
  and g_111462_(_049444_, out[763], _052874_);
  xor g_111463_(out[410], out[762], _052875_);
  xor g_111464_(out[406], out[758], _052877_);
  xor g_111465_(out[405], out[757], _052878_);
  xor g_111466_(out[403], out[755], _052879_);
  xor g_111467_(out[413], out[765], _052880_);
  xor g_111468_(out[414], out[766], _052881_);
  xor g_111469_(out[401], out[753], _052882_);
  xor g_111470_(out[402], out[754], _052883_);
  and g_111471_(out[411], _049686_, _052884_);
  xor g_111472_(out[400], out[752], _052885_);
  xor g_111473_(out[415], out[767], _052886_);
  xor g_111474_(out[408], out[760], _052888_);
  or g_111475_(_052880_, _052888_, _052889_);
  xor g_111476_(out[409], out[761], _052890_);
  or g_111477_(_052875_, _052883_, _052891_);
  or g_111478_(_052889_, _052891_, _052892_);
  or g_111479_(_052879_, _052890_, _052893_);
  or g_111480_(_052878_, _052893_, _052894_);
  or g_111481_(_052892_, _052894_, _052895_);
  or g_111482_(_052872_, _052881_, _052896_);
  or g_111483_(_052895_, _052896_, _052897_);
  or g_111484_(_052873_, _052874_, _052899_);
  xor g_111485_(out[407], out[759], _052900_);
  or g_111486_(_052877_, _052900_, _052901_);
  or g_111487_(_052899_, _052901_, _052902_);
  or g_111488_(_052882_, _052884_, _052903_);
  or g_111489_(_052886_, _052903_, _052904_);
  or g_111490_(_052902_, _052904_, _052905_);
  or g_111491_(_052885_, _052905_, _052906_);
  or g_111492_(_052897_, _052906_, _052907_);
  xor g_111493_(out[391], out[759], _052908_);
  and g_111494_(_049433_, out[763], _052910_);
  xor g_111495_(out[398], out[766], _052911_);
  xor g_111496_(out[392], out[760], _052912_);
  xor g_111497_(out[385], out[753], _052913_);
  xor g_111498_(out[397], out[765], _052914_);
  xor g_111499_(out[393], out[761], _052915_);
  xor g_111500_(out[388], out[756], _052916_);
  xor g_111501_(out[386], out[754], _052917_);
  and g_111502_(out[395], _049686_, _052918_);
  xor g_111503_(out[387], out[755], _052919_);
  xor g_111504_(out[390], out[758], _052921_);
  xor g_111505_(out[399], out[767], _052922_);
  xor g_111506_(out[394], out[762], _052923_);
  xor g_111507_(out[389], out[757], _052924_);
  xor g_111508_(out[384], out[752], _052925_);
  or g_111509_(_052911_, _052916_, _052926_);
  or g_111510_(_052912_, _052914_, _052927_);
  or g_111511_(_052917_, _052923_, _052928_);
  or g_111512_(_052927_, _052928_, _052929_);
  or g_111513_(_052915_, _052919_, _052930_);
  or g_111514_(_052924_, _052925_, _052932_);
  or g_111515_(_052930_, _052932_, _052933_);
  or g_111516_(_052929_, _052933_, _052934_);
  xor g_111517_(out[396], out[764], _052935_);
  or g_111518_(_052910_, _052935_, _052936_);
  or g_111519_(_052908_, _052921_, _052937_);
  or g_111520_(_052936_, _052937_, _052938_);
  or g_111521_(_052913_, _052918_, _052939_);
  or g_111522_(_052922_, _052939_, _052940_);
  or g_111523_(_052938_, _052940_, _052941_);
  or g_111524_(_052934_, _052941_, _052943_);
  or g_111525_(_052926_, _052943_, _052944_);
  xor g_111526_(out[371], out[755], _052945_);
  xor g_111527_(out[372], out[756], _052946_);
  xor g_111528_(out[382], out[766], _052947_);
  xor g_111529_(out[370], out[754], _052948_);
  xor g_111530_(out[373], out[757], _052949_);
  xor g_111531_(out[377], out[761], _052950_);
  xor g_111532_(out[376], out[760], _052951_);
  xor g_111533_(out[383], out[767], _052952_);
  xor g_111534_(out[378], out[762], _052954_);
  xor g_111535_(out[374], out[758], _052955_);
  xor g_111536_(out[368], out[752], _052956_);
  and g_111537_(_049422_, out[763], _052957_);
  and g_111538_(out[379], _049686_, _052958_);
  xor g_111539_(out[381], out[765], _052959_);
  or g_111540_(_052951_, _052959_, _052960_);
  xor g_111541_(out[369], out[753], _052961_);
  or g_111542_(_052948_, _052954_, _052962_);
  or g_111543_(_052960_, _052962_, _052963_);
  or g_111544_(_052945_, _052950_, _052965_);
  or g_111545_(_052949_, _052965_, _052966_);
  or g_111546_(_052963_, _052966_, _052967_);
  or g_111547_(_052946_, _052947_, _052968_);
  or g_111548_(_052967_, _052968_, _052969_);
  xor g_111549_(out[380], out[764], _052970_);
  or g_111550_(_052957_, _052970_, _052971_);
  xor g_111551_(out[375], out[759], _052972_);
  or g_111552_(_052955_, _052972_, _052973_);
  or g_111553_(_052971_, _052973_, _052974_);
  or g_111554_(_052958_, _052961_, _052976_);
  or g_111555_(_052952_, _052976_, _052977_);
  or g_111556_(_052974_, _052977_, _052978_);
  or g_111557_(_052956_, _052978_, _052979_);
  or g_111558_(_052969_, _052979_, _052980_);
  xor g_111559_(out[359], out[759], _052981_);
  and g_111560_(_049411_, out[763], _052982_);
  xor g_111561_(out[366], out[766], _052983_);
  xor g_111562_(out[360], out[760], _052984_);
  xor g_111563_(out[353], out[753], _052985_);
  xor g_111564_(out[365], out[765], _052987_);
  xor g_111565_(out[361], out[761], _052988_);
  xor g_111566_(out[356], out[756], _052989_);
  xor g_111567_(out[354], out[754], _052990_);
  and g_111568_(out[363], _049686_, _052991_);
  xor g_111569_(out[355], out[755], _052992_);
  xor g_111570_(out[358], out[758], _052993_);
  xor g_111571_(out[367], out[767], _052994_);
  xor g_111572_(out[362], out[762], _052995_);
  xor g_111573_(out[357], out[757], _052996_);
  xor g_111574_(out[352], out[752], _052998_);
  or g_111575_(_052983_, _052989_, _052999_);
  or g_111576_(_052984_, _052987_, _053000_);
  or g_111577_(_052990_, _052995_, _053001_);
  or g_111578_(_053000_, _053001_, _053002_);
  or g_111579_(_052988_, _052992_, _053003_);
  or g_111580_(_052996_, _052998_, _053004_);
  or g_111581_(_053003_, _053004_, _053005_);
  or g_111582_(_053002_, _053005_, _053006_);
  xor g_111583_(out[364], out[764], _053007_);
  or g_111584_(_052982_, _053007_, _053009_);
  or g_111585_(_052981_, _052993_, _053010_);
  or g_111586_(_053009_, _053010_, _053011_);
  or g_111587_(_052985_, _052991_, _053012_);
  or g_111588_(_052994_, _053012_, _053013_);
  or g_111589_(_053011_, _053013_, _053014_);
  or g_111590_(_053006_, _053014_, _053015_);
  or g_111591_(_052999_, _053015_, _053016_);
  xor g_111592_(out[337], out[753], _053017_);
  and g_111593_(out[347], _049686_, _053018_);
  xor g_111594_(out[345], out[761], _053020_);
  xor g_111595_(out[336], out[752], _053021_);
  xor g_111596_(out[350], out[766], _053022_);
  xor g_111597_(out[340], out[756], _053023_);
  or g_111598_(_053022_, _053023_, _053024_);
  xor g_111599_(out[349], out[765], _053025_);
  xor g_111600_(out[339], out[755], _053026_);
  and g_111601_(_049400_, out[763], _053027_);
  xor g_111602_(out[342], out[758], _053028_);
  xor g_111603_(out[346], out[762], _053029_);
  xor g_111604_(out[341], out[757], _053031_);
  xor g_111605_(out[351], out[767], _053032_);
  xor g_111606_(out[344], out[760], _053033_);
  or g_111607_(_053025_, _053033_, _053034_);
  xor g_111608_(out[338], out[754], _053035_);
  or g_111609_(_053029_, _053035_, _053036_);
  or g_111610_(_053034_, _053036_, _053037_);
  or g_111611_(_053020_, _053026_, _053038_);
  or g_111612_(_053031_, _053038_, _053039_);
  or g_111613_(_053037_, _053039_, _053040_);
  or g_111614_(_053024_, _053040_, _053042_);
  xor g_111615_(out[348], out[764], _053043_);
  or g_111616_(_053027_, _053043_, _053044_);
  xor g_111617_(out[343], out[759], _053045_);
  or g_111618_(_053028_, _053045_, _053046_);
  or g_111619_(_053044_, _053046_, _053047_);
  or g_111620_(_053017_, _053018_, _053048_);
  or g_111621_(_053032_, _053048_, _053049_);
  or g_111622_(_053047_, _053049_, _053050_);
  or g_111623_(_053021_, _053050_, _053051_);
  or g_111624_(_053042_, _053051_, _053053_);
  xor g_111625_(out[327], out[759], _053054_);
  and g_111626_(_098294_, out[763], _053055_);
  xor g_111627_(out[334], out[766], _053056_);
  xor g_111628_(out[328], out[760], _053057_);
  xor g_111629_(out[321], out[753], _053058_);
  xor g_111630_(out[333], out[765], _053059_);
  xor g_111631_(out[329], out[761], _053060_);
  xor g_111632_(out[324], out[756], _053061_);
  xor g_111633_(out[322], out[754], _053062_);
  and g_111634_(out[331], _049686_, _053064_);
  xor g_111635_(out[323], out[755], _053065_);
  xor g_111636_(out[326], out[758], _053066_);
  xor g_111637_(out[335], out[767], _053067_);
  xor g_111638_(out[330], out[762], _053068_);
  xor g_111639_(out[325], out[757], _053069_);
  xor g_111640_(out[320], out[752], _053070_);
  or g_111641_(_053056_, _053061_, _053071_);
  or g_111642_(_053057_, _053059_, _053072_);
  or g_111643_(_053062_, _053068_, _053073_);
  or g_111644_(_053072_, _053073_, _053075_);
  or g_111645_(_053060_, _053065_, _053076_);
  or g_111646_(_053069_, _053070_, _053077_);
  or g_111647_(_053076_, _053077_, _053078_);
  or g_111648_(_053075_, _053078_, _053079_);
  xor g_111649_(out[332], out[764], _053080_);
  or g_111650_(_053055_, _053080_, _053081_);
  or g_111651_(_053054_, _053066_, _053082_);
  or g_111652_(_053081_, _053082_, _053083_);
  or g_111653_(_053058_, _053064_, _053084_);
  or g_111654_(_053067_, _053084_, _053086_);
  or g_111655_(_053083_, _053086_, _053087_);
  or g_111656_(_053079_, _053087_, _053088_);
  or g_111657_(_053071_, _053088_, _053089_);
  not g_111658_(_053089_, _053090_);
  xor g_111659_(out[305], out[753], _053091_);
  and g_111660_(out[315], _049686_, _053092_);
  xor g_111661_(out[318], out[766], _053093_);
  xor g_111662_(out[307], out[755], _053094_);
  xor g_111663_(out[308], out[756], _053095_);
  xor g_111664_(out[306], out[754], _053097_);
  xor g_111665_(out[313], out[761], _053098_);
  xor g_111666_(out[304], out[752], _053099_);
  and g_111667_(_098283_, out[763], _053100_);
  xor g_111668_(out[310], out[758], _053101_);
  xor g_111669_(out[314], out[762], _053102_);
  xor g_111670_(out[309], out[757], _053103_);
  xor g_111671_(out[319], out[767], _053104_);
  xor g_111672_(out[317], out[765], _053105_);
  xor g_111673_(out[312], out[760], _053106_);
  or g_111674_(_053093_, _053095_, _053108_);
  or g_111675_(_053105_, _053106_, _053109_);
  or g_111676_(_053097_, _053102_, _053110_);
  or g_111677_(_053109_, _053110_, _053111_);
  or g_111678_(_053094_, _053098_, _053112_);
  or g_111679_(_053099_, _053103_, _053113_);
  or g_111680_(_053112_, _053113_, _053114_);
  or g_111681_(_053111_, _053114_, _053115_);
  xor g_111682_(out[316], out[764], _053116_);
  or g_111683_(_053100_, _053116_, _053117_);
  xor g_111684_(out[311], out[759], _053119_);
  or g_111685_(_053101_, _053119_, _053120_);
  or g_111686_(_053117_, _053120_, _053121_);
  or g_111687_(_053091_, _053092_, _053122_);
  or g_111688_(_053104_, _053122_, _053123_);
  or g_111689_(_053121_, _053123_, _053124_);
  or g_111690_(_053115_, _053124_, _053125_);
  or g_111691_(_053108_, _053125_, _053126_);
  xor g_111692_(out[295], out[759], _053127_);
  and g_111693_(_098272_, out[763], _053128_);
  xor g_111694_(out[302], out[766], _053130_);
  xor g_111695_(out[296], out[760], _053131_);
  xor g_111696_(out[289], out[753], _053132_);
  xor g_111697_(out[301], out[765], _053133_);
  xor g_111698_(out[297], out[761], _053134_);
  xor g_111699_(out[292], out[756], _053135_);
  xor g_111700_(out[290], out[754], _053136_);
  and g_111701_(out[299], _049686_, _053137_);
  xor g_111702_(out[291], out[755], _053138_);
  xor g_111703_(out[294], out[758], _053139_);
  xor g_111704_(out[303], out[767], _053141_);
  xor g_111705_(out[298], out[762], _053142_);
  xor g_111706_(out[293], out[757], _053143_);
  xor g_111707_(out[288], out[752], _053144_);
  or g_111708_(_053130_, _053135_, _053145_);
  or g_111709_(_053131_, _053133_, _053146_);
  or g_111710_(_053136_, _053142_, _053147_);
  or g_111711_(_053146_, _053147_, _053148_);
  or g_111712_(_053134_, _053138_, _053149_);
  or g_111713_(_053143_, _053144_, _053150_);
  or g_111714_(_053149_, _053150_, _053152_);
  or g_111715_(_053148_, _053152_, _053153_);
  xor g_111716_(out[300], out[764], _053154_);
  or g_111717_(_053128_, _053154_, _053155_);
  or g_111718_(_053127_, _053139_, _053156_);
  or g_111719_(_053155_, _053156_, _053157_);
  or g_111720_(_053132_, _053137_, _053158_);
  or g_111721_(_053141_, _053158_, _053159_);
  or g_111722_(_053157_, _053159_, _053160_);
  or g_111723_(_053153_, _053160_, _053161_);
  or g_111724_(_053145_, _053161_, _053163_);
  and g_111725_(out[283], _049686_, _053164_);
  and g_111726_(_098261_, out[763], _053165_);
  xor g_111727_(out[285], out[765], _053166_);
  xor g_111728_(out[282], out[762], _053167_);
  xor g_111729_(out[277], out[757], _053168_);
  xor g_111730_(out[284], out[764], _053169_);
  xor g_111731_(out[272], out[752], _053170_);
  xor g_111732_(out[274], out[754], _053171_);
  xor g_111733_(out[275], out[755], _053172_);
  xor g_111734_(out[281], out[761], _053174_);
  xor g_111735_(out[286], out[766], _053175_);
  xor g_111736_(out[287], out[767], _053176_);
  xor g_111737_(out[273], out[753], _053177_);
  xor g_111738_(out[278], out[758], _053178_);
  xor g_111739_(out[276], out[756], _053179_);
  xor g_111740_(out[280], out[760], _053180_);
  or g_111741_(_053166_, _053180_, _053181_);
  or g_111742_(_053167_, _053171_, _053182_);
  or g_111743_(_053181_, _053182_, _053183_);
  or g_111744_(_053172_, _053174_, _053185_);
  or g_111745_(_053168_, _053185_, _053186_);
  or g_111746_(_053183_, _053186_, _053187_);
  or g_111747_(_053175_, _053179_, _053188_);
  or g_111748_(_053187_, _053188_, _053189_);
  or g_111749_(_053165_, _053169_, _053190_);
  xor g_111750_(out[279], out[759], _053191_);
  or g_111751_(_053178_, _053191_, _053192_);
  or g_111752_(_053190_, _053192_, _053193_);
  or g_111753_(_053164_, _053177_, _053194_);
  or g_111754_(_053176_, _053194_, _053196_);
  or g_111755_(_053193_, _053196_, _053197_);
  or g_111756_(_053170_, _053197_, _053198_);
  or g_111757_(_053189_, _053198_, _053199_);
  not g_111758_(_053199_, _053200_);
  xor g_111759_(out[263], out[759], _053201_);
  and g_111760_(_098250_, out[763], _053202_);
  xor g_111761_(out[270], out[766], _053203_);
  xor g_111762_(out[264], out[760], _053204_);
  xor g_111763_(out[257], out[753], _053205_);
  xor g_111764_(out[269], out[765], _053207_);
  xor g_111765_(out[265], out[761], _053208_);
  xor g_111766_(out[260], out[756], _053209_);
  xor g_111767_(out[258], out[754], _053210_);
  and g_111768_(out[267], _049686_, _053211_);
  xor g_111769_(out[259], out[755], _053212_);
  xor g_111770_(out[262], out[758], _053213_);
  xor g_111771_(out[271], out[767], _053214_);
  xor g_111772_(out[266], out[762], _053215_);
  xor g_111773_(out[261], out[757], _053216_);
  xor g_111774_(out[256], out[752], _053218_);
  or g_111775_(_053203_, _053209_, _053219_);
  or g_111776_(_053204_, _053207_, _053220_);
  or g_111777_(_053210_, _053215_, _053221_);
  or g_111778_(_053220_, _053221_, _053222_);
  or g_111779_(_053208_, _053212_, _053223_);
  or g_111780_(_053216_, _053218_, _053224_);
  or g_111781_(_053223_, _053224_, _053225_);
  or g_111782_(_053222_, _053225_, _053226_);
  xor g_111783_(out[268], out[764], _053227_);
  or g_111784_(_053202_, _053227_, _053229_);
  or g_111785_(_053201_, _053213_, _053230_);
  or g_111786_(_053229_, _053230_, _053231_);
  or g_111787_(_053205_, _053211_, _053232_);
  or g_111788_(_053214_, _053232_, _053233_);
  or g_111789_(_053231_, _053233_, _053234_);
  or g_111790_(_053226_, _053234_, _053235_);
  or g_111791_(_053219_, _053235_, _053236_);
  not g_111792_(_053236_, _053237_);
  xor g_111793_(out[241], out[753], _053238_);
  and g_111794_(out[251], _049686_, _053240_);
  xor g_111795_(out[249], out[761], _053241_);
  xor g_111796_(out[240], out[752], _053242_);
  xor g_111797_(out[254], out[766], _053243_);
  xor g_111798_(out[244], out[756], _053244_);
  or g_111799_(_053243_, _053244_, _053245_);
  xor g_111800_(out[253], out[765], _053246_);
  xor g_111801_(out[243], out[755], _053247_);
  and g_111802_(_098239_, out[763], _053248_);
  xor g_111803_(out[246], out[758], _053249_);
  xor g_111804_(out[250], out[762], _053251_);
  xor g_111805_(out[245], out[757], _053252_);
  xor g_111806_(out[255], out[767], _053253_);
  xor g_111807_(out[248], out[760], _053254_);
  or g_111808_(_053246_, _053254_, _053255_);
  xor g_111809_(out[242], out[754], _053256_);
  or g_111810_(_053251_, _053256_, _053257_);
  or g_111811_(_053255_, _053257_, _053258_);
  or g_111812_(_053241_, _053247_, _053259_);
  or g_111813_(_053252_, _053259_, _053260_);
  or g_111814_(_053258_, _053260_, _053262_);
  or g_111815_(_053245_, _053262_, _053263_);
  xor g_111816_(out[252], out[764], _053264_);
  or g_111817_(_053248_, _053264_, _053265_);
  xor g_111818_(out[247], out[759], _053266_);
  or g_111819_(_053249_, _053266_, _053267_);
  or g_111820_(_053265_, _053267_, _053268_);
  or g_111821_(_053238_, _053240_, _053269_);
  or g_111822_(_053253_, _053269_, _053270_);
  or g_111823_(_053268_, _053270_, _053271_);
  or g_111824_(_053242_, _053271_, _053273_);
  or g_111825_(_053263_, _053273_, _053274_);
  xor g_111826_(out[231], out[759], _053275_);
  and g_111827_(_098228_, out[763], _053276_);
  xor g_111828_(out[238], out[766], _053277_);
  xor g_111829_(out[232], out[760], _053278_);
  xor g_111830_(out[225], out[753], _053279_);
  xor g_111831_(out[237], out[765], _053280_);
  xor g_111832_(out[233], out[761], _053281_);
  xor g_111833_(out[228], out[756], _053282_);
  xor g_111834_(out[226], out[754], _053284_);
  and g_111835_(out[235], _049686_, _053285_);
  xor g_111836_(out[227], out[755], _053286_);
  xor g_111837_(out[230], out[758], _053287_);
  xor g_111838_(out[239], out[767], _053288_);
  xor g_111839_(out[234], out[762], _053289_);
  xor g_111840_(out[229], out[757], _053290_);
  xor g_111841_(out[224], out[752], _053291_);
  or g_111842_(_053277_, _053282_, _053292_);
  or g_111843_(_053278_, _053280_, _053293_);
  or g_111844_(_053284_, _053289_, _053295_);
  or g_111845_(_053293_, _053295_, _053296_);
  or g_111846_(_053281_, _053286_, _053297_);
  or g_111847_(_053290_, _053291_, _053298_);
  or g_111848_(_053297_, _053298_, _053299_);
  or g_111849_(_053296_, _053299_, _053300_);
  xor g_111850_(out[236], out[764], _053301_);
  or g_111851_(_053276_, _053301_, _053302_);
  or g_111852_(_053275_, _053287_, _053303_);
  or g_111853_(_053302_, _053303_, _053304_);
  or g_111854_(_053279_, _053285_, _053306_);
  or g_111855_(_053288_, _053306_, _053307_);
  or g_111856_(_053304_, _053307_, _053308_);
  or g_111857_(_053300_, _053308_, _053309_);
  or g_111858_(_053292_, _053309_, _053310_);
  xor g_111859_(out[218], out[762], _053311_);
  xor g_111860_(out[210], out[754], _053312_);
  xor g_111861_(out[209], out[753], _053313_);
  and g_111862_(_098217_, out[763], _053314_);
  and g_111863_(out[219], _049686_, _053315_);
  xor g_111864_(out[221], out[765], _053317_);
  xor g_111865_(out[211], out[755], _053318_);
  xor g_111866_(out[222], out[766], _053319_);
  xor g_111867_(out[220], out[764], _053320_);
  xor g_111868_(out[216], out[760], _053321_);
  xor g_111869_(out[223], out[767], _053322_);
  xor g_111870_(out[213], out[757], _053323_);
  xor g_111871_(out[214], out[758], _053324_);
  xor g_111872_(out[208], out[752], _053325_);
  xor g_111873_(out[212], out[756], _053326_);
  or g_111874_(_053317_, _053321_, _053328_);
  xor g_111875_(out[217], out[761], _053329_);
  or g_111876_(_053311_, _053312_, _053330_);
  or g_111877_(_053328_, _053330_, _053331_);
  or g_111878_(_053318_, _053329_, _053332_);
  or g_111879_(_053323_, _053332_, _053333_);
  or g_111880_(_053331_, _053333_, _053334_);
  or g_111881_(_053319_, _053326_, _053335_);
  or g_111882_(_053334_, _053335_, _053336_);
  or g_111883_(_053314_, _053320_, _053337_);
  xor g_111884_(out[215], out[759], _053339_);
  or g_111885_(_053324_, _053339_, _053340_);
  or g_111886_(_053337_, _053340_, _053341_);
  or g_111887_(_053313_, _053315_, _053342_);
  or g_111888_(_053322_, _053342_, _053343_);
  or g_111889_(_053341_, _053343_, _053344_);
  or g_111890_(_053325_, _053344_, _053345_);
  or g_111891_(_053336_, _053345_, _053346_);
  not g_111892_(_053346_, _053347_);
  xor g_111893_(out[199], out[759], _053348_);
  and g_111894_(_098206_, out[763], _053350_);
  xor g_111895_(out[206], out[766], _053351_);
  xor g_111896_(out[200], out[760], _053352_);
  xor g_111897_(out[193], out[753], _053353_);
  xor g_111898_(out[205], out[765], _053354_);
  xor g_111899_(out[201], out[761], _053355_);
  xor g_111900_(out[196], out[756], _053356_);
  xor g_111901_(out[194], out[754], _053357_);
  and g_111902_(out[203], _049686_, _053358_);
  xor g_111903_(out[195], out[755], _053359_);
  xor g_111904_(out[198], out[758], _053361_);
  xor g_111905_(out[207], out[767], _053362_);
  xor g_111906_(out[202], out[762], _053363_);
  xor g_111907_(out[197], out[757], _053364_);
  xor g_111908_(out[192], out[752], _053365_);
  or g_111909_(_053351_, _053356_, _053366_);
  or g_111910_(_053352_, _053354_, _053367_);
  or g_111911_(_053357_, _053363_, _053368_);
  or g_111912_(_053367_, _053368_, _053369_);
  or g_111913_(_053355_, _053359_, _053370_);
  or g_111914_(_053364_, _053365_, _053372_);
  or g_111915_(_053370_, _053372_, _053373_);
  or g_111916_(_053369_, _053373_, _053374_);
  xor g_111917_(out[204], out[764], _053375_);
  or g_111918_(_053350_, _053375_, _053376_);
  or g_111919_(_053348_, _053361_, _053377_);
  or g_111920_(_053376_, _053377_, _053378_);
  or g_111921_(_053353_, _053358_, _053379_);
  or g_111922_(_053362_, _053379_, _053380_);
  or g_111923_(_053378_, _053380_, _053381_);
  or g_111924_(_053374_, _053381_, _053383_);
  or g_111925_(_053366_, _053383_, _053384_);
  xor g_111926_(out[188], out[764], _053385_);
  and g_111927_(_098195_, out[763], _053386_);
  xor g_111928_(out[184], out[760], _053387_);
  xor g_111929_(out[182], out[758], _053388_);
  xor g_111930_(out[189], out[765], _053389_);
  xor g_111931_(out[190], out[766], _053390_);
  xor g_111932_(out[178], out[754], _053391_);
  xor g_111933_(out[185], out[761], _053392_);
  xor g_111934_(out[181], out[757], _053394_);
  xor g_111935_(out[177], out[753], _053395_);
  and g_111936_(out[187], _049686_, _053396_);
  or g_111937_(_053387_, _053389_, _053397_);
  xor g_111938_(out[191], out[767], _053398_);
  xor g_111939_(out[186], out[762], _053399_);
  xor g_111940_(out[180], out[756], _053400_);
  xor g_111941_(out[179], out[755], _053401_);
  xor g_111942_(out[176], out[752], _053402_);
  or g_111943_(_053391_, _053399_, _053403_);
  or g_111944_(_053397_, _053403_, _053405_);
  or g_111945_(_053392_, _053401_, _053406_);
  or g_111946_(_053394_, _053406_, _053407_);
  or g_111947_(_053405_, _053407_, _053408_);
  or g_111948_(_053390_, _053400_, _053409_);
  or g_111949_(_053408_, _053409_, _053410_);
  or g_111950_(_053385_, _053386_, _053411_);
  xor g_111951_(out[183], out[759], _053412_);
  or g_111952_(_053388_, _053412_, _053413_);
  or g_111953_(_053411_, _053413_, _053414_);
  or g_111954_(_053395_, _053396_, _053416_);
  or g_111955_(_053398_, _053416_, _053417_);
  or g_111956_(_053414_, _053417_, _053418_);
  or g_111957_(_053402_, _053418_, _053419_);
  or g_111958_(_053410_, _053419_, _053420_);
  xor g_111959_(out[167], out[759], _053421_);
  and g_111960_(_098184_, out[763], _053422_);
  xor g_111961_(out[174], out[766], _053423_);
  xor g_111962_(out[168], out[760], _053424_);
  xor g_111963_(out[161], out[753], _053425_);
  xor g_111964_(out[173], out[765], _053427_);
  xor g_111965_(out[169], out[761], _053428_);
  xor g_111966_(out[164], out[756], _053429_);
  xor g_111967_(out[162], out[754], _053430_);
  and g_111968_(out[171], _049686_, _053431_);
  xor g_111969_(out[163], out[755], _053432_);
  xor g_111970_(out[166], out[758], _053433_);
  xor g_111971_(out[175], out[767], _053434_);
  xor g_111972_(out[170], out[762], _053435_);
  xor g_111973_(out[165], out[757], _053436_);
  xor g_111974_(out[160], out[752], _053438_);
  or g_111975_(_053423_, _053429_, _053439_);
  or g_111976_(_053424_, _053427_, _053440_);
  or g_111977_(_053430_, _053435_, _053441_);
  or g_111978_(_053440_, _053441_, _053442_);
  or g_111979_(_053428_, _053432_, _053443_);
  or g_111980_(_053436_, _053438_, _053444_);
  or g_111981_(_053443_, _053444_, _053445_);
  or g_111982_(_053442_, _053445_, _053446_);
  xor g_111983_(out[172], out[764], _053447_);
  or g_111984_(_053422_, _053447_, _053449_);
  or g_111985_(_053421_, _053433_, _053450_);
  or g_111986_(_053449_, _053450_, _053451_);
  or g_111987_(_053425_, _053431_, _053452_);
  or g_111988_(_053434_, _053452_, _053453_);
  or g_111989_(_053451_, _053453_, _053454_);
  or g_111990_(_053446_, _053454_, _053455_);
  or g_111991_(_053439_, _053455_, _053456_);
  not g_111992_(_053456_, _053457_);
  xor g_111993_(out[145], out[753], _053458_);
  and g_111994_(_098173_, out[763], _053460_);
  and g_111995_(out[155], _049686_, _053461_);
  xor g_111996_(out[153], out[761], _053462_);
  xor g_111997_(out[144], out[752], _053463_);
  xor g_111998_(out[158], out[766], _053464_);
  xor g_111999_(out[148], out[756], _053465_);
  or g_112000_(_053464_, _053465_, _053466_);
  xor g_112001_(out[157], out[765], _053467_);
  xor g_112002_(out[147], out[755], _053468_);
  xor g_112003_(out[156], out[764], _053469_);
  xor g_112004_(out[150], out[758], _053471_);
  xor g_112005_(out[154], out[762], _053472_);
  xor g_112006_(out[149], out[757], _053473_);
  xor g_112007_(out[159], out[767], _053474_);
  xor g_112008_(out[152], out[760], _053475_);
  or g_112009_(_053467_, _053475_, _053476_);
  xor g_112010_(out[146], out[754], _053477_);
  or g_112011_(_053472_, _053477_, _053478_);
  or g_112012_(_053476_, _053478_, _053479_);
  or g_112013_(_053462_, _053468_, _053480_);
  or g_112014_(_053473_, _053480_, _053482_);
  or g_112015_(_053479_, _053482_, _053483_);
  or g_112016_(_053466_, _053483_, _053484_);
  or g_112017_(_053460_, _053469_, _053485_);
  xor g_112018_(out[151], out[759], _053486_);
  or g_112019_(_053471_, _053486_, _053487_);
  or g_112020_(_053485_, _053487_, _053488_);
  or g_112021_(_053458_, _053461_, _053489_);
  or g_112022_(_053474_, _053489_, _053490_);
  or g_112023_(_053488_, _053490_, _053491_);
  or g_112024_(_053463_, _053491_, _053493_);
  or g_112025_(_053484_, _053493_, _053494_);
  not g_112026_(_053494_, _053495_);
  xor g_112027_(out[135], out[759], _053496_);
  and g_112028_(_098162_, out[763], _053497_);
  xor g_112029_(out[142], out[766], _053498_);
  xor g_112030_(out[136], out[760], _053499_);
  xor g_112031_(out[129], out[753], _053500_);
  xor g_112032_(out[141], out[765], _053501_);
  xor g_112033_(out[137], out[761], _053502_);
  xor g_112034_(out[132], out[756], _053504_);
  xor g_112035_(out[130], out[754], _053505_);
  and g_112036_(out[139], _049686_, _053506_);
  xor g_112037_(out[131], out[755], _053507_);
  xor g_112038_(out[134], out[758], _053508_);
  xor g_112039_(out[143], out[767], _053509_);
  xor g_112040_(out[138], out[762], _053510_);
  xor g_112041_(out[133], out[757], _053511_);
  xor g_112042_(out[128], out[752], _053512_);
  or g_112043_(_053498_, _053504_, _053513_);
  or g_112044_(_053499_, _053501_, _053515_);
  or g_112045_(_053505_, _053510_, _053516_);
  or g_112046_(_053515_, _053516_, _053517_);
  or g_112047_(_053502_, _053507_, _053518_);
  or g_112048_(_053511_, _053512_, _053519_);
  or g_112049_(_053518_, _053519_, _053520_);
  or g_112050_(_053517_, _053520_, _053521_);
  xor g_112051_(out[140], out[764], _053522_);
  or g_112052_(_053497_, _053522_, _053523_);
  or g_112053_(_053496_, _053508_, _053524_);
  or g_112054_(_053523_, _053524_, _053526_);
  or g_112055_(_053500_, _053506_, _053527_);
  or g_112056_(_053509_, _053527_, _053528_);
  or g_112057_(_053526_, _053528_, _053529_);
  or g_112058_(_053521_, _053529_, _053530_);
  or g_112059_(_053513_, _053530_, _053531_);
  xor g_112060_(out[120], out[760], _053532_);
  xor g_112061_(out[117], out[757], _053533_);
  xor g_112062_(out[115], out[755], _053534_);
  xor g_112063_(out[126], out[766], _053535_);
  xor g_112064_(out[125], out[765], _053537_);
  xor g_112065_(out[114], out[754], _053538_);
  xor g_112066_(out[121], out[761], _053539_);
  xor g_112067_(out[118], out[758], _053540_);
  xor g_112068_(out[127], out[767], _053541_);
  xor g_112069_(out[122], out[762], _053542_);
  xor g_112070_(out[116], out[756], _053543_);
  xor g_112071_(out[112], out[752], _053544_);
  and g_112072_(_098151_, out[763], _053545_);
  and g_112073_(out[123], _049686_, _053546_);
  or g_112074_(_053532_, _053537_, _053548_);
  xor g_112075_(out[113], out[753], _053549_);
  or g_112076_(_053538_, _053542_, _053550_);
  or g_112077_(_053548_, _053550_, _053551_);
  or g_112078_(_053534_, _053539_, _053552_);
  or g_112079_(_053533_, _053552_, _053553_);
  or g_112080_(_053551_, _053553_, _053554_);
  or g_112081_(_053535_, _053543_, _053555_);
  or g_112082_(_053554_, _053555_, _053556_);
  xor g_112083_(out[124], out[764], _053557_);
  or g_112084_(_053545_, _053557_, _053559_);
  xor g_112085_(out[119], out[759], _053560_);
  or g_112086_(_053540_, _053560_, _053561_);
  or g_112087_(_053559_, _053561_, _053562_);
  or g_112088_(_053546_, _053549_, _053563_);
  or g_112089_(_053541_, _053563_, _053564_);
  or g_112090_(_053562_, _053564_, _053565_);
  or g_112091_(_053544_, _053565_, _053566_);
  or g_112092_(_053556_, _053566_, _053567_);
  xor g_112093_(out[103], out[759], _053568_);
  and g_112094_(_098140_, out[763], _053570_);
  xor g_112095_(out[110], out[766], _053571_);
  xor g_112096_(out[104], out[760], _053572_);
  xor g_112097_(out[97], out[753], _053573_);
  xor g_112098_(out[109], out[765], _053574_);
  xor g_112099_(out[105], out[761], _053575_);
  xor g_112100_(out[100], out[756], _053576_);
  xor g_112101_(out[98], out[754], _053577_);
  and g_112102_(out[107], _049686_, _053578_);
  xor g_112103_(out[99], out[755], _053579_);
  xor g_112104_(out[102], out[758], _053581_);
  xor g_112105_(out[111], out[767], _053582_);
  xor g_112106_(out[106], out[762], _053583_);
  xor g_112107_(out[101], out[757], _053584_);
  xor g_112108_(out[96], out[752], _053585_);
  or g_112109_(_053571_, _053576_, _053586_);
  or g_112110_(_053572_, _053574_, _053587_);
  or g_112111_(_053577_, _053583_, _053588_);
  or g_112112_(_053587_, _053588_, _053589_);
  or g_112113_(_053575_, _053579_, _053590_);
  or g_112114_(_053584_, _053585_, _053592_);
  or g_112115_(_053590_, _053592_, _053593_);
  or g_112116_(_053589_, _053593_, _053594_);
  xor g_112117_(out[108], out[764], _053595_);
  or g_112118_(_053570_, _053595_, _053596_);
  or g_112119_(_053568_, _053581_, _053597_);
  or g_112120_(_053596_, _053597_, _053598_);
  or g_112121_(_053573_, _053578_, _053599_);
  or g_112122_(_053582_, _053599_, _053600_);
  or g_112123_(_053598_, _053600_, _053601_);
  or g_112124_(_053594_, _053601_, _053603_);
  or g_112125_(_053586_, _053603_, _053604_);
  xor g_112126_(out[92], out[764], _053605_);
  and g_112127_(_098129_, out[763], _053606_);
  xor g_112128_(out[93], out[765], _053607_);
  xor g_112129_(out[86], out[758], _053608_);
  xor g_112130_(out[88], out[760], _053609_);
  xor g_112131_(out[89], out[761], _053610_);
  xor g_112132_(out[94], out[766], _053611_);
  xor g_112133_(out[84], out[756], _053612_);
  or g_112134_(_053611_, _053612_, _053614_);
  xor g_112135_(out[85], out[757], _053615_);
  xor g_112136_(out[81], out[753], _053616_);
  and g_112137_(out[91], _049686_, _053617_);
  xor g_112138_(out[95], out[767], _053618_);
  xor g_112139_(out[90], out[762], _053619_);
  xor g_112140_(out[80], out[752], _053620_);
  xor g_112141_(out[82], out[754], _053621_);
  xor g_112142_(out[83], out[755], _053622_);
  or g_112143_(_053607_, _053609_, _053623_);
  or g_112144_(_053619_, _053621_, _053625_);
  or g_112145_(_053623_, _053625_, _053626_);
  or g_112146_(_053610_, _053622_, _053627_);
  or g_112147_(_053615_, _053620_, _053628_);
  or g_112148_(_053627_, _053628_, _053629_);
  or g_112149_(_053626_, _053629_, _053630_);
  or g_112150_(_053605_, _053606_, _053631_);
  xor g_112151_(out[87], out[759], _053632_);
  or g_112152_(_053608_, _053632_, _053633_);
  or g_112153_(_053631_, _053633_, _053634_);
  or g_112154_(_053616_, _053617_, _053636_);
  or g_112155_(_053618_, _053636_, _053637_);
  or g_112156_(_053634_, _053637_, _053638_);
  or g_112157_(_053630_, _053638_, _053639_);
  or g_112158_(_053614_, _053639_, _053640_);
  xor g_112159_(out[71], out[759], _053641_);
  and g_112160_(_098118_, out[763], _053642_);
  xor g_112161_(out[78], out[766], _053643_);
  xor g_112162_(out[72], out[760], _053644_);
  xor g_112163_(out[65], out[753], _053645_);
  xor g_112164_(out[77], out[765], _053647_);
  xor g_112165_(out[73], out[761], _053648_);
  xor g_112166_(out[68], out[756], _053649_);
  xor g_112167_(out[66], out[754], _053650_);
  and g_112168_(out[75], _049686_, _053651_);
  xor g_112169_(out[67], out[755], _053652_);
  xor g_112170_(out[70], out[758], _053653_);
  xor g_112171_(out[79], out[767], _053654_);
  xor g_112172_(out[74], out[762], _053655_);
  xor g_112173_(out[69], out[757], _053656_);
  xor g_112174_(out[64], out[752], _053658_);
  or g_112175_(_053643_, _053649_, _053659_);
  or g_112176_(_053644_, _053647_, _053660_);
  or g_112177_(_053650_, _053655_, _053661_);
  or g_112178_(_053660_, _053661_, _053662_);
  or g_112179_(_053648_, _053652_, _053663_);
  or g_112180_(_053656_, _053658_, _053664_);
  or g_112181_(_053663_, _053664_, _053665_);
  or g_112182_(_053662_, _053665_, _053666_);
  xor g_112183_(out[76], out[764], _053667_);
  or g_112184_(_053642_, _053667_, _053669_);
  or g_112185_(_053641_, _053653_, _053670_);
  or g_112186_(_053669_, _053670_, _053671_);
  or g_112187_(_053645_, _053651_, _053672_);
  or g_112188_(_053654_, _053672_, _053673_);
  or g_112189_(_053671_, _053673_, _053674_);
  or g_112190_(_053666_, _053674_, _053675_);
  or g_112191_(_053659_, _053675_, _053676_);
  xor g_112192_(out[49], out[753], _053677_);
  and g_112193_(_098107_, out[763], _053678_);
  and g_112194_(out[59], _049686_, _053680_);
  xor g_112195_(out[62], out[766], _053681_);
  xor g_112196_(out[51], out[755], _053682_);
  xor g_112197_(out[52], out[756], _053683_);
  xor g_112198_(out[50], out[754], _053684_);
  xor g_112199_(out[57], out[761], _053685_);
  xor g_112200_(out[48], out[752], _053686_);
  xor g_112201_(out[60], out[764], _053687_);
  xor g_112202_(out[54], out[758], _053688_);
  xor g_112203_(out[58], out[762], _053689_);
  xor g_112204_(out[53], out[757], _053691_);
  xor g_112205_(out[63], out[767], _053692_);
  xor g_112206_(out[61], out[765], _053693_);
  xor g_112207_(out[56], out[760], _053694_);
  or g_112208_(_053681_, _053683_, _053695_);
  or g_112209_(_053693_, _053694_, _053696_);
  or g_112210_(_053684_, _053689_, _053697_);
  or g_112211_(_053696_, _053697_, _053698_);
  or g_112212_(_053682_, _053685_, _053699_);
  or g_112213_(_053686_, _053691_, _053700_);
  or g_112214_(_053699_, _053700_, _053702_);
  or g_112215_(_053698_, _053702_, _053703_);
  or g_112216_(_053678_, _053687_, _053704_);
  xor g_112217_(out[55], out[759], _053705_);
  or g_112218_(_053688_, _053705_, _053706_);
  or g_112219_(_053704_, _053706_, _053707_);
  or g_112220_(_053677_, _053680_, _053708_);
  or g_112221_(_053692_, _053708_, _053709_);
  or g_112222_(_053707_, _053709_, _053710_);
  or g_112223_(_053703_, _053710_, _053711_);
  or g_112224_(_053695_, _053711_, _053713_);
  not g_112225_(_053713_, _053714_);
  xor g_112226_(out[39], out[759], _053715_);
  and g_112227_(_098096_, out[763], _053716_);
  xor g_112228_(out[46], out[766], _053717_);
  xor g_112229_(out[40], out[760], _053718_);
  xor g_112230_(out[33], out[753], _053719_);
  xor g_112231_(out[45], out[765], _053720_);
  xor g_112232_(out[41], out[761], _053721_);
  xor g_112233_(out[36], out[756], _053722_);
  xor g_112234_(out[34], out[754], _053724_);
  and g_112235_(out[43], _049686_, _053725_);
  xor g_112236_(out[35], out[755], _053726_);
  xor g_112237_(out[38], out[758], _053727_);
  xor g_112238_(out[47], out[767], _053728_);
  xor g_112239_(out[42], out[762], _053729_);
  xor g_112240_(out[37], out[757], _053730_);
  xor g_112241_(out[32], out[752], _053731_);
  or g_112242_(_053717_, _053722_, _053732_);
  or g_112243_(_053718_, _053720_, _053733_);
  or g_112244_(_053724_, _053729_, _053735_);
  or g_112245_(_053733_, _053735_, _053736_);
  or g_112246_(_053721_, _053726_, _053737_);
  or g_112247_(_053730_, _053731_, _053738_);
  or g_112248_(_053737_, _053738_, _053739_);
  or g_112249_(_053736_, _053739_, _053740_);
  xor g_112250_(out[44], out[764], _053741_);
  or g_112251_(_053716_, _053741_, _053742_);
  or g_112252_(_053715_, _053727_, _053743_);
  or g_112253_(_053742_, _053743_, _053744_);
  or g_112254_(_053719_, _053725_, _053746_);
  or g_112255_(_053728_, _053746_, _053747_);
  or g_112256_(_053744_, _053747_, _053748_);
  or g_112257_(_053740_, _053748_, _053749_);
  or g_112258_(_053732_, _053749_, _053750_);
  not g_112259_(_053750_, _053751_);
  xor g_112260_(out[19], out[755], _053752_);
  xor g_112261_(out[20], out[756], _053753_);
  xor g_112262_(out[30], out[766], _053754_);
  xor g_112263_(out[18], out[754], _053755_);
  xor g_112264_(out[21], out[757], _053757_);
  xor g_112265_(out[25], out[761], _053758_);
  xor g_112266_(out[24], out[760], _053759_);
  xor g_112267_(out[31], out[767], _053760_);
  xor g_112268_(out[26], out[762], _053761_);
  xor g_112269_(out[22], out[758], _053762_);
  xor g_112270_(out[16], out[752], _053763_);
  and g_112271_(_098063_, out[763], _053764_);
  and g_112272_(out[27], _049686_, _053765_);
  xor g_112273_(out[29], out[765], _053766_);
  or g_112274_(_053759_, _053766_, _053768_);
  xor g_112275_(out[17], out[753], _053769_);
  or g_112276_(_053755_, _053761_, _053770_);
  or g_112277_(_053768_, _053770_, _053771_);
  or g_112278_(_053752_, _053758_, _053772_);
  or g_112279_(_053757_, _053772_, _053773_);
  or g_112280_(_053771_, _053773_, _053774_);
  or g_112281_(_053753_, _053754_, _053775_);
  or g_112282_(_053774_, _053775_, _053776_);
  xor g_112283_(out[28], out[764], _053777_);
  or g_112284_(_053764_, _053777_, _053779_);
  xor g_112285_(out[23], out[759], _053780_);
  or g_112286_(_053762_, _053780_, _053781_);
  or g_112287_(_053779_, _053781_, _053782_);
  or g_112288_(_053765_, _053769_, _053783_);
  or g_112289_(_053760_, _053783_, _053784_);
  or g_112290_(_053782_, _053784_, _053785_);
  or g_112291_(_053763_, _053785_, _053786_);
  or g_112292_(_053776_, _053786_, _053787_);
  and g_112293_(out[11], _049686_, _053788_);
  and g_112294_(_098041_, out[763], _053790_);
  xor g_112295_(out[8], out[760], _053791_);
  xor g_112296_(out[15], out[767], _053792_);
  xor g_112297_(out[1], out[753], _053793_);
  xor g_112298_(out[2], out[754], _053794_);
  xor g_112299_(out[4], out[756], _053795_);
  xor g_112300_(out[13], out[765], _053796_);
  xor g_112301_(out[9], out[761], _053797_);
  xor g_112302_(out[3], out[755], _053798_);
  xor g_112303_(out[5], out[757], _053799_);
  xor g_112304_(out[14], out[766], _053801_);
  xor g_112305_(out[0], out[752], _053802_);
  xor g_112306_(out[10], out[762], _053803_);
  or g_112307_(_053791_, _053796_, _053804_);
  xor g_112308_(out[6], out[758], _053805_);
  or g_112309_(_053794_, _053803_, _053806_);
  or g_112310_(_053804_, _053806_, _053807_);
  or g_112311_(_053797_, _053798_, _053808_);
  or g_112312_(_053799_, _053808_, _053809_);
  or g_112313_(_053807_, _053809_, _053810_);
  or g_112314_(_053795_, _053801_, _053812_);
  or g_112315_(_053810_, _053812_, _053813_);
  xor g_112316_(out[12], out[764], _053814_);
  or g_112317_(_053790_, _053814_, _053815_);
  xor g_112318_(out[7], out[759], _053816_);
  or g_112319_(_053805_, _053816_, _053817_);
  or g_112320_(_053815_, _053817_, _053818_);
  or g_112321_(_053788_, _053793_, _053819_);
  or g_112322_(_053792_, _053819_, _053820_);
  or g_112323_(_053818_, _053820_, _053821_);
  or g_112324_(_053802_, _053821_, _053823_);
  or g_112325_(_053813_, _053823_, _053824_);
  xor g_112326_(out[471], out[743], _053825_);
  and g_112327_(_049499_, out[747], _053826_);
  xor g_112328_(out[478], out[750], _053827_);
  xor g_112329_(out[472], out[744], _053828_);
  xor g_112330_(out[465], out[737], _053829_);
  xor g_112331_(out[477], out[749], _053830_);
  xor g_112332_(out[473], out[745], _053831_);
  xor g_112333_(out[468], out[740], _053832_);
  xor g_112334_(out[466], out[738], _053834_);
  and g_112335_(out[475], _049675_, _053835_);
  xor g_112336_(out[467], out[739], _053836_);
  xor g_112337_(out[470], out[742], _053837_);
  xor g_112338_(out[479], out[751], _053838_);
  xor g_112339_(out[474], out[746], _053839_);
  xor g_112340_(out[469], out[741], _053840_);
  xor g_112341_(out[464], out[736], _053841_);
  or g_112342_(_053827_, _053832_, _053842_);
  or g_112343_(_053828_, _053830_, _053843_);
  or g_112344_(_053834_, _053839_, _053845_);
  or g_112345_(_053843_, _053845_, _053846_);
  or g_112346_(_053831_, _053836_, _053847_);
  or g_112347_(_053840_, _053841_, _053848_);
  or g_112348_(_053847_, _053848_, _053849_);
  or g_112349_(_053846_, _053849_, _053850_);
  xor g_112350_(out[476], out[748], _053851_);
  or g_112351_(_053826_, _053851_, _053852_);
  or g_112352_(_053825_, _053837_, _053853_);
  or g_112353_(_053852_, _053853_, _053854_);
  or g_112354_(_053829_, _053835_, _053856_);
  or g_112355_(_053838_, _053856_, _053857_);
  or g_112356_(_053854_, _053857_, _053858_);
  or g_112357_(_053850_, _053858_, _053859_);
  or g_112358_(_053842_, _053859_, _053860_);
  xor g_112359_(out[460], out[748], _053861_);
  and g_112360_(_049477_, out[747], _053862_);
  xor g_112361_(out[456], out[744], _053863_);
  xor g_112362_(out[454], out[742], _053864_);
  xor g_112363_(out[461], out[749], _053865_);
  xor g_112364_(out[462], out[750], _053867_);
  xor g_112365_(out[450], out[738], _053868_);
  xor g_112366_(out[457], out[745], _053869_);
  xor g_112367_(out[453], out[741], _053870_);
  xor g_112368_(out[449], out[737], _053871_);
  and g_112369_(out[459], _049675_, _053872_);
  or g_112370_(_053863_, _053865_, _053873_);
  xor g_112371_(out[463], out[751], _053874_);
  xor g_112372_(out[458], out[746], _053875_);
  xor g_112373_(out[452], out[740], _053876_);
  xor g_112374_(out[451], out[739], _053878_);
  xor g_112375_(out[448], out[736], _053879_);
  or g_112376_(_053868_, _053875_, _053880_);
  or g_112377_(_053873_, _053880_, _053881_);
  or g_112378_(_053869_, _053878_, _053882_);
  or g_112379_(_053870_, _053882_, _053883_);
  or g_112380_(_053881_, _053883_, _053884_);
  or g_112381_(_053867_, _053876_, _053885_);
  or g_112382_(_053884_, _053885_, _053886_);
  or g_112383_(_053861_, _053862_, _053887_);
  xor g_112384_(out[455], out[743], _053889_);
  or g_112385_(_053864_, _053889_, _053890_);
  or g_112386_(_053887_, _053890_, _053891_);
  or g_112387_(_053871_, _053872_, _053892_);
  or g_112388_(_053874_, _053892_, _053893_);
  or g_112389_(_053891_, _053893_, _053894_);
  or g_112390_(_053879_, _053894_, _053895_);
  or g_112391_(_053886_, _053895_, _053896_);
  xor g_112392_(out[439], out[743], _053897_);
  and g_112393_(_049466_, out[747], _053898_);
  xor g_112394_(out[446], out[750], _053900_);
  xor g_112395_(out[440], out[744], _053901_);
  xor g_112396_(out[433], out[737], _053902_);
  xor g_112397_(out[445], out[749], _053903_);
  xor g_112398_(out[441], out[745], _053904_);
  xor g_112399_(out[436], out[740], _053905_);
  xor g_112400_(out[434], out[738], _053906_);
  and g_112401_(out[443], _049675_, _053907_);
  xor g_112402_(out[435], out[739], _053908_);
  xor g_112403_(out[438], out[742], _053909_);
  xor g_112404_(out[447], out[751], _053911_);
  xor g_112405_(out[442], out[746], _053912_);
  xor g_112406_(out[437], out[741], _053913_);
  xor g_112407_(out[432], out[736], _053914_);
  or g_112408_(_053900_, _053905_, _053915_);
  or g_112409_(_053901_, _053903_, _053916_);
  or g_112410_(_053906_, _053912_, _053917_);
  or g_112411_(_053916_, _053917_, _053918_);
  or g_112412_(_053904_, _053908_, _053919_);
  or g_112413_(_053913_, _053914_, _053920_);
  or g_112414_(_053919_, _053920_, _053922_);
  or g_112415_(_053918_, _053922_, _053923_);
  xor g_112416_(out[444], out[748], _053924_);
  or g_112417_(_053898_, _053924_, _053925_);
  or g_112418_(_053897_, _053909_, _053926_);
  or g_112419_(_053925_, _053926_, _053927_);
  or g_112420_(_053902_, _053907_, _053928_);
  or g_112421_(_053911_, _053928_, _053929_);
  or g_112422_(_053927_, _053929_, _053930_);
  or g_112423_(_053923_, _053930_, _053931_);
  or g_112424_(_053915_, _053931_, _053933_);
  not g_112425_(_053933_, _053934_);
  and g_112426_(out[427], _049675_, _053935_);
  xor g_112427_(out[420], out[740], _053936_);
  xor g_112428_(out[430], out[750], _053937_);
  or g_112429_(_053936_, _053937_, _053938_);
  xor g_112430_(out[429], out[749], _053939_);
  xor g_112431_(out[419], out[739], _053940_);
  xor g_112432_(out[416], out[736], _053941_);
  and g_112433_(_049455_, out[747], _053942_);
  xor g_112434_(out[426], out[746], _053944_);
  xor g_112435_(out[431], out[751], _053945_);
  xor g_112436_(out[422], out[742], _053946_);
  xor g_112437_(out[421], out[741], _053947_);
  xor g_112438_(out[424], out[744], _053948_);
  or g_112439_(_053939_, _053948_, _053949_);
  xor g_112440_(out[418], out[738], _053950_);
  xor g_112441_(out[425], out[745], _053951_);
  xor g_112442_(out[417], out[737], _053952_);
  or g_112443_(_053944_, _053950_, _053953_);
  or g_112444_(_053949_, _053953_, _053955_);
  or g_112445_(_053940_, _053951_, _053956_);
  or g_112446_(_053947_, _053956_, _053957_);
  or g_112447_(_053955_, _053957_, _053958_);
  or g_112448_(_053938_, _053958_, _053959_);
  xor g_112449_(out[428], out[748], _053960_);
  or g_112450_(_053942_, _053960_, _053961_);
  xor g_112451_(out[423], out[743], _053962_);
  or g_112452_(_053946_, _053962_, _053963_);
  or g_112453_(_053961_, _053963_, _053964_);
  or g_112454_(_053935_, _053952_, _053966_);
  or g_112455_(_053945_, _053966_, _053967_);
  or g_112456_(_053964_, _053967_, _053968_);
  or g_112457_(_053941_, _053968_, _053969_);
  or g_112458_(_053959_, _053969_, _053970_);
  not g_112459_(_053970_, _053971_);
  xor g_112460_(out[407], out[743], _053972_);
  and g_112461_(_049444_, out[747], _053973_);
  xor g_112462_(out[414], out[750], _053974_);
  xor g_112463_(out[408], out[744], _053975_);
  xor g_112464_(out[401], out[737], _053977_);
  xor g_112465_(out[413], out[749], _053978_);
  xor g_112466_(out[409], out[745], _053979_);
  xor g_112467_(out[404], out[740], _053980_);
  xor g_112468_(out[402], out[738], _053981_);
  and g_112469_(out[411], _049675_, _053982_);
  xor g_112470_(out[403], out[739], _053983_);
  xor g_112471_(out[406], out[742], _053984_);
  xor g_112472_(out[415], out[751], _053985_);
  xor g_112473_(out[410], out[746], _053986_);
  xor g_112474_(out[405], out[741], _053988_);
  xor g_112475_(out[400], out[736], _053989_);
  or g_112476_(_053974_, _053980_, _053990_);
  or g_112477_(_053975_, _053978_, _053991_);
  or g_112478_(_053981_, _053986_, _053992_);
  or g_112479_(_053991_, _053992_, _053993_);
  or g_112480_(_053979_, _053983_, _053994_);
  or g_112481_(_053988_, _053989_, _053995_);
  or g_112482_(_053994_, _053995_, _053996_);
  or g_112483_(_053993_, _053996_, _053997_);
  xor g_112484_(out[412], out[748], _053999_);
  or g_112485_(_053973_, _053999_, _054000_);
  or g_112486_(_053972_, _053984_, _054001_);
  or g_112487_(_054000_, _054001_, _054002_);
  or g_112488_(_053977_, _053982_, _054003_);
  or g_112489_(_053985_, _054003_, _054004_);
  or g_112490_(_054002_, _054004_, _054005_);
  or g_112491_(_053997_, _054005_, _054006_);
  or g_112492_(_053990_, _054006_, _054007_);
  xor g_112493_(out[394], out[746], _054008_);
  xor g_112494_(out[392], out[744], _054010_);
  xor g_112495_(out[385], out[737], _054011_);
  and g_112496_(_049433_, out[747], _054012_);
  and g_112497_(out[395], _049675_, _054013_);
  xor g_112498_(out[386], out[738], _054014_);
  xor g_112499_(out[389], out[741], _054015_);
  xor g_112500_(out[393], out[745], _054016_);
  xor g_112501_(out[396], out[748], _054017_);
  xor g_112502_(out[397], out[749], _054018_);
  xor g_112503_(out[399], out[751], _054019_);
  xor g_112504_(out[388], out[740], _054021_);
  xor g_112505_(out[390], out[742], _054022_);
  xor g_112506_(out[387], out[739], _054023_);
  xor g_112507_(out[384], out[736], _054024_);
  xor g_112508_(out[398], out[750], _054025_);
  or g_112509_(_054021_, _054025_, _054026_);
  or g_112510_(_054010_, _054018_, _054027_);
  or g_112511_(_054008_, _054014_, _054028_);
  or g_112512_(_054027_, _054028_, _054029_);
  or g_112513_(_054016_, _054023_, _054030_);
  or g_112514_(_054015_, _054024_, _054032_);
  or g_112515_(_054030_, _054032_, _054033_);
  or g_112516_(_054029_, _054033_, _054034_);
  or g_112517_(_054012_, _054017_, _054035_);
  xor g_112518_(out[391], out[743], _054036_);
  or g_112519_(_054022_, _054036_, _054037_);
  or g_112520_(_054035_, _054037_, _054038_);
  or g_112521_(_054011_, _054013_, _054039_);
  or g_112522_(_054019_, _054039_, _054040_);
  or g_112523_(_054038_, _054040_, _054041_);
  or g_112524_(_054034_, _054041_, _054043_);
  or g_112525_(_054026_, _054043_, _054044_);
  xor g_112526_(out[375], out[743], _054045_);
  and g_112527_(_049422_, out[747], _054046_);
  xor g_112528_(out[382], out[750], _054047_);
  xor g_112529_(out[376], out[744], _054048_);
  xor g_112530_(out[369], out[737], _054049_);
  xor g_112531_(out[381], out[749], _054050_);
  xor g_112532_(out[377], out[745], _054051_);
  xor g_112533_(out[372], out[740], _054052_);
  xor g_112534_(out[370], out[738], _054054_);
  and g_112535_(out[379], _049675_, _054055_);
  xor g_112536_(out[371], out[739], _054056_);
  xor g_112537_(out[374], out[742], _054057_);
  xor g_112538_(out[383], out[751], _054058_);
  xor g_112539_(out[378], out[746], _054059_);
  xor g_112540_(out[373], out[741], _054060_);
  xor g_112541_(out[368], out[736], _054061_);
  or g_112542_(_054047_, _054052_, _054062_);
  or g_112543_(_054048_, _054050_, _054063_);
  or g_112544_(_054054_, _054059_, _054065_);
  or g_112545_(_054063_, _054065_, _054066_);
  or g_112546_(_054051_, _054056_, _054067_);
  or g_112547_(_054060_, _054061_, _054068_);
  or g_112548_(_054067_, _054068_, _054069_);
  or g_112549_(_054066_, _054069_, _054070_);
  xor g_112550_(out[380], out[748], _054071_);
  or g_112551_(_054046_, _054071_, _054072_);
  or g_112552_(_054045_, _054057_, _054073_);
  or g_112553_(_054072_, _054073_, _054074_);
  or g_112554_(_054049_, _054055_, _054076_);
  or g_112555_(_054058_, _054076_, _054077_);
  or g_112556_(_054074_, _054077_, _054078_);
  or g_112557_(_054070_, _054078_, _054079_);
  or g_112558_(_054062_, _054079_, _054080_);
  not g_112559_(_054080_, _054081_);
  xor g_112560_(out[353], out[737], _054082_);
  and g_112561_(out[363], _049675_, _054083_);
  xor g_112562_(out[361], out[745], _054084_);
  xor g_112563_(out[352], out[736], _054085_);
  xor g_112564_(out[366], out[750], _054087_);
  xor g_112565_(out[356], out[740], _054088_);
  or g_112566_(_054087_, _054088_, _054089_);
  xor g_112567_(out[365], out[749], _054090_);
  xor g_112568_(out[355], out[739], _054091_);
  and g_112569_(_049411_, out[747], _054092_);
  xor g_112570_(out[358], out[742], _054093_);
  xor g_112571_(out[362], out[746], _054094_);
  xor g_112572_(out[357], out[741], _054095_);
  xor g_112573_(out[367], out[751], _054096_);
  xor g_112574_(out[360], out[744], _054098_);
  or g_112575_(_054090_, _054098_, _054099_);
  xor g_112576_(out[354], out[738], _054100_);
  or g_112577_(_054094_, _054100_, _054101_);
  or g_112578_(_054099_, _054101_, _054102_);
  or g_112579_(_054084_, _054091_, _054103_);
  or g_112580_(_054095_, _054103_, _054104_);
  or g_112581_(_054102_, _054104_, _054105_);
  or g_112582_(_054089_, _054105_, _054106_);
  xor g_112583_(out[364], out[748], _054107_);
  or g_112584_(_054092_, _054107_, _054109_);
  xor g_112585_(out[359], out[743], _054110_);
  or g_112586_(_054093_, _054110_, _054111_);
  or g_112587_(_054109_, _054111_, _054112_);
  or g_112588_(_054082_, _054083_, _054113_);
  or g_112589_(_054096_, _054113_, _054114_);
  or g_112590_(_054112_, _054114_, _054115_);
  or g_112591_(_054085_, _054115_, _054116_);
  or g_112592_(_054106_, _054116_, _054117_);
  xor g_112593_(out[343], out[743], _054118_);
  and g_112594_(_049400_, out[747], _054120_);
  xor g_112595_(out[350], out[750], _054121_);
  xor g_112596_(out[344], out[744], _054122_);
  xor g_112597_(out[337], out[737], _054123_);
  xor g_112598_(out[349], out[749], _054124_);
  xor g_112599_(out[345], out[745], _054125_);
  xor g_112600_(out[340], out[740], _054126_);
  xor g_112601_(out[338], out[738], _054127_);
  and g_112602_(out[347], _049675_, _054128_);
  xor g_112603_(out[339], out[739], _054129_);
  xor g_112604_(out[342], out[742], _054131_);
  xor g_112605_(out[351], out[751], _054132_);
  xor g_112606_(out[346], out[746], _054133_);
  xor g_112607_(out[341], out[741], _054134_);
  xor g_112608_(out[336], out[736], _054135_);
  or g_112609_(_054121_, _054126_, _054136_);
  or g_112610_(_054122_, _054124_, _054137_);
  or g_112611_(_054127_, _054133_, _054138_);
  or g_112612_(_054137_, _054138_, _054139_);
  or g_112613_(_054125_, _054129_, _054140_);
  or g_112614_(_054134_, _054135_, _054142_);
  or g_112615_(_054140_, _054142_, _054143_);
  or g_112616_(_054139_, _054143_, _054144_);
  xor g_112617_(out[348], out[748], _054145_);
  or g_112618_(_054120_, _054145_, _054146_);
  or g_112619_(_054118_, _054131_, _054147_);
  or g_112620_(_054146_, _054147_, _054148_);
  or g_112621_(_054123_, _054128_, _054149_);
  or g_112622_(_054132_, _054149_, _054150_);
  or g_112623_(_054148_, _054150_, _054151_);
  or g_112624_(_054144_, _054151_, _054153_);
  or g_112625_(_054136_, _054153_, _054154_);
  xor g_112626_(out[328], out[744], _054155_);
  xor g_112627_(out[325], out[741], _054156_);
  xor g_112628_(out[323], out[739], _054157_);
  xor g_112629_(out[334], out[750], _054158_);
  xor g_112630_(out[333], out[749], _054159_);
  xor g_112631_(out[322], out[738], _054160_);
  xor g_112632_(out[329], out[745], _054161_);
  xor g_112633_(out[326], out[742], _054162_);
  xor g_112634_(out[335], out[751], _054164_);
  xor g_112635_(out[330], out[746], _054165_);
  xor g_112636_(out[324], out[740], _054166_);
  xor g_112637_(out[320], out[736], _054167_);
  and g_112638_(_098294_, out[747], _054168_);
  and g_112639_(out[331], _049675_, _054169_);
  or g_112640_(_054155_, _054159_, _054170_);
  xor g_112641_(out[321], out[737], _054171_);
  or g_112642_(_054160_, _054165_, _054172_);
  or g_112643_(_054170_, _054172_, _054173_);
  or g_112644_(_054157_, _054161_, _054175_);
  or g_112645_(_054156_, _054175_, _054176_);
  or g_112646_(_054173_, _054176_, _054177_);
  or g_112647_(_054158_, _054166_, _054178_);
  or g_112648_(_054177_, _054178_, _054179_);
  xor g_112649_(out[332], out[748], _054180_);
  or g_112650_(_054168_, _054180_, _054181_);
  xor g_112651_(out[327], out[743], _054182_);
  or g_112652_(_054162_, _054182_, _054183_);
  or g_112653_(_054181_, _054183_, _054184_);
  or g_112654_(_054169_, _054171_, _054186_);
  or g_112655_(_054164_, _054186_, _054187_);
  or g_112656_(_054184_, _054187_, _054188_);
  or g_112657_(_054167_, _054188_, _054189_);
  or g_112658_(_054179_, _054189_, _054190_);
  not g_112659_(_054190_, _054191_);
  xor g_112660_(out[311], out[743], _054192_);
  and g_112661_(_098283_, out[747], _054193_);
  xor g_112662_(out[318], out[750], _054194_);
  xor g_112663_(out[312], out[744], _054195_);
  xor g_112664_(out[305], out[737], _054197_);
  xor g_112665_(out[317], out[749], _054198_);
  xor g_112666_(out[313], out[745], _054199_);
  xor g_112667_(out[308], out[740], _054200_);
  xor g_112668_(out[306], out[738], _054201_);
  and g_112669_(out[315], _049675_, _054202_);
  xor g_112670_(out[307], out[739], _054203_);
  xor g_112671_(out[310], out[742], _054204_);
  xor g_112672_(out[319], out[751], _054205_);
  xor g_112673_(out[314], out[746], _054206_);
  xor g_112674_(out[309], out[741], _054208_);
  xor g_112675_(out[304], out[736], _054209_);
  or g_112676_(_054194_, _054200_, _054210_);
  or g_112677_(_054195_, _054198_, _054211_);
  or g_112678_(_054201_, _054206_, _054212_);
  or g_112679_(_054211_, _054212_, _054213_);
  or g_112680_(_054199_, _054203_, _054214_);
  or g_112681_(_054208_, _054209_, _054215_);
  or g_112682_(_054214_, _054215_, _054216_);
  or g_112683_(_054213_, _054216_, _054217_);
  xor g_112684_(out[316], out[748], _054219_);
  or g_112685_(_054193_, _054219_, _054220_);
  or g_112686_(_054192_, _054204_, _054221_);
  or g_112687_(_054220_, _054221_, _054222_);
  or g_112688_(_054197_, _054202_, _054223_);
  or g_112689_(_054205_, _054223_, _054224_);
  or g_112690_(_054222_, _054224_, _054225_);
  or g_112691_(_054217_, _054225_, _054226_);
  or g_112692_(_054210_, _054226_, _054227_);
  not g_112693_(_054227_, _054228_);
  xor g_112694_(out[289], out[737], _054230_);
  and g_112695_(out[299], _049675_, _054231_);
  xor g_112696_(out[297], out[745], _054232_);
  xor g_112697_(out[288], out[736], _054233_);
  xor g_112698_(out[302], out[750], _054234_);
  xor g_112699_(out[292], out[740], _054235_);
  or g_112700_(_054234_, _054235_, _054236_);
  xor g_112701_(out[301], out[749], _054237_);
  xor g_112702_(out[291], out[739], _054238_);
  and g_112703_(_098272_, out[747], _054239_);
  xor g_112704_(out[294], out[742], _054241_);
  xor g_112705_(out[298], out[746], _054242_);
  xor g_112706_(out[293], out[741], _054243_);
  xor g_112707_(out[303], out[751], _054244_);
  xor g_112708_(out[296], out[744], _054245_);
  or g_112709_(_054237_, _054245_, _054246_);
  xor g_112710_(out[290], out[738], _054247_);
  or g_112711_(_054242_, _054247_, _054248_);
  or g_112712_(_054246_, _054248_, _054249_);
  or g_112713_(_054232_, _054238_, _054250_);
  or g_112714_(_054243_, _054250_, _054252_);
  or g_112715_(_054249_, _054252_, _054253_);
  or g_112716_(_054236_, _054253_, _054254_);
  xor g_112717_(out[300], out[748], _054255_);
  or g_112718_(_054239_, _054255_, _054256_);
  xor g_112719_(out[295], out[743], _054257_);
  or g_112720_(_054241_, _054257_, _054258_);
  or g_112721_(_054256_, _054258_, _054259_);
  or g_112722_(_054230_, _054231_, _054260_);
  or g_112723_(_054244_, _054260_, _054261_);
  or g_112724_(_054259_, _054261_, _054263_);
  or g_112725_(_054233_, _054263_, _054264_);
  or g_112726_(_054254_, _054264_, _054265_);
  xor g_112727_(out[279], out[743], _054266_);
  and g_112728_(_098261_, out[747], _054267_);
  xor g_112729_(out[286], out[750], _054268_);
  xor g_112730_(out[280], out[744], _054269_);
  xor g_112731_(out[273], out[737], _054270_);
  xor g_112732_(out[285], out[749], _054271_);
  xor g_112733_(out[281], out[745], _054272_);
  xor g_112734_(out[276], out[740], _054274_);
  xor g_112735_(out[274], out[738], _054275_);
  and g_112736_(out[283], _049675_, _054276_);
  xor g_112737_(out[275], out[739], _054277_);
  xor g_112738_(out[278], out[742], _054278_);
  xor g_112739_(out[287], out[751], _054279_);
  xor g_112740_(out[282], out[746], _054280_);
  xor g_112741_(out[277], out[741], _054281_);
  xor g_112742_(out[272], out[736], _054282_);
  or g_112743_(_054268_, _054274_, _054283_);
  or g_112744_(_054269_, _054271_, _054285_);
  or g_112745_(_054275_, _054280_, _054286_);
  or g_112746_(_054285_, _054286_, _054287_);
  or g_112747_(_054272_, _054277_, _054288_);
  or g_112748_(_054281_, _054282_, _054289_);
  or g_112749_(_054288_, _054289_, _054290_);
  or g_112750_(_054287_, _054290_, _054291_);
  xor g_112751_(out[284], out[748], _054292_);
  or g_112752_(_054267_, _054292_, _054293_);
  or g_112753_(_054266_, _054278_, _054294_);
  or g_112754_(_054293_, _054294_, _054296_);
  or g_112755_(_054270_, _054276_, _054297_);
  or g_112756_(_054279_, _054297_, _054298_);
  or g_112757_(_054296_, _054298_, _054299_);
  or g_112758_(_054291_, _054299_, _054300_);
  or g_112759_(_054283_, _054300_, _054301_);
  xor g_112760_(out[264], out[744], _054302_);
  xor g_112761_(out[261], out[741], _054303_);
  xor g_112762_(out[259], out[739], _054304_);
  xor g_112763_(out[270], out[750], _054305_);
  xor g_112764_(out[269], out[749], _054307_);
  xor g_112765_(out[258], out[738], _054308_);
  xor g_112766_(out[265], out[745], _054309_);
  xor g_112767_(out[262], out[742], _054310_);
  xor g_112768_(out[271], out[751], _054311_);
  xor g_112769_(out[266], out[746], _054312_);
  xor g_112770_(out[260], out[740], _054313_);
  xor g_112771_(out[256], out[736], _054314_);
  and g_112772_(_098250_, out[747], _054315_);
  and g_112773_(out[267], _049675_, _054316_);
  or g_112774_(_054302_, _054307_, _054318_);
  xor g_112775_(out[257], out[737], _054319_);
  or g_112776_(_054308_, _054312_, _054320_);
  or g_112777_(_054318_, _054320_, _054321_);
  or g_112778_(_054304_, _054309_, _054322_);
  or g_112779_(_054303_, _054322_, _054323_);
  or g_112780_(_054321_, _054323_, _054324_);
  or g_112781_(_054305_, _054313_, _054325_);
  or g_112782_(_054324_, _054325_, _054326_);
  xor g_112783_(out[268], out[748], _054327_);
  or g_112784_(_054315_, _054327_, _054329_);
  xor g_112785_(out[263], out[743], _054330_);
  or g_112786_(_054310_, _054330_, _054331_);
  or g_112787_(_054329_, _054331_, _054332_);
  or g_112788_(_054316_, _054319_, _054333_);
  or g_112789_(_054311_, _054333_, _054334_);
  or g_112790_(_054332_, _054334_, _054335_);
  or g_112791_(_054314_, _054335_, _054336_);
  or g_112792_(_054326_, _054336_, _054337_);
  not g_112793_(_054337_, _054338_);
  xor g_112794_(out[247], out[743], _054340_);
  and g_112795_(_098239_, out[747], _054341_);
  xor g_112796_(out[254], out[750], _054342_);
  xor g_112797_(out[248], out[744], _054343_);
  xor g_112798_(out[241], out[737], _054344_);
  xor g_112799_(out[253], out[749], _054345_);
  xor g_112800_(out[249], out[745], _054346_);
  xor g_112801_(out[244], out[740], _054347_);
  xor g_112802_(out[242], out[738], _054348_);
  and g_112803_(out[251], _049675_, _054349_);
  xor g_112804_(out[243], out[739], _054351_);
  xor g_112805_(out[246], out[742], _054352_);
  xor g_112806_(out[255], out[751], _054353_);
  xor g_112807_(out[250], out[746], _054354_);
  xor g_112808_(out[245], out[741], _054355_);
  xor g_112809_(out[240], out[736], _054356_);
  or g_112810_(_054342_, _054347_, _054357_);
  or g_112811_(_054343_, _054345_, _054358_);
  or g_112812_(_054348_, _054354_, _054359_);
  or g_112813_(_054358_, _054359_, _054360_);
  or g_112814_(_054346_, _054351_, _054362_);
  or g_112815_(_054355_, _054356_, _054363_);
  or g_112816_(_054362_, _054363_, _054364_);
  or g_112817_(_054360_, _054364_, _054365_);
  xor g_112818_(out[252], out[748], _054366_);
  or g_112819_(_054341_, _054366_, _054367_);
  or g_112820_(_054340_, _054352_, _054368_);
  or g_112821_(_054367_, _054368_, _054369_);
  or g_112822_(_054344_, _054349_, _054370_);
  or g_112823_(_054353_, _054370_, _054371_);
  or g_112824_(_054369_, _054371_, _054373_);
  or g_112825_(_054365_, _054373_, _054374_);
  or g_112826_(_054357_, _054374_, _054375_);
  xor g_112827_(out[236], out[748], _054376_);
  and g_112828_(_098228_, out[747], _054377_);
  xor g_112829_(out[232], out[744], _054378_);
  xor g_112830_(out[230], out[742], _054379_);
  xor g_112831_(out[237], out[749], _054380_);
  xor g_112832_(out[238], out[750], _054381_);
  xor g_112833_(out[226], out[738], _054382_);
  xor g_112834_(out[233], out[745], _054384_);
  xor g_112835_(out[229], out[741], _054385_);
  xor g_112836_(out[225], out[737], _054386_);
  and g_112837_(out[235], _049675_, _054387_);
  or g_112838_(_054378_, _054380_, _054388_);
  xor g_112839_(out[239], out[751], _054389_);
  xor g_112840_(out[234], out[746], _054390_);
  xor g_112841_(out[228], out[740], _054391_);
  xor g_112842_(out[227], out[739], _054392_);
  xor g_112843_(out[224], out[736], _054393_);
  or g_112844_(_054382_, _054390_, _054395_);
  or g_112845_(_054388_, _054395_, _054396_);
  or g_112846_(_054384_, _054392_, _054397_);
  or g_112847_(_054385_, _054397_, _054398_);
  or g_112848_(_054396_, _054398_, _054399_);
  or g_112849_(_054381_, _054391_, _054400_);
  or g_112850_(_054399_, _054400_, _054401_);
  or g_112851_(_054376_, _054377_, _054402_);
  xor g_112852_(out[231], out[743], _054403_);
  or g_112853_(_054379_, _054403_, _054404_);
  or g_112854_(_054402_, _054404_, _054406_);
  or g_112855_(_054386_, _054387_, _054407_);
  or g_112856_(_054389_, _054407_, _054408_);
  or g_112857_(_054406_, _054408_, _054409_);
  or g_112858_(_054393_, _054409_, _054410_);
  or g_112859_(_054401_, _054410_, _054411_);
  xor g_112860_(out[215], out[743], _054412_);
  and g_112861_(_098217_, out[747], _054413_);
  xor g_112862_(out[222], out[750], _054414_);
  xor g_112863_(out[216], out[744], _054415_);
  xor g_112864_(out[209], out[737], _054417_);
  xor g_112865_(out[221], out[749], _054418_);
  xor g_112866_(out[217], out[745], _054419_);
  xor g_112867_(out[212], out[740], _054420_);
  xor g_112868_(out[210], out[738], _054421_);
  and g_112869_(out[219], _049675_, _054422_);
  xor g_112870_(out[211], out[739], _054423_);
  xor g_112871_(out[214], out[742], _054424_);
  xor g_112872_(out[223], out[751], _054425_);
  xor g_112873_(out[218], out[746], _054426_);
  xor g_112874_(out[213], out[741], _054428_);
  xor g_112875_(out[208], out[736], _054429_);
  or g_112876_(_054414_, _054420_, _054430_);
  or g_112877_(_054415_, _054418_, _054431_);
  or g_112878_(_054421_, _054426_, _054432_);
  or g_112879_(_054431_, _054432_, _054433_);
  or g_112880_(_054419_, _054423_, _054434_);
  or g_112881_(_054428_, _054429_, _054435_);
  or g_112882_(_054434_, _054435_, _054436_);
  or g_112883_(_054433_, _054436_, _054437_);
  xor g_112884_(out[220], out[748], _054439_);
  or g_112885_(_054413_, _054439_, _054440_);
  or g_112886_(_054412_, _054424_, _054441_);
  or g_112887_(_054440_, _054441_, _054442_);
  or g_112888_(_054417_, _054422_, _054443_);
  or g_112889_(_054425_, _054443_, _054444_);
  or g_112890_(_054442_, _054444_, _054445_);
  or g_112891_(_054437_, _054445_, _054446_);
  or g_112892_(_054430_, _054446_, _054447_);
  and g_112893_(out[203], _049675_, _054448_);
  and g_112894_(_098206_, out[747], _054450_);
  xor g_112895_(out[200], out[744], _054451_);
  xor g_112896_(out[207], out[751], _054452_);
  xor g_112897_(out[193], out[737], _054453_);
  xor g_112898_(out[194], out[738], _054454_);
  xor g_112899_(out[196], out[740], _054455_);
  xor g_112900_(out[205], out[749], _054456_);
  xor g_112901_(out[201], out[745], _054457_);
  xor g_112902_(out[195], out[739], _054458_);
  xor g_112903_(out[197], out[741], _054459_);
  xor g_112904_(out[206], out[750], _054461_);
  xor g_112905_(out[192], out[736], _054462_);
  xor g_112906_(out[202], out[746], _054463_);
  or g_112907_(_054451_, _054456_, _054464_);
  xor g_112908_(out[198], out[742], _054465_);
  or g_112909_(_054454_, _054463_, _054466_);
  or g_112910_(_054464_, _054466_, _054467_);
  or g_112911_(_054457_, _054458_, _054468_);
  or g_112912_(_054459_, _054468_, _054469_);
  or g_112913_(_054467_, _054469_, _054470_);
  or g_112914_(_054455_, _054461_, _054472_);
  or g_112915_(_054470_, _054472_, _054473_);
  xor g_112916_(out[204], out[748], _054474_);
  or g_112917_(_054450_, _054474_, _054475_);
  xor g_112918_(out[199], out[743], _054476_);
  or g_112919_(_054465_, _054476_, _054477_);
  or g_112920_(_054475_, _054477_, _054478_);
  or g_112921_(_054448_, _054453_, _054479_);
  or g_112922_(_054452_, _054479_, _054480_);
  or g_112923_(_054478_, _054480_, _054481_);
  or g_112924_(_054462_, _054481_, _054483_);
  or g_112925_(_054473_, _054483_, _054484_);
  xor g_112926_(out[183], out[743], _054485_);
  and g_112927_(_098195_, out[747], _054486_);
  xor g_112928_(out[190], out[750], _054487_);
  xor g_112929_(out[184], out[744], _054488_);
  xor g_112930_(out[177], out[737], _054489_);
  xor g_112931_(out[189], out[749], _054490_);
  xor g_112932_(out[185], out[745], _054491_);
  xor g_112933_(out[180], out[740], _054492_);
  xor g_112934_(out[178], out[738], _054494_);
  and g_112935_(out[187], _049675_, _054495_);
  xor g_112936_(out[179], out[739], _054496_);
  xor g_112937_(out[182], out[742], _054497_);
  xor g_112938_(out[191], out[751], _054498_);
  xor g_112939_(out[186], out[746], _054499_);
  xor g_112940_(out[181], out[741], _054500_);
  xor g_112941_(out[176], out[736], _054501_);
  or g_112942_(_054487_, _054492_, _054502_);
  or g_112943_(_054488_, _054490_, _054503_);
  or g_112944_(_054494_, _054499_, _054505_);
  or g_112945_(_054503_, _054505_, _054506_);
  or g_112946_(_054491_, _054496_, _054507_);
  or g_112947_(_054500_, _054501_, _054508_);
  or g_112948_(_054507_, _054508_, _054509_);
  or g_112949_(_054506_, _054509_, _054510_);
  xor g_112950_(out[188], out[748], _054511_);
  or g_112951_(_054486_, _054511_, _054512_);
  or g_112952_(_054485_, _054497_, _054513_);
  or g_112953_(_054512_, _054513_, _054514_);
  or g_112954_(_054489_, _054495_, _054516_);
  or g_112955_(_054498_, _054516_, _054517_);
  or g_112956_(_054514_, _054517_, _054518_);
  or g_112957_(_054510_, _054518_, _054519_);
  or g_112958_(_054502_, _054519_, _054520_);
  xor g_112959_(out[170], out[746], _054521_);
  xor g_112960_(out[162], out[738], _054522_);
  xor g_112961_(out[161], out[737], _054523_);
  and g_112962_(_098184_, out[747], _054524_);
  and g_112963_(out[171], _049675_, _054525_);
  xor g_112964_(out[173], out[749], _054527_);
  xor g_112965_(out[163], out[739], _054528_);
  xor g_112966_(out[174], out[750], _054529_);
  xor g_112967_(out[172], out[748], _054530_);
  xor g_112968_(out[168], out[744], _054531_);
  xor g_112969_(out[175], out[751], _054532_);
  xor g_112970_(out[165], out[741], _054533_);
  xor g_112971_(out[166], out[742], _054534_);
  xor g_112972_(out[160], out[736], _054535_);
  xor g_112973_(out[164], out[740], _054536_);
  or g_112974_(_054527_, _054531_, _054538_);
  xor g_112975_(out[169], out[745], _054539_);
  or g_112976_(_054521_, _054522_, _054540_);
  or g_112977_(_054538_, _054540_, _054541_);
  or g_112978_(_054528_, _054539_, _054542_);
  or g_112979_(_054533_, _054542_, _054543_);
  or g_112980_(_054541_, _054543_, _054544_);
  or g_112981_(_054529_, _054536_, _054545_);
  or g_112982_(_054544_, _054545_, _054546_);
  or g_112983_(_054524_, _054530_, _054547_);
  xor g_112984_(out[167], out[743], _054549_);
  or g_112985_(_054534_, _054549_, _054550_);
  or g_112986_(_054547_, _054550_, _054551_);
  or g_112987_(_054523_, _054525_, _054552_);
  or g_112988_(_054532_, _054552_, _054553_);
  or g_112989_(_054551_, _054553_, _054554_);
  or g_112990_(_054535_, _054554_, _054555_);
  or g_112991_(_054546_, _054555_, _054556_);
  xor g_112992_(out[151], out[743], _054557_);
  and g_112993_(_098173_, out[747], _054558_);
  xor g_112994_(out[158], out[750], _054560_);
  xor g_112995_(out[152], out[744], _054561_);
  xor g_112996_(out[145], out[737], _054562_);
  xor g_112997_(out[157], out[749], _054563_);
  xor g_112998_(out[153], out[745], _054564_);
  xor g_112999_(out[148], out[740], _054565_);
  xor g_113000_(out[146], out[738], _054566_);
  and g_113001_(out[155], _049675_, _054567_);
  xor g_113002_(out[147], out[739], _054568_);
  xor g_113003_(out[150], out[742], _054569_);
  xor g_113004_(out[159], out[751], _054571_);
  xor g_113005_(out[154], out[746], _054572_);
  xor g_113006_(out[149], out[741], _054573_);
  xor g_113007_(out[144], out[736], _054574_);
  or g_113008_(_054560_, _054565_, _054575_);
  or g_113009_(_054561_, _054563_, _054576_);
  or g_113010_(_054566_, _054572_, _054577_);
  or g_113011_(_054576_, _054577_, _054578_);
  or g_113012_(_054564_, _054568_, _054579_);
  or g_113013_(_054573_, _054574_, _054580_);
  or g_113014_(_054579_, _054580_, _054582_);
  or g_113015_(_054578_, _054582_, _054583_);
  xor g_113016_(out[156], out[748], _054584_);
  or g_113017_(_054558_, _054584_, _054585_);
  or g_113018_(_054557_, _054569_, _054586_);
  or g_113019_(_054585_, _054586_, _054587_);
  or g_113020_(_054562_, _054567_, _054588_);
  or g_113021_(_054571_, _054588_, _054589_);
  or g_113022_(_054587_, _054589_, _054590_);
  or g_113023_(_054583_, _054590_, _054591_);
  or g_113024_(_054575_, _054591_, _054593_);
  xor g_113025_(out[131], out[739], _054594_);
  xor g_113026_(out[132], out[740], _054595_);
  xor g_113027_(out[142], out[750], _054596_);
  xor g_113028_(out[130], out[738], _054597_);
  xor g_113029_(out[133], out[741], _054598_);
  xor g_113030_(out[137], out[745], _054599_);
  xor g_113031_(out[136], out[744], _054600_);
  xor g_113032_(out[143], out[751], _054601_);
  xor g_113033_(out[138], out[746], _054602_);
  xor g_113034_(out[134], out[742], _054604_);
  xor g_113035_(out[128], out[736], _054605_);
  and g_113036_(_098162_, out[747], _054606_);
  and g_113037_(out[139], _049675_, _054607_);
  xor g_113038_(out[141], out[749], _054608_);
  or g_113039_(_054600_, _054608_, _054609_);
  xor g_113040_(out[129], out[737], _054610_);
  or g_113041_(_054597_, _054602_, _054611_);
  or g_113042_(_054609_, _054611_, _054612_);
  or g_113043_(_054594_, _054599_, _054613_);
  or g_113044_(_054598_, _054613_, _054615_);
  or g_113045_(_054612_, _054615_, _054616_);
  or g_113046_(_054595_, _054596_, _054617_);
  or g_113047_(_054616_, _054617_, _054618_);
  xor g_113048_(out[140], out[748], _054619_);
  or g_113049_(_054606_, _054619_, _054620_);
  xor g_113050_(out[135], out[743], _054621_);
  or g_113051_(_054604_, _054621_, _054622_);
  or g_113052_(_054620_, _054622_, _054623_);
  or g_113053_(_054607_, _054610_, _054624_);
  or g_113054_(_054601_, _054624_, _054626_);
  or g_113055_(_054623_, _054626_, _054627_);
  or g_113056_(_054605_, _054627_, _054628_);
  or g_113057_(_054618_, _054628_, _054629_);
  xor g_113058_(out[119], out[743], _054630_);
  and g_113059_(_098151_, out[747], _054631_);
  xor g_113060_(out[126], out[750], _054632_);
  xor g_113061_(out[120], out[744], _054633_);
  xor g_113062_(out[113], out[737], _054634_);
  xor g_113063_(out[125], out[749], _054635_);
  xor g_113064_(out[121], out[745], _054637_);
  xor g_113065_(out[116], out[740], _054638_);
  xor g_113066_(out[114], out[738], _054639_);
  and g_113067_(out[123], _049675_, _054640_);
  xor g_113068_(out[115], out[739], _054641_);
  xor g_113069_(out[118], out[742], _054642_);
  xor g_113070_(out[127], out[751], _054643_);
  xor g_113071_(out[122], out[746], _054644_);
  xor g_113072_(out[117], out[741], _054645_);
  xor g_113073_(out[112], out[736], _054646_);
  or g_113074_(_054632_, _054638_, _054648_);
  or g_113075_(_054633_, _054635_, _054649_);
  or g_113076_(_054639_, _054644_, _054650_);
  or g_113077_(_054649_, _054650_, _054651_);
  or g_113078_(_054637_, _054641_, _054652_);
  or g_113079_(_054645_, _054646_, _054653_);
  or g_113080_(_054652_, _054653_, _054654_);
  or g_113081_(_054651_, _054654_, _054655_);
  xor g_113082_(out[124], out[748], _054656_);
  or g_113083_(_054631_, _054656_, _054657_);
  or g_113084_(_054630_, _054642_, _054659_);
  or g_113085_(_054657_, _054659_, _054660_);
  or g_113086_(_054634_, _054640_, _054661_);
  or g_113087_(_054643_, _054661_, _054662_);
  or g_113088_(_054660_, _054662_, _054663_);
  or g_113089_(_054655_, _054663_, _054664_);
  or g_113090_(_054648_, _054664_, _054665_);
  xor g_113091_(out[106], out[746], _054666_);
  xor g_113092_(out[104], out[744], _054667_);
  xor g_113093_(out[97], out[737], _054668_);
  and g_113094_(_098140_, out[747], _054670_);
  and g_113095_(out[107], _049675_, _054671_);
  xor g_113096_(out[98], out[738], _054672_);
  xor g_113097_(out[101], out[741], _054673_);
  xor g_113098_(out[105], out[745], _054674_);
  xor g_113099_(out[108], out[748], _054675_);
  xor g_113100_(out[109], out[749], _054676_);
  xor g_113101_(out[111], out[751], _054677_);
  xor g_113102_(out[100], out[740], _054678_);
  xor g_113103_(out[102], out[742], _054679_);
  xor g_113104_(out[99], out[739], _054681_);
  xor g_113105_(out[96], out[736], _054682_);
  xor g_113106_(out[110], out[750], _054683_);
  or g_113107_(_054678_, _054683_, _054684_);
  or g_113108_(_054667_, _054676_, _054685_);
  or g_113109_(_054666_, _054672_, _054686_);
  or g_113110_(_054685_, _054686_, _054687_);
  or g_113111_(_054674_, _054681_, _054688_);
  or g_113112_(_054673_, _054682_, _054689_);
  or g_113113_(_054688_, _054689_, _054690_);
  or g_113114_(_054687_, _054690_, _054692_);
  or g_113115_(_054670_, _054675_, _054693_);
  xor g_113116_(out[103], out[743], _054694_);
  or g_113117_(_054679_, _054694_, _054695_);
  or g_113118_(_054693_, _054695_, _054696_);
  or g_113119_(_054668_, _054671_, _054697_);
  or g_113120_(_054677_, _054697_, _054698_);
  or g_113121_(_054696_, _054698_, _054699_);
  or g_113122_(_054692_, _054699_, _054700_);
  or g_113123_(_054684_, _054700_, _054701_);
  xor g_113124_(out[87], out[743], _054703_);
  and g_113125_(_098129_, out[747], _054704_);
  xor g_113126_(out[94], out[750], _054705_);
  xor g_113127_(out[88], out[744], _054706_);
  xor g_113128_(out[81], out[737], _054707_);
  xor g_113129_(out[93], out[749], _054708_);
  xor g_113130_(out[89], out[745], _054709_);
  xor g_113131_(out[84], out[740], _054710_);
  xor g_113132_(out[82], out[738], _054711_);
  and g_113133_(out[91], _049675_, _054712_);
  xor g_113134_(out[83], out[739], _054714_);
  xor g_113135_(out[86], out[742], _054715_);
  xor g_113136_(out[95], out[751], _054716_);
  xor g_113137_(out[90], out[746], _054717_);
  xor g_113138_(out[85], out[741], _054718_);
  xor g_113139_(out[80], out[736], _054719_);
  or g_113140_(_054705_, _054710_, _054720_);
  or g_113141_(_054706_, _054708_, _054721_);
  or g_113142_(_054711_, _054717_, _054722_);
  or g_113143_(_054721_, _054722_, _054723_);
  or g_113144_(_054709_, _054714_, _054725_);
  or g_113145_(_054718_, _054719_, _054726_);
  or g_113146_(_054725_, _054726_, _054727_);
  or g_113147_(_054723_, _054727_, _054728_);
  xor g_113148_(out[92], out[748], _054729_);
  or g_113149_(_054704_, _054729_, _054730_);
  or g_113150_(_054703_, _054715_, _054731_);
  or g_113151_(_054730_, _054731_, _054732_);
  or g_113152_(_054707_, _054712_, _054733_);
  or g_113153_(_054716_, _054733_, _054734_);
  or g_113154_(_054732_, _054734_, _054736_);
  or g_113155_(_054728_, _054736_, _054737_);
  or g_113156_(_054720_, _054737_, _054738_);
  xor g_113157_(out[72], out[744], _054739_);
  xor g_113158_(out[69], out[741], _054740_);
  xor g_113159_(out[67], out[739], _054741_);
  xor g_113160_(out[78], out[750], _054742_);
  xor g_113161_(out[77], out[749], _054743_);
  xor g_113162_(out[66], out[738], _054744_);
  xor g_113163_(out[73], out[745], _054745_);
  xor g_113164_(out[70], out[742], _054747_);
  xor g_113165_(out[79], out[751], _054748_);
  xor g_113166_(out[74], out[746], _054749_);
  xor g_113167_(out[68], out[740], _054750_);
  xor g_113168_(out[64], out[736], _054751_);
  and g_113169_(_098118_, out[747], _054752_);
  and g_113170_(out[75], _049675_, _054753_);
  or g_113171_(_054739_, _054743_, _054754_);
  xor g_113172_(out[65], out[737], _054755_);
  or g_113173_(_054744_, _054749_, _054756_);
  or g_113174_(_054754_, _054756_, _054758_);
  or g_113175_(_054741_, _054745_, _054759_);
  or g_113176_(_054740_, _054759_, _054760_);
  or g_113177_(_054758_, _054760_, _054761_);
  or g_113178_(_054742_, _054750_, _054762_);
  or g_113179_(_054761_, _054762_, _054763_);
  xor g_113180_(out[76], out[748], _054764_);
  or g_113181_(_054752_, _054764_, _054765_);
  xor g_113182_(out[71], out[743], _054766_);
  or g_113183_(_054747_, _054766_, _054767_);
  or g_113184_(_054765_, _054767_, _054769_);
  or g_113185_(_054753_, _054755_, _054770_);
  or g_113186_(_054748_, _054770_, _054771_);
  or g_113187_(_054769_, _054771_, _054772_);
  or g_113188_(_054751_, _054772_, _054773_);
  or g_113189_(_054763_, _054773_, _054774_);
  xor g_113190_(out[55], out[743], _054775_);
  and g_113191_(_098107_, out[747], _054776_);
  xor g_113192_(out[62], out[750], _054777_);
  xor g_113193_(out[56], out[744], _054778_);
  xor g_113194_(out[49], out[737], _054780_);
  xor g_113195_(out[61], out[749], _054781_);
  xor g_113196_(out[57], out[745], _054782_);
  xor g_113197_(out[52], out[740], _054783_);
  xor g_113198_(out[50], out[738], _054784_);
  and g_113199_(out[59], _049675_, _054785_);
  xor g_113200_(out[51], out[739], _054786_);
  xor g_113201_(out[54], out[742], _054787_);
  xor g_113202_(out[63], out[751], _054788_);
  xor g_113203_(out[58], out[746], _054789_);
  xor g_113204_(out[53], out[741], _054791_);
  xor g_113205_(out[48], out[736], _054792_);
  or g_113206_(_054777_, _054783_, _054793_);
  or g_113207_(_054778_, _054781_, _054794_);
  or g_113208_(_054784_, _054789_, _054795_);
  or g_113209_(_054794_, _054795_, _054796_);
  or g_113210_(_054782_, _054786_, _054797_);
  or g_113211_(_054791_, _054792_, _054798_);
  or g_113212_(_054797_, _054798_, _054799_);
  or g_113213_(_054796_, _054799_, _054800_);
  xor g_113214_(out[60], out[748], _054802_);
  or g_113215_(_054776_, _054802_, _054803_);
  or g_113216_(_054775_, _054787_, _054804_);
  or g_113217_(_054803_, _054804_, _054805_);
  or g_113218_(_054780_, _054785_, _054806_);
  or g_113219_(_054788_, _054806_, _054807_);
  or g_113220_(_054805_, _054807_, _054808_);
  or g_113221_(_054800_, _054808_, _054809_);
  or g_113222_(_054793_, _054809_, _054810_);
  not g_113223_(_054810_, _054811_);
  and g_113224_(out[43], _049675_, _054813_);
  xor g_113225_(out[36], out[740], _054814_);
  xor g_113226_(out[46], out[750], _054815_);
  or g_113227_(_054814_, _054815_, _054816_);
  xor g_113228_(out[45], out[749], _054817_);
  xor g_113229_(out[35], out[739], _054818_);
  xor g_113230_(out[32], out[736], _054819_);
  and g_113231_(_098096_, out[747], _054820_);
  xor g_113232_(out[42], out[746], _054821_);
  xor g_113233_(out[47], out[751], _054822_);
  xor g_113234_(out[38], out[742], _054824_);
  xor g_113235_(out[37], out[741], _054825_);
  xor g_113236_(out[40], out[744], _054826_);
  or g_113237_(_054817_, _054826_, _054827_);
  xor g_113238_(out[34], out[738], _054828_);
  xor g_113239_(out[41], out[745], _054829_);
  xor g_113240_(out[33], out[737], _054830_);
  or g_113241_(_054821_, _054828_, _054831_);
  or g_113242_(_054827_, _054831_, _054832_);
  or g_113243_(_054818_, _054829_, _054833_);
  or g_113244_(_054825_, _054833_, _054835_);
  or g_113245_(_054832_, _054835_, _054836_);
  or g_113246_(_054816_, _054836_, _054837_);
  xor g_113247_(out[44], out[748], _054838_);
  or g_113248_(_054820_, _054838_, _054839_);
  xor g_113249_(out[39], out[743], _054840_);
  or g_113250_(_054824_, _054840_, _054841_);
  or g_113251_(_054839_, _054841_, _054842_);
  or g_113252_(_054813_, _054830_, _054843_);
  or g_113253_(_054822_, _054843_, _054844_);
  or g_113254_(_054842_, _054844_, _054846_);
  or g_113255_(_054819_, _054846_, _054847_);
  or g_113256_(_054837_, _054847_, _054848_);
  xor g_113257_(out[23], out[743], _054849_);
  and g_113258_(_098063_, out[747], _054850_);
  xor g_113259_(out[30], out[750], _054851_);
  xor g_113260_(out[24], out[744], _054852_);
  xor g_113261_(out[17], out[737], _054853_);
  xor g_113262_(out[29], out[749], _054854_);
  xor g_113263_(out[25], out[745], _054855_);
  xor g_113264_(out[20], out[740], _054857_);
  xor g_113265_(out[18], out[738], _054858_);
  and g_113266_(out[27], _049675_, _054859_);
  xor g_113267_(out[19], out[739], _054860_);
  xor g_113268_(out[22], out[742], _054861_);
  xor g_113269_(out[31], out[751], _054862_);
  xor g_113270_(out[26], out[746], _054863_);
  xor g_113271_(out[21], out[741], _054864_);
  xor g_113272_(out[16], out[736], _054865_);
  or g_113273_(_054851_, _054857_, _054866_);
  or g_113274_(_054852_, _054854_, _054868_);
  or g_113275_(_054858_, _054863_, _054869_);
  or g_113276_(_054868_, _054869_, _054870_);
  or g_113277_(_054855_, _054860_, _054871_);
  or g_113278_(_054864_, _054865_, _054872_);
  or g_113279_(_054871_, _054872_, _054873_);
  or g_113280_(_054870_, _054873_, _054874_);
  xor g_113281_(out[28], out[748], _054875_);
  or g_113282_(_054850_, _054875_, _054876_);
  or g_113283_(_054849_, _054861_, _054877_);
  or g_113284_(_054876_, _054877_, _054879_);
  or g_113285_(_054853_, _054859_, _054880_);
  or g_113286_(_054862_, _054880_, _054881_);
  or g_113287_(_054879_, _054881_, _054882_);
  or g_113288_(_054874_, _054882_, _054883_);
  or g_113289_(_054866_, _054883_, _054884_);
  not g_113290_(_054884_, _054885_);
  xor g_113291_(out[10], out[746], _054886_);
  xor g_113292_(out[2], out[738], _054887_);
  xor g_113293_(out[1], out[737], _054888_);
  and g_113294_(_098041_, out[747], _054890_);
  and g_113295_(out[11], _049675_, _054891_);
  xor g_113296_(out[13], out[749], _054892_);
  xor g_113297_(out[3], out[739], _054893_);
  xor g_113298_(out[14], out[750], _054894_);
  xor g_113299_(out[12], out[748], _054895_);
  xor g_113300_(out[8], out[744], _054896_);
  xor g_113301_(out[15], out[751], _054897_);
  xor g_113302_(out[5], out[741], _054898_);
  xor g_113303_(out[6], out[742], _054899_);
  xor g_113304_(out[0], out[736], _054901_);
  xor g_113305_(out[4], out[740], _054902_);
  or g_113306_(_054892_, _054896_, _054903_);
  xor g_113307_(out[9], out[745], _054904_);
  or g_113308_(_054886_, _054887_, _054905_);
  or g_113309_(_054903_, _054905_, _054906_);
  or g_113310_(_054893_, _054904_, _054907_);
  or g_113311_(_054898_, _054907_, _054908_);
  or g_113312_(_054906_, _054908_, _054909_);
  or g_113313_(_054894_, _054902_, _054910_);
  or g_113314_(_054909_, _054910_, _054912_);
  or g_113315_(_054890_, _054895_, _054913_);
  xor g_113316_(out[7], out[743], _054914_);
  or g_113317_(_054899_, _054914_, _054915_);
  or g_113318_(_054913_, _054915_, _054916_);
  or g_113319_(_054888_, _054891_, _054917_);
  or g_113320_(_054897_, _054917_, _054918_);
  or g_113321_(_054916_, _054918_, _054919_);
  or g_113322_(_054901_, _054919_, _054920_);
  or g_113323_(_054912_, _054920_, _054921_);
  xor g_113324_(out[465], out[721], _054923_);
  and g_113325_(out[475], _049664_, _054924_);
  xor g_113326_(out[473], out[729], _054925_);
  xor g_113327_(out[464], out[720], _054926_);
  xor g_113328_(out[478], out[734], _054927_);
  xor g_113329_(out[468], out[724], _054928_);
  or g_113330_(_054927_, _054928_, _054929_);
  xor g_113331_(out[477], out[733], _054930_);
  xor g_113332_(out[467], out[723], _054931_);
  and g_113333_(_049499_, out[731], _054932_);
  xor g_113334_(out[470], out[726], _054934_);
  xor g_113335_(out[474], out[730], _054935_);
  xor g_113336_(out[469], out[725], _054936_);
  xor g_113337_(out[479], out[735], _054937_);
  xor g_113338_(out[472], out[728], _054938_);
  or g_113339_(_054930_, _054938_, _054939_);
  xor g_113340_(out[466], out[722], _054940_);
  or g_113341_(_054935_, _054940_, _054941_);
  or g_113342_(_054939_, _054941_, _054942_);
  or g_113343_(_054925_, _054931_, _054943_);
  or g_113344_(_054936_, _054943_, _054945_);
  or g_113345_(_054942_, _054945_, _054946_);
  or g_113346_(_054929_, _054946_, _054947_);
  xor g_113347_(out[476], out[732], _054948_);
  or g_113348_(_054932_, _054948_, _054949_);
  xor g_113349_(out[471], out[727], _054950_);
  or g_113350_(_054934_, _054950_, _054951_);
  or g_113351_(_054949_, _054951_, _054952_);
  or g_113352_(_054923_, _054924_, _054953_);
  or g_113353_(_054937_, _054953_, _054954_);
  or g_113354_(_054952_, _054954_, _054956_);
  or g_113355_(_054926_, _054956_, _054957_);
  or g_113356_(_054947_, _054957_, _054958_);
  xor g_113357_(out[455], out[727], _054959_);
  and g_113358_(_049477_, out[731], _054960_);
  xor g_113359_(out[462], out[734], _054961_);
  xor g_113360_(out[456], out[728], _054962_);
  xor g_113361_(out[449], out[721], _054963_);
  xor g_113362_(out[461], out[733], _054964_);
  xor g_113363_(out[457], out[729], _054965_);
  xor g_113364_(out[452], out[724], _054967_);
  xor g_113365_(out[450], out[722], _054968_);
  and g_113366_(out[459], _049664_, _054969_);
  xor g_113367_(out[451], out[723], _054970_);
  xor g_113368_(out[454], out[726], _054971_);
  xor g_113369_(out[463], out[735], _054972_);
  xor g_113370_(out[458], out[730], _054973_);
  xor g_113371_(out[453], out[725], _054974_);
  xor g_113372_(out[448], out[720], _054975_);
  or g_113373_(_054961_, _054967_, _054976_);
  or g_113374_(_054962_, _054964_, _054978_);
  or g_113375_(_054968_, _054973_, _054979_);
  or g_113376_(_054978_, _054979_, _054980_);
  or g_113377_(_054965_, _054970_, _054981_);
  or g_113378_(_054974_, _054975_, _054982_);
  or g_113379_(_054981_, _054982_, _054983_);
  or g_113380_(_054980_, _054983_, _054984_);
  xor g_113381_(out[460], out[732], _054985_);
  or g_113382_(_054960_, _054985_, _054986_);
  or g_113383_(_054959_, _054971_, _054987_);
  or g_113384_(_054986_, _054987_, _054989_);
  or g_113385_(_054963_, _054969_, _054990_);
  or g_113386_(_054972_, _054990_, _054991_);
  or g_113387_(_054989_, _054991_, _054992_);
  or g_113388_(_054984_, _054992_, _054993_);
  or g_113389_(_054976_, _054993_, _054994_);
  and g_113390_(out[443], _049664_, _054995_);
  and g_113391_(_049466_, out[731], _054996_);
  xor g_113392_(out[436], out[724], _054997_);
  xor g_113393_(out[433], out[721], _054998_);
  xor g_113394_(out[437], out[725], _055000_);
  xor g_113395_(out[441], out[729], _055001_);
  xor g_113396_(out[445], out[733], _055002_);
  xor g_113397_(out[442], out[730], _055003_);
  xor g_113398_(out[438], out[726], _055004_);
  xor g_113399_(out[440], out[728], _055005_);
  or g_113400_(_055002_, _055005_, _055006_);
  xor g_113401_(out[434], out[722], _055007_);
  xor g_113402_(out[447], out[735], _055008_);
  xor g_113403_(out[435], out[723], _055009_);
  xor g_113404_(out[446], out[734], _055011_);
  xor g_113405_(out[432], out[720], _055012_);
  or g_113406_(_055003_, _055007_, _055013_);
  or g_113407_(_055006_, _055013_, _055014_);
  or g_113408_(_055001_, _055009_, _055015_);
  or g_113409_(_055000_, _055015_, _055016_);
  or g_113410_(_055014_, _055016_, _055017_);
  or g_113411_(_054997_, _055011_, _055018_);
  or g_113412_(_055017_, _055018_, _055019_);
  xor g_113413_(out[444], out[732], _055020_);
  or g_113414_(_054996_, _055020_, _055022_);
  xor g_113415_(out[439], out[727], _055023_);
  or g_113416_(_055004_, _055023_, _055024_);
  or g_113417_(_055022_, _055024_, _055025_);
  or g_113418_(_054995_, _054998_, _055026_);
  or g_113419_(_055008_, _055026_, _055027_);
  or g_113420_(_055025_, _055027_, _055028_);
  or g_113421_(_055012_, _055028_, _055029_);
  or g_113422_(_055019_, _055029_, _055030_);
  xor g_113423_(out[423], out[727], _055031_);
  and g_113424_(_049455_, out[731], _055033_);
  xor g_113425_(out[430], out[734], _055034_);
  xor g_113426_(out[424], out[728], _055035_);
  xor g_113427_(out[417], out[721], _055036_);
  xor g_113428_(out[429], out[733], _055037_);
  xor g_113429_(out[425], out[729], _055038_);
  xor g_113430_(out[420], out[724], _055039_);
  xor g_113431_(out[418], out[722], _055040_);
  and g_113432_(out[427], _049664_, _055041_);
  xor g_113433_(out[419], out[723], _055042_);
  xor g_113434_(out[422], out[726], _055044_);
  xor g_113435_(out[431], out[735], _055045_);
  xor g_113436_(out[426], out[730], _055046_);
  xor g_113437_(out[421], out[725], _055047_);
  xor g_113438_(out[416], out[720], _055048_);
  or g_113439_(_055034_, _055039_, _055049_);
  or g_113440_(_055035_, _055037_, _055050_);
  or g_113441_(_055040_, _055046_, _055051_);
  or g_113442_(_055050_, _055051_, _055052_);
  or g_113443_(_055038_, _055042_, _055053_);
  or g_113444_(_055047_, _055048_, _055055_);
  or g_113445_(_055053_, _055055_, _055056_);
  or g_113446_(_055052_, _055056_, _055057_);
  xor g_113447_(out[428], out[732], _055058_);
  or g_113448_(_055033_, _055058_, _055059_);
  or g_113449_(_055031_, _055044_, _055060_);
  or g_113450_(_055059_, _055060_, _055061_);
  or g_113451_(_055036_, _055041_, _055062_);
  or g_113452_(_055045_, _055062_, _055063_);
  or g_113453_(_055061_, _055063_, _055064_);
  or g_113454_(_055057_, _055064_, _055066_);
  or g_113455_(_055049_, _055066_, _055067_);
  xor g_113456_(out[408], out[728], _055068_);
  xor g_113457_(out[405], out[725], _055069_);
  xor g_113458_(out[403], out[723], _055070_);
  xor g_113459_(out[414], out[734], _055071_);
  xor g_113460_(out[413], out[733], _055072_);
  xor g_113461_(out[402], out[722], _055073_);
  xor g_113462_(out[409], out[729], _055074_);
  xor g_113463_(out[406], out[726], _055075_);
  xor g_113464_(out[415], out[735], _055077_);
  xor g_113465_(out[410], out[730], _055078_);
  xor g_113466_(out[404], out[724], _055079_);
  xor g_113467_(out[400], out[720], _055080_);
  and g_113468_(_049444_, out[731], _055081_);
  and g_113469_(out[411], _049664_, _055082_);
  or g_113470_(_055068_, _055072_, _055083_);
  xor g_113471_(out[401], out[721], _055084_);
  or g_113472_(_055073_, _055078_, _055085_);
  or g_113473_(_055083_, _055085_, _055086_);
  or g_113474_(_055070_, _055074_, _055088_);
  or g_113475_(_055069_, _055088_, _055089_);
  or g_113476_(_055086_, _055089_, _055090_);
  or g_113477_(_055071_, _055079_, _055091_);
  or g_113478_(_055090_, _055091_, _055092_);
  xor g_113479_(out[412], out[732], _055093_);
  or g_113480_(_055081_, _055093_, _055094_);
  xor g_113481_(out[407], out[727], _055095_);
  or g_113482_(_055075_, _055095_, _055096_);
  or g_113483_(_055094_, _055096_, _055097_);
  or g_113484_(_055082_, _055084_, _055099_);
  or g_113485_(_055077_, _055099_, _055100_);
  or g_113486_(_055097_, _055100_, _055101_);
  or g_113487_(_055080_, _055101_, _055102_);
  or g_113488_(_055092_, _055102_, _055103_);
  xor g_113489_(out[391], out[727], _055104_);
  and g_113490_(_049433_, out[731], _055105_);
  xor g_113491_(out[398], out[734], _055106_);
  xor g_113492_(out[392], out[728], _055107_);
  xor g_113493_(out[385], out[721], _055108_);
  xor g_113494_(out[397], out[733], _055110_);
  xor g_113495_(out[393], out[729], _055111_);
  xor g_113496_(out[388], out[724], _055112_);
  xor g_113497_(out[386], out[722], _055113_);
  and g_113498_(out[395], _049664_, _055114_);
  xor g_113499_(out[387], out[723], _055115_);
  xor g_113500_(out[390], out[726], _055116_);
  xor g_113501_(out[399], out[735], _055117_);
  xor g_113502_(out[394], out[730], _055118_);
  xor g_113503_(out[389], out[725], _055119_);
  xor g_113504_(out[384], out[720], _055121_);
  or g_113505_(_055106_, _055112_, _055122_);
  or g_113506_(_055107_, _055110_, _055123_);
  or g_113507_(_055113_, _055118_, _055124_);
  or g_113508_(_055123_, _055124_, _055125_);
  or g_113509_(_055111_, _055115_, _055126_);
  or g_113510_(_055119_, _055121_, _055127_);
  or g_113511_(_055126_, _055127_, _055128_);
  or g_113512_(_055125_, _055128_, _055129_);
  xor g_113513_(out[396], out[732], _055130_);
  or g_113514_(_055105_, _055130_, _055132_);
  or g_113515_(_055104_, _055116_, _055133_);
  or g_113516_(_055132_, _055133_, _055134_);
  or g_113517_(_055108_, _055114_, _055135_);
  or g_113518_(_055117_, _055135_, _055136_);
  or g_113519_(_055134_, _055136_, _055137_);
  or g_113520_(_055129_, _055137_, _055138_);
  or g_113521_(_055122_, _055138_, _055139_);
  and g_113522_(_049422_, out[731], _055140_);
  and g_113523_(out[379], _049664_, _055141_);
  xor g_113524_(out[377], out[729], _055143_);
  xor g_113525_(out[371], out[723], _055144_);
  or g_113526_(_055143_, _055144_, _055145_);
  xor g_113527_(out[378], out[730], _055146_);
  xor g_113528_(out[383], out[735], _055147_);
  xor g_113529_(out[376], out[728], _055148_);
  xor g_113530_(out[370], out[722], _055149_);
  xor g_113531_(out[382], out[734], _055150_);
  xor g_113532_(out[369], out[721], _055151_);
  xor g_113533_(out[373], out[725], _055152_);
  xor g_113534_(out[374], out[726], _055154_);
  xor g_113535_(out[368], out[720], _055155_);
  xor g_113536_(out[372], out[724], _055156_);
  xor g_113537_(out[381], out[733], _055157_);
  or g_113538_(_055150_, _055156_, _055158_);
  or g_113539_(_055148_, _055157_, _055159_);
  or g_113540_(_055146_, _055149_, _055160_);
  or g_113541_(_055159_, _055160_, _055161_);
  or g_113542_(_055152_, _055155_, _055162_);
  or g_113543_(_055145_, _055162_, _055163_);
  or g_113544_(_055161_, _055163_, _055165_);
  xor g_113545_(out[380], out[732], _055166_);
  or g_113546_(_055140_, _055166_, _055167_);
  xor g_113547_(out[375], out[727], _055168_);
  or g_113548_(_055154_, _055168_, _055169_);
  or g_113549_(_055167_, _055169_, _055170_);
  or g_113550_(_055141_, _055151_, _055171_);
  or g_113551_(_055147_, _055171_, _055172_);
  or g_113552_(_055170_, _055172_, _055173_);
  or g_113553_(_055165_, _055173_, _055174_);
  or g_113554_(_055158_, _055174_, _055176_);
  xor g_113555_(out[359], out[727], _055177_);
  and g_113556_(_049411_, out[731], _055178_);
  xor g_113557_(out[366], out[734], _055179_);
  xor g_113558_(out[360], out[728], _055180_);
  xor g_113559_(out[353], out[721], _055181_);
  xor g_113560_(out[365], out[733], _055182_);
  xor g_113561_(out[361], out[729], _055183_);
  xor g_113562_(out[356], out[724], _055184_);
  xor g_113563_(out[354], out[722], _055185_);
  and g_113564_(out[363], _049664_, _055187_);
  xor g_113565_(out[355], out[723], _055188_);
  xor g_113566_(out[358], out[726], _055189_);
  xor g_113567_(out[367], out[735], _055190_);
  xor g_113568_(out[362], out[730], _055191_);
  xor g_113569_(out[357], out[725], _055192_);
  xor g_113570_(out[352], out[720], _055193_);
  or g_113571_(_055179_, _055184_, _055194_);
  or g_113572_(_055180_, _055182_, _055195_);
  or g_113573_(_055185_, _055191_, _055196_);
  or g_113574_(_055195_, _055196_, _055198_);
  or g_113575_(_055183_, _055188_, _055199_);
  or g_113576_(_055192_, _055193_, _055200_);
  or g_113577_(_055199_, _055200_, _055201_);
  or g_113578_(_055198_, _055201_, _055202_);
  xor g_113579_(out[364], out[732], _055203_);
  or g_113580_(_055178_, _055203_, _055204_);
  or g_113581_(_055177_, _055189_, _055205_);
  or g_113582_(_055204_, _055205_, _055206_);
  or g_113583_(_055181_, _055187_, _055207_);
  or g_113584_(_055190_, _055207_, _055209_);
  or g_113585_(_055206_, _055209_, _055210_);
  or g_113586_(_055202_, _055210_, _055211_);
  or g_113587_(_055194_, _055211_, _055212_);
  and g_113588_(_049400_, out[731], _055213_);
  and g_113589_(out[347], _049664_, _055214_);
  xor g_113590_(out[340], out[724], _055215_);
  xor g_113591_(out[350], out[734], _055216_);
  or g_113592_(_055215_, _055216_, _055217_);
  xor g_113593_(out[349], out[733], _055218_);
  xor g_113594_(out[339], out[723], _055220_);
  xor g_113595_(out[336], out[720], _055221_);
  xor g_113596_(out[346], out[730], _055222_);
  xor g_113597_(out[351], out[735], _055223_);
  xor g_113598_(out[342], out[726], _055224_);
  xor g_113599_(out[341], out[725], _055225_);
  xor g_113600_(out[344], out[728], _055226_);
  or g_113601_(_055218_, _055226_, _055227_);
  xor g_113602_(out[338], out[722], _055228_);
  xor g_113603_(out[345], out[729], _055229_);
  xor g_113604_(out[337], out[721], _055231_);
  or g_113605_(_055222_, _055228_, _055232_);
  or g_113606_(_055227_, _055232_, _055233_);
  or g_113607_(_055220_, _055229_, _055234_);
  or g_113608_(_055225_, _055234_, _055235_);
  or g_113609_(_055233_, _055235_, _055236_);
  or g_113610_(_055217_, _055236_, _055237_);
  xor g_113611_(out[348], out[732], _055238_);
  or g_113612_(_055213_, _055238_, _055239_);
  xor g_113613_(out[343], out[727], _055240_);
  or g_113614_(_055224_, _055240_, _055242_);
  or g_113615_(_055239_, _055242_, _055243_);
  or g_113616_(_055214_, _055231_, _055244_);
  or g_113617_(_055223_, _055244_, _055245_);
  or g_113618_(_055243_, _055245_, _055246_);
  or g_113619_(_055221_, _055246_, _055247_);
  or g_113620_(_055237_, _055247_, _055248_);
  xor g_113621_(out[327], out[727], _055249_);
  and g_113622_(_098294_, out[731], _055250_);
  xor g_113623_(out[334], out[734], _055251_);
  xor g_113624_(out[328], out[728], _055253_);
  xor g_113625_(out[321], out[721], _055254_);
  xor g_113626_(out[333], out[733], _055255_);
  xor g_113627_(out[329], out[729], _055256_);
  xor g_113628_(out[324], out[724], _055257_);
  xor g_113629_(out[322], out[722], _055258_);
  and g_113630_(out[331], _049664_, _055259_);
  xor g_113631_(out[323], out[723], _055260_);
  xor g_113632_(out[326], out[726], _055261_);
  xor g_113633_(out[335], out[735], _055262_);
  xor g_113634_(out[330], out[730], _055264_);
  xor g_113635_(out[325], out[725], _055265_);
  xor g_113636_(out[320], out[720], _055266_);
  or g_113637_(_055251_, _055257_, _055267_);
  or g_113638_(_055253_, _055255_, _055268_);
  or g_113639_(_055258_, _055264_, _055269_);
  or g_113640_(_055268_, _055269_, _055270_);
  or g_113641_(_055256_, _055260_, _055271_);
  or g_113642_(_055265_, _055266_, _055272_);
  or g_113643_(_055271_, _055272_, _055273_);
  or g_113644_(_055270_, _055273_, _055275_);
  xor g_113645_(out[332], out[732], _055276_);
  or g_113646_(_055250_, _055276_, _055277_);
  or g_113647_(_055249_, _055261_, _055278_);
  or g_113648_(_055277_, _055278_, _055279_);
  or g_113649_(_055254_, _055259_, _055280_);
  or g_113650_(_055262_, _055280_, _055281_);
  or g_113651_(_055279_, _055281_, _055282_);
  or g_113652_(_055275_, _055282_, _055283_);
  or g_113653_(_055267_, _055283_, _055284_);
  xor g_113654_(out[312], out[728], _055286_);
  xor g_113655_(out[309], out[725], _055287_);
  xor g_113656_(out[307], out[723], _055288_);
  xor g_113657_(out[318], out[734], _055289_);
  xor g_113658_(out[317], out[733], _055290_);
  xor g_113659_(out[306], out[722], _055291_);
  xor g_113660_(out[313], out[729], _055292_);
  xor g_113661_(out[310], out[726], _055293_);
  xor g_113662_(out[319], out[735], _055294_);
  xor g_113663_(out[314], out[730], _055295_);
  xor g_113664_(out[308], out[724], _055297_);
  xor g_113665_(out[304], out[720], _055298_);
  and g_113666_(_098283_, out[731], _055299_);
  and g_113667_(out[315], _049664_, _055300_);
  or g_113668_(_055286_, _055290_, _055301_);
  xor g_113669_(out[305], out[721], _055302_);
  or g_113670_(_055291_, _055295_, _055303_);
  or g_113671_(_055301_, _055303_, _055304_);
  or g_113672_(_055288_, _055292_, _055305_);
  or g_113673_(_055287_, _055305_, _055306_);
  or g_113674_(_055304_, _055306_, _055308_);
  or g_113675_(_055289_, _055297_, _055309_);
  or g_113676_(_055308_, _055309_, _055310_);
  xor g_113677_(out[316], out[732], _055311_);
  or g_113678_(_055299_, _055311_, _055312_);
  xor g_113679_(out[311], out[727], _055313_);
  or g_113680_(_055293_, _055313_, _055314_);
  or g_113681_(_055312_, _055314_, _055315_);
  or g_113682_(_055300_, _055302_, _055316_);
  or g_113683_(_055294_, _055316_, _055317_);
  or g_113684_(_055315_, _055317_, _055319_);
  or g_113685_(_055298_, _055319_, _055320_);
  or g_113686_(_055310_, _055320_, _055321_);
  not g_113687_(_055321_, _055322_);
  xor g_113688_(out[295], out[727], _055323_);
  and g_113689_(_098272_, out[731], _055324_);
  xor g_113690_(out[302], out[734], _055325_);
  xor g_113691_(out[296], out[728], _055326_);
  xor g_113692_(out[289], out[721], _055327_);
  xor g_113693_(out[301], out[733], _055328_);
  xor g_113694_(out[297], out[729], _055330_);
  xor g_113695_(out[292], out[724], _055331_);
  xor g_113696_(out[290], out[722], _055332_);
  and g_113697_(out[299], _049664_, _055333_);
  xor g_113698_(out[291], out[723], _055334_);
  xor g_113699_(out[294], out[726], _055335_);
  xor g_113700_(out[303], out[735], _055336_);
  xor g_113701_(out[298], out[730], _055337_);
  xor g_113702_(out[293], out[725], _055338_);
  xor g_113703_(out[288], out[720], _055339_);
  or g_113704_(_055325_, _055331_, _055341_);
  or g_113705_(_055326_, _055328_, _055342_);
  or g_113706_(_055332_, _055337_, _055343_);
  or g_113707_(_055342_, _055343_, _055344_);
  or g_113708_(_055330_, _055334_, _055345_);
  or g_113709_(_055338_, _055339_, _055346_);
  or g_113710_(_055345_, _055346_, _055347_);
  or g_113711_(_055344_, _055347_, _055348_);
  xor g_113712_(out[300], out[732], _055349_);
  or g_113713_(_055324_, _055349_, _055350_);
  or g_113714_(_055323_, _055335_, _055352_);
  or g_113715_(_055350_, _055352_, _055353_);
  or g_113716_(_055327_, _055333_, _055354_);
  or g_113717_(_055336_, _055354_, _055355_);
  or g_113718_(_055353_, _055355_, _055356_);
  or g_113719_(_055348_, _055356_, _055357_);
  or g_113720_(_055341_, _055357_, _055358_);
  not g_113721_(_055358_, _055359_);
  and g_113722_(out[283], _049664_, _055360_);
  xor g_113723_(out[276], out[724], _055361_);
  xor g_113724_(out[286], out[734], _055363_);
  or g_113725_(_055361_, _055363_, _055364_);
  xor g_113726_(out[285], out[733], _055365_);
  xor g_113727_(out[275], out[723], _055366_);
  xor g_113728_(out[272], out[720], _055367_);
  and g_113729_(_098261_, out[731], _055368_);
  xor g_113730_(out[282], out[730], _055369_);
  xor g_113731_(out[287], out[735], _055370_);
  xor g_113732_(out[278], out[726], _055371_);
  xor g_113733_(out[277], out[725], _055372_);
  xor g_113734_(out[280], out[728], _055374_);
  or g_113735_(_055365_, _055374_, _055375_);
  xor g_113736_(out[274], out[722], _055376_);
  xor g_113737_(out[281], out[729], _055377_);
  xor g_113738_(out[273], out[721], _055378_);
  or g_113739_(_055369_, _055376_, _055379_);
  or g_113740_(_055375_, _055379_, _055380_);
  or g_113741_(_055366_, _055377_, _055381_);
  or g_113742_(_055372_, _055381_, _055382_);
  or g_113743_(_055380_, _055382_, _055383_);
  or g_113744_(_055364_, _055383_, _055385_);
  xor g_113745_(out[284], out[732], _055386_);
  or g_113746_(_055368_, _055386_, _055387_);
  xor g_113747_(out[279], out[727], _055388_);
  or g_113748_(_055371_, _055388_, _055389_);
  or g_113749_(_055387_, _055389_, _055390_);
  or g_113750_(_055360_, _055378_, _055391_);
  or g_113751_(_055370_, _055391_, _055392_);
  or g_113752_(_055390_, _055392_, _055393_);
  or g_113753_(_055367_, _055393_, _055394_);
  or g_113754_(_055385_, _055394_, _055396_);
  xor g_113755_(out[263], out[727], _055397_);
  and g_113756_(_098250_, out[731], _055398_);
  xor g_113757_(out[270], out[734], _055399_);
  xor g_113758_(out[264], out[728], _055400_);
  xor g_113759_(out[257], out[721], _055401_);
  xor g_113760_(out[269], out[733], _055402_);
  xor g_113761_(out[265], out[729], _055403_);
  xor g_113762_(out[260], out[724], _055404_);
  xor g_113763_(out[258], out[722], _055405_);
  and g_113764_(out[267], _049664_, _055407_);
  xor g_113765_(out[259], out[723], _055408_);
  xor g_113766_(out[262], out[726], _055409_);
  xor g_113767_(out[271], out[735], _055410_);
  xor g_113768_(out[266], out[730], _055411_);
  xor g_113769_(out[261], out[725], _055412_);
  xor g_113770_(out[256], out[720], _055413_);
  or g_113771_(_055399_, _055404_, _055414_);
  or g_113772_(_055400_, _055402_, _055415_);
  or g_113773_(_055405_, _055411_, _055416_);
  or g_113774_(_055415_, _055416_, _055418_);
  or g_113775_(_055403_, _055408_, _055419_);
  or g_113776_(_055412_, _055413_, _055420_);
  or g_113777_(_055419_, _055420_, _055421_);
  or g_113778_(_055418_, _055421_, _055422_);
  xor g_113779_(out[268], out[732], _055423_);
  or g_113780_(_055398_, _055423_, _055424_);
  or g_113781_(_055397_, _055409_, _055425_);
  or g_113782_(_055424_, _055425_, _055426_);
  or g_113783_(_055401_, _055407_, _055427_);
  or g_113784_(_055410_, _055427_, _055429_);
  or g_113785_(_055426_, _055429_, _055430_);
  or g_113786_(_055422_, _055430_, _055431_);
  or g_113787_(_055414_, _055431_, _055432_);
  xor g_113788_(out[253], out[733], _055433_);
  xor g_113789_(out[242], out[722], _055434_);
  xor g_113790_(out[245], out[725], _055435_);
  xor g_113791_(out[249], out[729], _055436_);
  xor g_113792_(out[244], out[724], _055437_);
  xor g_113793_(out[248], out[728], _055438_);
  xor g_113794_(out[254], out[734], _055440_);
  xor g_113795_(out[246], out[726], _055441_);
  xor g_113796_(out[255], out[735], _055442_);
  xor g_113797_(out[250], out[730], _055443_);
  xor g_113798_(out[240], out[720], _055444_);
  xor g_113799_(out[243], out[723], _055445_);
  and g_113800_(_098239_, out[731], _055446_);
  and g_113801_(out[251], _049664_, _055447_);
  xor g_113802_(out[241], out[721], _055448_);
  or g_113803_(_055437_, _055440_, _055449_);
  or g_113804_(_055433_, _055438_, _055451_);
  or g_113805_(_055434_, _055443_, _055452_);
  or g_113806_(_055451_, _055452_, _055453_);
  or g_113807_(_055436_, _055445_, _055454_);
  or g_113808_(_055435_, _055444_, _055455_);
  or g_113809_(_055454_, _055455_, _055456_);
  or g_113810_(_055453_, _055456_, _055457_);
  xor g_113811_(out[252], out[732], _055458_);
  or g_113812_(_055446_, _055458_, _055459_);
  xor g_113813_(out[247], out[727], _055460_);
  or g_113814_(_055441_, _055460_, _055462_);
  or g_113815_(_055459_, _055462_, _055463_);
  or g_113816_(_055447_, _055448_, _055464_);
  or g_113817_(_055442_, _055464_, _055465_);
  or g_113818_(_055463_, _055465_, _055466_);
  or g_113819_(_055457_, _055466_, _055467_);
  or g_113820_(_055449_, _055467_, _055468_);
  not g_113821_(_055468_, _055469_);
  xor g_113822_(out[231], out[727], _055470_);
  and g_113823_(_098228_, out[731], _055471_);
  xor g_113824_(out[238], out[734], _055473_);
  xor g_113825_(out[232], out[728], _055474_);
  xor g_113826_(out[225], out[721], _055475_);
  xor g_113827_(out[237], out[733], _055476_);
  xor g_113828_(out[233], out[729], _055477_);
  xor g_113829_(out[228], out[724], _055478_);
  xor g_113830_(out[226], out[722], _055479_);
  and g_113831_(out[235], _049664_, _055480_);
  xor g_113832_(out[227], out[723], _055481_);
  xor g_113833_(out[230], out[726], _055482_);
  xor g_113834_(out[239], out[735], _055484_);
  xor g_113835_(out[234], out[730], _055485_);
  xor g_113836_(out[229], out[725], _055486_);
  xor g_113837_(out[224], out[720], _055487_);
  or g_113838_(_055473_, _055478_, _055488_);
  or g_113839_(_055474_, _055476_, _055489_);
  or g_113840_(_055479_, _055485_, _055490_);
  or g_113841_(_055489_, _055490_, _055491_);
  or g_113842_(_055477_, _055481_, _055492_);
  or g_113843_(_055486_, _055487_, _055493_);
  or g_113844_(_055492_, _055493_, _055495_);
  or g_113845_(_055491_, _055495_, _055496_);
  xor g_113846_(out[236], out[732], _055497_);
  or g_113847_(_055471_, _055497_, _055498_);
  or g_113848_(_055470_, _055482_, _055499_);
  or g_113849_(_055498_, _055499_, _055500_);
  or g_113850_(_055475_, _055480_, _055501_);
  or g_113851_(_055484_, _055501_, _055502_);
  or g_113852_(_055500_, _055502_, _055503_);
  or g_113853_(_055496_, _055503_, _055504_);
  or g_113854_(_055488_, _055504_, _055506_);
  not g_113855_(_055506_, _055507_);
  xor g_113856_(out[209], out[721], _055508_);
  and g_113857_(out[219], _049664_, _055509_);
  xor g_113858_(out[217], out[729], _055510_);
  xor g_113859_(out[208], out[720], _055511_);
  xor g_113860_(out[222], out[734], _055512_);
  xor g_113861_(out[212], out[724], _055513_);
  or g_113862_(_055512_, _055513_, _055514_);
  xor g_113863_(out[221], out[733], _055515_);
  xor g_113864_(out[211], out[723], _055517_);
  and g_113865_(_098217_, out[731], _055518_);
  xor g_113866_(out[214], out[726], _055519_);
  xor g_113867_(out[218], out[730], _055520_);
  xor g_113868_(out[213], out[725], _055521_);
  xor g_113869_(out[223], out[735], _055522_);
  xor g_113870_(out[216], out[728], _055523_);
  or g_113871_(_055515_, _055523_, _055524_);
  xor g_113872_(out[210], out[722], _055525_);
  or g_113873_(_055520_, _055525_, _055526_);
  or g_113874_(_055524_, _055526_, _055528_);
  or g_113875_(_055510_, _055517_, _055529_);
  or g_113876_(_055521_, _055529_, _055530_);
  or g_113877_(_055528_, _055530_, _055531_);
  or g_113878_(_055514_, _055531_, _055532_);
  xor g_113879_(out[220], out[732], _055533_);
  or g_113880_(_055518_, _055533_, _055534_);
  xor g_113881_(out[215], out[727], _055535_);
  or g_113882_(_055519_, _055535_, _055536_);
  or g_113883_(_055534_, _055536_, _055537_);
  or g_113884_(_055508_, _055509_, _055539_);
  or g_113885_(_055522_, _055539_, _055540_);
  or g_113886_(_055537_, _055540_, _055541_);
  or g_113887_(_055511_, _055541_, _055542_);
  or g_113888_(_055532_, _055542_, _055543_);
  xor g_113889_(out[199], out[727], _055544_);
  and g_113890_(_098206_, out[731], _055545_);
  xor g_113891_(out[206], out[734], _055546_);
  xor g_113892_(out[200], out[728], _055547_);
  xor g_113893_(out[193], out[721], _055548_);
  xor g_113894_(out[205], out[733], _055550_);
  xor g_113895_(out[201], out[729], _055551_);
  xor g_113896_(out[196], out[724], _055552_);
  xor g_113897_(out[194], out[722], _055553_);
  and g_113898_(out[203], _049664_, _055554_);
  xor g_113899_(out[195], out[723], _055555_);
  xor g_113900_(out[198], out[726], _055556_);
  xor g_113901_(out[207], out[735], _055557_);
  xor g_113902_(out[202], out[730], _055558_);
  xor g_113903_(out[197], out[725], _055559_);
  xor g_113904_(out[192], out[720], _055561_);
  or g_113905_(_055546_, _055552_, _055562_);
  or g_113906_(_055547_, _055550_, _055563_);
  or g_113907_(_055553_, _055558_, _055564_);
  or g_113908_(_055563_, _055564_, _055565_);
  or g_113909_(_055551_, _055555_, _055566_);
  or g_113910_(_055559_, _055561_, _055567_);
  or g_113911_(_055566_, _055567_, _055568_);
  or g_113912_(_055565_, _055568_, _055569_);
  xor g_113913_(out[204], out[732], _055570_);
  or g_113914_(_055545_, _055570_, _055572_);
  or g_113915_(_055544_, _055556_, _055573_);
  or g_113916_(_055572_, _055573_, _055574_);
  or g_113917_(_055548_, _055554_, _055575_);
  or g_113918_(_055557_, _055575_, _055576_);
  or g_113919_(_055574_, _055576_, _055577_);
  or g_113920_(_055569_, _055577_, _055578_);
  or g_113921_(_055562_, _055578_, _055579_);
  xor g_113922_(out[177], out[721], _055580_);
  and g_113923_(out[187], _049664_, _055581_);
  xor g_113924_(out[185], out[729], _055583_);
  xor g_113925_(out[176], out[720], _055584_);
  xor g_113926_(out[190], out[734], _055585_);
  xor g_113927_(out[180], out[724], _055586_);
  or g_113928_(_055585_, _055586_, _055587_);
  xor g_113929_(out[189], out[733], _055588_);
  xor g_113930_(out[179], out[723], _055589_);
  and g_113931_(_098195_, out[731], _055590_);
  xor g_113932_(out[182], out[726], _055591_);
  xor g_113933_(out[186], out[730], _055592_);
  xor g_113934_(out[181], out[725], _055594_);
  xor g_113935_(out[191], out[735], _055595_);
  xor g_113936_(out[184], out[728], _055596_);
  or g_113937_(_055588_, _055596_, _055597_);
  xor g_113938_(out[178], out[722], _055598_);
  or g_113939_(_055592_, _055598_, _055599_);
  or g_113940_(_055597_, _055599_, _055600_);
  or g_113941_(_055583_, _055589_, _055601_);
  or g_113942_(_055594_, _055601_, _055602_);
  or g_113943_(_055600_, _055602_, _055603_);
  or g_113944_(_055587_, _055603_, _055605_);
  xor g_113945_(out[188], out[732], _055606_);
  or g_113946_(_055590_, _055606_, _055607_);
  xor g_113947_(out[183], out[727], _055608_);
  or g_113948_(_055591_, _055608_, _055609_);
  or g_113949_(_055607_, _055609_, _055610_);
  or g_113950_(_055580_, _055581_, _055611_);
  or g_113951_(_055595_, _055611_, _055612_);
  or g_113952_(_055610_, _055612_, _055613_);
  or g_113953_(_055584_, _055613_, _055614_);
  or g_113954_(_055605_, _055614_, _055616_);
  xor g_113955_(out[167], out[727], _055617_);
  and g_113956_(_098184_, out[731], _055618_);
  xor g_113957_(out[174], out[734], _055619_);
  xor g_113958_(out[168], out[728], _055620_);
  xor g_113959_(out[161], out[721], _055621_);
  xor g_113960_(out[173], out[733], _055622_);
  xor g_113961_(out[169], out[729], _055623_);
  xor g_113962_(out[164], out[724], _055624_);
  xor g_113963_(out[162], out[722], _055625_);
  and g_113964_(out[171], _049664_, _055627_);
  xor g_113965_(out[163], out[723], _055628_);
  xor g_113966_(out[166], out[726], _055629_);
  xor g_113967_(out[175], out[735], _055630_);
  xor g_113968_(out[170], out[730], _055631_);
  xor g_113969_(out[165], out[725], _055632_);
  xor g_113970_(out[160], out[720], _055633_);
  or g_113971_(_055619_, _055624_, _055634_);
  or g_113972_(_055620_, _055622_, _055635_);
  or g_113973_(_055625_, _055631_, _055636_);
  or g_113974_(_055635_, _055636_, _055638_);
  or g_113975_(_055623_, _055628_, _055639_);
  or g_113976_(_055632_, _055633_, _055640_);
  or g_113977_(_055639_, _055640_, _055641_);
  or g_113978_(_055638_, _055641_, _055642_);
  xor g_113979_(out[172], out[732], _055643_);
  or g_113980_(_055618_, _055643_, _055644_);
  or g_113981_(_055617_, _055629_, _055645_);
  or g_113982_(_055644_, _055645_, _055646_);
  or g_113983_(_055621_, _055627_, _055647_);
  or g_113984_(_055630_, _055647_, _055649_);
  or g_113985_(_055646_, _055649_, _055650_);
  or g_113986_(_055642_, _055650_, _055651_);
  or g_113987_(_055634_, _055651_, _055652_);
  and g_113988_(out[155], _049664_, _055653_);
  xor g_113989_(out[148], out[724], _055654_);
  xor g_113990_(out[158], out[734], _055655_);
  or g_113991_(_055654_, _055655_, _055656_);
  xor g_113992_(out[157], out[733], _055657_);
  xor g_113993_(out[147], out[723], _055658_);
  xor g_113994_(out[144], out[720], _055660_);
  and g_113995_(_098173_, out[731], _055661_);
  xor g_113996_(out[154], out[730], _055662_);
  xor g_113997_(out[159], out[735], _055663_);
  xor g_113998_(out[150], out[726], _055664_);
  xor g_113999_(out[149], out[725], _055665_);
  xor g_114000_(out[152], out[728], _055666_);
  or g_114001_(_055657_, _055666_, _055667_);
  xor g_114002_(out[146], out[722], _055668_);
  xor g_114003_(out[153], out[729], _055669_);
  xor g_114004_(out[145], out[721], _055671_);
  or g_114005_(_055662_, _055668_, _055672_);
  or g_114006_(_055667_, _055672_, _055673_);
  or g_114007_(_055658_, _055669_, _055674_);
  or g_114008_(_055665_, _055674_, _055675_);
  or g_114009_(_055673_, _055675_, _055676_);
  or g_114010_(_055656_, _055676_, _055677_);
  xor g_114011_(out[156], out[732], _055678_);
  or g_114012_(_055661_, _055678_, _055679_);
  xor g_114013_(out[151], out[727], _055680_);
  or g_114014_(_055664_, _055680_, _055682_);
  or g_114015_(_055679_, _055682_, _055683_);
  or g_114016_(_055653_, _055671_, _055684_);
  or g_114017_(_055663_, _055684_, _055685_);
  or g_114018_(_055683_, _055685_, _055686_);
  or g_114019_(_055660_, _055686_, _055687_);
  or g_114020_(_055677_, _055687_, _055688_);
  xor g_114021_(out[135], out[727], _055689_);
  and g_114022_(_098162_, out[731], _055690_);
  xor g_114023_(out[142], out[734], _055691_);
  xor g_114024_(out[136], out[728], _055693_);
  xor g_114025_(out[129], out[721], _055694_);
  xor g_114026_(out[141], out[733], _055695_);
  xor g_114027_(out[137], out[729], _055696_);
  xor g_114028_(out[132], out[724], _055697_);
  xor g_114029_(out[130], out[722], _055698_);
  and g_114030_(out[139], _049664_, _055699_);
  xor g_114031_(out[131], out[723], _055700_);
  xor g_114032_(out[134], out[726], _055701_);
  xor g_114033_(out[143], out[735], _055702_);
  xor g_114034_(out[138], out[730], _055704_);
  xor g_114035_(out[133], out[725], _055705_);
  xor g_114036_(out[128], out[720], _055706_);
  or g_114037_(_055691_, _055697_, _055707_);
  or g_114038_(_055693_, _055695_, _055708_);
  or g_114039_(_055698_, _055704_, _055709_);
  or g_114040_(_055708_, _055709_, _055710_);
  or g_114041_(_055696_, _055700_, _055711_);
  or g_114042_(_055705_, _055706_, _055712_);
  or g_114043_(_055711_, _055712_, _055713_);
  or g_114044_(_055710_, _055713_, _055715_);
  xor g_114045_(out[140], out[732], _055716_);
  or g_114046_(_055690_, _055716_, _055717_);
  or g_114047_(_055689_, _055701_, _055718_);
  or g_114048_(_055717_, _055718_, _055719_);
  or g_114049_(_055694_, _055699_, _055720_);
  or g_114050_(_055702_, _055720_, _055721_);
  or g_114051_(_055719_, _055721_, _055722_);
  or g_114052_(_055715_, _055722_, _055723_);
  or g_114053_(_055707_, _055723_, _055724_);
  xor g_114054_(out[125], out[733], _055726_);
  xor g_114055_(out[122], out[730], _055727_);
  xor g_114056_(out[117], out[725], _055728_);
  and g_114057_(_098151_, out[731], _055729_);
  xor g_114058_(out[112], out[720], _055730_);
  and g_114059_(out[123], _049664_, _055731_);
  xor g_114060_(out[114], out[722], _055732_);
  xor g_114061_(out[115], out[723], _055733_);
  xor g_114062_(out[121], out[729], _055734_);
  xor g_114063_(out[113], out[721], _055735_);
  xor g_114064_(out[127], out[735], _055737_);
  xor g_114065_(out[126], out[734], _055738_);
  xor g_114066_(out[118], out[726], _055739_);
  xor g_114067_(out[116], out[724], _055740_);
  xor g_114068_(out[120], out[728], _055741_);
  or g_114069_(_055726_, _055741_, _055742_);
  or g_114070_(_055727_, _055732_, _055743_);
  or g_114071_(_055742_, _055743_, _055744_);
  or g_114072_(_055733_, _055734_, _055745_);
  or g_114073_(_055728_, _055745_, _055746_);
  or g_114074_(_055744_, _055746_, _055748_);
  or g_114075_(_055738_, _055740_, _055749_);
  or g_114076_(_055748_, _055749_, _055750_);
  xor g_114077_(out[124], out[732], _055751_);
  or g_114078_(_055729_, _055751_, _055752_);
  xor g_114079_(out[119], out[727], _055753_);
  or g_114080_(_055739_, _055753_, _055754_);
  or g_114081_(_055752_, _055754_, _055755_);
  or g_114082_(_055731_, _055735_, _055756_);
  or g_114083_(_055737_, _055756_, _055757_);
  or g_114084_(_055755_, _055757_, _055759_);
  or g_114085_(_055730_, _055759_, _055760_);
  or g_114086_(_055750_, _055760_, _055761_);
  xor g_114087_(out[103], out[727], _055762_);
  and g_114088_(_098140_, out[731], _055763_);
  xor g_114089_(out[110], out[734], _055764_);
  xor g_114090_(out[104], out[728], _055765_);
  xor g_114091_(out[97], out[721], _055766_);
  xor g_114092_(out[109], out[733], _055767_);
  xor g_114093_(out[105], out[729], _055768_);
  xor g_114094_(out[100], out[724], _055770_);
  xor g_114095_(out[98], out[722], _055771_);
  and g_114096_(out[107], _049664_, _055772_);
  xor g_114097_(out[99], out[723], _055773_);
  xor g_114098_(out[102], out[726], _055774_);
  xor g_114099_(out[111], out[735], _055775_);
  xor g_114100_(out[106], out[730], _055776_);
  xor g_114101_(out[101], out[725], _055777_);
  xor g_114102_(out[96], out[720], _055778_);
  or g_114103_(_055764_, _055770_, _055779_);
  or g_114104_(_055765_, _055767_, _055781_);
  or g_114105_(_055771_, _055776_, _055782_);
  or g_114106_(_055781_, _055782_, _055783_);
  or g_114107_(_055768_, _055773_, _055784_);
  or g_114108_(_055777_, _055778_, _055785_);
  or g_114109_(_055784_, _055785_, _055786_);
  or g_114110_(_055783_, _055786_, _055787_);
  xor g_114111_(out[108], out[732], _055788_);
  or g_114112_(_055763_, _055788_, _055789_);
  or g_114113_(_055762_, _055774_, _055790_);
  or g_114114_(_055789_, _055790_, _055792_);
  or g_114115_(_055766_, _055772_, _055793_);
  or g_114116_(_055775_, _055793_, _055794_);
  or g_114117_(_055792_, _055794_, _055795_);
  or g_114118_(_055787_, _055795_, _055796_);
  or g_114119_(_055779_, _055796_, _055797_);
  xor g_114120_(out[81], out[721], _055798_);
  and g_114121_(_098129_, out[731], _055799_);
  and g_114122_(out[91], _049664_, _055800_);
  xor g_114123_(out[89], out[729], _055801_);
  xor g_114124_(out[80], out[720], _055803_);
  xor g_114125_(out[94], out[734], _055804_);
  xor g_114126_(out[84], out[724], _055805_);
  or g_114127_(_055804_, _055805_, _055806_);
  xor g_114128_(out[93], out[733], _055807_);
  xor g_114129_(out[83], out[723], _055808_);
  xor g_114130_(out[92], out[732], _055809_);
  xor g_114131_(out[86], out[726], _055810_);
  xor g_114132_(out[90], out[730], _055811_);
  xor g_114133_(out[85], out[725], _055812_);
  xor g_114134_(out[95], out[735], _055814_);
  xor g_114135_(out[88], out[728], _055815_);
  or g_114136_(_055807_, _055815_, _055816_);
  xor g_114137_(out[82], out[722], _055817_);
  or g_114138_(_055811_, _055817_, _055818_);
  or g_114139_(_055816_, _055818_, _055819_);
  or g_114140_(_055801_, _055808_, _055820_);
  or g_114141_(_055812_, _055820_, _055821_);
  or g_114142_(_055819_, _055821_, _055822_);
  or g_114143_(_055806_, _055822_, _055823_);
  or g_114144_(_055799_, _055809_, _055825_);
  xor g_114145_(out[87], out[727], _055826_);
  or g_114146_(_055810_, _055826_, _055827_);
  or g_114147_(_055825_, _055827_, _055828_);
  or g_114148_(_055798_, _055800_, _055829_);
  or g_114149_(_055814_, _055829_, _055830_);
  or g_114150_(_055828_, _055830_, _055831_);
  or g_114151_(_055803_, _055831_, _055832_);
  or g_114152_(_055823_, _055832_, _055833_);
  xor g_114153_(out[71], out[727], _055834_);
  and g_114154_(_098118_, out[731], _055836_);
  xor g_114155_(out[78], out[734], _055837_);
  xor g_114156_(out[72], out[728], _055838_);
  xor g_114157_(out[65], out[721], _055839_);
  xor g_114158_(out[77], out[733], _055840_);
  xor g_114159_(out[73], out[729], _055841_);
  xor g_114160_(out[68], out[724], _055842_);
  xor g_114161_(out[66], out[722], _055843_);
  and g_114162_(out[75], _049664_, _055844_);
  xor g_114163_(out[67], out[723], _055845_);
  xor g_114164_(out[70], out[726], _055847_);
  xor g_114165_(out[79], out[735], _055848_);
  xor g_114166_(out[74], out[730], _055849_);
  xor g_114167_(out[69], out[725], _055850_);
  xor g_114168_(out[64], out[720], _055851_);
  or g_114169_(_055837_, _055842_, _055852_);
  or g_114170_(_055838_, _055840_, _055853_);
  or g_114171_(_055843_, _055849_, _055854_);
  or g_114172_(_055853_, _055854_, _055855_);
  or g_114173_(_055841_, _055845_, _055856_);
  or g_114174_(_055850_, _055851_, _055858_);
  or g_114175_(_055856_, _055858_, _055859_);
  or g_114176_(_055855_, _055859_, _055860_);
  xor g_114177_(out[76], out[732], _055861_);
  or g_114178_(_055836_, _055861_, _055862_);
  or g_114179_(_055834_, _055847_, _055863_);
  or g_114180_(_055862_, _055863_, _055864_);
  or g_114181_(_055839_, _055844_, _055865_);
  or g_114182_(_055848_, _055865_, _055866_);
  or g_114183_(_055864_, _055866_, _055867_);
  or g_114184_(_055860_, _055867_, _055869_);
  or g_114185_(_055852_, _055869_, _055870_);
  xor g_114186_(out[49], out[721], _055871_);
  and g_114187_(out[59], _049664_, _055872_);
  xor g_114188_(out[62], out[734], _055873_);
  xor g_114189_(out[51], out[723], _055874_);
  xor g_114190_(out[52], out[724], _055875_);
  xor g_114191_(out[50], out[722], _055876_);
  xor g_114192_(out[57], out[729], _055877_);
  xor g_114193_(out[48], out[720], _055878_);
  and g_114194_(_098107_, out[731], _055880_);
  xor g_114195_(out[54], out[726], _055881_);
  xor g_114196_(out[58], out[730], _055882_);
  xor g_114197_(out[53], out[725], _055883_);
  xor g_114198_(out[63], out[735], _055884_);
  xor g_114199_(out[61], out[733], _055885_);
  xor g_114200_(out[56], out[728], _055886_);
  or g_114201_(_055873_, _055875_, _055887_);
  or g_114202_(_055885_, _055886_, _055888_);
  or g_114203_(_055876_, _055882_, _055889_);
  or g_114204_(_055888_, _055889_, _055891_);
  or g_114205_(_055874_, _055877_, _055892_);
  or g_114206_(_055878_, _055883_, _055893_);
  or g_114207_(_055892_, _055893_, _055894_);
  or g_114208_(_055891_, _055894_, _055895_);
  xor g_114209_(out[60], out[732], _055896_);
  or g_114210_(_055880_, _055896_, _055897_);
  xor g_114211_(out[55], out[727], _055898_);
  or g_114212_(_055881_, _055898_, _055899_);
  or g_114213_(_055897_, _055899_, _055900_);
  or g_114214_(_055871_, _055872_, _055902_);
  or g_114215_(_055884_, _055902_, _055903_);
  or g_114216_(_055900_, _055903_, _055904_);
  or g_114217_(_055895_, _055904_, _055905_);
  or g_114218_(_055887_, _055905_, _055906_);
  xor g_114219_(out[39], out[727], _055907_);
  and g_114220_(_098096_, out[731], _055908_);
  xor g_114221_(out[46], out[734], _055909_);
  xor g_114222_(out[40], out[728], _055910_);
  xor g_114223_(out[33], out[721], _055911_);
  xor g_114224_(out[45], out[733], _055913_);
  xor g_114225_(out[41], out[729], _055914_);
  xor g_114226_(out[36], out[724], _055915_);
  xor g_114227_(out[34], out[722], _055916_);
  and g_114228_(out[43], _049664_, _055917_);
  xor g_114229_(out[35], out[723], _055918_);
  xor g_114230_(out[38], out[726], _055919_);
  xor g_114231_(out[47], out[735], _055920_);
  xor g_114232_(out[42], out[730], _055921_);
  xor g_114233_(out[37], out[725], _055922_);
  xor g_114234_(out[32], out[720], _055924_);
  or g_114235_(_055909_, _055915_, _055925_);
  or g_114236_(_055910_, _055913_, _055926_);
  or g_114237_(_055916_, _055921_, _055927_);
  or g_114238_(_055926_, _055927_, _055928_);
  or g_114239_(_055914_, _055918_, _055929_);
  or g_114240_(_055922_, _055924_, _055930_);
  or g_114241_(_055929_, _055930_, _055931_);
  or g_114242_(_055928_, _055931_, _055932_);
  xor g_114243_(out[44], out[732], _055933_);
  or g_114244_(_055908_, _055933_, _055935_);
  or g_114245_(_055907_, _055919_, _055936_);
  or g_114246_(_055935_, _055936_, _055937_);
  or g_114247_(_055911_, _055917_, _055938_);
  or g_114248_(_055920_, _055938_, _055939_);
  or g_114249_(_055937_, _055939_, _055940_);
  or g_114250_(_055932_, _055940_, _055941_);
  or g_114251_(_055925_, _055941_, _055942_);
  xor g_114252_(out[17], out[721], _055943_);
  and g_114253_(out[27], _049664_, _055944_);
  xor g_114254_(out[30], out[734], _055946_);
  xor g_114255_(out[19], out[723], _055947_);
  xor g_114256_(out[20], out[724], _055948_);
  xor g_114257_(out[18], out[722], _055949_);
  xor g_114258_(out[25], out[729], _055950_);
  xor g_114259_(out[16], out[720], _055951_);
  and g_114260_(_098063_, out[731], _055952_);
  xor g_114261_(out[22], out[726], _055953_);
  xor g_114262_(out[26], out[730], _055954_);
  xor g_114263_(out[21], out[725], _055955_);
  xor g_114264_(out[31], out[735], _055957_);
  xor g_114265_(out[29], out[733], _055958_);
  xor g_114266_(out[24], out[728], _055959_);
  or g_114267_(_055946_, _055948_, _055960_);
  or g_114268_(_055958_, _055959_, _055961_);
  or g_114269_(_055949_, _055954_, _055962_);
  or g_114270_(_055961_, _055962_, _055963_);
  or g_114271_(_055947_, _055950_, _055964_);
  or g_114272_(_055951_, _055955_, _055965_);
  or g_114273_(_055964_, _055965_, _055966_);
  or g_114274_(_055963_, _055966_, _055968_);
  xor g_114275_(out[28], out[732], _055969_);
  or g_114276_(_055952_, _055969_, _055970_);
  xor g_114277_(out[23], out[727], _055971_);
  or g_114278_(_055953_, _055971_, _055972_);
  or g_114279_(_055970_, _055972_, _055973_);
  or g_114280_(_055943_, _055944_, _055974_);
  or g_114281_(_055957_, _055974_, _055975_);
  or g_114282_(_055973_, _055975_, _055976_);
  or g_114283_(_055968_, _055976_, _055977_);
  or g_114284_(_055960_, _055977_, _055979_);
  xor g_114285_(out[1], out[721], _055980_);
  and g_114286_(_098041_, out[731], _055981_);
  and g_114287_(out[11], _049664_, _055982_);
  xor g_114288_(out[13], out[733], _055983_);
  xor g_114289_(out[10], out[730], _055984_);
  xor g_114290_(out[4], out[724], _055985_);
  xor g_114291_(out[14], out[734], _055986_);
  or g_114292_(_055985_, _055986_, _055987_);
  xor g_114293_(out[8], out[728], _055988_);
  xor g_114294_(out[0], out[720], _055990_);
  xor g_114295_(out[2], out[722], _055991_);
  xor g_114296_(out[9], out[729], _055992_);
  xor g_114297_(out[5], out[725], _055993_);
  xor g_114298_(out[3], out[723], _055994_);
  xor g_114299_(out[15], out[735], _055995_);
  xor g_114300_(out[6], out[726], _055996_);
  or g_114301_(_055983_, _055988_, _055997_);
  or g_114302_(_055984_, _055991_, _055998_);
  or g_114303_(_055997_, _055998_, _055999_);
  or g_114304_(_055992_, _055994_, _056001_);
  or g_114305_(_055990_, _055993_, _056002_);
  or g_114306_(_056001_, _056002_, _056003_);
  or g_114307_(_055999_, _056003_, _056004_);
  xor g_114308_(out[12], out[732], _056005_);
  or g_114309_(_055981_, _056005_, _056006_);
  xor g_114310_(out[7], out[727], _056007_);
  or g_114311_(_055996_, _056007_, _056008_);
  or g_114312_(_056006_, _056008_, _056009_);
  or g_114313_(_055980_, _055982_, _056010_);
  or g_114314_(_055995_, _056010_, _056012_);
  or g_114315_(_056009_, _056012_, _056013_);
  or g_114316_(_056004_, _056013_, _056014_);
  or g_114317_(_055987_, _056014_, _056015_);
  xor g_114318_(out[471], out[711], _056016_);
  and g_114319_(_049499_, out[715], _056017_);
  xor g_114320_(out[478], out[718], _056018_);
  xor g_114321_(out[472], out[712], _056019_);
  xor g_114322_(out[465], out[705], _056020_);
  xor g_114323_(out[477], out[717], _056021_);
  xor g_114324_(out[473], out[713], _056023_);
  xor g_114325_(out[468], out[708], _056024_);
  xor g_114326_(out[466], out[706], _056025_);
  and g_114327_(out[475], _049653_, _056026_);
  xor g_114328_(out[467], out[707], _056027_);
  xor g_114329_(out[470], out[710], _056028_);
  xor g_114330_(out[479], out[719], _056029_);
  xor g_114331_(out[474], out[714], _056030_);
  xor g_114332_(out[469], out[709], _056031_);
  xor g_114333_(out[464], out[704], _056032_);
  or g_114334_(_056018_, _056024_, _056034_);
  or g_114335_(_056019_, _056021_, _056035_);
  or g_114336_(_056025_, _056030_, _056036_);
  or g_114337_(_056035_, _056036_, _056037_);
  or g_114338_(_056023_, _056027_, _056038_);
  or g_114339_(_056031_, _056032_, _056039_);
  or g_114340_(_056038_, _056039_, _056040_);
  or g_114341_(_056037_, _056040_, _056041_);
  xor g_114342_(out[476], out[716], _056042_);
  or g_114343_(_056017_, _056042_, _056043_);
  or g_114344_(_056016_, _056028_, _056045_);
  or g_114345_(_056043_, _056045_, _056046_);
  or g_114346_(_056020_, _056026_, _056047_);
  or g_114347_(_056029_, _056047_, _056048_);
  or g_114348_(_056046_, _056048_, _056049_);
  or g_114349_(_056041_, _056049_, _056050_);
  or g_114350_(_056034_, _056050_, _056051_);
  xor g_114351_(out[456], out[712], _056052_);
  xor g_114352_(out[453], out[709], _056053_);
  xor g_114353_(out[451], out[707], _056054_);
  xor g_114354_(out[462], out[718], _056056_);
  xor g_114355_(out[461], out[717], _056057_);
  xor g_114356_(out[450], out[706], _056058_);
  xor g_114357_(out[457], out[713], _056059_);
  xor g_114358_(out[454], out[710], _056060_);
  xor g_114359_(out[463], out[719], _056061_);
  xor g_114360_(out[458], out[714], _056062_);
  xor g_114361_(out[452], out[708], _056063_);
  xor g_114362_(out[448], out[704], _056064_);
  and g_114363_(_049477_, out[715], _056065_);
  and g_114364_(out[459], _049653_, _056067_);
  or g_114365_(_056052_, _056057_, _056068_);
  xor g_114366_(out[449], out[705], _056069_);
  or g_114367_(_056058_, _056062_, _056070_);
  or g_114368_(_056068_, _056070_, _056071_);
  or g_114369_(_056054_, _056059_, _056072_);
  or g_114370_(_056053_, _056072_, _056073_);
  or g_114371_(_056071_, _056073_, _056074_);
  or g_114372_(_056056_, _056063_, _056075_);
  or g_114373_(_056074_, _056075_, _056076_);
  xor g_114374_(out[460], out[716], _056078_);
  or g_114375_(_056065_, _056078_, _056079_);
  xor g_114376_(out[455], out[711], _056080_);
  or g_114377_(_056060_, _056080_, _056081_);
  or g_114378_(_056079_, _056081_, _056082_);
  or g_114379_(_056067_, _056069_, _056083_);
  or g_114380_(_056061_, _056083_, _056084_);
  or g_114381_(_056082_, _056084_, _056085_);
  or g_114382_(_056064_, _056085_, _056086_);
  or g_114383_(_056076_, _056086_, _056087_);
  xor g_114384_(out[439], out[711], _056089_);
  and g_114385_(_049466_, out[715], _056090_);
  xor g_114386_(out[446], out[718], _056091_);
  xor g_114387_(out[440], out[712], _056092_);
  xor g_114388_(out[433], out[705], _056093_);
  xor g_114389_(out[445], out[717], _056094_);
  xor g_114390_(out[441], out[713], _056095_);
  xor g_114391_(out[436], out[708], _056096_);
  xor g_114392_(out[434], out[706], _056097_);
  and g_114393_(out[443], _049653_, _056098_);
  xor g_114394_(out[435], out[707], _056100_);
  xor g_114395_(out[438], out[710], _056101_);
  xor g_114396_(out[447], out[719], _056102_);
  xor g_114397_(out[442], out[714], _056103_);
  xor g_114398_(out[437], out[709], _056104_);
  xor g_114399_(out[432], out[704], _056105_);
  or g_114400_(_056091_, _056096_, _056106_);
  or g_114401_(_056092_, _056094_, _056107_);
  or g_114402_(_056097_, _056103_, _056108_);
  or g_114403_(_056107_, _056108_, _056109_);
  or g_114404_(_056095_, _056100_, _056111_);
  or g_114405_(_056104_, _056105_, _056112_);
  or g_114406_(_056111_, _056112_, _056113_);
  or g_114407_(_056109_, _056113_, _056114_);
  xor g_114408_(out[444], out[716], _056115_);
  or g_114409_(_056090_, _056115_, _056116_);
  or g_114410_(_056089_, _056101_, _056117_);
  or g_114411_(_056116_, _056117_, _056118_);
  or g_114412_(_056093_, _056098_, _056119_);
  or g_114413_(_056102_, _056119_, _056120_);
  or g_114414_(_056118_, _056120_, _056122_);
  or g_114415_(_056114_, _056122_, _056123_);
  or g_114416_(_056106_, _056123_, _056124_);
  xor g_114417_(out[417], out[705], _056125_);
  and g_114418_(out[427], _049653_, _056126_);
  xor g_114419_(out[430], out[718], _056127_);
  xor g_114420_(out[419], out[707], _056128_);
  xor g_114421_(out[420], out[708], _056129_);
  xor g_114422_(out[418], out[706], _056130_);
  xor g_114423_(out[425], out[713], _056131_);
  xor g_114424_(out[416], out[704], _056133_);
  and g_114425_(_049455_, out[715], _056134_);
  xor g_114426_(out[422], out[710], _056135_);
  xor g_114427_(out[426], out[714], _056136_);
  xor g_114428_(out[421], out[709], _056137_);
  xor g_114429_(out[431], out[719], _056138_);
  xor g_114430_(out[429], out[717], _056139_);
  xor g_114431_(out[424], out[712], _056140_);
  or g_114432_(_056127_, _056129_, _056141_);
  or g_114433_(_056139_, _056140_, _056142_);
  or g_114434_(_056130_, _056136_, _056144_);
  or g_114435_(_056142_, _056144_, _056145_);
  or g_114436_(_056128_, _056131_, _056146_);
  or g_114437_(_056133_, _056137_, _056147_);
  or g_114438_(_056146_, _056147_, _056148_);
  or g_114439_(_056145_, _056148_, _056149_);
  xor g_114440_(out[428], out[716], _056150_);
  or g_114441_(_056134_, _056150_, _056151_);
  xor g_114442_(out[423], out[711], _056152_);
  or g_114443_(_056135_, _056152_, _056153_);
  or g_114444_(_056151_, _056153_, _056155_);
  or g_114445_(_056125_, _056126_, _056156_);
  or g_114446_(_056138_, _056156_, _056157_);
  or g_114447_(_056155_, _056157_, _056158_);
  or g_114448_(_056149_, _056158_, _056159_);
  or g_114449_(_056141_, _056159_, _056160_);
  xor g_114450_(out[407], out[711], _056161_);
  and g_114451_(_049444_, out[715], _056162_);
  xor g_114452_(out[414], out[718], _056163_);
  xor g_114453_(out[408], out[712], _056164_);
  xor g_114454_(out[401], out[705], _056166_);
  xor g_114455_(out[413], out[717], _056167_);
  xor g_114456_(out[409], out[713], _056168_);
  xor g_114457_(out[404], out[708], _056169_);
  xor g_114458_(out[402], out[706], _056170_);
  and g_114459_(out[411], _049653_, _056171_);
  xor g_114460_(out[403], out[707], _056172_);
  xor g_114461_(out[406], out[710], _056173_);
  xor g_114462_(out[415], out[719], _056174_);
  xor g_114463_(out[410], out[714], _056175_);
  xor g_114464_(out[405], out[709], _056177_);
  xor g_114465_(out[400], out[704], _056178_);
  or g_114466_(_056163_, _056169_, _056179_);
  or g_114467_(_056164_, _056167_, _056180_);
  or g_114468_(_056170_, _056175_, _056181_);
  or g_114469_(_056180_, _056181_, _056182_);
  or g_114470_(_056168_, _056172_, _056183_);
  or g_114471_(_056177_, _056178_, _056184_);
  or g_114472_(_056183_, _056184_, _056185_);
  or g_114473_(_056182_, _056185_, _056186_);
  xor g_114474_(out[412], out[716], _056188_);
  or g_114475_(_056162_, _056188_, _056189_);
  or g_114476_(_056161_, _056173_, _056190_);
  or g_114477_(_056189_, _056190_, _056191_);
  or g_114478_(_056166_, _056171_, _056192_);
  or g_114479_(_056174_, _056192_, _056193_);
  or g_114480_(_056191_, _056193_, _056194_);
  or g_114481_(_056186_, _056194_, _056195_);
  or g_114482_(_056179_, _056195_, _056196_);
  xor g_114483_(out[385], out[705], _056197_);
  and g_114484_(out[395], _049653_, _056199_);
  xor g_114485_(out[393], out[713], _056200_);
  xor g_114486_(out[384], out[704], _056201_);
  xor g_114487_(out[398], out[718], _056202_);
  xor g_114488_(out[388], out[708], _056203_);
  or g_114489_(_056202_, _056203_, _056204_);
  xor g_114490_(out[397], out[717], _056205_);
  xor g_114491_(out[387], out[707], _056206_);
  and g_114492_(_049433_, out[715], _056207_);
  xor g_114493_(out[390], out[710], _056208_);
  xor g_114494_(out[394], out[714], _056210_);
  xor g_114495_(out[389], out[709], _056211_);
  xor g_114496_(out[399], out[719], _056212_);
  xor g_114497_(out[392], out[712], _056213_);
  or g_114498_(_056205_, _056213_, _056214_);
  xor g_114499_(out[386], out[706], _056215_);
  or g_114500_(_056210_, _056215_, _056216_);
  or g_114501_(_056214_, _056216_, _056217_);
  or g_114502_(_056200_, _056206_, _056218_);
  or g_114503_(_056211_, _056218_, _056219_);
  or g_114504_(_056217_, _056219_, _056221_);
  or g_114505_(_056204_, _056221_, _056222_);
  xor g_114506_(out[396], out[716], _056223_);
  or g_114507_(_056207_, _056223_, _056224_);
  xor g_114508_(out[391], out[711], _056225_);
  or g_114509_(_056208_, _056225_, _056226_);
  or g_114510_(_056224_, _056226_, _056227_);
  or g_114511_(_056197_, _056199_, _056228_);
  or g_114512_(_056212_, _056228_, _056229_);
  or g_114513_(_056227_, _056229_, _056230_);
  or g_114514_(_056201_, _056230_, _056232_);
  or g_114515_(_056222_, _056232_, _056233_);
  xor g_114516_(out[375], out[711], _056234_);
  and g_114517_(_049422_, out[715], _056235_);
  xor g_114518_(out[382], out[718], _056236_);
  xor g_114519_(out[376], out[712], _056237_);
  xor g_114520_(out[369], out[705], _056238_);
  xor g_114521_(out[381], out[717], _056239_);
  xor g_114522_(out[377], out[713], _056240_);
  xor g_114523_(out[372], out[708], _056241_);
  xor g_114524_(out[370], out[706], _056243_);
  and g_114525_(out[379], _049653_, _056244_);
  xor g_114526_(out[371], out[707], _056245_);
  xor g_114527_(out[374], out[710], _056246_);
  xor g_114528_(out[383], out[719], _056247_);
  xor g_114529_(out[378], out[714], _056248_);
  xor g_114530_(out[373], out[709], _056249_);
  xor g_114531_(out[368], out[704], _056250_);
  or g_114532_(_056236_, _056241_, _056251_);
  or g_114533_(_056237_, _056239_, _056252_);
  or g_114534_(_056243_, _056248_, _056254_);
  or g_114535_(_056252_, _056254_, _056255_);
  or g_114536_(_056240_, _056245_, _056256_);
  or g_114537_(_056249_, _056250_, _056257_);
  or g_114538_(_056256_, _056257_, _056258_);
  or g_114539_(_056255_, _056258_, _056259_);
  xor g_114540_(out[380], out[716], _056260_);
  or g_114541_(_056235_, _056260_, _056261_);
  or g_114542_(_056234_, _056246_, _056262_);
  or g_114543_(_056261_, _056262_, _056263_);
  or g_114544_(_056238_, _056244_, _056265_);
  or g_114545_(_056247_, _056265_, _056266_);
  or g_114546_(_056263_, _056266_, _056267_);
  or g_114547_(_056259_, _056267_, _056268_);
  or g_114548_(_056251_, _056268_, _056269_);
  xor g_114549_(out[353], out[705], _056270_);
  and g_114550_(out[363], _049653_, _056271_);
  xor g_114551_(out[361], out[713], _056272_);
  xor g_114552_(out[352], out[704], _056273_);
  xor g_114553_(out[366], out[718], _056274_);
  xor g_114554_(out[356], out[708], _056276_);
  or g_114555_(_056274_, _056276_, _056277_);
  xor g_114556_(out[365], out[717], _056278_);
  xor g_114557_(out[355], out[707], _056279_);
  and g_114558_(_049411_, out[715], _056280_);
  xor g_114559_(out[358], out[710], _056281_);
  xor g_114560_(out[362], out[714], _056282_);
  xor g_114561_(out[357], out[709], _056283_);
  xor g_114562_(out[367], out[719], _056284_);
  xor g_114563_(out[360], out[712], _056285_);
  or g_114564_(_056278_, _056285_, _056287_);
  xor g_114565_(out[354], out[706], _056288_);
  or g_114566_(_056282_, _056288_, _056289_);
  or g_114567_(_056287_, _056289_, _056290_);
  or g_114568_(_056272_, _056279_, _056291_);
  or g_114569_(_056283_, _056291_, _056292_);
  or g_114570_(_056290_, _056292_, _056293_);
  or g_114571_(_056277_, _056293_, _056294_);
  xor g_114572_(out[364], out[716], _056295_);
  or g_114573_(_056280_, _056295_, _056296_);
  xor g_114574_(out[359], out[711], _056298_);
  or g_114575_(_056281_, _056298_, _056299_);
  or g_114576_(_056296_, _056299_, _056300_);
  or g_114577_(_056270_, _056271_, _056301_);
  or g_114578_(_056284_, _056301_, _056302_);
  or g_114579_(_056300_, _056302_, _056303_);
  or g_114580_(_056273_, _056303_, _056304_);
  or g_114581_(_056294_, _056304_, _056305_);
  xor g_114582_(out[343], out[711], _056306_);
  and g_114583_(_049400_, out[715], _056307_);
  xor g_114584_(out[350], out[718], _056309_);
  xor g_114585_(out[344], out[712], _056310_);
  xor g_114586_(out[337], out[705], _056311_);
  xor g_114587_(out[349], out[717], _056312_);
  xor g_114588_(out[345], out[713], _056313_);
  xor g_114589_(out[340], out[708], _056314_);
  xor g_114590_(out[338], out[706], _056315_);
  and g_114591_(out[347], _049653_, _056316_);
  xor g_114592_(out[339], out[707], _056317_);
  xor g_114593_(out[342], out[710], _056318_);
  xor g_114594_(out[351], out[719], _056320_);
  xor g_114595_(out[346], out[714], _056321_);
  xor g_114596_(out[341], out[709], _056322_);
  xor g_114597_(out[336], out[704], _056323_);
  or g_114598_(_056309_, _056314_, _056324_);
  or g_114599_(_056310_, _056312_, _056325_);
  or g_114600_(_056315_, _056321_, _056326_);
  or g_114601_(_056325_, _056326_, _056327_);
  or g_114602_(_056313_, _056317_, _056328_);
  or g_114603_(_056322_, _056323_, _056329_);
  or g_114604_(_056328_, _056329_, _056331_);
  or g_114605_(_056327_, _056331_, _056332_);
  xor g_114606_(out[348], out[716], _056333_);
  or g_114607_(_056307_, _056333_, _056334_);
  or g_114608_(_056306_, _056318_, _056335_);
  or g_114609_(_056334_, _056335_, _056336_);
  or g_114610_(_056311_, _056316_, _056337_);
  or g_114611_(_056320_, _056337_, _056338_);
  or g_114612_(_056336_, _056338_, _056339_);
  or g_114613_(_056332_, _056339_, _056340_);
  or g_114614_(_056324_, _056340_, _056342_);
  xor g_114615_(out[332], out[716], _056343_);
  and g_114616_(_098294_, out[715], _056344_);
  xor g_114617_(out[333], out[717], _056345_);
  xor g_114618_(out[326], out[710], _056346_);
  xor g_114619_(out[328], out[712], _056347_);
  xor g_114620_(out[329], out[713], _056348_);
  xor g_114621_(out[334], out[718], _056349_);
  xor g_114622_(out[324], out[708], _056350_);
  or g_114623_(_056349_, _056350_, _056351_);
  xor g_114624_(out[325], out[709], _056353_);
  xor g_114625_(out[321], out[705], _056354_);
  and g_114626_(out[331], _049653_, _056355_);
  xor g_114627_(out[335], out[719], _056356_);
  xor g_114628_(out[330], out[714], _056357_);
  xor g_114629_(out[320], out[704], _056358_);
  xor g_114630_(out[322], out[706], _056359_);
  xor g_114631_(out[323], out[707], _056360_);
  or g_114632_(_056345_, _056347_, _056361_);
  or g_114633_(_056357_, _056359_, _056362_);
  or g_114634_(_056361_, _056362_, _056364_);
  or g_114635_(_056348_, _056360_, _056365_);
  or g_114636_(_056353_, _056358_, _056366_);
  or g_114637_(_056365_, _056366_, _056367_);
  or g_114638_(_056364_, _056367_, _056368_);
  or g_114639_(_056343_, _056344_, _056369_);
  xor g_114640_(out[327], out[711], _056370_);
  or g_114641_(_056346_, _056370_, _056371_);
  or g_114642_(_056369_, _056371_, _056372_);
  or g_114643_(_056354_, _056355_, _056373_);
  or g_114644_(_056356_, _056373_, _056375_);
  or g_114645_(_056372_, _056375_, _056376_);
  or g_114646_(_056368_, _056376_, _056377_);
  or g_114647_(_056351_, _056377_, _056378_);
  not g_114648_(_056378_, _056379_);
  xor g_114649_(out[311], out[711], _056380_);
  and g_114650_(_098283_, out[715], _056381_);
  xor g_114651_(out[318], out[718], _056382_);
  xor g_114652_(out[312], out[712], _056383_);
  xor g_114653_(out[305], out[705], _056384_);
  xor g_114654_(out[317], out[717], _056386_);
  xor g_114655_(out[313], out[713], _056387_);
  xor g_114656_(out[308], out[708], _056388_);
  xor g_114657_(out[306], out[706], _056389_);
  and g_114658_(out[315], _049653_, _056390_);
  xor g_114659_(out[307], out[707], _056391_);
  xor g_114660_(out[310], out[710], _056392_);
  xor g_114661_(out[319], out[719], _056393_);
  xor g_114662_(out[314], out[714], _056394_);
  xor g_114663_(out[309], out[709], _056395_);
  xor g_114664_(out[304], out[704], _056397_);
  or g_114665_(_056382_, _056388_, _056398_);
  or g_114666_(_056383_, _056386_, _056399_);
  or g_114667_(_056389_, _056394_, _056400_);
  or g_114668_(_056399_, _056400_, _056401_);
  or g_114669_(_056387_, _056391_, _056402_);
  or g_114670_(_056395_, _056397_, _056403_);
  or g_114671_(_056402_, _056403_, _056404_);
  or g_114672_(_056401_, _056404_, _056405_);
  xor g_114673_(out[316], out[716], _056406_);
  or g_114674_(_056381_, _056406_, _056408_);
  or g_114675_(_056380_, _056392_, _056409_);
  or g_114676_(_056408_, _056409_, _056410_);
  or g_114677_(_056384_, _056390_, _056411_);
  or g_114678_(_056393_, _056411_, _056412_);
  or g_114679_(_056410_, _056412_, _056413_);
  or g_114680_(_056405_, _056413_, _056414_);
  or g_114681_(_056398_, _056414_, _056415_);
  not g_114682_(_056415_, _056416_);
  xor g_114683_(out[291], out[707], _056417_);
  xor g_114684_(out[292], out[708], _056419_);
  xor g_114685_(out[302], out[718], _056420_);
  xor g_114686_(out[290], out[706], _056421_);
  xor g_114687_(out[293], out[709], _056422_);
  xor g_114688_(out[297], out[713], _056423_);
  xor g_114689_(out[296], out[712], _056424_);
  xor g_114690_(out[303], out[719], _056425_);
  xor g_114691_(out[298], out[714], _056426_);
  xor g_114692_(out[294], out[710], _056427_);
  xor g_114693_(out[288], out[704], _056428_);
  and g_114694_(_098272_, out[715], _056430_);
  and g_114695_(out[299], _049653_, _056431_);
  xor g_114696_(out[301], out[717], _056432_);
  or g_114697_(_056424_, _056432_, _056433_);
  xor g_114698_(out[289], out[705], _056434_);
  or g_114699_(_056421_, _056426_, _056435_);
  or g_114700_(_056433_, _056435_, _056436_);
  or g_114701_(_056417_, _056423_, _056437_);
  or g_114702_(_056422_, _056437_, _056438_);
  or g_114703_(_056436_, _056438_, _056439_);
  or g_114704_(_056419_, _056420_, _056441_);
  or g_114705_(_056439_, _056441_, _056442_);
  xor g_114706_(out[300], out[716], _056443_);
  or g_114707_(_056430_, _056443_, _056444_);
  xor g_114708_(out[295], out[711], _056445_);
  or g_114709_(_056427_, _056445_, _056446_);
  or g_114710_(_056444_, _056446_, _056447_);
  or g_114711_(_056431_, _056434_, _056448_);
  or g_114712_(_056425_, _056448_, _056449_);
  or g_114713_(_056447_, _056449_, _056450_);
  or g_114714_(_056428_, _056450_, _056452_);
  or g_114715_(_056442_, _056452_, _056453_);
  xor g_114716_(out[279], out[711], _056454_);
  and g_114717_(_098261_, out[715], _056455_);
  xor g_114718_(out[286], out[718], _056456_);
  xor g_114719_(out[280], out[712], _056457_);
  xor g_114720_(out[273], out[705], _056458_);
  xor g_114721_(out[285], out[717], _056459_);
  xor g_114722_(out[281], out[713], _056460_);
  xor g_114723_(out[276], out[708], _056461_);
  xor g_114724_(out[274], out[706], _056463_);
  and g_114725_(out[283], _049653_, _056464_);
  xor g_114726_(out[275], out[707], _056465_);
  xor g_114727_(out[278], out[710], _056466_);
  xor g_114728_(out[287], out[719], _056467_);
  xor g_114729_(out[282], out[714], _056468_);
  xor g_114730_(out[277], out[709], _056469_);
  xor g_114731_(out[272], out[704], _056470_);
  or g_114732_(_056456_, _056461_, _056471_);
  or g_114733_(_056457_, _056459_, _056472_);
  or g_114734_(_056463_, _056468_, _056474_);
  or g_114735_(_056472_, _056474_, _056475_);
  or g_114736_(_056460_, _056465_, _056476_);
  or g_114737_(_056469_, _056470_, _056477_);
  or g_114738_(_056476_, _056477_, _056478_);
  or g_114739_(_056475_, _056478_, _056479_);
  xor g_114740_(out[284], out[716], _056480_);
  or g_114741_(_056455_, _056480_, _056481_);
  or g_114742_(_056454_, _056466_, _056482_);
  or g_114743_(_056481_, _056482_, _056483_);
  or g_114744_(_056458_, _056464_, _056485_);
  or g_114745_(_056467_, _056485_, _056486_);
  or g_114746_(_056483_, _056486_, _056487_);
  or g_114747_(_056479_, _056487_, _056488_);
  or g_114748_(_056471_, _056488_, _056489_);
  xor g_114749_(out[257], out[705], _056490_);
  and g_114750_(out[267], _049653_, _056491_);
  xor g_114751_(out[265], out[713], _056492_);
  xor g_114752_(out[256], out[704], _056493_);
  xor g_114753_(out[270], out[718], _056494_);
  xor g_114754_(out[260], out[708], _056496_);
  or g_114755_(_056494_, _056496_, _056497_);
  xor g_114756_(out[269], out[717], _056498_);
  xor g_114757_(out[259], out[707], _056499_);
  and g_114758_(_098250_, out[715], _056500_);
  xor g_114759_(out[262], out[710], _056501_);
  xor g_114760_(out[266], out[714], _056502_);
  xor g_114761_(out[261], out[709], _056503_);
  xor g_114762_(out[271], out[719], _056504_);
  xor g_114763_(out[264], out[712], _056505_);
  or g_114764_(_056498_, _056505_, _056507_);
  xor g_114765_(out[258], out[706], _056508_);
  or g_114766_(_056502_, _056508_, _056509_);
  or g_114767_(_056507_, _056509_, _056510_);
  or g_114768_(_056492_, _056499_, _056511_);
  or g_114769_(_056503_, _056511_, _056512_);
  or g_114770_(_056510_, _056512_, _056513_);
  or g_114771_(_056497_, _056513_, _056514_);
  xor g_114772_(out[268], out[716], _056515_);
  or g_114773_(_056500_, _056515_, _056516_);
  xor g_114774_(out[263], out[711], _056518_);
  or g_114775_(_056501_, _056518_, _056519_);
  or g_114776_(_056516_, _056519_, _056520_);
  or g_114777_(_056490_, _056491_, _056521_);
  or g_114778_(_056504_, _056521_, _056522_);
  or g_114779_(_056520_, _056522_, _056523_);
  or g_114780_(_056493_, _056523_, _056524_);
  or g_114781_(_056514_, _056524_, _056525_);
  xor g_114782_(out[247], out[711], _056526_);
  and g_114783_(_098239_, out[715], _056527_);
  xor g_114784_(out[254], out[718], _056529_);
  xor g_114785_(out[248], out[712], _056530_);
  xor g_114786_(out[241], out[705], _056531_);
  xor g_114787_(out[253], out[717], _056532_);
  xor g_114788_(out[249], out[713], _056533_);
  xor g_114789_(out[244], out[708], _056534_);
  xor g_114790_(out[242], out[706], _056535_);
  and g_114791_(out[251], _049653_, _056536_);
  xor g_114792_(out[243], out[707], _056537_);
  xor g_114793_(out[246], out[710], _056538_);
  xor g_114794_(out[255], out[719], _056540_);
  xor g_114795_(out[250], out[714], _056541_);
  xor g_114796_(out[245], out[709], _056542_);
  xor g_114797_(out[240], out[704], _056543_);
  or g_114798_(_056529_, _056534_, _056544_);
  or g_114799_(_056530_, _056532_, _056545_);
  or g_114800_(_056535_, _056541_, _056546_);
  or g_114801_(_056545_, _056546_, _056547_);
  or g_114802_(_056533_, _056537_, _056548_);
  or g_114803_(_056542_, _056543_, _056549_);
  or g_114804_(_056548_, _056549_, _056551_);
  or g_114805_(_056547_, _056551_, _056552_);
  xor g_114806_(out[252], out[716], _056553_);
  or g_114807_(_056527_, _056553_, _056554_);
  or g_114808_(_056526_, _056538_, _056555_);
  or g_114809_(_056554_, _056555_, _056556_);
  or g_114810_(_056531_, _056536_, _056557_);
  or g_114811_(_056540_, _056557_, _056558_);
  or g_114812_(_056556_, _056558_, _056559_);
  or g_114813_(_056552_, _056559_, _056560_);
  or g_114814_(_056544_, _056560_, _056562_);
  xor g_114815_(out[226], out[706], _056563_);
  xor g_114816_(out[224], out[704], _056564_);
  xor g_114817_(out[233], out[713], _056565_);
  xor g_114818_(out[232], out[712], _056566_);
  xor g_114819_(out[229], out[709], _056567_);
  xor g_114820_(out[238], out[718], _056568_);
  xor g_114821_(out[237], out[717], _056569_);
  xor g_114822_(out[239], out[719], _056570_);
  xor g_114823_(out[234], out[714], _056571_);
  xor g_114824_(out[230], out[710], _056573_);
  xor g_114825_(out[227], out[707], _056574_);
  and g_114826_(_098228_, out[715], _056575_);
  and g_114827_(out[235], _049653_, _056576_);
  xor g_114828_(out[228], out[708], _056577_);
  xor g_114829_(out[225], out[705], _056578_);
  or g_114830_(_056568_, _056577_, _056579_);
  or g_114831_(_056566_, _056569_, _056580_);
  or g_114832_(_056563_, _056571_, _056581_);
  or g_114833_(_056580_, _056581_, _056582_);
  or g_114834_(_056565_, _056574_, _056584_);
  or g_114835_(_056564_, _056567_, _056585_);
  or g_114836_(_056584_, _056585_, _056586_);
  or g_114837_(_056582_, _056586_, _056587_);
  xor g_114838_(out[236], out[716], _056588_);
  or g_114839_(_056575_, _056588_, _056589_);
  xor g_114840_(out[231], out[711], _056590_);
  or g_114841_(_056573_, _056590_, _056591_);
  or g_114842_(_056589_, _056591_, _056592_);
  or g_114843_(_056576_, _056578_, _056593_);
  or g_114844_(_056570_, _056593_, _056595_);
  or g_114845_(_056592_, _056595_, _056596_);
  or g_114846_(_056587_, _056596_, _056597_);
  or g_114847_(_056579_, _056597_, _056598_);
  not g_114848_(_056598_, _056599_);
  xor g_114849_(out[215], out[711], _056600_);
  and g_114850_(_098217_, out[715], _056601_);
  xor g_114851_(out[222], out[718], _056602_);
  xor g_114852_(out[216], out[712], _056603_);
  xor g_114853_(out[209], out[705], _056604_);
  xor g_114854_(out[221], out[717], _056606_);
  xor g_114855_(out[217], out[713], _056607_);
  xor g_114856_(out[212], out[708], _056608_);
  xor g_114857_(out[210], out[706], _056609_);
  and g_114858_(out[219], _049653_, _056610_);
  xor g_114859_(out[211], out[707], _056611_);
  xor g_114860_(out[214], out[710], _056612_);
  xor g_114861_(out[223], out[719], _056613_);
  xor g_114862_(out[218], out[714], _056614_);
  xor g_114863_(out[213], out[709], _056615_);
  xor g_114864_(out[208], out[704], _056617_);
  or g_114865_(_056602_, _056608_, _056618_);
  or g_114866_(_056603_, _056606_, _056619_);
  or g_114867_(_056609_, _056614_, _056620_);
  or g_114868_(_056619_, _056620_, _056621_);
  or g_114869_(_056607_, _056611_, _056622_);
  or g_114870_(_056615_, _056617_, _056623_);
  or g_114871_(_056622_, _056623_, _056624_);
  or g_114872_(_056621_, _056624_, _056625_);
  xor g_114873_(out[220], out[716], _056626_);
  or g_114874_(_056601_, _056626_, _056628_);
  or g_114875_(_056600_, _056612_, _056629_);
  or g_114876_(_056628_, _056629_, _056630_);
  or g_114877_(_056604_, _056610_, _056631_);
  or g_114878_(_056613_, _056631_, _056632_);
  or g_114879_(_056630_, _056632_, _056633_);
  or g_114880_(_056625_, _056633_, _056634_);
  or g_114881_(_056618_, _056634_, _056635_);
  xor g_114882_(out[204], out[716], _056636_);
  and g_114883_(_098206_, out[715], _056637_);
  xor g_114884_(out[200], out[712], _056639_);
  xor g_114885_(out[198], out[710], _056640_);
  xor g_114886_(out[205], out[717], _056641_);
  xor g_114887_(out[206], out[718], _056642_);
  xor g_114888_(out[194], out[706], _056643_);
  xor g_114889_(out[201], out[713], _056644_);
  xor g_114890_(out[197], out[709], _056645_);
  xor g_114891_(out[193], out[705], _056646_);
  and g_114892_(out[203], _049653_, _056647_);
  or g_114893_(_056639_, _056641_, _056648_);
  xor g_114894_(out[207], out[719], _056650_);
  xor g_114895_(out[202], out[714], _056651_);
  xor g_114896_(out[196], out[708], _056652_);
  xor g_114897_(out[195], out[707], _056653_);
  xor g_114898_(out[192], out[704], _056654_);
  or g_114899_(_056643_, _056651_, _056655_);
  or g_114900_(_056648_, _056655_, _056656_);
  or g_114901_(_056644_, _056653_, _056657_);
  or g_114902_(_056645_, _056657_, _056658_);
  or g_114903_(_056656_, _056658_, _056659_);
  or g_114904_(_056642_, _056652_, _056661_);
  or g_114905_(_056659_, _056661_, _056662_);
  or g_114906_(_056636_, _056637_, _056663_);
  xor g_114907_(out[199], out[711], _056664_);
  or g_114908_(_056640_, _056664_, _056665_);
  or g_114909_(_056663_, _056665_, _056666_);
  or g_114910_(_056646_, _056647_, _056667_);
  or g_114911_(_056650_, _056667_, _056668_);
  or g_114912_(_056666_, _056668_, _056669_);
  or g_114913_(_056654_, _056669_, _056670_);
  or g_114914_(_056662_, _056670_, _056672_);
  not g_114915_(_056672_, _056673_);
  xor g_114916_(out[183], out[711], _056674_);
  and g_114917_(_098195_, out[715], _056675_);
  xor g_114918_(out[190], out[718], _056676_);
  xor g_114919_(out[184], out[712], _056677_);
  xor g_114920_(out[177], out[705], _056678_);
  xor g_114921_(out[189], out[717], _056679_);
  xor g_114922_(out[185], out[713], _056680_);
  xor g_114923_(out[180], out[708], _056681_);
  xor g_114924_(out[178], out[706], _056683_);
  and g_114925_(out[187], _049653_, _056684_);
  xor g_114926_(out[179], out[707], _056685_);
  xor g_114927_(out[182], out[710], _056686_);
  xor g_114928_(out[191], out[719], _056687_);
  xor g_114929_(out[186], out[714], _056688_);
  xor g_114930_(out[181], out[709], _056689_);
  xor g_114931_(out[176], out[704], _056690_);
  or g_114932_(_056676_, _056681_, _056691_);
  or g_114933_(_056677_, _056679_, _056692_);
  or g_114934_(_056683_, _056688_, _056694_);
  or g_114935_(_056692_, _056694_, _056695_);
  or g_114936_(_056680_, _056685_, _056696_);
  or g_114937_(_056689_, _056690_, _056697_);
  or g_114938_(_056696_, _056697_, _056698_);
  or g_114939_(_056695_, _056698_, _056699_);
  xor g_114940_(out[188], out[716], _056700_);
  or g_114941_(_056675_, _056700_, _056701_);
  or g_114942_(_056674_, _056686_, _056702_);
  or g_114943_(_056701_, _056702_, _056703_);
  or g_114944_(_056678_, _056684_, _056705_);
  or g_114945_(_056687_, _056705_, _056706_);
  or g_114946_(_056703_, _056706_, _056707_);
  or g_114947_(_056699_, _056707_, _056708_);
  or g_114948_(_056691_, _056708_, _056709_);
  not g_114949_(_056709_, _056710_);
  xor g_114950_(out[172], out[716], _056711_);
  and g_114951_(_098184_, out[715], _056712_);
  xor g_114952_(out[168], out[712], _056713_);
  xor g_114953_(out[166], out[710], _056714_);
  xor g_114954_(out[173], out[717], _056716_);
  xor g_114955_(out[174], out[718], _056717_);
  xor g_114956_(out[162], out[706], _056718_);
  xor g_114957_(out[169], out[713], _056719_);
  xor g_114958_(out[165], out[709], _056720_);
  xor g_114959_(out[161], out[705], _056721_);
  and g_114960_(out[171], _049653_, _056722_);
  or g_114961_(_056713_, _056716_, _056723_);
  xor g_114962_(out[175], out[719], _056724_);
  xor g_114963_(out[170], out[714], _056725_);
  xor g_114964_(out[164], out[708], _056727_);
  xor g_114965_(out[163], out[707], _056728_);
  xor g_114966_(out[160], out[704], _056729_);
  or g_114967_(_056718_, _056725_, _056730_);
  or g_114968_(_056723_, _056730_, _056731_);
  or g_114969_(_056719_, _056728_, _056732_);
  or g_114970_(_056720_, _056732_, _056733_);
  or g_114971_(_056731_, _056733_, _056734_);
  or g_114972_(_056717_, _056727_, _056735_);
  or g_114973_(_056734_, _056735_, _056736_);
  or g_114974_(_056711_, _056712_, _056738_);
  xor g_114975_(out[167], out[711], _056739_);
  or g_114976_(_056714_, _056739_, _056740_);
  or g_114977_(_056738_, _056740_, _056741_);
  or g_114978_(_056721_, _056722_, _056742_);
  or g_114979_(_056724_, _056742_, _056743_);
  or g_114980_(_056741_, _056743_, _056744_);
  or g_114981_(_056729_, _056744_, _056745_);
  or g_114982_(_056736_, _056745_, _056746_);
  not g_114983_(_056746_, _056747_);
  xor g_114984_(out[151], out[711], _056749_);
  and g_114985_(_098173_, out[715], _056750_);
  xor g_114986_(out[158], out[718], _056751_);
  xor g_114987_(out[152], out[712], _056752_);
  xor g_114988_(out[145], out[705], _056753_);
  xor g_114989_(out[157], out[717], _056754_);
  xor g_114990_(out[153], out[713], _056755_);
  xor g_114991_(out[148], out[708], _056756_);
  xor g_114992_(out[146], out[706], _056757_);
  and g_114993_(out[155], _049653_, _056758_);
  xor g_114994_(out[147], out[707], _056760_);
  xor g_114995_(out[150], out[710], _056761_);
  xor g_114996_(out[159], out[719], _056762_);
  xor g_114997_(out[154], out[714], _056763_);
  xor g_114998_(out[149], out[709], _056764_);
  xor g_114999_(out[144], out[704], _056765_);
  or g_115000_(_056751_, _056756_, _056766_);
  or g_115001_(_056752_, _056754_, _056767_);
  or g_115002_(_056757_, _056763_, _056768_);
  or g_115003_(_056767_, _056768_, _056769_);
  or g_115004_(_056755_, _056760_, _056771_);
  or g_115005_(_056764_, _056765_, _056772_);
  or g_115006_(_056771_, _056772_, _056773_);
  or g_115007_(_056769_, _056773_, _056774_);
  xor g_115008_(out[156], out[716], _056775_);
  or g_115009_(_056750_, _056775_, _056776_);
  or g_115010_(_056749_, _056761_, _056777_);
  or g_115011_(_056776_, _056777_, _056778_);
  or g_115012_(_056753_, _056758_, _056779_);
  or g_115013_(_056762_, _056779_, _056780_);
  or g_115014_(_056778_, _056780_, _056782_);
  or g_115015_(_056774_, _056782_, _056783_);
  or g_115016_(_056766_, _056783_, _056784_);
  not g_115017_(_056784_, _056785_);
  xor g_115018_(out[129], out[705], _056786_);
  and g_115019_(out[139], _049653_, _056787_);
  xor g_115020_(out[142], out[718], _056788_);
  xor g_115021_(out[131], out[707], _056789_);
  xor g_115022_(out[132], out[708], _056790_);
  xor g_115023_(out[130], out[706], _056791_);
  xor g_115024_(out[137], out[713], _056793_);
  xor g_115025_(out[128], out[704], _056794_);
  and g_115026_(_098162_, out[715], _056795_);
  xor g_115027_(out[134], out[710], _056796_);
  xor g_115028_(out[138], out[714], _056797_);
  xor g_115029_(out[133], out[709], _056798_);
  xor g_115030_(out[143], out[719], _056799_);
  xor g_115031_(out[141], out[717], _056800_);
  xor g_115032_(out[136], out[712], _056801_);
  or g_115033_(_056788_, _056790_, _056802_);
  or g_115034_(_056800_, _056801_, _056804_);
  or g_115035_(_056791_, _056797_, _056805_);
  or g_115036_(_056804_, _056805_, _056806_);
  or g_115037_(_056789_, _056793_, _056807_);
  or g_115038_(_056794_, _056798_, _056808_);
  or g_115039_(_056807_, _056808_, _056809_);
  or g_115040_(_056806_, _056809_, _056810_);
  xor g_115041_(out[140], out[716], _056811_);
  or g_115042_(_056795_, _056811_, _056812_);
  xor g_115043_(out[135], out[711], _056813_);
  or g_115044_(_056796_, _056813_, _056815_);
  or g_115045_(_056812_, _056815_, _056816_);
  or g_115046_(_056786_, _056787_, _056817_);
  or g_115047_(_056799_, _056817_, _056818_);
  or g_115048_(_056816_, _056818_, _056819_);
  or g_115049_(_056810_, _056819_, _056820_);
  or g_115050_(_056802_, _056820_, _056821_);
  not g_115051_(_056821_, _056822_);
  xor g_115052_(out[119], out[711], _056823_);
  and g_115053_(_098151_, out[715], _056824_);
  xor g_115054_(out[126], out[718], _056826_);
  xor g_115055_(out[120], out[712], _056827_);
  xor g_115056_(out[113], out[705], _056828_);
  xor g_115057_(out[125], out[717], _056829_);
  xor g_115058_(out[121], out[713], _056830_);
  xor g_115059_(out[116], out[708], _056831_);
  xor g_115060_(out[114], out[706], _056832_);
  and g_115061_(out[123], _049653_, _056833_);
  xor g_115062_(out[115], out[707], _056834_);
  xor g_115063_(out[118], out[710], _056835_);
  xor g_115064_(out[127], out[719], _056837_);
  xor g_115065_(out[122], out[714], _056838_);
  xor g_115066_(out[117], out[709], _056839_);
  xor g_115067_(out[112], out[704], _056840_);
  or g_115068_(_056826_, _056831_, _056841_);
  or g_115069_(_056827_, _056829_, _056842_);
  or g_115070_(_056832_, _056838_, _056843_);
  or g_115071_(_056842_, _056843_, _056844_);
  or g_115072_(_056830_, _056834_, _056845_);
  or g_115073_(_056839_, _056840_, _056846_);
  or g_115074_(_056845_, _056846_, _056848_);
  or g_115075_(_056844_, _056848_, _056849_);
  xor g_115076_(out[124], out[716], _056850_);
  or g_115077_(_056824_, _056850_, _056851_);
  or g_115078_(_056823_, _056835_, _056852_);
  or g_115079_(_056851_, _056852_, _056853_);
  or g_115080_(_056828_, _056833_, _056854_);
  or g_115081_(_056837_, _056854_, _056855_);
  or g_115082_(_056853_, _056855_, _056856_);
  or g_115083_(_056849_, _056856_, _056857_);
  or g_115084_(_056841_, _056857_, _056859_);
  not g_115085_(_056859_, _056860_);
  xor g_115086_(out[97], out[705], _056861_);
  and g_115087_(out[107], _049653_, _056862_);
  xor g_115088_(out[105], out[713], _056863_);
  xor g_115089_(out[96], out[704], _056864_);
  xor g_115090_(out[110], out[718], _056865_);
  xor g_115091_(out[100], out[708], _056866_);
  or g_115092_(_056865_, _056866_, _056867_);
  xor g_115093_(out[109], out[717], _056868_);
  xor g_115094_(out[99], out[707], _056870_);
  and g_115095_(_098140_, out[715], _056871_);
  xor g_115096_(out[102], out[710], _056872_);
  xor g_115097_(out[106], out[714], _056873_);
  xor g_115098_(out[101], out[709], _056874_);
  xor g_115099_(out[111], out[719], _056875_);
  xor g_115100_(out[104], out[712], _056876_);
  or g_115101_(_056868_, _056876_, _056877_);
  xor g_115102_(out[98], out[706], _056878_);
  or g_115103_(_056873_, _056878_, _056879_);
  or g_115104_(_056877_, _056879_, _056881_);
  or g_115105_(_056863_, _056870_, _056882_);
  or g_115106_(_056874_, _056882_, _056883_);
  or g_115107_(_056881_, _056883_, _056884_);
  or g_115108_(_056867_, _056884_, _056885_);
  xor g_115109_(out[108], out[716], _056886_);
  or g_115110_(_056871_, _056886_, _056887_);
  xor g_115111_(out[103], out[711], _056888_);
  or g_115112_(_056872_, _056888_, _056889_);
  or g_115113_(_056887_, _056889_, _056890_);
  or g_115114_(_056861_, _056862_, _056892_);
  or g_115115_(_056875_, _056892_, _056893_);
  or g_115116_(_056890_, _056893_, _056894_);
  or g_115117_(_056864_, _056894_, _056895_);
  or g_115118_(_056885_, _056895_, _056896_);
  xor g_115119_(out[87], out[711], _056897_);
  and g_115120_(_098129_, out[715], _056898_);
  xor g_115121_(out[94], out[718], _056899_);
  xor g_115122_(out[88], out[712], _056900_);
  xor g_115123_(out[81], out[705], _056901_);
  xor g_115124_(out[93], out[717], _056903_);
  xor g_115125_(out[89], out[713], _056904_);
  xor g_115126_(out[84], out[708], _056905_);
  xor g_115127_(out[82], out[706], _056906_);
  and g_115128_(out[91], _049653_, _056907_);
  xor g_115129_(out[83], out[707], _056908_);
  xor g_115130_(out[86], out[710], _056909_);
  xor g_115131_(out[95], out[719], _056910_);
  xor g_115132_(out[90], out[714], _056911_);
  xor g_115133_(out[85], out[709], _056912_);
  xor g_115134_(out[80], out[704], _056914_);
  or g_115135_(_056899_, _056905_, _056915_);
  or g_115136_(_056900_, _056903_, _056916_);
  or g_115137_(_056906_, _056911_, _056917_);
  or g_115138_(_056916_, _056917_, _056918_);
  or g_115139_(_056904_, _056908_, _056919_);
  or g_115140_(_056912_, _056914_, _056920_);
  or g_115141_(_056919_, _056920_, _056921_);
  or g_115142_(_056918_, _056921_, _056922_);
  xor g_115143_(out[92], out[716], _056923_);
  or g_115144_(_056898_, _056923_, _056925_);
  or g_115145_(_056897_, _056909_, _056926_);
  or g_115146_(_056925_, _056926_, _056927_);
  or g_115147_(_056901_, _056907_, _056928_);
  or g_115148_(_056910_, _056928_, _056929_);
  or g_115149_(_056927_, _056929_, _056930_);
  or g_115150_(_056922_, _056930_, _056931_);
  or g_115151_(_056915_, _056931_, _056932_);
  xor g_115152_(out[72], out[712], _056933_);
  xor g_115153_(out[69], out[709], _056934_);
  xor g_115154_(out[67], out[707], _056936_);
  xor g_115155_(out[78], out[718], _056937_);
  xor g_115156_(out[77], out[717], _056938_);
  xor g_115157_(out[66], out[706], _056939_);
  xor g_115158_(out[73], out[713], _056940_);
  xor g_115159_(out[70], out[710], _056941_);
  xor g_115160_(out[79], out[719], _056942_);
  xor g_115161_(out[74], out[714], _056943_);
  xor g_115162_(out[68], out[708], _056944_);
  xor g_115163_(out[64], out[704], _056945_);
  and g_115164_(_098118_, out[715], _056947_);
  and g_115165_(out[75], _049653_, _056948_);
  or g_115166_(_056933_, _056938_, _056949_);
  xor g_115167_(out[65], out[705], _056950_);
  or g_115168_(_056939_, _056943_, _056951_);
  or g_115169_(_056949_, _056951_, _056952_);
  or g_115170_(_056936_, _056940_, _056953_);
  or g_115171_(_056934_, _056953_, _056954_);
  or g_115172_(_056952_, _056954_, _056955_);
  or g_115173_(_056937_, _056944_, _056956_);
  or g_115174_(_056955_, _056956_, _056958_);
  xor g_115175_(out[76], out[716], _056959_);
  or g_115176_(_056947_, _056959_, _056960_);
  xor g_115177_(out[71], out[711], _056961_);
  or g_115178_(_056941_, _056961_, _056962_);
  or g_115179_(_056960_, _056962_, _056963_);
  or g_115180_(_056948_, _056950_, _056964_);
  or g_115181_(_056942_, _056964_, _056965_);
  or g_115182_(_056963_, _056965_, _056966_);
  or g_115183_(_056945_, _056966_, _056967_);
  or g_115184_(_056958_, _056967_, _056969_);
  not g_115185_(_056969_, _056970_);
  xor g_115186_(out[55], out[711], _056971_);
  and g_115187_(_098107_, out[715], _056972_);
  xor g_115188_(out[62], out[718], _056973_);
  xor g_115189_(out[56], out[712], _056974_);
  xor g_115190_(out[49], out[705], _056975_);
  xor g_115191_(out[61], out[717], _056976_);
  xor g_115192_(out[57], out[713], _056977_);
  xor g_115193_(out[52], out[708], _056978_);
  xor g_115194_(out[50], out[706], _056980_);
  and g_115195_(out[59], _049653_, _056981_);
  xor g_115196_(out[51], out[707], _056982_);
  xor g_115197_(out[54], out[710], _056983_);
  xor g_115198_(out[63], out[719], _056984_);
  xor g_115199_(out[58], out[714], _056985_);
  xor g_115200_(out[53], out[709], _056986_);
  xor g_115201_(out[48], out[704], _056987_);
  or g_115202_(_056973_, _056978_, _056988_);
  or g_115203_(_056974_, _056976_, _056989_);
  or g_115204_(_056980_, _056985_, _056991_);
  or g_115205_(_056989_, _056991_, _056992_);
  or g_115206_(_056977_, _056982_, _056993_);
  or g_115207_(_056986_, _056987_, _056994_);
  or g_115208_(_056993_, _056994_, _056995_);
  or g_115209_(_056992_, _056995_, _056996_);
  xor g_115210_(out[60], out[716], _056997_);
  or g_115211_(_056972_, _056997_, _056998_);
  or g_115212_(_056971_, _056983_, _056999_);
  or g_115213_(_056998_, _056999_, _057000_);
  or g_115214_(_056975_, _056981_, _057002_);
  or g_115215_(_056984_, _057002_, _057003_);
  or g_115216_(_057000_, _057003_, _057004_);
  or g_115217_(_056996_, _057004_, _057005_);
  or g_115218_(_056988_, _057005_, _057006_);
  xor g_115219_(out[42], out[714], _057007_);
  xor g_115220_(out[40], out[712], _057008_);
  xor g_115221_(out[33], out[705], _057009_);
  and g_115222_(_098096_, out[715], _057010_);
  and g_115223_(out[43], _049653_, _057011_);
  xor g_115224_(out[34], out[706], _057013_);
  xor g_115225_(out[37], out[709], _057014_);
  xor g_115226_(out[41], out[713], _057015_);
  xor g_115227_(out[44], out[716], _057016_);
  xor g_115228_(out[45], out[717], _057017_);
  xor g_115229_(out[47], out[719], _057018_);
  xor g_115230_(out[36], out[708], _057019_);
  xor g_115231_(out[38], out[710], _057020_);
  xor g_115232_(out[35], out[707], _057021_);
  xor g_115233_(out[32], out[704], _057022_);
  xor g_115234_(out[46], out[718], _057024_);
  or g_115235_(_057019_, _057024_, _057025_);
  or g_115236_(_057008_, _057017_, _057026_);
  or g_115237_(_057007_, _057013_, _057027_);
  or g_115238_(_057026_, _057027_, _057028_);
  or g_115239_(_057015_, _057021_, _057029_);
  or g_115240_(_057014_, _057022_, _057030_);
  or g_115241_(_057029_, _057030_, _057031_);
  or g_115242_(_057028_, _057031_, _057032_);
  or g_115243_(_057010_, _057016_, _057033_);
  xor g_115244_(out[39], out[711], _057035_);
  or g_115245_(_057020_, _057035_, _057036_);
  or g_115246_(_057033_, _057036_, _057037_);
  or g_115247_(_057009_, _057011_, _057038_);
  or g_115248_(_057018_, _057038_, _057039_);
  or g_115249_(_057037_, _057039_, _057040_);
  or g_115250_(_057032_, _057040_, _057041_);
  or g_115251_(_057025_, _057041_, _057042_);
  xor g_115252_(out[23], out[711], _057043_);
  and g_115253_(_098063_, out[715], _057044_);
  xor g_115254_(out[30], out[718], _057046_);
  xor g_115255_(out[24], out[712], _057047_);
  xor g_115256_(out[17], out[705], _057048_);
  xor g_115257_(out[29], out[717], _057049_);
  xor g_115258_(out[25], out[713], _057050_);
  xor g_115259_(out[20], out[708], _057051_);
  xor g_115260_(out[18], out[706], _057052_);
  and g_115261_(out[27], _049653_, _057053_);
  xor g_115262_(out[19], out[707], _057054_);
  xor g_115263_(out[22], out[710], _057055_);
  xor g_115264_(out[31], out[719], _057057_);
  xor g_115265_(out[26], out[714], _057058_);
  xor g_115266_(out[21], out[709], _057059_);
  xor g_115267_(out[16], out[704], _057060_);
  or g_115268_(_057046_, _057051_, _057061_);
  or g_115269_(_057047_, _057049_, _057062_);
  or g_115270_(_057052_, _057058_, _057063_);
  or g_115271_(_057062_, _057063_, _057064_);
  or g_115272_(_057050_, _057054_, _057065_);
  or g_115273_(_057059_, _057060_, _057066_);
  or g_115274_(_057065_, _057066_, _057068_);
  or g_115275_(_057064_, _057068_, _057069_);
  xor g_115276_(out[28], out[716], _057070_);
  or g_115277_(_057044_, _057070_, _057071_);
  or g_115278_(_057043_, _057055_, _057072_);
  or g_115279_(_057071_, _057072_, _057073_);
  or g_115280_(_057048_, _057053_, _057074_);
  or g_115281_(_057057_, _057074_, _057075_);
  or g_115282_(_057073_, _057075_, _057076_);
  or g_115283_(_057069_, _057076_, _057077_);
  or g_115284_(_057061_, _057077_, _057079_);
  and g_115285_(out[11], _049653_, _057080_);
  and g_115286_(_098041_, out[715], _057081_);
  xor g_115287_(out[8], out[712], _057082_);
  xor g_115288_(out[15], out[719], _057083_);
  xor g_115289_(out[1], out[705], _057084_);
  xor g_115290_(out[2], out[706], _057085_);
  xor g_115291_(out[4], out[708], _057086_);
  xor g_115292_(out[5], out[709], _057087_);
  xor g_115293_(out[9], out[713], _057088_);
  xor g_115294_(out[3], out[707], _057090_);
  xor g_115295_(out[14], out[718], _057091_);
  xor g_115296_(out[0], out[704], _057092_);
  xor g_115297_(out[10], out[714], _057093_);
  xor g_115298_(out[13], out[717], _057094_);
  or g_115299_(_057082_, _057094_, _057095_);
  xor g_115300_(out[6], out[710], _057096_);
  or g_115301_(_057085_, _057093_, _057097_);
  or g_115302_(_057095_, _057097_, _057098_);
  or g_115303_(_057088_, _057090_, _057099_);
  or g_115304_(_057087_, _057099_, _057101_);
  or g_115305_(_057098_, _057101_, _057102_);
  or g_115306_(_057086_, _057091_, _057103_);
  or g_115307_(_057102_, _057103_, _057104_);
  xor g_115308_(out[12], out[716], _057105_);
  or g_115309_(_057081_, _057105_, _057106_);
  xor g_115310_(out[7], out[711], _057107_);
  or g_115311_(_057096_, _057107_, _057108_);
  or g_115312_(_057106_, _057108_, _057109_);
  or g_115313_(_057080_, _057084_, _057110_);
  or g_115314_(_057083_, _057110_, _057112_);
  or g_115315_(_057109_, _057112_, _057113_);
  or g_115316_(_057092_, _057113_, _057114_);
  or g_115317_(_057104_, _057114_, _057115_);
  xor g_115318_(out[465], out[689], _057116_);
  and g_115319_(out[475], _049642_, _057117_);
  xor g_115320_(out[473], out[697], _057118_);
  xor g_115321_(out[464], out[688], _057119_);
  xor g_115322_(out[478], out[702], _057120_);
  xor g_115323_(out[468], out[692], _057121_);
  or g_115324_(_057120_, _057121_, _057123_);
  xor g_115325_(out[477], out[701], _057124_);
  xor g_115326_(out[467], out[691], _057125_);
  and g_115327_(_049499_, out[699], _057126_);
  xor g_115328_(out[470], out[694], _057127_);
  xor g_115329_(out[474], out[698], _057128_);
  xor g_115330_(out[469], out[693], _057129_);
  xor g_115331_(out[479], out[703], _057130_);
  xor g_115332_(out[472], out[696], _057131_);
  or g_115333_(_057124_, _057131_, _057132_);
  xor g_115334_(out[466], out[690], _057134_);
  or g_115335_(_057128_, _057134_, _057135_);
  or g_115336_(_057132_, _057135_, _057136_);
  or g_115337_(_057118_, _057125_, _057137_);
  or g_115338_(_057129_, _057137_, _057138_);
  or g_115339_(_057136_, _057138_, _057139_);
  or g_115340_(_057123_, _057139_, _057140_);
  xor g_115341_(out[476], out[700], _057141_);
  or g_115342_(_057126_, _057141_, _057142_);
  xor g_115343_(out[471], out[695], _057143_);
  or g_115344_(_057127_, _057143_, _057145_);
  or g_115345_(_057142_, _057145_, _057146_);
  or g_115346_(_057116_, _057117_, _057147_);
  or g_115347_(_057130_, _057147_, _057148_);
  or g_115348_(_057146_, _057148_, _057149_);
  or g_115349_(_057119_, _057149_, _057150_);
  or g_115350_(_057140_, _057150_, _057151_);
  xor g_115351_(out[455], out[695], _057152_);
  and g_115352_(_049477_, out[699], _057153_);
  xor g_115353_(out[462], out[702], _057154_);
  xor g_115354_(out[456], out[696], _057156_);
  xor g_115355_(out[449], out[689], _057157_);
  xor g_115356_(out[461], out[701], _057158_);
  xor g_115357_(out[457], out[697], _057159_);
  xor g_115358_(out[452], out[692], _057160_);
  xor g_115359_(out[450], out[690], _057161_);
  and g_115360_(out[459], _049642_, _057162_);
  xor g_115361_(out[451], out[691], _057163_);
  xor g_115362_(out[454], out[694], _057164_);
  xor g_115363_(out[463], out[703], _057165_);
  xor g_115364_(out[458], out[698], _057167_);
  xor g_115365_(out[453], out[693], _057168_);
  xor g_115366_(out[448], out[688], _057169_);
  or g_115367_(_057154_, _057160_, _057170_);
  or g_115368_(_057156_, _057158_, _057171_);
  or g_115369_(_057161_, _057167_, _057172_);
  or g_115370_(_057171_, _057172_, _057173_);
  or g_115371_(_057159_, _057163_, _057174_);
  or g_115372_(_057168_, _057169_, _057175_);
  or g_115373_(_057174_, _057175_, _057176_);
  or g_115374_(_057173_, _057176_, _057178_);
  xor g_115375_(out[460], out[700], _057179_);
  or g_115376_(_057153_, _057179_, _057180_);
  or g_115377_(_057152_, _057164_, _057181_);
  or g_115378_(_057180_, _057181_, _057182_);
  or g_115379_(_057157_, _057162_, _057183_);
  or g_115380_(_057165_, _057183_, _057184_);
  or g_115381_(_057182_, _057184_, _057185_);
  or g_115382_(_057178_, _057185_, _057186_);
  or g_115383_(_057170_, _057186_, _057187_);
  not g_115384_(_057187_, _057189_);
  xor g_115385_(out[433], out[689], _057190_);
  and g_115386_(_049466_, out[699], _057191_);
  and g_115387_(out[443], _049642_, _057192_);
  xor g_115388_(out[445], out[701], _057193_);
  xor g_115389_(out[442], out[698], _057194_);
  xor g_115390_(out[436], out[692], _057195_);
  xor g_115391_(out[446], out[702], _057196_);
  or g_115392_(_057195_, _057196_, _057197_);
  xor g_115393_(out[440], out[696], _057198_);
  xor g_115394_(out[432], out[688], _057200_);
  xor g_115395_(out[434], out[690], _057201_);
  xor g_115396_(out[441], out[697], _057202_);
  xor g_115397_(out[437], out[693], _057203_);
  xor g_115398_(out[435], out[691], _057204_);
  xor g_115399_(out[447], out[703], _057205_);
  xor g_115400_(out[438], out[694], _057206_);
  or g_115401_(_057193_, _057198_, _057207_);
  or g_115402_(_057194_, _057201_, _057208_);
  or g_115403_(_057207_, _057208_, _057209_);
  or g_115404_(_057202_, _057204_, _057211_);
  or g_115405_(_057200_, _057203_, _057212_);
  or g_115406_(_057211_, _057212_, _057213_);
  or g_115407_(_057209_, _057213_, _057214_);
  xor g_115408_(out[444], out[700], _057215_);
  or g_115409_(_057191_, _057215_, _057216_);
  xor g_115410_(out[439], out[695], _057217_);
  or g_115411_(_057206_, _057217_, _057218_);
  or g_115412_(_057216_, _057218_, _057219_);
  or g_115413_(_057190_, _057192_, _057220_);
  or g_115414_(_057205_, _057220_, _057222_);
  or g_115415_(_057219_, _057222_, _057223_);
  or g_115416_(_057214_, _057223_, _057224_);
  or g_115417_(_057197_, _057224_, _057225_);
  not g_115418_(_057225_, _057226_);
  xor g_115419_(out[423], out[695], _057227_);
  and g_115420_(_049455_, out[699], _057228_);
  xor g_115421_(out[430], out[702], _057229_);
  xor g_115422_(out[424], out[696], _057230_);
  xor g_115423_(out[417], out[689], _057231_);
  xor g_115424_(out[429], out[701], _057233_);
  xor g_115425_(out[425], out[697], _057234_);
  xor g_115426_(out[420], out[692], _057235_);
  xor g_115427_(out[418], out[690], _057236_);
  and g_115428_(out[427], _049642_, _057237_);
  xor g_115429_(out[419], out[691], _057238_);
  xor g_115430_(out[422], out[694], _057239_);
  xor g_115431_(out[431], out[703], _057240_);
  xor g_115432_(out[426], out[698], _057241_);
  xor g_115433_(out[421], out[693], _057242_);
  xor g_115434_(out[416], out[688], _057244_);
  or g_115435_(_057229_, _057235_, _057245_);
  or g_115436_(_057230_, _057233_, _057246_);
  or g_115437_(_057236_, _057241_, _057247_);
  or g_115438_(_057246_, _057247_, _057248_);
  or g_115439_(_057234_, _057238_, _057249_);
  or g_115440_(_057242_, _057244_, _057250_);
  or g_115441_(_057249_, _057250_, _057251_);
  or g_115442_(_057248_, _057251_, _057252_);
  xor g_115443_(out[428], out[700], _057253_);
  or g_115444_(_057228_, _057253_, _057255_);
  or g_115445_(_057227_, _057239_, _057256_);
  or g_115446_(_057255_, _057256_, _057257_);
  or g_115447_(_057231_, _057237_, _057258_);
  or g_115448_(_057240_, _057258_, _057259_);
  or g_115449_(_057257_, _057259_, _057260_);
  or g_115450_(_057252_, _057260_, _057261_);
  or g_115451_(_057245_, _057261_, _057262_);
  xor g_115452_(out[410], out[698], _057263_);
  xor g_115453_(out[402], out[690], _057264_);
  xor g_115454_(out[401], out[689], _057266_);
  and g_115455_(_049444_, out[699], _057267_);
  and g_115456_(out[411], _049642_, _057268_);
  xor g_115457_(out[413], out[701], _057269_);
  xor g_115458_(out[403], out[691], _057270_);
  xor g_115459_(out[414], out[702], _057271_);
  xor g_115460_(out[412], out[700], _057272_);
  xor g_115461_(out[408], out[696], _057273_);
  xor g_115462_(out[415], out[703], _057274_);
  xor g_115463_(out[405], out[693], _057275_);
  xor g_115464_(out[406], out[694], _057277_);
  xor g_115465_(out[400], out[688], _057278_);
  xor g_115466_(out[404], out[692], _057279_);
  or g_115467_(_057269_, _057273_, _057280_);
  xor g_115468_(out[409], out[697], _057281_);
  or g_115469_(_057263_, _057264_, _057282_);
  or g_115470_(_057280_, _057282_, _057283_);
  or g_115471_(_057270_, _057281_, _057284_);
  or g_115472_(_057275_, _057284_, _057285_);
  or g_115473_(_057283_, _057285_, _057286_);
  or g_115474_(_057271_, _057279_, _057288_);
  or g_115475_(_057286_, _057288_, _057289_);
  or g_115476_(_057267_, _057272_, _057290_);
  xor g_115477_(out[407], out[695], _057291_);
  or g_115478_(_057277_, _057291_, _057292_);
  or g_115479_(_057290_, _057292_, _057293_);
  or g_115480_(_057266_, _057268_, _057294_);
  or g_115481_(_057274_, _057294_, _057295_);
  or g_115482_(_057293_, _057295_, _057296_);
  or g_115483_(_057278_, _057296_, _057297_);
  or g_115484_(_057289_, _057297_, _057299_);
  xor g_115485_(out[391], out[695], _057300_);
  and g_115486_(_049433_, out[699], _057301_);
  xor g_115487_(out[398], out[702], _057302_);
  xor g_115488_(out[392], out[696], _057303_);
  xor g_115489_(out[385], out[689], _057304_);
  xor g_115490_(out[397], out[701], _057305_);
  xor g_115491_(out[393], out[697], _057306_);
  xor g_115492_(out[388], out[692], _057307_);
  xor g_115493_(out[386], out[690], _057308_);
  and g_115494_(out[395], _049642_, _057310_);
  xor g_115495_(out[387], out[691], _057311_);
  xor g_115496_(out[390], out[694], _057312_);
  xor g_115497_(out[399], out[703], _057313_);
  xor g_115498_(out[394], out[698], _057314_);
  xor g_115499_(out[389], out[693], _057315_);
  xor g_115500_(out[384], out[688], _057316_);
  or g_115501_(_057302_, _057307_, _057317_);
  or g_115502_(_057303_, _057305_, _057318_);
  or g_115503_(_057308_, _057314_, _057319_);
  or g_115504_(_057318_, _057319_, _057321_);
  or g_115505_(_057306_, _057311_, _057322_);
  or g_115506_(_057315_, _057316_, _057323_);
  or g_115507_(_057322_, _057323_, _057324_);
  or g_115508_(_057321_, _057324_, _057325_);
  xor g_115509_(out[396], out[700], _057326_);
  or g_115510_(_057301_, _057326_, _057327_);
  or g_115511_(_057300_, _057312_, _057328_);
  or g_115512_(_057327_, _057328_, _057329_);
  or g_115513_(_057304_, _057310_, _057330_);
  or g_115514_(_057313_, _057330_, _057332_);
  or g_115515_(_057329_, _057332_, _057333_);
  or g_115516_(_057325_, _057333_, _057334_);
  or g_115517_(_057317_, _057334_, _057335_);
  xor g_115518_(out[369], out[689], _057336_);
  and g_115519_(_049422_, out[699], _057337_);
  and g_115520_(out[379], _049642_, _057338_);
  xor g_115521_(out[376], out[696], _057339_);
  xor g_115522_(out[378], out[698], _057340_);
  xor g_115523_(out[370], out[690], _057341_);
  xor g_115524_(out[372], out[692], _057343_);
  xor g_115525_(out[381], out[701], _057344_);
  xor g_115526_(out[377], out[697], _057345_);
  xor g_115527_(out[371], out[691], _057346_);
  xor g_115528_(out[373], out[693], _057347_);
  xor g_115529_(out[382], out[702], _057348_);
  xor g_115530_(out[368], out[688], _057349_);
  xor g_115531_(out[383], out[703], _057350_);
  or g_115532_(_057339_, _057344_, _057351_);
  xor g_115533_(out[374], out[694], _057352_);
  or g_115534_(_057340_, _057341_, _057354_);
  or g_115535_(_057351_, _057354_, _057355_);
  or g_115536_(_057345_, _057346_, _057356_);
  or g_115537_(_057347_, _057356_, _057357_);
  or g_115538_(_057355_, _057357_, _057358_);
  or g_115539_(_057343_, _057348_, _057359_);
  or g_115540_(_057358_, _057359_, _057360_);
  xor g_115541_(out[380], out[700], _057361_);
  or g_115542_(_057337_, _057361_, _057362_);
  xor g_115543_(out[375], out[695], _057363_);
  or g_115544_(_057352_, _057363_, _057365_);
  or g_115545_(_057362_, _057365_, _057366_);
  or g_115546_(_057336_, _057338_, _057367_);
  or g_115547_(_057350_, _057367_, _057368_);
  or g_115548_(_057366_, _057368_, _057369_);
  or g_115549_(_057349_, _057369_, _057370_);
  or g_115550_(_057360_, _057370_, _057371_);
  xor g_115551_(out[359], out[695], _057372_);
  and g_115552_(_049411_, out[699], _057373_);
  xor g_115553_(out[366], out[702], _057374_);
  xor g_115554_(out[360], out[696], _057376_);
  xor g_115555_(out[353], out[689], _057377_);
  xor g_115556_(out[365], out[701], _057378_);
  xor g_115557_(out[361], out[697], _057379_);
  xor g_115558_(out[356], out[692], _057380_);
  xor g_115559_(out[354], out[690], _057381_);
  and g_115560_(out[363], _049642_, _057382_);
  xor g_115561_(out[355], out[691], _057383_);
  xor g_115562_(out[358], out[694], _057384_);
  xor g_115563_(out[367], out[703], _057385_);
  xor g_115564_(out[362], out[698], _057387_);
  xor g_115565_(out[357], out[693], _057388_);
  xor g_115566_(out[352], out[688], _057389_);
  or g_115567_(_057374_, _057380_, _057390_);
  or g_115568_(_057376_, _057378_, _057391_);
  or g_115569_(_057381_, _057387_, _057392_);
  or g_115570_(_057391_, _057392_, _057393_);
  or g_115571_(_057379_, _057383_, _057394_);
  or g_115572_(_057388_, _057389_, _057395_);
  or g_115573_(_057394_, _057395_, _057396_);
  or g_115574_(_057393_, _057396_, _057398_);
  xor g_115575_(out[364], out[700], _057399_);
  or g_115576_(_057373_, _057399_, _057400_);
  or g_115577_(_057372_, _057384_, _057401_);
  or g_115578_(_057400_, _057401_, _057402_);
  or g_115579_(_057377_, _057382_, _057403_);
  or g_115580_(_057385_, _057403_, _057404_);
  or g_115581_(_057402_, _057404_, _057405_);
  or g_115582_(_057398_, _057405_, _057406_);
  or g_115583_(_057390_, _057406_, _057407_);
  xor g_115584_(out[346], out[698], _057409_);
  xor g_115585_(out[338], out[690], _057410_);
  xor g_115586_(out[337], out[689], _057411_);
  and g_115587_(_049400_, out[699], _057412_);
  and g_115588_(out[347], _049642_, _057413_);
  xor g_115589_(out[349], out[701], _057414_);
  xor g_115590_(out[339], out[691], _057415_);
  xor g_115591_(out[350], out[702], _057416_);
  xor g_115592_(out[348], out[700], _057417_);
  xor g_115593_(out[344], out[696], _057418_);
  xor g_115594_(out[351], out[703], _057420_);
  xor g_115595_(out[341], out[693], _057421_);
  xor g_115596_(out[342], out[694], _057422_);
  xor g_115597_(out[336], out[688], _057423_);
  xor g_115598_(out[340], out[692], _057424_);
  or g_115599_(_057414_, _057418_, _057425_);
  xor g_115600_(out[345], out[697], _057426_);
  or g_115601_(_057409_, _057410_, _057427_);
  or g_115602_(_057425_, _057427_, _057428_);
  or g_115603_(_057415_, _057426_, _057429_);
  or g_115604_(_057421_, _057429_, _057431_);
  or g_115605_(_057428_, _057431_, _057432_);
  or g_115606_(_057416_, _057424_, _057433_);
  or g_115607_(_057432_, _057433_, _057434_);
  or g_115608_(_057412_, _057417_, _057435_);
  xor g_115609_(out[343], out[695], _057436_);
  or g_115610_(_057422_, _057436_, _057437_);
  or g_115611_(_057435_, _057437_, _057438_);
  or g_115612_(_057411_, _057413_, _057439_);
  or g_115613_(_057420_, _057439_, _057440_);
  or g_115614_(_057438_, _057440_, _057442_);
  or g_115615_(_057423_, _057442_, _057443_);
  or g_115616_(_057434_, _057443_, _057444_);
  xor g_115617_(out[327], out[695], _057445_);
  and g_115618_(_098294_, out[699], _057446_);
  xor g_115619_(out[334], out[702], _057447_);
  xor g_115620_(out[328], out[696], _057448_);
  xor g_115621_(out[321], out[689], _057449_);
  xor g_115622_(out[333], out[701], _057450_);
  xor g_115623_(out[329], out[697], _057451_);
  xor g_115624_(out[324], out[692], _057453_);
  xor g_115625_(out[322], out[690], _057454_);
  and g_115626_(out[331], _049642_, _057455_);
  xor g_115627_(out[323], out[691], _057456_);
  xor g_115628_(out[326], out[694], _057457_);
  xor g_115629_(out[335], out[703], _057458_);
  xor g_115630_(out[330], out[698], _057459_);
  xor g_115631_(out[325], out[693], _057460_);
  xor g_115632_(out[320], out[688], _057461_);
  or g_115633_(_057447_, _057453_, _057462_);
  or g_115634_(_057448_, _057450_, _057464_);
  or g_115635_(_057454_, _057459_, _057465_);
  or g_115636_(_057464_, _057465_, _057466_);
  or g_115637_(_057451_, _057456_, _057467_);
  or g_115638_(_057460_, _057461_, _057468_);
  or g_115639_(_057467_, _057468_, _057469_);
  or g_115640_(_057466_, _057469_, _057470_);
  xor g_115641_(out[332], out[700], _057471_);
  or g_115642_(_057446_, _057471_, _057472_);
  or g_115643_(_057445_, _057457_, _057473_);
  or g_115644_(_057472_, _057473_, _057475_);
  or g_115645_(_057449_, _057455_, _057476_);
  or g_115646_(_057458_, _057476_, _057477_);
  or g_115647_(_057475_, _057477_, _057478_);
  or g_115648_(_057470_, _057478_, _057479_);
  or g_115649_(_057462_, _057479_, _057480_);
  xor g_115650_(out[316], out[700], _057481_);
  and g_115651_(_098283_, out[699], _057482_);
  xor g_115652_(out[312], out[696], _057483_);
  xor g_115653_(out[310], out[694], _057484_);
  xor g_115654_(out[317], out[701], _057486_);
  xor g_115655_(out[318], out[702], _057487_);
  xor g_115656_(out[306], out[690], _057488_);
  xor g_115657_(out[313], out[697], _057489_);
  xor g_115658_(out[309], out[693], _057490_);
  xor g_115659_(out[305], out[689], _057491_);
  and g_115660_(out[315], _049642_, _057492_);
  or g_115661_(_057483_, _057486_, _057493_);
  xor g_115662_(out[319], out[703], _057494_);
  xor g_115663_(out[314], out[698], _057495_);
  xor g_115664_(out[308], out[692], _057497_);
  xor g_115665_(out[307], out[691], _057498_);
  xor g_115666_(out[304], out[688], _057499_);
  or g_115667_(_057488_, _057495_, _057500_);
  or g_115668_(_057493_, _057500_, _057501_);
  or g_115669_(_057489_, _057498_, _057502_);
  or g_115670_(_057490_, _057502_, _057503_);
  or g_115671_(_057501_, _057503_, _057504_);
  or g_115672_(_057487_, _057497_, _057505_);
  or g_115673_(_057504_, _057505_, _057506_);
  or g_115674_(_057481_, _057482_, _057508_);
  xor g_115675_(out[311], out[695], _057509_);
  or g_115676_(_057484_, _057509_, _057510_);
  or g_115677_(_057508_, _057510_, _057511_);
  or g_115678_(_057491_, _057492_, _057512_);
  or g_115679_(_057494_, _057512_, _057513_);
  or g_115680_(_057511_, _057513_, _057514_);
  or g_115681_(_057499_, _057514_, _057515_);
  or g_115682_(_057506_, _057515_, _057516_);
  xor g_115683_(out[295], out[695], _057517_);
  and g_115684_(_098272_, out[699], _057519_);
  xor g_115685_(out[302], out[702], _057520_);
  xor g_115686_(out[296], out[696], _057521_);
  xor g_115687_(out[289], out[689], _057522_);
  xor g_115688_(out[301], out[701], _057523_);
  xor g_115689_(out[297], out[697], _057524_);
  xor g_115690_(out[292], out[692], _057525_);
  xor g_115691_(out[290], out[690], _057526_);
  and g_115692_(out[299], _049642_, _057527_);
  xor g_115693_(out[291], out[691], _057528_);
  xor g_115694_(out[294], out[694], _057530_);
  xor g_115695_(out[303], out[703], _057531_);
  xor g_115696_(out[298], out[698], _057532_);
  xor g_115697_(out[293], out[693], _057533_);
  xor g_115698_(out[288], out[688], _057534_);
  or g_115699_(_057520_, _057525_, _057535_);
  or g_115700_(_057521_, _057523_, _057536_);
  or g_115701_(_057526_, _057532_, _057537_);
  or g_115702_(_057536_, _057537_, _057538_);
  or g_115703_(_057524_, _057528_, _057539_);
  or g_115704_(_057533_, _057534_, _057541_);
  or g_115705_(_057539_, _057541_, _057542_);
  or g_115706_(_057538_, _057542_, _057543_);
  xor g_115707_(out[300], out[700], _057544_);
  or g_115708_(_057519_, _057544_, _057545_);
  or g_115709_(_057517_, _057530_, _057546_);
  or g_115710_(_057545_, _057546_, _057547_);
  or g_115711_(_057522_, _057527_, _057548_);
  or g_115712_(_057531_, _057548_, _057549_);
  or g_115713_(_057547_, _057549_, _057550_);
  or g_115714_(_057543_, _057550_, _057552_);
  or g_115715_(_057535_, _057552_, _057553_);
  xor g_115716_(out[273], out[689], _057554_);
  and g_115717_(_098261_, out[699], _057555_);
  and g_115718_(out[283], _049642_, _057556_);
  xor g_115719_(out[281], out[697], _057557_);
  xor g_115720_(out[272], out[688], _057558_);
  xor g_115721_(out[286], out[702], _057559_);
  xor g_115722_(out[276], out[692], _057560_);
  or g_115723_(_057559_, _057560_, _057561_);
  xor g_115724_(out[285], out[701], _057563_);
  xor g_115725_(out[275], out[691], _057564_);
  xor g_115726_(out[284], out[700], _057565_);
  xor g_115727_(out[278], out[694], _057566_);
  xor g_115728_(out[282], out[698], _057567_);
  xor g_115729_(out[277], out[693], _057568_);
  xor g_115730_(out[287], out[703], _057569_);
  xor g_115731_(out[280], out[696], _057570_);
  or g_115732_(_057563_, _057570_, _057571_);
  xor g_115733_(out[274], out[690], _057572_);
  or g_115734_(_057567_, _057572_, _057574_);
  or g_115735_(_057571_, _057574_, _057575_);
  or g_115736_(_057557_, _057564_, _057576_);
  or g_115737_(_057568_, _057576_, _057577_);
  or g_115738_(_057575_, _057577_, _057578_);
  or g_115739_(_057561_, _057578_, _057579_);
  or g_115740_(_057555_, _057565_, _057580_);
  xor g_115741_(out[279], out[695], _057581_);
  or g_115742_(_057566_, _057581_, _057582_);
  or g_115743_(_057580_, _057582_, _057583_);
  or g_115744_(_057554_, _057556_, _057585_);
  or g_115745_(_057569_, _057585_, _057586_);
  or g_115746_(_057583_, _057586_, _057587_);
  or g_115747_(_057558_, _057587_, _057588_);
  or g_115748_(_057579_, _057588_, _057589_);
  xor g_115749_(out[263], out[695], _057590_);
  and g_115750_(_098250_, out[699], _057591_);
  xor g_115751_(out[270], out[702], _057592_);
  xor g_115752_(out[264], out[696], _057593_);
  xor g_115753_(out[257], out[689], _057594_);
  xor g_115754_(out[269], out[701], _057596_);
  xor g_115755_(out[265], out[697], _057597_);
  xor g_115756_(out[260], out[692], _057598_);
  xor g_115757_(out[258], out[690], _057599_);
  and g_115758_(out[267], _049642_, _057600_);
  xor g_115759_(out[259], out[691], _057601_);
  xor g_115760_(out[262], out[694], _057602_);
  xor g_115761_(out[271], out[703], _057603_);
  xor g_115762_(out[266], out[698], _057604_);
  xor g_115763_(out[261], out[693], _057605_);
  xor g_115764_(out[256], out[688], _057607_);
  or g_115765_(_057592_, _057598_, _057608_);
  or g_115766_(_057593_, _057596_, _057609_);
  or g_115767_(_057599_, _057604_, _057610_);
  or g_115768_(_057609_, _057610_, _057611_);
  or g_115769_(_057597_, _057601_, _057612_);
  or g_115770_(_057605_, _057607_, _057613_);
  or g_115771_(_057612_, _057613_, _057614_);
  or g_115772_(_057611_, _057614_, _057615_);
  xor g_115773_(out[268], out[700], _057616_);
  or g_115774_(_057591_, _057616_, _057618_);
  or g_115775_(_057590_, _057602_, _057619_);
  or g_115776_(_057618_, _057619_, _057620_);
  or g_115777_(_057594_, _057600_, _057621_);
  or g_115778_(_057603_, _057621_, _057622_);
  or g_115779_(_057620_, _057622_, _057623_);
  or g_115780_(_057615_, _057623_, _057624_);
  or g_115781_(_057608_, _057624_, _057625_);
  not g_115782_(_057625_, _057626_);
  xor g_115783_(out[241], out[689], _057627_);
  and g_115784_(out[251], _049642_, _057629_);
  xor g_115785_(out[254], out[702], _057630_);
  xor g_115786_(out[243], out[691], _057631_);
  xor g_115787_(out[244], out[692], _057632_);
  xor g_115788_(out[242], out[690], _057633_);
  xor g_115789_(out[249], out[697], _057634_);
  xor g_115790_(out[240], out[688], _057635_);
  and g_115791_(_098239_, out[699], _057636_);
  xor g_115792_(out[246], out[694], _057637_);
  xor g_115793_(out[250], out[698], _057638_);
  xor g_115794_(out[245], out[693], _057640_);
  xor g_115795_(out[255], out[703], _057641_);
  xor g_115796_(out[253], out[701], _057642_);
  xor g_115797_(out[248], out[696], _057643_);
  or g_115798_(_057630_, _057632_, _057644_);
  or g_115799_(_057642_, _057643_, _057645_);
  or g_115800_(_057633_, _057638_, _057646_);
  or g_115801_(_057645_, _057646_, _057647_);
  or g_115802_(_057631_, _057634_, _057648_);
  or g_115803_(_057635_, _057640_, _057649_);
  or g_115804_(_057648_, _057649_, _057651_);
  or g_115805_(_057647_, _057651_, _057652_);
  xor g_115806_(out[252], out[700], _057653_);
  or g_115807_(_057636_, _057653_, _057654_);
  xor g_115808_(out[247], out[695], _057655_);
  or g_115809_(_057637_, _057655_, _057656_);
  or g_115810_(_057654_, _057656_, _057657_);
  or g_115811_(_057627_, _057629_, _057658_);
  or g_115812_(_057641_, _057658_, _057659_);
  or g_115813_(_057657_, _057659_, _057660_);
  or g_115814_(_057652_, _057660_, _057662_);
  or g_115815_(_057644_, _057662_, _057663_);
  xor g_115816_(out[231], out[695], _057664_);
  and g_115817_(_098228_, out[699], _057665_);
  xor g_115818_(out[238], out[702], _057666_);
  xor g_115819_(out[232], out[696], _057667_);
  xor g_115820_(out[225], out[689], _057668_);
  xor g_115821_(out[237], out[701], _057669_);
  xor g_115822_(out[233], out[697], _057670_);
  xor g_115823_(out[228], out[692], _057671_);
  xor g_115824_(out[226], out[690], _057673_);
  and g_115825_(out[235], _049642_, _057674_);
  xor g_115826_(out[227], out[691], _057675_);
  xor g_115827_(out[230], out[694], _057676_);
  xor g_115828_(out[239], out[703], _057677_);
  xor g_115829_(out[234], out[698], _057678_);
  xor g_115830_(out[229], out[693], _057679_);
  xor g_115831_(out[224], out[688], _057680_);
  or g_115832_(_057666_, _057671_, _057681_);
  or g_115833_(_057667_, _057669_, _057682_);
  or g_115834_(_057673_, _057678_, _057684_);
  or g_115835_(_057682_, _057684_, _057685_);
  or g_115836_(_057670_, _057675_, _057686_);
  or g_115837_(_057679_, _057680_, _057687_);
  or g_115838_(_057686_, _057687_, _057688_);
  or g_115839_(_057685_, _057688_, _057689_);
  xor g_115840_(out[236], out[700], _057690_);
  or g_115841_(_057665_, _057690_, _057691_);
  or g_115842_(_057664_, _057676_, _057692_);
  or g_115843_(_057691_, _057692_, _057693_);
  or g_115844_(_057668_, _057674_, _057695_);
  or g_115845_(_057677_, _057695_, _057696_);
  or g_115846_(_057693_, _057696_, _057697_);
  or g_115847_(_057689_, _057697_, _057698_);
  or g_115848_(_057681_, _057698_, _057699_);
  xor g_115849_(out[209], out[689], _057700_);
  and g_115850_(out[219], _049642_, _057701_);
  xor g_115851_(out[217], out[697], _057702_);
  xor g_115852_(out[208], out[688], _057703_);
  xor g_115853_(out[222], out[702], _057704_);
  xor g_115854_(out[212], out[692], _057706_);
  or g_115855_(_057704_, _057706_, _057707_);
  xor g_115856_(out[221], out[701], _057708_);
  xor g_115857_(out[211], out[691], _057709_);
  and g_115858_(_098217_, out[699], _057710_);
  xor g_115859_(out[214], out[694], _057711_);
  xor g_115860_(out[218], out[698], _057712_);
  xor g_115861_(out[213], out[693], _057713_);
  xor g_115862_(out[223], out[703], _057714_);
  xor g_115863_(out[216], out[696], _057715_);
  or g_115864_(_057708_, _057715_, _057717_);
  xor g_115865_(out[210], out[690], _057718_);
  or g_115866_(_057712_, _057718_, _057719_);
  or g_115867_(_057717_, _057719_, _057720_);
  or g_115868_(_057702_, _057709_, _057721_);
  or g_115869_(_057713_, _057721_, _057722_);
  or g_115870_(_057720_, _057722_, _057723_);
  or g_115871_(_057707_, _057723_, _057724_);
  xor g_115872_(out[220], out[700], _057725_);
  or g_115873_(_057710_, _057725_, _057726_);
  xor g_115874_(out[215], out[695], _057728_);
  or g_115875_(_057711_, _057728_, _057729_);
  or g_115876_(_057726_, _057729_, _057730_);
  or g_115877_(_057700_, _057701_, _057731_);
  or g_115878_(_057714_, _057731_, _057732_);
  or g_115879_(_057730_, _057732_, _057733_);
  or g_115880_(_057703_, _057733_, _057734_);
  or g_115881_(_057724_, _057734_, _057735_);
  xor g_115882_(out[199], out[695], _057736_);
  and g_115883_(_098206_, out[699], _057737_);
  xor g_115884_(out[206], out[702], _057739_);
  xor g_115885_(out[200], out[696], _057740_);
  xor g_115886_(out[193], out[689], _057741_);
  xor g_115887_(out[205], out[701], _057742_);
  xor g_115888_(out[201], out[697], _057743_);
  xor g_115889_(out[196], out[692], _057744_);
  xor g_115890_(out[194], out[690], _057745_);
  and g_115891_(out[203], _049642_, _057746_);
  xor g_115892_(out[195], out[691], _057747_);
  xor g_115893_(out[198], out[694], _057748_);
  xor g_115894_(out[207], out[703], _057750_);
  xor g_115895_(out[202], out[698], _057751_);
  xor g_115896_(out[197], out[693], _057752_);
  xor g_115897_(out[192], out[688], _057753_);
  or g_115898_(_057739_, _057744_, _057754_);
  or g_115899_(_057740_, _057742_, _057755_);
  or g_115900_(_057745_, _057751_, _057756_);
  or g_115901_(_057755_, _057756_, _057757_);
  or g_115902_(_057743_, _057747_, _057758_);
  or g_115903_(_057752_, _057753_, _057759_);
  or g_115904_(_057758_, _057759_, _057761_);
  or g_115905_(_057757_, _057761_, _057762_);
  xor g_115906_(out[204], out[700], _057763_);
  or g_115907_(_057737_, _057763_, _057764_);
  or g_115908_(_057736_, _057748_, _057765_);
  or g_115909_(_057764_, _057765_, _057766_);
  or g_115910_(_057741_, _057746_, _057767_);
  or g_115911_(_057750_, _057767_, _057768_);
  or g_115912_(_057766_, _057768_, _057769_);
  or g_115913_(_057762_, _057769_, _057770_);
  or g_115914_(_057754_, _057770_, _057772_);
  xor g_115915_(out[189], out[701], _057773_);
  xor g_115916_(out[178], out[690], _057774_);
  xor g_115917_(out[181], out[693], _057775_);
  xor g_115918_(out[185], out[697], _057776_);
  xor g_115919_(out[180], out[692], _057777_);
  xor g_115920_(out[184], out[696], _057778_);
  xor g_115921_(out[190], out[702], _057779_);
  xor g_115922_(out[182], out[694], _057780_);
  xor g_115923_(out[191], out[703], _057781_);
  xor g_115924_(out[186], out[698], _057783_);
  xor g_115925_(out[176], out[688], _057784_);
  xor g_115926_(out[179], out[691], _057785_);
  and g_115927_(_098195_, out[699], _057786_);
  and g_115928_(out[187], _049642_, _057787_);
  xor g_115929_(out[177], out[689], _057788_);
  or g_115930_(_057777_, _057779_, _057789_);
  or g_115931_(_057773_, _057778_, _057790_);
  or g_115932_(_057774_, _057783_, _057791_);
  or g_115933_(_057790_, _057791_, _057792_);
  or g_115934_(_057776_, _057785_, _057794_);
  or g_115935_(_057775_, _057784_, _057795_);
  or g_115936_(_057794_, _057795_, _057796_);
  or g_115937_(_057792_, _057796_, _057797_);
  xor g_115938_(out[188], out[700], _057798_);
  or g_115939_(_057786_, _057798_, _057799_);
  xor g_115940_(out[183], out[695], _057800_);
  or g_115941_(_057780_, _057800_, _057801_);
  or g_115942_(_057799_, _057801_, _057802_);
  or g_115943_(_057787_, _057788_, _057803_);
  or g_115944_(_057781_, _057803_, _057805_);
  or g_115945_(_057802_, _057805_, _057806_);
  or g_115946_(_057797_, _057806_, _057807_);
  or g_115947_(_057789_, _057807_, _057808_);
  not g_115948_(_057808_, _057809_);
  xor g_115949_(out[167], out[695], _057810_);
  and g_115950_(_098184_, out[699], _057811_);
  xor g_115951_(out[174], out[702], _057812_);
  xor g_115952_(out[168], out[696], _057813_);
  xor g_115953_(out[161], out[689], _057814_);
  xor g_115954_(out[173], out[701], _057816_);
  xor g_115955_(out[169], out[697], _057817_);
  xor g_115956_(out[164], out[692], _057818_);
  xor g_115957_(out[162], out[690], _057819_);
  and g_115958_(out[171], _049642_, _057820_);
  xor g_115959_(out[163], out[691], _057821_);
  xor g_115960_(out[166], out[694], _057822_);
  xor g_115961_(out[175], out[703], _057823_);
  xor g_115962_(out[170], out[698], _057824_);
  xor g_115963_(out[165], out[693], _057825_);
  xor g_115964_(out[160], out[688], _057827_);
  or g_115965_(_057812_, _057818_, _057828_);
  not g_115966_(_057828_, _057829_);
  or g_115967_(_057813_, _057816_, _057830_);
  or g_115968_(_057819_, _057824_, _057831_);
  or g_115969_(_057830_, _057831_, _057832_);
  or g_115970_(_057817_, _057821_, _057833_);
  or g_115971_(_057825_, _057827_, _057834_);
  or g_115972_(_057833_, _057834_, _057835_);
  or g_115973_(_057832_, _057835_, _057836_);
  xor g_115974_(out[172], out[700], _057838_);
  or g_115975_(_057811_, _057838_, _057839_);
  or g_115976_(_057810_, _057822_, _057840_);
  or g_115977_(_057839_, _057840_, _057841_);
  or g_115978_(_057814_, _057820_, _057842_);
  or g_115979_(_057823_, _057842_, _057843_);
  or g_115980_(_057841_, _057843_, _057844_);
  or g_115981_(_057836_, _057844_, _057845_);
  not g_115982_(_057845_, _057846_);
  and g_115983_(_057829_, _057846_, _057847_);
  not g_115984_(_057847_, _057849_);
  xor g_115985_(out[145], out[689], _057850_);
  and g_115986_(out[155], _049642_, _057851_);
  xor g_115987_(out[153], out[697], _057852_);
  xor g_115988_(out[144], out[688], _057853_);
  xor g_115989_(out[158], out[702], _057854_);
  xor g_115990_(out[148], out[692], _057855_);
  or g_115991_(_057854_, _057855_, _057856_);
  xor g_115992_(out[157], out[701], _057857_);
  xor g_115993_(out[147], out[691], _057858_);
  and g_115994_(_098173_, out[699], _057860_);
  xor g_115995_(out[150], out[694], _057861_);
  xor g_115996_(out[154], out[698], _057862_);
  xor g_115997_(out[149], out[693], _057863_);
  xor g_115998_(out[159], out[703], _057864_);
  xor g_115999_(out[152], out[696], _057865_);
  or g_116000_(_057857_, _057865_, _057866_);
  xor g_116001_(out[146], out[690], _057867_);
  or g_116002_(_057862_, _057867_, _057868_);
  or g_116003_(_057866_, _057868_, _057869_);
  or g_116004_(_057852_, _057858_, _057871_);
  or g_116005_(_057863_, _057871_, _057872_);
  or g_116006_(_057869_, _057872_, _057873_);
  or g_116007_(_057856_, _057873_, _057874_);
  xor g_116008_(out[156], out[700], _057875_);
  or g_116009_(_057860_, _057875_, _057876_);
  xor g_116010_(out[151], out[695], _057877_);
  or g_116011_(_057861_, _057877_, _057878_);
  or g_116012_(_057876_, _057878_, _057879_);
  or g_116013_(_057850_, _057851_, _057880_);
  or g_116014_(_057864_, _057880_, _057882_);
  or g_116015_(_057879_, _057882_, _057883_);
  or g_116016_(_057853_, _057883_, _057884_);
  or g_116017_(_057874_, _057884_, _057885_);
  xor g_116018_(out[135], out[695], _057886_);
  and g_116019_(_098162_, out[699], _057887_);
  xor g_116020_(out[142], out[702], _057888_);
  xor g_116021_(out[136], out[696], _057889_);
  xor g_116022_(out[129], out[689], _057890_);
  xor g_116023_(out[141], out[701], _057891_);
  xor g_116024_(out[137], out[697], _057893_);
  xor g_116025_(out[132], out[692], _057894_);
  xor g_116026_(out[130], out[690], _057895_);
  and g_116027_(out[139], _049642_, _057896_);
  xor g_116028_(out[131], out[691], _057897_);
  xor g_116029_(out[134], out[694], _057898_);
  xor g_116030_(out[143], out[703], _057899_);
  xor g_116031_(out[138], out[698], _057900_);
  xor g_116032_(out[133], out[693], _057901_);
  xor g_116033_(out[128], out[688], _057902_);
  or g_116034_(_057888_, _057894_, _057904_);
  or g_116035_(_057889_, _057891_, _057905_);
  or g_116036_(_057895_, _057900_, _057906_);
  or g_116037_(_057905_, _057906_, _057907_);
  or g_116038_(_057893_, _057897_, _057908_);
  or g_116039_(_057901_, _057902_, _057909_);
  or g_116040_(_057908_, _057909_, _057910_);
  or g_116041_(_057907_, _057910_, _057911_);
  xor g_116042_(out[140], out[700], _057912_);
  or g_116043_(_057887_, _057912_, _057913_);
  or g_116044_(_057886_, _057898_, _057915_);
  or g_116045_(_057913_, _057915_, _057916_);
  or g_116046_(_057890_, _057896_, _057917_);
  or g_116047_(_057899_, _057917_, _057918_);
  or g_116048_(_057916_, _057918_, _057919_);
  or g_116049_(_057911_, _057919_, _057920_);
  or g_116050_(_057904_, _057920_, _057921_);
  xor g_116051_(out[113], out[689], _057922_);
  and g_116052_(out[123], _049642_, _057923_);
  xor g_116053_(out[121], out[697], _057924_);
  xor g_116054_(out[112], out[688], _057926_);
  xor g_116055_(out[126], out[702], _057927_);
  xor g_116056_(out[116], out[692], _057928_);
  or g_116057_(_057927_, _057928_, _057929_);
  xor g_116058_(out[125], out[701], _057930_);
  xor g_116059_(out[115], out[691], _057931_);
  and g_116060_(_098151_, out[699], _057932_);
  xor g_116061_(out[118], out[694], _057933_);
  xor g_116062_(out[122], out[698], _057934_);
  xor g_116063_(out[117], out[693], _057935_);
  xor g_116064_(out[127], out[703], _057937_);
  xor g_116065_(out[120], out[696], _057938_);
  or g_116066_(_057930_, _057938_, _057939_);
  xor g_116067_(out[114], out[690], _057940_);
  or g_116068_(_057934_, _057940_, _057941_);
  or g_116069_(_057939_, _057941_, _057942_);
  or g_116070_(_057924_, _057931_, _057943_);
  or g_116071_(_057935_, _057943_, _057944_);
  or g_116072_(_057942_, _057944_, _057945_);
  or g_116073_(_057929_, _057945_, _057946_);
  xor g_116074_(out[124], out[700], _057948_);
  or g_116075_(_057932_, _057948_, _057949_);
  xor g_116076_(out[119], out[695], _057950_);
  or g_116077_(_057933_, _057950_, _057951_);
  or g_116078_(_057949_, _057951_, _057952_);
  or g_116079_(_057922_, _057923_, _057953_);
  or g_116080_(_057937_, _057953_, _057954_);
  or g_116081_(_057952_, _057954_, _057955_);
  or g_116082_(_057926_, _057955_, _057956_);
  or g_116083_(_057946_, _057956_, _057957_);
  xor g_116084_(out[103], out[695], _057959_);
  and g_116085_(_098140_, out[699], _057960_);
  xor g_116086_(out[110], out[702], _057961_);
  xor g_116087_(out[104], out[696], _057962_);
  xor g_116088_(out[97], out[689], _057963_);
  xor g_116089_(out[109], out[701], _057964_);
  xor g_116090_(out[105], out[697], _057965_);
  xor g_116091_(out[100], out[692], _057966_);
  xor g_116092_(out[98], out[690], _057967_);
  and g_116093_(out[107], _049642_, _057968_);
  xor g_116094_(out[99], out[691], _057970_);
  xor g_116095_(out[102], out[694], _057971_);
  xor g_116096_(out[111], out[703], _057972_);
  xor g_116097_(out[106], out[698], _057973_);
  xor g_116098_(out[101], out[693], _057974_);
  xor g_116099_(out[96], out[688], _057975_);
  or g_116100_(_057961_, _057966_, _057976_);
  or g_116101_(_057962_, _057964_, _057977_);
  or g_116102_(_057967_, _057973_, _057978_);
  or g_116103_(_057977_, _057978_, _057979_);
  or g_116104_(_057965_, _057970_, _057981_);
  or g_116105_(_057974_, _057975_, _057982_);
  or g_116106_(_057981_, _057982_, _057983_);
  or g_116107_(_057979_, _057983_, _057984_);
  xor g_116108_(out[108], out[700], _057985_);
  or g_116109_(_057960_, _057985_, _057986_);
  or g_116110_(_057959_, _057971_, _057987_);
  or g_116111_(_057986_, _057987_, _057988_);
  or g_116112_(_057963_, _057968_, _057989_);
  or g_116113_(_057972_, _057989_, _057990_);
  or g_116114_(_057988_, _057990_, _057992_);
  or g_116115_(_057984_, _057992_, _057993_);
  or g_116116_(_057976_, _057993_, _057994_);
  and g_116117_(out[91], _049642_, _057995_);
  xor g_116118_(out[84], out[692], _057996_);
  xor g_116119_(out[94], out[702], _057997_);
  or g_116120_(_057996_, _057997_, _057998_);
  xor g_116121_(out[93], out[701], _057999_);
  xor g_116122_(out[83], out[691], _058000_);
  xor g_116123_(out[80], out[688], _058001_);
  and g_116124_(_098129_, out[699], _058003_);
  xor g_116125_(out[90], out[698], _058004_);
  xor g_116126_(out[95], out[703], _058005_);
  xor g_116127_(out[86], out[694], _058006_);
  xor g_116128_(out[85], out[693], _058007_);
  xor g_116129_(out[88], out[696], _058008_);
  or g_116130_(_057999_, _058008_, _058009_);
  xor g_116131_(out[82], out[690], _058010_);
  xor g_116132_(out[89], out[697], _058011_);
  xor g_116133_(out[81], out[689], _058012_);
  or g_116134_(_058004_, _058010_, _058014_);
  or g_116135_(_058009_, _058014_, _058015_);
  or g_116136_(_058000_, _058011_, _058016_);
  or g_116137_(_058007_, _058016_, _058017_);
  or g_116138_(_058015_, _058017_, _058018_);
  or g_116139_(_057998_, _058018_, _058019_);
  xor g_116140_(out[92], out[700], _058020_);
  or g_116141_(_058003_, _058020_, _058021_);
  xor g_116142_(out[87], out[695], _058022_);
  or g_116143_(_058006_, _058022_, _058023_);
  or g_116144_(_058021_, _058023_, _058025_);
  or g_116145_(_057995_, _058012_, _058026_);
  or g_116146_(_058005_, _058026_, _058027_);
  or g_116147_(_058025_, _058027_, _058028_);
  or g_116148_(_058001_, _058028_, _058029_);
  or g_116149_(_058019_, _058029_, _058030_);
  xor g_116150_(out[71], out[695], _058031_);
  and g_116151_(_098118_, out[699], _058032_);
  xor g_116152_(out[78], out[702], _058033_);
  xor g_116153_(out[72], out[696], _058034_);
  xor g_116154_(out[65], out[689], _058036_);
  xor g_116155_(out[77], out[701], _058037_);
  xor g_116156_(out[73], out[697], _058038_);
  xor g_116157_(out[68], out[692], _058039_);
  xor g_116158_(out[66], out[690], _058040_);
  and g_116159_(out[75], _049642_, _058041_);
  xor g_116160_(out[67], out[691], _058042_);
  xor g_116161_(out[70], out[694], _058043_);
  xor g_116162_(out[79], out[703], _058044_);
  xor g_116163_(out[74], out[698], _058045_);
  xor g_116164_(out[69], out[693], _058047_);
  xor g_116165_(out[64], out[688], _058048_);
  or g_116166_(_058033_, _058039_, _058049_);
  or g_116167_(_058034_, _058037_, _058050_);
  or g_116168_(_058040_, _058045_, _058051_);
  or g_116169_(_058050_, _058051_, _058052_);
  or g_116170_(_058038_, _058042_, _058053_);
  or g_116171_(_058047_, _058048_, _058054_);
  or g_116172_(_058053_, _058054_, _058055_);
  or g_116173_(_058052_, _058055_, _058056_);
  xor g_116174_(out[76], out[700], _058058_);
  or g_116175_(_058032_, _058058_, _058059_);
  or g_116176_(_058031_, _058043_, _058060_);
  or g_116177_(_058059_, _058060_, _058061_);
  or g_116178_(_058036_, _058041_, _058062_);
  or g_116179_(_058044_, _058062_, _058063_);
  or g_116180_(_058061_, _058063_, _058064_);
  or g_116181_(_058056_, _058064_, _058065_);
  or g_116182_(_058049_, _058065_, _058066_);
  not g_116183_(_058066_, _058067_);
  xor g_116184_(out[49], out[689], _058069_);
  and g_116185_(out[59], _049642_, _058070_);
  xor g_116186_(out[62], out[702], _058071_);
  xor g_116187_(out[51], out[691], _058072_);
  xor g_116188_(out[52], out[692], _058073_);
  xor g_116189_(out[50], out[690], _058074_);
  xor g_116190_(out[57], out[697], _058075_);
  xor g_116191_(out[48], out[688], _058076_);
  and g_116192_(_098107_, out[699], _058077_);
  xor g_116193_(out[54], out[694], _058078_);
  xor g_116194_(out[58], out[698], _058080_);
  xor g_116195_(out[53], out[693], _058081_);
  xor g_116196_(out[63], out[703], _058082_);
  xor g_116197_(out[61], out[701], _058083_);
  xor g_116198_(out[56], out[696], _058084_);
  or g_116199_(_058071_, _058073_, _058085_);
  or g_116200_(_058083_, _058084_, _058086_);
  or g_116201_(_058074_, _058080_, _058087_);
  or g_116202_(_058086_, _058087_, _058088_);
  or g_116203_(_058072_, _058075_, _058089_);
  or g_116204_(_058076_, _058081_, _058091_);
  or g_116205_(_058089_, _058091_, _058092_);
  or g_116206_(_058088_, _058092_, _058093_);
  xor g_116207_(out[60], out[700], _058094_);
  or g_116208_(_058077_, _058094_, _058095_);
  xor g_116209_(out[55], out[695], _058096_);
  or g_116210_(_058078_, _058096_, _058097_);
  or g_116211_(_058095_, _058097_, _058098_);
  or g_116212_(_058069_, _058070_, _058099_);
  or g_116213_(_058082_, _058099_, _058100_);
  or g_116214_(_058098_, _058100_, _058102_);
  or g_116215_(_058093_, _058102_, _058103_);
  or g_116216_(_058085_, _058103_, _058104_);
  xor g_116217_(out[39], out[695], _058105_);
  and g_116218_(_098096_, out[699], _058106_);
  xor g_116219_(out[46], out[702], _058107_);
  xor g_116220_(out[40], out[696], _058108_);
  xor g_116221_(out[33], out[689], _058109_);
  xor g_116222_(out[45], out[701], _058110_);
  xor g_116223_(out[41], out[697], _058111_);
  xor g_116224_(out[36], out[692], _058113_);
  xor g_116225_(out[34], out[690], _058114_);
  and g_116226_(out[43], _049642_, _058115_);
  xor g_116227_(out[35], out[691], _058116_);
  xor g_116228_(out[38], out[694], _058117_);
  xor g_116229_(out[47], out[703], _058118_);
  xor g_116230_(out[42], out[698], _058119_);
  xor g_116231_(out[37], out[693], _058120_);
  xor g_116232_(out[32], out[688], _058121_);
  or g_116233_(_058107_, _058113_, _058122_);
  or g_116234_(_058108_, _058110_, _058124_);
  or g_116235_(_058114_, _058119_, _058125_);
  or g_116236_(_058124_, _058125_, _058126_);
  or g_116237_(_058111_, _058116_, _058127_);
  or g_116238_(_058120_, _058121_, _058128_);
  or g_116239_(_058127_, _058128_, _058129_);
  or g_116240_(_058126_, _058129_, _058130_);
  xor g_116241_(out[44], out[700], _058131_);
  or g_116242_(_058106_, _058131_, _058132_);
  or g_116243_(_058105_, _058117_, _058133_);
  or g_116244_(_058132_, _058133_, _058135_);
  or g_116245_(_058109_, _058115_, _058136_);
  or g_116246_(_058118_, _058136_, _058137_);
  or g_116247_(_058135_, _058137_, _058138_);
  or g_116248_(_058130_, _058138_, _058139_);
  or g_116249_(_058122_, _058139_, _058140_);
  xor g_116250_(out[29], out[701], _058141_);
  xor g_116251_(out[18], out[690], _058142_);
  xor g_116252_(out[21], out[693], _058143_);
  xor g_116253_(out[25], out[697], _058144_);
  xor g_116254_(out[20], out[692], _058146_);
  xor g_116255_(out[24], out[696], _058147_);
  xor g_116256_(out[30], out[702], _058148_);
  xor g_116257_(out[22], out[694], _058149_);
  xor g_116258_(out[31], out[703], _058150_);
  xor g_116259_(out[26], out[698], _058151_);
  xor g_116260_(out[16], out[688], _058152_);
  xor g_116261_(out[19], out[691], _058153_);
  and g_116262_(_098063_, out[699], _058154_);
  and g_116263_(out[27], _049642_, _058155_);
  xor g_116264_(out[17], out[689], _058157_);
  or g_116265_(_058146_, _058148_, _058158_);
  or g_116266_(_058141_, _058147_, _058159_);
  or g_116267_(_058142_, _058151_, _058160_);
  or g_116268_(_058159_, _058160_, _058161_);
  or g_116269_(_058144_, _058153_, _058162_);
  or g_116270_(_058143_, _058152_, _058163_);
  or g_116271_(_058162_, _058163_, _058164_);
  or g_116272_(_058161_, _058164_, _058165_);
  xor g_116273_(out[28], out[700], _058166_);
  or g_116274_(_058154_, _058166_, _058168_);
  xor g_116275_(out[23], out[695], _058169_);
  or g_116276_(_058149_, _058169_, _058170_);
  or g_116277_(_058168_, _058170_, _058171_);
  or g_116278_(_058155_, _058157_, _058172_);
  or g_116279_(_058150_, _058172_, _058173_);
  or g_116280_(_058171_, _058173_, _058174_);
  or g_116281_(_058165_, _058174_, _058175_);
  or g_116282_(_058158_, _058175_, _058176_);
  not g_116283_(_058176_, _058177_);
  and g_116284_(out[11], _049642_, _058179_);
  xor g_116285_(out[4], out[692], _058180_);
  xor g_116286_(out[14], out[702], _058181_);
  or g_116287_(_058180_, _058181_, _058182_);
  xor g_116288_(out[13], out[701], _058183_);
  xor g_116289_(out[3], out[691], _058184_);
  xor g_116290_(out[0], out[688], _058185_);
  and g_116291_(_098041_, out[699], _058186_);
  xor g_116292_(out[10], out[698], _058187_);
  xor g_116293_(out[15], out[703], _058188_);
  xor g_116294_(out[6], out[694], _058190_);
  xor g_116295_(out[5], out[693], _058191_);
  xor g_116296_(out[8], out[696], _058192_);
  or g_116297_(_058183_, _058192_, _058193_);
  xor g_116298_(out[2], out[690], _058194_);
  xor g_116299_(out[9], out[697], _058195_);
  xor g_116300_(out[1], out[689], _058196_);
  or g_116301_(_058187_, _058194_, _058197_);
  or g_116302_(_058193_, _058197_, _058198_);
  or g_116303_(_058184_, _058195_, _058199_);
  or g_116304_(_058191_, _058199_, _058201_);
  or g_116305_(_058198_, _058201_, _058202_);
  or g_116306_(_058182_, _058202_, _058203_);
  xor g_116307_(out[12], out[700], _058204_);
  or g_116308_(_058186_, _058204_, _058205_);
  xor g_116309_(out[7], out[695], _058206_);
  or g_116310_(_058190_, _058206_, _058207_);
  or g_116311_(_058205_, _058207_, _058208_);
  or g_116312_(_058179_, _058196_, _058209_);
  or g_116313_(_058188_, _058209_, _058210_);
  or g_116314_(_058208_, _058210_, _058212_);
  or g_116315_(_058185_, _058212_, _058213_);
  or g_116316_(_058203_, _058213_, _058214_);
  xor g_116317_(out[471], out[679], _058215_);
  and g_116318_(_049499_, out[683], _058216_);
  xor g_116319_(out[478], out[686], _058217_);
  xor g_116320_(out[472], out[680], _058218_);
  xor g_116321_(out[465], out[673], _058219_);
  xor g_116322_(out[477], out[685], _058220_);
  xor g_116323_(out[473], out[681], _058221_);
  xor g_116324_(out[468], out[676], _058223_);
  xor g_116325_(out[466], out[674], _058224_);
  and g_116326_(out[475], _049631_, _058225_);
  xor g_116327_(out[467], out[675], _058226_);
  xor g_116328_(out[470], out[678], _058227_);
  xor g_116329_(out[479], out[687], _058228_);
  xor g_116330_(out[474], out[682], _058229_);
  xor g_116331_(out[469], out[677], _058230_);
  xor g_116332_(out[464], out[672], _058231_);
  or g_116333_(_058217_, _058223_, _058232_);
  or g_116334_(_058218_, _058220_, _058234_);
  or g_116335_(_058224_, _058229_, _058235_);
  or g_116336_(_058234_, _058235_, _058236_);
  or g_116337_(_058221_, _058226_, _058237_);
  or g_116338_(_058230_, _058231_, _058238_);
  or g_116339_(_058237_, _058238_, _058239_);
  or g_116340_(_058236_, _058239_, _058240_);
  xor g_116341_(out[476], out[684], _058241_);
  or g_116342_(_058216_, _058241_, _058242_);
  or g_116343_(_058215_, _058227_, _058243_);
  or g_116344_(_058242_, _058243_, _058245_);
  or g_116345_(_058219_, _058225_, _058246_);
  or g_116346_(_058228_, _058246_, _058247_);
  or g_116347_(_058245_, _058247_, _058248_);
  or g_116348_(_058240_, _058248_, _058249_);
  or g_116349_(_058232_, _058249_, _058250_);
  xor g_116350_(out[451], out[675], _058251_);
  xor g_116351_(out[452], out[676], _058252_);
  xor g_116352_(out[462], out[686], _058253_);
  xor g_116353_(out[450], out[674], _058254_);
  xor g_116354_(out[453], out[677], _058256_);
  xor g_116355_(out[457], out[681], _058257_);
  xor g_116356_(out[456], out[680], _058258_);
  xor g_116357_(out[463], out[687], _058259_);
  xor g_116358_(out[458], out[682], _058260_);
  xor g_116359_(out[454], out[678], _058261_);
  xor g_116360_(out[448], out[672], _058262_);
  and g_116361_(_049477_, out[683], _058263_);
  and g_116362_(out[459], _049631_, _058264_);
  xor g_116363_(out[461], out[685], _058265_);
  or g_116364_(_058258_, _058265_, _058267_);
  xor g_116365_(out[449], out[673], _058268_);
  or g_116366_(_058254_, _058260_, _058269_);
  or g_116367_(_058267_, _058269_, _058270_);
  or g_116368_(_058251_, _058257_, _058271_);
  or g_116369_(_058256_, _058271_, _058272_);
  or g_116370_(_058270_, _058272_, _058273_);
  or g_116371_(_058252_, _058253_, _058274_);
  or g_116372_(_058273_, _058274_, _058275_);
  xor g_116373_(out[460], out[684], _058276_);
  or g_116374_(_058263_, _058276_, _058278_);
  xor g_116375_(out[455], out[679], _058279_);
  or g_116376_(_058261_, _058279_, _058280_);
  or g_116377_(_058278_, _058280_, _058281_);
  or g_116378_(_058264_, _058268_, _058282_);
  or g_116379_(_058259_, _058282_, _058283_);
  or g_116380_(_058281_, _058283_, _058284_);
  or g_116381_(_058262_, _058284_, _058285_);
  or g_116382_(_058275_, _058285_, _058286_);
  not g_116383_(_058286_, _058287_);
  xor g_116384_(out[439], out[679], _058289_);
  and g_116385_(_049466_, out[683], _058290_);
  xor g_116386_(out[446], out[686], _058291_);
  xor g_116387_(out[440], out[680], _058292_);
  xor g_116388_(out[433], out[673], _058293_);
  xor g_116389_(out[445], out[685], _058294_);
  xor g_116390_(out[441], out[681], _058295_);
  xor g_116391_(out[436], out[676], _058296_);
  xor g_116392_(out[434], out[674], _058297_);
  and g_116393_(out[443], _049631_, _058298_);
  xor g_116394_(out[435], out[675], _058300_);
  xor g_116395_(out[438], out[678], _058301_);
  xor g_116396_(out[447], out[687], _058302_);
  xor g_116397_(out[442], out[682], _058303_);
  xor g_116398_(out[437], out[677], _058304_);
  xor g_116399_(out[432], out[672], _058305_);
  or g_116400_(_058291_, _058296_, _058306_);
  or g_116401_(_058292_, _058294_, _058307_);
  or g_116402_(_058297_, _058303_, _058308_);
  or g_116403_(_058307_, _058308_, _058309_);
  or g_116404_(_058295_, _058300_, _058311_);
  or g_116405_(_058304_, _058305_, _058312_);
  or g_116406_(_058311_, _058312_, _058313_);
  or g_116407_(_058309_, _058313_, _058314_);
  xor g_116408_(out[444], out[684], _058315_);
  or g_116409_(_058290_, _058315_, _058316_);
  or g_116410_(_058289_, _058301_, _058317_);
  or g_116411_(_058316_, _058317_, _058318_);
  or g_116412_(_058293_, _058298_, _058319_);
  or g_116413_(_058302_, _058319_, _058320_);
  or g_116414_(_058318_, _058320_, _058322_);
  or g_116415_(_058314_, _058322_, _058323_);
  or g_116416_(_058306_, _058323_, _058324_);
  xor g_116417_(out[417], out[673], _058325_);
  and g_116418_(out[427], _049631_, _058326_);
  xor g_116419_(out[425], out[681], _058327_);
  xor g_116420_(out[416], out[672], _058328_);
  xor g_116421_(out[430], out[686], _058329_);
  xor g_116422_(out[420], out[676], _058330_);
  or g_116423_(_058329_, _058330_, _058331_);
  xor g_116424_(out[429], out[685], _058333_);
  xor g_116425_(out[419], out[675], _058334_);
  and g_116426_(_049455_, out[683], _058335_);
  xor g_116427_(out[422], out[678], _058336_);
  xor g_116428_(out[426], out[682], _058337_);
  xor g_116429_(out[421], out[677], _058338_);
  xor g_116430_(out[431], out[687], _058339_);
  xor g_116431_(out[424], out[680], _058340_);
  or g_116432_(_058333_, _058340_, _058341_);
  xor g_116433_(out[418], out[674], _058342_);
  or g_116434_(_058337_, _058342_, _058344_);
  or g_116435_(_058341_, _058344_, _058345_);
  or g_116436_(_058327_, _058334_, _058346_);
  or g_116437_(_058338_, _058346_, _058347_);
  or g_116438_(_058345_, _058347_, _058348_);
  or g_116439_(_058331_, _058348_, _058349_);
  xor g_116440_(out[428], out[684], _058350_);
  or g_116441_(_058335_, _058350_, _058351_);
  xor g_116442_(out[423], out[679], _058352_);
  or g_116443_(_058336_, _058352_, _058353_);
  or g_116444_(_058351_, _058353_, _058355_);
  or g_116445_(_058325_, _058326_, _058356_);
  or g_116446_(_058339_, _058356_, _058357_);
  or g_116447_(_058355_, _058357_, _058358_);
  or g_116448_(_058328_, _058358_, _058359_);
  or g_116449_(_058349_, _058359_, _058360_);
  xor g_116450_(out[407], out[679], _058361_);
  and g_116451_(_049444_, out[683], _058362_);
  xor g_116452_(out[414], out[686], _058363_);
  xor g_116453_(out[408], out[680], _058364_);
  xor g_116454_(out[401], out[673], _058366_);
  xor g_116455_(out[413], out[685], _058367_);
  xor g_116456_(out[409], out[681], _058368_);
  xor g_116457_(out[404], out[676], _058369_);
  xor g_116458_(out[402], out[674], _058370_);
  and g_116459_(out[411], _049631_, _058371_);
  xor g_116460_(out[403], out[675], _058372_);
  xor g_116461_(out[406], out[678], _058373_);
  xor g_116462_(out[415], out[687], _058374_);
  xor g_116463_(out[410], out[682], _058375_);
  xor g_116464_(out[405], out[677], _058377_);
  xor g_116465_(out[400], out[672], _058378_);
  or g_116466_(_058363_, _058369_, _058379_);
  or g_116467_(_058364_, _058367_, _058380_);
  or g_116468_(_058370_, _058375_, _058381_);
  or g_116469_(_058380_, _058381_, _058382_);
  or g_116470_(_058368_, _058372_, _058383_);
  or g_116471_(_058377_, _058378_, _058384_);
  or g_116472_(_058383_, _058384_, _058385_);
  or g_116473_(_058382_, _058385_, _058386_);
  xor g_116474_(out[412], out[684], _058388_);
  or g_116475_(_058362_, _058388_, _058389_);
  or g_116476_(_058361_, _058373_, _058390_);
  or g_116477_(_058389_, _058390_, _058391_);
  or g_116478_(_058366_, _058371_, _058392_);
  or g_116479_(_058374_, _058392_, _058393_);
  or g_116480_(_058391_, _058393_, _058394_);
  or g_116481_(_058386_, _058394_, _058395_);
  or g_116482_(_058379_, _058395_, _058396_);
  and g_116483_(out[395], _049631_, _058397_);
  and g_116484_(_049433_, out[683], _058399_);
  xor g_116485_(out[392], out[680], _058400_);
  xor g_116486_(out[399], out[687], _058401_);
  xor g_116487_(out[385], out[673], _058402_);
  xor g_116488_(out[386], out[674], _058403_);
  xor g_116489_(out[388], out[676], _058404_);
  xor g_116490_(out[389], out[677], _058405_);
  xor g_116491_(out[393], out[681], _058406_);
  xor g_116492_(out[387], out[675], _058407_);
  xor g_116493_(out[398], out[686], _058408_);
  xor g_116494_(out[384], out[672], _058410_);
  xor g_116495_(out[394], out[682], _058411_);
  xor g_116496_(out[397], out[685], _058412_);
  or g_116497_(_058400_, _058412_, _058413_);
  xor g_116498_(out[390], out[678], _058414_);
  or g_116499_(_058403_, _058411_, _058415_);
  or g_116500_(_058413_, _058415_, _058416_);
  or g_116501_(_058406_, _058407_, _058417_);
  or g_116502_(_058405_, _058417_, _058418_);
  or g_116503_(_058416_, _058418_, _058419_);
  or g_116504_(_058404_, _058408_, _058421_);
  or g_116505_(_058419_, _058421_, _058422_);
  xor g_116506_(out[396], out[684], _058423_);
  or g_116507_(_058399_, _058423_, _058424_);
  xor g_116508_(out[391], out[679], _058425_);
  or g_116509_(_058414_, _058425_, _058426_);
  or g_116510_(_058424_, _058426_, _058427_);
  or g_116511_(_058397_, _058402_, _058428_);
  or g_116512_(_058401_, _058428_, _058429_);
  or g_116513_(_058427_, _058429_, _058430_);
  or g_116514_(_058410_, _058430_, _058432_);
  or g_116515_(_058422_, _058432_, _058433_);
  xor g_116516_(out[375], out[679], _058434_);
  and g_116517_(_049422_, out[683], _058435_);
  xor g_116518_(out[382], out[686], _058436_);
  xor g_116519_(out[376], out[680], _058437_);
  xor g_116520_(out[369], out[673], _058438_);
  xor g_116521_(out[381], out[685], _058439_);
  xor g_116522_(out[377], out[681], _058440_);
  xor g_116523_(out[372], out[676], _058441_);
  xor g_116524_(out[370], out[674], _058443_);
  and g_116525_(out[379], _049631_, _058444_);
  xor g_116526_(out[371], out[675], _058445_);
  xor g_116527_(out[374], out[678], _058446_);
  xor g_116528_(out[383], out[687], _058447_);
  xor g_116529_(out[378], out[682], _058448_);
  xor g_116530_(out[373], out[677], _058449_);
  xor g_116531_(out[368], out[672], _058450_);
  or g_116532_(_058436_, _058441_, _058451_);
  or g_116533_(_058437_, _058439_, _058452_);
  or g_116534_(_058443_, _058448_, _058454_);
  or g_116535_(_058452_, _058454_, _058455_);
  or g_116536_(_058440_, _058445_, _058456_);
  or g_116537_(_058449_, _058450_, _058457_);
  or g_116538_(_058456_, _058457_, _058458_);
  or g_116539_(_058455_, _058458_, _058459_);
  xor g_116540_(out[380], out[684], _058460_);
  or g_116541_(_058435_, _058460_, _058461_);
  or g_116542_(_058434_, _058446_, _058462_);
  or g_116543_(_058461_, _058462_, _058463_);
  or g_116544_(_058438_, _058444_, _058465_);
  or g_116545_(_058447_, _058465_, _058466_);
  or g_116546_(_058463_, _058466_, _058467_);
  or g_116547_(_058459_, _058467_, _058468_);
  or g_116548_(_058451_, _058468_, _058469_);
  xor g_116549_(out[353], out[673], _058470_);
  and g_116550_(out[363], _049631_, _058471_);
  xor g_116551_(out[361], out[681], _058472_);
  xor g_116552_(out[352], out[672], _058473_);
  xor g_116553_(out[366], out[686], _058474_);
  xor g_116554_(out[356], out[676], _058476_);
  or g_116555_(_058474_, _058476_, _058477_);
  xor g_116556_(out[365], out[685], _058478_);
  xor g_116557_(out[355], out[675], _058479_);
  and g_116558_(_049411_, out[683], _058480_);
  xor g_116559_(out[358], out[678], _058481_);
  xor g_116560_(out[362], out[682], _058482_);
  xor g_116561_(out[357], out[677], _058483_);
  xor g_116562_(out[367], out[687], _058484_);
  xor g_116563_(out[360], out[680], _058485_);
  or g_116564_(_058478_, _058485_, _058487_);
  xor g_116565_(out[354], out[674], _058488_);
  or g_116566_(_058482_, _058488_, _058489_);
  or g_116567_(_058487_, _058489_, _058490_);
  or g_116568_(_058472_, _058479_, _058491_);
  or g_116569_(_058483_, _058491_, _058492_);
  or g_116570_(_058490_, _058492_, _058493_);
  or g_116571_(_058477_, _058493_, _058494_);
  xor g_116572_(out[364], out[684], _058495_);
  or g_116573_(_058480_, _058495_, _058496_);
  xor g_116574_(out[359], out[679], _058498_);
  or g_116575_(_058481_, _058498_, _058499_);
  or g_116576_(_058496_, _058499_, _058500_);
  or g_116577_(_058470_, _058471_, _058501_);
  or g_116578_(_058484_, _058501_, _058502_);
  or g_116579_(_058500_, _058502_, _058503_);
  or g_116580_(_058473_, _058503_, _058504_);
  or g_116581_(_058494_, _058504_, _058505_);
  xor g_116582_(out[343], out[679], _058506_);
  and g_116583_(_049400_, out[683], _058507_);
  xor g_116584_(out[350], out[686], _058509_);
  xor g_116585_(out[344], out[680], _058510_);
  xor g_116586_(out[337], out[673], _058511_);
  xor g_116587_(out[349], out[685], _058512_);
  xor g_116588_(out[345], out[681], _058513_);
  xor g_116589_(out[340], out[676], _058514_);
  xor g_116590_(out[338], out[674], _058515_);
  and g_116591_(out[347], _049631_, _058516_);
  xor g_116592_(out[339], out[675], _058517_);
  xor g_116593_(out[342], out[678], _058518_);
  xor g_116594_(out[351], out[687], _058520_);
  xor g_116595_(out[346], out[682], _058521_);
  xor g_116596_(out[341], out[677], _058522_);
  xor g_116597_(out[336], out[672], _058523_);
  or g_116598_(_058509_, _058514_, _058524_);
  or g_116599_(_058510_, _058512_, _058525_);
  or g_116600_(_058515_, _058521_, _058526_);
  or g_116601_(_058525_, _058526_, _058527_);
  or g_116602_(_058513_, _058517_, _058528_);
  or g_116603_(_058522_, _058523_, _058529_);
  or g_116604_(_058528_, _058529_, _058531_);
  or g_116605_(_058527_, _058531_, _058532_);
  xor g_116606_(out[348], out[684], _058533_);
  or g_116607_(_058507_, _058533_, _058534_);
  or g_116608_(_058506_, _058518_, _058535_);
  or g_116609_(_058534_, _058535_, _058536_);
  or g_116610_(_058511_, _058516_, _058537_);
  or g_116611_(_058520_, _058537_, _058538_);
  or g_116612_(_058536_, _058538_, _058539_);
  or g_116613_(_058532_, _058539_, _058540_);
  or g_116614_(_058524_, _058540_, _058542_);
  not g_116615_(_058542_, _058543_);
  xor g_116616_(out[321], out[673], _058544_);
  and g_116617_(out[331], _049631_, _058545_);
  xor g_116618_(out[329], out[681], _058546_);
  xor g_116619_(out[320], out[672], _058547_);
  xor g_116620_(out[334], out[686], _058548_);
  xor g_116621_(out[324], out[676], _058549_);
  or g_116622_(_058548_, _058549_, _058550_);
  xor g_116623_(out[333], out[685], _058551_);
  xor g_116624_(out[323], out[675], _058553_);
  and g_116625_(_098294_, out[683], _058554_);
  xor g_116626_(out[326], out[678], _058555_);
  xor g_116627_(out[330], out[682], _058556_);
  xor g_116628_(out[325], out[677], _058557_);
  xor g_116629_(out[335], out[687], _058558_);
  xor g_116630_(out[328], out[680], _058559_);
  or g_116631_(_058551_, _058559_, _058560_);
  xor g_116632_(out[322], out[674], _058561_);
  or g_116633_(_058556_, _058561_, _058562_);
  or g_116634_(_058560_, _058562_, _058564_);
  or g_116635_(_058546_, _058553_, _058565_);
  or g_116636_(_058557_, _058565_, _058566_);
  or g_116637_(_058564_, _058566_, _058567_);
  or g_116638_(_058550_, _058567_, _058568_);
  xor g_116639_(out[332], out[684], _058569_);
  or g_116640_(_058554_, _058569_, _058570_);
  xor g_116641_(out[327], out[679], _058571_);
  or g_116642_(_058555_, _058571_, _058572_);
  or g_116643_(_058570_, _058572_, _058573_);
  or g_116644_(_058544_, _058545_, _058575_);
  or g_116645_(_058558_, _058575_, _058576_);
  or g_116646_(_058573_, _058576_, _058577_);
  or g_116647_(_058547_, _058577_, _058578_);
  or g_116648_(_058568_, _058578_, _058579_);
  xor g_116649_(out[311], out[679], _058580_);
  and g_116650_(_098283_, out[683], _058581_);
  xor g_116651_(out[318], out[686], _058582_);
  xor g_116652_(out[312], out[680], _058583_);
  xor g_116653_(out[305], out[673], _058584_);
  xor g_116654_(out[317], out[685], _058586_);
  xor g_116655_(out[313], out[681], _058587_);
  xor g_116656_(out[308], out[676], _058588_);
  xor g_116657_(out[306], out[674], _058589_);
  and g_116658_(out[315], _049631_, _058590_);
  xor g_116659_(out[307], out[675], _058591_);
  xor g_116660_(out[310], out[678], _058592_);
  xor g_116661_(out[319], out[687], _058593_);
  xor g_116662_(out[314], out[682], _058594_);
  xor g_116663_(out[309], out[677], _058595_);
  xor g_116664_(out[304], out[672], _058597_);
  or g_116665_(_058582_, _058588_, _058598_);
  or g_116666_(_058583_, _058586_, _058599_);
  or g_116667_(_058589_, _058594_, _058600_);
  or g_116668_(_058599_, _058600_, _058601_);
  or g_116669_(_058587_, _058591_, _058602_);
  or g_116670_(_058595_, _058597_, _058603_);
  or g_116671_(_058602_, _058603_, _058604_);
  or g_116672_(_058601_, _058604_, _058605_);
  xor g_116673_(out[316], out[684], _058606_);
  or g_116674_(_058581_, _058606_, _058608_);
  or g_116675_(_058580_, _058592_, _058609_);
  or g_116676_(_058608_, _058609_, _058610_);
  or g_116677_(_058584_, _058590_, _058611_);
  or g_116678_(_058593_, _058611_, _058612_);
  or g_116679_(_058610_, _058612_, _058613_);
  or g_116680_(_058605_, _058613_, _058614_);
  or g_116681_(_058598_, _058614_, _058615_);
  xor g_116682_(out[300], out[684], _058616_);
  and g_116683_(_098272_, out[683], _058617_);
  xor g_116684_(out[301], out[685], _058619_);
  xor g_116685_(out[294], out[678], _058620_);
  xor g_116686_(out[296], out[680], _058621_);
  xor g_116687_(out[297], out[681], _058622_);
  xor g_116688_(out[302], out[686], _058623_);
  xor g_116689_(out[292], out[676], _058624_);
  or g_116690_(_058623_, _058624_, _058625_);
  xor g_116691_(out[293], out[677], _058626_);
  xor g_116692_(out[289], out[673], _058627_);
  and g_116693_(out[299], _049631_, _058628_);
  xor g_116694_(out[303], out[687], _058630_);
  xor g_116695_(out[298], out[682], _058631_);
  xor g_116696_(out[288], out[672], _058632_);
  xor g_116697_(out[290], out[674], _058633_);
  xor g_116698_(out[291], out[675], _058634_);
  or g_116699_(_058619_, _058621_, _058635_);
  or g_116700_(_058631_, _058633_, _058636_);
  or g_116701_(_058635_, _058636_, _058637_);
  or g_116702_(_058622_, _058634_, _058638_);
  or g_116703_(_058626_, _058632_, _058639_);
  or g_116704_(_058638_, _058639_, _058641_);
  or g_116705_(_058637_, _058641_, _058642_);
  or g_116706_(_058616_, _058617_, _058643_);
  xor g_116707_(out[295], out[679], _058644_);
  or g_116708_(_058620_, _058644_, _058645_);
  or g_116709_(_058643_, _058645_, _058646_);
  or g_116710_(_058627_, _058628_, _058647_);
  or g_116711_(_058630_, _058647_, _058648_);
  or g_116712_(_058646_, _058648_, _058649_);
  or g_116713_(_058642_, _058649_, _058650_);
  or g_116714_(_058625_, _058650_, _058652_);
  not g_116715_(_058652_, _058653_);
  xor g_116716_(out[279], out[679], _058654_);
  and g_116717_(_098261_, out[683], _058655_);
  xor g_116718_(out[286], out[686], _058656_);
  xor g_116719_(out[280], out[680], _058657_);
  xor g_116720_(out[273], out[673], _058658_);
  xor g_116721_(out[285], out[685], _058659_);
  xor g_116722_(out[281], out[681], _058660_);
  xor g_116723_(out[276], out[676], _058661_);
  xor g_116724_(out[274], out[674], _058663_);
  and g_116725_(out[283], _049631_, _058664_);
  xor g_116726_(out[275], out[675], _058665_);
  xor g_116727_(out[278], out[678], _058666_);
  xor g_116728_(out[287], out[687], _058667_);
  xor g_116729_(out[282], out[682], _058668_);
  xor g_116730_(out[277], out[677], _058669_);
  xor g_116731_(out[272], out[672], _058670_);
  or g_116732_(_058656_, _058661_, _058671_);
  or g_116733_(_058657_, _058659_, _058672_);
  or g_116734_(_058663_, _058668_, _058674_);
  or g_116735_(_058672_, _058674_, _058675_);
  or g_116736_(_058660_, _058665_, _058676_);
  or g_116737_(_058669_, _058670_, _058677_);
  or g_116738_(_058676_, _058677_, _058678_);
  or g_116739_(_058675_, _058678_, _058679_);
  xor g_116740_(out[284], out[684], _058680_);
  or g_116741_(_058655_, _058680_, _058681_);
  or g_116742_(_058654_, _058666_, _058682_);
  or g_116743_(_058681_, _058682_, _058683_);
  or g_116744_(_058658_, _058664_, _058685_);
  or g_116745_(_058667_, _058685_, _058686_);
  or g_116746_(_058683_, _058686_, _058687_);
  or g_116747_(_058679_, _058687_, _058688_);
  or g_116748_(_058671_, _058688_, _058689_);
  xor g_116749_(out[268], out[684], _058690_);
  and g_116750_(_098250_, out[683], _058691_);
  xor g_116751_(out[269], out[685], _058692_);
  xor g_116752_(out[262], out[678], _058693_);
  xor g_116753_(out[264], out[680], _058694_);
  xor g_116754_(out[265], out[681], _058696_);
  xor g_116755_(out[270], out[686], _058697_);
  xor g_116756_(out[260], out[676], _058698_);
  or g_116757_(_058697_, _058698_, _058699_);
  xor g_116758_(out[261], out[677], _058700_);
  xor g_116759_(out[257], out[673], _058701_);
  and g_116760_(out[267], _049631_, _058702_);
  xor g_116761_(out[271], out[687], _058703_);
  xor g_116762_(out[266], out[682], _058704_);
  xor g_116763_(out[256], out[672], _058705_);
  xor g_116764_(out[258], out[674], _058707_);
  xor g_116765_(out[259], out[675], _058708_);
  or g_116766_(_058692_, _058694_, _058709_);
  or g_116767_(_058704_, _058707_, _058710_);
  or g_116768_(_058709_, _058710_, _058711_);
  or g_116769_(_058696_, _058708_, _058712_);
  or g_116770_(_058700_, _058705_, _058713_);
  or g_116771_(_058712_, _058713_, _058714_);
  or g_116772_(_058711_, _058714_, _058715_);
  or g_116773_(_058690_, _058691_, _058716_);
  xor g_116774_(out[263], out[679], _058718_);
  or g_116775_(_058693_, _058718_, _058719_);
  or g_116776_(_058716_, _058719_, _058720_);
  or g_116777_(_058701_, _058702_, _058721_);
  or g_116778_(_058703_, _058721_, _058722_);
  or g_116779_(_058720_, _058722_, _058723_);
  or g_116780_(_058715_, _058723_, _058724_);
  or g_116781_(_058699_, _058724_, _058725_);
  xor g_116782_(out[247], out[679], _058726_);
  and g_116783_(_098239_, out[683], _058727_);
  xor g_116784_(out[254], out[686], _058729_);
  xor g_116785_(out[248], out[680], _058730_);
  xor g_116786_(out[241], out[673], _058731_);
  xor g_116787_(out[253], out[685], _058732_);
  xor g_116788_(out[249], out[681], _058733_);
  xor g_116789_(out[244], out[676], _058734_);
  xor g_116790_(out[242], out[674], _058735_);
  and g_116791_(out[251], _049631_, _058736_);
  xor g_116792_(out[243], out[675], _058737_);
  xor g_116793_(out[246], out[678], _058738_);
  xor g_116794_(out[255], out[687], _058740_);
  xor g_116795_(out[250], out[682], _058741_);
  xor g_116796_(out[245], out[677], _058742_);
  xor g_116797_(out[240], out[672], _058743_);
  or g_116798_(_058729_, _058734_, _058744_);
  or g_116799_(_058730_, _058732_, _058745_);
  or g_116800_(_058735_, _058741_, _058746_);
  or g_116801_(_058745_, _058746_, _058747_);
  or g_116802_(_058733_, _058737_, _058748_);
  or g_116803_(_058742_, _058743_, _058749_);
  or g_116804_(_058748_, _058749_, _058751_);
  or g_116805_(_058747_, _058751_, _058752_);
  xor g_116806_(out[252], out[684], _058753_);
  or g_116807_(_058727_, _058753_, _058754_);
  or g_116808_(_058726_, _058738_, _058755_);
  or g_116809_(_058754_, _058755_, _058756_);
  or g_116810_(_058731_, _058736_, _058757_);
  or g_116811_(_058740_, _058757_, _058758_);
  or g_116812_(_058756_, _058758_, _058759_);
  or g_116813_(_058752_, _058759_, _058760_);
  or g_116814_(_058744_, _058760_, _058762_);
  xor g_116815_(out[227], out[675], _058763_);
  xor g_116816_(out[228], out[676], _058764_);
  xor g_116817_(out[238], out[686], _058765_);
  xor g_116818_(out[226], out[674], _058766_);
  xor g_116819_(out[229], out[677], _058767_);
  xor g_116820_(out[233], out[681], _058768_);
  xor g_116821_(out[232], out[680], _058769_);
  xor g_116822_(out[239], out[687], _058770_);
  xor g_116823_(out[234], out[682], _058771_);
  xor g_116824_(out[230], out[678], _058773_);
  xor g_116825_(out[224], out[672], _058774_);
  and g_116826_(_098228_, out[683], _058775_);
  and g_116827_(out[235], _049631_, _058776_);
  xor g_116828_(out[237], out[685], _058777_);
  or g_116829_(_058769_, _058777_, _058778_);
  xor g_116830_(out[225], out[673], _058779_);
  or g_116831_(_058766_, _058771_, _058780_);
  or g_116832_(_058778_, _058780_, _058781_);
  or g_116833_(_058763_, _058768_, _058782_);
  or g_116834_(_058767_, _058782_, _058784_);
  or g_116835_(_058781_, _058784_, _058785_);
  or g_116836_(_058764_, _058765_, _058786_);
  or g_116837_(_058785_, _058786_, _058787_);
  xor g_116838_(out[236], out[684], _058788_);
  or g_116839_(_058775_, _058788_, _058789_);
  xor g_116840_(out[231], out[679], _058790_);
  or g_116841_(_058773_, _058790_, _058791_);
  or g_116842_(_058789_, _058791_, _058792_);
  or g_116843_(_058776_, _058779_, _058793_);
  or g_116844_(_058770_, _058793_, _058795_);
  or g_116845_(_058792_, _058795_, _058796_);
  or g_116846_(_058774_, _058796_, _058797_);
  or g_116847_(_058787_, _058797_, _058798_);
  xor g_116848_(out[215], out[679], _058799_);
  and g_116849_(_098217_, out[683], _058800_);
  xor g_116850_(out[222], out[686], _058801_);
  xor g_116851_(out[216], out[680], _058802_);
  xor g_116852_(out[209], out[673], _058803_);
  xor g_116853_(out[221], out[685], _058804_);
  xor g_116854_(out[217], out[681], _058806_);
  xor g_116855_(out[212], out[676], _058807_);
  xor g_116856_(out[210], out[674], _058808_);
  and g_116857_(out[219], _049631_, _058809_);
  xor g_116858_(out[211], out[675], _058810_);
  xor g_116859_(out[214], out[678], _058811_);
  xor g_116860_(out[223], out[687], _058812_);
  xor g_116861_(out[218], out[682], _058813_);
  xor g_116862_(out[213], out[677], _058814_);
  xor g_116863_(out[208], out[672], _058815_);
  or g_116864_(_058801_, _058807_, _058817_);
  or g_116865_(_058802_, _058804_, _058818_);
  or g_116866_(_058808_, _058813_, _058819_);
  or g_116867_(_058818_, _058819_, _058820_);
  or g_116868_(_058806_, _058810_, _058821_);
  or g_116869_(_058814_, _058815_, _058822_);
  or g_116870_(_058821_, _058822_, _058823_);
  or g_116871_(_058820_, _058823_, _058824_);
  xor g_116872_(out[220], out[684], _058825_);
  or g_116873_(_058800_, _058825_, _058826_);
  or g_116874_(_058799_, _058811_, _058828_);
  or g_116875_(_058826_, _058828_, _058829_);
  or g_116876_(_058803_, _058809_, _058830_);
  or g_116877_(_058812_, _058830_, _058831_);
  or g_116878_(_058829_, _058831_, _058832_);
  or g_116879_(_058824_, _058832_, _058833_);
  or g_116880_(_058817_, _058833_, _058834_);
  not g_116881_(_058834_, _058835_);
  xor g_116882_(out[193], out[673], _058836_);
  and g_116883_(out[203], _049631_, _058837_);
  xor g_116884_(out[201], out[681], _058839_);
  xor g_116885_(out[192], out[672], _058840_);
  xor g_116886_(out[206], out[686], _058841_);
  xor g_116887_(out[196], out[676], _058842_);
  or g_116888_(_058841_, _058842_, _058843_);
  xor g_116889_(out[205], out[685], _058844_);
  xor g_116890_(out[195], out[675], _058845_);
  and g_116891_(_098206_, out[683], _058846_);
  xor g_116892_(out[198], out[678], _058847_);
  xor g_116893_(out[202], out[682], _058848_);
  xor g_116894_(out[197], out[677], _058850_);
  xor g_116895_(out[207], out[687], _058851_);
  xor g_116896_(out[200], out[680], _058852_);
  or g_116897_(_058844_, _058852_, _058853_);
  xor g_116898_(out[194], out[674], _058854_);
  or g_116899_(_058848_, _058854_, _058855_);
  or g_116900_(_058853_, _058855_, _058856_);
  or g_116901_(_058839_, _058845_, _058857_);
  or g_116902_(_058850_, _058857_, _058858_);
  or g_116903_(_058856_, _058858_, _058859_);
  or g_116904_(_058843_, _058859_, _058861_);
  xor g_116905_(out[204], out[684], _058862_);
  or g_116906_(_058846_, _058862_, _058863_);
  xor g_116907_(out[199], out[679], _058864_);
  or g_116908_(_058847_, _058864_, _058865_);
  or g_116909_(_058863_, _058865_, _058866_);
  or g_116910_(_058836_, _058837_, _058867_);
  or g_116911_(_058851_, _058867_, _058868_);
  or g_116912_(_058866_, _058868_, _058869_);
  or g_116913_(_058840_, _058869_, _058870_);
  or g_116914_(_058861_, _058870_, _058872_);
  not g_116915_(_058872_, _058873_);
  xor g_116916_(out[183], out[679], _058874_);
  and g_116917_(_098195_, out[683], _058875_);
  xor g_116918_(out[190], out[686], _058876_);
  xor g_116919_(out[184], out[680], _058877_);
  xor g_116920_(out[177], out[673], _058878_);
  xor g_116921_(out[189], out[685], _058879_);
  xor g_116922_(out[185], out[681], _058880_);
  xor g_116923_(out[180], out[676], _058881_);
  xor g_116924_(out[178], out[674], _058883_);
  and g_116925_(out[187], _049631_, _058884_);
  xor g_116926_(out[179], out[675], _058885_);
  xor g_116927_(out[182], out[678], _058886_);
  xor g_116928_(out[191], out[687], _058887_);
  xor g_116929_(out[186], out[682], _058888_);
  xor g_116930_(out[181], out[677], _058889_);
  xor g_116931_(out[176], out[672], _058890_);
  or g_116932_(_058876_, _058881_, _058891_);
  or g_116933_(_058877_, _058879_, _058892_);
  or g_116934_(_058883_, _058888_, _058894_);
  or g_116935_(_058892_, _058894_, _058895_);
  or g_116936_(_058880_, _058885_, _058896_);
  or g_116937_(_058889_, _058890_, _058897_);
  or g_116938_(_058896_, _058897_, _058898_);
  or g_116939_(_058895_, _058898_, _058899_);
  xor g_116940_(out[188], out[684], _058900_);
  or g_116941_(_058875_, _058900_, _058901_);
  or g_116942_(_058874_, _058886_, _058902_);
  or g_116943_(_058901_, _058902_, _058903_);
  or g_116944_(_058878_, _058884_, _058905_);
  or g_116945_(_058887_, _058905_, _058906_);
  or g_116946_(_058903_, _058906_, _058907_);
  or g_116947_(_058899_, _058907_, _058908_);
  or g_116948_(_058891_, _058908_, _058909_);
  not g_116949_(_058909_, _058910_);
  xor g_116950_(out[168], out[680], _058911_);
  xor g_116951_(out[165], out[677], _058912_);
  xor g_116952_(out[163], out[675], _058913_);
  xor g_116953_(out[174], out[686], _058914_);
  xor g_116954_(out[173], out[685], _058916_);
  xor g_116955_(out[162], out[674], _058917_);
  xor g_116956_(out[169], out[681], _058918_);
  xor g_116957_(out[166], out[678], _058919_);
  xor g_116958_(out[175], out[687], _058920_);
  xor g_116959_(out[170], out[682], _058921_);
  xor g_116960_(out[164], out[676], _058922_);
  xor g_116961_(out[160], out[672], _058923_);
  and g_116962_(_098184_, out[683], _058924_);
  and g_116963_(out[171], _049631_, _058925_);
  or g_116964_(_058911_, _058916_, _058927_);
  xor g_116965_(out[161], out[673], _058928_);
  or g_116966_(_058917_, _058921_, _058929_);
  or g_116967_(_058927_, _058929_, _058930_);
  or g_116968_(_058913_, _058918_, _058931_);
  or g_116969_(_058912_, _058931_, _058932_);
  or g_116970_(_058930_, _058932_, _058933_);
  or g_116971_(_058914_, _058922_, _058934_);
  or g_116972_(_058933_, _058934_, _058935_);
  xor g_116973_(out[172], out[684], _058936_);
  or g_116974_(_058924_, _058936_, _058938_);
  xor g_116975_(out[167], out[679], _058939_);
  or g_116976_(_058919_, _058939_, _058940_);
  or g_116977_(_058938_, _058940_, _058941_);
  or g_116978_(_058925_, _058928_, _058942_);
  or g_116979_(_058920_, _058942_, _058943_);
  or g_116980_(_058941_, _058943_, _058944_);
  or g_116981_(_058923_, _058944_, _058945_);
  or g_116982_(_058935_, _058945_, _058946_);
  xor g_116983_(out[151], out[679], _058947_);
  and g_116984_(_098173_, out[683], _058949_);
  xor g_116985_(out[158], out[686], _058950_);
  xor g_116986_(out[152], out[680], _058951_);
  xor g_116987_(out[145], out[673], _058952_);
  xor g_116988_(out[157], out[685], _058953_);
  xor g_116989_(out[153], out[681], _058954_);
  xor g_116990_(out[148], out[676], _058955_);
  xor g_116991_(out[146], out[674], _058956_);
  and g_116992_(out[155], _049631_, _058957_);
  xor g_116993_(out[147], out[675], _058958_);
  xor g_116994_(out[150], out[678], _058960_);
  xor g_116995_(out[159], out[687], _058961_);
  xor g_116996_(out[154], out[682], _058962_);
  xor g_116997_(out[149], out[677], _058963_);
  xor g_116998_(out[144], out[672], _058964_);
  or g_116999_(_058950_, _058955_, _058965_);
  or g_117000_(_058951_, _058953_, _058966_);
  or g_117001_(_058956_, _058962_, _058967_);
  or g_117002_(_058966_, _058967_, _058968_);
  or g_117003_(_058954_, _058958_, _058969_);
  or g_117004_(_058963_, _058964_, _058971_);
  or g_117005_(_058969_, _058971_, _058972_);
  or g_117006_(_058968_, _058972_, _058973_);
  xor g_117007_(out[156], out[684], _058974_);
  or g_117008_(_058949_, _058974_, _058975_);
  or g_117009_(_058947_, _058960_, _058976_);
  or g_117010_(_058975_, _058976_, _058977_);
  or g_117011_(_058952_, _058957_, _058978_);
  or g_117012_(_058961_, _058978_, _058979_);
  or g_117013_(_058977_, _058979_, _058980_);
  or g_117014_(_058973_, _058980_, _058982_);
  or g_117015_(_058965_, _058982_, _058983_);
  not g_117016_(_058983_, _058984_);
  xor g_117017_(out[129], out[673], _058985_);
  and g_117018_(out[139], _049631_, _058986_);
  xor g_117019_(out[137], out[681], _058987_);
  xor g_117020_(out[128], out[672], _058988_);
  xor g_117021_(out[142], out[686], _058989_);
  xor g_117022_(out[132], out[676], _058990_);
  or g_117023_(_058989_, _058990_, _058991_);
  xor g_117024_(out[141], out[685], _058993_);
  xor g_117025_(out[131], out[675], _058994_);
  and g_117026_(_098162_, out[683], _058995_);
  xor g_117027_(out[134], out[678], _058996_);
  xor g_117028_(out[138], out[682], _058997_);
  xor g_117029_(out[133], out[677], _058998_);
  xor g_117030_(out[143], out[687], _058999_);
  xor g_117031_(out[136], out[680], _059000_);
  or g_117032_(_058993_, _059000_, _059001_);
  xor g_117033_(out[130], out[674], _059002_);
  or g_117034_(_058997_, _059002_, _059004_);
  or g_117035_(_059001_, _059004_, _059005_);
  or g_117036_(_058987_, _058994_, _059006_);
  or g_117037_(_058998_, _059006_, _059007_);
  or g_117038_(_059005_, _059007_, _059008_);
  or g_117039_(_058991_, _059008_, _059009_);
  xor g_117040_(out[140], out[684], _059010_);
  or g_117041_(_058995_, _059010_, _059011_);
  xor g_117042_(out[135], out[679], _059012_);
  or g_117043_(_058996_, _059012_, _059013_);
  or g_117044_(_059011_, _059013_, _059015_);
  or g_117045_(_058985_, _058986_, _059016_);
  or g_117046_(_058999_, _059016_, _059017_);
  or g_117047_(_059015_, _059017_, _059018_);
  or g_117048_(_058988_, _059018_, _059019_);
  or g_117049_(_059009_, _059019_, _059020_);
  xor g_117050_(out[119], out[679], _059021_);
  and g_117051_(_098151_, out[683], _059022_);
  xor g_117052_(out[126], out[686], _059023_);
  xor g_117053_(out[120], out[680], _059024_);
  xor g_117054_(out[113], out[673], _059026_);
  xor g_117055_(out[125], out[685], _059027_);
  xor g_117056_(out[121], out[681], _059028_);
  xor g_117057_(out[116], out[676], _059029_);
  xor g_117058_(out[114], out[674], _059030_);
  and g_117059_(out[123], _049631_, _059031_);
  xor g_117060_(out[115], out[675], _059032_);
  xor g_117061_(out[118], out[678], _059033_);
  xor g_117062_(out[127], out[687], _059034_);
  xor g_117063_(out[122], out[682], _059035_);
  xor g_117064_(out[117], out[677], _059037_);
  xor g_117065_(out[112], out[672], _059038_);
  or g_117066_(_059023_, _059029_, _059039_);
  or g_117067_(_059024_, _059027_, _059040_);
  or g_117068_(_059030_, _059035_, _059041_);
  or g_117069_(_059040_, _059041_, _059042_);
  or g_117070_(_059028_, _059032_, _059043_);
  or g_117071_(_059037_, _059038_, _059044_);
  or g_117072_(_059043_, _059044_, _059045_);
  or g_117073_(_059042_, _059045_, _059046_);
  xor g_117074_(out[124], out[684], _059048_);
  or g_117075_(_059022_, _059048_, _059049_);
  or g_117076_(_059021_, _059033_, _059050_);
  or g_117077_(_059049_, _059050_, _059051_);
  or g_117078_(_059026_, _059031_, _059052_);
  or g_117079_(_059034_, _059052_, _059053_);
  or g_117080_(_059051_, _059053_, _059054_);
  or g_117081_(_059046_, _059054_, _059055_);
  or g_117082_(_059039_, _059055_, _059056_);
  xor g_117083_(out[97], out[673], _059057_);
  and g_117084_(out[107], _049631_, _059059_);
  xor g_117085_(out[105], out[681], _059060_);
  xor g_117086_(out[96], out[672], _059061_);
  xor g_117087_(out[110], out[686], _059062_);
  xor g_117088_(out[100], out[676], _059063_);
  or g_117089_(_059062_, _059063_, _059064_);
  xor g_117090_(out[109], out[685], _059065_);
  xor g_117091_(out[99], out[675], _059066_);
  and g_117092_(_098140_, out[683], _059067_);
  xor g_117093_(out[102], out[678], _059068_);
  xor g_117094_(out[106], out[682], _059070_);
  xor g_117095_(out[101], out[677], _059071_);
  xor g_117096_(out[111], out[687], _059072_);
  xor g_117097_(out[104], out[680], _059073_);
  or g_117098_(_059065_, _059073_, _059074_);
  xor g_117099_(out[98], out[674], _059075_);
  or g_117100_(_059070_, _059075_, _059076_);
  or g_117101_(_059074_, _059076_, _059077_);
  or g_117102_(_059060_, _059066_, _059078_);
  or g_117103_(_059071_, _059078_, _059079_);
  or g_117104_(_059077_, _059079_, _059081_);
  or g_117105_(_059064_, _059081_, _059082_);
  xor g_117106_(out[108], out[684], _059083_);
  or g_117107_(_059067_, _059083_, _059084_);
  xor g_117108_(out[103], out[679], _059085_);
  or g_117109_(_059068_, _059085_, _059086_);
  or g_117110_(_059084_, _059086_, _059087_);
  or g_117111_(_059057_, _059059_, _059088_);
  or g_117112_(_059072_, _059088_, _059089_);
  or g_117113_(_059087_, _059089_, _059090_);
  or g_117114_(_059061_, _059090_, _059092_);
  or g_117115_(_059082_, _059092_, _059093_);
  xor g_117116_(out[87], out[679], _059094_);
  and g_117117_(_098129_, out[683], _059095_);
  xor g_117118_(out[94], out[686], _059096_);
  xor g_117119_(out[88], out[680], _059097_);
  xor g_117120_(out[81], out[673], _059098_);
  xor g_117121_(out[93], out[685], _059099_);
  xor g_117122_(out[89], out[681], _059100_);
  xor g_117123_(out[84], out[676], _059101_);
  xor g_117124_(out[82], out[674], _059103_);
  and g_117125_(out[91], _049631_, _059104_);
  xor g_117126_(out[83], out[675], _059105_);
  xor g_117127_(out[86], out[678], _059106_);
  xor g_117128_(out[95], out[687], _059107_);
  xor g_117129_(out[90], out[682], _059108_);
  xor g_117130_(out[85], out[677], _059109_);
  xor g_117131_(out[80], out[672], _059110_);
  or g_117132_(_059096_, _059101_, _059111_);
  or g_117133_(_059097_, _059099_, _059112_);
  or g_117134_(_059103_, _059108_, _059114_);
  or g_117135_(_059112_, _059114_, _059115_);
  or g_117136_(_059100_, _059105_, _059116_);
  or g_117137_(_059109_, _059110_, _059117_);
  or g_117138_(_059116_, _059117_, _059118_);
  or g_117139_(_059115_, _059118_, _059119_);
  xor g_117140_(out[92], out[684], _059120_);
  or g_117141_(_059095_, _059120_, _059121_);
  or g_117142_(_059094_, _059106_, _059122_);
  or g_117143_(_059121_, _059122_, _059123_);
  or g_117144_(_059098_, _059104_, _059125_);
  or g_117145_(_059107_, _059125_, _059126_);
  or g_117146_(_059123_, _059126_, _059127_);
  or g_117147_(_059119_, _059127_, _059128_);
  or g_117148_(_059111_, _059128_, _059129_);
  xor g_117149_(out[76], out[684], _059130_);
  and g_117150_(_098118_, out[683], _059131_);
  xor g_117151_(out[72], out[680], _059132_);
  xor g_117152_(out[70], out[678], _059133_);
  xor g_117153_(out[77], out[685], _059134_);
  xor g_117154_(out[78], out[686], _059136_);
  xor g_117155_(out[66], out[674], _059137_);
  xor g_117156_(out[73], out[681], _059138_);
  xor g_117157_(out[69], out[677], _059139_);
  xor g_117158_(out[65], out[673], _059140_);
  and g_117159_(out[75], _049631_, _059141_);
  or g_117160_(_059132_, _059134_, _059142_);
  xor g_117161_(out[79], out[687], _059143_);
  xor g_117162_(out[74], out[682], _059144_);
  xor g_117163_(out[68], out[676], _059145_);
  xor g_117164_(out[67], out[675], _059147_);
  xor g_117165_(out[64], out[672], _059148_);
  or g_117166_(_059137_, _059144_, _059149_);
  or g_117167_(_059142_, _059149_, _059150_);
  or g_117168_(_059138_, _059147_, _059151_);
  or g_117169_(_059139_, _059151_, _059152_);
  or g_117170_(_059150_, _059152_, _059153_);
  or g_117171_(_059136_, _059145_, _059154_);
  or g_117172_(_059153_, _059154_, _059155_);
  or g_117173_(_059130_, _059131_, _059156_);
  xor g_117174_(out[71], out[679], _059158_);
  or g_117175_(_059133_, _059158_, _059159_);
  or g_117176_(_059156_, _059159_, _059160_);
  or g_117177_(_059140_, _059141_, _059161_);
  or g_117178_(_059143_, _059161_, _059162_);
  or g_117179_(_059160_, _059162_, _059163_);
  or g_117180_(_059148_, _059163_, _059164_);
  or g_117181_(_059155_, _059164_, _059165_);
  not g_117182_(_059165_, _059166_);
  xor g_117183_(out[55], out[679], _059167_);
  and g_117184_(_098107_, out[683], _059169_);
  xor g_117185_(out[62], out[686], _059170_);
  xor g_117186_(out[56], out[680], _059171_);
  xor g_117187_(out[49], out[673], _059172_);
  xor g_117188_(out[61], out[685], _059173_);
  xor g_117189_(out[57], out[681], _059174_);
  xor g_117190_(out[52], out[676], _059175_);
  xor g_117191_(out[50], out[674], _059176_);
  and g_117192_(out[59], _049631_, _059177_);
  xor g_117193_(out[51], out[675], _059178_);
  xor g_117194_(out[54], out[678], _059180_);
  xor g_117195_(out[63], out[687], _059181_);
  xor g_117196_(out[58], out[682], _059182_);
  xor g_117197_(out[53], out[677], _059183_);
  xor g_117198_(out[48], out[672], _059184_);
  or g_117199_(_059170_, _059175_, _059185_);
  or g_117200_(_059171_, _059173_, _059186_);
  or g_117201_(_059176_, _059182_, _059187_);
  or g_117202_(_059186_, _059187_, _059188_);
  or g_117203_(_059174_, _059178_, _059189_);
  or g_117204_(_059183_, _059184_, _059191_);
  or g_117205_(_059189_, _059191_, _059192_);
  or g_117206_(_059188_, _059192_, _059193_);
  xor g_117207_(out[60], out[684], _059194_);
  or g_117208_(_059169_, _059194_, _059195_);
  or g_117209_(_059167_, _059180_, _059196_);
  or g_117210_(_059195_, _059196_, _059197_);
  or g_117211_(_059172_, _059177_, _059198_);
  or g_117212_(_059181_, _059198_, _059199_);
  or g_117213_(_059197_, _059199_, _059200_);
  or g_117214_(_059193_, _059200_, _059202_);
  or g_117215_(_059185_, _059202_, _059203_);
  not g_117216_(_059203_, _059204_);
  xor g_117217_(out[33], out[673], _059205_);
  and g_117218_(out[43], _049631_, _059206_);
  xor g_117219_(out[41], out[681], _059207_);
  xor g_117220_(out[32], out[672], _059208_);
  xor g_117221_(out[46], out[686], _059209_);
  xor g_117222_(out[36], out[676], _059210_);
  or g_117223_(_059209_, _059210_, _059211_);
  xor g_117224_(out[45], out[685], _059213_);
  xor g_117225_(out[35], out[675], _059214_);
  and g_117226_(_098096_, out[683], _059215_);
  xor g_117227_(out[38], out[678], _059216_);
  xor g_117228_(out[42], out[682], _059217_);
  xor g_117229_(out[37], out[677], _059218_);
  xor g_117230_(out[47], out[687], _059219_);
  xor g_117231_(out[40], out[680], _059220_);
  or g_117232_(_059213_, _059220_, _059221_);
  xor g_117233_(out[34], out[674], _059222_);
  or g_117234_(_059217_, _059222_, _059224_);
  or g_117235_(_059221_, _059224_, _059225_);
  or g_117236_(_059207_, _059214_, _059226_);
  or g_117237_(_059218_, _059226_, _059227_);
  or g_117238_(_059225_, _059227_, _059228_);
  or g_117239_(_059211_, _059228_, _059229_);
  xor g_117240_(out[44], out[684], _059230_);
  or g_117241_(_059215_, _059230_, _059231_);
  xor g_117242_(out[39], out[679], _059232_);
  or g_117243_(_059216_, _059232_, _059233_);
  or g_117244_(_059231_, _059233_, _059235_);
  or g_117245_(_059205_, _059206_, _059236_);
  or g_117246_(_059219_, _059236_, _059237_);
  or g_117247_(_059235_, _059237_, _059238_);
  or g_117248_(_059208_, _059238_, _059239_);
  or g_117249_(_059229_, _059239_, _059240_);
  xor g_117250_(out[23], out[679], _059241_);
  and g_117251_(_098063_, out[683], _059242_);
  xor g_117252_(out[30], out[686], _059243_);
  xor g_117253_(out[24], out[680], _059244_);
  xor g_117254_(out[17], out[673], _059246_);
  xor g_117255_(out[29], out[685], _059247_);
  xor g_117256_(out[25], out[681], _059248_);
  xor g_117257_(out[20], out[676], _059249_);
  xor g_117258_(out[18], out[674], _059250_);
  and g_117259_(out[27], _049631_, _059251_);
  xor g_117260_(out[19], out[675], _059252_);
  xor g_117261_(out[22], out[678], _059253_);
  xor g_117262_(out[31], out[687], _059254_);
  xor g_117263_(out[26], out[682], _059255_);
  xor g_117264_(out[21], out[677], _059257_);
  xor g_117265_(out[16], out[672], _059258_);
  or g_117266_(_059243_, _059249_, _059259_);
  or g_117267_(_059244_, _059247_, _059260_);
  or g_117268_(_059250_, _059255_, _059261_);
  or g_117269_(_059260_, _059261_, _059262_);
  or g_117270_(_059248_, _059252_, _059263_);
  or g_117271_(_059257_, _059258_, _059264_);
  or g_117272_(_059263_, _059264_, _059265_);
  or g_117273_(_059262_, _059265_, _059266_);
  xor g_117274_(out[28], out[684], _059268_);
  or g_117275_(_059242_, _059268_, _059269_);
  or g_117276_(_059241_, _059253_, _059270_);
  or g_117277_(_059269_, _059270_, _059271_);
  or g_117278_(_059246_, _059251_, _059272_);
  or g_117279_(_059254_, _059272_, _059273_);
  or g_117280_(_059271_, _059273_, _059274_);
  or g_117281_(_059266_, _059274_, _059275_);
  or g_117282_(_059259_, _059275_, _059276_);
  and g_117283_(_098041_, out[683], _059277_);
  and g_117284_(out[11], _049631_, _059279_);
  xor g_117285_(out[4], out[676], _059280_);
  xor g_117286_(out[14], out[686], _059281_);
  or g_117287_(_059280_, _059281_, _059282_);
  xor g_117288_(out[13], out[685], _059283_);
  xor g_117289_(out[3], out[675], _059284_);
  xor g_117290_(out[0], out[672], _059285_);
  xor g_117291_(out[10], out[682], _059286_);
  xor g_117292_(out[15], out[687], _059287_);
  xor g_117293_(out[6], out[678], _059288_);
  xor g_117294_(out[5], out[677], _059290_);
  xor g_117295_(out[8], out[680], _059291_);
  or g_117296_(_059283_, _059291_, _059292_);
  xor g_117297_(out[2], out[674], _059293_);
  xor g_117298_(out[9], out[681], _059294_);
  xor g_117299_(out[1], out[673], _059295_);
  or g_117300_(_059286_, _059293_, _059296_);
  or g_117301_(_059292_, _059296_, _059297_);
  or g_117302_(_059284_, _059294_, _059298_);
  or g_117303_(_059290_, _059298_, _059299_);
  or g_117304_(_059297_, _059299_, _059301_);
  or g_117305_(_059282_, _059301_, _059302_);
  xor g_117306_(out[12], out[684], _059303_);
  or g_117307_(_059277_, _059303_, _059304_);
  xor g_117308_(out[7], out[679], _059305_);
  or g_117309_(_059288_, _059305_, _059306_);
  or g_117310_(_059304_, _059306_, _059307_);
  or g_117311_(_059279_, _059295_, _059308_);
  or g_117312_(_059287_, _059308_, _059309_);
  or g_117313_(_059307_, _059309_, _059310_);
  or g_117314_(_059285_, _059310_, _059312_);
  or g_117315_(_059302_, _059312_, _059313_);
  xor g_117316_(out[465], out[657], _059314_);
  and g_117317_(_049499_, out[667], _059315_);
  and g_117318_(out[475], _049620_, _059316_);
  xor g_117319_(out[473], out[665], _059317_);
  xor g_117320_(out[464], out[656], _059318_);
  xor g_117321_(out[478], out[670], _059319_);
  xor g_117322_(out[468], out[660], _059320_);
  or g_117323_(_059319_, _059320_, _059321_);
  xor g_117324_(out[477], out[669], _059323_);
  xor g_117325_(out[467], out[659], _059324_);
  xor g_117326_(out[476], out[668], _059325_);
  xor g_117327_(out[470], out[662], _059326_);
  xor g_117328_(out[474], out[666], _059327_);
  xor g_117329_(out[469], out[661], _059328_);
  xor g_117330_(out[479], out[671], _059329_);
  xor g_117331_(out[472], out[664], _059330_);
  or g_117332_(_059323_, _059330_, _059331_);
  xor g_117333_(out[466], out[658], _059332_);
  or g_117334_(_059327_, _059332_, _059334_);
  or g_117335_(_059331_, _059334_, _059335_);
  or g_117336_(_059317_, _059324_, _059336_);
  or g_117337_(_059328_, _059336_, _059337_);
  or g_117338_(_059335_, _059337_, _059338_);
  or g_117339_(_059321_, _059338_, _059339_);
  or g_117340_(_059315_, _059325_, _059340_);
  xor g_117341_(out[471], out[663], _059341_);
  or g_117342_(_059326_, _059341_, _059342_);
  or g_117343_(_059340_, _059342_, _059343_);
  or g_117344_(_059314_, _059316_, _059345_);
  or g_117345_(_059329_, _059345_, _059346_);
  or g_117346_(_059343_, _059346_, _059347_);
  or g_117347_(_059318_, _059347_, _059348_);
  or g_117348_(_059339_, _059348_, _059349_);
  xor g_117349_(out[455], out[663], _059350_);
  and g_117350_(_049477_, out[667], _059351_);
  xor g_117351_(out[462], out[670], _059352_);
  xor g_117352_(out[456], out[664], _059353_);
  xor g_117353_(out[449], out[657], _059354_);
  xor g_117354_(out[461], out[669], _059356_);
  xor g_117355_(out[457], out[665], _059357_);
  xor g_117356_(out[452], out[660], _059358_);
  xor g_117357_(out[450], out[658], _059359_);
  and g_117358_(out[459], _049620_, _059360_);
  xor g_117359_(out[451], out[659], _059361_);
  xor g_117360_(out[454], out[662], _059362_);
  xor g_117361_(out[463], out[671], _059363_);
  xor g_117362_(out[458], out[666], _059364_);
  xor g_117363_(out[453], out[661], _059365_);
  xor g_117364_(out[448], out[656], _059367_);
  or g_117365_(_059352_, _059358_, _059368_);
  or g_117366_(_059353_, _059356_, _059369_);
  or g_117367_(_059359_, _059364_, _059370_);
  or g_117368_(_059369_, _059370_, _059371_);
  or g_117369_(_059357_, _059361_, _059372_);
  or g_117370_(_059365_, _059367_, _059373_);
  or g_117371_(_059372_, _059373_, _059374_);
  or g_117372_(_059371_, _059374_, _059375_);
  xor g_117373_(out[460], out[668], _059376_);
  or g_117374_(_059351_, _059376_, _059378_);
  or g_117375_(_059350_, _059362_, _059379_);
  or g_117376_(_059378_, _059379_, _059380_);
  or g_117377_(_059354_, _059360_, _059381_);
  or g_117378_(_059363_, _059381_, _059382_);
  or g_117379_(_059380_, _059382_, _059383_);
  or g_117380_(_059375_, _059383_, _059384_);
  or g_117381_(_059368_, _059384_, _059385_);
  xor g_117382_(out[433], out[657], _059386_);
  and g_117383_(out[443], _049620_, _059387_);
  xor g_117384_(out[441], out[665], _059389_);
  xor g_117385_(out[432], out[656], _059390_);
  xor g_117386_(out[446], out[670], _059391_);
  xor g_117387_(out[436], out[660], _059392_);
  or g_117388_(_059391_, _059392_, _059393_);
  xor g_117389_(out[445], out[669], _059394_);
  xor g_117390_(out[435], out[659], _059395_);
  and g_117391_(_049466_, out[667], _059396_);
  xor g_117392_(out[438], out[662], _059397_);
  xor g_117393_(out[442], out[666], _059398_);
  xor g_117394_(out[437], out[661], _059400_);
  xor g_117395_(out[447], out[671], _059401_);
  xor g_117396_(out[440], out[664], _059402_);
  or g_117397_(_059394_, _059402_, _059403_);
  xor g_117398_(out[434], out[658], _059404_);
  or g_117399_(_059398_, _059404_, _059405_);
  or g_117400_(_059403_, _059405_, _059406_);
  or g_117401_(_059389_, _059395_, _059407_);
  or g_117402_(_059400_, _059407_, _059408_);
  or g_117403_(_059406_, _059408_, _059409_);
  or g_117404_(_059393_, _059409_, _059411_);
  xor g_117405_(out[444], out[668], _059412_);
  or g_117406_(_059396_, _059412_, _059413_);
  xor g_117407_(out[439], out[663], _059414_);
  or g_117408_(_059397_, _059414_, _059415_);
  or g_117409_(_059413_, _059415_, _059416_);
  or g_117410_(_059386_, _059387_, _059417_);
  or g_117411_(_059401_, _059417_, _059418_);
  or g_117412_(_059416_, _059418_, _059419_);
  or g_117413_(_059390_, _059419_, _059420_);
  or g_117414_(_059411_, _059420_, _059422_);
  xor g_117415_(out[423], out[663], _059423_);
  and g_117416_(_049455_, out[667], _059424_);
  xor g_117417_(out[430], out[670], _059425_);
  xor g_117418_(out[424], out[664], _059426_);
  xor g_117419_(out[417], out[657], _059427_);
  xor g_117420_(out[429], out[669], _059428_);
  xor g_117421_(out[425], out[665], _059429_);
  xor g_117422_(out[420], out[660], _059430_);
  xor g_117423_(out[418], out[658], _059431_);
  and g_117424_(out[427], _049620_, _059433_);
  xor g_117425_(out[419], out[659], _059434_);
  xor g_117426_(out[422], out[662], _059435_);
  xor g_117427_(out[431], out[671], _059436_);
  xor g_117428_(out[426], out[666], _059437_);
  xor g_117429_(out[421], out[661], _059438_);
  xor g_117430_(out[416], out[656], _059439_);
  or g_117431_(_059425_, _059430_, _059440_);
  or g_117432_(_059426_, _059428_, _059441_);
  or g_117433_(_059431_, _059437_, _059442_);
  or g_117434_(_059441_, _059442_, _059444_);
  or g_117435_(_059429_, _059434_, _059445_);
  or g_117436_(_059438_, _059439_, _059446_);
  or g_117437_(_059445_, _059446_, _059447_);
  or g_117438_(_059444_, _059447_, _059448_);
  xor g_117439_(out[428], out[668], _059449_);
  or g_117440_(_059424_, _059449_, _059450_);
  or g_117441_(_059423_, _059435_, _059451_);
  or g_117442_(_059450_, _059451_, _059452_);
  or g_117443_(_059427_, _059433_, _059453_);
  or g_117444_(_059436_, _059453_, _059455_);
  or g_117445_(_059452_, _059455_, _059456_);
  or g_117446_(_059448_, _059456_, _059457_);
  or g_117447_(_059440_, _059457_, _059458_);
  xor g_117448_(out[401], out[657], _059459_);
  and g_117449_(out[411], _049620_, _059460_);
  xor g_117450_(out[409], out[665], _059461_);
  xor g_117451_(out[400], out[656], _059462_);
  xor g_117452_(out[414], out[670], _059463_);
  xor g_117453_(out[404], out[660], _059464_);
  or g_117454_(_059463_, _059464_, _059466_);
  xor g_117455_(out[413], out[669], _059467_);
  xor g_117456_(out[403], out[659], _059468_);
  and g_117457_(_049444_, out[667], _059469_);
  xor g_117458_(out[406], out[662], _059470_);
  xor g_117459_(out[410], out[666], _059471_);
  xor g_117460_(out[405], out[661], _059472_);
  xor g_117461_(out[415], out[671], _059473_);
  xor g_117462_(out[408], out[664], _059474_);
  or g_117463_(_059467_, _059474_, _059475_);
  xor g_117464_(out[402], out[658], _059477_);
  or g_117465_(_059471_, _059477_, _059478_);
  or g_117466_(_059475_, _059478_, _059479_);
  or g_117467_(_059461_, _059468_, _059480_);
  or g_117468_(_059472_, _059480_, _059481_);
  or g_117469_(_059479_, _059481_, _059482_);
  or g_117470_(_059466_, _059482_, _059483_);
  xor g_117471_(out[412], out[668], _059484_);
  or g_117472_(_059469_, _059484_, _059485_);
  xor g_117473_(out[407], out[663], _059486_);
  or g_117474_(_059470_, _059486_, _059488_);
  or g_117475_(_059485_, _059488_, _059489_);
  or g_117476_(_059459_, _059460_, _059490_);
  or g_117477_(_059473_, _059490_, _059491_);
  or g_117478_(_059489_, _059491_, _059492_);
  or g_117479_(_059462_, _059492_, _059493_);
  or g_117480_(_059483_, _059493_, _059494_);
  xor g_117481_(out[391], out[663], _059495_);
  and g_117482_(_049433_, out[667], _059496_);
  xor g_117483_(out[398], out[670], _059497_);
  xor g_117484_(out[392], out[664], _059499_);
  xor g_117485_(out[385], out[657], _059500_);
  xor g_117486_(out[397], out[669], _059501_);
  xor g_117487_(out[393], out[665], _059502_);
  xor g_117488_(out[388], out[660], _059503_);
  xor g_117489_(out[386], out[658], _059504_);
  and g_117490_(out[395], _049620_, _059505_);
  xor g_117491_(out[387], out[659], _059506_);
  xor g_117492_(out[390], out[662], _059507_);
  xor g_117493_(out[399], out[671], _059508_);
  xor g_117494_(out[394], out[666], _059510_);
  xor g_117495_(out[389], out[661], _059511_);
  xor g_117496_(out[384], out[656], _059512_);
  or g_117497_(_059497_, _059503_, _059513_);
  or g_117498_(_059499_, _059501_, _059514_);
  or g_117499_(_059504_, _059510_, _059515_);
  or g_117500_(_059514_, _059515_, _059516_);
  or g_117501_(_059502_, _059506_, _059517_);
  or g_117502_(_059511_, _059512_, _059518_);
  or g_117503_(_059517_, _059518_, _059519_);
  or g_117504_(_059516_, _059519_, _059521_);
  xor g_117505_(out[396], out[668], _059522_);
  or g_117506_(_059496_, _059522_, _059523_);
  or g_117507_(_059495_, _059507_, _059524_);
  or g_117508_(_059523_, _059524_, _059525_);
  or g_117509_(_059500_, _059505_, _059526_);
  or g_117510_(_059508_, _059526_, _059527_);
  or g_117511_(_059525_, _059527_, _059528_);
  or g_117512_(_059521_, _059528_, _059529_);
  or g_117513_(_059513_, _059529_, _059530_);
  xor g_117514_(out[369], out[657], _059532_);
  and g_117515_(out[379], _049620_, _059533_);
  xor g_117516_(out[382], out[670], _059534_);
  xor g_117517_(out[371], out[659], _059535_);
  xor g_117518_(out[372], out[660], _059536_);
  xor g_117519_(out[370], out[658], _059537_);
  xor g_117520_(out[377], out[665], _059538_);
  xor g_117521_(out[368], out[656], _059539_);
  and g_117522_(_049422_, out[667], _059540_);
  xor g_117523_(out[374], out[662], _059541_);
  xor g_117524_(out[378], out[666], _059543_);
  xor g_117525_(out[373], out[661], _059544_);
  xor g_117526_(out[383], out[671], _059545_);
  xor g_117527_(out[381], out[669], _059546_);
  xor g_117528_(out[376], out[664], _059547_);
  or g_117529_(_059534_, _059536_, _059548_);
  or g_117530_(_059546_, _059547_, _059549_);
  or g_117531_(_059537_, _059543_, _059550_);
  or g_117532_(_059549_, _059550_, _059551_);
  or g_117533_(_059535_, _059538_, _059552_);
  or g_117534_(_059539_, _059544_, _059554_);
  or g_117535_(_059552_, _059554_, _059555_);
  or g_117536_(_059551_, _059555_, _059556_);
  xor g_117537_(out[380], out[668], _059557_);
  or g_117538_(_059540_, _059557_, _059558_);
  xor g_117539_(out[375], out[663], _059559_);
  or g_117540_(_059541_, _059559_, _059560_);
  or g_117541_(_059558_, _059560_, _059561_);
  or g_117542_(_059532_, _059533_, _059562_);
  or g_117543_(_059545_, _059562_, _059563_);
  or g_117544_(_059561_, _059563_, _059565_);
  or g_117545_(_059556_, _059565_, _059566_);
  or g_117546_(_059548_, _059566_, _059567_);
  xor g_117547_(out[359], out[663], _059568_);
  and g_117548_(_049411_, out[667], _059569_);
  xor g_117549_(out[366], out[670], _059570_);
  xor g_117550_(out[360], out[664], _059571_);
  xor g_117551_(out[353], out[657], _059572_);
  xor g_117552_(out[365], out[669], _059573_);
  xor g_117553_(out[361], out[665], _059574_);
  xor g_117554_(out[356], out[660], _059576_);
  xor g_117555_(out[354], out[658], _059577_);
  and g_117556_(out[363], _049620_, _059578_);
  xor g_117557_(out[355], out[659], _059579_);
  xor g_117558_(out[358], out[662], _059580_);
  xor g_117559_(out[367], out[671], _059581_);
  xor g_117560_(out[362], out[666], _059582_);
  xor g_117561_(out[357], out[661], _059583_);
  xor g_117562_(out[352], out[656], _059584_);
  or g_117563_(_059570_, _059576_, _059585_);
  or g_117564_(_059571_, _059573_, _059587_);
  or g_117565_(_059577_, _059582_, _059588_);
  or g_117566_(_059587_, _059588_, _059589_);
  or g_117567_(_059574_, _059579_, _059590_);
  or g_117568_(_059583_, _059584_, _059591_);
  or g_117569_(_059590_, _059591_, _059592_);
  or g_117570_(_059589_, _059592_, _059593_);
  xor g_117571_(out[364], out[668], _059594_);
  or g_117572_(_059569_, _059594_, _059595_);
  or g_117573_(_059568_, _059580_, _059596_);
  or g_117574_(_059595_, _059596_, _059598_);
  or g_117575_(_059572_, _059578_, _059599_);
  or g_117576_(_059581_, _059599_, _059600_);
  or g_117577_(_059598_, _059600_, _059601_);
  or g_117578_(_059593_, _059601_, _059602_);
  or g_117579_(_059585_, _059602_, _059603_);
  not g_117580_(_059603_, _059604_);
  xor g_117581_(out[340], out[660], _059605_);
  xor g_117582_(out[348], out[668], _059606_);
  and g_117583_(_049400_, out[667], _059607_);
  xor g_117584_(out[346], out[666], _059609_);
  xor g_117585_(out[342], out[662], _059610_);
  xor g_117586_(out[341], out[661], _059611_);
  xor g_117587_(out[339], out[659], _059612_);
  xor g_117588_(out[349], out[669], _059613_);
  xor g_117589_(out[350], out[670], _059614_);
  xor g_117590_(out[337], out[657], _059615_);
  xor g_117591_(out[338], out[658], _059616_);
  and g_117592_(out[347], _049620_, _059617_);
  xor g_117593_(out[336], out[656], _059618_);
  xor g_117594_(out[351], out[671], _059620_);
  xor g_117595_(out[344], out[664], _059621_);
  or g_117596_(_059613_, _059621_, _059622_);
  xor g_117597_(out[345], out[665], _059623_);
  or g_117598_(_059609_, _059616_, _059624_);
  or g_117599_(_059622_, _059624_, _059625_);
  or g_117600_(_059612_, _059623_, _059626_);
  or g_117601_(_059611_, _059626_, _059627_);
  or g_117602_(_059625_, _059627_, _059628_);
  or g_117603_(_059605_, _059614_, _059629_);
  or g_117604_(_059628_, _059629_, _059631_);
  or g_117605_(_059606_, _059607_, _059632_);
  xor g_117606_(out[343], out[663], _059633_);
  or g_117607_(_059610_, _059633_, _059634_);
  or g_117608_(_059632_, _059634_, _059635_);
  or g_117609_(_059615_, _059617_, _059636_);
  or g_117610_(_059620_, _059636_, _059637_);
  or g_117611_(_059635_, _059637_, _059638_);
  or g_117612_(_059618_, _059638_, _059639_);
  or g_117613_(_059631_, _059639_, _059640_);
  not g_117614_(_059640_, _059642_);
  xor g_117615_(out[327], out[663], _059643_);
  and g_117616_(_098294_, out[667], _059644_);
  xor g_117617_(out[334], out[670], _059645_);
  xor g_117618_(out[328], out[664], _059646_);
  xor g_117619_(out[321], out[657], _059647_);
  xor g_117620_(out[333], out[669], _059648_);
  xor g_117621_(out[329], out[665], _059649_);
  xor g_117622_(out[324], out[660], _059650_);
  xor g_117623_(out[322], out[658], _059651_);
  and g_117624_(out[331], _049620_, _059653_);
  xor g_117625_(out[323], out[659], _059654_);
  xor g_117626_(out[326], out[662], _059655_);
  xor g_117627_(out[335], out[671], _059656_);
  xor g_117628_(out[330], out[666], _059657_);
  xor g_117629_(out[325], out[661], _059658_);
  xor g_117630_(out[320], out[656], _059659_);
  or g_117631_(_059645_, _059650_, _059660_);
  or g_117632_(_059646_, _059648_, _059661_);
  or g_117633_(_059651_, _059657_, _059662_);
  or g_117634_(_059661_, _059662_, _059664_);
  or g_117635_(_059649_, _059654_, _059665_);
  or g_117636_(_059658_, _059659_, _059666_);
  or g_117637_(_059665_, _059666_, _059667_);
  or g_117638_(_059664_, _059667_, _059668_);
  xor g_117639_(out[332], out[668], _059669_);
  or g_117640_(_059644_, _059669_, _059670_);
  or g_117641_(_059643_, _059655_, _059671_);
  or g_117642_(_059670_, _059671_, _059672_);
  or g_117643_(_059647_, _059653_, _059673_);
  or g_117644_(_059656_, _059673_, _059675_);
  or g_117645_(_059672_, _059675_, _059676_);
  or g_117646_(_059668_, _059676_, _059677_);
  or g_117647_(_059660_, _059677_, _059678_);
  xor g_117648_(out[312], out[664], _059679_);
  xor g_117649_(out[309], out[661], _059680_);
  xor g_117650_(out[307], out[659], _059681_);
  xor g_117651_(out[318], out[670], _059682_);
  xor g_117652_(out[317], out[669], _059683_);
  xor g_117653_(out[306], out[658], _059684_);
  xor g_117654_(out[313], out[665], _059686_);
  xor g_117655_(out[310], out[662], _059687_);
  xor g_117656_(out[319], out[671], _059688_);
  xor g_117657_(out[314], out[666], _059689_);
  xor g_117658_(out[308], out[660], _059690_);
  xor g_117659_(out[304], out[656], _059691_);
  and g_117660_(_098283_, out[667], _059692_);
  and g_117661_(out[315], _049620_, _059693_);
  or g_117662_(_059679_, _059683_, _059694_);
  xor g_117663_(out[305], out[657], _059695_);
  or g_117664_(_059684_, _059689_, _059697_);
  or g_117665_(_059694_, _059697_, _059698_);
  or g_117666_(_059681_, _059686_, _059699_);
  or g_117667_(_059680_, _059699_, _059700_);
  or g_117668_(_059698_, _059700_, _059701_);
  or g_117669_(_059682_, _059690_, _059702_);
  or g_117670_(_059701_, _059702_, _059703_);
  xor g_117671_(out[316], out[668], _059704_);
  or g_117672_(_059692_, _059704_, _059705_);
  xor g_117673_(out[311], out[663], _059706_);
  or g_117674_(_059687_, _059706_, _059708_);
  or g_117675_(_059705_, _059708_, _059709_);
  or g_117676_(_059693_, _059695_, _059710_);
  or g_117677_(_059688_, _059710_, _059711_);
  or g_117678_(_059709_, _059711_, _059712_);
  or g_117679_(_059691_, _059712_, _059713_);
  or g_117680_(_059703_, _059713_, _059714_);
  xor g_117681_(out[295], out[663], _059715_);
  and g_117682_(_098272_, out[667], _059716_);
  xor g_117683_(out[302], out[670], _059717_);
  xor g_117684_(out[296], out[664], _059719_);
  xor g_117685_(out[289], out[657], _059720_);
  xor g_117686_(out[301], out[669], _059721_);
  xor g_117687_(out[297], out[665], _059722_);
  xor g_117688_(out[292], out[660], _059723_);
  xor g_117689_(out[290], out[658], _059724_);
  and g_117690_(out[299], _049620_, _059725_);
  xor g_117691_(out[291], out[659], _059726_);
  xor g_117692_(out[294], out[662], _059727_);
  xor g_117693_(out[303], out[671], _059728_);
  xor g_117694_(out[298], out[666], _059730_);
  xor g_117695_(out[293], out[661], _059731_);
  xor g_117696_(out[288], out[656], _059732_);
  or g_117697_(_059717_, _059723_, _059733_);
  or g_117698_(_059719_, _059721_, _059734_);
  or g_117699_(_059724_, _059730_, _059735_);
  or g_117700_(_059734_, _059735_, _059736_);
  or g_117701_(_059722_, _059726_, _059737_);
  or g_117702_(_059731_, _059732_, _059738_);
  or g_117703_(_059737_, _059738_, _059739_);
  or g_117704_(_059736_, _059739_, _059741_);
  xor g_117705_(out[300], out[668], _059742_);
  or g_117706_(_059716_, _059742_, _059743_);
  or g_117707_(_059715_, _059727_, _059744_);
  or g_117708_(_059743_, _059744_, _059745_);
  or g_117709_(_059720_, _059725_, _059746_);
  or g_117710_(_059728_, _059746_, _059747_);
  or g_117711_(_059745_, _059747_, _059748_);
  or g_117712_(_059741_, _059748_, _059749_);
  or g_117713_(_059733_, _059749_, _059750_);
  not g_117714_(_059750_, _059752_);
  and g_117715_(out[283], _049620_, _059753_);
  xor g_117716_(out[276], out[660], _059754_);
  xor g_117717_(out[286], out[670], _059755_);
  or g_117718_(_059754_, _059755_, _059756_);
  xor g_117719_(out[285], out[669], _059757_);
  xor g_117720_(out[275], out[659], _059758_);
  xor g_117721_(out[272], out[656], _059759_);
  and g_117722_(_098261_, out[667], _059760_);
  xor g_117723_(out[282], out[666], _059761_);
  xor g_117724_(out[287], out[671], _059763_);
  xor g_117725_(out[278], out[662], _059764_);
  xor g_117726_(out[277], out[661], _059765_);
  xor g_117727_(out[280], out[664], _059766_);
  or g_117728_(_059757_, _059766_, _059767_);
  xor g_117729_(out[274], out[658], _059768_);
  xor g_117730_(out[281], out[665], _059769_);
  xor g_117731_(out[273], out[657], _059770_);
  or g_117732_(_059761_, _059768_, _059771_);
  or g_117733_(_059767_, _059771_, _059772_);
  or g_117734_(_059758_, _059769_, _059774_);
  or g_117735_(_059765_, _059774_, _059775_);
  or g_117736_(_059772_, _059775_, _059776_);
  or g_117737_(_059756_, _059776_, _059777_);
  xor g_117738_(out[284], out[668], _059778_);
  or g_117739_(_059760_, _059778_, _059779_);
  xor g_117740_(out[279], out[663], _059780_);
  or g_117741_(_059764_, _059780_, _059781_);
  or g_117742_(_059779_, _059781_, _059782_);
  or g_117743_(_059753_, _059770_, _059783_);
  or g_117744_(_059763_, _059783_, _059785_);
  or g_117745_(_059782_, _059785_, _059786_);
  or g_117746_(_059759_, _059786_, _059787_);
  or g_117747_(_059777_, _059787_, _059788_);
  xor g_117748_(out[263], out[663], _059789_);
  and g_117749_(_098250_, out[667], _059790_);
  xor g_117750_(out[270], out[670], _059791_);
  xor g_117751_(out[264], out[664], _059792_);
  xor g_117752_(out[257], out[657], _059793_);
  xor g_117753_(out[269], out[669], _059794_);
  xor g_117754_(out[265], out[665], _059796_);
  xor g_117755_(out[260], out[660], _059797_);
  xor g_117756_(out[258], out[658], _059798_);
  and g_117757_(out[267], _049620_, _059799_);
  xor g_117758_(out[259], out[659], _059800_);
  xor g_117759_(out[262], out[662], _059801_);
  xor g_117760_(out[271], out[671], _059802_);
  xor g_117761_(out[266], out[666], _059803_);
  xor g_117762_(out[261], out[661], _059804_);
  xor g_117763_(out[256], out[656], _059805_);
  or g_117764_(_059791_, _059797_, _059807_);
  or g_117765_(_059792_, _059794_, _059808_);
  or g_117766_(_059798_, _059803_, _059809_);
  or g_117767_(_059808_, _059809_, _059810_);
  or g_117768_(_059796_, _059800_, _059811_);
  or g_117769_(_059804_, _059805_, _059812_);
  or g_117770_(_059811_, _059812_, _059813_);
  or g_117771_(_059810_, _059813_, _059814_);
  xor g_117772_(out[268], out[668], _059815_);
  or g_117773_(_059790_, _059815_, _059816_);
  or g_117774_(_059789_, _059801_, _059818_);
  or g_117775_(_059816_, _059818_, _059819_);
  or g_117776_(_059793_, _059799_, _059820_);
  or g_117777_(_059802_, _059820_, _059821_);
  or g_117778_(_059819_, _059821_, _059822_);
  or g_117779_(_059814_, _059822_, _059823_);
  or g_117780_(_059807_, _059823_, _059824_);
  xor g_117781_(out[248], out[664], _059825_);
  xor g_117782_(out[245], out[661], _059826_);
  xor g_117783_(out[243], out[659], _059827_);
  xor g_117784_(out[254], out[670], _059829_);
  xor g_117785_(out[253], out[669], _059830_);
  xor g_117786_(out[242], out[658], _059831_);
  xor g_117787_(out[249], out[665], _059832_);
  xor g_117788_(out[246], out[662], _059833_);
  xor g_117789_(out[255], out[671], _059834_);
  xor g_117790_(out[250], out[666], _059835_);
  xor g_117791_(out[244], out[660], _059836_);
  xor g_117792_(out[240], out[656], _059837_);
  and g_117793_(_098239_, out[667], _059838_);
  and g_117794_(out[251], _049620_, _059840_);
  or g_117795_(_059825_, _059830_, _059841_);
  xor g_117796_(out[241], out[657], _059842_);
  or g_117797_(_059831_, _059835_, _059843_);
  or g_117798_(_059841_, _059843_, _059844_);
  or g_117799_(_059827_, _059832_, _059845_);
  or g_117800_(_059826_, _059845_, _059846_);
  or g_117801_(_059844_, _059846_, _059847_);
  or g_117802_(_059829_, _059836_, _059848_);
  or g_117803_(_059847_, _059848_, _059849_);
  xor g_117804_(out[252], out[668], _059851_);
  or g_117805_(_059838_, _059851_, _059852_);
  xor g_117806_(out[247], out[663], _059853_);
  or g_117807_(_059833_, _059853_, _059854_);
  or g_117808_(_059852_, _059854_, _059855_);
  or g_117809_(_059840_, _059842_, _059856_);
  or g_117810_(_059834_, _059856_, _059857_);
  or g_117811_(_059855_, _059857_, _059858_);
  or g_117812_(_059837_, _059858_, _059859_);
  or g_117813_(_059849_, _059859_, _059860_);
  not g_117814_(_059860_, _059862_);
  xor g_117815_(out[231], out[663], _059863_);
  and g_117816_(_098228_, out[667], _059864_);
  xor g_117817_(out[238], out[670], _059865_);
  xor g_117818_(out[232], out[664], _059866_);
  xor g_117819_(out[225], out[657], _059867_);
  xor g_117820_(out[237], out[669], _059868_);
  xor g_117821_(out[233], out[665], _059869_);
  xor g_117822_(out[228], out[660], _059870_);
  xor g_117823_(out[226], out[658], _059871_);
  and g_117824_(out[235], _049620_, _059873_);
  xor g_117825_(out[227], out[659], _059874_);
  xor g_117826_(out[230], out[662], _059875_);
  xor g_117827_(out[239], out[671], _059876_);
  xor g_117828_(out[234], out[666], _059877_);
  xor g_117829_(out[229], out[661], _059878_);
  xor g_117830_(out[224], out[656], _059879_);
  or g_117831_(_059865_, _059870_, _059880_);
  or g_117832_(_059866_, _059868_, _059881_);
  or g_117833_(_059871_, _059877_, _059882_);
  or g_117834_(_059881_, _059882_, _059884_);
  or g_117835_(_059869_, _059874_, _059885_);
  or g_117836_(_059878_, _059879_, _059886_);
  or g_117837_(_059885_, _059886_, _059887_);
  or g_117838_(_059884_, _059887_, _059888_);
  xor g_117839_(out[236], out[668], _059889_);
  or g_117840_(_059864_, _059889_, _059890_);
  or g_117841_(_059863_, _059875_, _059891_);
  or g_117842_(_059890_, _059891_, _059892_);
  or g_117843_(_059867_, _059873_, _059893_);
  or g_117844_(_059876_, _059893_, _059895_);
  or g_117845_(_059892_, _059895_, _059896_);
  or g_117846_(_059888_, _059896_, _059897_);
  or g_117847_(_059880_, _059897_, _059898_);
  xor g_117848_(out[218], out[666], _059899_);
  xor g_117849_(out[210], out[658], _059900_);
  xor g_117850_(out[209], out[657], _059901_);
  and g_117851_(_098217_, out[667], _059902_);
  and g_117852_(out[219], _049620_, _059903_);
  xor g_117853_(out[221], out[669], _059904_);
  xor g_117854_(out[211], out[659], _059906_);
  xor g_117855_(out[222], out[670], _059907_);
  xor g_117856_(out[220], out[668], _059908_);
  xor g_117857_(out[216], out[664], _059909_);
  xor g_117858_(out[223], out[671], _059910_);
  xor g_117859_(out[213], out[661], _059911_);
  xor g_117860_(out[214], out[662], _059912_);
  xor g_117861_(out[208], out[656], _059913_);
  xor g_117862_(out[212], out[660], _059914_);
  or g_117863_(_059904_, _059909_, _059915_);
  xor g_117864_(out[217], out[665], _059917_);
  or g_117865_(_059899_, _059900_, _059918_);
  or g_117866_(_059915_, _059918_, _059919_);
  or g_117867_(_059906_, _059917_, _059920_);
  or g_117868_(_059911_, _059920_, _059921_);
  or g_117869_(_059919_, _059921_, _059922_);
  or g_117870_(_059907_, _059914_, _059923_);
  or g_117871_(_059922_, _059923_, _059924_);
  or g_117872_(_059902_, _059908_, _059925_);
  xor g_117873_(out[215], out[663], _059926_);
  or g_117874_(_059912_, _059926_, _059928_);
  or g_117875_(_059925_, _059928_, _059929_);
  or g_117876_(_059901_, _059903_, _059930_);
  or g_117877_(_059910_, _059930_, _059931_);
  or g_117878_(_059929_, _059931_, _059932_);
  or g_117879_(_059913_, _059932_, _059933_);
  or g_117880_(_059924_, _059933_, _059934_);
  xor g_117881_(out[199], out[663], _059935_);
  and g_117882_(_098206_, out[667], _059936_);
  xor g_117883_(out[206], out[670], _059937_);
  xor g_117884_(out[200], out[664], _059939_);
  xor g_117885_(out[193], out[657], _059940_);
  xor g_117886_(out[205], out[669], _059941_);
  xor g_117887_(out[201], out[665], _059942_);
  xor g_117888_(out[196], out[660], _059943_);
  xor g_117889_(out[194], out[658], _059944_);
  and g_117890_(out[203], _049620_, _059945_);
  xor g_117891_(out[195], out[659], _059946_);
  xor g_117892_(out[198], out[662], _059947_);
  xor g_117893_(out[207], out[671], _059948_);
  xor g_117894_(out[202], out[666], _059950_);
  xor g_117895_(out[197], out[661], _059951_);
  xor g_117896_(out[192], out[656], _059952_);
  or g_117897_(_059937_, _059943_, _059953_);
  or g_117898_(_059939_, _059941_, _059954_);
  or g_117899_(_059944_, _059950_, _059955_);
  or g_117900_(_059954_, _059955_, _059956_);
  or g_117901_(_059942_, _059946_, _059957_);
  or g_117902_(_059951_, _059952_, _059958_);
  or g_117903_(_059957_, _059958_, _059959_);
  or g_117904_(_059956_, _059959_, _059961_);
  xor g_117905_(out[204], out[668], _059962_);
  or g_117906_(_059936_, _059962_, _059963_);
  or g_117907_(_059935_, _059947_, _059964_);
  or g_117908_(_059963_, _059964_, _059965_);
  or g_117909_(_059940_, _059945_, _059966_);
  or g_117910_(_059948_, _059966_, _059967_);
  or g_117911_(_059965_, _059967_, _059968_);
  or g_117912_(_059961_, _059968_, _059969_);
  or g_117913_(_059953_, _059969_, _059970_);
  xor g_117914_(out[184], out[664], _059972_);
  xor g_117915_(out[181], out[661], _059973_);
  xor g_117916_(out[179], out[659], _059974_);
  xor g_117917_(out[190], out[670], _059975_);
  xor g_117918_(out[189], out[669], _059976_);
  xor g_117919_(out[178], out[658], _059977_);
  xor g_117920_(out[185], out[665], _059978_);
  xor g_117921_(out[182], out[662], _059979_);
  xor g_117922_(out[191], out[671], _059980_);
  xor g_117923_(out[186], out[666], _059981_);
  xor g_117924_(out[180], out[660], _059983_);
  xor g_117925_(out[176], out[656], _059984_);
  and g_117926_(_098195_, out[667], _059985_);
  and g_117927_(out[187], _049620_, _059986_);
  or g_117928_(_059972_, _059976_, _059987_);
  xor g_117929_(out[177], out[657], _059988_);
  or g_117930_(_059977_, _059981_, _059989_);
  or g_117931_(_059987_, _059989_, _059990_);
  or g_117932_(_059974_, _059978_, _059991_);
  or g_117933_(_059973_, _059991_, _059992_);
  or g_117934_(_059990_, _059992_, _059994_);
  or g_117935_(_059975_, _059983_, _059995_);
  or g_117936_(_059994_, _059995_, _059996_);
  xor g_117937_(out[188], out[668], _059997_);
  or g_117938_(_059985_, _059997_, _059998_);
  xor g_117939_(out[183], out[663], _059999_);
  or g_117940_(_059979_, _059999_, _060000_);
  or g_117941_(_059998_, _060000_, _060001_);
  or g_117942_(_059986_, _059988_, _060002_);
  or g_117943_(_059980_, _060002_, _060003_);
  or g_117944_(_060001_, _060003_, _060005_);
  or g_117945_(_059984_, _060005_, _060006_);
  or g_117946_(_059996_, _060006_, _060007_);
  xor g_117947_(out[167], out[663], _060008_);
  and g_117948_(_098184_, out[667], _060009_);
  xor g_117949_(out[174], out[670], _060010_);
  xor g_117950_(out[168], out[664], _060011_);
  xor g_117951_(out[161], out[657], _060012_);
  xor g_117952_(out[173], out[669], _060013_);
  xor g_117953_(out[169], out[665], _060014_);
  xor g_117954_(out[164], out[660], _060016_);
  xor g_117955_(out[162], out[658], _060017_);
  and g_117956_(out[171], _049620_, _060018_);
  xor g_117957_(out[163], out[659], _060019_);
  xor g_117958_(out[166], out[662], _060020_);
  xor g_117959_(out[175], out[671], _060021_);
  xor g_117960_(out[170], out[666], _060022_);
  xor g_117961_(out[165], out[661], _060023_);
  xor g_117962_(out[160], out[656], _060024_);
  or g_117963_(_060010_, _060016_, _060025_);
  or g_117964_(_060011_, _060013_, _060027_);
  or g_117965_(_060017_, _060022_, _060028_);
  or g_117966_(_060027_, _060028_, _060029_);
  or g_117967_(_060014_, _060019_, _060030_);
  or g_117968_(_060023_, _060024_, _060031_);
  or g_117969_(_060030_, _060031_, _060032_);
  or g_117970_(_060029_, _060032_, _060033_);
  xor g_117971_(out[172], out[668], _060034_);
  or g_117972_(_060009_, _060034_, _060035_);
  or g_117973_(_060008_, _060020_, _060036_);
  or g_117974_(_060035_, _060036_, _060038_);
  or g_117975_(_060012_, _060018_, _060039_);
  or g_117976_(_060021_, _060039_, _060040_);
  or g_117977_(_060038_, _060040_, _060041_);
  or g_117978_(_060033_, _060041_, _060042_);
  or g_117979_(_060025_, _060042_, _060043_);
  not g_117980_(_060043_, _060044_);
  xor g_117981_(out[145], out[657], _060045_);
  and g_117982_(out[155], _049620_, _060046_);
  xor g_117983_(out[158], out[670], _060047_);
  xor g_117984_(out[147], out[659], _060049_);
  xor g_117985_(out[148], out[660], _060050_);
  xor g_117986_(out[146], out[658], _060051_);
  xor g_117987_(out[153], out[665], _060052_);
  xor g_117988_(out[144], out[656], _060053_);
  and g_117989_(_098173_, out[667], _060054_);
  xor g_117990_(out[150], out[662], _060055_);
  xor g_117991_(out[154], out[666], _060056_);
  xor g_117992_(out[149], out[661], _060057_);
  xor g_117993_(out[159], out[671], _060058_);
  xor g_117994_(out[157], out[669], _060060_);
  xor g_117995_(out[152], out[664], _060061_);
  or g_117996_(_060047_, _060050_, _060062_);
  or g_117997_(_060060_, _060061_, _060063_);
  or g_117998_(_060051_, _060056_, _060064_);
  or g_117999_(_060063_, _060064_, _060065_);
  or g_118000_(_060049_, _060052_, _060066_);
  or g_118001_(_060053_, _060057_, _060067_);
  or g_118002_(_060066_, _060067_, _060068_);
  or g_118003_(_060065_, _060068_, _060069_);
  xor g_118004_(out[156], out[668], _060071_);
  or g_118005_(_060054_, _060071_, _060072_);
  xor g_118006_(out[151], out[663], _060073_);
  or g_118007_(_060055_, _060073_, _060074_);
  or g_118008_(_060072_, _060074_, _060075_);
  or g_118009_(_060045_, _060046_, _060076_);
  or g_118010_(_060058_, _060076_, _060077_);
  or g_118011_(_060075_, _060077_, _060078_);
  or g_118012_(_060069_, _060078_, _060079_);
  or g_118013_(_060062_, _060079_, _060080_);
  xor g_118014_(out[135], out[663], _060082_);
  and g_118015_(_098162_, out[667], _060083_);
  xor g_118016_(out[142], out[670], _060084_);
  xor g_118017_(out[136], out[664], _060085_);
  xor g_118018_(out[129], out[657], _060086_);
  xor g_118019_(out[141], out[669], _060087_);
  xor g_118020_(out[137], out[665], _060088_);
  xor g_118021_(out[132], out[660], _060089_);
  xor g_118022_(out[130], out[658], _060090_);
  and g_118023_(out[139], _049620_, _060091_);
  xor g_118024_(out[131], out[659], _060093_);
  xor g_118025_(out[134], out[662], _060094_);
  xor g_118026_(out[143], out[671], _060095_);
  xor g_118027_(out[138], out[666], _060096_);
  xor g_118028_(out[133], out[661], _060097_);
  xor g_118029_(out[128], out[656], _060098_);
  or g_118030_(_060084_, _060089_, _060099_);
  or g_118031_(_060085_, _060087_, _060100_);
  or g_118032_(_060090_, _060096_, _060101_);
  or g_118033_(_060100_, _060101_, _060102_);
  or g_118034_(_060088_, _060093_, _060104_);
  or g_118035_(_060097_, _060098_, _060105_);
  or g_118036_(_060104_, _060105_, _060106_);
  or g_118037_(_060102_, _060106_, _060107_);
  xor g_118038_(out[140], out[668], _060108_);
  or g_118039_(_060083_, _060108_, _060109_);
  or g_118040_(_060082_, _060094_, _060110_);
  or g_118041_(_060109_, _060110_, _060111_);
  or g_118042_(_060086_, _060091_, _060112_);
  or g_118043_(_060095_, _060112_, _060113_);
  or g_118044_(_060111_, _060113_, _060115_);
  or g_118045_(_060107_, _060115_, _060116_);
  or g_118046_(_060099_, _060116_, _060117_);
  xor g_118047_(out[113], out[657], _060118_);
  and g_118048_(out[123], _049620_, _060119_);
  xor g_118049_(out[126], out[670], _060120_);
  xor g_118050_(out[115], out[659], _060121_);
  xor g_118051_(out[116], out[660], _060122_);
  xor g_118052_(out[114], out[658], _060123_);
  xor g_118053_(out[121], out[665], _060124_);
  xor g_118054_(out[112], out[656], _060126_);
  and g_118055_(_098151_, out[667], _060127_);
  xor g_118056_(out[118], out[662], _060128_);
  xor g_118057_(out[122], out[666], _060129_);
  xor g_118058_(out[117], out[661], _060130_);
  xor g_118059_(out[127], out[671], _060131_);
  xor g_118060_(out[125], out[669], _060132_);
  xor g_118061_(out[120], out[664], _060133_);
  or g_118062_(_060120_, _060122_, _060134_);
  or g_118063_(_060132_, _060133_, _060135_);
  or g_118064_(_060123_, _060129_, _060137_);
  or g_118065_(_060135_, _060137_, _060138_);
  or g_118066_(_060121_, _060124_, _060139_);
  or g_118067_(_060126_, _060130_, _060140_);
  or g_118068_(_060139_, _060140_, _060141_);
  or g_118069_(_060138_, _060141_, _060142_);
  xor g_118070_(out[124], out[668], _060143_);
  or g_118071_(_060127_, _060143_, _060144_);
  xor g_118072_(out[119], out[663], _060145_);
  or g_118073_(_060128_, _060145_, _060146_);
  or g_118074_(_060144_, _060146_, _060148_);
  or g_118075_(_060118_, _060119_, _060149_);
  or g_118076_(_060131_, _060149_, _060150_);
  or g_118077_(_060148_, _060150_, _060151_);
  or g_118078_(_060142_, _060151_, _060152_);
  or g_118079_(_060134_, _060152_, _060153_);
  xor g_118080_(out[103], out[663], _060154_);
  and g_118081_(_098140_, out[667], _060155_);
  xor g_118082_(out[110], out[670], _060156_);
  xor g_118083_(out[104], out[664], _060157_);
  xor g_118084_(out[97], out[657], _060159_);
  xor g_118085_(out[109], out[669], _060160_);
  xor g_118086_(out[105], out[665], _060161_);
  xor g_118087_(out[100], out[660], _060162_);
  xor g_118088_(out[98], out[658], _060163_);
  and g_118089_(out[107], _049620_, _060164_);
  xor g_118090_(out[99], out[659], _060165_);
  xor g_118091_(out[102], out[662], _060166_);
  xor g_118092_(out[111], out[671], _060167_);
  xor g_118093_(out[106], out[666], _060168_);
  xor g_118094_(out[101], out[661], _060170_);
  xor g_118095_(out[96], out[656], _060171_);
  or g_118096_(_060156_, _060162_, _060172_);
  or g_118097_(_060157_, _060160_, _060173_);
  or g_118098_(_060163_, _060168_, _060174_);
  or g_118099_(_060173_, _060174_, _060175_);
  or g_118100_(_060161_, _060165_, _060176_);
  or g_118101_(_060170_, _060171_, _060177_);
  or g_118102_(_060176_, _060177_, _060178_);
  or g_118103_(_060175_, _060178_, _060179_);
  xor g_118104_(out[108], out[668], _060181_);
  or g_118105_(_060155_, _060181_, _060182_);
  or g_118106_(_060154_, _060166_, _060183_);
  or g_118107_(_060182_, _060183_, _060184_);
  or g_118108_(_060159_, _060164_, _060185_);
  or g_118109_(_060167_, _060185_, _060186_);
  or g_118110_(_060184_, _060186_, _060187_);
  or g_118111_(_060179_, _060187_, _060188_);
  or g_118112_(_060172_, _060188_, _060189_);
  xor g_118113_(out[83], out[659], _060190_);
  xor g_118114_(out[84], out[660], _060192_);
  xor g_118115_(out[94], out[670], _060193_);
  xor g_118116_(out[82], out[658], _060194_);
  xor g_118117_(out[85], out[661], _060195_);
  xor g_118118_(out[89], out[665], _060196_);
  xor g_118119_(out[88], out[664], _060197_);
  xor g_118120_(out[95], out[671], _060198_);
  xor g_118121_(out[90], out[666], _060199_);
  xor g_118122_(out[86], out[662], _060200_);
  xor g_118123_(out[80], out[656], _060201_);
  and g_118124_(_098129_, out[667], _060203_);
  and g_118125_(out[91], _049620_, _060204_);
  xor g_118126_(out[93], out[669], _060205_);
  or g_118127_(_060197_, _060205_, _060206_);
  xor g_118128_(out[81], out[657], _060207_);
  or g_118129_(_060194_, _060199_, _060208_);
  or g_118130_(_060206_, _060208_, _060209_);
  or g_118131_(_060190_, _060196_, _060210_);
  or g_118132_(_060195_, _060210_, _060211_);
  or g_118133_(_060209_, _060211_, _060212_);
  or g_118134_(_060192_, _060193_, _060214_);
  or g_118135_(_060212_, _060214_, _060215_);
  xor g_118136_(out[92], out[668], _060216_);
  or g_118137_(_060203_, _060216_, _060217_);
  xor g_118138_(out[87], out[663], _060218_);
  or g_118139_(_060200_, _060218_, _060219_);
  or g_118140_(_060217_, _060219_, _060220_);
  or g_118141_(_060204_, _060207_, _060221_);
  or g_118142_(_060198_, _060221_, _060222_);
  or g_118143_(_060220_, _060222_, _060223_);
  or g_118144_(_060201_, _060223_, _060225_);
  or g_118145_(_060215_, _060225_, _060226_);
  not g_118146_(_060226_, _060227_);
  xor g_118147_(out[71], out[663], _060228_);
  and g_118148_(_098118_, out[667], _060229_);
  xor g_118149_(out[78], out[670], _060230_);
  xor g_118150_(out[72], out[664], _060231_);
  xor g_118151_(out[65], out[657], _060232_);
  xor g_118152_(out[77], out[669], _060233_);
  xor g_118153_(out[73], out[665], _060234_);
  xor g_118154_(out[68], out[660], _060236_);
  xor g_118155_(out[66], out[658], _060237_);
  and g_118156_(out[75], _049620_, _060238_);
  xor g_118157_(out[67], out[659], _060239_);
  xor g_118158_(out[70], out[662], _060240_);
  xor g_118159_(out[79], out[671], _060241_);
  xor g_118160_(out[74], out[666], _060242_);
  xor g_118161_(out[69], out[661], _060243_);
  xor g_118162_(out[64], out[656], _060244_);
  or g_118163_(_060230_, _060236_, _060245_);
  or g_118164_(_060231_, _060233_, _060247_);
  or g_118165_(_060237_, _060242_, _060248_);
  or g_118166_(_060247_, _060248_, _060249_);
  or g_118167_(_060234_, _060239_, _060250_);
  or g_118168_(_060243_, _060244_, _060251_);
  or g_118169_(_060250_, _060251_, _060252_);
  or g_118170_(_060249_, _060252_, _060253_);
  xor g_118171_(out[76], out[668], _060254_);
  or g_118172_(_060229_, _060254_, _060255_);
  or g_118173_(_060228_, _060240_, _060256_);
  or g_118174_(_060255_, _060256_, _060258_);
  or g_118175_(_060232_, _060238_, _060259_);
  or g_118176_(_060241_, _060259_, _060260_);
  or g_118177_(_060258_, _060260_, _060261_);
  or g_118178_(_060253_, _060261_, _060262_);
  or g_118179_(_060245_, _060262_, _060263_);
  xor g_118180_(out[60], out[668], _060264_);
  and g_118181_(_098107_, out[667], _060265_);
  xor g_118182_(out[56], out[664], _060266_);
  xor g_118183_(out[54], out[662], _060267_);
  xor g_118184_(out[61], out[669], _060269_);
  xor g_118185_(out[62], out[670], _060270_);
  xor g_118186_(out[50], out[658], _060271_);
  xor g_118187_(out[57], out[665], _060272_);
  xor g_118188_(out[53], out[661], _060273_);
  xor g_118189_(out[49], out[657], _060274_);
  and g_118190_(out[59], _049620_, _060275_);
  or g_118191_(_060266_, _060269_, _060276_);
  xor g_118192_(out[63], out[671], _060277_);
  xor g_118193_(out[58], out[666], _060278_);
  xor g_118194_(out[52], out[660], _060280_);
  xor g_118195_(out[51], out[659], _060281_);
  xor g_118196_(out[48], out[656], _060282_);
  or g_118197_(_060271_, _060278_, _060283_);
  or g_118198_(_060276_, _060283_, _060284_);
  or g_118199_(_060272_, _060281_, _060285_);
  or g_118200_(_060273_, _060285_, _060286_);
  or g_118201_(_060284_, _060286_, _060287_);
  or g_118202_(_060270_, _060280_, _060288_);
  or g_118203_(_060287_, _060288_, _060289_);
  or g_118204_(_060264_, _060265_, _060291_);
  xor g_118205_(out[55], out[663], _060292_);
  or g_118206_(_060267_, _060292_, _060293_);
  or g_118207_(_060291_, _060293_, _060294_);
  or g_118208_(_060274_, _060275_, _060295_);
  or g_118209_(_060277_, _060295_, _060296_);
  or g_118210_(_060294_, _060296_, _060297_);
  or g_118211_(_060282_, _060297_, _060298_);
  or g_118212_(_060289_, _060298_, _060299_);
  xor g_118213_(out[39], out[663], _060300_);
  and g_118214_(_098096_, out[667], _060302_);
  xor g_118215_(out[46], out[670], _060303_);
  xor g_118216_(out[40], out[664], _060304_);
  xor g_118217_(out[33], out[657], _060305_);
  xor g_118218_(out[45], out[669], _060306_);
  xor g_118219_(out[41], out[665], _060307_);
  xor g_118220_(out[36], out[660], _060308_);
  xor g_118221_(out[34], out[658], _060309_);
  and g_118222_(out[43], _049620_, _060310_);
  xor g_118223_(out[35], out[659], _060311_);
  xor g_118224_(out[38], out[662], _060313_);
  xor g_118225_(out[47], out[671], _060314_);
  xor g_118226_(out[42], out[666], _060315_);
  xor g_118227_(out[37], out[661], _060316_);
  xor g_118228_(out[32], out[656], _060317_);
  or g_118229_(_060303_, _060308_, _060318_);
  or g_118230_(_060304_, _060306_, _060319_);
  or g_118231_(_060309_, _060315_, _060320_);
  or g_118232_(_060319_, _060320_, _060321_);
  or g_118233_(_060307_, _060311_, _060322_);
  or g_118234_(_060316_, _060317_, _060324_);
  or g_118235_(_060322_, _060324_, _060325_);
  or g_118236_(_060321_, _060325_, _060326_);
  xor g_118237_(out[44], out[668], _060327_);
  or g_118238_(_060302_, _060327_, _060328_);
  or g_118239_(_060300_, _060313_, _060329_);
  or g_118240_(_060328_, _060329_, _060330_);
  or g_118241_(_060305_, _060310_, _060331_);
  or g_118242_(_060314_, _060331_, _060332_);
  or g_118243_(_060330_, _060332_, _060333_);
  or g_118244_(_060326_, _060333_, _060335_);
  or g_118245_(_060318_, _060335_, _060336_);
  not g_118246_(_060336_, _060337_);
  xor g_118247_(out[24], out[664], _060338_);
  xor g_118248_(out[21], out[661], _060339_);
  xor g_118249_(out[19], out[659], _060340_);
  xor g_118250_(out[30], out[670], _060341_);
  xor g_118251_(out[29], out[669], _060342_);
  xor g_118252_(out[18], out[658], _060343_);
  xor g_118253_(out[25], out[665], _060344_);
  xor g_118254_(out[22], out[662], _060346_);
  xor g_118255_(out[31], out[671], _060347_);
  xor g_118256_(out[26], out[666], _060348_);
  xor g_118257_(out[20], out[660], _060349_);
  xor g_118258_(out[16], out[656], _060350_);
  and g_118259_(_098063_, out[667], _060351_);
  and g_118260_(out[27], _049620_, _060352_);
  or g_118261_(_060338_, _060342_, _060353_);
  xor g_118262_(out[17], out[657], _060354_);
  or g_118263_(_060343_, _060348_, _060355_);
  or g_118264_(_060353_, _060355_, _060357_);
  or g_118265_(_060340_, _060344_, _060358_);
  or g_118266_(_060339_, _060358_, _060359_);
  or g_118267_(_060357_, _060359_, _060360_);
  or g_118268_(_060341_, _060349_, _060361_);
  or g_118269_(_060360_, _060361_, _060362_);
  xor g_118270_(out[28], out[668], _060363_);
  or g_118271_(_060351_, _060363_, _060364_);
  xor g_118272_(out[23], out[663], _060365_);
  or g_118273_(_060346_, _060365_, _060366_);
  or g_118274_(_060364_, _060366_, _060368_);
  or g_118275_(_060352_, _060354_, _060369_);
  or g_118276_(_060347_, _060369_, _060370_);
  or g_118277_(_060368_, _060370_, _060371_);
  or g_118278_(_060350_, _060371_, _060372_);
  or g_118279_(_060362_, _060372_, _060373_);
  not g_118280_(_060373_, _060374_);
  and g_118281_(out[11], _049620_, _060375_);
  and g_118282_(_098041_, out[667], _060376_);
  xor g_118283_(out[13], out[669], _060377_);
  xor g_118284_(out[15], out[671], _060379_);
  xor g_118285_(out[1], out[657], _060380_);
  xor g_118286_(out[4], out[660], _060381_);
  xor g_118287_(out[14], out[670], _060382_);
  or g_118288_(_060381_, _060382_, _060383_);
  xor g_118289_(out[8], out[664], _060384_);
  xor g_118290_(out[0], out[656], _060385_);
  xor g_118291_(out[2], out[658], _060386_);
  xor g_118292_(out[9], out[665], _060387_);
  xor g_118293_(out[5], out[661], _060388_);
  xor g_118294_(out[3], out[659], _060390_);
  xor g_118295_(out[10], out[666], _060391_);
  xor g_118296_(out[6], out[662], _060392_);
  or g_118297_(_060377_, _060384_, _060393_);
  or g_118298_(_060386_, _060391_, _060394_);
  or g_118299_(_060393_, _060394_, _060395_);
  or g_118300_(_060387_, _060390_, _060396_);
  or g_118301_(_060385_, _060388_, _060397_);
  or g_118302_(_060396_, _060397_, _060398_);
  or g_118303_(_060395_, _060398_, _060399_);
  xor g_118304_(out[12], out[668], _060401_);
  or g_118305_(_060376_, _060401_, _060402_);
  xor g_118306_(out[7], out[663], _060403_);
  or g_118307_(_060392_, _060403_, _060404_);
  or g_118308_(_060402_, _060404_, _060405_);
  or g_118309_(_060375_, _060380_, _060406_);
  or g_118310_(_060379_, _060406_, _060407_);
  or g_118311_(_060405_, _060407_, _060408_);
  or g_118312_(_060399_, _060408_, _060409_);
  or g_118313_(_060383_, _060409_, _060410_);
  not g_118314_(_060410_, _060412_);
  xor g_118315_(out[471], out[647], _060413_);
  and g_118316_(_049499_, out[651], _060414_);
  xor g_118317_(out[478], out[654], _060415_);
  xor g_118318_(out[472], out[648], _060416_);
  xor g_118319_(out[465], out[641], _060417_);
  xor g_118320_(out[477], out[653], _060418_);
  xor g_118321_(out[473], out[649], _060419_);
  xor g_118322_(out[468], out[644], _060420_);
  xor g_118323_(out[466], out[642], _060421_);
  and g_118324_(out[475], _049609_, _060423_);
  xor g_118325_(out[467], out[643], _060424_);
  xor g_118326_(out[470], out[646], _060425_);
  xor g_118327_(out[479], out[655], _060426_);
  xor g_118328_(out[474], out[650], _060427_);
  xor g_118329_(out[469], out[645], _060428_);
  xor g_118330_(out[464], out[640], _060429_);
  or g_118331_(_060415_, _060420_, _060430_);
  or g_118332_(_060416_, _060418_, _060431_);
  or g_118333_(_060421_, _060427_, _060432_);
  or g_118334_(_060431_, _060432_, _060434_);
  or g_118335_(_060419_, _060424_, _060435_);
  or g_118336_(_060428_, _060429_, _060436_);
  or g_118337_(_060435_, _060436_, _060437_);
  or g_118338_(_060434_, _060437_, _060438_);
  xor g_118339_(out[476], out[652], _060439_);
  or g_118340_(_060414_, _060439_, _060440_);
  or g_118341_(_060413_, _060425_, _060441_);
  or g_118342_(_060440_, _060441_, _060442_);
  or g_118343_(_060417_, _060423_, _060443_);
  or g_118344_(_060426_, _060443_, _060445_);
  or g_118345_(_060442_, _060445_, _060446_);
  or g_118346_(_060438_, _060446_, _060447_);
  or g_118347_(_060430_, _060447_, _060448_);
  xor g_118348_(out[460], out[652], _060449_);
  and g_118349_(_049477_, out[651], _060450_);
  xor g_118350_(out[456], out[648], _060451_);
  xor g_118351_(out[454], out[646], _060452_);
  xor g_118352_(out[461], out[653], _060453_);
  xor g_118353_(out[462], out[654], _060454_);
  xor g_118354_(out[450], out[642], _060456_);
  xor g_118355_(out[457], out[649], _060457_);
  xor g_118356_(out[453], out[645], _060458_);
  xor g_118357_(out[449], out[641], _060459_);
  and g_118358_(out[459], _049609_, _060460_);
  or g_118359_(_060451_, _060453_, _060461_);
  xor g_118360_(out[463], out[655], _060462_);
  xor g_118361_(out[458], out[650], _060463_);
  xor g_118362_(out[452], out[644], _060464_);
  xor g_118363_(out[451], out[643], _060465_);
  xor g_118364_(out[448], out[640], _060467_);
  or g_118365_(_060456_, _060463_, _060468_);
  or g_118366_(_060461_, _060468_, _060469_);
  or g_118367_(_060457_, _060465_, _060470_);
  or g_118368_(_060458_, _060470_, _060471_);
  or g_118369_(_060469_, _060471_, _060472_);
  or g_118370_(_060454_, _060464_, _060473_);
  or g_118371_(_060472_, _060473_, _060474_);
  or g_118372_(_060449_, _060450_, _060475_);
  xor g_118373_(out[455], out[647], _060476_);
  or g_118374_(_060452_, _060476_, _060478_);
  or g_118375_(_060475_, _060478_, _060479_);
  or g_118376_(_060459_, _060460_, _060480_);
  or g_118377_(_060462_, _060480_, _060481_);
  or g_118378_(_060479_, _060481_, _060482_);
  or g_118379_(_060467_, _060482_, _060483_);
  or g_118380_(_060474_, _060483_, _060484_);
  xor g_118381_(out[439], out[647], _060485_);
  and g_118382_(_049466_, out[651], _060486_);
  xor g_118383_(out[446], out[654], _060487_);
  xor g_118384_(out[440], out[648], _060489_);
  xor g_118385_(out[433], out[641], _060490_);
  xor g_118386_(out[445], out[653], _060491_);
  xor g_118387_(out[441], out[649], _060492_);
  xor g_118388_(out[436], out[644], _060493_);
  xor g_118389_(out[434], out[642], _060494_);
  and g_118390_(out[443], _049609_, _060495_);
  xor g_118391_(out[435], out[643], _060496_);
  xor g_118392_(out[438], out[646], _060497_);
  xor g_118393_(out[447], out[655], _060498_);
  xor g_118394_(out[442], out[650], _060500_);
  xor g_118395_(out[437], out[645], _060501_);
  xor g_118396_(out[432], out[640], _060502_);
  or g_118397_(_060487_, _060493_, _060503_);
  or g_118398_(_060489_, _060491_, _060504_);
  or g_118399_(_060494_, _060500_, _060505_);
  or g_118400_(_060504_, _060505_, _060506_);
  or g_118401_(_060492_, _060496_, _060507_);
  or g_118402_(_060501_, _060502_, _060508_);
  or g_118403_(_060507_, _060508_, _060509_);
  or g_118404_(_060506_, _060509_, _060511_);
  xor g_118405_(out[444], out[652], _060512_);
  or g_118406_(_060486_, _060512_, _060513_);
  or g_118407_(_060485_, _060497_, _060514_);
  or g_118408_(_060513_, _060514_, _060515_);
  or g_118409_(_060490_, _060495_, _060516_);
  or g_118410_(_060498_, _060516_, _060517_);
  or g_118411_(_060515_, _060517_, _060518_);
  or g_118412_(_060511_, _060518_, _060519_);
  or g_118413_(_060503_, _060519_, _060520_);
  not g_118414_(_060520_, _060522_);
  xor g_118415_(out[417], out[641], _060523_);
  and g_118416_(out[427], _049609_, _060524_);
  xor g_118417_(out[425], out[649], _060525_);
  xor g_118418_(out[416], out[640], _060526_);
  xor g_118419_(out[430], out[654], _060527_);
  xor g_118420_(out[420], out[644], _060528_);
  or g_118421_(_060527_, _060528_, _060529_);
  xor g_118422_(out[429], out[653], _060530_);
  xor g_118423_(out[419], out[643], _060531_);
  and g_118424_(_049455_, out[651], _060533_);
  xor g_118425_(out[422], out[646], _060534_);
  xor g_118426_(out[426], out[650], _060535_);
  xor g_118427_(out[421], out[645], _060536_);
  xor g_118428_(out[431], out[655], _060537_);
  xor g_118429_(out[424], out[648], _060538_);
  or g_118430_(_060530_, _060538_, _060539_);
  xor g_118431_(out[418], out[642], _060540_);
  or g_118432_(_060535_, _060540_, _060541_);
  or g_118433_(_060539_, _060541_, _060542_);
  or g_118434_(_060525_, _060531_, _060544_);
  or g_118435_(_060536_, _060544_, _060545_);
  or g_118436_(_060542_, _060545_, _060546_);
  or g_118437_(_060529_, _060546_, _060547_);
  xor g_118438_(out[428], out[652], _060548_);
  or g_118439_(_060533_, _060548_, _060549_);
  xor g_118440_(out[423], out[647], _060550_);
  or g_118441_(_060534_, _060550_, _060551_);
  or g_118442_(_060549_, _060551_, _060552_);
  or g_118443_(_060523_, _060524_, _060553_);
  or g_118444_(_060537_, _060553_, _060555_);
  or g_118445_(_060552_, _060555_, _060556_);
  or g_118446_(_060526_, _060556_, _060557_);
  or g_118447_(_060547_, _060557_, _060558_);
  xor g_118448_(out[407], out[647], _060559_);
  and g_118449_(_049444_, out[651], _060560_);
  xor g_118450_(out[414], out[654], _060561_);
  xor g_118451_(out[408], out[648], _060562_);
  xor g_118452_(out[401], out[641], _060563_);
  xor g_118453_(out[413], out[653], _060564_);
  xor g_118454_(out[409], out[649], _060566_);
  xor g_118455_(out[404], out[644], _060567_);
  xor g_118456_(out[402], out[642], _060568_);
  and g_118457_(out[411], _049609_, _060569_);
  xor g_118458_(out[403], out[643], _060570_);
  xor g_118459_(out[406], out[646], _060571_);
  xor g_118460_(out[415], out[655], _060572_);
  xor g_118461_(out[410], out[650], _060573_);
  xor g_118462_(out[405], out[645], _060574_);
  xor g_118463_(out[400], out[640], _060575_);
  or g_118464_(_060561_, _060567_, _060577_);
  or g_118465_(_060562_, _060564_, _060578_);
  or g_118466_(_060568_, _060573_, _060579_);
  or g_118467_(_060578_, _060579_, _060580_);
  or g_118468_(_060566_, _060570_, _060581_);
  or g_118469_(_060574_, _060575_, _060582_);
  or g_118470_(_060581_, _060582_, _060583_);
  or g_118471_(_060580_, _060583_, _060584_);
  xor g_118472_(out[412], out[652], _060585_);
  or g_118473_(_060560_, _060585_, _060586_);
  or g_118474_(_060559_, _060571_, _060588_);
  or g_118475_(_060586_, _060588_, _060589_);
  or g_118476_(_060563_, _060569_, _060590_);
  or g_118477_(_060572_, _060590_, _060591_);
  or g_118478_(_060589_, _060591_, _060592_);
  or g_118479_(_060584_, _060592_, _060593_);
  or g_118480_(_060577_, _060593_, _060594_);
  xor g_118481_(out[392], out[648], _060595_);
  xor g_118482_(out[389], out[645], _060596_);
  xor g_118483_(out[387], out[643], _060597_);
  xor g_118484_(out[398], out[654], _060599_);
  xor g_118485_(out[397], out[653], _060600_);
  xor g_118486_(out[386], out[642], _060601_);
  xor g_118487_(out[393], out[649], _060602_);
  xor g_118488_(out[390], out[646], _060603_);
  xor g_118489_(out[399], out[655], _060604_);
  xor g_118490_(out[394], out[650], _060605_);
  xor g_118491_(out[388], out[644], _060606_);
  xor g_118492_(out[384], out[640], _060607_);
  and g_118493_(_049433_, out[651], _060608_);
  and g_118494_(out[395], _049609_, _060610_);
  or g_118495_(_060595_, _060600_, _060611_);
  xor g_118496_(out[385], out[641], _060612_);
  or g_118497_(_060601_, _060605_, _060613_);
  or g_118498_(_060611_, _060613_, _060614_);
  or g_118499_(_060597_, _060602_, _060615_);
  or g_118500_(_060596_, _060615_, _060616_);
  or g_118501_(_060614_, _060616_, _060617_);
  or g_118502_(_060599_, _060606_, _060618_);
  or g_118503_(_060617_, _060618_, _060619_);
  xor g_118504_(out[396], out[652], _060621_);
  or g_118505_(_060608_, _060621_, _060622_);
  xor g_118506_(out[391], out[647], _060623_);
  or g_118507_(_060603_, _060623_, _060624_);
  or g_118508_(_060622_, _060624_, _060625_);
  or g_118509_(_060610_, _060612_, _060626_);
  or g_118510_(_060604_, _060626_, _060627_);
  or g_118511_(_060625_, _060627_, _060628_);
  or g_118512_(_060607_, _060628_, _060629_);
  or g_118513_(_060619_, _060629_, _060630_);
  not g_118514_(_060630_, _060632_);
  xor g_118515_(out[375], out[647], _060633_);
  and g_118516_(_049422_, out[651], _060634_);
  xor g_118517_(out[382], out[654], _060635_);
  xor g_118518_(out[376], out[648], _060636_);
  xor g_118519_(out[369], out[641], _060637_);
  xor g_118520_(out[381], out[653], _060638_);
  xor g_118521_(out[377], out[649], _060639_);
  xor g_118522_(out[372], out[644], _060640_);
  xor g_118523_(out[370], out[642], _060641_);
  and g_118524_(out[379], _049609_, _060643_);
  xor g_118525_(out[371], out[643], _060644_);
  xor g_118526_(out[374], out[646], _060645_);
  xor g_118527_(out[383], out[655], _060646_);
  xor g_118528_(out[378], out[650], _060647_);
  xor g_118529_(out[373], out[645], _060648_);
  xor g_118530_(out[368], out[640], _060649_);
  or g_118531_(_060635_, _060640_, _060650_);
  or g_118532_(_060636_, _060638_, _060651_);
  or g_118533_(_060641_, _060647_, _060652_);
  or g_118534_(_060651_, _060652_, _060654_);
  or g_118535_(_060639_, _060644_, _060655_);
  or g_118536_(_060648_, _060649_, _060656_);
  or g_118537_(_060655_, _060656_, _060657_);
  or g_118538_(_060654_, _060657_, _060658_);
  xor g_118539_(out[380], out[652], _060659_);
  or g_118540_(_060634_, _060659_, _060660_);
  or g_118541_(_060633_, _060645_, _060661_);
  or g_118542_(_060660_, _060661_, _060662_);
  or g_118543_(_060637_, _060643_, _060663_);
  or g_118544_(_060646_, _060663_, _060665_);
  or g_118545_(_060662_, _060665_, _060666_);
  or g_118546_(_060658_, _060666_, _060667_);
  or g_118547_(_060650_, _060667_, _060668_);
  xor g_118548_(out[353], out[641], _060669_);
  and g_118549_(out[363], _049609_, _060670_);
  xor g_118550_(out[361], out[649], _060671_);
  xor g_118551_(out[352], out[640], _060672_);
  xor g_118552_(out[366], out[654], _060673_);
  xor g_118553_(out[356], out[644], _060674_);
  or g_118554_(_060673_, _060674_, _060676_);
  xor g_118555_(out[365], out[653], _060677_);
  xor g_118556_(out[355], out[643], _060678_);
  and g_118557_(_049411_, out[651], _060679_);
  xor g_118558_(out[358], out[646], _060680_);
  xor g_118559_(out[362], out[650], _060681_);
  xor g_118560_(out[357], out[645], _060682_);
  xor g_118561_(out[367], out[655], _060683_);
  xor g_118562_(out[360], out[648], _060684_);
  or g_118563_(_060677_, _060684_, _060685_);
  xor g_118564_(out[354], out[642], _060687_);
  or g_118565_(_060681_, _060687_, _060688_);
  or g_118566_(_060685_, _060688_, _060689_);
  or g_118567_(_060671_, _060678_, _060690_);
  or g_118568_(_060682_, _060690_, _060691_);
  or g_118569_(_060689_, _060691_, _060692_);
  or g_118570_(_060676_, _060692_, _060693_);
  xor g_118571_(out[364], out[652], _060694_);
  or g_118572_(_060679_, _060694_, _060695_);
  xor g_118573_(out[359], out[647], _060696_);
  or g_118574_(_060680_, _060696_, _060698_);
  or g_118575_(_060695_, _060698_, _060699_);
  or g_118576_(_060669_, _060670_, _060700_);
  or g_118577_(_060683_, _060700_, _060701_);
  or g_118578_(_060699_, _060701_, _060702_);
  or g_118579_(_060672_, _060702_, _060703_);
  or g_118580_(_060693_, _060703_, _060704_);
  xor g_118581_(out[343], out[647], _060705_);
  and g_118582_(_049400_, out[651], _060706_);
  xor g_118583_(out[350], out[654], _060707_);
  xor g_118584_(out[344], out[648], _060709_);
  xor g_118585_(out[337], out[641], _060710_);
  xor g_118586_(out[349], out[653], _060711_);
  xor g_118587_(out[345], out[649], _060712_);
  xor g_118588_(out[340], out[644], _060713_);
  xor g_118589_(out[338], out[642], _060714_);
  and g_118590_(out[347], _049609_, _060715_);
  xor g_118591_(out[339], out[643], _060716_);
  xor g_118592_(out[342], out[646], _060717_);
  xor g_118593_(out[351], out[655], _060718_);
  xor g_118594_(out[346], out[650], _060720_);
  xor g_118595_(out[341], out[645], _060721_);
  xor g_118596_(out[336], out[640], _060722_);
  or g_118597_(_060707_, _060713_, _060723_);
  or g_118598_(_060709_, _060711_, _060724_);
  or g_118599_(_060714_, _060720_, _060725_);
  or g_118600_(_060724_, _060725_, _060726_);
  or g_118601_(_060712_, _060716_, _060727_);
  or g_118602_(_060721_, _060722_, _060728_);
  or g_118603_(_060727_, _060728_, _060729_);
  or g_118604_(_060726_, _060729_, _060731_);
  xor g_118605_(out[348], out[652], _060732_);
  or g_118606_(_060706_, _060732_, _060733_);
  or g_118607_(_060705_, _060717_, _060734_);
  or g_118608_(_060733_, _060734_, _060735_);
  or g_118609_(_060710_, _060715_, _060736_);
  or g_118610_(_060718_, _060736_, _060737_);
  or g_118611_(_060735_, _060737_, _060738_);
  or g_118612_(_060731_, _060738_, _060739_);
  or g_118613_(_060723_, _060739_, _060740_);
  not g_118614_(_060740_, _060742_);
  xor g_118615_(out[321], out[641], _060743_);
  and g_118616_(out[331], _049609_, _060744_);
  xor g_118617_(out[329], out[649], _060745_);
  xor g_118618_(out[320], out[640], _060746_);
  xor g_118619_(out[334], out[654], _060747_);
  xor g_118620_(out[324], out[644], _060748_);
  or g_118621_(_060747_, _060748_, _060749_);
  xor g_118622_(out[333], out[653], _060750_);
  xor g_118623_(out[323], out[643], _060751_);
  and g_118624_(_098294_, out[651], _060753_);
  xor g_118625_(out[326], out[646], _060754_);
  xor g_118626_(out[330], out[650], _060755_);
  xor g_118627_(out[325], out[645], _060756_);
  xor g_118628_(out[335], out[655], _060757_);
  xor g_118629_(out[328], out[648], _060758_);
  or g_118630_(_060750_, _060758_, _060759_);
  xor g_118631_(out[322], out[642], _060760_);
  or g_118632_(_060755_, _060760_, _060761_);
  or g_118633_(_060759_, _060761_, _060762_);
  or g_118634_(_060745_, _060751_, _060764_);
  or g_118635_(_060756_, _060764_, _060765_);
  or g_118636_(_060762_, _060765_, _060766_);
  or g_118637_(_060749_, _060766_, _060767_);
  xor g_118638_(out[332], out[652], _060768_);
  or g_118639_(_060753_, _060768_, _060769_);
  xor g_118640_(out[327], out[647], _060770_);
  or g_118641_(_060754_, _060770_, _060771_);
  or g_118642_(_060769_, _060771_, _060772_);
  or g_118643_(_060743_, _060744_, _060773_);
  or g_118644_(_060757_, _060773_, _060775_);
  or g_118645_(_060772_, _060775_, _060776_);
  or g_118646_(_060746_, _060776_, _060777_);
  or g_118647_(_060767_, _060777_, _060778_);
  xor g_118648_(out[311], out[647], _060779_);
  and g_118649_(_098283_, out[651], _060780_);
  xor g_118650_(out[318], out[654], _060781_);
  xor g_118651_(out[312], out[648], _060782_);
  xor g_118652_(out[305], out[641], _060783_);
  xor g_118653_(out[317], out[653], _060784_);
  xor g_118654_(out[313], out[649], _060786_);
  xor g_118655_(out[308], out[644], _060787_);
  xor g_118656_(out[306], out[642], _060788_);
  and g_118657_(out[315], _049609_, _060789_);
  xor g_118658_(out[307], out[643], _060790_);
  xor g_118659_(out[310], out[646], _060791_);
  xor g_118660_(out[319], out[655], _060792_);
  xor g_118661_(out[314], out[650], _060793_);
  xor g_118662_(out[309], out[645], _060794_);
  xor g_118663_(out[304], out[640], _060795_);
  or g_118664_(_060781_, _060787_, _060797_);
  or g_118665_(_060782_, _060784_, _060798_);
  or g_118666_(_060788_, _060793_, _060799_);
  or g_118667_(_060798_, _060799_, _060800_);
  or g_118668_(_060786_, _060790_, _060801_);
  or g_118669_(_060794_, _060795_, _060802_);
  or g_118670_(_060801_, _060802_, _060803_);
  or g_118671_(_060800_, _060803_, _060804_);
  xor g_118672_(out[316], out[652], _060805_);
  or g_118673_(_060780_, _060805_, _060806_);
  or g_118674_(_060779_, _060791_, _060808_);
  or g_118675_(_060806_, _060808_, _060809_);
  or g_118676_(_060783_, _060789_, _060810_);
  or g_118677_(_060792_, _060810_, _060811_);
  or g_118678_(_060809_, _060811_, _060812_);
  or g_118679_(_060804_, _060812_, _060813_);
  or g_118680_(_060797_, _060813_, _060814_);
  xor g_118681_(out[289], out[641], _060815_);
  and g_118682_(out[299], _049609_, _060816_);
  xor g_118683_(out[297], out[649], _060817_);
  xor g_118684_(out[288], out[640], _060819_);
  xor g_118685_(out[302], out[654], _060820_);
  xor g_118686_(out[292], out[644], _060821_);
  or g_118687_(_060820_, _060821_, _060822_);
  xor g_118688_(out[301], out[653], _060823_);
  xor g_118689_(out[291], out[643], _060824_);
  and g_118690_(_098272_, out[651], _060825_);
  xor g_118691_(out[294], out[646], _060826_);
  xor g_118692_(out[298], out[650], _060827_);
  xor g_118693_(out[293], out[645], _060828_);
  xor g_118694_(out[303], out[655], _060830_);
  xor g_118695_(out[296], out[648], _060831_);
  or g_118696_(_060823_, _060831_, _060832_);
  xor g_118697_(out[290], out[642], _060833_);
  or g_118698_(_060827_, _060833_, _060834_);
  or g_118699_(_060832_, _060834_, _060835_);
  or g_118700_(_060817_, _060824_, _060836_);
  or g_118701_(_060828_, _060836_, _060837_);
  or g_118702_(_060835_, _060837_, _060838_);
  or g_118703_(_060822_, _060838_, _060839_);
  xor g_118704_(out[300], out[652], _060841_);
  or g_118705_(_060825_, _060841_, _060842_);
  xor g_118706_(out[295], out[647], _060843_);
  or g_118707_(_060826_, _060843_, _060844_);
  or g_118708_(_060842_, _060844_, _060845_);
  or g_118709_(_060815_, _060816_, _060846_);
  or g_118710_(_060830_, _060846_, _060847_);
  or g_118711_(_060845_, _060847_, _060848_);
  or g_118712_(_060819_, _060848_, _060849_);
  or g_118713_(_060839_, _060849_, _060850_);
  xor g_118714_(out[279], out[647], _060852_);
  and g_118715_(_098261_, out[651], _060853_);
  xor g_118716_(out[286], out[654], _060854_);
  xor g_118717_(out[280], out[648], _060855_);
  xor g_118718_(out[273], out[641], _060856_);
  xor g_118719_(out[285], out[653], _060857_);
  xor g_118720_(out[281], out[649], _060858_);
  xor g_118721_(out[276], out[644], _060859_);
  xor g_118722_(out[274], out[642], _060860_);
  and g_118723_(out[283], _049609_, _060861_);
  xor g_118724_(out[275], out[643], _060863_);
  xor g_118725_(out[278], out[646], _060864_);
  xor g_118726_(out[287], out[655], _060865_);
  xor g_118727_(out[282], out[650], _060866_);
  xor g_118728_(out[277], out[645], _060867_);
  xor g_118729_(out[272], out[640], _060868_);
  or g_118730_(_060854_, _060859_, _060869_);
  or g_118731_(_060855_, _060857_, _060870_);
  or g_118732_(_060860_, _060866_, _060871_);
  or g_118733_(_060870_, _060871_, _060872_);
  or g_118734_(_060858_, _060863_, _060874_);
  or g_118735_(_060867_, _060868_, _060875_);
  or g_118736_(_060874_, _060875_, _060876_);
  or g_118737_(_060872_, _060876_, _060877_);
  xor g_118738_(out[284], out[652], _060878_);
  or g_118739_(_060853_, _060878_, _060879_);
  or g_118740_(_060852_, _060864_, _060880_);
  or g_118741_(_060879_, _060880_, _060881_);
  or g_118742_(_060856_, _060861_, _060882_);
  or g_118743_(_060865_, _060882_, _060883_);
  or g_118744_(_060881_, _060883_, _060885_);
  or g_118745_(_060877_, _060885_, _060886_);
  or g_118746_(_060869_, _060886_, _060887_);
  and g_118747_(out[267], _049609_, _060888_);
  xor g_118748_(out[260], out[644], _060889_);
  xor g_118749_(out[270], out[654], _060890_);
  or g_118750_(_060889_, _060890_, _060891_);
  xor g_118751_(out[269], out[653], _060892_);
  xor g_118752_(out[259], out[643], _060893_);
  xor g_118753_(out[256], out[640], _060894_);
  and g_118754_(_098250_, out[651], _060896_);
  xor g_118755_(out[266], out[650], _060897_);
  xor g_118756_(out[271], out[655], _060898_);
  xor g_118757_(out[262], out[646], _060899_);
  xor g_118758_(out[261], out[645], _060900_);
  xor g_118759_(out[264], out[648], _060901_);
  or g_118760_(_060892_, _060901_, _060902_);
  xor g_118761_(out[258], out[642], _060903_);
  xor g_118762_(out[265], out[649], _060904_);
  xor g_118763_(out[257], out[641], _060905_);
  or g_118764_(_060897_, _060903_, _060907_);
  or g_118765_(_060902_, _060907_, _060908_);
  or g_118766_(_060893_, _060904_, _060909_);
  or g_118767_(_060900_, _060909_, _060910_);
  or g_118768_(_060908_, _060910_, _060911_);
  or g_118769_(_060891_, _060911_, _060912_);
  xor g_118770_(out[268], out[652], _060913_);
  or g_118771_(_060896_, _060913_, _060914_);
  xor g_118772_(out[263], out[647], _060915_);
  or g_118773_(_060899_, _060915_, _060916_);
  or g_118774_(_060914_, _060916_, _060918_);
  or g_118775_(_060888_, _060905_, _060919_);
  or g_118776_(_060898_, _060919_, _060920_);
  or g_118777_(_060918_, _060920_, _060921_);
  or g_118778_(_060894_, _060921_, _060922_);
  or g_118779_(_060912_, _060922_, _060923_);
  xor g_118780_(out[247], out[647], _060924_);
  and g_118781_(_098239_, out[651], _060925_);
  xor g_118782_(out[254], out[654], _060926_);
  xor g_118783_(out[248], out[648], _060927_);
  xor g_118784_(out[241], out[641], _060929_);
  xor g_118785_(out[253], out[653], _060930_);
  xor g_118786_(out[249], out[649], _060931_);
  xor g_118787_(out[244], out[644], _060932_);
  xor g_118788_(out[242], out[642], _060933_);
  and g_118789_(out[251], _049609_, _060934_);
  xor g_118790_(out[243], out[643], _060935_);
  xor g_118791_(out[246], out[646], _060936_);
  xor g_118792_(out[255], out[655], _060937_);
  xor g_118793_(out[250], out[650], _060938_);
  xor g_118794_(out[245], out[645], _060940_);
  xor g_118795_(out[240], out[640], _060941_);
  or g_118796_(_060926_, _060932_, _060942_);
  or g_118797_(_060927_, _060930_, _060943_);
  or g_118798_(_060933_, _060938_, _060944_);
  or g_118799_(_060943_, _060944_, _060945_);
  or g_118800_(_060931_, _060935_, _060946_);
  or g_118801_(_060940_, _060941_, _060947_);
  or g_118802_(_060946_, _060947_, _060948_);
  or g_118803_(_060945_, _060948_, _060949_);
  xor g_118804_(out[252], out[652], _060951_);
  or g_118805_(_060925_, _060951_, _060952_);
  or g_118806_(_060924_, _060936_, _060953_);
  or g_118807_(_060952_, _060953_, _060954_);
  or g_118808_(_060929_, _060934_, _060955_);
  or g_118809_(_060937_, _060955_, _060956_);
  or g_118810_(_060954_, _060956_, _060957_);
  or g_118811_(_060949_, _060957_, _060958_);
  or g_118812_(_060942_, _060958_, _060959_);
  xor g_118813_(out[225], out[641], _060960_);
  and g_118814_(out[235], _049609_, _060962_);
  xor g_118815_(out[233], out[649], _060963_);
  xor g_118816_(out[224], out[640], _060964_);
  xor g_118817_(out[238], out[654], _060965_);
  xor g_118818_(out[228], out[644], _060966_);
  or g_118819_(_060965_, _060966_, _060967_);
  xor g_118820_(out[237], out[653], _060968_);
  xor g_118821_(out[227], out[643], _060969_);
  and g_118822_(_098228_, out[651], _060970_);
  xor g_118823_(out[230], out[646], _060971_);
  xor g_118824_(out[234], out[650], _060973_);
  xor g_118825_(out[229], out[645], _060974_);
  xor g_118826_(out[239], out[655], _060975_);
  xor g_118827_(out[232], out[648], _060976_);
  or g_118828_(_060968_, _060976_, _060977_);
  xor g_118829_(out[226], out[642], _060978_);
  or g_118830_(_060973_, _060978_, _060979_);
  or g_118831_(_060977_, _060979_, _060980_);
  or g_118832_(_060963_, _060969_, _060981_);
  or g_118833_(_060974_, _060981_, _060982_);
  or g_118834_(_060980_, _060982_, _060984_);
  or g_118835_(_060967_, _060984_, _060985_);
  xor g_118836_(out[236], out[652], _060986_);
  or g_118837_(_060970_, _060986_, _060987_);
  xor g_118838_(out[231], out[647], _060988_);
  or g_118839_(_060971_, _060988_, _060989_);
  or g_118840_(_060987_, _060989_, _060990_);
  or g_118841_(_060960_, _060962_, _060991_);
  or g_118842_(_060975_, _060991_, _060992_);
  or g_118843_(_060990_, _060992_, _060993_);
  or g_118844_(_060964_, _060993_, _060995_);
  or g_118845_(_060985_, _060995_, _060996_);
  xor g_118846_(out[215], out[647], _060997_);
  and g_118847_(_098217_, out[651], _060998_);
  xor g_118848_(out[222], out[654], _060999_);
  xor g_118849_(out[216], out[648], _061000_);
  xor g_118850_(out[209], out[641], _061001_);
  xor g_118851_(out[221], out[653], _061002_);
  xor g_118852_(out[217], out[649], _061003_);
  xor g_118853_(out[212], out[644], _061004_);
  xor g_118854_(out[210], out[642], _061006_);
  and g_118855_(out[219], _049609_, _061007_);
  xor g_118856_(out[211], out[643], _061008_);
  xor g_118857_(out[214], out[646], _061009_);
  xor g_118858_(out[223], out[655], _061010_);
  xor g_118859_(out[218], out[650], _061011_);
  xor g_118860_(out[213], out[645], _061012_);
  xor g_118861_(out[208], out[640], _061013_);
  or g_118862_(_060999_, _061004_, _061014_);
  or g_118863_(_061000_, _061002_, _061015_);
  or g_118864_(_061006_, _061011_, _061017_);
  or g_118865_(_061015_, _061017_, _061018_);
  or g_118866_(_061003_, _061008_, _061019_);
  or g_118867_(_061012_, _061013_, _061020_);
  or g_118868_(_061019_, _061020_, _061021_);
  or g_118869_(_061018_, _061021_, _061022_);
  xor g_118870_(out[220], out[652], _061023_);
  or g_118871_(_060998_, _061023_, _061024_);
  or g_118872_(_060997_, _061009_, _061025_);
  or g_118873_(_061024_, _061025_, _061026_);
  or g_118874_(_061001_, _061007_, _061028_);
  or g_118875_(_061010_, _061028_, _061029_);
  or g_118876_(_061026_, _061029_, _061030_);
  or g_118877_(_061022_, _061030_, _061031_);
  or g_118878_(_061014_, _061031_, _061032_);
  xor g_118879_(out[193], out[641], _061033_);
  and g_118880_(out[203], _049609_, _061034_);
  xor g_118881_(out[206], out[654], _061035_);
  xor g_118882_(out[195], out[643], _061036_);
  xor g_118883_(out[196], out[644], _061037_);
  xor g_118884_(out[194], out[642], _061039_);
  xor g_118885_(out[201], out[649], _061040_);
  xor g_118886_(out[192], out[640], _061041_);
  and g_118887_(_098206_, out[651], _061042_);
  xor g_118888_(out[198], out[646], _061043_);
  xor g_118889_(out[202], out[650], _061044_);
  xor g_118890_(out[197], out[645], _061045_);
  xor g_118891_(out[207], out[655], _061046_);
  xor g_118892_(out[205], out[653], _061047_);
  xor g_118893_(out[200], out[648], _061048_);
  or g_118894_(_061035_, _061037_, _061050_);
  or g_118895_(_061047_, _061048_, _061051_);
  or g_118896_(_061039_, _061044_, _061052_);
  or g_118897_(_061051_, _061052_, _061053_);
  or g_118898_(_061036_, _061040_, _061054_);
  or g_118899_(_061041_, _061045_, _061055_);
  or g_118900_(_061054_, _061055_, _061056_);
  or g_118901_(_061053_, _061056_, _061057_);
  xor g_118902_(out[204], out[652], _061058_);
  or g_118903_(_061042_, _061058_, _061059_);
  xor g_118904_(out[199], out[647], _061061_);
  or g_118905_(_061043_, _061061_, _061062_);
  or g_118906_(_061059_, _061062_, _061063_);
  or g_118907_(_061033_, _061034_, _061064_);
  or g_118908_(_061046_, _061064_, _061065_);
  or g_118909_(_061063_, _061065_, _061066_);
  or g_118910_(_061057_, _061066_, _061067_);
  or g_118911_(_061050_, _061067_, _061068_);
  xor g_118912_(out[183], out[647], _061069_);
  and g_118913_(_098195_, out[651], _061070_);
  xor g_118914_(out[190], out[654], _061072_);
  xor g_118915_(out[184], out[648], _061073_);
  xor g_118916_(out[177], out[641], _061074_);
  xor g_118917_(out[189], out[653], _061075_);
  xor g_118918_(out[185], out[649], _061076_);
  xor g_118919_(out[180], out[644], _061077_);
  xor g_118920_(out[178], out[642], _061078_);
  and g_118921_(out[187], _049609_, _061079_);
  xor g_118922_(out[179], out[643], _061080_);
  xor g_118923_(out[182], out[646], _061081_);
  xor g_118924_(out[191], out[655], _061083_);
  xor g_118925_(out[186], out[650], _061084_);
  xor g_118926_(out[181], out[645], _061085_);
  xor g_118927_(out[176], out[640], _061086_);
  or g_118928_(_061072_, _061077_, _061087_);
  or g_118929_(_061073_, _061075_, _061088_);
  or g_118930_(_061078_, _061084_, _061089_);
  or g_118931_(_061088_, _061089_, _061090_);
  or g_118932_(_061076_, _061080_, _061091_);
  or g_118933_(_061085_, _061086_, _061092_);
  or g_118934_(_061091_, _061092_, _061094_);
  or g_118935_(_061090_, _061094_, _061095_);
  xor g_118936_(out[188], out[652], _061096_);
  or g_118937_(_061070_, _061096_, _061097_);
  or g_118938_(_061069_, _061081_, _061098_);
  or g_118939_(_061097_, _061098_, _061099_);
  or g_118940_(_061074_, _061079_, _061100_);
  or g_118941_(_061083_, _061100_, _061101_);
  or g_118942_(_061099_, _061101_, _061102_);
  or g_118943_(_061095_, _061102_, _061103_);
  or g_118944_(_061087_, _061103_, _061105_);
  xor g_118945_(out[172], out[652], _061106_);
  and g_118946_(_098184_, out[651], _061107_);
  xor g_118947_(out[168], out[648], _061108_);
  xor g_118948_(out[166], out[646], _061109_);
  xor g_118949_(out[173], out[653], _061110_);
  xor g_118950_(out[174], out[654], _061111_);
  xor g_118951_(out[162], out[642], _061112_);
  xor g_118952_(out[169], out[649], _061113_);
  xor g_118953_(out[165], out[645], _061114_);
  xor g_118954_(out[161], out[641], _061116_);
  and g_118955_(out[171], _049609_, _061117_);
  or g_118956_(_061108_, _061110_, _061118_);
  xor g_118957_(out[175], out[655], _061119_);
  xor g_118958_(out[170], out[650], _061120_);
  xor g_118959_(out[164], out[644], _061121_);
  xor g_118960_(out[163], out[643], _061122_);
  xor g_118961_(out[160], out[640], _061123_);
  or g_118962_(_061112_, _061120_, _061124_);
  or g_118963_(_061118_, _061124_, _061125_);
  or g_118964_(_061113_, _061122_, _061127_);
  or g_118965_(_061114_, _061127_, _061128_);
  or g_118966_(_061125_, _061128_, _061129_);
  or g_118967_(_061111_, _061121_, _061130_);
  or g_118968_(_061129_, _061130_, _061131_);
  or g_118969_(_061106_, _061107_, _061132_);
  xor g_118970_(out[167], out[647], _061133_);
  or g_118971_(_061109_, _061133_, _061134_);
  or g_118972_(_061132_, _061134_, _061135_);
  or g_118973_(_061116_, _061117_, _061136_);
  or g_118974_(_061119_, _061136_, _061138_);
  or g_118975_(_061135_, _061138_, _061139_);
  or g_118976_(_061123_, _061139_, _061140_);
  or g_118977_(_061131_, _061140_, _061141_);
  not g_118978_(_061141_, _061142_);
  xor g_118979_(out[151], out[647], _061143_);
  and g_118980_(_098173_, out[651], _061144_);
  xor g_118981_(out[158], out[654], _061145_);
  xor g_118982_(out[152], out[648], _061146_);
  xor g_118983_(out[145], out[641], _061147_);
  xor g_118984_(out[157], out[653], _061149_);
  xor g_118985_(out[153], out[649], _061150_);
  xor g_118986_(out[148], out[644], _061151_);
  xor g_118987_(out[146], out[642], _061152_);
  and g_118988_(out[155], _049609_, _061153_);
  xor g_118989_(out[147], out[643], _061154_);
  xor g_118990_(out[150], out[646], _061155_);
  xor g_118991_(out[159], out[655], _061156_);
  xor g_118992_(out[154], out[650], _061157_);
  xor g_118993_(out[149], out[645], _061158_);
  xor g_118994_(out[144], out[640], _061160_);
  or g_118995_(_061145_, _061151_, _061161_);
  or g_118996_(_061146_, _061149_, _061162_);
  or g_118997_(_061152_, _061157_, _061163_);
  or g_118998_(_061162_, _061163_, _061164_);
  or g_118999_(_061150_, _061154_, _061165_);
  or g_119000_(_061158_, _061160_, _061166_);
  or g_119001_(_061165_, _061166_, _061167_);
  or g_119002_(_061164_, _061167_, _061168_);
  xor g_119003_(out[156], out[652], _061169_);
  or g_119004_(_061144_, _061169_, _061171_);
  or g_119005_(_061143_, _061155_, _061172_);
  or g_119006_(_061171_, _061172_, _061173_);
  or g_119007_(_061147_, _061153_, _061174_);
  or g_119008_(_061156_, _061174_, _061175_);
  or g_119009_(_061173_, _061175_, _061176_);
  or g_119010_(_061168_, _061176_, _061177_);
  or g_119011_(_061161_, _061177_, _061178_);
  not g_119012_(_061178_, _061179_);
  and g_119013_(out[139], _049609_, _061180_);
  xor g_119014_(out[132], out[644], _061182_);
  xor g_119015_(out[142], out[654], _061183_);
  or g_119016_(_061182_, _061183_, _061184_);
  xor g_119017_(out[141], out[653], _061185_);
  xor g_119018_(out[131], out[643], _061186_);
  xor g_119019_(out[128], out[640], _061187_);
  and g_119020_(_098162_, out[651], _061188_);
  xor g_119021_(out[138], out[650], _061189_);
  xor g_119022_(out[143], out[655], _061190_);
  xor g_119023_(out[134], out[646], _061191_);
  xor g_119024_(out[133], out[645], _061193_);
  xor g_119025_(out[136], out[648], _061194_);
  or g_119026_(_061185_, _061194_, _061195_);
  xor g_119027_(out[130], out[642], _061196_);
  xor g_119028_(out[137], out[649], _061197_);
  xor g_119029_(out[129], out[641], _061198_);
  or g_119030_(_061189_, _061196_, _061199_);
  or g_119031_(_061195_, _061199_, _061200_);
  or g_119032_(_061186_, _061197_, _061201_);
  or g_119033_(_061193_, _061201_, _061202_);
  or g_119034_(_061200_, _061202_, _061204_);
  or g_119035_(_061184_, _061204_, _061205_);
  xor g_119036_(out[140], out[652], _061206_);
  or g_119037_(_061188_, _061206_, _061207_);
  xor g_119038_(out[135], out[647], _061208_);
  or g_119039_(_061191_, _061208_, _061209_);
  or g_119040_(_061207_, _061209_, _061210_);
  or g_119041_(_061180_, _061198_, _061211_);
  or g_119042_(_061190_, _061211_, _061212_);
  or g_119043_(_061210_, _061212_, _061213_);
  or g_119044_(_061187_, _061213_, _061215_);
  or g_119045_(_061205_, _061215_, _061216_);
  xor g_119046_(out[119], out[647], _061217_);
  and g_119047_(_098151_, out[651], _061218_);
  xor g_119048_(out[126], out[654], _061219_);
  xor g_119049_(out[120], out[648], _061220_);
  xor g_119050_(out[113], out[641], _061221_);
  xor g_119051_(out[125], out[653], _061222_);
  xor g_119052_(out[121], out[649], _061223_);
  xor g_119053_(out[116], out[644], _061224_);
  xor g_119054_(out[114], out[642], _061226_);
  and g_119055_(out[123], _049609_, _061227_);
  xor g_119056_(out[115], out[643], _061228_);
  xor g_119057_(out[118], out[646], _061229_);
  xor g_119058_(out[127], out[655], _061230_);
  xor g_119059_(out[122], out[650], _061231_);
  xor g_119060_(out[117], out[645], _061232_);
  xor g_119061_(out[112], out[640], _061233_);
  or g_119062_(_061219_, _061224_, _061234_);
  or g_119063_(_061220_, _061222_, _061235_);
  or g_119064_(_061226_, _061231_, _061237_);
  or g_119065_(_061235_, _061237_, _061238_);
  or g_119066_(_061223_, _061228_, _061239_);
  or g_119067_(_061232_, _061233_, _061240_);
  or g_119068_(_061239_, _061240_, _061241_);
  or g_119069_(_061238_, _061241_, _061242_);
  xor g_119070_(out[124], out[652], _061243_);
  or g_119071_(_061218_, _061243_, _061244_);
  or g_119072_(_061217_, _061229_, _061245_);
  or g_119073_(_061244_, _061245_, _061246_);
  or g_119074_(_061221_, _061227_, _061248_);
  or g_119075_(_061230_, _061248_, _061249_);
  or g_119076_(_061246_, _061249_, _061250_);
  or g_119077_(_061242_, _061250_, _061251_);
  or g_119078_(_061234_, _061251_, _061252_);
  xor g_119079_(out[97], out[641], _061253_);
  and g_119080_(out[107], _049609_, _061254_);
  xor g_119081_(out[105], out[649], _061255_);
  xor g_119082_(out[96], out[640], _061256_);
  xor g_119083_(out[110], out[654], _061257_);
  xor g_119084_(out[100], out[644], _061259_);
  or g_119085_(_061257_, _061259_, _061260_);
  xor g_119086_(out[109], out[653], _061261_);
  xor g_119087_(out[99], out[643], _061262_);
  and g_119088_(_098140_, out[651], _061263_);
  xor g_119089_(out[102], out[646], _061264_);
  xor g_119090_(out[106], out[650], _061265_);
  xor g_119091_(out[101], out[645], _061266_);
  xor g_119092_(out[111], out[655], _061267_);
  xor g_119093_(out[104], out[648], _061268_);
  or g_119094_(_061261_, _061268_, _061270_);
  xor g_119095_(out[98], out[642], _061271_);
  or g_119096_(_061265_, _061271_, _061272_);
  or g_119097_(_061270_, _061272_, _061273_);
  or g_119098_(_061255_, _061262_, _061274_);
  or g_119099_(_061266_, _061274_, _061275_);
  or g_119100_(_061273_, _061275_, _061276_);
  or g_119101_(_061260_, _061276_, _061277_);
  xor g_119102_(out[108], out[652], _061278_);
  or g_119103_(_061263_, _061278_, _061279_);
  xor g_119104_(out[103], out[647], _061281_);
  or g_119105_(_061264_, _061281_, _061282_);
  or g_119106_(_061279_, _061282_, _061283_);
  or g_119107_(_061253_, _061254_, _061284_);
  or g_119108_(_061267_, _061284_, _061285_);
  or g_119109_(_061283_, _061285_, _061286_);
  or g_119110_(_061256_, _061286_, _061287_);
  or g_119111_(_061277_, _061287_, _061288_);
  xor g_119112_(out[87], out[647], _061289_);
  and g_119113_(_098129_, out[651], _061290_);
  xor g_119114_(out[94], out[654], _061292_);
  xor g_119115_(out[88], out[648], _061293_);
  xor g_119116_(out[81], out[641], _061294_);
  xor g_119117_(out[93], out[653], _061295_);
  xor g_119118_(out[89], out[649], _061296_);
  xor g_119119_(out[84], out[644], _061297_);
  xor g_119120_(out[82], out[642], _061298_);
  and g_119121_(out[91], _049609_, _061299_);
  xor g_119122_(out[83], out[643], _061300_);
  xor g_119123_(out[86], out[646], _061301_);
  xor g_119124_(out[95], out[655], _061303_);
  xor g_119125_(out[90], out[650], _061304_);
  xor g_119126_(out[85], out[645], _061305_);
  xor g_119127_(out[80], out[640], _061306_);
  or g_119128_(_061292_, _061297_, _061307_);
  or g_119129_(_061293_, _061295_, _061308_);
  or g_119130_(_061298_, _061304_, _061309_);
  or g_119131_(_061308_, _061309_, _061310_);
  or g_119132_(_061296_, _061300_, _061311_);
  or g_119133_(_061305_, _061306_, _061312_);
  or g_119134_(_061311_, _061312_, _061314_);
  or g_119135_(_061310_, _061314_, _061315_);
  xor g_119136_(out[92], out[652], _061316_);
  or g_119137_(_061290_, _061316_, _061317_);
  or g_119138_(_061289_, _061301_, _061318_);
  or g_119139_(_061317_, _061318_, _061319_);
  or g_119140_(_061294_, _061299_, _061320_);
  or g_119141_(_061303_, _061320_, _061321_);
  or g_119142_(_061319_, _061321_, _061322_);
  or g_119143_(_061315_, _061322_, _061323_);
  or g_119144_(_061307_, _061323_, _061325_);
  xor g_119145_(out[65], out[641], _061326_);
  and g_119146_(out[75], _049609_, _061327_);
  xor g_119147_(out[73], out[649], _061328_);
  xor g_119148_(out[64], out[640], _061329_);
  xor g_119149_(out[78], out[654], _061330_);
  xor g_119150_(out[68], out[644], _061331_);
  or g_119151_(_061330_, _061331_, _061332_);
  xor g_119152_(out[77], out[653], _061333_);
  xor g_119153_(out[67], out[643], _061334_);
  and g_119154_(_098118_, out[651], _061336_);
  xor g_119155_(out[70], out[646], _061337_);
  xor g_119156_(out[74], out[650], _061338_);
  xor g_119157_(out[69], out[645], _061339_);
  xor g_119158_(out[79], out[655], _061340_);
  xor g_119159_(out[72], out[648], _061341_);
  or g_119160_(_061333_, _061341_, _061342_);
  xor g_119161_(out[66], out[642], _061343_);
  or g_119162_(_061338_, _061343_, _061344_);
  or g_119163_(_061342_, _061344_, _061345_);
  or g_119164_(_061328_, _061334_, _061347_);
  or g_119165_(_061339_, _061347_, _061348_);
  or g_119166_(_061345_, _061348_, _061349_);
  or g_119167_(_061332_, _061349_, _061350_);
  xor g_119168_(out[76], out[652], _061351_);
  or g_119169_(_061336_, _061351_, _061352_);
  xor g_119170_(out[71], out[647], _061353_);
  or g_119171_(_061337_, _061353_, _061354_);
  or g_119172_(_061352_, _061354_, _061355_);
  or g_119173_(_061326_, _061327_, _061356_);
  or g_119174_(_061340_, _061356_, _061358_);
  or g_119175_(_061355_, _061358_, _061359_);
  or g_119176_(_061329_, _061359_, _061360_);
  or g_119177_(_061350_, _061360_, _061361_);
  xor g_119178_(out[55], out[647], _061362_);
  and g_119179_(_098107_, out[651], _061363_);
  xor g_119180_(out[62], out[654], _061364_);
  xor g_119181_(out[56], out[648], _061365_);
  xor g_119182_(out[49], out[641], _061366_);
  xor g_119183_(out[61], out[653], _061367_);
  xor g_119184_(out[57], out[649], _061369_);
  xor g_119185_(out[52], out[644], _061370_);
  xor g_119186_(out[50], out[642], _061371_);
  and g_119187_(out[59], _049609_, _061372_);
  xor g_119188_(out[51], out[643], _061373_);
  xor g_119189_(out[54], out[646], _061374_);
  xor g_119190_(out[63], out[655], _061375_);
  xor g_119191_(out[58], out[650], _061376_);
  xor g_119192_(out[53], out[645], _061377_);
  xor g_119193_(out[48], out[640], _061378_);
  or g_119194_(_061364_, _061370_, _061380_);
  or g_119195_(_061365_, _061367_, _061381_);
  or g_119196_(_061371_, _061376_, _061382_);
  or g_119197_(_061381_, _061382_, _061383_);
  or g_119198_(_061369_, _061373_, _061384_);
  or g_119199_(_061377_, _061378_, _061385_);
  or g_119200_(_061384_, _061385_, _061386_);
  or g_119201_(_061383_, _061386_, _061387_);
  xor g_119202_(out[60], out[652], _061388_);
  or g_119203_(_061363_, _061388_, _061389_);
  or g_119204_(_061362_, _061374_, _061391_);
  or g_119205_(_061389_, _061391_, _061392_);
  or g_119206_(_061366_, _061372_, _061393_);
  or g_119207_(_061375_, _061393_, _061394_);
  or g_119208_(_061392_, _061394_, _061395_);
  or g_119209_(_061387_, _061395_, _061396_);
  or g_119210_(_061380_, _061396_, _061397_);
  xor g_119211_(out[33], out[641], _061398_);
  and g_119212_(out[43], _049609_, _061399_);
  xor g_119213_(out[41], out[649], _061400_);
  xor g_119214_(out[32], out[640], _061402_);
  xor g_119215_(out[46], out[654], _061403_);
  xor g_119216_(out[36], out[644], _061404_);
  or g_119217_(_061403_, _061404_, _061405_);
  xor g_119218_(out[45], out[653], _061406_);
  xor g_119219_(out[35], out[643], _061407_);
  and g_119220_(_098096_, out[651], _061408_);
  xor g_119221_(out[38], out[646], _061409_);
  xor g_119222_(out[42], out[650], _061410_);
  xor g_119223_(out[37], out[645], _061411_);
  xor g_119224_(out[47], out[655], _061413_);
  xor g_119225_(out[40], out[648], _061414_);
  or g_119226_(_061406_, _061414_, _061415_);
  xor g_119227_(out[34], out[642], _061416_);
  or g_119228_(_061410_, _061416_, _061417_);
  or g_119229_(_061415_, _061417_, _061418_);
  or g_119230_(_061400_, _061407_, _061419_);
  or g_119231_(_061411_, _061419_, _061420_);
  or g_119232_(_061418_, _061420_, _061421_);
  or g_119233_(_061405_, _061421_, _061422_);
  xor g_119234_(out[44], out[652], _061424_);
  or g_119235_(_061408_, _061424_, _061425_);
  xor g_119236_(out[39], out[647], _061426_);
  or g_119237_(_061409_, _061426_, _061427_);
  or g_119238_(_061425_, _061427_, _061428_);
  or g_119239_(_061398_, _061399_, _061429_);
  or g_119240_(_061413_, _061429_, _061430_);
  or g_119241_(_061428_, _061430_, _061431_);
  or g_119242_(_061402_, _061431_, _061432_);
  or g_119243_(_061422_, _061432_, _061433_);
  xor g_119244_(out[23], out[647], _061435_);
  and g_119245_(_098063_, out[651], _061436_);
  xor g_119246_(out[30], out[654], _061437_);
  xor g_119247_(out[24], out[648], _061438_);
  xor g_119248_(out[17], out[641], _061439_);
  xor g_119249_(out[29], out[653], _061440_);
  xor g_119250_(out[25], out[649], _061441_);
  xor g_119251_(out[20], out[644], _061442_);
  xor g_119252_(out[18], out[642], _061443_);
  and g_119253_(out[27], _049609_, _061444_);
  xor g_119254_(out[19], out[643], _061446_);
  xor g_119255_(out[22], out[646], _061447_);
  xor g_119256_(out[31], out[655], _061448_);
  xor g_119257_(out[26], out[650], _061449_);
  xor g_119258_(out[21], out[645], _061450_);
  xor g_119259_(out[16], out[640], _061451_);
  or g_119260_(_061437_, _061442_, _061452_);
  or g_119261_(_061438_, _061440_, _061453_);
  or g_119262_(_061443_, _061449_, _061454_);
  or g_119263_(_061453_, _061454_, _061455_);
  or g_119264_(_061441_, _061446_, _061457_);
  or g_119265_(_061450_, _061451_, _061458_);
  or g_119266_(_061457_, _061458_, _061459_);
  or g_119267_(_061455_, _061459_, _061460_);
  xor g_119268_(out[28], out[652], _061461_);
  or g_119269_(_061436_, _061461_, _061462_);
  or g_119270_(_061435_, _061447_, _061463_);
  or g_119271_(_061462_, _061463_, _061464_);
  or g_119272_(_061439_, _061444_, _061465_);
  or g_119273_(_061448_, _061465_, _061466_);
  or g_119274_(_061464_, _061466_, _061468_);
  or g_119275_(_061460_, _061468_, _061469_);
  or g_119276_(_061452_, _061469_, _061470_);
  xor g_119277_(out[1], out[641], _061471_);
  and g_119278_(out[11], _049609_, _061472_);
  xor g_119279_(out[14], out[654], _061473_);
  xor g_119280_(out[3], out[643], _061474_);
  xor g_119281_(out[4], out[644], _061475_);
  xor g_119282_(out[2], out[642], _061476_);
  xor g_119283_(out[9], out[649], _061477_);
  xor g_119284_(out[0], out[640], _061479_);
  and g_119285_(_098041_, out[651], _061480_);
  xor g_119286_(out[6], out[646], _061481_);
  xor g_119287_(out[10], out[650], _061482_);
  xor g_119288_(out[5], out[645], _061483_);
  xor g_119289_(out[15], out[655], _061484_);
  xor g_119290_(out[13], out[653], _061485_);
  xor g_119291_(out[8], out[648], _061486_);
  or g_119292_(_061473_, _061475_, _061487_);
  or g_119293_(_061485_, _061486_, _061488_);
  or g_119294_(_061476_, _061482_, _061490_);
  or g_119295_(_061488_, _061490_, _061491_);
  or g_119296_(_061474_, _061477_, _061492_);
  or g_119297_(_061479_, _061483_, _061493_);
  or g_119298_(_061492_, _061493_, _061494_);
  or g_119299_(_061491_, _061494_, _061495_);
  xor g_119300_(out[12], out[652], _061496_);
  or g_119301_(_061480_, _061496_, _061497_);
  xor g_119302_(out[7], out[647], _061498_);
  or g_119303_(_061481_, _061498_, _061499_);
  or g_119304_(_061497_, _061499_, _061501_);
  or g_119305_(_061471_, _061472_, _061502_);
  or g_119306_(_061484_, _061502_, _061503_);
  or g_119307_(_061501_, _061503_, _061504_);
  or g_119308_(_061495_, _061504_, _061505_);
  or g_119309_(_061487_, _061505_, _061506_);
  xor g_119310_(out[476], out[636], _061507_);
  and g_119311_(_049499_, out[635], _061508_);
  xor g_119312_(out[472], out[632], _061509_);
  xor g_119313_(out[470], out[630], _061510_);
  xor g_119314_(out[477], out[637], _061512_);
  xor g_119315_(out[478], out[638], _061513_);
  xor g_119316_(out[466], out[626], _061514_);
  xor g_119317_(out[473], out[633], _061515_);
  xor g_119318_(out[469], out[629], _061516_);
  xor g_119319_(out[465], out[625], _061517_);
  and g_119320_(out[475], _049598_, _061518_);
  or g_119321_(_061509_, _061512_, _061519_);
  xor g_119322_(out[479], out[639], _061520_);
  xor g_119323_(out[474], out[634], _061521_);
  xor g_119324_(out[468], out[628], _061523_);
  xor g_119325_(out[467], out[627], _061524_);
  xor g_119326_(out[464], out[624], _061525_);
  or g_119327_(_061514_, _061521_, _061526_);
  or g_119328_(_061519_, _061526_, _061527_);
  or g_119329_(_061515_, _061524_, _061528_);
  or g_119330_(_061516_, _061528_, _061529_);
  or g_119331_(_061527_, _061529_, _061530_);
  or g_119332_(_061513_, _061523_, _061531_);
  or g_119333_(_061530_, _061531_, _061532_);
  or g_119334_(_061507_, _061508_, _061534_);
  xor g_119335_(out[471], out[631], _061535_);
  or g_119336_(_061510_, _061535_, _061536_);
  or g_119337_(_061534_, _061536_, _061537_);
  or g_119338_(_061517_, _061518_, _061538_);
  or g_119339_(_061520_, _061538_, _061539_);
  or g_119340_(_061537_, _061539_, _061540_);
  or g_119341_(_061525_, _061540_, _061541_);
  or g_119342_(_061532_, _061541_, _061542_);
  xor g_119343_(out[455], out[631], _061543_);
  and g_119344_(_049477_, out[635], _061545_);
  xor g_119345_(out[462], out[638], _061546_);
  xor g_119346_(out[456], out[632], _061547_);
  xor g_119347_(out[449], out[625], _061548_);
  xor g_119348_(out[461], out[637], _061549_);
  xor g_119349_(out[457], out[633], _061550_);
  xor g_119350_(out[452], out[628], _061551_);
  xor g_119351_(out[450], out[626], _061552_);
  and g_119352_(out[459], _049598_, _061553_);
  xor g_119353_(out[451], out[627], _061554_);
  xor g_119354_(out[454], out[630], _061556_);
  xor g_119355_(out[463], out[639], _061557_);
  xor g_119356_(out[458], out[634], _061558_);
  xor g_119357_(out[453], out[629], _061559_);
  xor g_119358_(out[448], out[624], _061560_);
  or g_119359_(_061546_, _061551_, _061561_);
  or g_119360_(_061547_, _061549_, _061562_);
  or g_119361_(_061552_, _061558_, _061563_);
  or g_119362_(_061562_, _061563_, _061564_);
  or g_119363_(_061550_, _061554_, _061565_);
  or g_119364_(_061559_, _061560_, _061567_);
  or g_119365_(_061565_, _061567_, _061568_);
  or g_119366_(_061564_, _061568_, _061569_);
  xor g_119367_(out[460], out[636], _061570_);
  or g_119368_(_061545_, _061570_, _061571_);
  or g_119369_(_061543_, _061556_, _061572_);
  or g_119370_(_061571_, _061572_, _061573_);
  or g_119371_(_061548_, _061553_, _061574_);
  or g_119372_(_061557_, _061574_, _061575_);
  or g_119373_(_061573_, _061575_, _061576_);
  or g_119374_(_061569_, _061576_, _061578_);
  or g_119375_(_061561_, _061578_, _061579_);
  not g_119376_(_061579_, _061580_);
  xor g_119377_(out[440], out[632], _061581_);
  xor g_119378_(out[437], out[629], _061582_);
  xor g_119379_(out[435], out[627], _061583_);
  xor g_119380_(out[446], out[638], _061584_);
  xor g_119381_(out[445], out[637], _061585_);
  xor g_119382_(out[434], out[626], _061586_);
  xor g_119383_(out[441], out[633], _061587_);
  xor g_119384_(out[438], out[630], _061589_);
  xor g_119385_(out[447], out[639], _061590_);
  xor g_119386_(out[442], out[634], _061591_);
  xor g_119387_(out[436], out[628], _061592_);
  xor g_119388_(out[432], out[624], _061593_);
  and g_119389_(_049466_, out[635], _061594_);
  and g_119390_(out[443], _049598_, _061595_);
  or g_119391_(_061581_, _061585_, _061596_);
  xor g_119392_(out[433], out[625], _061597_);
  or g_119393_(_061586_, _061591_, _061598_);
  or g_119394_(_061596_, _061598_, _061600_);
  or g_119395_(_061583_, _061587_, _061601_);
  or g_119396_(_061582_, _061601_, _061602_);
  or g_119397_(_061600_, _061602_, _061603_);
  or g_119398_(_061584_, _061592_, _061604_);
  or g_119399_(_061603_, _061604_, _061605_);
  xor g_119400_(out[444], out[636], _061606_);
  or g_119401_(_061594_, _061606_, _061607_);
  xor g_119402_(out[439], out[631], _061608_);
  or g_119403_(_061589_, _061608_, _061609_);
  or g_119404_(_061607_, _061609_, _061611_);
  or g_119405_(_061595_, _061597_, _061612_);
  or g_119406_(_061590_, _061612_, _061613_);
  or g_119407_(_061611_, _061613_, _061614_);
  or g_119408_(_061593_, _061614_, _061615_);
  or g_119409_(_061605_, _061615_, _061616_);
  not g_119410_(_061616_, _061617_);
  xor g_119411_(out[423], out[631], _061618_);
  and g_119412_(_049455_, out[635], _061619_);
  xor g_119413_(out[430], out[638], _061620_);
  xor g_119414_(out[424], out[632], _061622_);
  xor g_119415_(out[417], out[625], _061623_);
  xor g_119416_(out[429], out[637], _061624_);
  xor g_119417_(out[425], out[633], _061625_);
  xor g_119418_(out[420], out[628], _061626_);
  xor g_119419_(out[418], out[626], _061627_);
  and g_119420_(out[427], _049598_, _061628_);
  xor g_119421_(out[419], out[627], _061629_);
  xor g_119422_(out[422], out[630], _061630_);
  xor g_119423_(out[431], out[639], _061631_);
  xor g_119424_(out[426], out[634], _061633_);
  xor g_119425_(out[421], out[629], _061634_);
  xor g_119426_(out[416], out[624], _061635_);
  or g_119427_(_061620_, _061626_, _061636_);
  or g_119428_(_061622_, _061624_, _061637_);
  or g_119429_(_061627_, _061633_, _061638_);
  or g_119430_(_061637_, _061638_, _061639_);
  or g_119431_(_061625_, _061629_, _061640_);
  or g_119432_(_061634_, _061635_, _061641_);
  or g_119433_(_061640_, _061641_, _061642_);
  or g_119434_(_061639_, _061642_, _061644_);
  xor g_119435_(out[428], out[636], _061645_);
  or g_119436_(_061619_, _061645_, _061646_);
  or g_119437_(_061618_, _061630_, _061647_);
  or g_119438_(_061646_, _061647_, _061648_);
  or g_119439_(_061623_, _061628_, _061649_);
  or g_119440_(_061631_, _061649_, _061650_);
  or g_119441_(_061648_, _061650_, _061651_);
  or g_119442_(_061644_, _061651_, _061652_);
  or g_119443_(_061636_, _061652_, _061653_);
  xor g_119444_(out[410], out[634], _061655_);
  xor g_119445_(out[402], out[626], _061656_);
  xor g_119446_(out[401], out[625], _061657_);
  and g_119447_(_049444_, out[635], _061658_);
  and g_119448_(out[411], _049598_, _061659_);
  xor g_119449_(out[413], out[637], _061660_);
  xor g_119450_(out[403], out[627], _061661_);
  xor g_119451_(out[414], out[638], _061662_);
  xor g_119452_(out[412], out[636], _061663_);
  xor g_119453_(out[408], out[632], _061664_);
  xor g_119454_(out[415], out[639], _061666_);
  xor g_119455_(out[405], out[629], _061667_);
  xor g_119456_(out[406], out[630], _061668_);
  xor g_119457_(out[400], out[624], _061669_);
  xor g_119458_(out[404], out[628], _061670_);
  or g_119459_(_061660_, _061664_, _061671_);
  xor g_119460_(out[409], out[633], _061672_);
  or g_119461_(_061655_, _061656_, _061673_);
  or g_119462_(_061671_, _061673_, _061674_);
  or g_119463_(_061661_, _061672_, _061675_);
  or g_119464_(_061667_, _061675_, _061677_);
  or g_119465_(_061674_, _061677_, _061678_);
  or g_119466_(_061662_, _061670_, _061679_);
  or g_119467_(_061678_, _061679_, _061680_);
  or g_119468_(_061658_, _061663_, _061681_);
  xor g_119469_(out[407], out[631], _061682_);
  or g_119470_(_061668_, _061682_, _061683_);
  or g_119471_(_061681_, _061683_, _061684_);
  or g_119472_(_061657_, _061659_, _061685_);
  or g_119473_(_061666_, _061685_, _061686_);
  or g_119474_(_061684_, _061686_, _061688_);
  or g_119475_(_061669_, _061688_, _061689_);
  or g_119476_(_061680_, _061689_, _061690_);
  xor g_119477_(out[391], out[631], _061691_);
  and g_119478_(_049433_, out[635], _061692_);
  xor g_119479_(out[398], out[638], _061693_);
  xor g_119480_(out[392], out[632], _061694_);
  xor g_119481_(out[385], out[625], _061695_);
  xor g_119482_(out[397], out[637], _061696_);
  xor g_119483_(out[393], out[633], _061697_);
  xor g_119484_(out[388], out[628], _061699_);
  xor g_119485_(out[386], out[626], _061700_);
  and g_119486_(out[395], _049598_, _061701_);
  xor g_119487_(out[387], out[627], _061702_);
  xor g_119488_(out[390], out[630], _061703_);
  xor g_119489_(out[399], out[639], _061704_);
  xor g_119490_(out[394], out[634], _061705_);
  xor g_119491_(out[389], out[629], _061706_);
  xor g_119492_(out[384], out[624], _061707_);
  or g_119493_(_061693_, _061699_, _061708_);
  or g_119494_(_061694_, _061696_, _061710_);
  or g_119495_(_061700_, _061705_, _061711_);
  or g_119496_(_061710_, _061711_, _061712_);
  or g_119497_(_061697_, _061702_, _061713_);
  or g_119498_(_061706_, _061707_, _061714_);
  or g_119499_(_061713_, _061714_, _061715_);
  or g_119500_(_061712_, _061715_, _061716_);
  xor g_119501_(out[396], out[636], _061717_);
  or g_119502_(_061692_, _061717_, _061718_);
  or g_119503_(_061691_, _061703_, _061719_);
  or g_119504_(_061718_, _061719_, _061721_);
  or g_119505_(_061695_, _061701_, _061722_);
  or g_119506_(_061704_, _061722_, _061723_);
  or g_119507_(_061721_, _061723_, _061724_);
  or g_119508_(_061716_, _061724_, _061725_);
  or g_119509_(_061708_, _061725_, _061726_);
  not g_119510_(_061726_, _061727_);
  xor g_119511_(out[376], out[632], _061728_);
  xor g_119512_(out[373], out[629], _061729_);
  xor g_119513_(out[371], out[627], _061730_);
  xor g_119514_(out[382], out[638], _061732_);
  xor g_119515_(out[381], out[637], _061733_);
  xor g_119516_(out[370], out[626], _061734_);
  xor g_119517_(out[377], out[633], _061735_);
  xor g_119518_(out[374], out[630], _061736_);
  xor g_119519_(out[383], out[639], _061737_);
  xor g_119520_(out[378], out[634], _061738_);
  xor g_119521_(out[372], out[628], _061739_);
  xor g_119522_(out[368], out[624], _061740_);
  and g_119523_(_049422_, out[635], _061741_);
  and g_119524_(out[379], _049598_, _061743_);
  or g_119525_(_061728_, _061733_, _061744_);
  xor g_119526_(out[369], out[625], _061745_);
  or g_119527_(_061734_, _061738_, _061746_);
  or g_119528_(_061744_, _061746_, _061747_);
  or g_119529_(_061730_, _061735_, _061748_);
  or g_119530_(_061729_, _061748_, _061749_);
  or g_119531_(_061747_, _061749_, _061750_);
  or g_119532_(_061732_, _061739_, _061751_);
  or g_119533_(_061750_, _061751_, _061752_);
  xor g_119534_(out[380], out[636], _061754_);
  or g_119535_(_061741_, _061754_, _061755_);
  xor g_119536_(out[375], out[631], _061756_);
  or g_119537_(_061736_, _061756_, _061757_);
  or g_119538_(_061755_, _061757_, _061758_);
  or g_119539_(_061743_, _061745_, _061759_);
  or g_119540_(_061737_, _061759_, _061760_);
  or g_119541_(_061758_, _061760_, _061761_);
  or g_119542_(_061740_, _061761_, _061762_);
  or g_119543_(_061752_, _061762_, _061763_);
  not g_119544_(_061763_, _061765_);
  xor g_119545_(out[359], out[631], _061766_);
  and g_119546_(_049411_, out[635], _061767_);
  xor g_119547_(out[366], out[638], _061768_);
  xor g_119548_(out[360], out[632], _061769_);
  xor g_119549_(out[353], out[625], _061770_);
  xor g_119550_(out[365], out[637], _061771_);
  xor g_119551_(out[361], out[633], _061772_);
  xor g_119552_(out[356], out[628], _061773_);
  xor g_119553_(out[354], out[626], _061774_);
  and g_119554_(out[363], _049598_, _061776_);
  xor g_119555_(out[355], out[627], _061777_);
  xor g_119556_(out[358], out[630], _061778_);
  xor g_119557_(out[367], out[639], _061779_);
  xor g_119558_(out[362], out[634], _061780_);
  xor g_119559_(out[357], out[629], _061781_);
  xor g_119560_(out[352], out[624], _061782_);
  or g_119561_(_061768_, _061773_, _061783_);
  or g_119562_(_061769_, _061771_, _061784_);
  or g_119563_(_061774_, _061780_, _061785_);
  or g_119564_(_061784_, _061785_, _061787_);
  or g_119565_(_061772_, _061777_, _061788_);
  or g_119566_(_061781_, _061782_, _061789_);
  or g_119567_(_061788_, _061789_, _061790_);
  or g_119568_(_061787_, _061790_, _061791_);
  xor g_119569_(out[364], out[636], _061792_);
  or g_119570_(_061767_, _061792_, _061793_);
  or g_119571_(_061766_, _061778_, _061794_);
  or g_119572_(_061793_, _061794_, _061795_);
  or g_119573_(_061770_, _061776_, _061796_);
  or g_119574_(_061779_, _061796_, _061798_);
  or g_119575_(_061795_, _061798_, _061799_);
  or g_119576_(_061791_, _061799_, _061800_);
  or g_119577_(_061783_, _061800_, _061801_);
  xor g_119578_(out[346], out[634], _061802_);
  xor g_119579_(out[338], out[626], _061803_);
  xor g_119580_(out[337], out[625], _061804_);
  and g_119581_(_049400_, out[635], _061805_);
  and g_119582_(out[347], _049598_, _061806_);
  xor g_119583_(out[349], out[637], _061807_);
  xor g_119584_(out[339], out[627], _061809_);
  xor g_119585_(out[350], out[638], _061810_);
  xor g_119586_(out[348], out[636], _061811_);
  xor g_119587_(out[344], out[632], _061812_);
  xor g_119588_(out[351], out[639], _061813_);
  xor g_119589_(out[341], out[629], _061814_);
  xor g_119590_(out[342], out[630], _061815_);
  xor g_119591_(out[336], out[624], _061816_);
  xor g_119592_(out[340], out[628], _061817_);
  or g_119593_(_061807_, _061812_, _061818_);
  xor g_119594_(out[345], out[633], _061820_);
  or g_119595_(_061802_, _061803_, _061821_);
  or g_119596_(_061818_, _061821_, _061822_);
  or g_119597_(_061809_, _061820_, _061823_);
  or g_119598_(_061814_, _061823_, _061824_);
  or g_119599_(_061822_, _061824_, _061825_);
  or g_119600_(_061810_, _061817_, _061826_);
  or g_119601_(_061825_, _061826_, _061827_);
  or g_119602_(_061805_, _061811_, _061828_);
  xor g_119603_(out[343], out[631], _061829_);
  or g_119604_(_061815_, _061829_, _061831_);
  or g_119605_(_061828_, _061831_, _061832_);
  or g_119606_(_061804_, _061806_, _061833_);
  or g_119607_(_061813_, _061833_, _061834_);
  or g_119608_(_061832_, _061834_, _061835_);
  or g_119609_(_061816_, _061835_, _061836_);
  or g_119610_(_061827_, _061836_, _061837_);
  xor g_119611_(out[327], out[631], _061838_);
  and g_119612_(_098294_, out[635], _061839_);
  xor g_119613_(out[334], out[638], _061840_);
  xor g_119614_(out[328], out[632], _061842_);
  xor g_119615_(out[321], out[625], _061843_);
  xor g_119616_(out[333], out[637], _061844_);
  xor g_119617_(out[329], out[633], _061845_);
  xor g_119618_(out[324], out[628], _061846_);
  xor g_119619_(out[322], out[626], _061847_);
  and g_119620_(out[331], _049598_, _061848_);
  xor g_119621_(out[323], out[627], _061849_);
  xor g_119622_(out[326], out[630], _061850_);
  xor g_119623_(out[335], out[639], _061851_);
  xor g_119624_(out[330], out[634], _061853_);
  xor g_119625_(out[325], out[629], _061854_);
  xor g_119626_(out[320], out[624], _061855_);
  or g_119627_(_061840_, _061846_, _061856_);
  or g_119628_(_061842_, _061844_, _061857_);
  or g_119629_(_061847_, _061853_, _061858_);
  or g_119630_(_061857_, _061858_, _061859_);
  or g_119631_(_061845_, _061849_, _061860_);
  or g_119632_(_061854_, _061855_, _061861_);
  or g_119633_(_061860_, _061861_, _061862_);
  or g_119634_(_061859_, _061862_, _061864_);
  xor g_119635_(out[332], out[636], _061865_);
  or g_119636_(_061839_, _061865_, _061866_);
  or g_119637_(_061838_, _061850_, _061867_);
  or g_119638_(_061866_, _061867_, _061868_);
  or g_119639_(_061843_, _061848_, _061869_);
  or g_119640_(_061851_, _061869_, _061870_);
  or g_119641_(_061868_, _061870_, _061871_);
  or g_119642_(_061864_, _061871_, _061872_);
  or g_119643_(_061856_, _061872_, _061873_);
  xor g_119644_(out[317], out[637], _061875_);
  xor g_119645_(out[306], out[626], _061876_);
  xor g_119646_(out[309], out[629], _061877_);
  xor g_119647_(out[313], out[633], _061878_);
  xor g_119648_(out[308], out[628], _061879_);
  xor g_119649_(out[312], out[632], _061880_);
  xor g_119650_(out[318], out[638], _061881_);
  xor g_119651_(out[310], out[630], _061882_);
  xor g_119652_(out[319], out[639], _061883_);
  xor g_119653_(out[314], out[634], _061884_);
  xor g_119654_(out[304], out[624], _061886_);
  xor g_119655_(out[307], out[627], _061887_);
  and g_119656_(_098283_, out[635], _061888_);
  and g_119657_(out[315], _049598_, _061889_);
  xor g_119658_(out[305], out[625], _061890_);
  or g_119659_(_061879_, _061881_, _061891_);
  or g_119660_(_061875_, _061880_, _061892_);
  or g_119661_(_061876_, _061884_, _061893_);
  or g_119662_(_061892_, _061893_, _061894_);
  or g_119663_(_061878_, _061887_, _061895_);
  or g_119664_(_061877_, _061886_, _061897_);
  or g_119665_(_061895_, _061897_, _061898_);
  or g_119666_(_061894_, _061898_, _061899_);
  xor g_119667_(out[316], out[636], _061900_);
  or g_119668_(_061888_, _061900_, _061901_);
  xor g_119669_(out[311], out[631], _061902_);
  or g_119670_(_061882_, _061902_, _061903_);
  or g_119671_(_061901_, _061903_, _061904_);
  or g_119672_(_061889_, _061890_, _061905_);
  or g_119673_(_061883_, _061905_, _061906_);
  or g_119674_(_061904_, _061906_, _061908_);
  or g_119675_(_061899_, _061908_, _061909_);
  or g_119676_(_061891_, _061909_, _061910_);
  xor g_119677_(out[295], out[631], _061911_);
  and g_119678_(_098272_, out[635], _061912_);
  xor g_119679_(out[302], out[638], _061913_);
  xor g_119680_(out[296], out[632], _061914_);
  xor g_119681_(out[289], out[625], _061915_);
  xor g_119682_(out[301], out[637], _061916_);
  xor g_119683_(out[297], out[633], _061917_);
  xor g_119684_(out[292], out[628], _061919_);
  xor g_119685_(out[290], out[626], _061920_);
  and g_119686_(out[299], _049598_, _061921_);
  xor g_119687_(out[291], out[627], _061922_);
  xor g_119688_(out[294], out[630], _061923_);
  xor g_119689_(out[303], out[639], _061924_);
  xor g_119690_(out[298], out[634], _061925_);
  xor g_119691_(out[293], out[629], _061926_);
  xor g_119692_(out[288], out[624], _061927_);
  or g_119693_(_061913_, _061919_, _061928_);
  or g_119694_(_061914_, _061916_, _061930_);
  or g_119695_(_061920_, _061925_, _061931_);
  or g_119696_(_061930_, _061931_, _061932_);
  or g_119697_(_061917_, _061922_, _061933_);
  or g_119698_(_061926_, _061927_, _061934_);
  or g_119699_(_061933_, _061934_, _061935_);
  or g_119700_(_061932_, _061935_, _061936_);
  xor g_119701_(out[300], out[636], _061937_);
  or g_119702_(_061912_, _061937_, _061938_);
  or g_119703_(_061911_, _061923_, _061939_);
  or g_119704_(_061938_, _061939_, _061941_);
  or g_119705_(_061915_, _061921_, _061942_);
  or g_119706_(_061924_, _061942_, _061943_);
  or g_119707_(_061941_, _061943_, _061944_);
  or g_119708_(_061936_, _061944_, _061945_);
  or g_119709_(_061928_, _061945_, _061946_);
  not g_119710_(_061946_, _061947_);
  xor g_119711_(out[273], out[625], _061948_);
  and g_119712_(out[283], _049598_, _061949_);
  xor g_119713_(out[281], out[633], _061950_);
  xor g_119714_(out[272], out[624], _061952_);
  xor g_119715_(out[286], out[638], _061953_);
  xor g_119716_(out[276], out[628], _061954_);
  or g_119717_(_061953_, _061954_, _061955_);
  xor g_119718_(out[285], out[637], _061956_);
  xor g_119719_(out[275], out[627], _061957_);
  and g_119720_(_098261_, out[635], _061958_);
  xor g_119721_(out[278], out[630], _061959_);
  xor g_119722_(out[282], out[634], _061960_);
  xor g_119723_(out[277], out[629], _061961_);
  xor g_119724_(out[287], out[639], _061963_);
  xor g_119725_(out[280], out[632], _061964_);
  or g_119726_(_061956_, _061964_, _061965_);
  xor g_119727_(out[274], out[626], _061966_);
  or g_119728_(_061960_, _061966_, _061967_);
  or g_119729_(_061965_, _061967_, _061968_);
  or g_119730_(_061950_, _061957_, _061969_);
  or g_119731_(_061961_, _061969_, _061970_);
  or g_119732_(_061968_, _061970_, _061971_);
  or g_119733_(_061955_, _061971_, _061972_);
  xor g_119734_(out[284], out[636], _061974_);
  or g_119735_(_061958_, _061974_, _061975_);
  xor g_119736_(out[279], out[631], _061976_);
  or g_119737_(_061959_, _061976_, _061977_);
  or g_119738_(_061975_, _061977_, _061978_);
  or g_119739_(_061948_, _061949_, _061979_);
  or g_119740_(_061963_, _061979_, _061980_);
  or g_119741_(_061978_, _061980_, _061981_);
  or g_119742_(_061952_, _061981_, _061982_);
  or g_119743_(_061972_, _061982_, _061983_);
  xor g_119744_(out[263], out[631], _061985_);
  and g_119745_(_098250_, out[635], _061986_);
  xor g_119746_(out[270], out[638], _061987_);
  xor g_119747_(out[264], out[632], _061988_);
  xor g_119748_(out[257], out[625], _061989_);
  xor g_119749_(out[269], out[637], _061990_);
  xor g_119750_(out[265], out[633], _061991_);
  xor g_119751_(out[260], out[628], _061992_);
  xor g_119752_(out[258], out[626], _061993_);
  and g_119753_(out[267], _049598_, _061994_);
  xor g_119754_(out[259], out[627], _061996_);
  xor g_119755_(out[262], out[630], _061997_);
  xor g_119756_(out[271], out[639], _061998_);
  xor g_119757_(out[266], out[634], _061999_);
  xor g_119758_(out[261], out[629], _062000_);
  xor g_119759_(out[256], out[624], _062001_);
  or g_119760_(_061987_, _061992_, _062002_);
  or g_119761_(_061988_, _061990_, _062003_);
  or g_119762_(_061993_, _061999_, _062004_);
  or g_119763_(_062003_, _062004_, _062005_);
  or g_119764_(_061991_, _061996_, _062007_);
  or g_119765_(_062000_, _062001_, _062008_);
  or g_119766_(_062007_, _062008_, _062009_);
  or g_119767_(_062005_, _062009_, _062010_);
  xor g_119768_(out[268], out[636], _062011_);
  or g_119769_(_061986_, _062011_, _062012_);
  or g_119770_(_061985_, _061997_, _062013_);
  or g_119771_(_062012_, _062013_, _062014_);
  or g_119772_(_061989_, _061994_, _062015_);
  or g_119773_(_061998_, _062015_, _062016_);
  or g_119774_(_062014_, _062016_, _062018_);
  or g_119775_(_062010_, _062018_, _062019_);
  or g_119776_(_062002_, _062019_, _062020_);
  xor g_119777_(out[241], out[625], _062021_);
  and g_119778_(out[251], _049598_, _062022_);
  xor g_119779_(out[249], out[633], _062023_);
  xor g_119780_(out[240], out[624], _062024_);
  xor g_119781_(out[254], out[638], _062025_);
  xor g_119782_(out[244], out[628], _062026_);
  or g_119783_(_062025_, _062026_, _062027_);
  xor g_119784_(out[253], out[637], _062029_);
  xor g_119785_(out[243], out[627], _062030_);
  and g_119786_(_098239_, out[635], _062031_);
  xor g_119787_(out[246], out[630], _062032_);
  xor g_119788_(out[250], out[634], _062033_);
  xor g_119789_(out[245], out[629], _062034_);
  xor g_119790_(out[255], out[639], _062035_);
  xor g_119791_(out[248], out[632], _062036_);
  or g_119792_(_062029_, _062036_, _062037_);
  xor g_119793_(out[242], out[626], _062038_);
  or g_119794_(_062033_, _062038_, _062040_);
  or g_119795_(_062037_, _062040_, _062041_);
  or g_119796_(_062023_, _062030_, _062042_);
  or g_119797_(_062034_, _062042_, _062043_);
  or g_119798_(_062041_, _062043_, _062044_);
  or g_119799_(_062027_, _062044_, _062045_);
  xor g_119800_(out[252], out[636], _062046_);
  or g_119801_(_062031_, _062046_, _062047_);
  xor g_119802_(out[247], out[631], _062048_);
  or g_119803_(_062032_, _062048_, _062049_);
  or g_119804_(_062047_, _062049_, _062051_);
  or g_119805_(_062021_, _062022_, _062052_);
  or g_119806_(_062035_, _062052_, _062053_);
  or g_119807_(_062051_, _062053_, _062054_);
  or g_119808_(_062024_, _062054_, _062055_);
  or g_119809_(_062045_, _062055_, _062056_);
  not g_119810_(_062056_, _062057_);
  xor g_119811_(out[231], out[631], _062058_);
  and g_119812_(_098228_, out[635], _062059_);
  xor g_119813_(out[238], out[638], _062060_);
  xor g_119814_(out[232], out[632], _062062_);
  xor g_119815_(out[225], out[625], _062063_);
  xor g_119816_(out[237], out[637], _062064_);
  xor g_119817_(out[233], out[633], _062065_);
  xor g_119818_(out[228], out[628], _062066_);
  xor g_119819_(out[226], out[626], _062067_);
  and g_119820_(out[235], _049598_, _062068_);
  xor g_119821_(out[227], out[627], _062069_);
  xor g_119822_(out[230], out[630], _062070_);
  xor g_119823_(out[239], out[639], _062071_);
  xor g_119824_(out[234], out[634], _062073_);
  xor g_119825_(out[229], out[629], _062074_);
  xor g_119826_(out[224], out[624], _062075_);
  or g_119827_(_062060_, _062066_, _062076_);
  or g_119828_(_062062_, _062064_, _062077_);
  or g_119829_(_062067_, _062073_, _062078_);
  or g_119830_(_062077_, _062078_, _062079_);
  or g_119831_(_062065_, _062069_, _062080_);
  or g_119832_(_062074_, _062075_, _062081_);
  or g_119833_(_062080_, _062081_, _062082_);
  or g_119834_(_062079_, _062082_, _062084_);
  xor g_119835_(out[236], out[636], _062085_);
  or g_119836_(_062059_, _062085_, _062086_);
  or g_119837_(_062058_, _062070_, _062087_);
  or g_119838_(_062086_, _062087_, _062088_);
  or g_119839_(_062063_, _062068_, _062089_);
  or g_119840_(_062071_, _062089_, _062090_);
  or g_119841_(_062088_, _062090_, _062091_);
  or g_119842_(_062084_, _062091_, _062092_);
  or g_119843_(_062076_, _062092_, _062093_);
  and g_119844_(out[219], _049598_, _062095_);
  xor g_119845_(out[212], out[628], _062096_);
  xor g_119846_(out[222], out[638], _062097_);
  or g_119847_(_062096_, _062097_, _062098_);
  xor g_119848_(out[221], out[637], _062099_);
  xor g_119849_(out[211], out[627], _062100_);
  xor g_119850_(out[208], out[624], _062101_);
  and g_119851_(_098217_, out[635], _062102_);
  xor g_119852_(out[218], out[634], _062103_);
  xor g_119853_(out[223], out[639], _062104_);
  xor g_119854_(out[214], out[630], _062106_);
  xor g_119855_(out[213], out[629], _062107_);
  xor g_119856_(out[216], out[632], _062108_);
  or g_119857_(_062099_, _062108_, _062109_);
  xor g_119858_(out[210], out[626], _062110_);
  xor g_119859_(out[217], out[633], _062111_);
  xor g_119860_(out[209], out[625], _062112_);
  or g_119861_(_062103_, _062110_, _062113_);
  or g_119862_(_062109_, _062113_, _062114_);
  or g_119863_(_062100_, _062111_, _062115_);
  or g_119864_(_062107_, _062115_, _062117_);
  or g_119865_(_062114_, _062117_, _062118_);
  or g_119866_(_062098_, _062118_, _062119_);
  xor g_119867_(out[220], out[636], _062120_);
  or g_119868_(_062102_, _062120_, _062121_);
  xor g_119869_(out[215], out[631], _062122_);
  or g_119870_(_062106_, _062122_, _062123_);
  or g_119871_(_062121_, _062123_, _062124_);
  or g_119872_(_062095_, _062112_, _062125_);
  or g_119873_(_062104_, _062125_, _062126_);
  or g_119874_(_062124_, _062126_, _062128_);
  or g_119875_(_062101_, _062128_, _062129_);
  or g_119876_(_062119_, _062129_, _062130_);
  xor g_119877_(out[199], out[631], _062131_);
  and g_119878_(_098206_, out[635], _062132_);
  xor g_119879_(out[206], out[638], _062133_);
  xor g_119880_(out[200], out[632], _062134_);
  xor g_119881_(out[193], out[625], _062135_);
  xor g_119882_(out[205], out[637], _062136_);
  xor g_119883_(out[201], out[633], _062137_);
  xor g_119884_(out[196], out[628], _062139_);
  xor g_119885_(out[194], out[626], _062140_);
  and g_119886_(out[203], _049598_, _062141_);
  xor g_119887_(out[195], out[627], _062142_);
  xor g_119888_(out[198], out[630], _062143_);
  xor g_119889_(out[207], out[639], _062144_);
  xor g_119890_(out[202], out[634], _062145_);
  xor g_119891_(out[197], out[629], _062146_);
  xor g_119892_(out[192], out[624], _062147_);
  or g_119893_(_062133_, _062139_, _062148_);
  or g_119894_(_062134_, _062136_, _062150_);
  or g_119895_(_062140_, _062145_, _062151_);
  or g_119896_(_062150_, _062151_, _062152_);
  or g_119897_(_062137_, _062142_, _062153_);
  or g_119898_(_062146_, _062147_, _062154_);
  or g_119899_(_062153_, _062154_, _062155_);
  or g_119900_(_062152_, _062155_, _062156_);
  xor g_119901_(out[204], out[636], _062157_);
  or g_119902_(_062132_, _062157_, _062158_);
  or g_119903_(_062131_, _062143_, _062159_);
  or g_119904_(_062158_, _062159_, _062161_);
  or g_119905_(_062135_, _062141_, _062162_);
  or g_119906_(_062144_, _062162_, _062163_);
  or g_119907_(_062161_, _062163_, _062164_);
  or g_119908_(_062156_, _062164_, _062165_);
  or g_119909_(_062148_, _062165_, _062166_);
  xor g_119910_(out[177], out[625], _062167_);
  and g_119911_(out[187], _049598_, _062168_);
  xor g_119912_(out[185], out[633], _062169_);
  xor g_119913_(out[176], out[624], _062170_);
  xor g_119914_(out[190], out[638], _062172_);
  xor g_119915_(out[180], out[628], _062173_);
  or g_119916_(_062172_, _062173_, _062174_);
  xor g_119917_(out[189], out[637], _062175_);
  xor g_119918_(out[179], out[627], _062176_);
  and g_119919_(_098195_, out[635], _062177_);
  xor g_119920_(out[182], out[630], _062178_);
  xor g_119921_(out[186], out[634], _062179_);
  xor g_119922_(out[181], out[629], _062180_);
  xor g_119923_(out[191], out[639], _062181_);
  xor g_119924_(out[184], out[632], _062183_);
  or g_119925_(_062175_, _062183_, _062184_);
  xor g_119926_(out[178], out[626], _062185_);
  or g_119927_(_062179_, _062185_, _062186_);
  or g_119928_(_062184_, _062186_, _062187_);
  or g_119929_(_062169_, _062176_, _062188_);
  or g_119930_(_062180_, _062188_, _062189_);
  or g_119931_(_062187_, _062189_, _062190_);
  or g_119932_(_062174_, _062190_, _062191_);
  xor g_119933_(out[188], out[636], _062192_);
  or g_119934_(_062177_, _062192_, _062194_);
  xor g_119935_(out[183], out[631], _062195_);
  or g_119936_(_062178_, _062195_, _062196_);
  or g_119937_(_062194_, _062196_, _062197_);
  or g_119938_(_062167_, _062168_, _062198_);
  or g_119939_(_062181_, _062198_, _062199_);
  or g_119940_(_062197_, _062199_, _062200_);
  or g_119941_(_062170_, _062200_, _062201_);
  or g_119942_(_062191_, _062201_, _062202_);
  xor g_119943_(out[167], out[631], _062203_);
  and g_119944_(_098184_, out[635], _062205_);
  xor g_119945_(out[174], out[638], _062206_);
  xor g_119946_(out[168], out[632], _062207_);
  xor g_119947_(out[161], out[625], _062208_);
  xor g_119948_(out[173], out[637], _062209_);
  xor g_119949_(out[169], out[633], _062210_);
  xor g_119950_(out[164], out[628], _062211_);
  xor g_119951_(out[162], out[626], _062212_);
  and g_119952_(out[171], _049598_, _062213_);
  xor g_119953_(out[163], out[627], _062214_);
  xor g_119954_(out[166], out[630], _062216_);
  xor g_119955_(out[175], out[639], _062217_);
  xor g_119956_(out[170], out[634], _062218_);
  xor g_119957_(out[165], out[629], _062219_);
  xor g_119958_(out[160], out[624], _062220_);
  or g_119959_(_062206_, _062211_, _062221_);
  or g_119960_(_062207_, _062209_, _062222_);
  or g_119961_(_062212_, _062218_, _062223_);
  or g_119962_(_062222_, _062223_, _062224_);
  or g_119963_(_062210_, _062214_, _062225_);
  or g_119964_(_062219_, _062220_, _062227_);
  or g_119965_(_062225_, _062227_, _062228_);
  or g_119966_(_062224_, _062228_, _062229_);
  xor g_119967_(out[172], out[636], _062230_);
  or g_119968_(_062205_, _062230_, _062231_);
  or g_119969_(_062203_, _062216_, _062232_);
  or g_119970_(_062231_, _062232_, _062233_);
  or g_119971_(_062208_, _062213_, _062234_);
  or g_119972_(_062217_, _062234_, _062235_);
  or g_119973_(_062233_, _062235_, _062236_);
  or g_119974_(_062229_, _062236_, _062238_);
  or g_119975_(_062221_, _062238_, _062239_);
  xor g_119976_(out[145], out[625], _062240_);
  and g_119977_(_098173_, out[635], _062241_);
  and g_119978_(out[155], _049598_, _062242_);
  xor g_119979_(out[153], out[633], _062243_);
  xor g_119980_(out[144], out[624], _062244_);
  xor g_119981_(out[158], out[638], _062245_);
  xor g_119982_(out[148], out[628], _062246_);
  or g_119983_(_062245_, _062246_, _062247_);
  xor g_119984_(out[157], out[637], _062249_);
  xor g_119985_(out[147], out[627], _062250_);
  xor g_119986_(out[156], out[636], _062251_);
  xor g_119987_(out[150], out[630], _062252_);
  xor g_119988_(out[154], out[634], _062253_);
  xor g_119989_(out[149], out[629], _062254_);
  xor g_119990_(out[159], out[639], _062255_);
  xor g_119991_(out[152], out[632], _062256_);
  or g_119992_(_062249_, _062256_, _062257_);
  xor g_119993_(out[146], out[626], _062258_);
  or g_119994_(_062253_, _062258_, _062260_);
  or g_119995_(_062257_, _062260_, _062261_);
  or g_119996_(_062243_, _062250_, _062262_);
  or g_119997_(_062254_, _062262_, _062263_);
  or g_119998_(_062261_, _062263_, _062264_);
  or g_119999_(_062247_, _062264_, _062265_);
  or g_120000_(_062241_, _062251_, _062266_);
  xor g_120001_(out[151], out[631], _062267_);
  or g_120002_(_062252_, _062267_, _062268_);
  or g_120003_(_062266_, _062268_, _062269_);
  or g_120004_(_062240_, _062242_, _062271_);
  or g_120005_(_062255_, _062271_, _062272_);
  or g_120006_(_062269_, _062272_, _062273_);
  or g_120007_(_062244_, _062273_, _062274_);
  or g_120008_(_062265_, _062274_, _062275_);
  not g_120009_(_062275_, _062276_);
  xor g_120010_(out[135], out[631], _062277_);
  and g_120011_(_098162_, out[635], _062278_);
  xor g_120012_(out[142], out[638], _062279_);
  xor g_120013_(out[136], out[632], _062280_);
  xor g_120014_(out[129], out[625], _062282_);
  xor g_120015_(out[141], out[637], _062283_);
  xor g_120016_(out[137], out[633], _062284_);
  xor g_120017_(out[132], out[628], _062285_);
  xor g_120018_(out[130], out[626], _062286_);
  and g_120019_(out[139], _049598_, _062287_);
  xor g_120020_(out[131], out[627], _062288_);
  xor g_120021_(out[134], out[630], _062289_);
  xor g_120022_(out[143], out[639], _062290_);
  xor g_120023_(out[138], out[634], _062291_);
  xor g_120024_(out[133], out[629], _062293_);
  xor g_120025_(out[128], out[624], _062294_);
  or g_120026_(_062279_, _062285_, _062295_);
  or g_120027_(_062280_, _062283_, _062296_);
  or g_120028_(_062286_, _062291_, _062297_);
  or g_120029_(_062296_, _062297_, _062298_);
  or g_120030_(_062284_, _062288_, _062299_);
  or g_120031_(_062293_, _062294_, _062300_);
  or g_120032_(_062299_, _062300_, _062301_);
  or g_120033_(_062298_, _062301_, _062302_);
  xor g_120034_(out[140], out[636], _062304_);
  or g_120035_(_062278_, _062304_, _062305_);
  or g_120036_(_062277_, _062289_, _062306_);
  or g_120037_(_062305_, _062306_, _062307_);
  or g_120038_(_062282_, _062287_, _062308_);
  or g_120039_(_062290_, _062308_, _062309_);
  or g_120040_(_062307_, _062309_, _062310_);
  or g_120041_(_062302_, _062310_, _062311_);
  or g_120042_(_062295_, _062311_, _062312_);
  xor g_120043_(out[113], out[625], _062313_);
  and g_120044_(out[123], _049598_, _062315_);
  xor g_120045_(out[121], out[633], _062316_);
  xor g_120046_(out[112], out[624], _062317_);
  xor g_120047_(out[126], out[638], _062318_);
  xor g_120048_(out[116], out[628], _062319_);
  or g_120049_(_062318_, _062319_, _062320_);
  xor g_120050_(out[125], out[637], _062321_);
  xor g_120051_(out[115], out[627], _062322_);
  and g_120052_(_098151_, out[635], _062323_);
  xor g_120053_(out[118], out[630], _062324_);
  xor g_120054_(out[122], out[634], _062326_);
  xor g_120055_(out[117], out[629], _062327_);
  xor g_120056_(out[127], out[639], _062328_);
  xor g_120057_(out[120], out[632], _062329_);
  or g_120058_(_062321_, _062329_, _062330_);
  xor g_120059_(out[114], out[626], _062331_);
  or g_120060_(_062326_, _062331_, _062332_);
  or g_120061_(_062330_, _062332_, _062333_);
  or g_120062_(_062316_, _062322_, _062334_);
  or g_120063_(_062327_, _062334_, _062335_);
  or g_120064_(_062333_, _062335_, _062337_);
  or g_120065_(_062320_, _062337_, _062338_);
  xor g_120066_(out[124], out[636], _062339_);
  or g_120067_(_062323_, _062339_, _062340_);
  xor g_120068_(out[119], out[631], _062341_);
  or g_120069_(_062324_, _062341_, _062342_);
  or g_120070_(_062340_, _062342_, _062343_);
  or g_120071_(_062313_, _062315_, _062344_);
  or g_120072_(_062328_, _062344_, _062345_);
  or g_120073_(_062343_, _062345_, _062346_);
  or g_120074_(_062317_, _062346_, _062348_);
  or g_120075_(_062338_, _062348_, _062349_);
  xor g_120076_(out[103], out[631], _062350_);
  and g_120077_(_098140_, out[635], _062351_);
  xor g_120078_(out[110], out[638], _062352_);
  xor g_120079_(out[104], out[632], _062353_);
  xor g_120080_(out[97], out[625], _062354_);
  xor g_120081_(out[109], out[637], _062355_);
  xor g_120082_(out[105], out[633], _062356_);
  xor g_120083_(out[100], out[628], _062357_);
  xor g_120084_(out[98], out[626], _062359_);
  and g_120085_(out[107], _049598_, _062360_);
  xor g_120086_(out[99], out[627], _062361_);
  xor g_120087_(out[102], out[630], _062362_);
  xor g_120088_(out[111], out[639], _062363_);
  xor g_120089_(out[106], out[634], _062364_);
  xor g_120090_(out[101], out[629], _062365_);
  xor g_120091_(out[96], out[624], _062366_);
  or g_120092_(_062352_, _062357_, _062367_);
  or g_120093_(_062353_, _062355_, _062368_);
  or g_120094_(_062359_, _062364_, _062370_);
  or g_120095_(_062368_, _062370_, _062371_);
  or g_120096_(_062356_, _062361_, _062372_);
  or g_120097_(_062365_, _062366_, _062373_);
  or g_120098_(_062372_, _062373_, _062374_);
  or g_120099_(_062371_, _062374_, _062375_);
  xor g_120100_(out[108], out[636], _062376_);
  or g_120101_(_062351_, _062376_, _062377_);
  or g_120102_(_062350_, _062362_, _062378_);
  or g_120103_(_062377_, _062378_, _062379_);
  or g_120104_(_062354_, _062360_, _062381_);
  or g_120105_(_062363_, _062381_, _062382_);
  or g_120106_(_062379_, _062382_, _062383_);
  or g_120107_(_062375_, _062383_, _062384_);
  or g_120108_(_062367_, _062384_, _062385_);
  xor g_120109_(out[81], out[625], _062386_);
  and g_120110_(out[91], _049598_, _062387_);
  xor g_120111_(out[94], out[638], _062388_);
  xor g_120112_(out[83], out[627], _062389_);
  xor g_120113_(out[84], out[628], _062390_);
  xor g_120114_(out[82], out[626], _062392_);
  xor g_120115_(out[89], out[633], _062393_);
  xor g_120116_(out[80], out[624], _062394_);
  and g_120117_(_098129_, out[635], _062395_);
  xor g_120118_(out[86], out[630], _062396_);
  xor g_120119_(out[90], out[634], _062397_);
  xor g_120120_(out[85], out[629], _062398_);
  xor g_120121_(out[95], out[639], _062399_);
  xor g_120122_(out[93], out[637], _062400_);
  xor g_120123_(out[88], out[632], _062401_);
  or g_120124_(_062388_, _062390_, _062403_);
  or g_120125_(_062400_, _062401_, _062404_);
  or g_120126_(_062392_, _062397_, _062405_);
  or g_120127_(_062404_, _062405_, _062406_);
  or g_120128_(_062389_, _062393_, _062407_);
  or g_120129_(_062394_, _062398_, _062408_);
  or g_120130_(_062407_, _062408_, _062409_);
  or g_120131_(_062406_, _062409_, _062410_);
  xor g_120132_(out[92], out[636], _062411_);
  or g_120133_(_062395_, _062411_, _062412_);
  xor g_120134_(out[87], out[631], _062414_);
  or g_120135_(_062396_, _062414_, _062415_);
  or g_120136_(_062412_, _062415_, _062416_);
  or g_120137_(_062386_, _062387_, _062417_);
  or g_120138_(_062399_, _062417_, _062418_);
  or g_120139_(_062416_, _062418_, _062419_);
  or g_120140_(_062410_, _062419_, _062420_);
  or g_120141_(_062403_, _062420_, _062421_);
  xor g_120142_(out[71], out[631], _062422_);
  and g_120143_(_098118_, out[635], _062423_);
  xor g_120144_(out[78], out[638], _062425_);
  xor g_120145_(out[72], out[632], _062426_);
  xor g_120146_(out[65], out[625], _062427_);
  xor g_120147_(out[77], out[637], _062428_);
  xor g_120148_(out[73], out[633], _062429_);
  xor g_120149_(out[68], out[628], _062430_);
  xor g_120150_(out[66], out[626], _062431_);
  and g_120151_(out[75], _049598_, _062432_);
  xor g_120152_(out[67], out[627], _062433_);
  xor g_120153_(out[70], out[630], _062434_);
  xor g_120154_(out[79], out[639], _062436_);
  xor g_120155_(out[74], out[634], _062437_);
  xor g_120156_(out[69], out[629], _062438_);
  xor g_120157_(out[64], out[624], _062439_);
  or g_120158_(_062425_, _062430_, _062440_);
  or g_120159_(_062426_, _062428_, _062441_);
  or g_120160_(_062431_, _062437_, _062442_);
  or g_120161_(_062441_, _062442_, _062443_);
  or g_120162_(_062429_, _062433_, _062444_);
  or g_120163_(_062438_, _062439_, _062445_);
  or g_120164_(_062444_, _062445_, _062447_);
  or g_120165_(_062443_, _062447_, _062448_);
  xor g_120166_(out[76], out[636], _062449_);
  or g_120167_(_062423_, _062449_, _062450_);
  or g_120168_(_062422_, _062434_, _062451_);
  or g_120169_(_062450_, _062451_, _062452_);
  or g_120170_(_062427_, _062432_, _062453_);
  or g_120171_(_062436_, _062453_, _062454_);
  or g_120172_(_062452_, _062454_, _062455_);
  or g_120173_(_062448_, _062455_, _062456_);
  or g_120174_(_062440_, _062456_, _062458_);
  xor g_120175_(out[58], out[634], _062459_);
  xor g_120176_(out[56], out[632], _062460_);
  xor g_120177_(out[49], out[625], _062461_);
  and g_120178_(_098107_, out[635], _062462_);
  and g_120179_(out[59], _049598_, _062463_);
  xor g_120180_(out[50], out[626], _062464_);
  xor g_120181_(out[53], out[629], _062465_);
  xor g_120182_(out[57], out[633], _062466_);
  xor g_120183_(out[60], out[636], _062467_);
  xor g_120184_(out[61], out[637], _062469_);
  xor g_120185_(out[63], out[639], _062470_);
  xor g_120186_(out[52], out[628], _062471_);
  xor g_120187_(out[54], out[630], _062472_);
  xor g_120188_(out[51], out[627], _062473_);
  xor g_120189_(out[48], out[624], _062474_);
  xor g_120190_(out[62], out[638], _062475_);
  or g_120191_(_062471_, _062475_, _062476_);
  or g_120192_(_062460_, _062469_, _062477_);
  or g_120193_(_062459_, _062464_, _062478_);
  or g_120194_(_062477_, _062478_, _062480_);
  or g_120195_(_062466_, _062473_, _062481_);
  or g_120196_(_062465_, _062474_, _062482_);
  or g_120197_(_062481_, _062482_, _062483_);
  or g_120198_(_062480_, _062483_, _062484_);
  or g_120199_(_062462_, _062467_, _062485_);
  xor g_120200_(out[55], out[631], _062486_);
  or g_120201_(_062472_, _062486_, _062487_);
  or g_120202_(_062485_, _062487_, _062488_);
  or g_120203_(_062461_, _062463_, _062489_);
  or g_120204_(_062470_, _062489_, _062491_);
  or g_120205_(_062488_, _062491_, _062492_);
  or g_120206_(_062484_, _062492_, _062493_);
  or g_120207_(_062476_, _062493_, _062494_);
  xor g_120208_(out[39], out[631], _062495_);
  and g_120209_(_098096_, out[635], _062496_);
  xor g_120210_(out[46], out[638], _062497_);
  xor g_120211_(out[40], out[632], _062498_);
  xor g_120212_(out[33], out[625], _062499_);
  xor g_120213_(out[45], out[637], _062500_);
  xor g_120214_(out[41], out[633], _062502_);
  xor g_120215_(out[36], out[628], _062503_);
  xor g_120216_(out[34], out[626], _062504_);
  and g_120217_(out[43], _049598_, _062505_);
  xor g_120218_(out[35], out[627], _062506_);
  xor g_120219_(out[38], out[630], _062507_);
  xor g_120220_(out[47], out[639], _062508_);
  xor g_120221_(out[42], out[634], _062509_);
  xor g_120222_(out[37], out[629], _062510_);
  xor g_120223_(out[32], out[624], _062511_);
  or g_120224_(_062497_, _062503_, _062513_);
  or g_120225_(_062498_, _062500_, _062514_);
  or g_120226_(_062504_, _062509_, _062515_);
  or g_120227_(_062514_, _062515_, _062516_);
  or g_120228_(_062502_, _062506_, _062517_);
  or g_120229_(_062510_, _062511_, _062518_);
  or g_120230_(_062517_, _062518_, _062519_);
  or g_120231_(_062516_, _062519_, _062520_);
  xor g_120232_(out[44], out[636], _062521_);
  or g_120233_(_062496_, _062521_, _062522_);
  or g_120234_(_062495_, _062507_, _062524_);
  or g_120235_(_062522_, _062524_, _062525_);
  or g_120236_(_062499_, _062505_, _062526_);
  or g_120237_(_062508_, _062526_, _062527_);
  or g_120238_(_062525_, _062527_, _062528_);
  or g_120239_(_062520_, _062528_, _062529_);
  or g_120240_(_062513_, _062529_, _062530_);
  xor g_120241_(out[19], out[627], _062531_);
  xor g_120242_(out[20], out[628], _062532_);
  xor g_120243_(out[30], out[638], _062533_);
  xor g_120244_(out[18], out[626], _062535_);
  xor g_120245_(out[21], out[629], _062536_);
  xor g_120246_(out[25], out[633], _062537_);
  xor g_120247_(out[24], out[632], _062538_);
  xor g_120248_(out[31], out[639], _062539_);
  xor g_120249_(out[26], out[634], _062540_);
  xor g_120250_(out[22], out[630], _062541_);
  xor g_120251_(out[16], out[624], _062542_);
  and g_120252_(_098063_, out[635], _062543_);
  and g_120253_(out[27], _049598_, _062544_);
  xor g_120254_(out[29], out[637], _062546_);
  or g_120255_(_062538_, _062546_, _062547_);
  xor g_120256_(out[17], out[625], _062548_);
  or g_120257_(_062535_, _062540_, _062549_);
  or g_120258_(_062547_, _062549_, _062550_);
  or g_120259_(_062531_, _062537_, _062551_);
  or g_120260_(_062536_, _062551_, _062552_);
  or g_120261_(_062550_, _062552_, _062553_);
  or g_120262_(_062532_, _062533_, _062554_);
  or g_120263_(_062553_, _062554_, _062555_);
  xor g_120264_(out[28], out[636], _062557_);
  or g_120265_(_062543_, _062557_, _062558_);
  xor g_120266_(out[23], out[631], _062559_);
  or g_120267_(_062541_, _062559_, _062560_);
  or g_120268_(_062558_, _062560_, _062561_);
  or g_120269_(_062544_, _062548_, _062562_);
  or g_120270_(_062539_, _062562_, _062563_);
  or g_120271_(_062561_, _062563_, _062564_);
  or g_120272_(_062542_, _062564_, _062565_);
  or g_120273_(_062555_, _062565_, _062566_);
  xor g_120274_(out[1], out[625], _062568_);
  and g_120275_(out[11], _049598_, _062569_);
  xor g_120276_(out[14], out[638], _062570_);
  xor g_120277_(out[3], out[627], _062571_);
  xor g_120278_(out[4], out[628], _062572_);
  xor g_120279_(out[2], out[626], _062573_);
  xor g_120280_(out[9], out[633], _062574_);
  xor g_120281_(out[0], out[624], _062575_);
  and g_120282_(_098041_, out[635], _062576_);
  xor g_120283_(out[6], out[630], _062577_);
  xor g_120284_(out[10], out[634], _062579_);
  xor g_120285_(out[5], out[629], _062580_);
  xor g_120286_(out[15], out[639], _062581_);
  xor g_120287_(out[13], out[637], _062582_);
  xor g_120288_(out[8], out[632], _062583_);
  or g_120289_(_062570_, _062572_, _062584_);
  or g_120290_(_062582_, _062583_, _062585_);
  or g_120291_(_062573_, _062579_, _062586_);
  or g_120292_(_062585_, _062586_, _062587_);
  or g_120293_(_062571_, _062574_, _062588_);
  or g_120294_(_062575_, _062580_, _062590_);
  or g_120295_(_062588_, _062590_, _062591_);
  or g_120296_(_062587_, _062591_, _062592_);
  xor g_120297_(out[12], out[636], _062593_);
  or g_120298_(_062576_, _062593_, _062594_);
  xor g_120299_(out[7], out[631], _062595_);
  or g_120300_(_062577_, _062595_, _062596_);
  or g_120301_(_062594_, _062596_, _062597_);
  or g_120302_(_062568_, _062569_, _062598_);
  or g_120303_(_062581_, _062598_, _062599_);
  or g_120304_(_062597_, _062599_, _062601_);
  or g_120305_(_062592_, _062601_, _062602_);
  or g_120306_(_062584_, _062602_, _062603_);
  not g_120307_(_062603_, _062604_);
  xor g_120308_(out[471], out[615], _062605_);
  and g_120309_(_049499_, out[619], _062606_);
  xor g_120310_(out[478], out[622], _062607_);
  xor g_120311_(out[472], out[616], _062608_);
  xor g_120312_(out[465], out[609], _062609_);
  xor g_120313_(out[477], out[621], _062610_);
  xor g_120314_(out[473], out[617], _062612_);
  xor g_120315_(out[468], out[612], _062613_);
  xor g_120316_(out[466], out[610], _062614_);
  and g_120317_(out[475], _049587_, _062615_);
  xor g_120318_(out[467], out[611], _062616_);
  xor g_120319_(out[470], out[614], _062617_);
  xor g_120320_(out[479], out[623], _062618_);
  xor g_120321_(out[474], out[618], _062619_);
  xor g_120322_(out[469], out[613], _062620_);
  xor g_120323_(out[464], out[608], _062621_);
  or g_120324_(_062607_, _062613_, _062623_);
  or g_120325_(_062608_, _062610_, _062624_);
  or g_120326_(_062614_, _062619_, _062625_);
  or g_120327_(_062624_, _062625_, _062626_);
  or g_120328_(_062612_, _062616_, _062627_);
  or g_120329_(_062620_, _062621_, _062628_);
  or g_120330_(_062627_, _062628_, _062629_);
  or g_120331_(_062626_, _062629_, _062630_);
  xor g_120332_(out[476], out[620], _062631_);
  or g_120333_(_062606_, _062631_, _062632_);
  or g_120334_(_062605_, _062617_, _062634_);
  or g_120335_(_062632_, _062634_, _062635_);
  or g_120336_(_062609_, _062615_, _062636_);
  or g_120337_(_062618_, _062636_, _062637_);
  or g_120338_(_062635_, _062637_, _062638_);
  or g_120339_(_062630_, _062638_, _062639_);
  or g_120340_(_062623_, _062639_, _062640_);
  xor g_120341_(out[449], out[609], _062641_);
  and g_120342_(out[459], _049587_, _062642_);
  xor g_120343_(out[462], out[622], _062643_);
  xor g_120344_(out[451], out[611], _062645_);
  xor g_120345_(out[452], out[612], _062646_);
  xor g_120346_(out[450], out[610], _062647_);
  xor g_120347_(out[457], out[617], _062648_);
  xor g_120348_(out[448], out[608], _062649_);
  and g_120349_(_049477_, out[619], _062650_);
  xor g_120350_(out[454], out[614], _062651_);
  xor g_120351_(out[458], out[618], _062652_);
  xor g_120352_(out[453], out[613], _062653_);
  xor g_120353_(out[463], out[623], _062654_);
  xor g_120354_(out[461], out[621], _062656_);
  xor g_120355_(out[456], out[616], _062657_);
  or g_120356_(_062643_, _062646_, _062658_);
  or g_120357_(_062656_, _062657_, _062659_);
  or g_120358_(_062647_, _062652_, _062660_);
  or g_120359_(_062659_, _062660_, _062661_);
  or g_120360_(_062645_, _062648_, _062662_);
  or g_120361_(_062649_, _062653_, _062663_);
  or g_120362_(_062662_, _062663_, _062664_);
  or g_120363_(_062661_, _062664_, _062665_);
  xor g_120364_(out[460], out[620], _062667_);
  or g_120365_(_062650_, _062667_, _062668_);
  xor g_120366_(out[455], out[615], _062669_);
  or g_120367_(_062651_, _062669_, _062670_);
  or g_120368_(_062668_, _062670_, _062671_);
  or g_120369_(_062641_, _062642_, _062672_);
  or g_120370_(_062654_, _062672_, _062673_);
  or g_120371_(_062671_, _062673_, _062674_);
  or g_120372_(_062665_, _062674_, _062675_);
  or g_120373_(_062658_, _062675_, _062676_);
  xor g_120374_(out[439], out[615], _062678_);
  and g_120375_(_049466_, out[619], _062679_);
  xor g_120376_(out[446], out[622], _062680_);
  xor g_120377_(out[440], out[616], _062681_);
  xor g_120378_(out[433], out[609], _062682_);
  xor g_120379_(out[445], out[621], _062683_);
  xor g_120380_(out[441], out[617], _062684_);
  xor g_120381_(out[436], out[612], _062685_);
  xor g_120382_(out[434], out[610], _062686_);
  and g_120383_(out[443], _049587_, _062687_);
  xor g_120384_(out[435], out[611], _062689_);
  xor g_120385_(out[438], out[614], _062690_);
  xor g_120386_(out[447], out[623], _062691_);
  xor g_120387_(out[442], out[618], _062692_);
  xor g_120388_(out[437], out[613], _062693_);
  xor g_120389_(out[432], out[608], _062694_);
  or g_120390_(_062680_, _062685_, _062695_);
  or g_120391_(_062681_, _062683_, _062696_);
  or g_120392_(_062686_, _062692_, _062697_);
  or g_120393_(_062696_, _062697_, _062698_);
  or g_120394_(_062684_, _062689_, _062700_);
  or g_120395_(_062693_, _062694_, _062701_);
  or g_120396_(_062700_, _062701_, _062702_);
  or g_120397_(_062698_, _062702_, _062703_);
  xor g_120398_(out[444], out[620], _062704_);
  or g_120399_(_062679_, _062704_, _062705_);
  or g_120400_(_062678_, _062690_, _062706_);
  or g_120401_(_062705_, _062706_, _062707_);
  or g_120402_(_062682_, _062687_, _062708_);
  or g_120403_(_062691_, _062708_, _062709_);
  or g_120404_(_062707_, _062709_, _062711_);
  or g_120405_(_062703_, _062711_, _062712_);
  or g_120406_(_062695_, _062712_, _062713_);
  xor g_120407_(out[417], out[609], _062714_);
  and g_120408_(out[427], _049587_, _062715_);
  xor g_120409_(out[425], out[617], _062716_);
  xor g_120410_(out[416], out[608], _062717_);
  xor g_120411_(out[430], out[622], _062718_);
  xor g_120412_(out[420], out[612], _062719_);
  or g_120413_(_062718_, _062719_, _062720_);
  xor g_120414_(out[429], out[621], _062722_);
  xor g_120415_(out[419], out[611], _062723_);
  and g_120416_(_049455_, out[619], _062724_);
  xor g_120417_(out[422], out[614], _062725_);
  xor g_120418_(out[426], out[618], _062726_);
  xor g_120419_(out[421], out[613], _062727_);
  xor g_120420_(out[431], out[623], _062728_);
  xor g_120421_(out[424], out[616], _062729_);
  or g_120422_(_062722_, _062729_, _062730_);
  xor g_120423_(out[418], out[610], _062731_);
  or g_120424_(_062726_, _062731_, _062733_);
  or g_120425_(_062730_, _062733_, _062734_);
  or g_120426_(_062716_, _062723_, _062735_);
  or g_120427_(_062727_, _062735_, _062736_);
  or g_120428_(_062734_, _062736_, _062737_);
  or g_120429_(_062720_, _062737_, _062738_);
  xor g_120430_(out[428], out[620], _062739_);
  or g_120431_(_062724_, _062739_, _062740_);
  xor g_120432_(out[423], out[615], _062741_);
  or g_120433_(_062725_, _062741_, _062742_);
  or g_120434_(_062740_, _062742_, _062744_);
  or g_120435_(_062714_, _062715_, _062745_);
  or g_120436_(_062728_, _062745_, _062746_);
  or g_120437_(_062744_, _062746_, _062747_);
  or g_120438_(_062717_, _062747_, _062748_);
  or g_120439_(_062738_, _062748_, _062749_);
  not g_120440_(_062749_, _062750_);
  xor g_120441_(out[407], out[615], _062751_);
  and g_120442_(_049444_, out[619], _062752_);
  xor g_120443_(out[414], out[622], _062753_);
  xor g_120444_(out[408], out[616], _062755_);
  xor g_120445_(out[401], out[609], _062756_);
  xor g_120446_(out[413], out[621], _062757_);
  xor g_120447_(out[409], out[617], _062758_);
  xor g_120448_(out[404], out[612], _062759_);
  xor g_120449_(out[402], out[610], _062760_);
  and g_120450_(out[411], _049587_, _062761_);
  xor g_120451_(out[403], out[611], _062762_);
  xor g_120452_(out[406], out[614], _062763_);
  xor g_120453_(out[415], out[623], _062764_);
  xor g_120454_(out[410], out[618], _062766_);
  xor g_120455_(out[405], out[613], _062767_);
  xor g_120456_(out[400], out[608], _062768_);
  or g_120457_(_062753_, _062759_, _062769_);
  or g_120458_(_062755_, _062757_, _062770_);
  or g_120459_(_062760_, _062766_, _062771_);
  or g_120460_(_062770_, _062771_, _062772_);
  or g_120461_(_062758_, _062762_, _062773_);
  or g_120462_(_062767_, _062768_, _062774_);
  or g_120463_(_062773_, _062774_, _062775_);
  or g_120464_(_062772_, _062775_, _062777_);
  xor g_120465_(out[412], out[620], _062778_);
  or g_120466_(_062752_, _062778_, _062779_);
  or g_120467_(_062751_, _062763_, _062780_);
  or g_120468_(_062779_, _062780_, _062781_);
  or g_120469_(_062756_, _062761_, _062782_);
  or g_120470_(_062764_, _062782_, _062783_);
  or g_120471_(_062781_, _062783_, _062784_);
  or g_120472_(_062777_, _062784_, _062785_);
  or g_120473_(_062769_, _062785_, _062786_);
  and g_120474_(out[395], _049587_, _062788_);
  xor g_120475_(out[388], out[612], _062789_);
  xor g_120476_(out[387], out[611], _062790_);
  xor g_120477_(out[391], out[615], _062791_);
  xor g_120478_(out[398], out[622], _062792_);
  and g_120479_(_049433_, out[619], _062793_);
  xor g_120480_(out[397], out[621], _062794_);
  xor g_120481_(out[386], out[610], _062795_);
  xor g_120482_(out[393], out[617], _062796_);
  xor g_120483_(out[384], out[608], _062797_);
  xor g_120484_(out[392], out[616], _062799_);
  xor g_120485_(out[390], out[614], _062800_);
  xor g_120486_(out[389], out[613], _062801_);
  xor g_120487_(out[399], out[623], _062802_);
  xor g_120488_(out[394], out[618], _062803_);
  or g_120489_(_062794_, _062799_, _062804_);
  xor g_120490_(out[385], out[609], _062805_);
  or g_120491_(_062795_, _062803_, _062806_);
  or g_120492_(_062804_, _062806_, _062807_);
  or g_120493_(_062790_, _062796_, _062808_);
  or g_120494_(_062801_, _062808_, _062810_);
  or g_120495_(_062807_, _062810_, _062811_);
  or g_120496_(_062789_, _062792_, _062812_);
  or g_120497_(_062811_, _062812_, _062813_);
  xor g_120498_(out[396], out[620], _062814_);
  or g_120499_(_062793_, _062814_, _062815_);
  or g_120500_(_062791_, _062800_, _062816_);
  or g_120501_(_062815_, _062816_, _062817_);
  or g_120502_(_062788_, _062805_, _062818_);
  or g_120503_(_062802_, _062818_, _062819_);
  or g_120504_(_062817_, _062819_, _062821_);
  or g_120505_(_062797_, _062821_, _062822_);
  or g_120506_(_062813_, _062822_, _062823_);
  not g_120507_(_062823_, _062824_);
  xor g_120508_(out[375], out[615], _062825_);
  and g_120509_(_049422_, out[619], _062826_);
  xor g_120510_(out[382], out[622], _062827_);
  xor g_120511_(out[376], out[616], _062828_);
  xor g_120512_(out[369], out[609], _062829_);
  xor g_120513_(out[381], out[621], _062830_);
  xor g_120514_(out[377], out[617], _062832_);
  xor g_120515_(out[372], out[612], _062833_);
  xor g_120516_(out[370], out[610], _062834_);
  and g_120517_(out[379], _049587_, _062835_);
  xor g_120518_(out[371], out[611], _062836_);
  xor g_120519_(out[374], out[614], _062837_);
  xor g_120520_(out[383], out[623], _062838_);
  xor g_120521_(out[378], out[618], _062839_);
  xor g_120522_(out[373], out[613], _062840_);
  xor g_120523_(out[368], out[608], _062841_);
  or g_120524_(_062827_, _062833_, _062843_);
  or g_120525_(_062828_, _062830_, _062844_);
  or g_120526_(_062834_, _062839_, _062845_);
  or g_120527_(_062844_, _062845_, _062846_);
  or g_120528_(_062832_, _062836_, _062847_);
  or g_120529_(_062840_, _062841_, _062848_);
  or g_120530_(_062847_, _062848_, _062849_);
  or g_120531_(_062846_, _062849_, _062850_);
  xor g_120532_(out[380], out[620], _062851_);
  or g_120533_(_062826_, _062851_, _062852_);
  or g_120534_(_062825_, _062837_, _062854_);
  or g_120535_(_062852_, _062854_, _062855_);
  or g_120536_(_062829_, _062835_, _062856_);
  or g_120537_(_062838_, _062856_, _062857_);
  or g_120538_(_062855_, _062857_, _062858_);
  or g_120539_(_062850_, _062858_, _062859_);
  or g_120540_(_062843_, _062859_, _062860_);
  xor g_120541_(out[362], out[618], _062861_);
  xor g_120542_(out[360], out[616], _062862_);
  xor g_120543_(out[353], out[609], _062863_);
  and g_120544_(_049411_, out[619], _062865_);
  and g_120545_(out[363], _049587_, _062866_);
  xor g_120546_(out[354], out[610], _062867_);
  xor g_120547_(out[357], out[613], _062868_);
  xor g_120548_(out[361], out[617], _062869_);
  xor g_120549_(out[364], out[620], _062870_);
  xor g_120550_(out[365], out[621], _062871_);
  xor g_120551_(out[367], out[623], _062872_);
  xor g_120552_(out[356], out[612], _062873_);
  xor g_120553_(out[358], out[614], _062874_);
  xor g_120554_(out[355], out[611], _062876_);
  xor g_120555_(out[352], out[608], _062877_);
  xor g_120556_(out[366], out[622], _062878_);
  or g_120557_(_062873_, _062878_, _062879_);
  or g_120558_(_062862_, _062871_, _062880_);
  or g_120559_(_062861_, _062867_, _062881_);
  or g_120560_(_062880_, _062881_, _062882_);
  or g_120561_(_062869_, _062876_, _062883_);
  or g_120562_(_062868_, _062877_, _062884_);
  or g_120563_(_062883_, _062884_, _062885_);
  or g_120564_(_062882_, _062885_, _062887_);
  or g_120565_(_062865_, _062870_, _062888_);
  xor g_120566_(out[359], out[615], _062889_);
  or g_120567_(_062874_, _062889_, _062890_);
  or g_120568_(_062888_, _062890_, _062891_);
  or g_120569_(_062863_, _062866_, _062892_);
  or g_120570_(_062872_, _062892_, _062893_);
  or g_120571_(_062891_, _062893_, _062894_);
  or g_120572_(_062887_, _062894_, _062895_);
  or g_120573_(_062879_, _062895_, _062896_);
  xor g_120574_(out[343], out[615], _062898_);
  and g_120575_(_049400_, out[619], _062899_);
  xor g_120576_(out[350], out[622], _062900_);
  xor g_120577_(out[344], out[616], _062901_);
  xor g_120578_(out[337], out[609], _062902_);
  xor g_120579_(out[349], out[621], _062903_);
  xor g_120580_(out[345], out[617], _062904_);
  xor g_120581_(out[340], out[612], _062905_);
  xor g_120582_(out[338], out[610], _062906_);
  and g_120583_(out[347], _049587_, _062907_);
  xor g_120584_(out[339], out[611], _062909_);
  xor g_120585_(out[342], out[614], _062910_);
  xor g_120586_(out[351], out[623], _062911_);
  xor g_120587_(out[346], out[618], _062912_);
  xor g_120588_(out[341], out[613], _062913_);
  xor g_120589_(out[336], out[608], _062914_);
  or g_120590_(_062900_, _062905_, _062915_);
  or g_120591_(_062901_, _062903_, _062916_);
  or g_120592_(_062906_, _062912_, _062917_);
  or g_120593_(_062916_, _062917_, _062918_);
  or g_120594_(_062904_, _062909_, _062920_);
  or g_120595_(_062913_, _062914_, _062921_);
  or g_120596_(_062920_, _062921_, _062922_);
  or g_120597_(_062918_, _062922_, _062923_);
  xor g_120598_(out[348], out[620], _062924_);
  or g_120599_(_062899_, _062924_, _062925_);
  or g_120600_(_062898_, _062910_, _062926_);
  or g_120601_(_062925_, _062926_, _062927_);
  or g_120602_(_062902_, _062907_, _062928_);
  or g_120603_(_062911_, _062928_, _062929_);
  or g_120604_(_062927_, _062929_, _062931_);
  or g_120605_(_062923_, _062931_, _062932_);
  or g_120606_(_062915_, _062932_, _062933_);
  xor g_120607_(out[332], out[620], _062934_);
  and g_120608_(_098294_, out[619], _062935_);
  xor g_120609_(out[328], out[616], _062936_);
  xor g_120610_(out[326], out[614], _062937_);
  xor g_120611_(out[333], out[621], _062938_);
  xor g_120612_(out[334], out[622], _062939_);
  xor g_120613_(out[322], out[610], _062940_);
  xor g_120614_(out[329], out[617], _062942_);
  xor g_120615_(out[325], out[613], _062943_);
  xor g_120616_(out[321], out[609], _062944_);
  and g_120617_(out[331], _049587_, _062945_);
  or g_120618_(_062936_, _062938_, _062946_);
  xor g_120619_(out[335], out[623], _062947_);
  xor g_120620_(out[330], out[618], _062948_);
  xor g_120621_(out[324], out[612], _062949_);
  xor g_120622_(out[323], out[611], _062950_);
  xor g_120623_(out[320], out[608], _062951_);
  or g_120624_(_062940_, _062948_, _062953_);
  or g_120625_(_062946_, _062953_, _062954_);
  or g_120626_(_062942_, _062950_, _062955_);
  or g_120627_(_062943_, _062955_, _062956_);
  or g_120628_(_062954_, _062956_, _062957_);
  or g_120629_(_062939_, _062949_, _062958_);
  or g_120630_(_062957_, _062958_, _062959_);
  or g_120631_(_062934_, _062935_, _062960_);
  xor g_120632_(out[327], out[615], _062961_);
  or g_120633_(_062937_, _062961_, _062962_);
  or g_120634_(_062960_, _062962_, _062964_);
  or g_120635_(_062944_, _062945_, _062965_);
  or g_120636_(_062947_, _062965_, _062966_);
  or g_120637_(_062964_, _062966_, _062967_);
  or g_120638_(_062951_, _062967_, _062968_);
  or g_120639_(_062959_, _062968_, _062969_);
  xor g_120640_(out[311], out[615], _062970_);
  and g_120641_(_098283_, out[619], _062971_);
  xor g_120642_(out[318], out[622], _062972_);
  xor g_120643_(out[312], out[616], _062973_);
  xor g_120644_(out[305], out[609], _062975_);
  xor g_120645_(out[317], out[621], _062976_);
  xor g_120646_(out[313], out[617], _062977_);
  xor g_120647_(out[308], out[612], _062978_);
  xor g_120648_(out[306], out[610], _062979_);
  and g_120649_(out[315], _049587_, _062980_);
  xor g_120650_(out[307], out[611], _062981_);
  xor g_120651_(out[310], out[614], _062982_);
  xor g_120652_(out[319], out[623], _062983_);
  xor g_120653_(out[314], out[618], _062984_);
  xor g_120654_(out[309], out[613], _062986_);
  xor g_120655_(out[304], out[608], _062987_);
  or g_120656_(_062972_, _062978_, _062988_);
  or g_120657_(_062973_, _062976_, _062989_);
  or g_120658_(_062979_, _062984_, _062990_);
  or g_120659_(_062989_, _062990_, _062991_);
  or g_120660_(_062977_, _062981_, _062992_);
  or g_120661_(_062986_, _062987_, _062993_);
  or g_120662_(_062992_, _062993_, _062994_);
  or g_120663_(_062991_, _062994_, _062995_);
  xor g_120664_(out[316], out[620], _062997_);
  or g_120665_(_062971_, _062997_, _062998_);
  or g_120666_(_062970_, _062982_, _062999_);
  or g_120667_(_062998_, _062999_, _063000_);
  or g_120668_(_062975_, _062980_, _063001_);
  or g_120669_(_062983_, _063001_, _063002_);
  or g_120670_(_063000_, _063002_, _063003_);
  or g_120671_(_062995_, _063003_, _063004_);
  or g_120672_(_062988_, _063004_, _063005_);
  not g_120673_(_063005_, _063006_);
  xor g_120674_(out[289], out[609], _063008_);
  and g_120675_(out[299], _049587_, _063009_);
  xor g_120676_(out[302], out[622], _063010_);
  xor g_120677_(out[291], out[611], _063011_);
  xor g_120678_(out[292], out[612], _063012_);
  xor g_120679_(out[290], out[610], _063013_);
  xor g_120680_(out[297], out[617], _063014_);
  xor g_120681_(out[288], out[608], _063015_);
  and g_120682_(_098272_, out[619], _063016_);
  xor g_120683_(out[294], out[614], _063017_);
  xor g_120684_(out[298], out[618], _063019_);
  xor g_120685_(out[293], out[613], _063020_);
  xor g_120686_(out[303], out[623], _063021_);
  xor g_120687_(out[301], out[621], _063022_);
  xor g_120688_(out[296], out[616], _063023_);
  or g_120689_(_063010_, _063012_, _063024_);
  or g_120690_(_063022_, _063023_, _063025_);
  or g_120691_(_063013_, _063019_, _063026_);
  or g_120692_(_063025_, _063026_, _063027_);
  or g_120693_(_063011_, _063014_, _063028_);
  or g_120694_(_063015_, _063020_, _063030_);
  or g_120695_(_063028_, _063030_, _063031_);
  or g_120696_(_063027_, _063031_, _063032_);
  xor g_120697_(out[300], out[620], _063033_);
  or g_120698_(_063016_, _063033_, _063034_);
  xor g_120699_(out[295], out[615], _063035_);
  or g_120700_(_063017_, _063035_, _063036_);
  or g_120701_(_063034_, _063036_, _063037_);
  or g_120702_(_063008_, _063009_, _063038_);
  or g_120703_(_063021_, _063038_, _063039_);
  or g_120704_(_063037_, _063039_, _063041_);
  or g_120705_(_063032_, _063041_, _063042_);
  or g_120706_(_063024_, _063042_, _063043_);
  xor g_120707_(out[279], out[615], _063044_);
  and g_120708_(_098261_, out[619], _063045_);
  xor g_120709_(out[286], out[622], _063046_);
  xor g_120710_(out[280], out[616], _063047_);
  xor g_120711_(out[273], out[609], _063048_);
  xor g_120712_(out[285], out[621], _063049_);
  xor g_120713_(out[281], out[617], _063050_);
  xor g_120714_(out[276], out[612], _063052_);
  xor g_120715_(out[274], out[610], _063053_);
  and g_120716_(out[283], _049587_, _063054_);
  xor g_120717_(out[275], out[611], _063055_);
  xor g_120718_(out[278], out[614], _063056_);
  xor g_120719_(out[287], out[623], _063057_);
  xor g_120720_(out[282], out[618], _063058_);
  xor g_120721_(out[277], out[613], _063059_);
  xor g_120722_(out[272], out[608], _063060_);
  or g_120723_(_063046_, _063052_, _063061_);
  or g_120724_(_063047_, _063049_, _063063_);
  or g_120725_(_063053_, _063058_, _063064_);
  or g_120726_(_063063_, _063064_, _063065_);
  or g_120727_(_063050_, _063055_, _063066_);
  or g_120728_(_063059_, _063060_, _063067_);
  or g_120729_(_063066_, _063067_, _063068_);
  or g_120730_(_063065_, _063068_, _063069_);
  xor g_120731_(out[284], out[620], _063070_);
  or g_120732_(_063045_, _063070_, _063071_);
  or g_120733_(_063044_, _063056_, _063072_);
  or g_120734_(_063071_, _063072_, _063074_);
  or g_120735_(_063048_, _063054_, _063075_);
  or g_120736_(_063057_, _063075_, _063076_);
  or g_120737_(_063074_, _063076_, _063077_);
  or g_120738_(_063069_, _063077_, _063078_);
  or g_120739_(_063061_, _063078_, _063079_);
  xor g_120740_(out[259], out[611], _063080_);
  xor g_120741_(out[260], out[612], _063081_);
  xor g_120742_(out[270], out[622], _063082_);
  xor g_120743_(out[258], out[610], _063083_);
  xor g_120744_(out[261], out[613], _063085_);
  xor g_120745_(out[265], out[617], _063086_);
  xor g_120746_(out[264], out[616], _063087_);
  xor g_120747_(out[271], out[623], _063088_);
  xor g_120748_(out[266], out[618], _063089_);
  xor g_120749_(out[262], out[614], _063090_);
  xor g_120750_(out[256], out[608], _063091_);
  and g_120751_(_098250_, out[619], _063092_);
  and g_120752_(out[267], _049587_, _063093_);
  xor g_120753_(out[269], out[621], _063094_);
  or g_120754_(_063087_, _063094_, _063096_);
  xor g_120755_(out[257], out[609], _063097_);
  or g_120756_(_063083_, _063089_, _063098_);
  or g_120757_(_063096_, _063098_, _063099_);
  or g_120758_(_063080_, _063086_, _063100_);
  or g_120759_(_063085_, _063100_, _063101_);
  or g_120760_(_063099_, _063101_, _063102_);
  or g_120761_(_063081_, _063082_, _063103_);
  or g_120762_(_063102_, _063103_, _063104_);
  xor g_120763_(out[268], out[620], _063105_);
  or g_120764_(_063092_, _063105_, _063107_);
  xor g_120765_(out[263], out[615], _063108_);
  or g_120766_(_063090_, _063108_, _063109_);
  or g_120767_(_063107_, _063109_, _063110_);
  or g_120768_(_063093_, _063097_, _063111_);
  or g_120769_(_063088_, _063111_, _063112_);
  or g_120770_(_063110_, _063112_, _063113_);
  or g_120771_(_063091_, _063113_, _063114_);
  or g_120772_(_063104_, _063114_, _063115_);
  not g_120773_(_063115_, _063116_);
  xor g_120774_(out[247], out[615], _063118_);
  and g_120775_(_098239_, out[619], _063119_);
  xor g_120776_(out[254], out[622], _063120_);
  xor g_120777_(out[248], out[616], _063121_);
  xor g_120778_(out[241], out[609], _063122_);
  xor g_120779_(out[253], out[621], _063123_);
  xor g_120780_(out[249], out[617], _063124_);
  xor g_120781_(out[244], out[612], _063125_);
  xor g_120782_(out[242], out[610], _063126_);
  and g_120783_(out[251], _049587_, _063127_);
  xor g_120784_(out[243], out[611], _063129_);
  xor g_120785_(out[246], out[614], _063130_);
  xor g_120786_(out[255], out[623], _063131_);
  xor g_120787_(out[250], out[618], _063132_);
  xor g_120788_(out[245], out[613], _063133_);
  xor g_120789_(out[240], out[608], _063134_);
  or g_120790_(_063120_, _063125_, _063135_);
  or g_120791_(_063121_, _063123_, _063136_);
  or g_120792_(_063126_, _063132_, _063137_);
  or g_120793_(_063136_, _063137_, _063138_);
  or g_120794_(_063124_, _063129_, _063140_);
  or g_120795_(_063133_, _063134_, _063141_);
  or g_120796_(_063140_, _063141_, _063142_);
  or g_120797_(_063138_, _063142_, _063143_);
  xor g_120798_(out[252], out[620], _063144_);
  or g_120799_(_063119_, _063144_, _063145_);
  or g_120800_(_063118_, _063130_, _063146_);
  or g_120801_(_063145_, _063146_, _063147_);
  or g_120802_(_063122_, _063127_, _063148_);
  or g_120803_(_063131_, _063148_, _063149_);
  or g_120804_(_063147_, _063149_, _063151_);
  or g_120805_(_063143_, _063151_, _063152_);
  or g_120806_(_063135_, _063152_, _063153_);
  not g_120807_(_063153_, _063154_);
  xor g_120808_(out[234], out[618], _063155_);
  xor g_120809_(out[226], out[610], _063156_);
  xor g_120810_(out[225], out[609], _063157_);
  and g_120811_(_098228_, out[619], _063158_);
  and g_120812_(out[235], _049587_, _063159_);
  xor g_120813_(out[237], out[621], _063160_);
  xor g_120814_(out[227], out[611], _063162_);
  xor g_120815_(out[238], out[622], _063163_);
  xor g_120816_(out[236], out[620], _063164_);
  xor g_120817_(out[232], out[616], _063165_);
  xor g_120818_(out[239], out[623], _063166_);
  xor g_120819_(out[229], out[613], _063167_);
  xor g_120820_(out[230], out[614], _063168_);
  xor g_120821_(out[224], out[608], _063169_);
  xor g_120822_(out[228], out[612], _063170_);
  or g_120823_(_063160_, _063165_, _063171_);
  xor g_120824_(out[233], out[617], _063173_);
  or g_120825_(_063155_, _063156_, _063174_);
  or g_120826_(_063171_, _063174_, _063175_);
  or g_120827_(_063162_, _063173_, _063176_);
  or g_120828_(_063167_, _063176_, _063177_);
  or g_120829_(_063175_, _063177_, _063178_);
  or g_120830_(_063163_, _063170_, _063179_);
  or g_120831_(_063178_, _063179_, _063180_);
  not g_120832_(_063180_, _063181_);
  or g_120833_(_063158_, _063164_, _063182_);
  xor g_120834_(out[231], out[615], _063184_);
  or g_120835_(_063168_, _063184_, _063185_);
  or g_120836_(_063182_, _063185_, _063186_);
  or g_120837_(_063157_, _063159_, _063187_);
  or g_120838_(_063166_, _063187_, _063188_);
  or g_120839_(_063186_, _063188_, _063189_);
  or g_120840_(_063169_, _063189_, _063190_);
  not g_120841_(_063190_, _063191_);
  and g_120842_(_063181_, _063191_, _063192_);
  or g_120843_(_063180_, _063190_, _063193_);
  xor g_120844_(out[215], out[615], _063195_);
  and g_120845_(_098217_, out[619], _063196_);
  xor g_120846_(out[222], out[622], _063197_);
  xor g_120847_(out[216], out[616], _063198_);
  xor g_120848_(out[209], out[609], _063199_);
  xor g_120849_(out[221], out[621], _063200_);
  xor g_120850_(out[217], out[617], _063201_);
  xor g_120851_(out[212], out[612], _063202_);
  xor g_120852_(out[210], out[610], _063203_);
  and g_120853_(out[219], _049587_, _063204_);
  xor g_120854_(out[211], out[611], _063206_);
  xor g_120855_(out[214], out[614], _063207_);
  xor g_120856_(out[223], out[623], _063208_);
  xor g_120857_(out[218], out[618], _063209_);
  xor g_120858_(out[213], out[613], _063210_);
  xor g_120859_(out[208], out[608], _063211_);
  or g_120860_(_063197_, _063202_, _063212_);
  or g_120861_(_063198_, _063200_, _063213_);
  or g_120862_(_063203_, _063209_, _063214_);
  or g_120863_(_063213_, _063214_, _063215_);
  or g_120864_(_063201_, _063206_, _063217_);
  or g_120865_(_063210_, _063211_, _063218_);
  or g_120866_(_063217_, _063218_, _063219_);
  or g_120867_(_063215_, _063219_, _063220_);
  xor g_120868_(out[220], out[620], _063221_);
  or g_120869_(_063196_, _063221_, _063222_);
  or g_120870_(_063195_, _063207_, _063223_);
  or g_120871_(_063222_, _063223_, _063224_);
  or g_120872_(_063199_, _063204_, _063225_);
  or g_120873_(_063208_, _063225_, _063226_);
  or g_120874_(_063224_, _063226_, _063228_);
  or g_120875_(_063220_, _063228_, _063229_);
  or g_120876_(_063212_, _063229_, _063230_);
  xor g_120877_(out[200], out[616], _063231_);
  xor g_120878_(out[197], out[613], _063232_);
  xor g_120879_(out[195], out[611], _063233_);
  xor g_120880_(out[206], out[622], _063234_);
  xor g_120881_(out[205], out[621], _063235_);
  xor g_120882_(out[194], out[610], _063236_);
  xor g_120883_(out[201], out[617], _063237_);
  xor g_120884_(out[198], out[614], _063239_);
  xor g_120885_(out[207], out[623], _063240_);
  xor g_120886_(out[202], out[618], _063241_);
  xor g_120887_(out[196], out[612], _063242_);
  xor g_120888_(out[192], out[608], _063243_);
  and g_120889_(_098206_, out[619], _063244_);
  and g_120890_(out[203], _049587_, _063245_);
  or g_120891_(_063231_, _063235_, _063246_);
  xor g_120892_(out[193], out[609], _063247_);
  or g_120893_(_063236_, _063241_, _063248_);
  or g_120894_(_063246_, _063248_, _063250_);
  or g_120895_(_063233_, _063237_, _063251_);
  or g_120896_(_063232_, _063251_, _063252_);
  or g_120897_(_063250_, _063252_, _063253_);
  or g_120898_(_063234_, _063242_, _063254_);
  or g_120899_(_063253_, _063254_, _063255_);
  xor g_120900_(out[204], out[620], _063256_);
  or g_120901_(_063244_, _063256_, _063257_);
  xor g_120902_(out[199], out[615], _063258_);
  or g_120903_(_063239_, _063258_, _063259_);
  or g_120904_(_063257_, _063259_, _063261_);
  or g_120905_(_063245_, _063247_, _063262_);
  or g_120906_(_063240_, _063262_, _063263_);
  or g_120907_(_063261_, _063263_, _063264_);
  or g_120908_(_063243_, _063264_, _063265_);
  or g_120909_(_063255_, _063265_, _063266_);
  xor g_120910_(out[183], out[615], _063267_);
  and g_120911_(_098195_, out[619], _063268_);
  xor g_120912_(out[190], out[622], _063269_);
  xor g_120913_(out[184], out[616], _063270_);
  xor g_120914_(out[177], out[609], _063272_);
  xor g_120915_(out[189], out[621], _063273_);
  xor g_120916_(out[185], out[617], _063274_);
  xor g_120917_(out[180], out[612], _063275_);
  xor g_120918_(out[178], out[610], _063276_);
  and g_120919_(out[187], _049587_, _063277_);
  xor g_120920_(out[179], out[611], _063278_);
  xor g_120921_(out[182], out[614], _063279_);
  xor g_120922_(out[191], out[623], _063280_);
  xor g_120923_(out[186], out[618], _063281_);
  xor g_120924_(out[181], out[613], _063283_);
  xor g_120925_(out[176], out[608], _063284_);
  or g_120926_(_063269_, _063275_, _063285_);
  or g_120927_(_063270_, _063273_, _063286_);
  or g_120928_(_063276_, _063281_, _063287_);
  or g_120929_(_063286_, _063287_, _063288_);
  or g_120930_(_063274_, _063278_, _063289_);
  or g_120931_(_063283_, _063284_, _063290_);
  or g_120932_(_063289_, _063290_, _063291_);
  or g_120933_(_063288_, _063291_, _063292_);
  xor g_120934_(out[188], out[620], _063294_);
  or g_120935_(_063268_, _063294_, _063295_);
  or g_120936_(_063267_, _063279_, _063296_);
  or g_120937_(_063295_, _063296_, _063297_);
  or g_120938_(_063272_, _063277_, _063298_);
  or g_120939_(_063280_, _063298_, _063299_);
  or g_120940_(_063297_, _063299_, _063300_);
  or g_120941_(_063292_, _063300_, _063301_);
  or g_120942_(_063285_, _063301_, _063302_);
  not g_120943_(_063302_, _063303_);
  and g_120944_(out[171], _049587_, _063305_);
  xor g_120945_(out[164], out[612], _063306_);
  xor g_120946_(out[162], out[610], _063307_);
  xor g_120947_(out[169], out[617], _063308_);
  xor g_120948_(out[160], out[608], _063309_);
  xor g_120949_(out[163], out[611], _063310_);
  and g_120950_(_098184_, out[619], _063311_);
  xor g_120951_(out[170], out[618], _063312_);
  xor g_120952_(out[175], out[623], _063313_);
  xor g_120953_(out[166], out[614], _063314_);
  xor g_120954_(out[165], out[613], _063316_);
  xor g_120955_(out[173], out[621], _063317_);
  xor g_120956_(out[174], out[622], _063318_);
  xor g_120957_(out[168], out[616], _063319_);
  xor g_120958_(out[161], out[609], _063320_);
  or g_120959_(_063306_, _063318_, _063321_);
  or g_120960_(_063317_, _063319_, _063322_);
  or g_120961_(_063307_, _063312_, _063323_);
  or g_120962_(_063322_, _063323_, _063324_);
  or g_120963_(_063308_, _063310_, _063325_);
  or g_120964_(_063309_, _063316_, _063327_);
  or g_120965_(_063325_, _063327_, _063328_);
  or g_120966_(_063324_, _063328_, _063329_);
  xor g_120967_(out[172], out[620], _063330_);
  or g_120968_(_063311_, _063330_, _063331_);
  xor g_120969_(out[167], out[615], _063332_);
  or g_120970_(_063314_, _063332_, _063333_);
  or g_120971_(_063331_, _063333_, _063334_);
  or g_120972_(_063305_, _063320_, _063335_);
  or g_120973_(_063313_, _063335_, _063336_);
  or g_120974_(_063334_, _063336_, _063338_);
  or g_120975_(_063329_, _063338_, _063339_);
  or g_120976_(_063321_, _063339_, _063340_);
  xor g_120977_(out[151], out[615], _063341_);
  and g_120978_(_098173_, out[619], _063342_);
  xor g_120979_(out[158], out[622], _063343_);
  xor g_120980_(out[152], out[616], _063344_);
  xor g_120981_(out[145], out[609], _063345_);
  xor g_120982_(out[157], out[621], _063346_);
  xor g_120983_(out[153], out[617], _063347_);
  xor g_120984_(out[148], out[612], _063349_);
  xor g_120985_(out[146], out[610], _063350_);
  and g_120986_(out[155], _049587_, _063351_);
  xor g_120987_(out[147], out[611], _063352_);
  xor g_120988_(out[150], out[614], _063353_);
  xor g_120989_(out[159], out[623], _063354_);
  xor g_120990_(out[154], out[618], _063355_);
  xor g_120991_(out[149], out[613], _063356_);
  xor g_120992_(out[144], out[608], _063357_);
  or g_120993_(_063343_, _063349_, _063358_);
  or g_120994_(_063344_, _063346_, _063360_);
  or g_120995_(_063350_, _063355_, _063361_);
  or g_120996_(_063360_, _063361_, _063362_);
  or g_120997_(_063347_, _063352_, _063363_);
  or g_120998_(_063356_, _063357_, _063364_);
  or g_120999_(_063363_, _063364_, _063365_);
  or g_121000_(_063362_, _063365_, _063366_);
  xor g_121001_(out[156], out[620], _063367_);
  or g_121002_(_063342_, _063367_, _063368_);
  or g_121003_(_063341_, _063353_, _063369_);
  or g_121004_(_063368_, _063369_, _063371_);
  or g_121005_(_063345_, _063351_, _063372_);
  or g_121006_(_063354_, _063372_, _063373_);
  or g_121007_(_063371_, _063373_, _063374_);
  or g_121008_(_063366_, _063374_, _063375_);
  or g_121009_(_063358_, _063375_, _063376_);
  and g_121010_(out[139], _049587_, _063377_);
  xor g_121011_(out[132], out[612], _063378_);
  xor g_121012_(out[142], out[622], _063379_);
  or g_121013_(_063378_, _063379_, _063380_);
  xor g_121014_(out[141], out[621], _063382_);
  xor g_121015_(out[131], out[611], _063383_);
  xor g_121016_(out[128], out[608], _063384_);
  and g_121017_(_098162_, out[619], _063385_);
  xor g_121018_(out[138], out[618], _063386_);
  xor g_121019_(out[143], out[623], _063387_);
  xor g_121020_(out[134], out[614], _063388_);
  xor g_121021_(out[133], out[613], _063389_);
  xor g_121022_(out[136], out[616], _063390_);
  or g_121023_(_063382_, _063390_, _063391_);
  xor g_121024_(out[130], out[610], _063393_);
  xor g_121025_(out[137], out[617], _063394_);
  xor g_121026_(out[129], out[609], _063395_);
  or g_121027_(_063386_, _063393_, _063396_);
  or g_121028_(_063391_, _063396_, _063397_);
  or g_121029_(_063383_, _063394_, _063398_);
  or g_121030_(_063389_, _063398_, _063399_);
  or g_121031_(_063397_, _063399_, _063400_);
  or g_121032_(_063380_, _063400_, _063401_);
  xor g_121033_(out[140], out[620], _063402_);
  or g_121034_(_063385_, _063402_, _063404_);
  xor g_121035_(out[135], out[615], _063405_);
  or g_121036_(_063388_, _063405_, _063406_);
  or g_121037_(_063404_, _063406_, _063407_);
  or g_121038_(_063377_, _063395_, _063408_);
  or g_121039_(_063387_, _063408_, _063409_);
  or g_121040_(_063407_, _063409_, _063410_);
  or g_121041_(_063384_, _063410_, _063411_);
  or g_121042_(_063401_, _063411_, _063412_);
  xor g_121043_(out[119], out[615], _063413_);
  and g_121044_(_098151_, out[619], _063415_);
  xor g_121045_(out[126], out[622], _063416_);
  xor g_121046_(out[120], out[616], _063417_);
  xor g_121047_(out[113], out[609], _063418_);
  xor g_121048_(out[125], out[621], _063419_);
  xor g_121049_(out[121], out[617], _063420_);
  xor g_121050_(out[116], out[612], _063421_);
  xor g_121051_(out[114], out[610], _063422_);
  and g_121052_(out[123], _049587_, _063423_);
  xor g_121053_(out[115], out[611], _063424_);
  xor g_121054_(out[118], out[614], _063426_);
  xor g_121055_(out[127], out[623], _063427_);
  xor g_121056_(out[122], out[618], _063428_);
  xor g_121057_(out[117], out[613], _063429_);
  xor g_121058_(out[112], out[608], _063430_);
  or g_121059_(_063416_, _063421_, _063431_);
  or g_121060_(_063417_, _063419_, _063432_);
  or g_121061_(_063422_, _063428_, _063433_);
  or g_121062_(_063432_, _063433_, _063434_);
  or g_121063_(_063420_, _063424_, _063435_);
  or g_121064_(_063429_, _063430_, _063437_);
  or g_121065_(_063435_, _063437_, _063438_);
  or g_121066_(_063434_, _063438_, _063439_);
  xor g_121067_(out[124], out[620], _063440_);
  or g_121068_(_063415_, _063440_, _063441_);
  or g_121069_(_063413_, _063426_, _063442_);
  or g_121070_(_063441_, _063442_, _063443_);
  or g_121071_(_063418_, _063423_, _063444_);
  or g_121072_(_063427_, _063444_, _063445_);
  or g_121073_(_063443_, _063445_, _063446_);
  or g_121074_(_063439_, _063446_, _063448_);
  or g_121075_(_063431_, _063448_, _063449_);
  xor g_121076_(out[97], out[609], _063450_);
  and g_121077_(_098140_, out[619], _063451_);
  and g_121078_(out[107], _049587_, _063452_);
  xor g_121079_(out[105], out[617], _063453_);
  xor g_121080_(out[96], out[608], _063454_);
  xor g_121081_(out[110], out[622], _063455_);
  xor g_121082_(out[100], out[612], _063456_);
  or g_121083_(_063455_, _063456_, _063457_);
  xor g_121084_(out[109], out[621], _063459_);
  xor g_121085_(out[99], out[611], _063460_);
  xor g_121086_(out[108], out[620], _063461_);
  xor g_121087_(out[102], out[614], _063462_);
  xor g_121088_(out[106], out[618], _063463_);
  xor g_121089_(out[101], out[613], _063464_);
  xor g_121090_(out[111], out[623], _063465_);
  xor g_121091_(out[104], out[616], _063466_);
  or g_121092_(_063459_, _063466_, _063467_);
  xor g_121093_(out[98], out[610], _063468_);
  or g_121094_(_063463_, _063468_, _063470_);
  or g_121095_(_063467_, _063470_, _063471_);
  or g_121096_(_063453_, _063460_, _063472_);
  or g_121097_(_063464_, _063472_, _063473_);
  or g_121098_(_063471_, _063473_, _063474_);
  or g_121099_(_063457_, _063474_, _063475_);
  or g_121100_(_063451_, _063461_, _063476_);
  xor g_121101_(out[103], out[615], _063477_);
  or g_121102_(_063462_, _063477_, _063478_);
  or g_121103_(_063476_, _063478_, _063479_);
  or g_121104_(_063450_, _063452_, _063481_);
  or g_121105_(_063465_, _063481_, _063482_);
  or g_121106_(_063479_, _063482_, _063483_);
  or g_121107_(_063454_, _063483_, _063484_);
  or g_121108_(_063475_, _063484_, _063485_);
  not g_121109_(_063485_, _063486_);
  xor g_121110_(out[87], out[615], _063487_);
  and g_121111_(_098129_, out[619], _063488_);
  xor g_121112_(out[94], out[622], _063489_);
  xor g_121113_(out[88], out[616], _063490_);
  xor g_121114_(out[81], out[609], _063492_);
  xor g_121115_(out[93], out[621], _063493_);
  xor g_121116_(out[89], out[617], _063494_);
  xor g_121117_(out[84], out[612], _063495_);
  xor g_121118_(out[82], out[610], _063496_);
  and g_121119_(out[91], _049587_, _063497_);
  xor g_121120_(out[83], out[611], _063498_);
  xor g_121121_(out[86], out[614], _063499_);
  xor g_121122_(out[95], out[623], _063500_);
  xor g_121123_(out[90], out[618], _063501_);
  xor g_121124_(out[85], out[613], _063503_);
  xor g_121125_(out[80], out[608], _063504_);
  or g_121126_(_063489_, _063495_, _063505_);
  or g_121127_(_063490_, _063493_, _063506_);
  or g_121128_(_063496_, _063501_, _063507_);
  or g_121129_(_063506_, _063507_, _063508_);
  or g_121130_(_063494_, _063498_, _063509_);
  or g_121131_(_063503_, _063504_, _063510_);
  or g_121132_(_063509_, _063510_, _063511_);
  or g_121133_(_063508_, _063511_, _063512_);
  xor g_121134_(out[92], out[620], _063514_);
  or g_121135_(_063488_, _063514_, _063515_);
  or g_121136_(_063487_, _063499_, _063516_);
  or g_121137_(_063515_, _063516_, _063517_);
  or g_121138_(_063492_, _063497_, _063518_);
  or g_121139_(_063500_, _063518_, _063519_);
  or g_121140_(_063517_, _063519_, _063520_);
  or g_121141_(_063512_, _063520_, _063521_);
  or g_121142_(_063505_, _063521_, _063522_);
  not g_121143_(_063522_, _063523_);
  xor g_121144_(out[65], out[609], _063525_);
  and g_121145_(out[75], _049587_, _063526_);
  xor g_121146_(out[78], out[622], _063527_);
  xor g_121147_(out[67], out[611], _063528_);
  xor g_121148_(out[68], out[612], _063529_);
  xor g_121149_(out[66], out[610], _063530_);
  xor g_121150_(out[73], out[617], _063531_);
  xor g_121151_(out[64], out[608], _063532_);
  and g_121152_(_098118_, out[619], _063533_);
  xor g_121153_(out[70], out[614], _063534_);
  xor g_121154_(out[74], out[618], _063536_);
  xor g_121155_(out[69], out[613], _063537_);
  xor g_121156_(out[79], out[623], _063538_);
  xor g_121157_(out[77], out[621], _063539_);
  xor g_121158_(out[72], out[616], _063540_);
  or g_121159_(_063527_, _063529_, _063541_);
  or g_121160_(_063539_, _063540_, _063542_);
  or g_121161_(_063530_, _063536_, _063543_);
  or g_121162_(_063542_, _063543_, _063544_);
  or g_121163_(_063528_, _063531_, _063545_);
  or g_121164_(_063532_, _063537_, _063547_);
  or g_121165_(_063545_, _063547_, _063548_);
  or g_121166_(_063544_, _063548_, _063549_);
  xor g_121167_(out[76], out[620], _063550_);
  or g_121168_(_063533_, _063550_, _063551_);
  xor g_121169_(out[71], out[615], _063552_);
  or g_121170_(_063534_, _063552_, _063553_);
  or g_121171_(_063551_, _063553_, _063554_);
  or g_121172_(_063525_, _063526_, _063555_);
  or g_121173_(_063538_, _063555_, _063556_);
  or g_121174_(_063554_, _063556_, _063558_);
  or g_121175_(_063549_, _063558_, _063559_);
  or g_121176_(_063541_, _063559_, _063560_);
  xor g_121177_(out[55], out[615], _063561_);
  and g_121178_(_098107_, out[619], _063562_);
  xor g_121179_(out[62], out[622], _063563_);
  xor g_121180_(out[56], out[616], _063564_);
  xor g_121181_(out[49], out[609], _063565_);
  xor g_121182_(out[61], out[621], _063566_);
  xor g_121183_(out[57], out[617], _063567_);
  xor g_121184_(out[52], out[612], _063569_);
  xor g_121185_(out[50], out[610], _063570_);
  and g_121186_(out[59], _049587_, _063571_);
  xor g_121187_(out[51], out[611], _063572_);
  xor g_121188_(out[54], out[614], _063573_);
  xor g_121189_(out[63], out[623], _063574_);
  xor g_121190_(out[58], out[618], _063575_);
  xor g_121191_(out[53], out[613], _063576_);
  xor g_121192_(out[48], out[608], _063577_);
  or g_121193_(_063563_, _063569_, _063578_);
  or g_121194_(_063564_, _063566_, _063580_);
  or g_121195_(_063570_, _063575_, _063581_);
  or g_121196_(_063580_, _063581_, _063582_);
  or g_121197_(_063567_, _063572_, _063583_);
  or g_121198_(_063576_, _063577_, _063584_);
  or g_121199_(_063583_, _063584_, _063585_);
  or g_121200_(_063582_, _063585_, _063586_);
  xor g_121201_(out[60], out[620], _063587_);
  or g_121202_(_063562_, _063587_, _063588_);
  or g_121203_(_063561_, _063573_, _063589_);
  or g_121204_(_063588_, _063589_, _063591_);
  or g_121205_(_063565_, _063571_, _063592_);
  or g_121206_(_063574_, _063592_, _063593_);
  or g_121207_(_063591_, _063593_, _063594_);
  or g_121208_(_063586_, _063594_, _063595_);
  or g_121209_(_063578_, _063595_, _063596_);
  and g_121210_(out[43], _049587_, _063597_);
  and g_121211_(_098096_, out[619], _063598_);
  xor g_121212_(out[40], out[616], _063599_);
  xor g_121213_(out[47], out[623], _063600_);
  xor g_121214_(out[33], out[609], _063602_);
  xor g_121215_(out[34], out[610], _063603_);
  xor g_121216_(out[36], out[612], _063604_);
  xor g_121217_(out[45], out[621], _063605_);
  xor g_121218_(out[41], out[617], _063606_);
  xor g_121219_(out[35], out[611], _063607_);
  xor g_121220_(out[37], out[613], _063608_);
  xor g_121221_(out[46], out[622], _063609_);
  xor g_121222_(out[32], out[608], _063610_);
  xor g_121223_(out[42], out[618], _063611_);
  or g_121224_(_063599_, _063605_, _063613_);
  xor g_121225_(out[38], out[614], _063614_);
  or g_121226_(_063603_, _063611_, _063615_);
  or g_121227_(_063613_, _063615_, _063616_);
  or g_121228_(_063606_, _063607_, _063617_);
  or g_121229_(_063608_, _063617_, _063618_);
  or g_121230_(_063616_, _063618_, _063619_);
  or g_121231_(_063604_, _063609_, _063620_);
  or g_121232_(_063619_, _063620_, _063621_);
  xor g_121233_(out[44], out[620], _063622_);
  or g_121234_(_063598_, _063622_, _063624_);
  xor g_121235_(out[39], out[615], _063625_);
  or g_121236_(_063614_, _063625_, _063626_);
  or g_121237_(_063624_, _063626_, _063627_);
  or g_121238_(_063597_, _063602_, _063628_);
  or g_121239_(_063600_, _063628_, _063629_);
  or g_121240_(_063627_, _063629_, _063630_);
  or g_121241_(_063610_, _063630_, _063631_);
  or g_121242_(_063621_, _063631_, _063632_);
  not g_121243_(_063632_, _063633_);
  xor g_121244_(out[23], out[615], _063635_);
  and g_121245_(_098063_, out[619], _063636_);
  xor g_121246_(out[30], out[622], _063637_);
  xor g_121247_(out[24], out[616], _063638_);
  xor g_121248_(out[17], out[609], _063639_);
  xor g_121249_(out[29], out[621], _063640_);
  xor g_121250_(out[25], out[617], _063641_);
  xor g_121251_(out[20], out[612], _063642_);
  xor g_121252_(out[18], out[610], _063643_);
  and g_121253_(out[27], _049587_, _063644_);
  xor g_121254_(out[19], out[611], _063646_);
  xor g_121255_(out[22], out[614], _063647_);
  xor g_121256_(out[31], out[623], _063648_);
  xor g_121257_(out[26], out[618], _063649_);
  xor g_121258_(out[21], out[613], _063650_);
  xor g_121259_(out[16], out[608], _063651_);
  or g_121260_(_063637_, _063642_, _063652_);
  or g_121261_(_063638_, _063640_, _063653_);
  or g_121262_(_063643_, _063649_, _063654_);
  or g_121263_(_063653_, _063654_, _063655_);
  or g_121264_(_063641_, _063646_, _063657_);
  or g_121265_(_063650_, _063651_, _063658_);
  or g_121266_(_063657_, _063658_, _063659_);
  or g_121267_(_063655_, _063659_, _063660_);
  xor g_121268_(out[28], out[620], _063661_);
  or g_121269_(_063636_, _063661_, _063662_);
  or g_121270_(_063635_, _063647_, _063663_);
  or g_121271_(_063662_, _063663_, _063664_);
  or g_121272_(_063639_, _063644_, _063665_);
  or g_121273_(_063648_, _063665_, _063666_);
  or g_121274_(_063664_, _063666_, _063668_);
  or g_121275_(_063660_, _063668_, _063669_);
  or g_121276_(_063652_, _063669_, _063670_);
  not g_121277_(_063670_, _063671_);
  xor g_121278_(out[1], out[609], _063672_);
  and g_121279_(out[11], _049587_, _063673_);
  xor g_121280_(out[9], out[617], _063674_);
  xor g_121281_(out[0], out[608], _063675_);
  xor g_121282_(out[14], out[622], _063676_);
  xor g_121283_(out[4], out[612], _063677_);
  or g_121284_(_063676_, _063677_, _063679_);
  xor g_121285_(out[13], out[621], _063680_);
  xor g_121286_(out[3], out[611], _063681_);
  and g_121287_(_098041_, out[619], _063682_);
  xor g_121288_(out[6], out[614], _063683_);
  xor g_121289_(out[10], out[618], _063684_);
  xor g_121290_(out[5], out[613], _063685_);
  xor g_121291_(out[15], out[623], _063686_);
  xor g_121292_(out[8], out[616], _063687_);
  or g_121293_(_063680_, _063687_, _063688_);
  xor g_121294_(out[2], out[610], _063690_);
  or g_121295_(_063684_, _063690_, _063691_);
  or g_121296_(_063688_, _063691_, _063692_);
  or g_121297_(_063674_, _063681_, _063693_);
  or g_121298_(_063685_, _063693_, _063694_);
  or g_121299_(_063692_, _063694_, _063695_);
  or g_121300_(_063679_, _063695_, _063696_);
  xor g_121301_(out[12], out[620], _063697_);
  or g_121302_(_063682_, _063697_, _063698_);
  xor g_121303_(out[7], out[615], _063699_);
  or g_121304_(_063683_, _063699_, _063701_);
  or g_121305_(_063698_, _063701_, _063702_);
  or g_121306_(_063672_, _063673_, _063703_);
  or g_121307_(_063686_, _063703_, _063704_);
  or g_121308_(_063702_, _063704_, _063705_);
  or g_121309_(_063675_, _063705_, _063706_);
  or g_121310_(_063696_, _063706_, _063707_);
  xor g_121311_(out[465], out[593], _063708_);
  and g_121312_(out[475], _049576_, _063709_);
  xor g_121313_(out[473], out[601], _063710_);
  xor g_121314_(out[464], out[592], _063712_);
  xor g_121315_(out[478], out[606], _063713_);
  xor g_121316_(out[468], out[596], _063714_);
  or g_121317_(_063713_, _063714_, _063715_);
  xor g_121318_(out[477], out[605], _063716_);
  xor g_121319_(out[467], out[595], _063717_);
  and g_121320_(_049499_, out[603], _063718_);
  xor g_121321_(out[470], out[598], _063719_);
  xor g_121322_(out[474], out[602], _063720_);
  xor g_121323_(out[469], out[597], _063721_);
  xor g_121324_(out[479], out[607], _063723_);
  xor g_121325_(out[472], out[600], _063724_);
  or g_121326_(_063716_, _063724_, _063725_);
  xor g_121327_(out[466], out[594], _063726_);
  or g_121328_(_063720_, _063726_, _063727_);
  or g_121329_(_063725_, _063727_, _063728_);
  or g_121330_(_063710_, _063717_, _063729_);
  or g_121331_(_063721_, _063729_, _063730_);
  or g_121332_(_063728_, _063730_, _063731_);
  or g_121333_(_063715_, _063731_, _063732_);
  xor g_121334_(out[476], out[604], _063734_);
  or g_121335_(_063718_, _063734_, _063735_);
  xor g_121336_(out[471], out[599], _063736_);
  or g_121337_(_063719_, _063736_, _063737_);
  or g_121338_(_063735_, _063737_, _063738_);
  or g_121339_(_063708_, _063709_, _063739_);
  or g_121340_(_063723_, _063739_, _063740_);
  or g_121341_(_063738_, _063740_, _063741_);
  or g_121342_(_063712_, _063741_, _063742_);
  or g_121343_(_063732_, _063742_, _063743_);
  xor g_121344_(out[455], out[599], _063745_);
  and g_121345_(_049477_, out[603], _063746_);
  xor g_121346_(out[462], out[606], _063747_);
  xor g_121347_(out[456], out[600], _063748_);
  xor g_121348_(out[449], out[593], _063749_);
  xor g_121349_(out[461], out[605], _063750_);
  xor g_121350_(out[457], out[601], _063751_);
  xor g_121351_(out[452], out[596], _063752_);
  xor g_121352_(out[450], out[594], _063753_);
  and g_121353_(out[459], _049576_, _063754_);
  xor g_121354_(out[451], out[595], _063756_);
  xor g_121355_(out[454], out[598], _063757_);
  xor g_121356_(out[463], out[607], _063758_);
  xor g_121357_(out[458], out[602], _063759_);
  xor g_121358_(out[453], out[597], _063760_);
  xor g_121359_(out[448], out[592], _063761_);
  or g_121360_(_063747_, _063752_, _063762_);
  or g_121361_(_063748_, _063750_, _063763_);
  or g_121362_(_063753_, _063759_, _063764_);
  or g_121363_(_063763_, _063764_, _063765_);
  or g_121364_(_063751_, _063756_, _063767_);
  or g_121365_(_063760_, _063761_, _063768_);
  or g_121366_(_063767_, _063768_, _063769_);
  or g_121367_(_063765_, _063769_, _063770_);
  xor g_121368_(out[460], out[604], _063771_);
  or g_121369_(_063746_, _063771_, _063772_);
  or g_121370_(_063745_, _063757_, _063773_);
  or g_121371_(_063772_, _063773_, _063774_);
  or g_121372_(_063749_, _063754_, _063775_);
  or g_121373_(_063758_, _063775_, _063776_);
  or g_121374_(_063774_, _063776_, _063778_);
  or g_121375_(_063770_, _063778_, _063779_);
  or g_121376_(_063762_, _063779_, _063780_);
  not g_121377_(_063780_, _063781_);
  xor g_121378_(out[433], out[593], _063782_);
  and g_121379_(out[443], _049576_, _063783_);
  xor g_121380_(out[441], out[601], _063784_);
  xor g_121381_(out[432], out[592], _063785_);
  xor g_121382_(out[446], out[606], _063786_);
  xor g_121383_(out[436], out[596], _063787_);
  or g_121384_(_063786_, _063787_, _063789_);
  xor g_121385_(out[445], out[605], _063790_);
  xor g_121386_(out[435], out[595], _063791_);
  and g_121387_(_049466_, out[603], _063792_);
  xor g_121388_(out[438], out[598], _063793_);
  xor g_121389_(out[442], out[602], _063794_);
  xor g_121390_(out[437], out[597], _063795_);
  xor g_121391_(out[447], out[607], _063796_);
  xor g_121392_(out[440], out[600], _063797_);
  or g_121393_(_063790_, _063797_, _063798_);
  xor g_121394_(out[434], out[594], _063800_);
  or g_121395_(_063794_, _063800_, _063801_);
  or g_121396_(_063798_, _063801_, _063802_);
  or g_121397_(_063784_, _063791_, _063803_);
  or g_121398_(_063795_, _063803_, _063804_);
  or g_121399_(_063802_, _063804_, _063805_);
  or g_121400_(_063789_, _063805_, _063806_);
  xor g_121401_(out[444], out[604], _063807_);
  or g_121402_(_063792_, _063807_, _063808_);
  xor g_121403_(out[439], out[599], _063809_);
  or g_121404_(_063793_, _063809_, _063811_);
  or g_121405_(_063808_, _063811_, _063812_);
  or g_121406_(_063782_, _063783_, _063813_);
  or g_121407_(_063796_, _063813_, _063814_);
  or g_121408_(_063812_, _063814_, _063815_);
  or g_121409_(_063785_, _063815_, _063816_);
  or g_121410_(_063806_, _063816_, _063817_);
  xor g_121411_(out[423], out[599], _063818_);
  and g_121412_(_049455_, out[603], _063819_);
  xor g_121413_(out[430], out[606], _063820_);
  xor g_121414_(out[424], out[600], _063822_);
  xor g_121415_(out[417], out[593], _063823_);
  xor g_121416_(out[429], out[605], _063824_);
  xor g_121417_(out[425], out[601], _063825_);
  xor g_121418_(out[420], out[596], _063826_);
  xor g_121419_(out[418], out[594], _063827_);
  and g_121420_(out[427], _049576_, _063828_);
  xor g_121421_(out[419], out[595], _063829_);
  xor g_121422_(out[422], out[598], _063830_);
  xor g_121423_(out[431], out[607], _063831_);
  xor g_121424_(out[426], out[602], _063833_);
  xor g_121425_(out[421], out[597], _063834_);
  xor g_121426_(out[416], out[592], _063835_);
  or g_121427_(_063820_, _063826_, _063836_);
  or g_121428_(_063822_, _063824_, _063837_);
  or g_121429_(_063827_, _063833_, _063838_);
  or g_121430_(_063837_, _063838_, _063839_);
  or g_121431_(_063825_, _063829_, _063840_);
  or g_121432_(_063834_, _063835_, _063841_);
  or g_121433_(_063840_, _063841_, _063842_);
  or g_121434_(_063839_, _063842_, _063844_);
  xor g_121435_(out[428], out[604], _063845_);
  or g_121436_(_063819_, _063845_, _063846_);
  or g_121437_(_063818_, _063830_, _063847_);
  or g_121438_(_063846_, _063847_, _063848_);
  or g_121439_(_063823_, _063828_, _063849_);
  or g_121440_(_063831_, _063849_, _063850_);
  or g_121441_(_063848_, _063850_, _063851_);
  or g_121442_(_063844_, _063851_, _063852_);
  or g_121443_(_063836_, _063852_, _063853_);
  xor g_121444_(out[401], out[593], _063855_);
  and g_121445_(out[411], _049576_, _063856_);
  xor g_121446_(out[409], out[601], _063857_);
  xor g_121447_(out[400], out[592], _063858_);
  xor g_121448_(out[414], out[606], _063859_);
  xor g_121449_(out[404], out[596], _063860_);
  or g_121450_(_063859_, _063860_, _063861_);
  xor g_121451_(out[413], out[605], _063862_);
  xor g_121452_(out[403], out[595], _063863_);
  and g_121453_(_049444_, out[603], _063864_);
  xor g_121454_(out[406], out[598], _063866_);
  xor g_121455_(out[410], out[602], _063867_);
  xor g_121456_(out[405], out[597], _063868_);
  xor g_121457_(out[415], out[607], _063869_);
  xor g_121458_(out[408], out[600], _063870_);
  or g_121459_(_063862_, _063870_, _063871_);
  xor g_121460_(out[402], out[594], _063872_);
  or g_121461_(_063867_, _063872_, _063873_);
  or g_121462_(_063871_, _063873_, _063874_);
  or g_121463_(_063857_, _063863_, _063875_);
  or g_121464_(_063868_, _063875_, _063877_);
  or g_121465_(_063874_, _063877_, _063878_);
  or g_121466_(_063861_, _063878_, _063879_);
  xor g_121467_(out[412], out[604], _063880_);
  or g_121468_(_063864_, _063880_, _063881_);
  xor g_121469_(out[407], out[599], _063882_);
  or g_121470_(_063866_, _063882_, _063883_);
  or g_121471_(_063881_, _063883_, _063884_);
  or g_121472_(_063855_, _063856_, _063885_);
  or g_121473_(_063869_, _063885_, _063886_);
  or g_121474_(_063884_, _063886_, _063888_);
  or g_121475_(_063858_, _063888_, _063889_);
  or g_121476_(_063879_, _063889_, _063890_);
  xor g_121477_(out[391], out[599], _063891_);
  and g_121478_(_049433_, out[603], _063892_);
  xor g_121479_(out[398], out[606], _063893_);
  xor g_121480_(out[392], out[600], _063894_);
  xor g_121481_(out[385], out[593], _063895_);
  xor g_121482_(out[397], out[605], _063896_);
  xor g_121483_(out[393], out[601], _063897_);
  xor g_121484_(out[388], out[596], _063899_);
  xor g_121485_(out[386], out[594], _063900_);
  and g_121486_(out[395], _049576_, _063901_);
  xor g_121487_(out[387], out[595], _063902_);
  xor g_121488_(out[390], out[598], _063903_);
  xor g_121489_(out[399], out[607], _063904_);
  xor g_121490_(out[394], out[602], _063905_);
  xor g_121491_(out[389], out[597], _063906_);
  xor g_121492_(out[384], out[592], _063907_);
  or g_121493_(_063893_, _063899_, _063908_);
  or g_121494_(_063894_, _063896_, _063910_);
  or g_121495_(_063900_, _063905_, _063911_);
  or g_121496_(_063910_, _063911_, _063912_);
  or g_121497_(_063897_, _063902_, _063913_);
  or g_121498_(_063906_, _063907_, _063914_);
  or g_121499_(_063913_, _063914_, _063915_);
  or g_121500_(_063912_, _063915_, _063916_);
  xor g_121501_(out[396], out[604], _063917_);
  or g_121502_(_063892_, _063917_, _063918_);
  or g_121503_(_063891_, _063903_, _063919_);
  or g_121504_(_063918_, _063919_, _063921_);
  or g_121505_(_063895_, _063901_, _063922_);
  or g_121506_(_063904_, _063922_, _063923_);
  or g_121507_(_063921_, _063923_, _063924_);
  or g_121508_(_063916_, _063924_, _063925_);
  or g_121509_(_063908_, _063925_, _063926_);
  xor g_121510_(out[369], out[593], _063927_);
  and g_121511_(out[379], _049576_, _063928_);
  xor g_121512_(out[382], out[606], _063929_);
  xor g_121513_(out[371], out[595], _063930_);
  xor g_121514_(out[372], out[596], _063932_);
  xor g_121515_(out[370], out[594], _063933_);
  xor g_121516_(out[377], out[601], _063934_);
  xor g_121517_(out[368], out[592], _063935_);
  and g_121518_(_049422_, out[603], _063936_);
  xor g_121519_(out[374], out[598], _063937_);
  xor g_121520_(out[378], out[602], _063938_);
  xor g_121521_(out[373], out[597], _063939_);
  xor g_121522_(out[383], out[607], _063940_);
  xor g_121523_(out[381], out[605], _063941_);
  xor g_121524_(out[376], out[600], _063943_);
  or g_121525_(_063929_, _063932_, _063944_);
  or g_121526_(_063941_, _063943_, _063945_);
  or g_121527_(_063933_, _063938_, _063946_);
  or g_121528_(_063945_, _063946_, _063947_);
  or g_121529_(_063930_, _063934_, _063948_);
  or g_121530_(_063935_, _063939_, _063949_);
  or g_121531_(_063948_, _063949_, _063950_);
  or g_121532_(_063947_, _063950_, _063951_);
  xor g_121533_(out[380], out[604], _063952_);
  or g_121534_(_063936_, _063952_, _063954_);
  xor g_121535_(out[375], out[599], _063955_);
  or g_121536_(_063937_, _063955_, _063956_);
  or g_121537_(_063954_, _063956_, _063957_);
  or g_121538_(_063927_, _063928_, _063958_);
  or g_121539_(_063940_, _063958_, _063959_);
  or g_121540_(_063957_, _063959_, _063960_);
  or g_121541_(_063951_, _063960_, _063961_);
  or g_121542_(_063944_, _063961_, _063962_);
  xor g_121543_(out[359], out[599], _063963_);
  and g_121544_(_049411_, out[603], _063965_);
  xor g_121545_(out[366], out[606], _063966_);
  xor g_121546_(out[360], out[600], _063967_);
  xor g_121547_(out[353], out[593], _063968_);
  xor g_121548_(out[365], out[605], _063969_);
  xor g_121549_(out[361], out[601], _063970_);
  xor g_121550_(out[356], out[596], _063971_);
  xor g_121551_(out[354], out[594], _063972_);
  and g_121552_(out[363], _049576_, _063973_);
  xor g_121553_(out[355], out[595], _063974_);
  xor g_121554_(out[358], out[598], _063976_);
  xor g_121555_(out[367], out[607], _063977_);
  xor g_121556_(out[362], out[602], _063978_);
  xor g_121557_(out[357], out[597], _063979_);
  xor g_121558_(out[352], out[592], _063980_);
  or g_121559_(_063966_, _063971_, _063981_);
  or g_121560_(_063967_, _063969_, _063982_);
  or g_121561_(_063972_, _063978_, _063983_);
  or g_121562_(_063982_, _063983_, _063984_);
  or g_121563_(_063970_, _063974_, _063985_);
  or g_121564_(_063979_, _063980_, _063987_);
  or g_121565_(_063985_, _063987_, _063988_);
  or g_121566_(_063984_, _063988_, _063989_);
  xor g_121567_(out[364], out[604], _063990_);
  or g_121568_(_063965_, _063990_, _063991_);
  or g_121569_(_063963_, _063976_, _063992_);
  or g_121570_(_063991_, _063992_, _063993_);
  or g_121571_(_063968_, _063973_, _063994_);
  or g_121572_(_063977_, _063994_, _063995_);
  or g_121573_(_063993_, _063995_, _063996_);
  or g_121574_(_063989_, _063996_, _063998_);
  or g_121575_(_063981_, _063998_, _063999_);
  xor g_121576_(out[337], out[593], _064000_);
  and g_121577_(out[347], _049576_, _064001_);
  xor g_121578_(out[350], out[606], _064002_);
  xor g_121579_(out[339], out[595], _064003_);
  xor g_121580_(out[340], out[596], _064004_);
  xor g_121581_(out[338], out[594], _064005_);
  xor g_121582_(out[345], out[601], _064006_);
  xor g_121583_(out[336], out[592], _064007_);
  and g_121584_(_049400_, out[603], _064009_);
  xor g_121585_(out[342], out[598], _064010_);
  xor g_121586_(out[346], out[602], _064011_);
  xor g_121587_(out[341], out[597], _064012_);
  xor g_121588_(out[351], out[607], _064013_);
  xor g_121589_(out[349], out[605], _064014_);
  xor g_121590_(out[344], out[600], _064015_);
  or g_121591_(_064002_, _064004_, _064016_);
  or g_121592_(_064014_, _064015_, _064017_);
  or g_121593_(_064005_, _064011_, _064018_);
  or g_121594_(_064017_, _064018_, _064020_);
  or g_121595_(_064003_, _064006_, _064021_);
  or g_121596_(_064007_, _064012_, _064022_);
  or g_121597_(_064021_, _064022_, _064023_);
  or g_121598_(_064020_, _064023_, _064024_);
  xor g_121599_(out[348], out[604], _064025_);
  or g_121600_(_064009_, _064025_, _064026_);
  xor g_121601_(out[343], out[599], _064027_);
  or g_121602_(_064010_, _064027_, _064028_);
  or g_121603_(_064026_, _064028_, _064029_);
  or g_121604_(_064000_, _064001_, _064031_);
  or g_121605_(_064013_, _064031_, _064032_);
  or g_121606_(_064029_, _064032_, _064033_);
  or g_121607_(_064024_, _064033_, _064034_);
  or g_121608_(_064016_, _064034_, _064035_);
  xor g_121609_(out[327], out[599], _064036_);
  and g_121610_(_098294_, out[603], _064037_);
  xor g_121611_(out[334], out[606], _064038_);
  xor g_121612_(out[328], out[600], _064039_);
  xor g_121613_(out[321], out[593], _064040_);
  xor g_121614_(out[333], out[605], _064042_);
  xor g_121615_(out[329], out[601], _064043_);
  xor g_121616_(out[324], out[596], _064044_);
  xor g_121617_(out[322], out[594], _064045_);
  and g_121618_(out[331], _049576_, _064046_);
  xor g_121619_(out[323], out[595], _064047_);
  xor g_121620_(out[326], out[598], _064048_);
  xor g_121621_(out[335], out[607], _064049_);
  xor g_121622_(out[330], out[602], _064050_);
  xor g_121623_(out[325], out[597], _064051_);
  xor g_121624_(out[320], out[592], _064053_);
  or g_121625_(_064038_, _064044_, _064054_);
  or g_121626_(_064039_, _064042_, _064055_);
  or g_121627_(_064045_, _064050_, _064056_);
  or g_121628_(_064055_, _064056_, _064057_);
  or g_121629_(_064043_, _064047_, _064058_);
  or g_121630_(_064051_, _064053_, _064059_);
  or g_121631_(_064058_, _064059_, _064060_);
  or g_121632_(_064057_, _064060_, _064061_);
  xor g_121633_(out[332], out[604], _064062_);
  or g_121634_(_064037_, _064062_, _064064_);
  or g_121635_(_064036_, _064048_, _064065_);
  or g_121636_(_064064_, _064065_, _064066_);
  or g_121637_(_064040_, _064046_, _064067_);
  or g_121638_(_064049_, _064067_, _064068_);
  or g_121639_(_064066_, _064068_, _064069_);
  or g_121640_(_064061_, _064069_, _064070_);
  or g_121641_(_064054_, _064070_, _064071_);
  xor g_121642_(out[305], out[593], _064072_);
  and g_121643_(out[315], _049576_, _064073_);
  xor g_121644_(out[313], out[601], _064075_);
  xor g_121645_(out[304], out[592], _064076_);
  xor g_121646_(out[318], out[606], _064077_);
  xor g_121647_(out[308], out[596], _064078_);
  or g_121648_(_064077_, _064078_, _064079_);
  xor g_121649_(out[317], out[605], _064080_);
  xor g_121650_(out[307], out[595], _064081_);
  and g_121651_(_098283_, out[603], _064082_);
  xor g_121652_(out[310], out[598], _064083_);
  xor g_121653_(out[314], out[602], _064084_);
  xor g_121654_(out[309], out[597], _064086_);
  xor g_121655_(out[319], out[607], _064087_);
  xor g_121656_(out[312], out[600], _064088_);
  or g_121657_(_064080_, _064088_, _064089_);
  xor g_121658_(out[306], out[594], _064090_);
  or g_121659_(_064084_, _064090_, _064091_);
  or g_121660_(_064089_, _064091_, _064092_);
  or g_121661_(_064075_, _064081_, _064093_);
  or g_121662_(_064086_, _064093_, _064094_);
  or g_121663_(_064092_, _064094_, _064095_);
  or g_121664_(_064079_, _064095_, _064097_);
  xor g_121665_(out[316], out[604], _064098_);
  or g_121666_(_064082_, _064098_, _064099_);
  xor g_121667_(out[311], out[599], _064100_);
  or g_121668_(_064083_, _064100_, _064101_);
  or g_121669_(_064099_, _064101_, _064102_);
  or g_121670_(_064072_, _064073_, _064103_);
  or g_121671_(_064087_, _064103_, _064104_);
  or g_121672_(_064102_, _064104_, _064105_);
  or g_121673_(_064076_, _064105_, _064106_);
  or g_121674_(_064097_, _064106_, _064108_);
  xor g_121675_(out[295], out[599], _064109_);
  and g_121676_(_098272_, out[603], _064110_);
  xor g_121677_(out[302], out[606], _064111_);
  xor g_121678_(out[296], out[600], _064112_);
  xor g_121679_(out[289], out[593], _064113_);
  xor g_121680_(out[301], out[605], _064114_);
  xor g_121681_(out[297], out[601], _064115_);
  xor g_121682_(out[292], out[596], _064116_);
  xor g_121683_(out[290], out[594], _064117_);
  and g_121684_(out[299], _049576_, _064119_);
  xor g_121685_(out[291], out[595], _064120_);
  xor g_121686_(out[294], out[598], _064121_);
  xor g_121687_(out[303], out[607], _064122_);
  xor g_121688_(out[298], out[602], _064123_);
  xor g_121689_(out[293], out[597], _064124_);
  xor g_121690_(out[288], out[592], _064125_);
  or g_121691_(_064111_, _064116_, _064126_);
  or g_121692_(_064112_, _064114_, _064127_);
  or g_121693_(_064117_, _064123_, _064128_);
  or g_121694_(_064127_, _064128_, _064130_);
  or g_121695_(_064115_, _064120_, _064131_);
  or g_121696_(_064124_, _064125_, _064132_);
  or g_121697_(_064131_, _064132_, _064133_);
  or g_121698_(_064130_, _064133_, _064134_);
  xor g_121699_(out[300], out[604], _064135_);
  or g_121700_(_064110_, _064135_, _064136_);
  or g_121701_(_064109_, _064121_, _064137_);
  or g_121702_(_064136_, _064137_, _064138_);
  or g_121703_(_064113_, _064119_, _064139_);
  or g_121704_(_064122_, _064139_, _064141_);
  or g_121705_(_064138_, _064141_, _064142_);
  or g_121706_(_064134_, _064142_, _064143_);
  or g_121707_(_064126_, _064143_, _064144_);
  not g_121708_(_064144_, _064145_);
  xor g_121709_(out[280], out[600], _064146_);
  xor g_121710_(out[277], out[597], _064147_);
  xor g_121711_(out[275], out[595], _064148_);
  xor g_121712_(out[286], out[606], _064149_);
  xor g_121713_(out[285], out[605], _064150_);
  xor g_121714_(out[274], out[594], _064152_);
  xor g_121715_(out[281], out[601], _064153_);
  xor g_121716_(out[278], out[598], _064154_);
  xor g_121717_(out[287], out[607], _064155_);
  xor g_121718_(out[282], out[602], _064156_);
  xor g_121719_(out[276], out[596], _064157_);
  xor g_121720_(out[272], out[592], _064158_);
  and g_121721_(_098261_, out[603], _064159_);
  and g_121722_(out[283], _049576_, _064160_);
  or g_121723_(_064146_, _064150_, _064161_);
  xor g_121724_(out[273], out[593], _064163_);
  or g_121725_(_064152_, _064156_, _064164_);
  or g_121726_(_064161_, _064164_, _064165_);
  or g_121727_(_064148_, _064153_, _064166_);
  or g_121728_(_064147_, _064166_, _064167_);
  or g_121729_(_064165_, _064167_, _064168_);
  or g_121730_(_064149_, _064157_, _064169_);
  or g_121731_(_064168_, _064169_, _064170_);
  xor g_121732_(out[284], out[604], _064171_);
  or g_121733_(_064159_, _064171_, _064172_);
  xor g_121734_(out[279], out[599], _064174_);
  or g_121735_(_064154_, _064174_, _064175_);
  or g_121736_(_064172_, _064175_, _064176_);
  or g_121737_(_064160_, _064163_, _064177_);
  or g_121738_(_064155_, _064177_, _064178_);
  or g_121739_(_064176_, _064178_, _064179_);
  or g_121740_(_064158_, _064179_, _064180_);
  or g_121741_(_064170_, _064180_, _064181_);
  xor g_121742_(out[263], out[599], _064182_);
  and g_121743_(_098250_, out[603], _064183_);
  xor g_121744_(out[270], out[606], _064185_);
  xor g_121745_(out[264], out[600], _064186_);
  xor g_121746_(out[257], out[593], _064187_);
  xor g_121747_(out[269], out[605], _064188_);
  xor g_121748_(out[265], out[601], _064189_);
  xor g_121749_(out[260], out[596], _064190_);
  xor g_121750_(out[258], out[594], _064191_);
  and g_121751_(out[267], _049576_, _064192_);
  xor g_121752_(out[259], out[595], _064193_);
  xor g_121753_(out[262], out[598], _064194_);
  xor g_121754_(out[271], out[607], _064196_);
  xor g_121755_(out[266], out[602], _064197_);
  xor g_121756_(out[261], out[597], _064198_);
  xor g_121757_(out[256], out[592], _064199_);
  or g_121758_(_064185_, _064190_, _064200_);
  or g_121759_(_064186_, _064188_, _064201_);
  or g_121760_(_064191_, _064197_, _064202_);
  or g_121761_(_064201_, _064202_, _064203_);
  or g_121762_(_064189_, _064193_, _064204_);
  or g_121763_(_064198_, _064199_, _064205_);
  or g_121764_(_064204_, _064205_, _064207_);
  or g_121765_(_064203_, _064207_, _064208_);
  xor g_121766_(out[268], out[604], _064209_);
  or g_121767_(_064183_, _064209_, _064210_);
  or g_121768_(_064182_, _064194_, _064211_);
  or g_121769_(_064210_, _064211_, _064212_);
  or g_121770_(_064187_, _064192_, _064213_);
  or g_121771_(_064196_, _064213_, _064214_);
  or g_121772_(_064212_, _064214_, _064215_);
  or g_121773_(_064208_, _064215_, _064216_);
  or g_121774_(_064200_, _064216_, _064218_);
  xor g_121775_(out[252], out[604], _064219_);
  and g_121776_(_098239_, out[603], _064220_);
  xor g_121777_(out[253], out[605], _064221_);
  xor g_121778_(out[246], out[598], _064222_);
  xor g_121779_(out[248], out[600], _064223_);
  xor g_121780_(out[249], out[601], _064224_);
  xor g_121781_(out[254], out[606], _064225_);
  xor g_121782_(out[244], out[596], _064226_);
  or g_121783_(_064225_, _064226_, _064227_);
  xor g_121784_(out[245], out[597], _064229_);
  xor g_121785_(out[241], out[593], _064230_);
  and g_121786_(out[251], _049576_, _064231_);
  xor g_121787_(out[255], out[607], _064232_);
  xor g_121788_(out[250], out[602], _064233_);
  xor g_121789_(out[240], out[592], _064234_);
  xor g_121790_(out[242], out[594], _064235_);
  xor g_121791_(out[243], out[595], _064236_);
  or g_121792_(_064221_, _064223_, _064237_);
  or g_121793_(_064233_, _064235_, _064238_);
  or g_121794_(_064237_, _064238_, _064240_);
  or g_121795_(_064224_, _064236_, _064241_);
  or g_121796_(_064229_, _064234_, _064242_);
  or g_121797_(_064241_, _064242_, _064243_);
  or g_121798_(_064240_, _064243_, _064244_);
  or g_121799_(_064219_, _064220_, _064245_);
  xor g_121800_(out[247], out[599], _064246_);
  or g_121801_(_064222_, _064246_, _064247_);
  or g_121802_(_064245_, _064247_, _064248_);
  or g_121803_(_064230_, _064231_, _064249_);
  or g_121804_(_064232_, _064249_, _064251_);
  or g_121805_(_064248_, _064251_, _064252_);
  or g_121806_(_064244_, _064252_, _064253_);
  or g_121807_(_064227_, _064253_, _064254_);
  xor g_121808_(out[231], out[599], _064255_);
  and g_121809_(_098228_, out[603], _064256_);
  xor g_121810_(out[238], out[606], _064257_);
  xor g_121811_(out[232], out[600], _064258_);
  xor g_121812_(out[225], out[593], _064259_);
  xor g_121813_(out[237], out[605], _064260_);
  xor g_121814_(out[233], out[601], _064262_);
  xor g_121815_(out[228], out[596], _064263_);
  xor g_121816_(out[226], out[594], _064264_);
  and g_121817_(out[235], _049576_, _064265_);
  xor g_121818_(out[227], out[595], _064266_);
  xor g_121819_(out[230], out[598], _064267_);
  xor g_121820_(out[239], out[607], _064268_);
  xor g_121821_(out[234], out[602], _064269_);
  xor g_121822_(out[229], out[597], _064270_);
  xor g_121823_(out[224], out[592], _064271_);
  or g_121824_(_064257_, _064263_, _064273_);
  or g_121825_(_064258_, _064260_, _064274_);
  or g_121826_(_064264_, _064269_, _064275_);
  or g_121827_(_064274_, _064275_, _064276_);
  or g_121828_(_064262_, _064266_, _064277_);
  or g_121829_(_064270_, _064271_, _064278_);
  or g_121830_(_064277_, _064278_, _064279_);
  or g_121831_(_064276_, _064279_, _064280_);
  xor g_121832_(out[236], out[604], _064281_);
  or g_121833_(_064256_, _064281_, _064282_);
  or g_121834_(_064255_, _064267_, _064284_);
  or g_121835_(_064282_, _064284_, _064285_);
  or g_121836_(_064259_, _064265_, _064286_);
  or g_121837_(_064268_, _064286_, _064287_);
  or g_121838_(_064285_, _064287_, _064288_);
  or g_121839_(_064280_, _064288_, _064289_);
  or g_121840_(_064273_, _064289_, _064290_);
  xor g_121841_(out[209], out[593], _064291_);
  and g_121842_(out[219], _049576_, _064292_);
  xor g_121843_(out[217], out[601], _064293_);
  xor g_121844_(out[208], out[592], _064295_);
  xor g_121845_(out[222], out[606], _064296_);
  xor g_121846_(out[212], out[596], _064297_);
  or g_121847_(_064296_, _064297_, _064298_);
  xor g_121848_(out[221], out[605], _064299_);
  xor g_121849_(out[211], out[595], _064300_);
  and g_121850_(_098217_, out[603], _064301_);
  xor g_121851_(out[214], out[598], _064302_);
  xor g_121852_(out[218], out[602], _064303_);
  xor g_121853_(out[213], out[597], _064304_);
  xor g_121854_(out[223], out[607], _064306_);
  xor g_121855_(out[216], out[600], _064307_);
  or g_121856_(_064299_, _064307_, _064308_);
  xor g_121857_(out[210], out[594], _064309_);
  or g_121858_(_064303_, _064309_, _064310_);
  or g_121859_(_064308_, _064310_, _064311_);
  or g_121860_(_064293_, _064300_, _064312_);
  or g_121861_(_064304_, _064312_, _064313_);
  or g_121862_(_064311_, _064313_, _064314_);
  or g_121863_(_064298_, _064314_, _064315_);
  xor g_121864_(out[220], out[604], _064317_);
  or g_121865_(_064301_, _064317_, _064318_);
  xor g_121866_(out[215], out[599], _064319_);
  or g_121867_(_064302_, _064319_, _064320_);
  or g_121868_(_064318_, _064320_, _064321_);
  or g_121869_(_064291_, _064292_, _064322_);
  or g_121870_(_064306_, _064322_, _064323_);
  or g_121871_(_064321_, _064323_, _064324_);
  or g_121872_(_064295_, _064324_, _064325_);
  or g_121873_(_064315_, _064325_, _064326_);
  xor g_121874_(out[199], out[599], _064328_);
  and g_121875_(_098206_, out[603], _064329_);
  xor g_121876_(out[206], out[606], _064330_);
  xor g_121877_(out[200], out[600], _064331_);
  xor g_121878_(out[193], out[593], _064332_);
  xor g_121879_(out[205], out[605], _064333_);
  xor g_121880_(out[201], out[601], _064334_);
  xor g_121881_(out[196], out[596], _064335_);
  xor g_121882_(out[194], out[594], _064336_);
  and g_121883_(out[203], _049576_, _064337_);
  xor g_121884_(out[195], out[595], _064339_);
  xor g_121885_(out[198], out[598], _064340_);
  xor g_121886_(out[207], out[607], _064341_);
  xor g_121887_(out[202], out[602], _064342_);
  xor g_121888_(out[197], out[597], _064343_);
  xor g_121889_(out[192], out[592], _064344_);
  or g_121890_(_064330_, _064335_, _064345_);
  or g_121891_(_064331_, _064333_, _064346_);
  or g_121892_(_064336_, _064342_, _064347_);
  or g_121893_(_064346_, _064347_, _064348_);
  or g_121894_(_064334_, _064339_, _064350_);
  or g_121895_(_064343_, _064344_, _064351_);
  or g_121896_(_064350_, _064351_, _064352_);
  or g_121897_(_064348_, _064352_, _064353_);
  xor g_121898_(out[204], out[604], _064354_);
  or g_121899_(_064329_, _064354_, _064355_);
  or g_121900_(_064328_, _064340_, _064356_);
  or g_121901_(_064355_, _064356_, _064357_);
  or g_121902_(_064332_, _064337_, _064358_);
  or g_121903_(_064341_, _064358_, _064359_);
  or g_121904_(_064357_, _064359_, _064361_);
  or g_121905_(_064353_, _064361_, _064362_);
  or g_121906_(_064345_, _064362_, _064363_);
  not g_121907_(_064363_, _064364_);
  xor g_121908_(out[177], out[593], _064365_);
  and g_121909_(out[187], _049576_, _064366_);
  xor g_121910_(out[185], out[601], _064367_);
  xor g_121911_(out[176], out[592], _064368_);
  xor g_121912_(out[190], out[606], _064369_);
  xor g_121913_(out[180], out[596], _064370_);
  or g_121914_(_064369_, _064370_, _064372_);
  xor g_121915_(out[189], out[605], _064373_);
  xor g_121916_(out[179], out[595], _064374_);
  and g_121917_(_098195_, out[603], _064375_);
  xor g_121918_(out[182], out[598], _064376_);
  xor g_121919_(out[186], out[602], _064377_);
  xor g_121920_(out[181], out[597], _064378_);
  xor g_121921_(out[191], out[607], _064379_);
  xor g_121922_(out[184], out[600], _064380_);
  or g_121923_(_064373_, _064380_, _064381_);
  xor g_121924_(out[178], out[594], _064383_);
  or g_121925_(_064377_, _064383_, _064384_);
  or g_121926_(_064381_, _064384_, _064385_);
  or g_121927_(_064367_, _064374_, _064386_);
  or g_121928_(_064378_, _064386_, _064387_);
  or g_121929_(_064385_, _064387_, _064388_);
  or g_121930_(_064372_, _064388_, _064389_);
  xor g_121931_(out[188], out[604], _064390_);
  or g_121932_(_064375_, _064390_, _064391_);
  xor g_121933_(out[183], out[599], _064392_);
  or g_121934_(_064376_, _064392_, _064394_);
  or g_121935_(_064391_, _064394_, _064395_);
  or g_121936_(_064365_, _064366_, _064396_);
  or g_121937_(_064379_, _064396_, _064397_);
  or g_121938_(_064395_, _064397_, _064398_);
  or g_121939_(_064368_, _064398_, _064399_);
  or g_121940_(_064389_, _064399_, _064400_);
  xor g_121941_(out[167], out[599], _064401_);
  and g_121942_(_098184_, out[603], _064402_);
  xor g_121943_(out[174], out[606], _064403_);
  xor g_121944_(out[168], out[600], _064405_);
  xor g_121945_(out[161], out[593], _064406_);
  xor g_121946_(out[173], out[605], _064407_);
  xor g_121947_(out[169], out[601], _064408_);
  xor g_121948_(out[164], out[596], _064409_);
  xor g_121949_(out[162], out[594], _064410_);
  and g_121950_(out[171], _049576_, _064411_);
  xor g_121951_(out[163], out[595], _064412_);
  xor g_121952_(out[166], out[598], _064413_);
  xor g_121953_(out[175], out[607], _064414_);
  xor g_121954_(out[170], out[602], _064416_);
  xor g_121955_(out[165], out[597], _064417_);
  xor g_121956_(out[160], out[592], _064418_);
  or g_121957_(_064403_, _064409_, _064419_);
  or g_121958_(_064405_, _064407_, _064420_);
  or g_121959_(_064410_, _064416_, _064421_);
  or g_121960_(_064420_, _064421_, _064422_);
  or g_121961_(_064408_, _064412_, _064423_);
  or g_121962_(_064417_, _064418_, _064424_);
  or g_121963_(_064423_, _064424_, _064425_);
  or g_121964_(_064422_, _064425_, _064427_);
  xor g_121965_(out[172], out[604], _064428_);
  or g_121966_(_064402_, _064428_, _064429_);
  or g_121967_(_064401_, _064413_, _064430_);
  or g_121968_(_064429_, _064430_, _064431_);
  or g_121969_(_064406_, _064411_, _064432_);
  or g_121970_(_064414_, _064432_, _064433_);
  or g_121971_(_064431_, _064433_, _064434_);
  or g_121972_(_064427_, _064434_, _064435_);
  or g_121973_(_064419_, _064435_, _064436_);
  xor g_121974_(out[145], out[593], _064438_);
  and g_121975_(out[155], _049576_, _064439_);
  xor g_121976_(out[153], out[601], _064440_);
  xor g_121977_(out[144], out[592], _064441_);
  xor g_121978_(out[158], out[606], _064442_);
  xor g_121979_(out[148], out[596], _064443_);
  or g_121980_(_064442_, _064443_, _064444_);
  xor g_121981_(out[157], out[605], _064445_);
  xor g_121982_(out[147], out[595], _064446_);
  and g_121983_(_098173_, out[603], _064447_);
  xor g_121984_(out[150], out[598], _064449_);
  xor g_121985_(out[154], out[602], _064450_);
  xor g_121986_(out[149], out[597], _064451_);
  xor g_121987_(out[159], out[607], _064452_);
  xor g_121988_(out[152], out[600], _064453_);
  or g_121989_(_064445_, _064453_, _064454_);
  xor g_121990_(out[146], out[594], _064455_);
  or g_121991_(_064450_, _064455_, _064456_);
  or g_121992_(_064454_, _064456_, _064457_);
  or g_121993_(_064440_, _064446_, _064458_);
  or g_121994_(_064451_, _064458_, _064460_);
  or g_121995_(_064457_, _064460_, _064461_);
  or g_121996_(_064444_, _064461_, _064462_);
  xor g_121997_(out[156], out[604], _064463_);
  or g_121998_(_064447_, _064463_, _064464_);
  xor g_121999_(out[151], out[599], _064465_);
  or g_122000_(_064449_, _064465_, _064466_);
  or g_122001_(_064464_, _064466_, _064467_);
  or g_122002_(_064438_, _064439_, _064468_);
  or g_122003_(_064452_, _064468_, _064469_);
  or g_122004_(_064467_, _064469_, _064471_);
  or g_122005_(_064441_, _064471_, _064472_);
  or g_122006_(_064462_, _064472_, _064473_);
  xor g_122007_(out[135], out[599], _064474_);
  and g_122008_(_098162_, out[603], _064475_);
  xor g_122009_(out[142], out[606], _064476_);
  xor g_122010_(out[136], out[600], _064477_);
  xor g_122011_(out[129], out[593], _064478_);
  xor g_122012_(out[141], out[605], _064479_);
  xor g_122013_(out[137], out[601], _064480_);
  xor g_122014_(out[132], out[596], _064482_);
  xor g_122015_(out[130], out[594], _064483_);
  and g_122016_(out[139], _049576_, _064484_);
  xor g_122017_(out[131], out[595], _064485_);
  xor g_122018_(out[134], out[598], _064486_);
  xor g_122019_(out[143], out[607], _064487_);
  xor g_122020_(out[138], out[602], _064488_);
  xor g_122021_(out[133], out[597], _064489_);
  xor g_122022_(out[128], out[592], _064490_);
  or g_122023_(_064476_, _064482_, _064491_);
  or g_122024_(_064477_, _064479_, _064493_);
  or g_122025_(_064483_, _064488_, _064494_);
  or g_122026_(_064493_, _064494_, _064495_);
  or g_122027_(_064480_, _064485_, _064496_);
  or g_122028_(_064489_, _064490_, _064497_);
  or g_122029_(_064496_, _064497_, _064498_);
  or g_122030_(_064495_, _064498_, _064499_);
  xor g_122031_(out[140], out[604], _064500_);
  or g_122032_(_064475_, _064500_, _064501_);
  or g_122033_(_064474_, _064486_, _064502_);
  or g_122034_(_064501_, _064502_, _064504_);
  or g_122035_(_064478_, _064484_, _064505_);
  or g_122036_(_064487_, _064505_, _064506_);
  or g_122037_(_064504_, _064506_, _064507_);
  or g_122038_(_064499_, _064507_, _064508_);
  or g_122039_(_064491_, _064508_, _064509_);
  xor g_122040_(out[122], out[602], _064510_);
  xor g_122041_(out[114], out[594], _064511_);
  xor g_122042_(out[113], out[593], _064512_);
  and g_122043_(_098151_, out[603], _064513_);
  and g_122044_(out[123], _049576_, _064515_);
  xor g_122045_(out[125], out[605], _064516_);
  xor g_122046_(out[115], out[595], _064517_);
  xor g_122047_(out[126], out[606], _064518_);
  xor g_122048_(out[124], out[604], _064519_);
  xor g_122049_(out[120], out[600], _064520_);
  xor g_122050_(out[127], out[607], _064521_);
  xor g_122051_(out[117], out[597], _064522_);
  xor g_122052_(out[118], out[598], _064523_);
  xor g_122053_(out[112], out[592], _064524_);
  xor g_122054_(out[116], out[596], _064526_);
  or g_122055_(_064516_, _064520_, _064527_);
  xor g_122056_(out[121], out[601], _064528_);
  or g_122057_(_064510_, _064511_, _064529_);
  or g_122058_(_064527_, _064529_, _064530_);
  or g_122059_(_064517_, _064528_, _064531_);
  or g_122060_(_064522_, _064531_, _064532_);
  or g_122061_(_064530_, _064532_, _064533_);
  or g_122062_(_064518_, _064526_, _064534_);
  or g_122063_(_064533_, _064534_, _064535_);
  or g_122064_(_064513_, _064519_, _064537_);
  xor g_122065_(out[119], out[599], _064538_);
  or g_122066_(_064523_, _064538_, _064539_);
  or g_122067_(_064537_, _064539_, _064540_);
  or g_122068_(_064512_, _064515_, _064541_);
  or g_122069_(_064521_, _064541_, _064542_);
  or g_122070_(_064540_, _064542_, _064543_);
  or g_122071_(_064524_, _064543_, _064544_);
  or g_122072_(_064535_, _064544_, _064545_);
  not g_122073_(_064545_, _064546_);
  xor g_122074_(out[103], out[599], _064548_);
  and g_122075_(_098140_, out[603], _064549_);
  xor g_122076_(out[110], out[606], _064550_);
  xor g_122077_(out[104], out[600], _064551_);
  xor g_122078_(out[97], out[593], _064552_);
  xor g_122079_(out[109], out[605], _064553_);
  xor g_122080_(out[105], out[601], _064554_);
  xor g_122081_(out[100], out[596], _064555_);
  xor g_122082_(out[98], out[594], _064556_);
  and g_122083_(out[107], _049576_, _064557_);
  xor g_122084_(out[99], out[595], _064559_);
  xor g_122085_(out[102], out[598], _064560_);
  xor g_122086_(out[111], out[607], _064561_);
  xor g_122087_(out[106], out[602], _064562_);
  xor g_122088_(out[101], out[597], _064563_);
  xor g_122089_(out[96], out[592], _064564_);
  or g_122090_(_064550_, _064555_, _064565_);
  not g_122091_(_064565_, _064566_);
  or g_122092_(_064551_, _064553_, _064567_);
  or g_122093_(_064556_, _064562_, _064568_);
  or g_122094_(_064567_, _064568_, _064570_);
  or g_122095_(_064554_, _064559_, _064571_);
  or g_122096_(_064563_, _064564_, _064572_);
  or g_122097_(_064571_, _064572_, _064573_);
  or g_122098_(_064570_, _064573_, _064574_);
  xor g_122099_(out[108], out[604], _064575_);
  or g_122100_(_064549_, _064575_, _064576_);
  or g_122101_(_064548_, _064560_, _064577_);
  or g_122102_(_064576_, _064577_, _064578_);
  or g_122103_(_064552_, _064557_, _064579_);
  or g_122104_(_064561_, _064579_, _064581_);
  or g_122105_(_064578_, _064581_, _064582_);
  or g_122106_(_064574_, _064582_, _064583_);
  not g_122107_(_064583_, _064584_);
  and g_122108_(_064566_, _064584_, _064585_);
  not g_122109_(_064585_, _064586_);
  xor g_122110_(out[81], out[593], _064587_);
  and g_122111_(out[91], _049576_, _064588_);
  xor g_122112_(out[94], out[606], _064589_);
  xor g_122113_(out[83], out[595], _064590_);
  xor g_122114_(out[84], out[596], _064592_);
  xor g_122115_(out[82], out[594], _064593_);
  xor g_122116_(out[89], out[601], _064594_);
  xor g_122117_(out[80], out[592], _064595_);
  and g_122118_(_098129_, out[603], _064596_);
  xor g_122119_(out[86], out[598], _064597_);
  xor g_122120_(out[90], out[602], _064598_);
  xor g_122121_(out[85], out[597], _064599_);
  xor g_122122_(out[95], out[607], _064600_);
  xor g_122123_(out[93], out[605], _064601_);
  xor g_122124_(out[88], out[600], _064603_);
  or g_122125_(_064589_, _064592_, _064604_);
  or g_122126_(_064601_, _064603_, _064605_);
  or g_122127_(_064593_, _064598_, _064606_);
  or g_122128_(_064605_, _064606_, _064607_);
  or g_122129_(_064590_, _064594_, _064608_);
  or g_122130_(_064595_, _064599_, _064609_);
  or g_122131_(_064608_, _064609_, _064610_);
  or g_122132_(_064607_, _064610_, _064611_);
  xor g_122133_(out[92], out[604], _064612_);
  or g_122134_(_064596_, _064612_, _064614_);
  xor g_122135_(out[87], out[599], _064615_);
  or g_122136_(_064597_, _064615_, _064616_);
  or g_122137_(_064614_, _064616_, _064617_);
  or g_122138_(_064587_, _064588_, _064618_);
  or g_122139_(_064600_, _064618_, _064619_);
  or g_122140_(_064617_, _064619_, _064620_);
  or g_122141_(_064611_, _064620_, _064621_);
  or g_122142_(_064604_, _064621_, _064622_);
  xor g_122143_(out[71], out[599], _064623_);
  and g_122144_(_098118_, out[603], _064625_);
  xor g_122145_(out[78], out[606], _064626_);
  xor g_122146_(out[72], out[600], _064627_);
  xor g_122147_(out[65], out[593], _064628_);
  xor g_122148_(out[77], out[605], _064629_);
  xor g_122149_(out[73], out[601], _064630_);
  xor g_122150_(out[68], out[596], _064631_);
  xor g_122151_(out[66], out[594], _064632_);
  and g_122152_(out[75], _049576_, _064633_);
  xor g_122153_(out[67], out[595], _064634_);
  xor g_122154_(out[70], out[598], _064636_);
  xor g_122155_(out[79], out[607], _064637_);
  xor g_122156_(out[74], out[602], _064638_);
  xor g_122157_(out[69], out[597], _064639_);
  xor g_122158_(out[64], out[592], _064640_);
  or g_122159_(_064626_, _064631_, _064641_);
  or g_122160_(_064627_, _064629_, _064642_);
  or g_122161_(_064632_, _064638_, _064643_);
  or g_122162_(_064642_, _064643_, _064644_);
  or g_122163_(_064630_, _064634_, _064645_);
  or g_122164_(_064639_, _064640_, _064647_);
  or g_122165_(_064645_, _064647_, _064648_);
  or g_122166_(_064644_, _064648_, _064649_);
  xor g_122167_(out[76], out[604], _064650_);
  or g_122168_(_064625_, _064650_, _064651_);
  or g_122169_(_064623_, _064636_, _064652_);
  or g_122170_(_064651_, _064652_, _064653_);
  or g_122171_(_064628_, _064633_, _064654_);
  or g_122172_(_064637_, _064654_, _064655_);
  or g_122173_(_064653_, _064655_, _064656_);
  or g_122174_(_064649_, _064656_, _064658_);
  or g_122175_(_064641_, _064658_, _064659_);
  xor g_122176_(out[49], out[593], _064660_);
  and g_122177_(out[59], _049576_, _064661_);
  xor g_122178_(out[57], out[601], _064662_);
  xor g_122179_(out[48], out[592], _064663_);
  xor g_122180_(out[62], out[606], _064664_);
  xor g_122181_(out[52], out[596], _064665_);
  or g_122182_(_064664_, _064665_, _064666_);
  xor g_122183_(out[61], out[605], _064667_);
  xor g_122184_(out[51], out[595], _064669_);
  and g_122185_(_098107_, out[603], _064670_);
  xor g_122186_(out[54], out[598], _064671_);
  xor g_122187_(out[58], out[602], _064672_);
  xor g_122188_(out[53], out[597], _064673_);
  xor g_122189_(out[63], out[607], _064674_);
  xor g_122190_(out[56], out[600], _064675_);
  or g_122191_(_064667_, _064675_, _064676_);
  xor g_122192_(out[50], out[594], _064677_);
  or g_122193_(_064672_, _064677_, _064678_);
  or g_122194_(_064676_, _064678_, _064680_);
  or g_122195_(_064662_, _064669_, _064681_);
  or g_122196_(_064673_, _064681_, _064682_);
  or g_122197_(_064680_, _064682_, _064683_);
  or g_122198_(_064666_, _064683_, _064684_);
  xor g_122199_(out[60], out[604], _064685_);
  or g_122200_(_064670_, _064685_, _064686_);
  xor g_122201_(out[55], out[599], _064687_);
  or g_122202_(_064671_, _064687_, _064688_);
  or g_122203_(_064686_, _064688_, _064689_);
  or g_122204_(_064660_, _064661_, _064691_);
  or g_122205_(_064674_, _064691_, _064692_);
  or g_122206_(_064689_, _064692_, _064693_);
  or g_122207_(_064663_, _064693_, _064694_);
  or g_122208_(_064684_, _064694_, _064695_);
  xor g_122209_(out[39], out[599], _064696_);
  and g_122210_(_098096_, out[603], _064697_);
  xor g_122211_(out[46], out[606], _064698_);
  xor g_122212_(out[40], out[600], _064699_);
  xor g_122213_(out[33], out[593], _064700_);
  xor g_122214_(out[45], out[605], _064702_);
  xor g_122215_(out[41], out[601], _064703_);
  xor g_122216_(out[36], out[596], _064704_);
  xor g_122217_(out[34], out[594], _064705_);
  and g_122218_(out[43], _049576_, _064706_);
  xor g_122219_(out[35], out[595], _064707_);
  xor g_122220_(out[38], out[598], _064708_);
  xor g_122221_(out[47], out[607], _064709_);
  xor g_122222_(out[42], out[602], _064710_);
  xor g_122223_(out[37], out[597], _064711_);
  xor g_122224_(out[32], out[592], _064713_);
  or g_122225_(_064698_, _064704_, _064714_);
  or g_122226_(_064699_, _064702_, _064715_);
  or g_122227_(_064705_, _064710_, _064716_);
  or g_122228_(_064715_, _064716_, _064717_);
  or g_122229_(_064703_, _064707_, _064718_);
  or g_122230_(_064711_, _064713_, _064719_);
  or g_122231_(_064718_, _064719_, _064720_);
  or g_122232_(_064717_, _064720_, _064721_);
  xor g_122233_(out[44], out[604], _064722_);
  or g_122234_(_064697_, _064722_, _064724_);
  or g_122235_(_064696_, _064708_, _064725_);
  or g_122236_(_064724_, _064725_, _064726_);
  or g_122237_(_064700_, _064706_, _064727_);
  or g_122238_(_064709_, _064727_, _064728_);
  or g_122239_(_064726_, _064728_, _064729_);
  or g_122240_(_064721_, _064729_, _064730_);
  or g_122241_(_064714_, _064730_, _064731_);
  xor g_122242_(out[17], out[593], _064732_);
  and g_122243_(out[27], _049576_, _064733_);
  xor g_122244_(out[25], out[601], _064735_);
  xor g_122245_(out[16], out[592], _064736_);
  xor g_122246_(out[30], out[606], _064737_);
  xor g_122247_(out[20], out[596], _064738_);
  or g_122248_(_064737_, _064738_, _064739_);
  xor g_122249_(out[29], out[605], _064740_);
  xor g_122250_(out[19], out[595], _064741_);
  and g_122251_(_098063_, out[603], _064742_);
  xor g_122252_(out[22], out[598], _064743_);
  xor g_122253_(out[26], out[602], _064744_);
  xor g_122254_(out[21], out[597], _064746_);
  xor g_122255_(out[31], out[607], _064747_);
  xor g_122256_(out[24], out[600], _064748_);
  or g_122257_(_064740_, _064748_, _064749_);
  xor g_122258_(out[18], out[594], _064750_);
  or g_122259_(_064744_, _064750_, _064751_);
  or g_122260_(_064749_, _064751_, _064752_);
  or g_122261_(_064735_, _064741_, _064753_);
  or g_122262_(_064746_, _064753_, _064754_);
  or g_122263_(_064752_, _064754_, _064755_);
  or g_122264_(_064739_, _064755_, _064757_);
  xor g_122265_(out[28], out[604], _064758_);
  or g_122266_(_064742_, _064758_, _064759_);
  xor g_122267_(out[23], out[599], _064760_);
  or g_122268_(_064743_, _064760_, _064761_);
  or g_122269_(_064759_, _064761_, _064762_);
  or g_122270_(_064732_, _064733_, _064763_);
  or g_122271_(_064747_, _064763_, _064764_);
  or g_122272_(_064762_, _064764_, _064765_);
  or g_122273_(_064736_, _064765_, _064766_);
  or g_122274_(_064757_, _064766_, _064768_);
  xor g_122275_(out[12], out[604], _064769_);
  and g_122276_(_098041_, out[603], _064770_);
  xor g_122277_(out[8], out[600], _064771_);
  xor g_122278_(out[6], out[598], _064772_);
  xor g_122279_(out[13], out[605], _064773_);
  xor g_122280_(out[14], out[606], _064774_);
  xor g_122281_(out[2], out[594], _064775_);
  xor g_122282_(out[9], out[601], _064776_);
  xor g_122283_(out[5], out[597], _064777_);
  xor g_122284_(out[1], out[593], _064779_);
  and g_122285_(out[11], _049576_, _064780_);
  or g_122286_(_064771_, _064773_, _064781_);
  xor g_122287_(out[15], out[607], _064782_);
  xor g_122288_(out[10], out[602], _064783_);
  xor g_122289_(out[4], out[596], _064784_);
  xor g_122290_(out[3], out[595], _064785_);
  xor g_122291_(out[0], out[592], _064786_);
  or g_122292_(_064775_, _064783_, _064787_);
  or g_122293_(_064781_, _064787_, _064788_);
  or g_122294_(_064776_, _064785_, _064790_);
  or g_122295_(_064777_, _064790_, _064791_);
  or g_122296_(_064788_, _064791_, _064792_);
  or g_122297_(_064774_, _064784_, _064793_);
  or g_122298_(_064792_, _064793_, _064794_);
  or g_122299_(_064769_, _064770_, _064795_);
  xor g_122300_(out[7], out[599], _064796_);
  or g_122301_(_064772_, _064796_, _064797_);
  or g_122302_(_064795_, _064797_, _064798_);
  or g_122303_(_064779_, _064780_, _064799_);
  or g_122304_(_064782_, _064799_, _064801_);
  or g_122305_(_064798_, _064801_, _064802_);
  or g_122306_(_064786_, _064802_, _064803_);
  or g_122307_(_064794_, _064803_, _064804_);
  xor g_122308_(out[471], out[583], _064805_);
  and g_122309_(_049499_, out[587], _064806_);
  xor g_122310_(out[478], out[590], _064807_);
  xor g_122311_(out[472], out[584], _064808_);
  xor g_122312_(out[465], out[577], _064809_);
  xor g_122313_(out[477], out[589], _064810_);
  xor g_122314_(out[473], out[585], _064812_);
  xor g_122315_(out[468], out[580], _064813_);
  xor g_122316_(out[466], out[578], _064814_);
  and g_122317_(out[475], _049565_, _064815_);
  xor g_122318_(out[467], out[579], _064816_);
  xor g_122319_(out[470], out[582], _064817_);
  xor g_122320_(out[479], out[591], _064818_);
  xor g_122321_(out[474], out[586], _064819_);
  xor g_122322_(out[469], out[581], _064820_);
  xor g_122323_(out[464], out[576], _064821_);
  or g_122324_(_064807_, _064813_, _064823_);
  or g_122325_(_064808_, _064810_, _064824_);
  or g_122326_(_064814_, _064819_, _064825_);
  or g_122327_(_064824_, _064825_, _064826_);
  or g_122328_(_064812_, _064816_, _064827_);
  or g_122329_(_064820_, _064821_, _064828_);
  or g_122330_(_064827_, _064828_, _064829_);
  or g_122331_(_064826_, _064829_, _064830_);
  xor g_122332_(out[476], out[588], _064831_);
  or g_122333_(_064806_, _064831_, _064832_);
  or g_122334_(_064805_, _064817_, _064834_);
  or g_122335_(_064832_, _064834_, _064835_);
  or g_122336_(_064809_, _064815_, _064836_);
  or g_122337_(_064818_, _064836_, _064837_);
  or g_122338_(_064835_, _064837_, _064838_);
  or g_122339_(_064830_, _064838_, _064839_);
  or g_122340_(_064823_, _064839_, _064840_);
  not g_122341_(_064840_, _064841_);
  xor g_122342_(out[460], out[588], _064842_);
  and g_122343_(_049477_, out[587], _064843_);
  xor g_122344_(out[456], out[584], _064845_);
  xor g_122345_(out[454], out[582], _064846_);
  xor g_122346_(out[461], out[589], _064847_);
  xor g_122347_(out[462], out[590], _064848_);
  xor g_122348_(out[450], out[578], _064849_);
  xor g_122349_(out[457], out[585], _064850_);
  xor g_122350_(out[453], out[581], _064851_);
  xor g_122351_(out[449], out[577], _064852_);
  and g_122352_(out[459], _049565_, _064853_);
  or g_122353_(_064845_, _064847_, _064854_);
  xor g_122354_(out[463], out[591], _064856_);
  xor g_122355_(out[458], out[586], _064857_);
  xor g_122356_(out[452], out[580], _064858_);
  xor g_122357_(out[451], out[579], _064859_);
  xor g_122358_(out[448], out[576], _064860_);
  or g_122359_(_064849_, _064857_, _064861_);
  or g_122360_(_064854_, _064861_, _064862_);
  or g_122361_(_064850_, _064859_, _064863_);
  or g_122362_(_064851_, _064863_, _064864_);
  or g_122363_(_064862_, _064864_, _064865_);
  or g_122364_(_064848_, _064858_, _064867_);
  or g_122365_(_064865_, _064867_, _064868_);
  or g_122366_(_064842_, _064843_, _064869_);
  xor g_122367_(out[455], out[583], _064870_);
  or g_122368_(_064846_, _064870_, _064871_);
  or g_122369_(_064869_, _064871_, _064872_);
  or g_122370_(_064852_, _064853_, _064873_);
  or g_122371_(_064856_, _064873_, _064874_);
  or g_122372_(_064872_, _064874_, _064875_);
  or g_122373_(_064860_, _064875_, _064876_);
  or g_122374_(_064868_, _064876_, _064878_);
  not g_122375_(_064878_, _064879_);
  xor g_122376_(out[439], out[583], _064880_);
  and g_122377_(_049466_, out[587], _064881_);
  xor g_122378_(out[446], out[590], _064882_);
  xor g_122379_(out[440], out[584], _064883_);
  xor g_122380_(out[433], out[577], _064884_);
  xor g_122381_(out[445], out[589], _064885_);
  xor g_122382_(out[441], out[585], _064886_);
  xor g_122383_(out[436], out[580], _064887_);
  xor g_122384_(out[434], out[578], _064889_);
  and g_122385_(out[443], _049565_, _064890_);
  xor g_122386_(out[435], out[579], _064891_);
  xor g_122387_(out[438], out[582], _064892_);
  xor g_122388_(out[447], out[591], _064893_);
  xor g_122389_(out[442], out[586], _064894_);
  xor g_122390_(out[437], out[581], _064895_);
  xor g_122391_(out[432], out[576], _064896_);
  or g_122392_(_064882_, _064887_, _064897_);
  or g_122393_(_064883_, _064885_, _064898_);
  or g_122394_(_064889_, _064894_, _064900_);
  or g_122395_(_064898_, _064900_, _064901_);
  or g_122396_(_064886_, _064891_, _064902_);
  or g_122397_(_064895_, _064896_, _064903_);
  or g_122398_(_064902_, _064903_, _064904_);
  or g_122399_(_064901_, _064904_, _064905_);
  xor g_122400_(out[444], out[588], _064906_);
  or g_122401_(_064881_, _064906_, _064907_);
  or g_122402_(_064880_, _064892_, _064908_);
  or g_122403_(_064907_, _064908_, _064909_);
  or g_122404_(_064884_, _064890_, _064911_);
  or g_122405_(_064893_, _064911_, _064912_);
  or g_122406_(_064909_, _064912_, _064913_);
  or g_122407_(_064905_, _064913_, _064914_);
  or g_122408_(_064897_, _064914_, _064915_);
  not g_122409_(_064915_, _064916_);
  xor g_122410_(out[417], out[577], _064917_);
  and g_122411_(out[427], _049565_, _064918_);
  xor g_122412_(out[425], out[585], _064919_);
  xor g_122413_(out[416], out[576], _064920_);
  xor g_122414_(out[430], out[590], _064922_);
  xor g_122415_(out[420], out[580], _064923_);
  or g_122416_(_064922_, _064923_, _064924_);
  xor g_122417_(out[429], out[589], _064925_);
  xor g_122418_(out[419], out[579], _064926_);
  and g_122419_(_049455_, out[587], _064927_);
  xor g_122420_(out[422], out[582], _064928_);
  xor g_122421_(out[426], out[586], _064929_);
  xor g_122422_(out[421], out[581], _064930_);
  xor g_122423_(out[431], out[591], _064931_);
  xor g_122424_(out[424], out[584], _064933_);
  or g_122425_(_064925_, _064933_, _064934_);
  xor g_122426_(out[418], out[578], _064935_);
  or g_122427_(_064929_, _064935_, _064936_);
  or g_122428_(_064934_, _064936_, _064937_);
  or g_122429_(_064919_, _064926_, _064938_);
  or g_122430_(_064930_, _064938_, _064939_);
  or g_122431_(_064937_, _064939_, _064940_);
  or g_122432_(_064924_, _064940_, _064941_);
  xor g_122433_(out[428], out[588], _064942_);
  or g_122434_(_064927_, _064942_, _064944_);
  xor g_122435_(out[423], out[583], _064945_);
  or g_122436_(_064928_, _064945_, _064946_);
  or g_122437_(_064944_, _064946_, _064947_);
  or g_122438_(_064917_, _064918_, _064948_);
  or g_122439_(_064931_, _064948_, _064949_);
  or g_122440_(_064947_, _064949_, _064950_);
  or g_122441_(_064920_, _064950_, _064951_);
  or g_122442_(_064941_, _064951_, _064952_);
  xor g_122443_(out[407], out[583], _064953_);
  and g_122444_(_049444_, out[587], _064955_);
  xor g_122445_(out[414], out[590], _064956_);
  xor g_122446_(out[408], out[584], _064957_);
  xor g_122447_(out[401], out[577], _064958_);
  xor g_122448_(out[413], out[589], _064959_);
  xor g_122449_(out[409], out[585], _064960_);
  xor g_122450_(out[404], out[580], _064961_);
  xor g_122451_(out[402], out[578], _064962_);
  and g_122452_(out[411], _049565_, _064963_);
  xor g_122453_(out[403], out[579], _064964_);
  xor g_122454_(out[406], out[582], _064966_);
  xor g_122455_(out[415], out[591], _064967_);
  xor g_122456_(out[410], out[586], _064968_);
  xor g_122457_(out[405], out[581], _064969_);
  xor g_122458_(out[400], out[576], _064970_);
  or g_122459_(_064956_, _064961_, _064971_);
  or g_122460_(_064957_, _064959_, _064972_);
  or g_122461_(_064962_, _064968_, _064973_);
  or g_122462_(_064972_, _064973_, _064974_);
  or g_122463_(_064960_, _064964_, _064975_);
  or g_122464_(_064969_, _064970_, _064977_);
  or g_122465_(_064975_, _064977_, _064978_);
  or g_122466_(_064974_, _064978_, _064979_);
  xor g_122467_(out[412], out[588], _064980_);
  or g_122468_(_064955_, _064980_, _064981_);
  or g_122469_(_064953_, _064966_, _064982_);
  or g_122470_(_064981_, _064982_, _064983_);
  or g_122471_(_064958_, _064963_, _064984_);
  or g_122472_(_064967_, _064984_, _064985_);
  or g_122473_(_064983_, _064985_, _064986_);
  or g_122474_(_064979_, _064986_, _064988_);
  or g_122475_(_064971_, _064988_, _064989_);
  xor g_122476_(out[385], out[577], _064990_);
  and g_122477_(out[395], _049565_, _064991_);
  xor g_122478_(out[393], out[585], _064992_);
  xor g_122479_(out[384], out[576], _064993_);
  xor g_122480_(out[398], out[590], _064994_);
  xor g_122481_(out[388], out[580], _064995_);
  or g_122482_(_064994_, _064995_, _064996_);
  xor g_122483_(out[397], out[589], _064997_);
  xor g_122484_(out[387], out[579], _064999_);
  and g_122485_(_049433_, out[587], _065000_);
  xor g_122486_(out[390], out[582], _065001_);
  xor g_122487_(out[394], out[586], _065002_);
  xor g_122488_(out[389], out[581], _065003_);
  xor g_122489_(out[399], out[591], _065004_);
  xor g_122490_(out[392], out[584], _065005_);
  or g_122491_(_064997_, _065005_, _065006_);
  xor g_122492_(out[386], out[578], _065007_);
  or g_122493_(_065002_, _065007_, _065008_);
  or g_122494_(_065006_, _065008_, _065010_);
  or g_122495_(_064992_, _064999_, _065011_);
  or g_122496_(_065003_, _065011_, _065012_);
  or g_122497_(_065010_, _065012_, _065013_);
  or g_122498_(_064996_, _065013_, _065014_);
  xor g_122499_(out[396], out[588], _065015_);
  or g_122500_(_065000_, _065015_, _065016_);
  xor g_122501_(out[391], out[583], _065017_);
  or g_122502_(_065001_, _065017_, _065018_);
  or g_122503_(_065016_, _065018_, _065019_);
  or g_122504_(_064990_, _064991_, _065021_);
  or g_122505_(_065004_, _065021_, _065022_);
  or g_122506_(_065019_, _065022_, _065023_);
  or g_122507_(_064993_, _065023_, _065024_);
  or g_122508_(_065014_, _065024_, _065025_);
  xor g_122509_(out[375], out[583], _065026_);
  and g_122510_(_049422_, out[587], _065027_);
  xor g_122511_(out[382], out[590], _065028_);
  xor g_122512_(out[376], out[584], _065029_);
  xor g_122513_(out[369], out[577], _065030_);
  xor g_122514_(out[381], out[589], _065032_);
  xor g_122515_(out[377], out[585], _065033_);
  xor g_122516_(out[372], out[580], _065034_);
  xor g_122517_(out[370], out[578], _065035_);
  and g_122518_(out[379], _049565_, _065036_);
  xor g_122519_(out[371], out[579], _065037_);
  xor g_122520_(out[374], out[582], _065038_);
  xor g_122521_(out[383], out[591], _065039_);
  xor g_122522_(out[378], out[586], _065040_);
  xor g_122523_(out[373], out[581], _065041_);
  xor g_122524_(out[368], out[576], _065043_);
  or g_122525_(_065028_, _065034_, _065044_);
  or g_122526_(_065029_, _065032_, _065045_);
  or g_122527_(_065035_, _065040_, _065046_);
  or g_122528_(_065045_, _065046_, _065047_);
  or g_122529_(_065033_, _065037_, _065048_);
  or g_122530_(_065041_, _065043_, _065049_);
  or g_122531_(_065048_, _065049_, _065050_);
  or g_122532_(_065047_, _065050_, _065051_);
  xor g_122533_(out[380], out[588], _065052_);
  or g_122534_(_065027_, _065052_, _065054_);
  or g_122535_(_065026_, _065038_, _065055_);
  or g_122536_(_065054_, _065055_, _065056_);
  or g_122537_(_065030_, _065036_, _065057_);
  or g_122538_(_065039_, _065057_, _065058_);
  or g_122539_(_065056_, _065058_, _065059_);
  or g_122540_(_065051_, _065059_, _065060_);
  or g_122541_(_065044_, _065060_, _065061_);
  and g_122542_(out[363], _049565_, _065062_);
  xor g_122543_(out[356], out[580], _065063_);
  xor g_122544_(out[366], out[590], _065065_);
  or g_122545_(_065063_, _065065_, _065066_);
  xor g_122546_(out[365], out[589], _065067_);
  xor g_122547_(out[355], out[579], _065068_);
  xor g_122548_(out[352], out[576], _065069_);
  and g_122549_(_049411_, out[587], _065070_);
  xor g_122550_(out[362], out[586], _065071_);
  xor g_122551_(out[367], out[591], _065072_);
  xor g_122552_(out[358], out[582], _065073_);
  xor g_122553_(out[357], out[581], _065074_);
  xor g_122554_(out[360], out[584], _065076_);
  or g_122555_(_065067_, _065076_, _065077_);
  xor g_122556_(out[354], out[578], _065078_);
  xor g_122557_(out[361], out[585], _065079_);
  xor g_122558_(out[353], out[577], _065080_);
  or g_122559_(_065071_, _065078_, _065081_);
  or g_122560_(_065077_, _065081_, _065082_);
  or g_122561_(_065068_, _065079_, _065083_);
  or g_122562_(_065074_, _065083_, _065084_);
  or g_122563_(_065082_, _065084_, _065085_);
  or g_122564_(_065066_, _065085_, _065087_);
  xor g_122565_(out[364], out[588], _065088_);
  or g_122566_(_065070_, _065088_, _065089_);
  xor g_122567_(out[359], out[583], _065090_);
  or g_122568_(_065073_, _065090_, _065091_);
  or g_122569_(_065089_, _065091_, _065092_);
  or g_122570_(_065062_, _065080_, _065093_);
  or g_122571_(_065072_, _065093_, _065094_);
  or g_122572_(_065092_, _065094_, _065095_);
  or g_122573_(_065069_, _065095_, _065096_);
  or g_122574_(_065087_, _065096_, _065098_);
  xor g_122575_(out[343], out[583], _065099_);
  and g_122576_(_049400_, out[587], _065100_);
  xor g_122577_(out[350], out[590], _065101_);
  xor g_122578_(out[344], out[584], _065102_);
  xor g_122579_(out[337], out[577], _065103_);
  xor g_122580_(out[349], out[589], _065104_);
  xor g_122581_(out[345], out[585], _065105_);
  xor g_122582_(out[340], out[580], _065106_);
  xor g_122583_(out[338], out[578], _065107_);
  and g_122584_(out[347], _049565_, _065109_);
  xor g_122585_(out[339], out[579], _065110_);
  xor g_122586_(out[342], out[582], _065111_);
  xor g_122587_(out[351], out[591], _065112_);
  xor g_122588_(out[346], out[586], _065113_);
  xor g_122589_(out[341], out[581], _065114_);
  xor g_122590_(out[336], out[576], _065115_);
  or g_122591_(_065101_, _065106_, _065116_);
  or g_122592_(_065102_, _065104_, _065117_);
  or g_122593_(_065107_, _065113_, _065118_);
  or g_122594_(_065117_, _065118_, _065120_);
  or g_122595_(_065105_, _065110_, _065121_);
  or g_122596_(_065114_, _065115_, _065122_);
  or g_122597_(_065121_, _065122_, _065123_);
  or g_122598_(_065120_, _065123_, _065124_);
  xor g_122599_(out[348], out[588], _065125_);
  or g_122600_(_065100_, _065125_, _065126_);
  or g_122601_(_065099_, _065111_, _065127_);
  or g_122602_(_065126_, _065127_, _065128_);
  or g_122603_(_065103_, _065109_, _065129_);
  or g_122604_(_065112_, _065129_, _065131_);
  or g_122605_(_065128_, _065131_, _065132_);
  or g_122606_(_065124_, _065132_, _065133_);
  or g_122607_(_065116_, _065133_, _065134_);
  xor g_122608_(out[321], out[577], _065135_);
  and g_122609_(out[331], _049565_, _065136_);
  xor g_122610_(out[329], out[585], _065137_);
  xor g_122611_(out[320], out[576], _065138_);
  xor g_122612_(out[334], out[590], _065139_);
  xor g_122613_(out[324], out[580], _065140_);
  or g_122614_(_065139_, _065140_, _065142_);
  xor g_122615_(out[333], out[589], _065143_);
  xor g_122616_(out[323], out[579], _065144_);
  and g_122617_(_098294_, out[587], _065145_);
  xor g_122618_(out[326], out[582], _065146_);
  xor g_122619_(out[330], out[586], _065147_);
  xor g_122620_(out[325], out[581], _065148_);
  xor g_122621_(out[335], out[591], _065149_);
  xor g_122622_(out[328], out[584], _065150_);
  or g_122623_(_065143_, _065150_, _065151_);
  xor g_122624_(out[322], out[578], _065153_);
  or g_122625_(_065147_, _065153_, _065154_);
  or g_122626_(_065151_, _065154_, _065155_);
  or g_122627_(_065137_, _065144_, _065156_);
  or g_122628_(_065148_, _065156_, _065157_);
  or g_122629_(_065155_, _065157_, _065158_);
  or g_122630_(_065142_, _065158_, _065159_);
  xor g_122631_(out[332], out[588], _065160_);
  or g_122632_(_065145_, _065160_, _065161_);
  xor g_122633_(out[327], out[583], _065162_);
  or g_122634_(_065146_, _065162_, _065164_);
  or g_122635_(_065161_, _065164_, _065165_);
  or g_122636_(_065135_, _065136_, _065166_);
  or g_122637_(_065149_, _065166_, _065167_);
  or g_122638_(_065165_, _065167_, _065168_);
  or g_122639_(_065138_, _065168_, _065169_);
  or g_122640_(_065159_, _065169_, _065170_);
  xor g_122641_(out[311], out[583], _065171_);
  and g_122642_(_098283_, out[587], _065172_);
  xor g_122643_(out[318], out[590], _065173_);
  xor g_122644_(out[312], out[584], _065175_);
  xor g_122645_(out[305], out[577], _065176_);
  xor g_122646_(out[317], out[589], _065177_);
  xor g_122647_(out[313], out[585], _065178_);
  xor g_122648_(out[308], out[580], _065179_);
  xor g_122649_(out[306], out[578], _065180_);
  and g_122650_(out[315], _049565_, _065181_);
  xor g_122651_(out[307], out[579], _065182_);
  xor g_122652_(out[310], out[582], _065183_);
  xor g_122653_(out[319], out[591], _065184_);
  xor g_122654_(out[314], out[586], _065186_);
  xor g_122655_(out[309], out[581], _065187_);
  xor g_122656_(out[304], out[576], _065188_);
  or g_122657_(_065173_, _065179_, _065189_);
  or g_122658_(_065175_, _065177_, _065190_);
  or g_122659_(_065180_, _065186_, _065191_);
  or g_122660_(_065190_, _065191_, _065192_);
  or g_122661_(_065178_, _065182_, _065193_);
  or g_122662_(_065187_, _065188_, _065194_);
  or g_122663_(_065193_, _065194_, _065195_);
  or g_122664_(_065192_, _065195_, _065197_);
  xor g_122665_(out[316], out[588], _065198_);
  or g_122666_(_065172_, _065198_, _065199_);
  or g_122667_(_065171_, _065183_, _065200_);
  or g_122668_(_065199_, _065200_, _065201_);
  or g_122669_(_065176_, _065181_, _065202_);
  or g_122670_(_065184_, _065202_, _065203_);
  or g_122671_(_065201_, _065203_, _065204_);
  or g_122672_(_065197_, _065204_, _065205_);
  or g_122673_(_065189_, _065205_, _065206_);
  xor g_122674_(out[289], out[577], _065208_);
  and g_122675_(_098272_, out[587], _065209_);
  and g_122676_(out[299], _049565_, _065210_);
  xor g_122677_(out[297], out[585], _065211_);
  xor g_122678_(out[288], out[576], _065212_);
  xor g_122679_(out[302], out[590], _065213_);
  xor g_122680_(out[292], out[580], _065214_);
  or g_122681_(_065213_, _065214_, _065215_);
  xor g_122682_(out[301], out[589], _065216_);
  xor g_122683_(out[291], out[579], _065217_);
  xor g_122684_(out[300], out[588], _065219_);
  xor g_122685_(out[294], out[582], _065220_);
  xor g_122686_(out[298], out[586], _065221_);
  xor g_122687_(out[293], out[581], _065222_);
  xor g_122688_(out[303], out[591], _065223_);
  xor g_122689_(out[296], out[584], _065224_);
  or g_122690_(_065216_, _065224_, _065225_);
  xor g_122691_(out[290], out[578], _065226_);
  or g_122692_(_065221_, _065226_, _065227_);
  or g_122693_(_065225_, _065227_, _065228_);
  or g_122694_(_065211_, _065217_, _065230_);
  or g_122695_(_065222_, _065230_, _065231_);
  or g_122696_(_065228_, _065231_, _065232_);
  or g_122697_(_065215_, _065232_, _065233_);
  or g_122698_(_065209_, _065219_, _065234_);
  xor g_122699_(out[295], out[583], _065235_);
  or g_122700_(_065220_, _065235_, _065236_);
  or g_122701_(_065234_, _065236_, _065237_);
  or g_122702_(_065208_, _065210_, _065238_);
  or g_122703_(_065223_, _065238_, _065239_);
  or g_122704_(_065237_, _065239_, _065241_);
  or g_122705_(_065212_, _065241_, _065242_);
  or g_122706_(_065233_, _065242_, _065243_);
  not g_122707_(_065243_, _065244_);
  xor g_122708_(out[279], out[583], _065245_);
  and g_122709_(_098261_, out[587], _065246_);
  xor g_122710_(out[286], out[590], _065247_);
  xor g_122711_(out[280], out[584], _065248_);
  xor g_122712_(out[273], out[577], _065249_);
  xor g_122713_(out[285], out[589], _065250_);
  xor g_122714_(out[281], out[585], _065252_);
  xor g_122715_(out[276], out[580], _065253_);
  xor g_122716_(out[274], out[578], _065254_);
  and g_122717_(out[283], _049565_, _065255_);
  xor g_122718_(out[275], out[579], _065256_);
  xor g_122719_(out[278], out[582], _065257_);
  xor g_122720_(out[287], out[591], _065258_);
  xor g_122721_(out[282], out[586], _065259_);
  xor g_122722_(out[277], out[581], _065260_);
  xor g_122723_(out[272], out[576], _065261_);
  or g_122724_(_065247_, _065253_, _065263_);
  or g_122725_(_065248_, _065250_, _065264_);
  or g_122726_(_065254_, _065259_, _065265_);
  or g_122727_(_065264_, _065265_, _065266_);
  or g_122728_(_065252_, _065256_, _065267_);
  or g_122729_(_065260_, _065261_, _065268_);
  or g_122730_(_065267_, _065268_, _065269_);
  or g_122731_(_065266_, _065269_, _065270_);
  xor g_122732_(out[284], out[588], _065271_);
  or g_122733_(_065246_, _065271_, _065272_);
  or g_122734_(_065245_, _065257_, _065274_);
  or g_122735_(_065272_, _065274_, _065275_);
  or g_122736_(_065249_, _065255_, _065276_);
  or g_122737_(_065258_, _065276_, _065277_);
  or g_122738_(_065275_, _065277_, _065278_);
  or g_122739_(_065270_, _065278_, _065279_);
  or g_122740_(_065263_, _065279_, _065280_);
  xor g_122741_(out[266], out[586], _065281_);
  xor g_122742_(out[264], out[584], _065282_);
  xor g_122743_(out[257], out[577], _065283_);
  and g_122744_(_098250_, out[587], _065285_);
  and g_122745_(out[267], _049565_, _065286_);
  xor g_122746_(out[258], out[578], _065287_);
  xor g_122747_(out[261], out[581], _065288_);
  xor g_122748_(out[265], out[585], _065289_);
  xor g_122749_(out[268], out[588], _065290_);
  xor g_122750_(out[269], out[589], _065291_);
  xor g_122751_(out[271], out[591], _065292_);
  xor g_122752_(out[260], out[580], _065293_);
  xor g_122753_(out[262], out[582], _065294_);
  xor g_122754_(out[259], out[579], _065296_);
  xor g_122755_(out[256], out[576], _065297_);
  xor g_122756_(out[270], out[590], _065298_);
  or g_122757_(_065293_, _065298_, _065299_);
  or g_122758_(_065282_, _065291_, _065300_);
  or g_122759_(_065281_, _065287_, _065301_);
  or g_122760_(_065300_, _065301_, _065302_);
  or g_122761_(_065289_, _065296_, _065303_);
  or g_122762_(_065288_, _065297_, _065304_);
  or g_122763_(_065303_, _065304_, _065305_);
  or g_122764_(_065302_, _065305_, _065307_);
  or g_122765_(_065285_, _065290_, _065308_);
  xor g_122766_(out[263], out[583], _065309_);
  or g_122767_(_065294_, _065309_, _065310_);
  or g_122768_(_065308_, _065310_, _065311_);
  or g_122769_(_065283_, _065286_, _065312_);
  or g_122770_(_065292_, _065312_, _065313_);
  or g_122771_(_065311_, _065313_, _065314_);
  or g_122772_(_065307_, _065314_, _065315_);
  or g_122773_(_065299_, _065315_, _065316_);
  xor g_122774_(out[247], out[583], _065318_);
  and g_122775_(_098239_, out[587], _065319_);
  xor g_122776_(out[254], out[590], _065320_);
  xor g_122777_(out[248], out[584], _065321_);
  xor g_122778_(out[241], out[577], _065322_);
  xor g_122779_(out[253], out[589], _065323_);
  xor g_122780_(out[249], out[585], _065324_);
  xor g_122781_(out[244], out[580], _065325_);
  xor g_122782_(out[242], out[578], _065326_);
  and g_122783_(out[251], _049565_, _065327_);
  xor g_122784_(out[243], out[579], _065329_);
  xor g_122785_(out[246], out[582], _065330_);
  xor g_122786_(out[255], out[591], _065331_);
  xor g_122787_(out[250], out[586], _065332_);
  xor g_122788_(out[245], out[581], _065333_);
  xor g_122789_(out[240], out[576], _065334_);
  or g_122790_(_065320_, _065325_, _065335_);
  or g_122791_(_065321_, _065323_, _065336_);
  or g_122792_(_065326_, _065332_, _065337_);
  or g_122793_(_065336_, _065337_, _065338_);
  or g_122794_(_065324_, _065329_, _065340_);
  or g_122795_(_065333_, _065334_, _065341_);
  or g_122796_(_065340_, _065341_, _065342_);
  or g_122797_(_065338_, _065342_, _065343_);
  xor g_122798_(out[252], out[588], _065344_);
  or g_122799_(_065319_, _065344_, _065345_);
  or g_122800_(_065318_, _065330_, _065346_);
  or g_122801_(_065345_, _065346_, _065347_);
  or g_122802_(_065322_, _065327_, _065348_);
  or g_122803_(_065331_, _065348_, _065349_);
  or g_122804_(_065347_, _065349_, _065351_);
  or g_122805_(_065343_, _065351_, _065352_);
  or g_122806_(_065335_, _065352_, _065353_);
  not g_122807_(_065353_, _065354_);
  xor g_122808_(out[225], out[577], _065355_);
  and g_122809_(out[235], _049565_, _065356_);
  xor g_122810_(out[233], out[585], _065357_);
  xor g_122811_(out[224], out[576], _065358_);
  xor g_122812_(out[238], out[590], _065359_);
  xor g_122813_(out[228], out[580], _065360_);
  or g_122814_(_065359_, _065360_, _065362_);
  xor g_122815_(out[237], out[589], _065363_);
  xor g_122816_(out[227], out[579], _065364_);
  and g_122817_(_098228_, out[587], _065365_);
  xor g_122818_(out[230], out[582], _065366_);
  xor g_122819_(out[234], out[586], _065367_);
  xor g_122820_(out[229], out[581], _065368_);
  xor g_122821_(out[239], out[591], _065369_);
  xor g_122822_(out[232], out[584], _065370_);
  or g_122823_(_065363_, _065370_, _065371_);
  xor g_122824_(out[226], out[578], _065373_);
  or g_122825_(_065367_, _065373_, _065374_);
  or g_122826_(_065371_, _065374_, _065375_);
  or g_122827_(_065357_, _065364_, _065376_);
  or g_122828_(_065368_, _065376_, _065377_);
  or g_122829_(_065375_, _065377_, _065378_);
  or g_122830_(_065362_, _065378_, _065379_);
  xor g_122831_(out[236], out[588], _065380_);
  or g_122832_(_065365_, _065380_, _065381_);
  xor g_122833_(out[231], out[583], _065382_);
  or g_122834_(_065366_, _065382_, _065384_);
  or g_122835_(_065381_, _065384_, _065385_);
  or g_122836_(_065355_, _065356_, _065386_);
  or g_122837_(_065369_, _065386_, _065387_);
  or g_122838_(_065385_, _065387_, _065388_);
  or g_122839_(_065358_, _065388_, _065389_);
  or g_122840_(_065379_, _065389_, _065390_);
  not g_122841_(_065390_, _065391_);
  xor g_122842_(out[215], out[583], _065392_);
  and g_122843_(_098217_, out[587], _065393_);
  xor g_122844_(out[222], out[590], _065395_);
  xor g_122845_(out[216], out[584], _065396_);
  xor g_122846_(out[209], out[577], _065397_);
  xor g_122847_(out[221], out[589], _065398_);
  xor g_122848_(out[217], out[585], _065399_);
  xor g_122849_(out[212], out[580], _065400_);
  xor g_122850_(out[210], out[578], _065401_);
  and g_122851_(out[219], _049565_, _065402_);
  xor g_122852_(out[211], out[579], _065403_);
  xor g_122853_(out[214], out[582], _065404_);
  xor g_122854_(out[223], out[591], _065406_);
  xor g_122855_(out[218], out[586], _065407_);
  xor g_122856_(out[213], out[581], _065408_);
  xor g_122857_(out[208], out[576], _065409_);
  or g_122858_(_065395_, _065400_, _065410_);
  or g_122859_(_065396_, _065398_, _065411_);
  or g_122860_(_065401_, _065407_, _065412_);
  or g_122861_(_065411_, _065412_, _065413_);
  or g_122862_(_065399_, _065403_, _065414_);
  or g_122863_(_065408_, _065409_, _065415_);
  or g_122864_(_065414_, _065415_, _065417_);
  or g_122865_(_065413_, _065417_, _065418_);
  xor g_122866_(out[220], out[588], _065419_);
  or g_122867_(_065393_, _065419_, _065420_);
  or g_122868_(_065392_, _065404_, _065421_);
  or g_122869_(_065420_, _065421_, _065422_);
  or g_122870_(_065397_, _065402_, _065423_);
  or g_122871_(_065406_, _065423_, _065424_);
  or g_122872_(_065422_, _065424_, _065425_);
  or g_122873_(_065418_, _065425_, _065426_);
  or g_122874_(_065410_, _065426_, _065428_);
  xor g_122875_(out[195], out[579], _065429_);
  xor g_122876_(out[196], out[580], _065430_);
  xor g_122877_(out[206], out[590], _065431_);
  xor g_122878_(out[194], out[578], _065432_);
  xor g_122879_(out[197], out[581], _065433_);
  xor g_122880_(out[201], out[585], _065434_);
  xor g_122881_(out[200], out[584], _065435_);
  xor g_122882_(out[207], out[591], _065436_);
  xor g_122883_(out[202], out[586], _065437_);
  xor g_122884_(out[198], out[582], _065439_);
  xor g_122885_(out[192], out[576], _065440_);
  and g_122886_(_098206_, out[587], _065441_);
  and g_122887_(out[203], _049565_, _065442_);
  xor g_122888_(out[205], out[589], _065443_);
  or g_122889_(_065435_, _065443_, _065444_);
  xor g_122890_(out[193], out[577], _065445_);
  or g_122891_(_065432_, _065437_, _065446_);
  or g_122892_(_065444_, _065446_, _065447_);
  or g_122893_(_065429_, _065434_, _065448_);
  or g_122894_(_065433_, _065448_, _065450_);
  or g_122895_(_065447_, _065450_, _065451_);
  or g_122896_(_065430_, _065431_, _065452_);
  or g_122897_(_065451_, _065452_, _065453_);
  xor g_122898_(out[204], out[588], _065454_);
  or g_122899_(_065441_, _065454_, _065455_);
  xor g_122900_(out[199], out[583], _065456_);
  or g_122901_(_065439_, _065456_, _065457_);
  or g_122902_(_065455_, _065457_, _065458_);
  or g_122903_(_065442_, _065445_, _065459_);
  or g_122904_(_065436_, _065459_, _065461_);
  or g_122905_(_065458_, _065461_, _065462_);
  or g_122906_(_065440_, _065462_, _065463_);
  or g_122907_(_065453_, _065463_, _065464_);
  not g_122908_(_065464_, _065465_);
  xor g_122909_(out[183], out[583], _065466_);
  and g_122910_(_098195_, out[587], _065467_);
  xor g_122911_(out[190], out[590], _065468_);
  xor g_122912_(out[184], out[584], _065469_);
  xor g_122913_(out[177], out[577], _065470_);
  xor g_122914_(out[189], out[589], _065472_);
  xor g_122915_(out[185], out[585], _065473_);
  xor g_122916_(out[180], out[580], _065474_);
  xor g_122917_(out[178], out[578], _065475_);
  and g_122918_(out[187], _049565_, _065476_);
  xor g_122919_(out[179], out[579], _065477_);
  xor g_122920_(out[182], out[582], _065478_);
  xor g_122921_(out[191], out[591], _065479_);
  xor g_122922_(out[186], out[586], _065480_);
  xor g_122923_(out[181], out[581], _065481_);
  xor g_122924_(out[176], out[576], _065483_);
  or g_122925_(_065468_, _065474_, _065484_);
  or g_122926_(_065469_, _065472_, _065485_);
  or g_122927_(_065475_, _065480_, _065486_);
  or g_122928_(_065485_, _065486_, _065487_);
  or g_122929_(_065473_, _065477_, _065488_);
  or g_122930_(_065481_, _065483_, _065489_);
  or g_122931_(_065488_, _065489_, _065490_);
  or g_122932_(_065487_, _065490_, _065491_);
  xor g_122933_(out[188], out[588], _065492_);
  or g_122934_(_065467_, _065492_, _065494_);
  or g_122935_(_065466_, _065478_, _065495_);
  or g_122936_(_065494_, _065495_, _065496_);
  or g_122937_(_065470_, _065476_, _065497_);
  or g_122938_(_065479_, _065497_, _065498_);
  or g_122939_(_065496_, _065498_, _065499_);
  or g_122940_(_065491_, _065499_, _065500_);
  or g_122941_(_065484_, _065500_, _065501_);
  xor g_122942_(out[172], out[588], _065502_);
  and g_122943_(_098184_, out[587], _065503_);
  xor g_122944_(out[173], out[589], _065505_);
  xor g_122945_(out[166], out[582], _065506_);
  xor g_122946_(out[168], out[584], _065507_);
  xor g_122947_(out[169], out[585], _065508_);
  xor g_122948_(out[174], out[590], _065509_);
  xor g_122949_(out[164], out[580], _065510_);
  or g_122950_(_065509_, _065510_, _065511_);
  xor g_122951_(out[165], out[581], _065512_);
  xor g_122952_(out[161], out[577], _065513_);
  and g_122953_(out[171], _049565_, _065514_);
  xor g_122954_(out[175], out[591], _065516_);
  xor g_122955_(out[170], out[586], _065517_);
  xor g_122956_(out[160], out[576], _065518_);
  xor g_122957_(out[162], out[578], _065519_);
  xor g_122958_(out[163], out[579], _065520_);
  or g_122959_(_065505_, _065507_, _065521_);
  or g_122960_(_065517_, _065519_, _065522_);
  or g_122961_(_065521_, _065522_, _065523_);
  or g_122962_(_065508_, _065520_, _065524_);
  or g_122963_(_065512_, _065518_, _065525_);
  or g_122964_(_065524_, _065525_, _065527_);
  or g_122965_(_065523_, _065527_, _065528_);
  or g_122966_(_065502_, _065503_, _065529_);
  xor g_122967_(out[167], out[583], _065530_);
  or g_122968_(_065506_, _065530_, _065531_);
  or g_122969_(_065529_, _065531_, _065532_);
  or g_122970_(_065513_, _065514_, _065533_);
  or g_122971_(_065516_, _065533_, _065534_);
  or g_122972_(_065532_, _065534_, _065535_);
  or g_122973_(_065528_, _065535_, _065536_);
  or g_122974_(_065511_, _065536_, _065538_);
  xor g_122975_(out[151], out[583], _065539_);
  and g_122976_(_098173_, out[587], _065540_);
  xor g_122977_(out[158], out[590], _065541_);
  xor g_122978_(out[152], out[584], _065542_);
  xor g_122979_(out[145], out[577], _065543_);
  xor g_122980_(out[157], out[589], _065544_);
  xor g_122981_(out[153], out[585], _065545_);
  xor g_122982_(out[148], out[580], _065546_);
  xor g_122983_(out[146], out[578], _065547_);
  and g_122984_(out[155], _049565_, _065549_);
  xor g_122985_(out[147], out[579], _065550_);
  xor g_122986_(out[150], out[582], _065551_);
  xor g_122987_(out[159], out[591], _065552_);
  xor g_122988_(out[154], out[586], _065553_);
  xor g_122989_(out[149], out[581], _065554_);
  xor g_122990_(out[144], out[576], _065555_);
  or g_122991_(_065541_, _065546_, _065556_);
  or g_122992_(_065542_, _065544_, _065557_);
  or g_122993_(_065547_, _065553_, _065558_);
  or g_122994_(_065557_, _065558_, _065560_);
  or g_122995_(_065545_, _065550_, _065561_);
  or g_122996_(_065554_, _065555_, _065562_);
  or g_122997_(_065561_, _065562_, _065563_);
  or g_122998_(_065560_, _065563_, _065564_);
  xor g_122999_(out[156], out[588], _065565_);
  or g_123000_(_065540_, _065565_, _065566_);
  or g_123001_(_065539_, _065551_, _065567_);
  or g_123002_(_065566_, _065567_, _065568_);
  or g_123003_(_065543_, _065549_, _065569_);
  or g_123004_(_065552_, _065569_, _065571_);
  or g_123005_(_065568_, _065571_, _065572_);
  or g_123006_(_065564_, _065572_, _065573_);
  or g_123007_(_065556_, _065573_, _065574_);
  xor g_123008_(out[136], out[584], _065575_);
  xor g_123009_(out[133], out[581], _065576_);
  xor g_123010_(out[131], out[579], _065577_);
  xor g_123011_(out[142], out[590], _065578_);
  xor g_123012_(out[141], out[589], _065579_);
  xor g_123013_(out[130], out[578], _065580_);
  xor g_123014_(out[137], out[585], _065582_);
  xor g_123015_(out[134], out[582], _065583_);
  xor g_123016_(out[143], out[591], _065584_);
  xor g_123017_(out[138], out[586], _065585_);
  xor g_123018_(out[132], out[580], _065586_);
  xor g_123019_(out[128], out[576], _065587_);
  and g_123020_(_098162_, out[587], _065588_);
  and g_123021_(out[139], _049565_, _065589_);
  or g_123022_(_065575_, _065579_, _065590_);
  xor g_123023_(out[129], out[577], _065591_);
  or g_123024_(_065580_, _065585_, _065593_);
  or g_123025_(_065590_, _065593_, _065594_);
  or g_123026_(_065577_, _065582_, _065595_);
  or g_123027_(_065576_, _065595_, _065596_);
  or g_123028_(_065594_, _065596_, _065597_);
  or g_123029_(_065578_, _065586_, _065598_);
  or g_123030_(_065597_, _065598_, _065599_);
  xor g_123031_(out[140], out[588], _065600_);
  or g_123032_(_065588_, _065600_, _065601_);
  xor g_123033_(out[135], out[583], _065602_);
  or g_123034_(_065583_, _065602_, _065604_);
  or g_123035_(_065601_, _065604_, _065605_);
  or g_123036_(_065589_, _065591_, _065606_);
  or g_123037_(_065584_, _065606_, _065607_);
  or g_123038_(_065605_, _065607_, _065608_);
  or g_123039_(_065587_, _065608_, _065609_);
  or g_123040_(_065599_, _065609_, _065610_);
  xor g_123041_(out[119], out[583], _065611_);
  and g_123042_(_098151_, out[587], _065612_);
  xor g_123043_(out[126], out[590], _065613_);
  xor g_123044_(out[120], out[584], _065615_);
  xor g_123045_(out[113], out[577], _065616_);
  xor g_123046_(out[125], out[589], _065617_);
  xor g_123047_(out[121], out[585], _065618_);
  xor g_123048_(out[116], out[580], _065619_);
  xor g_123049_(out[114], out[578], _065620_);
  and g_123050_(out[123], _049565_, _065621_);
  xor g_123051_(out[115], out[579], _065622_);
  xor g_123052_(out[118], out[582], _065623_);
  xor g_123053_(out[127], out[591], _065624_);
  xor g_123054_(out[122], out[586], _065626_);
  xor g_123055_(out[117], out[581], _065627_);
  xor g_123056_(out[112], out[576], _065628_);
  or g_123057_(_065613_, _065619_, _065629_);
  or g_123058_(_065615_, _065617_, _065630_);
  or g_123059_(_065620_, _065626_, _065631_);
  or g_123060_(_065630_, _065631_, _065632_);
  or g_123061_(_065618_, _065622_, _065633_);
  or g_123062_(_065627_, _065628_, _065634_);
  or g_123063_(_065633_, _065634_, _065635_);
  or g_123064_(_065632_, _065635_, _065637_);
  xor g_123065_(out[124], out[588], _065638_);
  or g_123066_(_065612_, _065638_, _065639_);
  or g_123067_(_065611_, _065623_, _065640_);
  or g_123068_(_065639_, _065640_, _065641_);
  or g_123069_(_065616_, _065621_, _065642_);
  or g_123070_(_065624_, _065642_, _065643_);
  or g_123071_(_065641_, _065643_, _065644_);
  or g_123072_(_065637_, _065644_, _065645_);
  or g_123073_(_065629_, _065645_, _065646_);
  xor g_123074_(out[108], out[588], _065648_);
  and g_123075_(_098140_, out[587], _065649_);
  xor g_123076_(out[104], out[584], _065650_);
  xor g_123077_(out[102], out[582], _065651_);
  xor g_123078_(out[109], out[589], _065652_);
  xor g_123079_(out[110], out[590], _065653_);
  xor g_123080_(out[98], out[578], _065654_);
  xor g_123081_(out[105], out[585], _065655_);
  xor g_123082_(out[101], out[581], _065656_);
  xor g_123083_(out[97], out[577], _065657_);
  and g_123084_(out[107], _049565_, _065659_);
  or g_123085_(_065650_, _065652_, _065660_);
  xor g_123086_(out[111], out[591], _065661_);
  xor g_123087_(out[106], out[586], _065662_);
  xor g_123088_(out[100], out[580], _065663_);
  xor g_123089_(out[99], out[579], _065664_);
  xor g_123090_(out[96], out[576], _065665_);
  or g_123091_(_065654_, _065662_, _065666_);
  or g_123092_(_065660_, _065666_, _065667_);
  or g_123093_(_065655_, _065664_, _065668_);
  or g_123094_(_065656_, _065668_, _065670_);
  or g_123095_(_065667_, _065670_, _065671_);
  or g_123096_(_065653_, _065663_, _065672_);
  or g_123097_(_065671_, _065672_, _065673_);
  or g_123098_(_065648_, _065649_, _065674_);
  xor g_123099_(out[103], out[583], _065675_);
  or g_123100_(_065651_, _065675_, _065676_);
  or g_123101_(_065674_, _065676_, _065677_);
  or g_123102_(_065657_, _065659_, _065678_);
  or g_123103_(_065661_, _065678_, _065679_);
  or g_123104_(_065677_, _065679_, _065681_);
  or g_123105_(_065665_, _065681_, _065682_);
  or g_123106_(_065673_, _065682_, _065683_);
  xor g_123107_(out[87], out[583], _065684_);
  and g_123108_(_098129_, out[587], _065685_);
  xor g_123109_(out[94], out[590], _065686_);
  xor g_123110_(out[88], out[584], _065687_);
  xor g_123111_(out[81], out[577], _065688_);
  xor g_123112_(out[93], out[589], _065689_);
  xor g_123113_(out[89], out[585], _065690_);
  xor g_123114_(out[84], out[580], _065692_);
  xor g_123115_(out[82], out[578], _065693_);
  and g_123116_(out[91], _049565_, _065694_);
  xor g_123117_(out[83], out[579], _065695_);
  xor g_123118_(out[86], out[582], _065696_);
  xor g_123119_(out[95], out[591], _065697_);
  xor g_123120_(out[90], out[586], _065698_);
  xor g_123121_(out[85], out[581], _065699_);
  xor g_123122_(out[80], out[576], _065700_);
  or g_123123_(_065686_, _065692_, _065701_);
  or g_123124_(_065687_, _065689_, _065703_);
  or g_123125_(_065693_, _065698_, _065704_);
  or g_123126_(_065703_, _065704_, _065705_);
  or g_123127_(_065690_, _065695_, _065706_);
  or g_123128_(_065699_, _065700_, _065707_);
  or g_123129_(_065706_, _065707_, _065708_);
  or g_123130_(_065705_, _065708_, _065709_);
  xor g_123131_(out[92], out[588], _065710_);
  or g_123132_(_065685_, _065710_, _065711_);
  or g_123133_(_065684_, _065696_, _065712_);
  or g_123134_(_065711_, _065712_, _065714_);
  or g_123135_(_065688_, _065694_, _065715_);
  or g_123136_(_065697_, _065715_, _065716_);
  or g_123137_(_065714_, _065716_, _065717_);
  or g_123138_(_065709_, _065717_, _065718_);
  or g_123139_(_065701_, _065718_, _065719_);
  not g_123140_(_065719_, _065720_);
  xor g_123141_(out[65], out[577], _065721_);
  and g_123142_(out[75], _049565_, _065722_);
  xor g_123143_(out[78], out[590], _065723_);
  xor g_123144_(out[67], out[579], _065725_);
  xor g_123145_(out[68], out[580], _065726_);
  xor g_123146_(out[66], out[578], _065727_);
  xor g_123147_(out[73], out[585], _065728_);
  xor g_123148_(out[64], out[576], _065729_);
  and g_123149_(_098118_, out[587], _065730_);
  xor g_123150_(out[70], out[582], _065731_);
  xor g_123151_(out[74], out[586], _065732_);
  xor g_123152_(out[69], out[581], _065733_);
  xor g_123153_(out[79], out[591], _065734_);
  xor g_123154_(out[77], out[589], _065736_);
  xor g_123155_(out[72], out[584], _065737_);
  or g_123156_(_065723_, _065726_, _065738_);
  or g_123157_(_065736_, _065737_, _065739_);
  or g_123158_(_065727_, _065732_, _065740_);
  or g_123159_(_065739_, _065740_, _065741_);
  or g_123160_(_065725_, _065728_, _065742_);
  or g_123161_(_065729_, _065733_, _065743_);
  or g_123162_(_065742_, _065743_, _065744_);
  or g_123163_(_065741_, _065744_, _065745_);
  xor g_123164_(out[76], out[588], _065747_);
  or g_123165_(_065730_, _065747_, _065748_);
  xor g_123166_(out[71], out[583], _065749_);
  or g_123167_(_065731_, _065749_, _065750_);
  or g_123168_(_065748_, _065750_, _065751_);
  or g_123169_(_065721_, _065722_, _065752_);
  or g_123170_(_065734_, _065752_, _065753_);
  or g_123171_(_065751_, _065753_, _065754_);
  or g_123172_(_065745_, _065754_, _065755_);
  or g_123173_(_065738_, _065755_, _065756_);
  xor g_123174_(out[55], out[583], _065758_);
  and g_123175_(_098107_, out[587], _065759_);
  xor g_123176_(out[62], out[590], _065760_);
  xor g_123177_(out[56], out[584], _065761_);
  xor g_123178_(out[49], out[577], _065762_);
  xor g_123179_(out[61], out[589], _065763_);
  xor g_123180_(out[57], out[585], _065764_);
  xor g_123181_(out[52], out[580], _065765_);
  xor g_123182_(out[50], out[578], _065766_);
  and g_123183_(out[59], _049565_, _065767_);
  xor g_123184_(out[51], out[579], _065769_);
  xor g_123185_(out[54], out[582], _065770_);
  xor g_123186_(out[63], out[591], _065771_);
  xor g_123187_(out[58], out[586], _065772_);
  xor g_123188_(out[53], out[581], _065773_);
  xor g_123189_(out[48], out[576], _065774_);
  or g_123190_(_065760_, _065765_, _065775_);
  or g_123191_(_065761_, _065763_, _065776_);
  or g_123192_(_065766_, _065772_, _065777_);
  or g_123193_(_065776_, _065777_, _065778_);
  or g_123194_(_065764_, _065769_, _065780_);
  or g_123195_(_065773_, _065774_, _065781_);
  or g_123196_(_065780_, _065781_, _065782_);
  or g_123197_(_065778_, _065782_, _065783_);
  xor g_123198_(out[60], out[588], _065784_);
  or g_123199_(_065759_, _065784_, _065785_);
  or g_123200_(_065758_, _065770_, _065786_);
  or g_123201_(_065785_, _065786_, _065787_);
  or g_123202_(_065762_, _065767_, _065788_);
  or g_123203_(_065771_, _065788_, _065789_);
  or g_123204_(_065787_, _065789_, _065791_);
  or g_123205_(_065783_, _065791_, _065792_);
  or g_123206_(_065775_, _065792_, _065793_);
  xor g_123207_(out[33], out[577], _065794_);
  and g_123208_(_098096_, out[587], _065795_);
  and g_123209_(out[43], _049565_, _065796_);
  xor g_123210_(out[41], out[585], _065797_);
  xor g_123211_(out[32], out[576], _065798_);
  xor g_123212_(out[46], out[590], _065799_);
  xor g_123213_(out[36], out[580], _065800_);
  or g_123214_(_065799_, _065800_, _065802_);
  xor g_123215_(out[45], out[589], _065803_);
  xor g_123216_(out[35], out[579], _065804_);
  xor g_123217_(out[44], out[588], _065805_);
  xor g_123218_(out[38], out[582], _065806_);
  xor g_123219_(out[42], out[586], _065807_);
  xor g_123220_(out[37], out[581], _065808_);
  xor g_123221_(out[47], out[591], _065809_);
  xor g_123222_(out[40], out[584], _065810_);
  or g_123223_(_065803_, _065810_, _065811_);
  xor g_123224_(out[34], out[578], _065813_);
  or g_123225_(_065807_, _065813_, _065814_);
  or g_123226_(_065811_, _065814_, _065815_);
  or g_123227_(_065797_, _065804_, _065816_);
  or g_123228_(_065808_, _065816_, _065817_);
  or g_123229_(_065815_, _065817_, _065818_);
  or g_123230_(_065802_, _065818_, _065819_);
  or g_123231_(_065795_, _065805_, _065820_);
  xor g_123232_(out[39], out[583], _065821_);
  or g_123233_(_065806_, _065821_, _065822_);
  or g_123234_(_065820_, _065822_, _065824_);
  or g_123235_(_065794_, _065796_, _065825_);
  or g_123236_(_065809_, _065825_, _065826_);
  or g_123237_(_065824_, _065826_, _065827_);
  or g_123238_(_065798_, _065827_, _065828_);
  or g_123239_(_065819_, _065828_, _065829_);
  not g_123240_(_065829_, _065830_);
  xor g_123241_(out[23], out[583], _065831_);
  and g_123242_(_098063_, out[587], _065832_);
  xor g_123243_(out[30], out[590], _065833_);
  xor g_123244_(out[24], out[584], _065835_);
  xor g_123245_(out[17], out[577], _065836_);
  xor g_123246_(out[29], out[589], _065837_);
  xor g_123247_(out[25], out[585], _065838_);
  xor g_123248_(out[20], out[580], _065839_);
  xor g_123249_(out[18], out[578], _065840_);
  and g_123250_(out[27], _049565_, _065841_);
  xor g_123251_(out[19], out[579], _065842_);
  xor g_123252_(out[22], out[582], _065843_);
  xor g_123253_(out[31], out[591], _065844_);
  xor g_123254_(out[26], out[586], _065846_);
  xor g_123255_(out[21], out[581], _065847_);
  xor g_123256_(out[16], out[576], _065848_);
  or g_123257_(_065833_, _065839_, _065849_);
  or g_123258_(_065835_, _065837_, _065850_);
  or g_123259_(_065840_, _065846_, _065851_);
  or g_123260_(_065850_, _065851_, _065852_);
  or g_123261_(_065838_, _065842_, _065853_);
  or g_123262_(_065847_, _065848_, _065854_);
  or g_123263_(_065853_, _065854_, _065855_);
  or g_123264_(_065852_, _065855_, _065857_);
  xor g_123265_(out[28], out[588], _065858_);
  or g_123266_(_065832_, _065858_, _065859_);
  or g_123267_(_065831_, _065843_, _065860_);
  or g_123268_(_065859_, _065860_, _065861_);
  or g_123269_(_065836_, _065841_, _065862_);
  or g_123270_(_065844_, _065862_, _065863_);
  or g_123271_(_065861_, _065863_, _065864_);
  or g_123272_(_065857_, _065864_, _065865_);
  or g_123273_(_065849_, _065865_, _065866_);
  xor g_123274_(out[1], out[577], _065868_);
  and g_123275_(_098041_, out[587], _065869_);
  and g_123276_(out[11], _049565_, _065870_);
  xor g_123277_(out[9], out[585], _065871_);
  xor g_123278_(out[0], out[576], _065872_);
  xor g_123279_(out[14], out[590], _065873_);
  xor g_123280_(out[4], out[580], _065874_);
  or g_123281_(_065873_, _065874_, _065875_);
  xor g_123282_(out[13], out[589], _065876_);
  xor g_123283_(out[3], out[579], _065877_);
  xor g_123284_(out[12], out[588], _065879_);
  xor g_123285_(out[6], out[582], _065880_);
  xor g_123286_(out[10], out[586], _065881_);
  xor g_123287_(out[5], out[581], _065882_);
  xor g_123288_(out[15], out[591], _065883_);
  xor g_123289_(out[8], out[584], _065884_);
  or g_123290_(_065876_, _065884_, _065885_);
  xor g_123291_(out[2], out[578], _065886_);
  or g_123292_(_065881_, _065886_, _065887_);
  or g_123293_(_065885_, _065887_, _065888_);
  or g_123294_(_065871_, _065877_, _065890_);
  or g_123295_(_065882_, _065890_, _065891_);
  or g_123296_(_065888_, _065891_, _065892_);
  or g_123297_(_065875_, _065892_, _065893_);
  or g_123298_(_065869_, _065879_, _065894_);
  xor g_123299_(out[7], out[583], _065895_);
  or g_123300_(_065880_, _065895_, _065896_);
  or g_123301_(_065894_, _065896_, _065897_);
  or g_123302_(_065868_, _065870_, _065898_);
  or g_123303_(_065883_, _065898_, _065899_);
  or g_123304_(_065897_, _065899_, _065901_);
  or g_123305_(_065872_, _065901_, _065902_);
  or g_123306_(_065893_, _065902_, _065903_);
  and g_123307_(out[475], _049554_, _065904_);
  xor g_123308_(out[468], out[564], _065905_);
  xor g_123309_(out[478], out[574], _065906_);
  or g_123310_(_065905_, _065906_, _065907_);
  xor g_123311_(out[477], out[573], _065908_);
  xor g_123312_(out[467], out[563], _065909_);
  xor g_123313_(out[464], out[560], _065910_);
  and g_123314_(_049499_, out[571], _065912_);
  xor g_123315_(out[474], out[570], _065913_);
  xor g_123316_(out[479], out[575], _065914_);
  xor g_123317_(out[470], out[566], _065915_);
  xor g_123318_(out[469], out[565], _065916_);
  xor g_123319_(out[472], out[568], _065917_);
  or g_123320_(_065908_, _065917_, _065918_);
  xor g_123321_(out[466], out[562], _065919_);
  xor g_123322_(out[473], out[569], _065920_);
  xor g_123323_(out[465], out[561], _065921_);
  or g_123324_(_065913_, _065919_, _065923_);
  or g_123325_(_065918_, _065923_, _065924_);
  or g_123326_(_065909_, _065920_, _065925_);
  or g_123327_(_065916_, _065925_, _065926_);
  or g_123328_(_065924_, _065926_, _065927_);
  or g_123329_(_065907_, _065927_, _065928_);
  xor g_123330_(out[476], out[572], _065929_);
  or g_123331_(_065912_, _065929_, _065930_);
  xor g_123332_(out[471], out[567], _065931_);
  or g_123333_(_065915_, _065931_, _065932_);
  or g_123334_(_065930_, _065932_, _065934_);
  or g_123335_(_065904_, _065921_, _065935_);
  or g_123336_(_065914_, _065935_, _065936_);
  or g_123337_(_065934_, _065936_, _065937_);
  or g_123338_(_065910_, _065937_, _065938_);
  or g_123339_(_065928_, _065938_, _065939_);
  xor g_123340_(out[455], out[567], _065940_);
  and g_123341_(_049477_, out[571], _065941_);
  xor g_123342_(out[462], out[574], _065942_);
  xor g_123343_(out[456], out[568], _065943_);
  xor g_123344_(out[449], out[561], _065945_);
  xor g_123345_(out[461], out[573], _065946_);
  xor g_123346_(out[457], out[569], _065947_);
  xor g_123347_(out[452], out[564], _065948_);
  xor g_123348_(out[450], out[562], _065949_);
  and g_123349_(out[459], _049554_, _065950_);
  xor g_123350_(out[451], out[563], _065951_);
  xor g_123351_(out[454], out[566], _065952_);
  xor g_123352_(out[463], out[575], _065953_);
  xor g_123353_(out[458], out[570], _065954_);
  xor g_123354_(out[453], out[565], _065956_);
  xor g_123355_(out[448], out[560], _065957_);
  or g_123356_(_065942_, _065948_, _065958_);
  or g_123357_(_065943_, _065946_, _065959_);
  or g_123358_(_065949_, _065954_, _065960_);
  or g_123359_(_065959_, _065960_, _065961_);
  or g_123360_(_065947_, _065951_, _065962_);
  or g_123361_(_065956_, _065957_, _065963_);
  or g_123362_(_065962_, _065963_, _065964_);
  or g_123363_(_065961_, _065964_, _065965_);
  xor g_123364_(out[460], out[572], _065967_);
  or g_123365_(_065941_, _065967_, _065968_);
  or g_123366_(_065940_, _065952_, _065969_);
  or g_123367_(_065968_, _065969_, _065970_);
  or g_123368_(_065945_, _065950_, _065971_);
  or g_123369_(_065953_, _065971_, _065972_);
  or g_123370_(_065970_, _065972_, _065973_);
  or g_123371_(_065965_, _065973_, _065974_);
  or g_123372_(_065958_, _065974_, _065975_);
  xor g_123373_(out[433], out[561], _065976_);
  and g_123374_(_049466_, out[571], _065978_);
  and g_123375_(out[443], _049554_, _065979_);
  xor g_123376_(out[445], out[573], _065980_);
  xor g_123377_(out[442], out[570], _065981_);
  xor g_123378_(out[436], out[564], _065982_);
  xor g_123379_(out[446], out[574], _065983_);
  or g_123380_(_065982_, _065983_, _065984_);
  xor g_123381_(out[440], out[568], _065985_);
  xor g_123382_(out[432], out[560], _065986_);
  xor g_123383_(out[434], out[562], _065987_);
  xor g_123384_(out[441], out[569], _065989_);
  xor g_123385_(out[437], out[565], _065990_);
  xor g_123386_(out[435], out[563], _065991_);
  xor g_123387_(out[447], out[575], _065992_);
  xor g_123388_(out[438], out[566], _065993_);
  or g_123389_(_065980_, _065985_, _065994_);
  or g_123390_(_065981_, _065987_, _065995_);
  or g_123391_(_065994_, _065995_, _065996_);
  or g_123392_(_065989_, _065991_, _065997_);
  or g_123393_(_065986_, _065990_, _065998_);
  or g_123394_(_065997_, _065998_, _066000_);
  or g_123395_(_065996_, _066000_, _066001_);
  xor g_123396_(out[444], out[572], _066002_);
  or g_123397_(_065978_, _066002_, _066003_);
  xor g_123398_(out[439], out[567], _066004_);
  or g_123399_(_065993_, _066004_, _066005_);
  or g_123400_(_066003_, _066005_, _066006_);
  or g_123401_(_065976_, _065979_, _066007_);
  or g_123402_(_065992_, _066007_, _066008_);
  or g_123403_(_066006_, _066008_, _066009_);
  or g_123404_(_066001_, _066009_, _066011_);
  or g_123405_(_065984_, _066011_, _066012_);
  not g_123406_(_066012_, _066013_);
  xor g_123407_(out[423], out[567], _066014_);
  and g_123408_(_049455_, out[571], _066015_);
  xor g_123409_(out[430], out[574], _066016_);
  xor g_123410_(out[424], out[568], _066017_);
  xor g_123411_(out[417], out[561], _066018_);
  xor g_123412_(out[429], out[573], _066019_);
  xor g_123413_(out[425], out[569], _066020_);
  xor g_123414_(out[420], out[564], _066022_);
  xor g_123415_(out[418], out[562], _066023_);
  and g_123416_(out[427], _049554_, _066024_);
  xor g_123417_(out[419], out[563], _066025_);
  xor g_123418_(out[422], out[566], _066026_);
  xor g_123419_(out[431], out[575], _066027_);
  xor g_123420_(out[426], out[570], _066028_);
  xor g_123421_(out[421], out[565], _066029_);
  xor g_123422_(out[416], out[560], _066030_);
  or g_123423_(_066016_, _066022_, _066031_);
  or g_123424_(_066017_, _066019_, _066033_);
  or g_123425_(_066023_, _066028_, _066034_);
  or g_123426_(_066033_, _066034_, _066035_);
  or g_123427_(_066020_, _066025_, _066036_);
  or g_123428_(_066029_, _066030_, _066037_);
  or g_123429_(_066036_, _066037_, _066038_);
  or g_123430_(_066035_, _066038_, _066039_);
  xor g_123431_(out[428], out[572], _066040_);
  or g_123432_(_066015_, _066040_, _066041_);
  or g_123433_(_066014_, _066026_, _066042_);
  or g_123434_(_066041_, _066042_, _066044_);
  or g_123435_(_066018_, _066024_, _066045_);
  or g_123436_(_066027_, _066045_, _066046_);
  or g_123437_(_066044_, _066046_, _066047_);
  or g_123438_(_066039_, _066047_, _066048_);
  or g_123439_(_066031_, _066048_, _066049_);
  not g_123440_(_066049_, _066050_);
  xor g_123441_(out[401], out[561], _066051_);
  and g_123442_(out[411], _049554_, _066052_);
  xor g_123443_(out[409], out[569], _066053_);
  xor g_123444_(out[400], out[560], _066055_);
  xor g_123445_(out[414], out[574], _066056_);
  xor g_123446_(out[404], out[564], _066057_);
  or g_123447_(_066056_, _066057_, _066058_);
  xor g_123448_(out[413], out[573], _066059_);
  xor g_123449_(out[403], out[563], _066060_);
  and g_123450_(_049444_, out[571], _066061_);
  xor g_123451_(out[406], out[566], _066062_);
  xor g_123452_(out[410], out[570], _066063_);
  xor g_123453_(out[405], out[565], _066064_);
  xor g_123454_(out[415], out[575], _066066_);
  xor g_123455_(out[408], out[568], _066067_);
  or g_123456_(_066059_, _066067_, _066068_);
  xor g_123457_(out[402], out[562], _066069_);
  or g_123458_(_066063_, _066069_, _066070_);
  or g_123459_(_066068_, _066070_, _066071_);
  or g_123460_(_066053_, _066060_, _066072_);
  or g_123461_(_066064_, _066072_, _066073_);
  or g_123462_(_066071_, _066073_, _066074_);
  or g_123463_(_066058_, _066074_, _066075_);
  xor g_123464_(out[412], out[572], _066077_);
  or g_123465_(_066061_, _066077_, _066078_);
  xor g_123466_(out[407], out[567], _066079_);
  or g_123467_(_066062_, _066079_, _066080_);
  or g_123468_(_066078_, _066080_, _066081_);
  or g_123469_(_066051_, _066052_, _066082_);
  or g_123470_(_066066_, _066082_, _066083_);
  or g_123471_(_066081_, _066083_, _066084_);
  or g_123472_(_066055_, _066084_, _066085_);
  or g_123473_(_066075_, _066085_, _066086_);
  xor g_123474_(out[391], out[567], _066088_);
  and g_123475_(_049433_, out[571], _066089_);
  xor g_123476_(out[398], out[574], _066090_);
  xor g_123477_(out[392], out[568], _066091_);
  xor g_123478_(out[385], out[561], _066092_);
  xor g_123479_(out[397], out[573], _066093_);
  xor g_123480_(out[393], out[569], _066094_);
  xor g_123481_(out[388], out[564], _066095_);
  xor g_123482_(out[386], out[562], _066096_);
  and g_123483_(out[395], _049554_, _066097_);
  xor g_123484_(out[387], out[563], _066099_);
  xor g_123485_(out[390], out[566], _066100_);
  xor g_123486_(out[399], out[575], _066101_);
  xor g_123487_(out[394], out[570], _066102_);
  xor g_123488_(out[389], out[565], _066103_);
  xor g_123489_(out[384], out[560], _066104_);
  or g_123490_(_066090_, _066095_, _066105_);
  or g_123491_(_066091_, _066093_, _066106_);
  or g_123492_(_066096_, _066102_, _066107_);
  or g_123493_(_066106_, _066107_, _066108_);
  or g_123494_(_066094_, _066099_, _066110_);
  or g_123495_(_066103_, _066104_, _066111_);
  or g_123496_(_066110_, _066111_, _066112_);
  or g_123497_(_066108_, _066112_, _066113_);
  xor g_123498_(out[396], out[572], _066114_);
  or g_123499_(_066089_, _066114_, _066115_);
  or g_123500_(_066088_, _066100_, _066116_);
  or g_123501_(_066115_, _066116_, _066117_);
  or g_123502_(_066092_, _066097_, _066118_);
  or g_123503_(_066101_, _066118_, _066119_);
  or g_123504_(_066117_, _066119_, _066121_);
  or g_123505_(_066113_, _066121_, _066122_);
  or g_123506_(_066105_, _066122_, _066123_);
  xor g_123507_(out[369], out[561], _066124_);
  and g_123508_(out[379], _049554_, _066125_);
  xor g_123509_(out[377], out[569], _066126_);
  xor g_123510_(out[368], out[560], _066127_);
  xor g_123511_(out[382], out[574], _066128_);
  xor g_123512_(out[372], out[564], _066129_);
  or g_123513_(_066128_, _066129_, _066130_);
  xor g_123514_(out[381], out[573], _066132_);
  xor g_123515_(out[371], out[563], _066133_);
  and g_123516_(_049422_, out[571], _066134_);
  xor g_123517_(out[374], out[566], _066135_);
  xor g_123518_(out[378], out[570], _066136_);
  xor g_123519_(out[373], out[565], _066137_);
  xor g_123520_(out[383], out[575], _066138_);
  xor g_123521_(out[376], out[568], _066139_);
  or g_123522_(_066132_, _066139_, _066140_);
  xor g_123523_(out[370], out[562], _066141_);
  or g_123524_(_066136_, _066141_, _066143_);
  or g_123525_(_066140_, _066143_, _066144_);
  or g_123526_(_066126_, _066133_, _066145_);
  or g_123527_(_066137_, _066145_, _066146_);
  or g_123528_(_066144_, _066146_, _066147_);
  or g_123529_(_066130_, _066147_, _066148_);
  xor g_123530_(out[380], out[572], _066149_);
  or g_123531_(_066134_, _066149_, _066150_);
  xor g_123532_(out[375], out[567], _066151_);
  or g_123533_(_066135_, _066151_, _066152_);
  or g_123534_(_066150_, _066152_, _066154_);
  or g_123535_(_066124_, _066125_, _066155_);
  or g_123536_(_066138_, _066155_, _066156_);
  or g_123537_(_066154_, _066156_, _066157_);
  or g_123538_(_066127_, _066157_, _066158_);
  or g_123539_(_066148_, _066158_, _066159_);
  not g_123540_(_066159_, _066160_);
  xor g_123541_(out[359], out[567], _066161_);
  and g_123542_(_049411_, out[571], _066162_);
  xor g_123543_(out[366], out[574], _066163_);
  xor g_123544_(out[360], out[568], _066165_);
  xor g_123545_(out[353], out[561], _066166_);
  xor g_123546_(out[365], out[573], _066167_);
  xor g_123547_(out[361], out[569], _066168_);
  xor g_123548_(out[356], out[564], _066169_);
  xor g_123549_(out[354], out[562], _066170_);
  and g_123550_(out[363], _049554_, _066171_);
  xor g_123551_(out[355], out[563], _066172_);
  xor g_123552_(out[358], out[566], _066173_);
  xor g_123553_(out[367], out[575], _066174_);
  xor g_123554_(out[362], out[570], _066176_);
  xor g_123555_(out[357], out[565], _066177_);
  xor g_123556_(out[352], out[560], _066178_);
  or g_123557_(_066163_, _066169_, _066179_);
  or g_123558_(_066165_, _066167_, _066180_);
  or g_123559_(_066170_, _066176_, _066181_);
  or g_123560_(_066180_, _066181_, _066182_);
  or g_123561_(_066168_, _066172_, _066183_);
  or g_123562_(_066177_, _066178_, _066184_);
  or g_123563_(_066183_, _066184_, _066185_);
  or g_123564_(_066182_, _066185_, _066187_);
  xor g_123565_(out[364], out[572], _066188_);
  or g_123566_(_066162_, _066188_, _066189_);
  or g_123567_(_066161_, _066173_, _066190_);
  or g_123568_(_066189_, _066190_, _066191_);
  or g_123569_(_066166_, _066171_, _066192_);
  or g_123570_(_066174_, _066192_, _066193_);
  or g_123571_(_066191_, _066193_, _066194_);
  or g_123572_(_066187_, _066194_, _066195_);
  or g_123573_(_066179_, _066195_, _066196_);
  not g_123574_(_066196_, _066198_);
  xor g_123575_(out[337], out[561], _066199_);
  and g_123576_(out[347], _049554_, _066200_);
  xor g_123577_(out[345], out[569], _066201_);
  xor g_123578_(out[336], out[560], _066202_);
  xor g_123579_(out[350], out[574], _066203_);
  xor g_123580_(out[340], out[564], _066204_);
  or g_123581_(_066203_, _066204_, _066205_);
  xor g_123582_(out[349], out[573], _066206_);
  xor g_123583_(out[339], out[563], _066207_);
  and g_123584_(_049400_, out[571], _066209_);
  xor g_123585_(out[342], out[566], _066210_);
  xor g_123586_(out[346], out[570], _066211_);
  xor g_123587_(out[341], out[565], _066212_);
  xor g_123588_(out[351], out[575], _066213_);
  xor g_123589_(out[344], out[568], _066214_);
  or g_123590_(_066206_, _066214_, _066215_);
  xor g_123591_(out[338], out[562], _066216_);
  or g_123592_(_066211_, _066216_, _066217_);
  or g_123593_(_066215_, _066217_, _066218_);
  or g_123594_(_066201_, _066207_, _066220_);
  or g_123595_(_066212_, _066220_, _066221_);
  or g_123596_(_066218_, _066221_, _066222_);
  or g_123597_(_066205_, _066222_, _066223_);
  xor g_123598_(out[348], out[572], _066224_);
  or g_123599_(_066209_, _066224_, _066225_);
  xor g_123600_(out[343], out[567], _066226_);
  or g_123601_(_066210_, _066226_, _066227_);
  or g_123602_(_066225_, _066227_, _066228_);
  or g_123603_(_066199_, _066200_, _066229_);
  or g_123604_(_066213_, _066229_, _066231_);
  or g_123605_(_066228_, _066231_, _066232_);
  or g_123606_(_066202_, _066232_, _066233_);
  or g_123607_(_066223_, _066233_, _066234_);
  xor g_123608_(out[327], out[567], _066235_);
  and g_123609_(_098294_, out[571], _066236_);
  xor g_123610_(out[334], out[574], _066237_);
  xor g_123611_(out[328], out[568], _066238_);
  xor g_123612_(out[321], out[561], _066239_);
  xor g_123613_(out[333], out[573], _066240_);
  xor g_123614_(out[329], out[569], _066242_);
  xor g_123615_(out[324], out[564], _066243_);
  xor g_123616_(out[322], out[562], _066244_);
  and g_123617_(out[331], _049554_, _066245_);
  xor g_123618_(out[323], out[563], _066246_);
  xor g_123619_(out[326], out[566], _066247_);
  xor g_123620_(out[335], out[575], _066248_);
  xor g_123621_(out[330], out[570], _066249_);
  xor g_123622_(out[325], out[565], _066250_);
  xor g_123623_(out[320], out[560], _066251_);
  or g_123624_(_066237_, _066243_, _066253_);
  or g_123625_(_066238_, _066240_, _066254_);
  or g_123626_(_066244_, _066249_, _066255_);
  or g_123627_(_066254_, _066255_, _066256_);
  or g_123628_(_066242_, _066246_, _066257_);
  or g_123629_(_066250_, _066251_, _066258_);
  or g_123630_(_066257_, _066258_, _066259_);
  or g_123631_(_066256_, _066259_, _066260_);
  xor g_123632_(out[332], out[572], _066261_);
  or g_123633_(_066236_, _066261_, _066262_);
  or g_123634_(_066235_, _066247_, _066264_);
  or g_123635_(_066262_, _066264_, _066265_);
  or g_123636_(_066239_, _066245_, _066266_);
  or g_123637_(_066248_, _066266_, _066267_);
  or g_123638_(_066265_, _066267_, _066268_);
  or g_123639_(_066260_, _066268_, _066269_);
  or g_123640_(_066253_, _066269_, _066270_);
  and g_123641_(out[315], _049554_, _066271_);
  xor g_123642_(out[308], out[564], _066272_);
  xor g_123643_(out[318], out[574], _066273_);
  or g_123644_(_066272_, _066273_, _066275_);
  xor g_123645_(out[317], out[573], _066276_);
  xor g_123646_(out[307], out[563], _066277_);
  xor g_123647_(out[304], out[560], _066278_);
  and g_123648_(_098283_, out[571], _066279_);
  xor g_123649_(out[314], out[570], _066280_);
  xor g_123650_(out[319], out[575], _066281_);
  xor g_123651_(out[310], out[566], _066282_);
  xor g_123652_(out[309], out[565], _066283_);
  xor g_123653_(out[312], out[568], _066284_);
  or g_123654_(_066276_, _066284_, _066286_);
  xor g_123655_(out[306], out[562], _066287_);
  xor g_123656_(out[313], out[569], _066288_);
  xor g_123657_(out[305], out[561], _066289_);
  or g_123658_(_066280_, _066287_, _066290_);
  or g_123659_(_066286_, _066290_, _066291_);
  or g_123660_(_066277_, _066288_, _066292_);
  or g_123661_(_066283_, _066292_, _066293_);
  or g_123662_(_066291_, _066293_, _066294_);
  or g_123663_(_066275_, _066294_, _066295_);
  xor g_123664_(out[316], out[572], _066297_);
  or g_123665_(_066279_, _066297_, _066298_);
  xor g_123666_(out[311], out[567], _066299_);
  or g_123667_(_066282_, _066299_, _066300_);
  or g_123668_(_066298_, _066300_, _066301_);
  or g_123669_(_066271_, _066289_, _066302_);
  or g_123670_(_066281_, _066302_, _066303_);
  or g_123671_(_066301_, _066303_, _066304_);
  or g_123672_(_066278_, _066304_, _066305_);
  or g_123673_(_066295_, _066305_, _066306_);
  xor g_123674_(out[295], out[567], _066308_);
  and g_123675_(_098272_, out[571], _066309_);
  xor g_123676_(out[302], out[574], _066310_);
  xor g_123677_(out[296], out[568], _066311_);
  xor g_123678_(out[289], out[561], _066312_);
  xor g_123679_(out[301], out[573], _066313_);
  xor g_123680_(out[297], out[569], _066314_);
  xor g_123681_(out[292], out[564], _066315_);
  xor g_123682_(out[290], out[562], _066316_);
  and g_123683_(out[299], _049554_, _066317_);
  xor g_123684_(out[291], out[563], _066319_);
  xor g_123685_(out[294], out[566], _066320_);
  xor g_123686_(out[303], out[575], _066321_);
  xor g_123687_(out[298], out[570], _066322_);
  xor g_123688_(out[293], out[565], _066323_);
  xor g_123689_(out[288], out[560], _066324_);
  or g_123690_(_066310_, _066315_, _066325_);
  or g_123691_(_066311_, _066313_, _066326_);
  or g_123692_(_066316_, _066322_, _066327_);
  or g_123693_(_066326_, _066327_, _066328_);
  or g_123694_(_066314_, _066319_, _066330_);
  or g_123695_(_066323_, _066324_, _066331_);
  or g_123696_(_066330_, _066331_, _066332_);
  or g_123697_(_066328_, _066332_, _066333_);
  xor g_123698_(out[300], out[572], _066334_);
  or g_123699_(_066309_, _066334_, _066335_);
  or g_123700_(_066308_, _066320_, _066336_);
  or g_123701_(_066335_, _066336_, _066337_);
  or g_123702_(_066312_, _066317_, _066338_);
  or g_123703_(_066321_, _066338_, _066339_);
  or g_123704_(_066337_, _066339_, _066341_);
  or g_123705_(_066333_, _066341_, _066342_);
  or g_123706_(_066325_, _066342_, _066343_);
  xor g_123707_(out[276], out[564], _066344_);
  xor g_123708_(out[284], out[572], _066345_);
  and g_123709_(_098261_, out[571], _066346_);
  xor g_123710_(out[282], out[570], _066347_);
  xor g_123711_(out[278], out[566], _066348_);
  xor g_123712_(out[277], out[565], _066349_);
  xor g_123713_(out[275], out[563], _066350_);
  xor g_123714_(out[285], out[573], _066352_);
  xor g_123715_(out[286], out[574], _066353_);
  xor g_123716_(out[273], out[561], _066354_);
  xor g_123717_(out[274], out[562], _066355_);
  and g_123718_(out[283], _049554_, _066356_);
  xor g_123719_(out[272], out[560], _066357_);
  xor g_123720_(out[287], out[575], _066358_);
  xor g_123721_(out[280], out[568], _066359_);
  or g_123722_(_066352_, _066359_, _066360_);
  xor g_123723_(out[281], out[569], _066361_);
  or g_123724_(_066347_, _066355_, _066363_);
  or g_123725_(_066360_, _066363_, _066364_);
  or g_123726_(_066350_, _066361_, _066365_);
  or g_123727_(_066349_, _066365_, _066366_);
  or g_123728_(_066364_, _066366_, _066367_);
  or g_123729_(_066344_, _066353_, _066368_);
  or g_123730_(_066367_, _066368_, _066369_);
  or g_123731_(_066345_, _066346_, _066370_);
  xor g_123732_(out[279], out[567], _066371_);
  or g_123733_(_066348_, _066371_, _066372_);
  or g_123734_(_066370_, _066372_, _066374_);
  or g_123735_(_066354_, _066356_, _066375_);
  or g_123736_(_066358_, _066375_, _066376_);
  or g_123737_(_066374_, _066376_, _066377_);
  or g_123738_(_066357_, _066377_, _066378_);
  or g_123739_(_066369_, _066378_, _066379_);
  not g_123740_(_066379_, _066380_);
  xor g_123741_(out[263], out[567], _066381_);
  and g_123742_(_098250_, out[571], _066382_);
  xor g_123743_(out[270], out[574], _066383_);
  xor g_123744_(out[264], out[568], _066385_);
  xor g_123745_(out[257], out[561], _066386_);
  xor g_123746_(out[269], out[573], _066387_);
  xor g_123747_(out[265], out[569], _066388_);
  xor g_123748_(out[260], out[564], _066389_);
  xor g_123749_(out[258], out[562], _066390_);
  and g_123750_(out[267], _049554_, _066391_);
  xor g_123751_(out[259], out[563], _066392_);
  xor g_123752_(out[262], out[566], _066393_);
  xor g_123753_(out[271], out[575], _066394_);
  xor g_123754_(out[266], out[570], _066396_);
  xor g_123755_(out[261], out[565], _066397_);
  xor g_123756_(out[256], out[560], _066398_);
  or g_123757_(_066383_, _066389_, _066399_);
  or g_123758_(_066385_, _066387_, _066400_);
  or g_123759_(_066390_, _066396_, _066401_);
  or g_123760_(_066400_, _066401_, _066402_);
  or g_123761_(_066388_, _066392_, _066403_);
  or g_123762_(_066397_, _066398_, _066404_);
  or g_123763_(_066403_, _066404_, _066405_);
  or g_123764_(_066402_, _066405_, _066407_);
  xor g_123765_(out[268], out[572], _066408_);
  or g_123766_(_066382_, _066408_, _066409_);
  or g_123767_(_066381_, _066393_, _066410_);
  or g_123768_(_066409_, _066410_, _066411_);
  or g_123769_(_066386_, _066391_, _066412_);
  or g_123770_(_066394_, _066412_, _066413_);
  or g_123771_(_066411_, _066413_, _066414_);
  or g_123772_(_066407_, _066414_, _066415_);
  or g_123773_(_066399_, _066415_, _066416_);
  xor g_123774_(out[241], out[561], _066418_);
  and g_123775_(out[251], _049554_, _066419_);
  xor g_123776_(out[249], out[569], _066420_);
  xor g_123777_(out[240], out[560], _066421_);
  xor g_123778_(out[254], out[574], _066422_);
  xor g_123779_(out[244], out[564], _066423_);
  or g_123780_(_066422_, _066423_, _066424_);
  xor g_123781_(out[253], out[573], _066425_);
  xor g_123782_(out[243], out[563], _066426_);
  and g_123783_(_098239_, out[571], _066427_);
  xor g_123784_(out[246], out[566], _066429_);
  xor g_123785_(out[250], out[570], _066430_);
  xor g_123786_(out[245], out[565], _066431_);
  xor g_123787_(out[255], out[575], _066432_);
  xor g_123788_(out[248], out[568], _066433_);
  or g_123789_(_066425_, _066433_, _066434_);
  xor g_123790_(out[242], out[562], _066435_);
  or g_123791_(_066430_, _066435_, _066436_);
  or g_123792_(_066434_, _066436_, _066437_);
  or g_123793_(_066420_, _066426_, _066438_);
  or g_123794_(_066431_, _066438_, _066440_);
  or g_123795_(_066437_, _066440_, _066441_);
  or g_123796_(_066424_, _066441_, _066442_);
  xor g_123797_(out[252], out[572], _066443_);
  or g_123798_(_066427_, _066443_, _066444_);
  xor g_123799_(out[247], out[567], _066445_);
  or g_123800_(_066429_, _066445_, _066446_);
  or g_123801_(_066444_, _066446_, _066447_);
  or g_123802_(_066418_, _066419_, _066448_);
  or g_123803_(_066432_, _066448_, _066449_);
  or g_123804_(_066447_, _066449_, _066451_);
  or g_123805_(_066421_, _066451_, _066452_);
  or g_123806_(_066442_, _066452_, _066453_);
  xor g_123807_(out[231], out[567], _066454_);
  and g_123808_(_098228_, out[571], _066455_);
  xor g_123809_(out[238], out[574], _066456_);
  xor g_123810_(out[232], out[568], _066457_);
  xor g_123811_(out[225], out[561], _066458_);
  xor g_123812_(out[237], out[573], _066459_);
  xor g_123813_(out[233], out[569], _066460_);
  xor g_123814_(out[228], out[564], _066462_);
  xor g_123815_(out[226], out[562], _066463_);
  and g_123816_(out[235], _049554_, _066464_);
  xor g_123817_(out[227], out[563], _066465_);
  xor g_123818_(out[230], out[566], _066466_);
  xor g_123819_(out[239], out[575], _066467_);
  xor g_123820_(out[234], out[570], _066468_);
  xor g_123821_(out[229], out[565], _066469_);
  xor g_123822_(out[224], out[560], _066470_);
  or g_123823_(_066456_, _066462_, _066471_);
  or g_123824_(_066457_, _066459_, _066473_);
  or g_123825_(_066463_, _066468_, _066474_);
  or g_123826_(_066473_, _066474_, _066475_);
  or g_123827_(_066460_, _066465_, _066476_);
  or g_123828_(_066469_, _066470_, _066477_);
  or g_123829_(_066476_, _066477_, _066478_);
  or g_123830_(_066475_, _066478_, _066479_);
  xor g_123831_(out[236], out[572], _066480_);
  or g_123832_(_066455_, _066480_, _066481_);
  or g_123833_(_066454_, _066466_, _066482_);
  or g_123834_(_066481_, _066482_, _066484_);
  or g_123835_(_066458_, _066464_, _066485_);
  or g_123836_(_066467_, _066485_, _066486_);
  or g_123837_(_066484_, _066486_, _066487_);
  or g_123838_(_066479_, _066487_, _066488_);
  or g_123839_(_066471_, _066488_, _066489_);
  xor g_123840_(out[218], out[570], _066490_);
  xor g_123841_(out[210], out[562], _066491_);
  xor g_123842_(out[209], out[561], _066492_);
  and g_123843_(_098217_, out[571], _066493_);
  and g_123844_(out[219], _049554_, _066495_);
  xor g_123845_(out[221], out[573], _066496_);
  xor g_123846_(out[211], out[563], _066497_);
  xor g_123847_(out[222], out[574], _066498_);
  xor g_123848_(out[220], out[572], _066499_);
  xor g_123849_(out[216], out[568], _066500_);
  xor g_123850_(out[223], out[575], _066501_);
  xor g_123851_(out[213], out[565], _066502_);
  xor g_123852_(out[214], out[566], _066503_);
  xor g_123853_(out[208], out[560], _066504_);
  xor g_123854_(out[212], out[564], _066506_);
  or g_123855_(_066496_, _066500_, _066507_);
  xor g_123856_(out[217], out[569], _066508_);
  or g_123857_(_066490_, _066491_, _066509_);
  or g_123858_(_066507_, _066509_, _066510_);
  or g_123859_(_066497_, _066508_, _066511_);
  or g_123860_(_066502_, _066511_, _066512_);
  or g_123861_(_066510_, _066512_, _066513_);
  or g_123862_(_066498_, _066506_, _066514_);
  or g_123863_(_066513_, _066514_, _066515_);
  or g_123864_(_066493_, _066499_, _066517_);
  xor g_123865_(out[215], out[567], _066518_);
  or g_123866_(_066503_, _066518_, _066519_);
  or g_123867_(_066517_, _066519_, _066520_);
  or g_123868_(_066492_, _066495_, _066521_);
  or g_123869_(_066501_, _066521_, _066522_);
  or g_123870_(_066520_, _066522_, _066523_);
  or g_123871_(_066504_, _066523_, _066524_);
  or g_123872_(_066515_, _066524_, _066525_);
  xor g_123873_(out[199], out[567], _066526_);
  and g_123874_(_098206_, out[571], _066528_);
  xor g_123875_(out[206], out[574], _066529_);
  xor g_123876_(out[200], out[568], _066530_);
  xor g_123877_(out[193], out[561], _066531_);
  xor g_123878_(out[205], out[573], _066532_);
  xor g_123879_(out[201], out[569], _066533_);
  xor g_123880_(out[196], out[564], _066534_);
  xor g_123881_(out[194], out[562], _066535_);
  and g_123882_(out[203], _049554_, _066536_);
  xor g_123883_(out[195], out[563], _066537_);
  xor g_123884_(out[198], out[566], _066539_);
  xor g_123885_(out[207], out[575], _066540_);
  xor g_123886_(out[202], out[570], _066541_);
  xor g_123887_(out[197], out[565], _066542_);
  xor g_123888_(out[192], out[560], _066543_);
  or g_123889_(_066529_, _066534_, _066544_);
  or g_123890_(_066530_, _066532_, _066545_);
  or g_123891_(_066535_, _066541_, _066546_);
  or g_123892_(_066545_, _066546_, _066547_);
  or g_123893_(_066533_, _066537_, _066548_);
  or g_123894_(_066542_, _066543_, _066550_);
  or g_123895_(_066548_, _066550_, _066551_);
  or g_123896_(_066547_, _066551_, _066552_);
  xor g_123897_(out[204], out[572], _066553_);
  or g_123898_(_066528_, _066553_, _066554_);
  or g_123899_(_066526_, _066539_, _066555_);
  or g_123900_(_066554_, _066555_, _066556_);
  or g_123901_(_066531_, _066536_, _066557_);
  or g_123902_(_066540_, _066557_, _066558_);
  or g_123903_(_066556_, _066558_, _066559_);
  or g_123904_(_066552_, _066559_, _066561_);
  or g_123905_(_066544_, _066561_, _066562_);
  xor g_123906_(out[189], out[573], _066563_);
  xor g_123907_(out[178], out[562], _066564_);
  xor g_123908_(out[181], out[565], _066565_);
  xor g_123909_(out[185], out[569], _066566_);
  xor g_123910_(out[180], out[564], _066567_);
  xor g_123911_(out[184], out[568], _066568_);
  xor g_123912_(out[190], out[574], _066569_);
  xor g_123913_(out[182], out[566], _066570_);
  xor g_123914_(out[191], out[575], _066572_);
  xor g_123915_(out[186], out[570], _066573_);
  xor g_123916_(out[176], out[560], _066574_);
  xor g_123917_(out[179], out[563], _066575_);
  and g_123918_(_098195_, out[571], _066576_);
  and g_123919_(out[187], _049554_, _066577_);
  xor g_123920_(out[177], out[561], _066578_);
  or g_123921_(_066567_, _066569_, _066579_);
  or g_123922_(_066563_, _066568_, _066580_);
  or g_123923_(_066564_, _066573_, _066581_);
  or g_123924_(_066580_, _066581_, _066583_);
  or g_123925_(_066566_, _066575_, _066584_);
  or g_123926_(_066565_, _066574_, _066585_);
  or g_123927_(_066584_, _066585_, _066586_);
  or g_123928_(_066583_, _066586_, _066587_);
  xor g_123929_(out[188], out[572], _066588_);
  or g_123930_(_066576_, _066588_, _066589_);
  xor g_123931_(out[183], out[567], _066590_);
  or g_123932_(_066570_, _066590_, _066591_);
  or g_123933_(_066589_, _066591_, _066592_);
  or g_123934_(_066577_, _066578_, _066594_);
  or g_123935_(_066572_, _066594_, _066595_);
  or g_123936_(_066592_, _066595_, _066596_);
  or g_123937_(_066587_, _066596_, _066597_);
  or g_123938_(_066579_, _066597_, _066598_);
  xor g_123939_(out[167], out[567], _066599_);
  and g_123940_(_098184_, out[571], _066600_);
  xor g_123941_(out[174], out[574], _066601_);
  xor g_123942_(out[168], out[568], _066602_);
  xor g_123943_(out[161], out[561], _066603_);
  xor g_123944_(out[173], out[573], _066605_);
  xor g_123945_(out[169], out[569], _066606_);
  xor g_123946_(out[164], out[564], _066607_);
  xor g_123947_(out[162], out[562], _066608_);
  and g_123948_(out[171], _049554_, _066609_);
  xor g_123949_(out[163], out[563], _066610_);
  xor g_123950_(out[166], out[566], _066611_);
  xor g_123951_(out[175], out[575], _066612_);
  xor g_123952_(out[170], out[570], _066613_);
  xor g_123953_(out[165], out[565], _066614_);
  xor g_123954_(out[160], out[560], _066616_);
  or g_123955_(_066601_, _066607_, _066617_);
  or g_123956_(_066602_, _066605_, _066618_);
  or g_123957_(_066608_, _066613_, _066619_);
  or g_123958_(_066618_, _066619_, _066620_);
  or g_123959_(_066606_, _066610_, _066621_);
  or g_123960_(_066614_, _066616_, _066622_);
  or g_123961_(_066621_, _066622_, _066623_);
  or g_123962_(_066620_, _066623_, _066624_);
  xor g_123963_(out[172], out[572], _066625_);
  or g_123964_(_066600_, _066625_, _066627_);
  or g_123965_(_066599_, _066611_, _066628_);
  or g_123966_(_066627_, _066628_, _066629_);
  or g_123967_(_066603_, _066609_, _066630_);
  or g_123968_(_066612_, _066630_, _066631_);
  or g_123969_(_066629_, _066631_, _066632_);
  or g_123970_(_066624_, _066632_, _066633_);
  or g_123971_(_066617_, _066633_, _066634_);
  not g_123972_(_066634_, _066635_);
  xor g_123973_(out[145], out[561], _066636_);
  and g_123974_(out[155], _049554_, _066638_);
  xor g_123975_(out[153], out[569], _066639_);
  xor g_123976_(out[144], out[560], _066640_);
  xor g_123977_(out[158], out[574], _066641_);
  xor g_123978_(out[148], out[564], _066642_);
  or g_123979_(_066641_, _066642_, _066643_);
  xor g_123980_(out[157], out[573], _066644_);
  xor g_123981_(out[147], out[563], _066645_);
  and g_123982_(_098173_, out[571], _066646_);
  xor g_123983_(out[150], out[566], _066647_);
  xor g_123984_(out[154], out[570], _066649_);
  xor g_123985_(out[149], out[565], _066650_);
  xor g_123986_(out[159], out[575], _066651_);
  xor g_123987_(out[152], out[568], _066652_);
  or g_123988_(_066644_, _066652_, _066653_);
  xor g_123989_(out[146], out[562], _066654_);
  or g_123990_(_066649_, _066654_, _066655_);
  or g_123991_(_066653_, _066655_, _066656_);
  or g_123992_(_066639_, _066645_, _066657_);
  or g_123993_(_066650_, _066657_, _066658_);
  or g_123994_(_066656_, _066658_, _066660_);
  or g_123995_(_066643_, _066660_, _066661_);
  xor g_123996_(out[156], out[572], _066662_);
  or g_123997_(_066646_, _066662_, _066663_);
  xor g_123998_(out[151], out[567], _066664_);
  or g_123999_(_066647_, _066664_, _066665_);
  or g_124000_(_066663_, _066665_, _066666_);
  or g_124001_(_066636_, _066638_, _066667_);
  or g_124002_(_066651_, _066667_, _066668_);
  or g_124003_(_066666_, _066668_, _066669_);
  or g_124004_(_066640_, _066669_, _066671_);
  or g_124005_(_066661_, _066671_, _066672_);
  xor g_124006_(out[135], out[567], _066673_);
  and g_124007_(_098162_, out[571], _066674_);
  xor g_124008_(out[142], out[574], _066675_);
  xor g_124009_(out[136], out[568], _066676_);
  xor g_124010_(out[129], out[561], _066677_);
  xor g_124011_(out[141], out[573], _066678_);
  xor g_124012_(out[137], out[569], _066679_);
  xor g_124013_(out[132], out[564], _066680_);
  xor g_124014_(out[130], out[562], _066682_);
  and g_124015_(out[139], _049554_, _066683_);
  xor g_124016_(out[131], out[563], _066684_);
  xor g_124017_(out[134], out[566], _066685_);
  xor g_124018_(out[143], out[575], _066686_);
  xor g_124019_(out[138], out[570], _066687_);
  xor g_124020_(out[133], out[565], _066688_);
  xor g_124021_(out[128], out[560], _066689_);
  or g_124022_(_066675_, _066680_, _066690_);
  or g_124023_(_066676_, _066678_, _066691_);
  or g_124024_(_066682_, _066687_, _066693_);
  or g_124025_(_066691_, _066693_, _066694_);
  or g_124026_(_066679_, _066684_, _066695_);
  or g_124027_(_066688_, _066689_, _066696_);
  or g_124028_(_066695_, _066696_, _066697_);
  or g_124029_(_066694_, _066697_, _066698_);
  xor g_124030_(out[140], out[572], _066699_);
  or g_124031_(_066674_, _066699_, _066700_);
  or g_124032_(_066673_, _066685_, _066701_);
  or g_124033_(_066700_, _066701_, _066702_);
  or g_124034_(_066677_, _066683_, _066704_);
  or g_124035_(_066686_, _066704_, _066705_);
  or g_124036_(_066702_, _066705_, _066706_);
  or g_124037_(_066698_, _066706_, _066707_);
  or g_124038_(_066690_, _066707_, _066708_);
  xor g_124039_(out[113], out[561], _066709_);
  and g_124040_(out[123], _049554_, _066710_);
  xor g_124041_(out[121], out[569], _066711_);
  xor g_124042_(out[112], out[560], _066712_);
  xor g_124043_(out[126], out[574], _066713_);
  xor g_124044_(out[116], out[564], _066715_);
  or g_124045_(_066713_, _066715_, _066716_);
  xor g_124046_(out[125], out[573], _066717_);
  xor g_124047_(out[115], out[563], _066718_);
  and g_124048_(_098151_, out[571], _066719_);
  xor g_124049_(out[118], out[566], _066720_);
  xor g_124050_(out[122], out[570], _066721_);
  xor g_124051_(out[117], out[565], _066722_);
  xor g_124052_(out[127], out[575], _066723_);
  xor g_124053_(out[120], out[568], _066724_);
  or g_124054_(_066717_, _066724_, _066726_);
  xor g_124055_(out[114], out[562], _066727_);
  or g_124056_(_066721_, _066727_, _066728_);
  or g_124057_(_066726_, _066728_, _066729_);
  or g_124058_(_066711_, _066718_, _066730_);
  or g_124059_(_066722_, _066730_, _066731_);
  or g_124060_(_066729_, _066731_, _066732_);
  or g_124061_(_066716_, _066732_, _066733_);
  xor g_124062_(out[124], out[572], _066734_);
  or g_124063_(_066719_, _066734_, _066735_);
  xor g_124064_(out[119], out[567], _066737_);
  or g_124065_(_066720_, _066737_, _066738_);
  or g_124066_(_066735_, _066738_, _066739_);
  or g_124067_(_066709_, _066710_, _066740_);
  or g_124068_(_066723_, _066740_, _066741_);
  or g_124069_(_066739_, _066741_, _066742_);
  or g_124070_(_066712_, _066742_, _066743_);
  or g_124071_(_066733_, _066743_, _066744_);
  xor g_124072_(out[103], out[567], _066745_);
  and g_124073_(_098140_, out[571], _066746_);
  xor g_124074_(out[110], out[574], _066748_);
  xor g_124075_(out[104], out[568], _066749_);
  xor g_124076_(out[97], out[561], _066750_);
  xor g_124077_(out[109], out[573], _066751_);
  xor g_124078_(out[105], out[569], _066752_);
  xor g_124079_(out[100], out[564], _066753_);
  xor g_124080_(out[98], out[562], _066754_);
  and g_124081_(out[107], _049554_, _066755_);
  xor g_124082_(out[99], out[563], _066756_);
  xor g_124083_(out[102], out[566], _066757_);
  xor g_124084_(out[111], out[575], _066759_);
  xor g_124085_(out[106], out[570], _066760_);
  xor g_124086_(out[101], out[565], _066761_);
  xor g_124087_(out[96], out[560], _066762_);
  or g_124088_(_066748_, _066753_, _066763_);
  or g_124089_(_066749_, _066751_, _066764_);
  or g_124090_(_066754_, _066760_, _066765_);
  or g_124091_(_066764_, _066765_, _066766_);
  or g_124092_(_066752_, _066756_, _066767_);
  or g_124093_(_066761_, _066762_, _066768_);
  or g_124094_(_066767_, _066768_, _066770_);
  or g_124095_(_066766_, _066770_, _066771_);
  xor g_124096_(out[108], out[572], _066772_);
  or g_124097_(_066746_, _066772_, _066773_);
  or g_124098_(_066745_, _066757_, _066774_);
  or g_124099_(_066773_, _066774_, _066775_);
  or g_124100_(_066750_, _066755_, _066776_);
  or g_124101_(_066759_, _066776_, _066777_);
  or g_124102_(_066775_, _066777_, _066778_);
  or g_124103_(_066771_, _066778_, _066779_);
  or g_124104_(_066763_, _066779_, _066781_);
  xor g_124105_(out[81], out[561], _066782_);
  and g_124106_(out[91], _049554_, _066783_);
  xor g_124107_(out[89], out[569], _066784_);
  xor g_124108_(out[80], out[560], _066785_);
  xor g_124109_(out[94], out[574], _066786_);
  xor g_124110_(out[84], out[564], _066787_);
  or g_124111_(_066786_, _066787_, _066788_);
  xor g_124112_(out[93], out[573], _066789_);
  xor g_124113_(out[83], out[563], _066790_);
  and g_124114_(_098129_, out[571], _066792_);
  xor g_124115_(out[86], out[566], _066793_);
  xor g_124116_(out[90], out[570], _066794_);
  xor g_124117_(out[85], out[565], _066795_);
  xor g_124118_(out[95], out[575], _066796_);
  xor g_124119_(out[88], out[568], _066797_);
  or g_124120_(_066789_, _066797_, _066798_);
  xor g_124121_(out[82], out[562], _066799_);
  or g_124122_(_066794_, _066799_, _066800_);
  or g_124123_(_066798_, _066800_, _066801_);
  or g_124124_(_066784_, _066790_, _066803_);
  or g_124125_(_066795_, _066803_, _066804_);
  or g_124126_(_066801_, _066804_, _066805_);
  or g_124127_(_066788_, _066805_, _066806_);
  xor g_124128_(out[92], out[572], _066807_);
  or g_124129_(_066792_, _066807_, _066808_);
  xor g_124130_(out[87], out[567], _066809_);
  or g_124131_(_066793_, _066809_, _066810_);
  or g_124132_(_066808_, _066810_, _066811_);
  or g_124133_(_066782_, _066783_, _066812_);
  or g_124134_(_066796_, _066812_, _066814_);
  or g_124135_(_066811_, _066814_, _066815_);
  or g_124136_(_066785_, _066815_, _066816_);
  or g_124137_(_066806_, _066816_, _066817_);
  xor g_124138_(out[71], out[567], _066818_);
  and g_124139_(_098118_, out[571], _066819_);
  xor g_124140_(out[78], out[574], _066820_);
  xor g_124141_(out[72], out[568], _066821_);
  xor g_124142_(out[65], out[561], _066822_);
  xor g_124143_(out[77], out[573], _066823_);
  xor g_124144_(out[73], out[569], _066825_);
  xor g_124145_(out[68], out[564], _066826_);
  xor g_124146_(out[66], out[562], _066827_);
  and g_124147_(out[75], _049554_, _066828_);
  xor g_124148_(out[67], out[563], _066829_);
  xor g_124149_(out[70], out[566], _066830_);
  xor g_124150_(out[79], out[575], _066831_);
  xor g_124151_(out[74], out[570], _066832_);
  xor g_124152_(out[69], out[565], _066833_);
  xor g_124153_(out[64], out[560], _066834_);
  or g_124154_(_066820_, _066826_, _066836_);
  or g_124155_(_066821_, _066823_, _066837_);
  or g_124156_(_066827_, _066832_, _066838_);
  or g_124157_(_066837_, _066838_, _066839_);
  or g_124158_(_066825_, _066829_, _066840_);
  or g_124159_(_066833_, _066834_, _066841_);
  or g_124160_(_066840_, _066841_, _066842_);
  or g_124161_(_066839_, _066842_, _066843_);
  xor g_124162_(out[76], out[572], _066844_);
  or g_124163_(_066819_, _066844_, _066845_);
  or g_124164_(_066818_, _066830_, _066847_);
  or g_124165_(_066845_, _066847_, _066848_);
  or g_124166_(_066822_, _066828_, _066849_);
  or g_124167_(_066831_, _066849_, _066850_);
  or g_124168_(_066848_, _066850_, _066851_);
  or g_124169_(_066843_, _066851_, _066852_);
  or g_124170_(_066836_, _066852_, _066853_);
  xor g_124171_(out[49], out[561], _066854_);
  and g_124172_(out[59], _049554_, _066855_);
  xor g_124173_(out[62], out[574], _066856_);
  xor g_124174_(out[51], out[563], _066858_);
  xor g_124175_(out[52], out[564], _066859_);
  xor g_124176_(out[50], out[562], _066860_);
  xor g_124177_(out[57], out[569], _066861_);
  xor g_124178_(out[48], out[560], _066862_);
  and g_124179_(_098107_, out[571], _066863_);
  xor g_124180_(out[54], out[566], _066864_);
  xor g_124181_(out[58], out[570], _066865_);
  xor g_124182_(out[53], out[565], _066866_);
  xor g_124183_(out[63], out[575], _066867_);
  xor g_124184_(out[61], out[573], _066869_);
  xor g_124185_(out[56], out[568], _066870_);
  or g_124186_(_066856_, _066859_, _066871_);
  or g_124187_(_066869_, _066870_, _066872_);
  or g_124188_(_066860_, _066865_, _066873_);
  or g_124189_(_066872_, _066873_, _066874_);
  or g_124190_(_066858_, _066861_, _066875_);
  or g_124191_(_066862_, _066866_, _066876_);
  or g_124192_(_066875_, _066876_, _066877_);
  or g_124193_(_066874_, _066877_, _066878_);
  xor g_124194_(out[60], out[572], _066880_);
  or g_124195_(_066863_, _066880_, _066881_);
  xor g_124196_(out[55], out[567], _066882_);
  or g_124197_(_066864_, _066882_, _066883_);
  or g_124198_(_066881_, _066883_, _066884_);
  or g_124199_(_066854_, _066855_, _066885_);
  or g_124200_(_066867_, _066885_, _066886_);
  or g_124201_(_066884_, _066886_, _066887_);
  or g_124202_(_066878_, _066887_, _066888_);
  or g_124203_(_066871_, _066888_, _066889_);
  xor g_124204_(out[39], out[567], _066891_);
  and g_124205_(_098096_, out[571], _066892_);
  xor g_124206_(out[46], out[574], _066893_);
  xor g_124207_(out[40], out[568], _066894_);
  xor g_124208_(out[33], out[561], _066895_);
  xor g_124209_(out[45], out[573], _066896_);
  xor g_124210_(out[41], out[569], _066897_);
  xor g_124211_(out[36], out[564], _066898_);
  xor g_124212_(out[34], out[562], _066899_);
  and g_124213_(out[43], _049554_, _066900_);
  xor g_124214_(out[35], out[563], _066902_);
  xor g_124215_(out[38], out[566], _066903_);
  xor g_124216_(out[47], out[575], _066904_);
  xor g_124217_(out[42], out[570], _066905_);
  xor g_124218_(out[37], out[565], _066906_);
  xor g_124219_(out[32], out[560], _066907_);
  or g_124220_(_066893_, _066898_, _066908_);
  or g_124221_(_066894_, _066896_, _066909_);
  or g_124222_(_066899_, _066905_, _066910_);
  or g_124223_(_066909_, _066910_, _066911_);
  or g_124224_(_066897_, _066902_, _066913_);
  or g_124225_(_066906_, _066907_, _066914_);
  or g_124226_(_066913_, _066914_, _066915_);
  or g_124227_(_066911_, _066915_, _066916_);
  xor g_124228_(out[44], out[572], _066917_);
  or g_124229_(_066892_, _066917_, _066918_);
  or g_124230_(_066891_, _066903_, _066919_);
  or g_124231_(_066918_, _066919_, _066920_);
  or g_124232_(_066895_, _066900_, _066921_);
  or g_124233_(_066904_, _066921_, _066922_);
  or g_124234_(_066920_, _066922_, _066924_);
  or g_124235_(_066916_, _066924_, _066925_);
  or g_124236_(_066908_, _066925_, _066926_);
  xor g_124237_(out[18], out[562], _066927_);
  xor g_124238_(out[16], out[560], _066928_);
  xor g_124239_(out[25], out[569], _066929_);
  xor g_124240_(out[24], out[568], _066930_);
  xor g_124241_(out[21], out[565], _066931_);
  xor g_124242_(out[30], out[574], _066932_);
  xor g_124243_(out[29], out[573], _066933_);
  xor g_124244_(out[31], out[575], _066935_);
  xor g_124245_(out[26], out[570], _066936_);
  xor g_124246_(out[22], out[566], _066937_);
  xor g_124247_(out[19], out[563], _066938_);
  and g_124248_(_098063_, out[571], _066939_);
  and g_124249_(out[27], _049554_, _066940_);
  xor g_124250_(out[20], out[564], _066941_);
  xor g_124251_(out[17], out[561], _066942_);
  or g_124252_(_066932_, _066941_, _066943_);
  or g_124253_(_066930_, _066933_, _066944_);
  or g_124254_(_066927_, _066936_, _066946_);
  or g_124255_(_066944_, _066946_, _066947_);
  or g_124256_(_066929_, _066938_, _066948_);
  or g_124257_(_066928_, _066931_, _066949_);
  or g_124258_(_066948_, _066949_, _066950_);
  or g_124259_(_066947_, _066950_, _066951_);
  xor g_124260_(out[28], out[572], _066952_);
  or g_124261_(_066939_, _066952_, _066953_);
  xor g_124262_(out[23], out[567], _066954_);
  or g_124263_(_066937_, _066954_, _066955_);
  or g_124264_(_066953_, _066955_, _066957_);
  or g_124265_(_066940_, _066942_, _066958_);
  or g_124266_(_066935_, _066958_, _066959_);
  or g_124267_(_066957_, _066959_, _066960_);
  or g_124268_(_066951_, _066960_, _066961_);
  or g_124269_(_066943_, _066961_, _066962_);
  not g_124270_(_066962_, _066963_);
  xor g_124271_(out[12], out[572], _066964_);
  and g_124272_(_098041_, out[571], _066965_);
  xor g_124273_(out[8], out[568], _066966_);
  xor g_124274_(out[6], out[566], _066968_);
  xor g_124275_(out[13], out[573], _066969_);
  xor g_124276_(out[14], out[574], _066970_);
  xor g_124277_(out[2], out[562], _066971_);
  xor g_124278_(out[9], out[569], _066972_);
  xor g_124279_(out[5], out[565], _066973_);
  xor g_124280_(out[1], out[561], _066974_);
  and g_124281_(out[11], _049554_, _066975_);
  or g_124282_(_066966_, _066969_, _066976_);
  xor g_124283_(out[15], out[575], _066977_);
  xor g_124284_(out[10], out[570], _066979_);
  xor g_124285_(out[4], out[564], _066980_);
  xor g_124286_(out[3], out[563], _066981_);
  xor g_124287_(out[0], out[560], _066982_);
  or g_124288_(_066971_, _066979_, _066983_);
  or g_124289_(_066976_, _066983_, _066984_);
  or g_124290_(_066972_, _066981_, _066985_);
  or g_124291_(_066973_, _066985_, _066986_);
  or g_124292_(_066984_, _066986_, _066987_);
  or g_124293_(_066970_, _066980_, _066988_);
  or g_124294_(_066987_, _066988_, _066990_);
  or g_124295_(_066964_, _066965_, _066991_);
  xor g_124296_(out[7], out[567], _066992_);
  or g_124297_(_066968_, _066992_, _066993_);
  or g_124298_(_066991_, _066993_, _066994_);
  or g_124299_(_066974_, _066975_, _066995_);
  or g_124300_(_066977_, _066995_, _066996_);
  or g_124301_(_066994_, _066996_, _066997_);
  or g_124302_(_066982_, _066997_, _066998_);
  or g_124303_(_066990_, _066998_, _066999_);
  not g_124304_(_066999_, _067001_);
  xor g_124305_(out[471], out[551], _067002_);
  and g_124306_(_049499_, out[555], _067003_);
  xor g_124307_(out[478], out[558], _067004_);
  xor g_124308_(out[472], out[552], _067005_);
  xor g_124309_(out[465], out[545], _067006_);
  xor g_124310_(out[477], out[557], _067007_);
  xor g_124311_(out[473], out[553], _067008_);
  xor g_124312_(out[468], out[548], _067009_);
  xor g_124313_(out[466], out[546], _067010_);
  and g_124314_(out[475], _049543_, _067012_);
  xor g_124315_(out[467], out[547], _067013_);
  xor g_124316_(out[470], out[550], _067014_);
  xor g_124317_(out[479], out[559], _067015_);
  xor g_124318_(out[474], out[554], _067016_);
  xor g_124319_(out[469], out[549], _067017_);
  xor g_124320_(out[464], out[544], _067018_);
  or g_124321_(_067004_, _067009_, _067019_);
  or g_124322_(_067005_, _067007_, _067020_);
  or g_124323_(_067010_, _067016_, _067021_);
  or g_124324_(_067020_, _067021_, _067023_);
  or g_124325_(_067008_, _067013_, _067024_);
  or g_124326_(_067017_, _067018_, _067025_);
  or g_124327_(_067024_, _067025_, _067026_);
  or g_124328_(_067023_, _067026_, _067027_);
  xor g_124329_(out[476], out[556], _067028_);
  or g_124330_(_067003_, _067028_, _067029_);
  or g_124331_(_067002_, _067014_, _067030_);
  or g_124332_(_067029_, _067030_, _067031_);
  or g_124333_(_067006_, _067012_, _067032_);
  or g_124334_(_067015_, _067032_, _067034_);
  or g_124335_(_067031_, _067034_, _067035_);
  or g_124336_(_067027_, _067035_, _067036_);
  or g_124337_(_067019_, _067036_, _067037_);
  not g_124338_(_067037_, _067038_);
  and g_124339_(out[459], _049543_, _067039_);
  xor g_124340_(out[452], out[548], _067040_);
  xor g_124341_(out[462], out[558], _067041_);
  or g_124342_(_067040_, _067041_, _067042_);
  xor g_124343_(out[461], out[557], _067043_);
  xor g_124344_(out[451], out[547], _067045_);
  xor g_124345_(out[448], out[544], _067046_);
  and g_124346_(_049477_, out[555], _067047_);
  xor g_124347_(out[458], out[554], _067048_);
  xor g_124348_(out[463], out[559], _067049_);
  xor g_124349_(out[454], out[550], _067050_);
  xor g_124350_(out[453], out[549], _067051_);
  xor g_124351_(out[456], out[552], _067052_);
  or g_124352_(_067043_, _067052_, _067053_);
  xor g_124353_(out[450], out[546], _067054_);
  xor g_124354_(out[457], out[553], _067056_);
  xor g_124355_(out[449], out[545], _067057_);
  or g_124356_(_067048_, _067054_, _067058_);
  or g_124357_(_067053_, _067058_, _067059_);
  or g_124358_(_067045_, _067056_, _067060_);
  or g_124359_(_067051_, _067060_, _067061_);
  or g_124360_(_067059_, _067061_, _067062_);
  or g_124361_(_067042_, _067062_, _067063_);
  xor g_124362_(out[460], out[556], _067064_);
  or g_124363_(_067047_, _067064_, _067065_);
  xor g_124364_(out[455], out[551], _067067_);
  or g_124365_(_067050_, _067067_, _067068_);
  or g_124366_(_067065_, _067068_, _067069_);
  or g_124367_(_067039_, _067057_, _067070_);
  or g_124368_(_067049_, _067070_, _067071_);
  or g_124369_(_067069_, _067071_, _067072_);
  or g_124370_(_067046_, _067072_, _067073_);
  or g_124371_(_067063_, _067073_, _067074_);
  not g_124372_(_067074_, _067075_);
  xor g_124373_(out[439], out[551], _067076_);
  and g_124374_(_049466_, out[555], _067078_);
  xor g_124375_(out[446], out[558], _067079_);
  xor g_124376_(out[440], out[552], _067080_);
  xor g_124377_(out[433], out[545], _067081_);
  xor g_124378_(out[445], out[557], _067082_);
  xor g_124379_(out[441], out[553], _067083_);
  xor g_124380_(out[436], out[548], _067084_);
  xor g_124381_(out[434], out[546], _067085_);
  and g_124382_(out[443], _049543_, _067086_);
  xor g_124383_(out[435], out[547], _067087_);
  xor g_124384_(out[438], out[550], _067089_);
  xor g_124385_(out[447], out[559], _067090_);
  xor g_124386_(out[442], out[554], _067091_);
  xor g_124387_(out[437], out[549], _067092_);
  xor g_124388_(out[432], out[544], _067093_);
  or g_124389_(_067079_, _067084_, _067094_);
  or g_124390_(_067080_, _067082_, _067095_);
  or g_124391_(_067085_, _067091_, _067096_);
  or g_124392_(_067095_, _067096_, _067097_);
  or g_124393_(_067083_, _067087_, _067098_);
  or g_124394_(_067092_, _067093_, _067100_);
  or g_124395_(_067098_, _067100_, _067101_);
  or g_124396_(_067097_, _067101_, _067102_);
  xor g_124397_(out[444], out[556], _067103_);
  or g_124398_(_067078_, _067103_, _067104_);
  or g_124399_(_067076_, _067089_, _067105_);
  or g_124400_(_067104_, _067105_, _067106_);
  or g_124401_(_067081_, _067086_, _067107_);
  or g_124402_(_067090_, _067107_, _067108_);
  or g_124403_(_067106_, _067108_, _067109_);
  or g_124404_(_067102_, _067109_, _067111_);
  or g_124405_(_067094_, _067111_, _067112_);
  xor g_124406_(out[417], out[545], _067113_);
  and g_124407_(out[427], _049543_, _067114_);
  xor g_124408_(out[425], out[553], _067115_);
  xor g_124409_(out[416], out[544], _067116_);
  xor g_124410_(out[430], out[558], _067117_);
  xor g_124411_(out[420], out[548], _067118_);
  or g_124412_(_067117_, _067118_, _067119_);
  xor g_124413_(out[429], out[557], _067120_);
  xor g_124414_(out[419], out[547], _067122_);
  and g_124415_(_049455_, out[555], _067123_);
  xor g_124416_(out[422], out[550], _067124_);
  xor g_124417_(out[426], out[554], _067125_);
  xor g_124418_(out[421], out[549], _067126_);
  xor g_124419_(out[431], out[559], _067127_);
  xor g_124420_(out[424], out[552], _067128_);
  or g_124421_(_067120_, _067128_, _067129_);
  xor g_124422_(out[418], out[546], _067130_);
  or g_124423_(_067125_, _067130_, _067131_);
  or g_124424_(_067129_, _067131_, _067133_);
  or g_124425_(_067115_, _067122_, _067134_);
  or g_124426_(_067126_, _067134_, _067135_);
  or g_124427_(_067133_, _067135_, _067136_);
  or g_124428_(_067119_, _067136_, _067137_);
  xor g_124429_(out[428], out[556], _067138_);
  or g_124430_(_067123_, _067138_, _067139_);
  xor g_124431_(out[423], out[551], _067140_);
  or g_124432_(_067124_, _067140_, _067141_);
  or g_124433_(_067139_, _067141_, _067142_);
  or g_124434_(_067113_, _067114_, _067144_);
  or g_124435_(_067127_, _067144_, _067145_);
  or g_124436_(_067142_, _067145_, _067146_);
  or g_124437_(_067116_, _067146_, _067147_);
  or g_124438_(_067137_, _067147_, _067148_);
  xor g_124439_(out[407], out[551], _067149_);
  and g_124440_(_049444_, out[555], _067150_);
  xor g_124441_(out[414], out[558], _067151_);
  xor g_124442_(out[408], out[552], _067152_);
  xor g_124443_(out[401], out[545], _067153_);
  xor g_124444_(out[413], out[557], _067155_);
  xor g_124445_(out[409], out[553], _067156_);
  xor g_124446_(out[404], out[548], _067157_);
  xor g_124447_(out[402], out[546], _067158_);
  and g_124448_(out[411], _049543_, _067159_);
  xor g_124449_(out[403], out[547], _067160_);
  xor g_124450_(out[406], out[550], _067161_);
  xor g_124451_(out[415], out[559], _067162_);
  xor g_124452_(out[410], out[554], _067163_);
  xor g_124453_(out[405], out[549], _067164_);
  xor g_124454_(out[400], out[544], _067166_);
  or g_124455_(_067151_, _067157_, _067167_);
  or g_124456_(_067152_, _067155_, _067168_);
  or g_124457_(_067158_, _067163_, _067169_);
  or g_124458_(_067168_, _067169_, _067170_);
  or g_124459_(_067156_, _067160_, _067171_);
  or g_124460_(_067164_, _067166_, _067172_);
  or g_124461_(_067171_, _067172_, _067173_);
  or g_124462_(_067170_, _067173_, _067174_);
  xor g_124463_(out[412], out[556], _067175_);
  or g_124464_(_067150_, _067175_, _067177_);
  or g_124465_(_067149_, _067161_, _067178_);
  or g_124466_(_067177_, _067178_, _067179_);
  or g_124467_(_067153_, _067159_, _067180_);
  or g_124468_(_067162_, _067180_, _067181_);
  or g_124469_(_067179_, _067181_, _067182_);
  or g_124470_(_067174_, _067182_, _067183_);
  or g_124471_(_067167_, _067183_, _067184_);
  xor g_124472_(out[385], out[545], _067185_);
  and g_124473_(_049433_, out[555], _067186_);
  and g_124474_(out[395], _049543_, _067188_);
  xor g_124475_(out[393], out[553], _067189_);
  xor g_124476_(out[384], out[544], _067190_);
  xor g_124477_(out[398], out[558], _067191_);
  xor g_124478_(out[388], out[548], _067192_);
  or g_124479_(_067191_, _067192_, _067193_);
  xor g_124480_(out[397], out[557], _067194_);
  xor g_124481_(out[387], out[547], _067195_);
  xor g_124482_(out[396], out[556], _067196_);
  xor g_124483_(out[390], out[550], _067197_);
  xor g_124484_(out[394], out[554], _067199_);
  xor g_124485_(out[389], out[549], _067200_);
  xor g_124486_(out[399], out[559], _067201_);
  xor g_124487_(out[392], out[552], _067202_);
  or g_124488_(_067194_, _067202_, _067203_);
  xor g_124489_(out[386], out[546], _067204_);
  or g_124490_(_067199_, _067204_, _067205_);
  or g_124491_(_067203_, _067205_, _067206_);
  or g_124492_(_067189_, _067195_, _067207_);
  or g_124493_(_067200_, _067207_, _067208_);
  or g_124494_(_067206_, _067208_, _067210_);
  or g_124495_(_067193_, _067210_, _067211_);
  or g_124496_(_067186_, _067196_, _067212_);
  xor g_124497_(out[391], out[551], _067213_);
  or g_124498_(_067197_, _067213_, _067214_);
  or g_124499_(_067212_, _067214_, _067215_);
  or g_124500_(_067185_, _067188_, _067216_);
  or g_124501_(_067201_, _067216_, _067217_);
  or g_124502_(_067215_, _067217_, _067218_);
  or g_124503_(_067190_, _067218_, _067219_);
  or g_124504_(_067211_, _067219_, _067221_);
  not g_124505_(_067221_, _067222_);
  xor g_124506_(out[375], out[551], _067223_);
  and g_124507_(_049422_, out[555], _067224_);
  xor g_124508_(out[382], out[558], _067225_);
  xor g_124509_(out[376], out[552], _067226_);
  xor g_124510_(out[369], out[545], _067227_);
  xor g_124511_(out[381], out[557], _067228_);
  xor g_124512_(out[377], out[553], _067229_);
  xor g_124513_(out[372], out[548], _067230_);
  xor g_124514_(out[370], out[546], _067232_);
  and g_124515_(out[379], _049543_, _067233_);
  xor g_124516_(out[371], out[547], _067234_);
  xor g_124517_(out[374], out[550], _067235_);
  xor g_124518_(out[383], out[559], _067236_);
  xor g_124519_(out[378], out[554], _067237_);
  xor g_124520_(out[373], out[549], _067238_);
  xor g_124521_(out[368], out[544], _067239_);
  or g_124522_(_067225_, _067230_, _067240_);
  or g_124523_(_067226_, _067228_, _067241_);
  or g_124524_(_067232_, _067237_, _067243_);
  or g_124525_(_067241_, _067243_, _067244_);
  or g_124526_(_067229_, _067234_, _067245_);
  or g_124527_(_067238_, _067239_, _067246_);
  or g_124528_(_067245_, _067246_, _067247_);
  or g_124529_(_067244_, _067247_, _067248_);
  xor g_124530_(out[380], out[556], _067249_);
  or g_124531_(_067224_, _067249_, _067250_);
  or g_124532_(_067223_, _067235_, _067251_);
  or g_124533_(_067250_, _067251_, _067252_);
  or g_124534_(_067227_, _067233_, _067254_);
  or g_124535_(_067236_, _067254_, _067255_);
  or g_124536_(_067252_, _067255_, _067256_);
  or g_124537_(_067248_, _067256_, _067257_);
  or g_124538_(_067240_, _067257_, _067258_);
  not g_124539_(_067258_, _067259_);
  xor g_124540_(out[353], out[545], _067260_);
  and g_124541_(out[363], _049543_, _067261_);
  xor g_124542_(out[361], out[553], _067262_);
  xor g_124543_(out[352], out[544], _067263_);
  xor g_124544_(out[366], out[558], _067265_);
  xor g_124545_(out[356], out[548], _067266_);
  or g_124546_(_067265_, _067266_, _067267_);
  xor g_124547_(out[365], out[557], _067268_);
  xor g_124548_(out[355], out[547], _067269_);
  and g_124549_(_049411_, out[555], _067270_);
  xor g_124550_(out[358], out[550], _067271_);
  xor g_124551_(out[362], out[554], _067272_);
  xor g_124552_(out[357], out[549], _067273_);
  xor g_124553_(out[367], out[559], _067274_);
  xor g_124554_(out[360], out[552], _067276_);
  or g_124555_(_067268_, _067276_, _067277_);
  xor g_124556_(out[354], out[546], _067278_);
  or g_124557_(_067272_, _067278_, _067279_);
  or g_124558_(_067277_, _067279_, _067280_);
  or g_124559_(_067262_, _067269_, _067281_);
  or g_124560_(_067273_, _067281_, _067282_);
  or g_124561_(_067280_, _067282_, _067283_);
  or g_124562_(_067267_, _067283_, _067284_);
  xor g_124563_(out[364], out[556], _067285_);
  or g_124564_(_067270_, _067285_, _067287_);
  xor g_124565_(out[359], out[551], _067288_);
  or g_124566_(_067271_, _067288_, _067289_);
  or g_124567_(_067287_, _067289_, _067290_);
  or g_124568_(_067260_, _067261_, _067291_);
  or g_124569_(_067274_, _067291_, _067292_);
  or g_124570_(_067290_, _067292_, _067293_);
  or g_124571_(_067263_, _067293_, _067294_);
  or g_124572_(_067284_, _067294_, _067295_);
  xor g_124573_(out[343], out[551], _067296_);
  and g_124574_(_049400_, out[555], _067298_);
  xor g_124575_(out[350], out[558], _067299_);
  xor g_124576_(out[344], out[552], _067300_);
  xor g_124577_(out[337], out[545], _067301_);
  xor g_124578_(out[349], out[557], _067302_);
  xor g_124579_(out[345], out[553], _067303_);
  xor g_124580_(out[340], out[548], _067304_);
  xor g_124581_(out[338], out[546], _067305_);
  and g_124582_(out[347], _049543_, _067306_);
  xor g_124583_(out[339], out[547], _067307_);
  xor g_124584_(out[342], out[550], _067309_);
  xor g_124585_(out[351], out[559], _067310_);
  xor g_124586_(out[346], out[554], _067311_);
  xor g_124587_(out[341], out[549], _067312_);
  xor g_124588_(out[336], out[544], _067313_);
  or g_124589_(_067299_, _067304_, _067314_);
  or g_124590_(_067300_, _067302_, _067315_);
  or g_124591_(_067305_, _067311_, _067316_);
  or g_124592_(_067315_, _067316_, _067317_);
  or g_124593_(_067303_, _067307_, _067318_);
  or g_124594_(_067312_, _067313_, _067320_);
  or g_124595_(_067318_, _067320_, _067321_);
  or g_124596_(_067317_, _067321_, _067322_);
  xor g_124597_(out[348], out[556], _067323_);
  or g_124598_(_067298_, _067323_, _067324_);
  or g_124599_(_067296_, _067309_, _067325_);
  or g_124600_(_067324_, _067325_, _067326_);
  or g_124601_(_067301_, _067306_, _067327_);
  or g_124602_(_067310_, _067327_, _067328_);
  or g_124603_(_067326_, _067328_, _067329_);
  or g_124604_(_067322_, _067329_, _067331_);
  or g_124605_(_067314_, _067331_, _067332_);
  xor g_124606_(out[321], out[545], _067333_);
  and g_124607_(out[331], _049543_, _067334_);
  xor g_124608_(out[329], out[553], _067335_);
  xor g_124609_(out[320], out[544], _067336_);
  xor g_124610_(out[334], out[558], _067337_);
  xor g_124611_(out[324], out[548], _067338_);
  or g_124612_(_067337_, _067338_, _067339_);
  xor g_124613_(out[333], out[557], _067340_);
  xor g_124614_(out[323], out[547], _067342_);
  and g_124615_(_098294_, out[555], _067343_);
  xor g_124616_(out[326], out[550], _067344_);
  xor g_124617_(out[330], out[554], _067345_);
  xor g_124618_(out[325], out[549], _067346_);
  xor g_124619_(out[335], out[559], _067347_);
  xor g_124620_(out[328], out[552], _067348_);
  or g_124621_(_067340_, _067348_, _067349_);
  xor g_124622_(out[322], out[546], _067350_);
  or g_124623_(_067345_, _067350_, _067351_);
  or g_124624_(_067349_, _067351_, _067353_);
  or g_124625_(_067335_, _067342_, _067354_);
  or g_124626_(_067346_, _067354_, _067355_);
  or g_124627_(_067353_, _067355_, _067356_);
  or g_124628_(_067339_, _067356_, _067357_);
  xor g_124629_(out[332], out[556], _067358_);
  or g_124630_(_067343_, _067358_, _067359_);
  xor g_124631_(out[327], out[551], _067360_);
  or g_124632_(_067344_, _067360_, _067361_);
  or g_124633_(_067359_, _067361_, _067362_);
  or g_124634_(_067333_, _067334_, _067364_);
  or g_124635_(_067347_, _067364_, _067365_);
  or g_124636_(_067362_, _067365_, _067366_);
  or g_124637_(_067336_, _067366_, _067367_);
  or g_124638_(_067357_, _067367_, _067368_);
  xor g_124639_(out[311], out[551], _067369_);
  and g_124640_(_098283_, out[555], _067370_);
  xor g_124641_(out[318], out[558], _067371_);
  xor g_124642_(out[312], out[552], _067372_);
  xor g_124643_(out[305], out[545], _067373_);
  xor g_124644_(out[317], out[557], _067375_);
  xor g_124645_(out[313], out[553], _067376_);
  xor g_124646_(out[308], out[548], _067377_);
  xor g_124647_(out[306], out[546], _067378_);
  and g_124648_(out[315], _049543_, _067379_);
  xor g_124649_(out[307], out[547], _067380_);
  xor g_124650_(out[310], out[550], _067381_);
  xor g_124651_(out[319], out[559], _067382_);
  xor g_124652_(out[314], out[554], _067383_);
  xor g_124653_(out[309], out[549], _067384_);
  xor g_124654_(out[304], out[544], _067386_);
  or g_124655_(_067371_, _067377_, _067387_);
  or g_124656_(_067372_, _067375_, _067388_);
  or g_124657_(_067378_, _067383_, _067389_);
  or g_124658_(_067388_, _067389_, _067390_);
  or g_124659_(_067376_, _067380_, _067391_);
  or g_124660_(_067384_, _067386_, _067392_);
  or g_124661_(_067391_, _067392_, _067393_);
  or g_124662_(_067390_, _067393_, _067394_);
  xor g_124663_(out[316], out[556], _067395_);
  or g_124664_(_067370_, _067395_, _067397_);
  or g_124665_(_067369_, _067381_, _067398_);
  or g_124666_(_067397_, _067398_, _067399_);
  or g_124667_(_067373_, _067379_, _067400_);
  or g_124668_(_067382_, _067400_, _067401_);
  or g_124669_(_067399_, _067401_, _067402_);
  or g_124670_(_067394_, _067402_, _067403_);
  or g_124671_(_067387_, _067403_, _067404_);
  and g_124672_(out[299], _049543_, _067405_);
  xor g_124673_(out[292], out[548], _067406_);
  xor g_124674_(out[290], out[546], _067408_);
  xor g_124675_(out[297], out[553], _067409_);
  xor g_124676_(out[288], out[544], _067410_);
  xor g_124677_(out[291], out[547], _067411_);
  and g_124678_(_098272_, out[555], _067412_);
  xor g_124679_(out[298], out[554], _067413_);
  xor g_124680_(out[303], out[559], _067414_);
  xor g_124681_(out[294], out[550], _067415_);
  xor g_124682_(out[293], out[549], _067416_);
  xor g_124683_(out[301], out[557], _067417_);
  xor g_124684_(out[302], out[558], _067419_);
  xor g_124685_(out[296], out[552], _067420_);
  xor g_124686_(out[289], out[545], _067421_);
  or g_124687_(_067406_, _067419_, _067422_);
  or g_124688_(_067417_, _067420_, _067423_);
  or g_124689_(_067408_, _067413_, _067424_);
  or g_124690_(_067423_, _067424_, _067425_);
  or g_124691_(_067409_, _067411_, _067426_);
  or g_124692_(_067410_, _067416_, _067427_);
  or g_124693_(_067426_, _067427_, _067428_);
  or g_124694_(_067425_, _067428_, _067430_);
  xor g_124695_(out[300], out[556], _067431_);
  or g_124696_(_067412_, _067431_, _067432_);
  xor g_124697_(out[295], out[551], _067433_);
  or g_124698_(_067415_, _067433_, _067434_);
  or g_124699_(_067432_, _067434_, _067435_);
  or g_124700_(_067405_, _067421_, _067436_);
  or g_124701_(_067414_, _067436_, _067437_);
  or g_124702_(_067435_, _067437_, _067438_);
  or g_124703_(_067430_, _067438_, _067439_);
  or g_124704_(_067422_, _067439_, _067441_);
  xor g_124705_(out[279], out[551], _067442_);
  and g_124706_(_098261_, out[555], _067443_);
  xor g_124707_(out[286], out[558], _067444_);
  xor g_124708_(out[280], out[552], _067445_);
  xor g_124709_(out[273], out[545], _067446_);
  xor g_124710_(out[285], out[557], _067447_);
  xor g_124711_(out[281], out[553], _067448_);
  xor g_124712_(out[276], out[548], _067449_);
  xor g_124713_(out[274], out[546], _067450_);
  and g_124714_(out[283], _049543_, _067452_);
  xor g_124715_(out[275], out[547], _067453_);
  xor g_124716_(out[278], out[550], _067454_);
  xor g_124717_(out[287], out[559], _067455_);
  xor g_124718_(out[282], out[554], _067456_);
  xor g_124719_(out[277], out[549], _067457_);
  xor g_124720_(out[272], out[544], _067458_);
  or g_124721_(_067444_, _067449_, _067459_);
  or g_124722_(_067445_, _067447_, _067460_);
  or g_124723_(_067450_, _067456_, _067461_);
  or g_124724_(_067460_, _067461_, _067463_);
  or g_124725_(_067448_, _067453_, _067464_);
  or g_124726_(_067457_, _067458_, _067465_);
  or g_124727_(_067464_, _067465_, _067466_);
  or g_124728_(_067463_, _067466_, _067467_);
  xor g_124729_(out[284], out[556], _067468_);
  or g_124730_(_067443_, _067468_, _067469_);
  or g_124731_(_067442_, _067454_, _067470_);
  or g_124732_(_067469_, _067470_, _067471_);
  or g_124733_(_067446_, _067452_, _067472_);
  or g_124734_(_067455_, _067472_, _067474_);
  or g_124735_(_067471_, _067474_, _067475_);
  or g_124736_(_067467_, _067475_, _067476_);
  or g_124737_(_067459_, _067476_, _067477_);
  xor g_124738_(out[258], out[546], _067478_);
  xor g_124739_(out[256], out[544], _067479_);
  xor g_124740_(out[265], out[553], _067480_);
  xor g_124741_(out[264], out[552], _067481_);
  xor g_124742_(out[261], out[549], _067482_);
  xor g_124743_(out[270], out[558], _067483_);
  xor g_124744_(out[269], out[557], _067485_);
  xor g_124745_(out[271], out[559], _067486_);
  xor g_124746_(out[266], out[554], _067487_);
  xor g_124747_(out[262], out[550], _067488_);
  xor g_124748_(out[259], out[547], _067489_);
  and g_124749_(_098250_, out[555], _067490_);
  and g_124750_(out[267], _049543_, _067491_);
  xor g_124751_(out[260], out[548], _067492_);
  xor g_124752_(out[257], out[545], _067493_);
  or g_124753_(_067483_, _067492_, _067494_);
  or g_124754_(_067481_, _067485_, _067496_);
  or g_124755_(_067478_, _067487_, _067497_);
  or g_124756_(_067496_, _067497_, _067498_);
  or g_124757_(_067480_, _067489_, _067499_);
  or g_124758_(_067479_, _067482_, _067500_);
  or g_124759_(_067499_, _067500_, _067501_);
  or g_124760_(_067498_, _067501_, _067502_);
  xor g_124761_(out[268], out[556], _067503_);
  or g_124762_(_067490_, _067503_, _067504_);
  xor g_124763_(out[263], out[551], _067505_);
  or g_124764_(_067488_, _067505_, _067507_);
  or g_124765_(_067504_, _067507_, _067508_);
  or g_124766_(_067491_, _067493_, _067509_);
  or g_124767_(_067486_, _067509_, _067510_);
  or g_124768_(_067508_, _067510_, _067511_);
  or g_124769_(_067502_, _067511_, _067512_);
  or g_124770_(_067494_, _067512_, _067513_);
  xor g_124771_(out[247], out[551], _067514_);
  and g_124772_(_098239_, out[555], _067515_);
  xor g_124773_(out[254], out[558], _067516_);
  xor g_124774_(out[248], out[552], _067518_);
  xor g_124775_(out[241], out[545], _067519_);
  xor g_124776_(out[253], out[557], _067520_);
  xor g_124777_(out[249], out[553], _067521_);
  xor g_124778_(out[244], out[548], _067522_);
  xor g_124779_(out[242], out[546], _067523_);
  and g_124780_(out[251], _049543_, _067524_);
  xor g_124781_(out[243], out[547], _067525_);
  xor g_124782_(out[246], out[550], _067526_);
  xor g_124783_(out[255], out[559], _067527_);
  xor g_124784_(out[250], out[554], _067529_);
  xor g_124785_(out[245], out[549], _067530_);
  xor g_124786_(out[240], out[544], _067531_);
  or g_124787_(_067516_, _067522_, _067532_);
  or g_124788_(_067518_, _067520_, _067533_);
  or g_124789_(_067523_, _067529_, _067534_);
  or g_124790_(_067533_, _067534_, _067535_);
  or g_124791_(_067521_, _067525_, _067536_);
  or g_124792_(_067530_, _067531_, _067537_);
  or g_124793_(_067536_, _067537_, _067538_);
  or g_124794_(_067535_, _067538_, _067540_);
  xor g_124795_(out[252], out[556], _067541_);
  or g_124796_(_067515_, _067541_, _067542_);
  or g_124797_(_067514_, _067526_, _067543_);
  or g_124798_(_067542_, _067543_, _067544_);
  or g_124799_(_067519_, _067524_, _067545_);
  or g_124800_(_067527_, _067545_, _067546_);
  or g_124801_(_067544_, _067546_, _067547_);
  or g_124802_(_067540_, _067547_, _067548_);
  or g_124803_(_067532_, _067548_, _067549_);
  xor g_124804_(out[236], out[556], _067551_);
  and g_124805_(_098228_, out[555], _067552_);
  xor g_124806_(out[232], out[552], _067553_);
  xor g_124807_(out[230], out[550], _067554_);
  xor g_124808_(out[237], out[557], _067555_);
  xor g_124809_(out[238], out[558], _067556_);
  xor g_124810_(out[226], out[546], _067557_);
  xor g_124811_(out[233], out[553], _067558_);
  xor g_124812_(out[229], out[549], _067559_);
  xor g_124813_(out[225], out[545], _067560_);
  and g_124814_(out[235], _049543_, _067562_);
  or g_124815_(_067553_, _067555_, _067563_);
  xor g_124816_(out[239], out[559], _067564_);
  xor g_124817_(out[234], out[554], _067565_);
  xor g_124818_(out[228], out[548], _067566_);
  xor g_124819_(out[227], out[547], _067567_);
  xor g_124820_(out[224], out[544], _067568_);
  or g_124821_(_067557_, _067565_, _067569_);
  or g_124822_(_067563_, _067569_, _067570_);
  or g_124823_(_067558_, _067567_, _067571_);
  or g_124824_(_067559_, _067571_, _067573_);
  or g_124825_(_067570_, _067573_, _067574_);
  or g_124826_(_067556_, _067566_, _067575_);
  or g_124827_(_067574_, _067575_, _067576_);
  or g_124828_(_067551_, _067552_, _067577_);
  xor g_124829_(out[231], out[551], _067578_);
  or g_124830_(_067554_, _067578_, _067579_);
  or g_124831_(_067577_, _067579_, _067580_);
  or g_124832_(_067560_, _067562_, _067581_);
  or g_124833_(_067564_, _067581_, _067582_);
  or g_124834_(_067580_, _067582_, _067584_);
  or g_124835_(_067568_, _067584_, _067585_);
  or g_124836_(_067576_, _067585_, _067586_);
  xor g_124837_(out[215], out[551], _067587_);
  and g_124838_(_098217_, out[555], _067588_);
  xor g_124839_(out[222], out[558], _067589_);
  xor g_124840_(out[216], out[552], _067590_);
  xor g_124841_(out[209], out[545], _067591_);
  xor g_124842_(out[221], out[557], _067592_);
  xor g_124843_(out[217], out[553], _067593_);
  xor g_124844_(out[212], out[548], _067595_);
  xor g_124845_(out[210], out[546], _067596_);
  and g_124846_(out[219], _049543_, _067597_);
  xor g_124847_(out[211], out[547], _067598_);
  xor g_124848_(out[214], out[550], _067599_);
  xor g_124849_(out[223], out[559], _067600_);
  xor g_124850_(out[218], out[554], _067601_);
  xor g_124851_(out[213], out[549], _067602_);
  xor g_124852_(out[208], out[544], _067603_);
  or g_124853_(_067589_, _067595_, _067604_);
  or g_124854_(_067590_, _067592_, _067606_);
  or g_124855_(_067596_, _067601_, _067607_);
  or g_124856_(_067606_, _067607_, _067608_);
  or g_124857_(_067593_, _067598_, _067609_);
  or g_124858_(_067602_, _067603_, _067610_);
  or g_124859_(_067609_, _067610_, _067611_);
  or g_124860_(_067608_, _067611_, _067612_);
  xor g_124861_(out[220], out[556], _067613_);
  or g_124862_(_067588_, _067613_, _067614_);
  or g_124863_(_067587_, _067599_, _067615_);
  or g_124864_(_067614_, _067615_, _067617_);
  or g_124865_(_067591_, _067597_, _067618_);
  or g_124866_(_067600_, _067618_, _067619_);
  or g_124867_(_067617_, _067619_, _067620_);
  or g_124868_(_067612_, _067620_, _067621_);
  or g_124869_(_067604_, _067621_, _067622_);
  xor g_124870_(out[193], out[545], _067623_);
  and g_124871_(out[203], _049543_, _067624_);
  xor g_124872_(out[201], out[553], _067625_);
  xor g_124873_(out[192], out[544], _067626_);
  xor g_124874_(out[206], out[558], _067628_);
  xor g_124875_(out[196], out[548], _067629_);
  or g_124876_(_067628_, _067629_, _067630_);
  xor g_124877_(out[205], out[557], _067631_);
  xor g_124878_(out[195], out[547], _067632_);
  and g_124879_(_098206_, out[555], _067633_);
  xor g_124880_(out[198], out[550], _067634_);
  xor g_124881_(out[202], out[554], _067635_);
  xor g_124882_(out[197], out[549], _067636_);
  xor g_124883_(out[207], out[559], _067637_);
  xor g_124884_(out[200], out[552], _067639_);
  or g_124885_(_067631_, _067639_, _067640_);
  xor g_124886_(out[194], out[546], _067641_);
  or g_124887_(_067635_, _067641_, _067642_);
  or g_124888_(_067640_, _067642_, _067643_);
  or g_124889_(_067625_, _067632_, _067644_);
  or g_124890_(_067636_, _067644_, _067645_);
  or g_124891_(_067643_, _067645_, _067646_);
  or g_124892_(_067630_, _067646_, _067647_);
  xor g_124893_(out[204], out[556], _067648_);
  or g_124894_(_067633_, _067648_, _067650_);
  xor g_124895_(out[199], out[551], _067651_);
  or g_124896_(_067634_, _067651_, _067652_);
  or g_124897_(_067650_, _067652_, _067653_);
  or g_124898_(_067623_, _067624_, _067654_);
  or g_124899_(_067637_, _067654_, _067655_);
  or g_124900_(_067653_, _067655_, _067656_);
  or g_124901_(_067626_, _067656_, _067657_);
  or g_124902_(_067647_, _067657_, _067658_);
  xor g_124903_(out[183], out[551], _067659_);
  and g_124904_(_098195_, out[555], _067661_);
  xor g_124905_(out[190], out[558], _067662_);
  xor g_124906_(out[184], out[552], _067663_);
  xor g_124907_(out[177], out[545], _067664_);
  xor g_124908_(out[189], out[557], _067665_);
  xor g_124909_(out[185], out[553], _067666_);
  xor g_124910_(out[180], out[548], _067667_);
  xor g_124911_(out[178], out[546], _067668_);
  and g_124912_(out[187], _049543_, _067669_);
  xor g_124913_(out[179], out[547], _067670_);
  xor g_124914_(out[182], out[550], _067672_);
  xor g_124915_(out[191], out[559], _067673_);
  xor g_124916_(out[186], out[554], _067674_);
  xor g_124917_(out[181], out[549], _067675_);
  xor g_124918_(out[176], out[544], _067676_);
  or g_124919_(_067662_, _067667_, _067677_);
  or g_124920_(_067663_, _067665_, _067678_);
  or g_124921_(_067668_, _067674_, _067679_);
  or g_124922_(_067678_, _067679_, _067680_);
  or g_124923_(_067666_, _067670_, _067681_);
  or g_124924_(_067675_, _067676_, _067683_);
  or g_124925_(_067681_, _067683_, _067684_);
  or g_124926_(_067680_, _067684_, _067685_);
  xor g_124927_(out[188], out[556], _067686_);
  or g_124928_(_067661_, _067686_, _067687_);
  or g_124929_(_067659_, _067672_, _067688_);
  or g_124930_(_067687_, _067688_, _067689_);
  or g_124931_(_067664_, _067669_, _067690_);
  or g_124932_(_067673_, _067690_, _067691_);
  or g_124933_(_067689_, _067691_, _067692_);
  or g_124934_(_067685_, _067692_, _067694_);
  or g_124935_(_067677_, _067694_, _067695_);
  xor g_124936_(out[161], out[545], _067696_);
  and g_124937_(out[171], _049543_, _067697_);
  xor g_124938_(out[169], out[553], _067698_);
  xor g_124939_(out[160], out[544], _067699_);
  xor g_124940_(out[174], out[558], _067700_);
  xor g_124941_(out[164], out[548], _067701_);
  or g_124942_(_067700_, _067701_, _067702_);
  xor g_124943_(out[173], out[557], _067703_);
  xor g_124944_(out[163], out[547], _067705_);
  and g_124945_(_098184_, out[555], _067706_);
  xor g_124946_(out[166], out[550], _067707_);
  xor g_124947_(out[170], out[554], _067708_);
  xor g_124948_(out[165], out[549], _067709_);
  xor g_124949_(out[175], out[559], _067710_);
  xor g_124950_(out[168], out[552], _067711_);
  or g_124951_(_067703_, _067711_, _067712_);
  xor g_124952_(out[162], out[546], _067713_);
  or g_124953_(_067708_, _067713_, _067714_);
  or g_124954_(_067712_, _067714_, _067716_);
  or g_124955_(_067698_, _067705_, _067717_);
  or g_124956_(_067709_, _067717_, _067718_);
  or g_124957_(_067716_, _067718_, _067719_);
  or g_124958_(_067702_, _067719_, _067720_);
  xor g_124959_(out[172], out[556], _067721_);
  or g_124960_(_067706_, _067721_, _067722_);
  xor g_124961_(out[167], out[551], _067723_);
  or g_124962_(_067707_, _067723_, _067724_);
  or g_124963_(_067722_, _067724_, _067725_);
  or g_124964_(_067696_, _067697_, _067727_);
  or g_124965_(_067710_, _067727_, _067728_);
  or g_124966_(_067725_, _067728_, _067729_);
  or g_124967_(_067699_, _067729_, _067730_);
  or g_124968_(_067720_, _067730_, _067731_);
  xor g_124969_(out[151], out[551], _067732_);
  and g_124970_(_098173_, out[555], _067733_);
  xor g_124971_(out[158], out[558], _067734_);
  xor g_124972_(out[152], out[552], _067735_);
  xor g_124973_(out[145], out[545], _067736_);
  xor g_124974_(out[157], out[557], _067738_);
  xor g_124975_(out[153], out[553], _067739_);
  xor g_124976_(out[148], out[548], _067740_);
  xor g_124977_(out[146], out[546], _067741_);
  and g_124978_(out[155], _049543_, _067742_);
  xor g_124979_(out[147], out[547], _067743_);
  xor g_124980_(out[150], out[550], _067744_);
  xor g_124981_(out[159], out[559], _067745_);
  xor g_124982_(out[154], out[554], _067746_);
  xor g_124983_(out[149], out[549], _067747_);
  xor g_124984_(out[144], out[544], _067749_);
  or g_124985_(_067734_, _067740_, _067750_);
  or g_124986_(_067735_, _067738_, _067751_);
  or g_124987_(_067741_, _067746_, _067752_);
  or g_124988_(_067751_, _067752_, _067753_);
  or g_124989_(_067739_, _067743_, _067754_);
  or g_124990_(_067747_, _067749_, _067755_);
  or g_124991_(_067754_, _067755_, _067756_);
  or g_124992_(_067753_, _067756_, _067757_);
  xor g_124993_(out[156], out[556], _067758_);
  or g_124994_(_067733_, _067758_, _067760_);
  or g_124995_(_067732_, _067744_, _067761_);
  or g_124996_(_067760_, _067761_, _067762_);
  or g_124997_(_067736_, _067742_, _067763_);
  or g_124998_(_067745_, _067763_, _067764_);
  or g_124999_(_067762_, _067764_, _067765_);
  or g_125000_(_067757_, _067765_, _067766_);
  or g_125001_(_067750_, _067766_, _067767_);
  and g_125002_(out[139], _049543_, _067768_);
  xor g_125003_(out[138], out[554], _067769_);
  xor g_125004_(out[143], out[559], _067771_);
  xor g_125005_(out[128], out[544], _067772_);
  xor g_125006_(out[129], out[545], _067773_);
  xor g_125007_(out[130], out[546], _067774_);
  xor g_125008_(out[131], out[547], _067775_);
  xor g_125009_(out[137], out[553], _067776_);
  xor g_125010_(out[142], out[558], _067777_);
  and g_125011_(_098162_, out[555], _067778_);
  xor g_125012_(out[133], out[549], _067779_);
  xor g_125013_(out[134], out[550], _067780_);
  xor g_125014_(out[132], out[548], _067782_);
  xor g_125015_(out[141], out[557], _067783_);
  xor g_125016_(out[136], out[552], _067784_);
  or g_125017_(_067783_, _067784_, _067785_);
  or g_125018_(_067769_, _067774_, _067786_);
  or g_125019_(_067785_, _067786_, _067787_);
  or g_125020_(_067775_, _067776_, _067788_);
  or g_125021_(_067779_, _067788_, _067789_);
  or g_125022_(_067787_, _067789_, _067790_);
  or g_125023_(_067777_, _067782_, _067791_);
  or g_125024_(_067790_, _067791_, _067793_);
  xor g_125025_(out[140], out[556], _067794_);
  or g_125026_(_067778_, _067794_, _067795_);
  xor g_125027_(out[135], out[551], _067796_);
  or g_125028_(_067780_, _067796_, _067797_);
  or g_125029_(_067795_, _067797_, _067798_);
  or g_125030_(_067768_, _067773_, _067799_);
  or g_125031_(_067771_, _067799_, _067800_);
  or g_125032_(_067798_, _067800_, _067801_);
  or g_125033_(_067772_, _067801_, _067802_);
  or g_125034_(_067793_, _067802_, _067804_);
  xor g_125035_(out[119], out[551], _067805_);
  and g_125036_(_098151_, out[555], _067806_);
  xor g_125037_(out[126], out[558], _067807_);
  xor g_125038_(out[120], out[552], _067808_);
  xor g_125039_(out[113], out[545], _067809_);
  xor g_125040_(out[125], out[557], _067810_);
  xor g_125041_(out[121], out[553], _067811_);
  xor g_125042_(out[116], out[548], _067812_);
  xor g_125043_(out[114], out[546], _067813_);
  and g_125044_(out[123], _049543_, _067815_);
  xor g_125045_(out[115], out[547], _067816_);
  xor g_125046_(out[118], out[550], _067817_);
  xor g_125047_(out[127], out[559], _067818_);
  xor g_125048_(out[122], out[554], _067819_);
  xor g_125049_(out[117], out[549], _067820_);
  xor g_125050_(out[112], out[544], _067821_);
  or g_125051_(_067807_, _067812_, _067822_);
  or g_125052_(_067808_, _067810_, _067823_);
  or g_125053_(_067813_, _067819_, _067824_);
  or g_125054_(_067823_, _067824_, _067826_);
  or g_125055_(_067811_, _067816_, _067827_);
  or g_125056_(_067820_, _067821_, _067828_);
  or g_125057_(_067827_, _067828_, _067829_);
  or g_125058_(_067826_, _067829_, _067830_);
  xor g_125059_(out[124], out[556], _067831_);
  or g_125060_(_067806_, _067831_, _067832_);
  or g_125061_(_067805_, _067817_, _067833_);
  or g_125062_(_067832_, _067833_, _067834_);
  or g_125063_(_067809_, _067815_, _067835_);
  or g_125064_(_067818_, _067835_, _067837_);
  or g_125065_(_067834_, _067837_, _067838_);
  or g_125066_(_067830_, _067838_, _067839_);
  or g_125067_(_067822_, _067839_, _067840_);
  xor g_125068_(out[97], out[545], _067841_);
  and g_125069_(out[107], _049543_, _067842_);
  xor g_125070_(out[105], out[553], _067843_);
  xor g_125071_(out[96], out[544], _067844_);
  xor g_125072_(out[110], out[558], _067845_);
  xor g_125073_(out[100], out[548], _067846_);
  or g_125074_(_067845_, _067846_, _067848_);
  xor g_125075_(out[109], out[557], _067849_);
  xor g_125076_(out[99], out[547], _067850_);
  and g_125077_(_098140_, out[555], _067851_);
  xor g_125078_(out[102], out[550], _067852_);
  xor g_125079_(out[106], out[554], _067853_);
  xor g_125080_(out[101], out[549], _067854_);
  xor g_125081_(out[111], out[559], _067855_);
  xor g_125082_(out[104], out[552], _067856_);
  or g_125083_(_067849_, _067856_, _067857_);
  xor g_125084_(out[98], out[546], _067859_);
  or g_125085_(_067853_, _067859_, _067860_);
  or g_125086_(_067857_, _067860_, _067861_);
  or g_125087_(_067843_, _067850_, _067862_);
  or g_125088_(_067854_, _067862_, _067863_);
  or g_125089_(_067861_, _067863_, _067864_);
  or g_125090_(_067848_, _067864_, _067865_);
  xor g_125091_(out[108], out[556], _067866_);
  or g_125092_(_067851_, _067866_, _067867_);
  xor g_125093_(out[103], out[551], _067868_);
  or g_125094_(_067852_, _067868_, _067870_);
  or g_125095_(_067867_, _067870_, _067871_);
  or g_125096_(_067841_, _067842_, _067872_);
  or g_125097_(_067855_, _067872_, _067873_);
  or g_125098_(_067871_, _067873_, _067874_);
  or g_125099_(_067844_, _067874_, _067875_);
  or g_125100_(_067865_, _067875_, _067876_);
  not g_125101_(_067876_, _067877_);
  xor g_125102_(out[87], out[551], _067878_);
  and g_125103_(_098129_, out[555], _067879_);
  xor g_125104_(out[94], out[558], _067881_);
  xor g_125105_(out[88], out[552], _067882_);
  xor g_125106_(out[81], out[545], _067883_);
  xor g_125107_(out[93], out[557], _067884_);
  xor g_125108_(out[89], out[553], _067885_);
  xor g_125109_(out[84], out[548], _067886_);
  xor g_125110_(out[82], out[546], _067887_);
  and g_125111_(out[91], _049543_, _067888_);
  xor g_125112_(out[83], out[547], _067889_);
  xor g_125113_(out[86], out[550], _067890_);
  xor g_125114_(out[95], out[559], _067892_);
  xor g_125115_(out[90], out[554], _067893_);
  xor g_125116_(out[85], out[549], _067894_);
  xor g_125117_(out[80], out[544], _067895_);
  or g_125118_(_067881_, _067886_, _067896_);
  or g_125119_(_067882_, _067884_, _067897_);
  or g_125120_(_067887_, _067893_, _067898_);
  or g_125121_(_067897_, _067898_, _067899_);
  or g_125122_(_067885_, _067889_, _067900_);
  or g_125123_(_067894_, _067895_, _067901_);
  or g_125124_(_067900_, _067901_, _067903_);
  or g_125125_(_067899_, _067903_, _067904_);
  xor g_125126_(out[92], out[556], _067905_);
  or g_125127_(_067879_, _067905_, _067906_);
  or g_125128_(_067878_, _067890_, _067907_);
  or g_125129_(_067906_, _067907_, _067908_);
  or g_125130_(_067883_, _067888_, _067909_);
  or g_125131_(_067892_, _067909_, _067910_);
  or g_125132_(_067908_, _067910_, _067911_);
  or g_125133_(_067904_, _067911_, _067912_);
  or g_125134_(_067896_, _067912_, _067914_);
  not g_125135_(_067914_, _067915_);
  xor g_125136_(out[65], out[545], _067916_);
  and g_125137_(out[75], _049543_, _067917_);
  xor g_125138_(out[73], out[553], _067918_);
  xor g_125139_(out[64], out[544], _067919_);
  xor g_125140_(out[78], out[558], _067920_);
  xor g_125141_(out[68], out[548], _067921_);
  or g_125142_(_067920_, _067921_, _067922_);
  xor g_125143_(out[77], out[557], _067923_);
  xor g_125144_(out[67], out[547], _067925_);
  and g_125145_(_098118_, out[555], _067926_);
  xor g_125146_(out[70], out[550], _067927_);
  xor g_125147_(out[74], out[554], _067928_);
  xor g_125148_(out[69], out[549], _067929_);
  xor g_125149_(out[79], out[559], _067930_);
  xor g_125150_(out[72], out[552], _067931_);
  or g_125151_(_067923_, _067931_, _067932_);
  xor g_125152_(out[66], out[546], _067933_);
  or g_125153_(_067928_, _067933_, _067934_);
  or g_125154_(_067932_, _067934_, _067936_);
  or g_125155_(_067918_, _067925_, _067937_);
  or g_125156_(_067929_, _067937_, _067938_);
  or g_125157_(_067936_, _067938_, _067939_);
  or g_125158_(_067922_, _067939_, _067940_);
  xor g_125159_(out[76], out[556], _067941_);
  or g_125160_(_067926_, _067941_, _067942_);
  xor g_125161_(out[71], out[551], _067943_);
  or g_125162_(_067927_, _067943_, _067944_);
  or g_125163_(_067942_, _067944_, _067945_);
  or g_125164_(_067916_, _067917_, _067947_);
  or g_125165_(_067930_, _067947_, _067948_);
  or g_125166_(_067945_, _067948_, _067949_);
  or g_125167_(_067919_, _067949_, _067950_);
  or g_125168_(_067940_, _067950_, _067951_);
  not g_125169_(_067951_, _067952_);
  xor g_125170_(out[55], out[551], _067953_);
  and g_125171_(_098107_, out[555], _067954_);
  xor g_125172_(out[62], out[558], _067955_);
  xor g_125173_(out[56], out[552], _067956_);
  xor g_125174_(out[49], out[545], _067958_);
  xor g_125175_(out[61], out[557], _067959_);
  xor g_125176_(out[57], out[553], _067960_);
  xor g_125177_(out[52], out[548], _067961_);
  xor g_125178_(out[50], out[546], _067962_);
  and g_125179_(out[59], _049543_, _067963_);
  xor g_125180_(out[51], out[547], _067964_);
  xor g_125181_(out[54], out[550], _067965_);
  xor g_125182_(out[63], out[559], _067966_);
  xor g_125183_(out[58], out[554], _067967_);
  xor g_125184_(out[53], out[549], _067969_);
  xor g_125185_(out[48], out[544], _067970_);
  or g_125186_(_067955_, _067961_, _067971_);
  or g_125187_(_067956_, _067959_, _067972_);
  or g_125188_(_067962_, _067967_, _067973_);
  or g_125189_(_067972_, _067973_, _067974_);
  or g_125190_(_067960_, _067964_, _067975_);
  or g_125191_(_067969_, _067970_, _067976_);
  or g_125192_(_067975_, _067976_, _067977_);
  or g_125193_(_067974_, _067977_, _067978_);
  xor g_125194_(out[60], out[556], _067980_);
  or g_125195_(_067954_, _067980_, _067981_);
  or g_125196_(_067953_, _067965_, _067982_);
  or g_125197_(_067981_, _067982_, _067983_);
  or g_125198_(_067958_, _067963_, _067984_);
  or g_125199_(_067966_, _067984_, _067985_);
  or g_125200_(_067983_, _067985_, _067986_);
  or g_125201_(_067978_, _067986_, _067987_);
  or g_125202_(_067971_, _067987_, _067988_);
  and g_125203_(out[43], _049543_, _067989_);
  xor g_125204_(out[36], out[548], _067991_);
  xor g_125205_(out[46], out[558], _067992_);
  or g_125206_(_067991_, _067992_, _067993_);
  xor g_125207_(out[45], out[557], _067994_);
  xor g_125208_(out[35], out[547], _067995_);
  xor g_125209_(out[32], out[544], _067996_);
  and g_125210_(_098096_, out[555], _067997_);
  xor g_125211_(out[42], out[554], _067998_);
  xor g_125212_(out[47], out[559], _067999_);
  xor g_125213_(out[38], out[550], _068000_);
  xor g_125214_(out[37], out[549], _068002_);
  xor g_125215_(out[40], out[552], _068003_);
  or g_125216_(_067994_, _068003_, _068004_);
  xor g_125217_(out[34], out[546], _068005_);
  xor g_125218_(out[41], out[553], _068006_);
  xor g_125219_(out[33], out[545], _068007_);
  or g_125220_(_067998_, _068005_, _068008_);
  or g_125221_(_068004_, _068008_, _068009_);
  or g_125222_(_067995_, _068006_, _068010_);
  or g_125223_(_068002_, _068010_, _068011_);
  or g_125224_(_068009_, _068011_, _068013_);
  or g_125225_(_067993_, _068013_, _068014_);
  xor g_125226_(out[44], out[556], _068015_);
  or g_125227_(_067997_, _068015_, _068016_);
  xor g_125228_(out[39], out[551], _068017_);
  or g_125229_(_068000_, _068017_, _068018_);
  or g_125230_(_068016_, _068018_, _068019_);
  or g_125231_(_067989_, _068007_, _068020_);
  or g_125232_(_067999_, _068020_, _068021_);
  or g_125233_(_068019_, _068021_, _068022_);
  or g_125234_(_067996_, _068022_, _068024_);
  or g_125235_(_068014_, _068024_, _068025_);
  not g_125236_(_068025_, _068026_);
  xor g_125237_(out[23], out[551], _068027_);
  and g_125238_(_098063_, out[555], _068028_);
  xor g_125239_(out[30], out[558], _068029_);
  xor g_125240_(out[24], out[552], _068030_);
  xor g_125241_(out[17], out[545], _068031_);
  xor g_125242_(out[29], out[557], _068032_);
  xor g_125243_(out[25], out[553], _068033_);
  xor g_125244_(out[20], out[548], _068035_);
  xor g_125245_(out[18], out[546], _068036_);
  and g_125246_(out[27], _049543_, _068037_);
  xor g_125247_(out[19], out[547], _068038_);
  xor g_125248_(out[22], out[550], _068039_);
  xor g_125249_(out[31], out[559], _068040_);
  xor g_125250_(out[26], out[554], _068041_);
  xor g_125251_(out[21], out[549], _068042_);
  xor g_125252_(out[16], out[544], _068043_);
  or g_125253_(_068029_, _068035_, _068044_);
  or g_125254_(_068030_, _068032_, _068046_);
  or g_125255_(_068036_, _068041_, _068047_);
  or g_125256_(_068046_, _068047_, _068048_);
  or g_125257_(_068033_, _068038_, _068049_);
  or g_125258_(_068042_, _068043_, _068050_);
  or g_125259_(_068049_, _068050_, _068051_);
  or g_125260_(_068048_, _068051_, _068052_);
  xor g_125261_(out[28], out[556], _068053_);
  or g_125262_(_068028_, _068053_, _068054_);
  or g_125263_(_068027_, _068039_, _068055_);
  or g_125264_(_068054_, _068055_, _068057_);
  or g_125265_(_068031_, _068037_, _068058_);
  or g_125266_(_068040_, _068058_, _068059_);
  or g_125267_(_068057_, _068059_, _068060_);
  or g_125268_(_068052_, _068060_, _068061_);
  or g_125269_(_068044_, _068061_, _068062_);
  xor g_125270_(out[1], out[545], _068063_);
  and g_125271_(out[11], _049543_, _068064_);
  xor g_125272_(out[9], out[553], _068065_);
  xor g_125273_(out[0], out[544], _068066_);
  xor g_125274_(out[14], out[558], _068068_);
  xor g_125275_(out[4], out[548], _068069_);
  or g_125276_(_068068_, _068069_, _068070_);
  xor g_125277_(out[13], out[557], _068071_);
  xor g_125278_(out[3], out[547], _068072_);
  and g_125279_(_098041_, out[555], _068073_);
  xor g_125280_(out[6], out[550], _068074_);
  xor g_125281_(out[10], out[554], _068075_);
  xor g_125282_(out[5], out[549], _068076_);
  xor g_125283_(out[15], out[559], _068077_);
  xor g_125284_(out[8], out[552], _068079_);
  or g_125285_(_068071_, _068079_, _068080_);
  xor g_125286_(out[2], out[546], _068081_);
  or g_125287_(_068075_, _068081_, _068082_);
  or g_125288_(_068080_, _068082_, _068083_);
  or g_125289_(_068065_, _068072_, _068084_);
  or g_125290_(_068076_, _068084_, _068085_);
  or g_125291_(_068083_, _068085_, _068086_);
  or g_125292_(_068070_, _068086_, _068087_);
  xor g_125293_(out[12], out[556], _068088_);
  or g_125294_(_068073_, _068088_, _068090_);
  xor g_125295_(out[7], out[551], _068091_);
  or g_125296_(_068074_, _068091_, _068092_);
  or g_125297_(_068090_, _068092_, _068093_);
  or g_125298_(_068063_, _068064_, _068094_);
  or g_125299_(_068077_, _068094_, _068095_);
  or g_125300_(_068093_, _068095_, _068096_);
  or g_125301_(_068066_, _068096_, _068097_);
  or g_125302_(_068087_, _068097_, _068098_);
  xor g_125303_(out[465], out[529], _068099_);
  and g_125304_(out[475], _049532_, _068101_);
  xor g_125305_(out[473], out[537], _068102_);
  xor g_125306_(out[464], out[528], _068103_);
  xor g_125307_(out[478], out[542], _068104_);
  xor g_125308_(out[468], out[532], _068105_);
  or g_125309_(_068104_, _068105_, _068106_);
  xor g_125310_(out[477], out[541], _068107_);
  xor g_125311_(out[467], out[531], _068108_);
  and g_125312_(_049499_, out[539], _068109_);
  xor g_125313_(out[470], out[534], _068110_);
  xor g_125314_(out[474], out[538], _068112_);
  xor g_125315_(out[469], out[533], _068113_);
  xor g_125316_(out[479], out[543], _068114_);
  xor g_125317_(out[472], out[536], _068115_);
  or g_125318_(_068107_, _068115_, _068116_);
  xor g_125319_(out[466], out[530], _068117_);
  or g_125320_(_068112_, _068117_, _068118_);
  or g_125321_(_068116_, _068118_, _068119_);
  or g_125322_(_068102_, _068108_, _068120_);
  or g_125323_(_068113_, _068120_, _068121_);
  or g_125324_(_068119_, _068121_, _068123_);
  or g_125325_(_068106_, _068123_, _068124_);
  xor g_125326_(out[476], out[540], _068125_);
  or g_125327_(_068109_, _068125_, _068126_);
  xor g_125328_(out[471], out[535], _068127_);
  or g_125329_(_068110_, _068127_, _068128_);
  or g_125330_(_068126_, _068128_, _068129_);
  or g_125331_(_068099_, _068101_, _068130_);
  or g_125332_(_068114_, _068130_, _068131_);
  or g_125333_(_068129_, _068131_, _068132_);
  or g_125334_(_068103_, _068132_, _068134_);
  or g_125335_(_068124_, _068134_, _068135_);
  not g_125336_(_068135_, _068136_);
  xor g_125337_(out[455], out[535], _068137_);
  and g_125338_(_049477_, out[539], _068138_);
  xor g_125339_(out[462], out[542], _068139_);
  xor g_125340_(out[456], out[536], _068140_);
  xor g_125341_(out[449], out[529], _068141_);
  xor g_125342_(out[461], out[541], _068142_);
  xor g_125343_(out[457], out[537], _068143_);
  xor g_125344_(out[452], out[532], _068145_);
  xor g_125345_(out[450], out[530], _068146_);
  and g_125346_(out[459], _049532_, _068147_);
  xor g_125347_(out[451], out[531], _068148_);
  xor g_125348_(out[454], out[534], _068149_);
  xor g_125349_(out[463], out[543], _068150_);
  xor g_125350_(out[458], out[538], _068151_);
  xor g_125351_(out[453], out[533], _068152_);
  xor g_125352_(out[448], out[528], _068153_);
  or g_125353_(_068139_, _068145_, _068154_);
  or g_125354_(_068140_, _068142_, _068156_);
  or g_125355_(_068146_, _068151_, _068157_);
  or g_125356_(_068156_, _068157_, _068158_);
  or g_125357_(_068143_, _068148_, _068159_);
  or g_125358_(_068152_, _068153_, _068160_);
  or g_125359_(_068159_, _068160_, _068161_);
  or g_125360_(_068158_, _068161_, _068162_);
  xor g_125361_(out[460], out[540], _068163_);
  or g_125362_(_068138_, _068163_, _068164_);
  or g_125363_(_068137_, _068149_, _068165_);
  or g_125364_(_068164_, _068165_, _068167_);
  or g_125365_(_068141_, _068147_, _068168_);
  or g_125366_(_068150_, _068168_, _068169_);
  or g_125367_(_068167_, _068169_, _068170_);
  or g_125368_(_068162_, _068170_, _068171_);
  or g_125369_(_068154_, _068171_, _068172_);
  not g_125370_(_068172_, _068173_);
  xor g_125371_(out[433], out[529], _068174_);
  and g_125372_(out[443], _049532_, _068175_);
  xor g_125373_(out[441], out[537], _068176_);
  xor g_125374_(out[432], out[528], _068178_);
  xor g_125375_(out[446], out[542], _068179_);
  xor g_125376_(out[436], out[532], _068180_);
  or g_125377_(_068179_, _068180_, _068181_);
  xor g_125378_(out[445], out[541], _068182_);
  xor g_125379_(out[435], out[531], _068183_);
  and g_125380_(_049466_, out[539], _068184_);
  xor g_125381_(out[438], out[534], _068185_);
  xor g_125382_(out[442], out[538], _068186_);
  xor g_125383_(out[437], out[533], _068187_);
  xor g_125384_(out[447], out[543], _068189_);
  xor g_125385_(out[440], out[536], _068190_);
  or g_125386_(_068182_, _068190_, _068191_);
  xor g_125387_(out[434], out[530], _068192_);
  or g_125388_(_068186_, _068192_, _068193_);
  or g_125389_(_068191_, _068193_, _068194_);
  or g_125390_(_068176_, _068183_, _068195_);
  or g_125391_(_068187_, _068195_, _068196_);
  or g_125392_(_068194_, _068196_, _068197_);
  or g_125393_(_068181_, _068197_, _068198_);
  xor g_125394_(out[444], out[540], _068200_);
  or g_125395_(_068184_, _068200_, _068201_);
  xor g_125396_(out[439], out[535], _068202_);
  or g_125397_(_068185_, _068202_, _068203_);
  or g_125398_(_068201_, _068203_, _068204_);
  or g_125399_(_068174_, _068175_, _068205_);
  or g_125400_(_068189_, _068205_, _068206_);
  or g_125401_(_068204_, _068206_, _068207_);
  or g_125402_(_068178_, _068207_, _068208_);
  or g_125403_(_068198_, _068208_, _068209_);
  xor g_125404_(out[423], out[535], _068211_);
  and g_125405_(_049455_, out[539], _068212_);
  xor g_125406_(out[430], out[542], _068213_);
  xor g_125407_(out[424], out[536], _068214_);
  xor g_125408_(out[417], out[529], _068215_);
  xor g_125409_(out[429], out[541], _068216_);
  xor g_125410_(out[425], out[537], _068217_);
  xor g_125411_(out[420], out[532], _068218_);
  xor g_125412_(out[418], out[530], _068219_);
  and g_125413_(out[427], _049532_, _068220_);
  xor g_125414_(out[419], out[531], _068222_);
  xor g_125415_(out[422], out[534], _068223_);
  xor g_125416_(out[431], out[543], _068224_);
  xor g_125417_(out[426], out[538], _068225_);
  xor g_125418_(out[421], out[533], _068226_);
  xor g_125419_(out[416], out[528], _068227_);
  or g_125420_(_068213_, _068218_, _068228_);
  or g_125421_(_068214_, _068216_, _068229_);
  or g_125422_(_068219_, _068225_, _068230_);
  or g_125423_(_068229_, _068230_, _068231_);
  or g_125424_(_068217_, _068222_, _068233_);
  or g_125425_(_068226_, _068227_, _068234_);
  or g_125426_(_068233_, _068234_, _068235_);
  or g_125427_(_068231_, _068235_, _068236_);
  xor g_125428_(out[428], out[540], _068237_);
  or g_125429_(_068212_, _068237_, _068238_);
  or g_125430_(_068211_, _068223_, _068239_);
  or g_125431_(_068238_, _068239_, _068240_);
  or g_125432_(_068215_, _068220_, _068241_);
  or g_125433_(_068224_, _068241_, _068242_);
  or g_125434_(_068240_, _068242_, _068244_);
  or g_125435_(_068236_, _068244_, _068245_);
  or g_125436_(_068228_, _068245_, _068246_);
  xor g_125437_(out[401], out[529], _068247_);
  and g_125438_(out[411], _049532_, _068248_);
  xor g_125439_(out[409], out[537], _068249_);
  xor g_125440_(out[400], out[528], _068250_);
  xor g_125441_(out[414], out[542], _068251_);
  xor g_125442_(out[404], out[532], _068252_);
  or g_125443_(_068251_, _068252_, _068253_);
  xor g_125444_(out[413], out[541], _068255_);
  xor g_125445_(out[403], out[531], _068256_);
  and g_125446_(_049444_, out[539], _068257_);
  xor g_125447_(out[406], out[534], _068258_);
  xor g_125448_(out[410], out[538], _068259_);
  xor g_125449_(out[405], out[533], _068260_);
  xor g_125450_(out[415], out[543], _068261_);
  xor g_125451_(out[408], out[536], _068262_);
  or g_125452_(_068255_, _068262_, _068263_);
  xor g_125453_(out[402], out[530], _068264_);
  or g_125454_(_068259_, _068264_, _068266_);
  or g_125455_(_068263_, _068266_, _068267_);
  or g_125456_(_068249_, _068256_, _068268_);
  or g_125457_(_068260_, _068268_, _068269_);
  or g_125458_(_068267_, _068269_, _068270_);
  or g_125459_(_068253_, _068270_, _068271_);
  xor g_125460_(out[412], out[540], _068272_);
  or g_125461_(_068257_, _068272_, _068273_);
  xor g_125462_(out[407], out[535], _068274_);
  or g_125463_(_068258_, _068274_, _068275_);
  or g_125464_(_068273_, _068275_, _068277_);
  or g_125465_(_068247_, _068248_, _068278_);
  or g_125466_(_068261_, _068278_, _068279_);
  or g_125467_(_068277_, _068279_, _068280_);
  or g_125468_(_068250_, _068280_, _068281_);
  or g_125469_(_068271_, _068281_, _068282_);
  xor g_125470_(out[391], out[535], _068283_);
  and g_125471_(_049433_, out[539], _068284_);
  xor g_125472_(out[398], out[542], _068285_);
  xor g_125473_(out[392], out[536], _068286_);
  xor g_125474_(out[385], out[529], _068288_);
  xor g_125475_(out[397], out[541], _068289_);
  xor g_125476_(out[393], out[537], _068290_);
  xor g_125477_(out[388], out[532], _068291_);
  xor g_125478_(out[386], out[530], _068292_);
  and g_125479_(out[395], _049532_, _068293_);
  xor g_125480_(out[387], out[531], _068294_);
  xor g_125481_(out[390], out[534], _068295_);
  xor g_125482_(out[399], out[543], _068296_);
  xor g_125483_(out[394], out[538], _068297_);
  xor g_125484_(out[389], out[533], _068299_);
  xor g_125485_(out[384], out[528], _068300_);
  or g_125486_(_068285_, _068291_, _068301_);
  or g_125487_(_068286_, _068289_, _068302_);
  or g_125488_(_068292_, _068297_, _068303_);
  or g_125489_(_068302_, _068303_, _068304_);
  or g_125490_(_068290_, _068294_, _068305_);
  or g_125491_(_068299_, _068300_, _068306_);
  or g_125492_(_068305_, _068306_, _068307_);
  or g_125493_(_068304_, _068307_, _068308_);
  xor g_125494_(out[396], out[540], _068310_);
  or g_125495_(_068284_, _068310_, _068311_);
  or g_125496_(_068283_, _068295_, _068312_);
  or g_125497_(_068311_, _068312_, _068313_);
  or g_125498_(_068288_, _068293_, _068314_);
  or g_125499_(_068296_, _068314_, _068315_);
  or g_125500_(_068313_, _068315_, _068316_);
  or g_125501_(_068308_, _068316_, _068317_);
  or g_125502_(_068301_, _068317_, _068318_);
  xor g_125503_(out[381], out[541], _068319_);
  xor g_125504_(out[370], out[530], _068321_);
  xor g_125505_(out[373], out[533], _068322_);
  xor g_125506_(out[377], out[537], _068323_);
  xor g_125507_(out[372], out[532], _068324_);
  xor g_125508_(out[376], out[536], _068325_);
  xor g_125509_(out[382], out[542], _068326_);
  xor g_125510_(out[374], out[534], _068327_);
  xor g_125511_(out[383], out[543], _068328_);
  xor g_125512_(out[378], out[538], _068329_);
  xor g_125513_(out[368], out[528], _068330_);
  xor g_125514_(out[371], out[531], _068332_);
  and g_125515_(_049422_, out[539], _068333_);
  and g_125516_(out[379], _049532_, _068334_);
  xor g_125517_(out[369], out[529], _068335_);
  or g_125518_(_068324_, _068326_, _068336_);
  or g_125519_(_068319_, _068325_, _068337_);
  or g_125520_(_068321_, _068329_, _068338_);
  or g_125521_(_068337_, _068338_, _068339_);
  or g_125522_(_068323_, _068332_, _068340_);
  or g_125523_(_068322_, _068330_, _068341_);
  or g_125524_(_068340_, _068341_, _068343_);
  or g_125525_(_068339_, _068343_, _068344_);
  xor g_125526_(out[380], out[540], _068345_);
  or g_125527_(_068333_, _068345_, _068346_);
  xor g_125528_(out[375], out[535], _068347_);
  or g_125529_(_068327_, _068347_, _068348_);
  or g_125530_(_068346_, _068348_, _068349_);
  or g_125531_(_068334_, _068335_, _068350_);
  or g_125532_(_068328_, _068350_, _068351_);
  or g_125533_(_068349_, _068351_, _068352_);
  or g_125534_(_068344_, _068352_, _068354_);
  or g_125535_(_068336_, _068354_, _068355_);
  not g_125536_(_068355_, _068356_);
  xor g_125537_(out[359], out[535], _068357_);
  and g_125538_(_049411_, out[539], _068358_);
  xor g_125539_(out[366], out[542], _068359_);
  xor g_125540_(out[360], out[536], _068360_);
  xor g_125541_(out[353], out[529], _068361_);
  xor g_125542_(out[365], out[541], _068362_);
  xor g_125543_(out[361], out[537], _068363_);
  xor g_125544_(out[356], out[532], _068365_);
  xor g_125545_(out[354], out[530], _068366_);
  and g_125546_(out[363], _049532_, _068367_);
  xor g_125547_(out[355], out[531], _068368_);
  xor g_125548_(out[358], out[534], _068369_);
  xor g_125549_(out[367], out[543], _068370_);
  xor g_125550_(out[362], out[538], _068371_);
  xor g_125551_(out[357], out[533], _068372_);
  xor g_125552_(out[352], out[528], _068373_);
  or g_125553_(_068359_, _068365_, _068374_);
  or g_125554_(_068360_, _068362_, _068376_);
  or g_125555_(_068366_, _068371_, _068377_);
  or g_125556_(_068376_, _068377_, _068378_);
  or g_125557_(_068363_, _068368_, _068379_);
  or g_125558_(_068372_, _068373_, _068380_);
  or g_125559_(_068379_, _068380_, _068381_);
  or g_125560_(_068378_, _068381_, _068382_);
  xor g_125561_(out[364], out[540], _068383_);
  or g_125562_(_068358_, _068383_, _068384_);
  or g_125563_(_068357_, _068369_, _068385_);
  or g_125564_(_068384_, _068385_, _068387_);
  or g_125565_(_068361_, _068367_, _068388_);
  or g_125566_(_068370_, _068388_, _068389_);
  or g_125567_(_068387_, _068389_, _068390_);
  or g_125568_(_068382_, _068390_, _068391_);
  or g_125569_(_068374_, _068391_, _068392_);
  xor g_125570_(out[346], out[538], _068393_);
  xor g_125571_(out[338], out[530], _068394_);
  xor g_125572_(out[337], out[529], _068395_);
  and g_125573_(_049400_, out[539], _068396_);
  and g_125574_(out[347], _049532_, _068398_);
  xor g_125575_(out[349], out[541], _068399_);
  xor g_125576_(out[339], out[531], _068400_);
  xor g_125577_(out[350], out[542], _068401_);
  xor g_125578_(out[348], out[540], _068402_);
  xor g_125579_(out[344], out[536], _068403_);
  xor g_125580_(out[351], out[543], _068404_);
  xor g_125581_(out[341], out[533], _068405_);
  xor g_125582_(out[342], out[534], _068406_);
  xor g_125583_(out[336], out[528], _068407_);
  xor g_125584_(out[340], out[532], _068409_);
  or g_125585_(_068399_, _068403_, _068410_);
  xor g_125586_(out[345], out[537], _068411_);
  or g_125587_(_068393_, _068394_, _068412_);
  or g_125588_(_068410_, _068412_, _068413_);
  or g_125589_(_068400_, _068411_, _068414_);
  or g_125590_(_068405_, _068414_, _068415_);
  or g_125591_(_068413_, _068415_, _068416_);
  or g_125592_(_068401_, _068409_, _068417_);
  or g_125593_(_068416_, _068417_, _068418_);
  or g_125594_(_068396_, _068402_, _068420_);
  xor g_125595_(out[343], out[535], _068421_);
  or g_125596_(_068406_, _068421_, _068422_);
  or g_125597_(_068420_, _068422_, _068423_);
  or g_125598_(_068395_, _068398_, _068424_);
  or g_125599_(_068404_, _068424_, _068425_);
  or g_125600_(_068423_, _068425_, _068426_);
  or g_125601_(_068407_, _068426_, _068427_);
  or g_125602_(_068418_, _068427_, _068428_);
  xor g_125603_(out[327], out[535], _068429_);
  and g_125604_(_098294_, out[539], _068431_);
  xor g_125605_(out[334], out[542], _068432_);
  xor g_125606_(out[328], out[536], _068433_);
  xor g_125607_(out[321], out[529], _068434_);
  xor g_125608_(out[333], out[541], _068435_);
  xor g_125609_(out[329], out[537], _068436_);
  xor g_125610_(out[324], out[532], _068437_);
  xor g_125611_(out[322], out[530], _068438_);
  and g_125612_(out[331], _049532_, _068439_);
  xor g_125613_(out[323], out[531], _068440_);
  xor g_125614_(out[326], out[534], _068442_);
  xor g_125615_(out[335], out[543], _068443_);
  xor g_125616_(out[330], out[538], _068444_);
  xor g_125617_(out[325], out[533], _068445_);
  xor g_125618_(out[320], out[528], _068446_);
  or g_125619_(_068432_, _068437_, _068447_);
  or g_125620_(_068433_, _068435_, _068448_);
  or g_125621_(_068438_, _068444_, _068449_);
  or g_125622_(_068448_, _068449_, _068450_);
  or g_125623_(_068436_, _068440_, _068451_);
  or g_125624_(_068445_, _068446_, _068453_);
  or g_125625_(_068451_, _068453_, _068454_);
  or g_125626_(_068450_, _068454_, _068455_);
  xor g_125627_(out[332], out[540], _068456_);
  or g_125628_(_068431_, _068456_, _068457_);
  or g_125629_(_068429_, _068442_, _068458_);
  or g_125630_(_068457_, _068458_, _068459_);
  or g_125631_(_068434_, _068439_, _068460_);
  or g_125632_(_068443_, _068460_, _068461_);
  or g_125633_(_068459_, _068461_, _068462_);
  or g_125634_(_068455_, _068462_, _068464_);
  or g_125635_(_068447_, _068464_, _068465_);
  xor g_125636_(out[312], out[536], _068466_);
  xor g_125637_(out[309], out[533], _068467_);
  xor g_125638_(out[307], out[531], _068468_);
  xor g_125639_(out[318], out[542], _068469_);
  xor g_125640_(out[317], out[541], _068470_);
  xor g_125641_(out[306], out[530], _068471_);
  xor g_125642_(out[313], out[537], _068472_);
  xor g_125643_(out[310], out[534], _068473_);
  xor g_125644_(out[319], out[543], _068475_);
  xor g_125645_(out[314], out[538], _068476_);
  xor g_125646_(out[308], out[532], _068477_);
  xor g_125647_(out[304], out[528], _068478_);
  and g_125648_(_098283_, out[539], _068479_);
  and g_125649_(out[315], _049532_, _068480_);
  or g_125650_(_068466_, _068470_, _068481_);
  xor g_125651_(out[305], out[529], _068482_);
  or g_125652_(_068471_, _068476_, _068483_);
  or g_125653_(_068481_, _068483_, _068484_);
  or g_125654_(_068468_, _068472_, _068486_);
  or g_125655_(_068467_, _068486_, _068487_);
  or g_125656_(_068484_, _068487_, _068488_);
  or g_125657_(_068469_, _068477_, _068489_);
  or g_125658_(_068488_, _068489_, _068490_);
  xor g_125659_(out[316], out[540], _068491_);
  or g_125660_(_068479_, _068491_, _068492_);
  xor g_125661_(out[311], out[535], _068493_);
  or g_125662_(_068473_, _068493_, _068494_);
  or g_125663_(_068492_, _068494_, _068495_);
  or g_125664_(_068480_, _068482_, _068497_);
  or g_125665_(_068475_, _068497_, _068498_);
  or g_125666_(_068495_, _068498_, _068499_);
  or g_125667_(_068478_, _068499_, _068500_);
  or g_125668_(_068490_, _068500_, _068501_);
  xor g_125669_(out[295], out[535], _068502_);
  and g_125670_(_098272_, out[539], _068503_);
  xor g_125671_(out[302], out[542], _068504_);
  xor g_125672_(out[296], out[536], _068505_);
  xor g_125673_(out[289], out[529], _068506_);
  xor g_125674_(out[301], out[541], _068508_);
  xor g_125675_(out[297], out[537], _068509_);
  xor g_125676_(out[292], out[532], _068510_);
  xor g_125677_(out[290], out[530], _068511_);
  and g_125678_(out[299], _049532_, _068512_);
  xor g_125679_(out[291], out[531], _068513_);
  xor g_125680_(out[294], out[534], _068514_);
  xor g_125681_(out[303], out[543], _068515_);
  xor g_125682_(out[298], out[538], _068516_);
  xor g_125683_(out[293], out[533], _068517_);
  xor g_125684_(out[288], out[528], _068519_);
  or g_125685_(_068504_, _068510_, _068520_);
  or g_125686_(_068505_, _068508_, _068521_);
  or g_125687_(_068511_, _068516_, _068522_);
  or g_125688_(_068521_, _068522_, _068523_);
  or g_125689_(_068509_, _068513_, _068524_);
  or g_125690_(_068517_, _068519_, _068525_);
  or g_125691_(_068524_, _068525_, _068526_);
  or g_125692_(_068523_, _068526_, _068527_);
  xor g_125693_(out[300], out[540], _068528_);
  or g_125694_(_068503_, _068528_, _068530_);
  or g_125695_(_068502_, _068514_, _068531_);
  or g_125696_(_068530_, _068531_, _068532_);
  or g_125697_(_068506_, _068512_, _068533_);
  or g_125698_(_068515_, _068533_, _068534_);
  or g_125699_(_068532_, _068534_, _068535_);
  or g_125700_(_068527_, _068535_, _068536_);
  or g_125701_(_068520_, _068536_, _068537_);
  xor g_125702_(out[284], out[540], _068538_);
  and g_125703_(_098261_, out[539], _068539_);
  xor g_125704_(out[280], out[536], _068541_);
  xor g_125705_(out[278], out[534], _068542_);
  xor g_125706_(out[285], out[541], _068543_);
  xor g_125707_(out[286], out[542], _068544_);
  xor g_125708_(out[274], out[530], _068545_);
  xor g_125709_(out[281], out[537], _068546_);
  xor g_125710_(out[277], out[533], _068547_);
  xor g_125711_(out[273], out[529], _068548_);
  and g_125712_(out[283], _049532_, _068549_);
  or g_125713_(_068541_, _068543_, _068550_);
  xor g_125714_(out[287], out[543], _068552_);
  xor g_125715_(out[282], out[538], _068553_);
  xor g_125716_(out[276], out[532], _068554_);
  xor g_125717_(out[275], out[531], _068555_);
  xor g_125718_(out[272], out[528], _068556_);
  or g_125719_(_068545_, _068553_, _068557_);
  or g_125720_(_068550_, _068557_, _068558_);
  or g_125721_(_068546_, _068555_, _068559_);
  or g_125722_(_068547_, _068559_, _068560_);
  or g_125723_(_068558_, _068560_, _068561_);
  or g_125724_(_068544_, _068554_, _068563_);
  or g_125725_(_068561_, _068563_, _068564_);
  or g_125726_(_068538_, _068539_, _068565_);
  xor g_125727_(out[279], out[535], _068566_);
  or g_125728_(_068542_, _068566_, _068567_);
  or g_125729_(_068565_, _068567_, _068568_);
  or g_125730_(_068548_, _068549_, _068569_);
  or g_125731_(_068552_, _068569_, _068570_);
  or g_125732_(_068568_, _068570_, _068571_);
  or g_125733_(_068556_, _068571_, _068572_);
  or g_125734_(_068564_, _068572_, _068574_);
  xor g_125735_(out[263], out[535], _068575_);
  and g_125736_(_098250_, out[539], _068576_);
  xor g_125737_(out[270], out[542], _068577_);
  xor g_125738_(out[264], out[536], _068578_);
  xor g_125739_(out[257], out[529], _068579_);
  xor g_125740_(out[269], out[541], _068580_);
  xor g_125741_(out[265], out[537], _068581_);
  xor g_125742_(out[260], out[532], _068582_);
  xor g_125743_(out[258], out[530], _068583_);
  and g_125744_(out[267], _049532_, _068585_);
  xor g_125745_(out[259], out[531], _068586_);
  xor g_125746_(out[262], out[534], _068587_);
  xor g_125747_(out[271], out[543], _068588_);
  xor g_125748_(out[266], out[538], _068589_);
  xor g_125749_(out[261], out[533], _068590_);
  xor g_125750_(out[256], out[528], _068591_);
  or g_125751_(_068577_, _068582_, _068592_);
  or g_125752_(_068578_, _068580_, _068593_);
  or g_125753_(_068583_, _068589_, _068594_);
  or g_125754_(_068593_, _068594_, _068596_);
  or g_125755_(_068581_, _068586_, _068597_);
  or g_125756_(_068590_, _068591_, _068598_);
  or g_125757_(_068597_, _068598_, _068599_);
  or g_125758_(_068596_, _068599_, _068600_);
  xor g_125759_(out[268], out[540], _068601_);
  or g_125760_(_068576_, _068601_, _068602_);
  or g_125761_(_068575_, _068587_, _068603_);
  or g_125762_(_068602_, _068603_, _068604_);
  or g_125763_(_068579_, _068585_, _068605_);
  or g_125764_(_068588_, _068605_, _068607_);
  or g_125765_(_068604_, _068607_, _068608_);
  or g_125766_(_068600_, _068608_, _068609_);
  or g_125767_(_068592_, _068609_, _068610_);
  not g_125768_(_068610_, _068611_);
  xor g_125769_(out[248], out[536], _068612_);
  xor g_125770_(out[245], out[533], _068613_);
  xor g_125771_(out[243], out[531], _068614_);
  xor g_125772_(out[254], out[542], _068615_);
  xor g_125773_(out[253], out[541], _068616_);
  xor g_125774_(out[242], out[530], _068618_);
  xor g_125775_(out[249], out[537], _068619_);
  xor g_125776_(out[246], out[534], _068620_);
  xor g_125777_(out[255], out[543], _068621_);
  xor g_125778_(out[250], out[538], _068622_);
  xor g_125779_(out[244], out[532], _068623_);
  xor g_125780_(out[240], out[528], _068624_);
  and g_125781_(_098239_, out[539], _068625_);
  and g_125782_(out[251], _049532_, _068626_);
  or g_125783_(_068612_, _068616_, _068627_);
  xor g_125784_(out[241], out[529], _068629_);
  or g_125785_(_068618_, _068622_, _068630_);
  or g_125786_(_068627_, _068630_, _068631_);
  or g_125787_(_068614_, _068619_, _068632_);
  or g_125788_(_068613_, _068632_, _068633_);
  or g_125789_(_068631_, _068633_, _068634_);
  or g_125790_(_068615_, _068623_, _068635_);
  or g_125791_(_068634_, _068635_, _068636_);
  xor g_125792_(out[252], out[540], _068637_);
  or g_125793_(_068625_, _068637_, _068638_);
  xor g_125794_(out[247], out[535], _068640_);
  or g_125795_(_068620_, _068640_, _068641_);
  or g_125796_(_068638_, _068641_, _068642_);
  or g_125797_(_068626_, _068629_, _068643_);
  or g_125798_(_068621_, _068643_, _068644_);
  or g_125799_(_068642_, _068644_, _068645_);
  or g_125800_(_068624_, _068645_, _068646_);
  or g_125801_(_068636_, _068646_, _068647_);
  not g_125802_(_068647_, _068648_);
  xor g_125803_(out[231], out[535], _068649_);
  and g_125804_(_098228_, out[539], _068651_);
  xor g_125805_(out[238], out[542], _068652_);
  xor g_125806_(out[232], out[536], _068653_);
  xor g_125807_(out[225], out[529], _068654_);
  xor g_125808_(out[237], out[541], _068655_);
  xor g_125809_(out[233], out[537], _068656_);
  xor g_125810_(out[228], out[532], _068657_);
  xor g_125811_(out[226], out[530], _068658_);
  and g_125812_(out[235], _049532_, _068659_);
  xor g_125813_(out[227], out[531], _068660_);
  xor g_125814_(out[230], out[534], _068662_);
  xor g_125815_(out[239], out[543], _068663_);
  xor g_125816_(out[234], out[538], _068664_);
  xor g_125817_(out[229], out[533], _068665_);
  xor g_125818_(out[224], out[528], _068666_);
  or g_125819_(_068652_, _068657_, _068667_);
  or g_125820_(_068653_, _068655_, _068668_);
  or g_125821_(_068658_, _068664_, _068669_);
  or g_125822_(_068668_, _068669_, _068670_);
  or g_125823_(_068656_, _068660_, _068671_);
  or g_125824_(_068665_, _068666_, _068673_);
  or g_125825_(_068671_, _068673_, _068674_);
  or g_125826_(_068670_, _068674_, _068675_);
  xor g_125827_(out[236], out[540], _068676_);
  or g_125828_(_068651_, _068676_, _068677_);
  or g_125829_(_068649_, _068662_, _068678_);
  or g_125830_(_068677_, _068678_, _068679_);
  or g_125831_(_068654_, _068659_, _068680_);
  or g_125832_(_068663_, _068680_, _068681_);
  or g_125833_(_068679_, _068681_, _068682_);
  or g_125834_(_068675_, _068682_, _068684_);
  or g_125835_(_068667_, _068684_, _068685_);
  xor g_125836_(out[212], out[532], _068686_);
  xor g_125837_(out[220], out[540], _068687_);
  and g_125838_(_098217_, out[539], _068688_);
  xor g_125839_(out[218], out[538], _068689_);
  xor g_125840_(out[214], out[534], _068690_);
  xor g_125841_(out[213], out[533], _068691_);
  xor g_125842_(out[211], out[531], _068692_);
  xor g_125843_(out[221], out[541], _068693_);
  xor g_125844_(out[222], out[542], _068695_);
  xor g_125845_(out[209], out[529], _068696_);
  xor g_125846_(out[210], out[530], _068697_);
  and g_125847_(out[219], _049532_, _068698_);
  xor g_125848_(out[208], out[528], _068699_);
  xor g_125849_(out[223], out[543], _068700_);
  xor g_125850_(out[216], out[536], _068701_);
  or g_125851_(_068693_, _068701_, _068702_);
  xor g_125852_(out[217], out[537], _068703_);
  or g_125853_(_068689_, _068697_, _068704_);
  or g_125854_(_068702_, _068704_, _068706_);
  or g_125855_(_068692_, _068703_, _068707_);
  or g_125856_(_068691_, _068707_, _068708_);
  or g_125857_(_068706_, _068708_, _068709_);
  or g_125858_(_068686_, _068695_, _068710_);
  or g_125859_(_068709_, _068710_, _068711_);
  or g_125860_(_068687_, _068688_, _068712_);
  xor g_125861_(out[215], out[535], _068713_);
  or g_125862_(_068690_, _068713_, _068714_);
  or g_125863_(_068712_, _068714_, _068715_);
  or g_125864_(_068696_, _068698_, _068717_);
  or g_125865_(_068700_, _068717_, _068718_);
  or g_125866_(_068715_, _068718_, _068719_);
  or g_125867_(_068699_, _068719_, _068720_);
  or g_125868_(_068711_, _068720_, _068721_);
  xor g_125869_(out[199], out[535], _068722_);
  and g_125870_(_098206_, out[539], _068723_);
  xor g_125871_(out[206], out[542], _068724_);
  xor g_125872_(out[200], out[536], _068725_);
  xor g_125873_(out[193], out[529], _068726_);
  xor g_125874_(out[205], out[541], _068728_);
  xor g_125875_(out[201], out[537], _068729_);
  xor g_125876_(out[196], out[532], _068730_);
  xor g_125877_(out[194], out[530], _068731_);
  and g_125878_(out[203], _049532_, _068732_);
  xor g_125879_(out[195], out[531], _068733_);
  xor g_125880_(out[198], out[534], _068734_);
  xor g_125881_(out[207], out[543], _068735_);
  xor g_125882_(out[202], out[538], _068736_);
  xor g_125883_(out[197], out[533], _068737_);
  xor g_125884_(out[192], out[528], _068739_);
  or g_125885_(_068724_, _068730_, _068740_);
  or g_125886_(_068725_, _068728_, _068741_);
  or g_125887_(_068731_, _068736_, _068742_);
  or g_125888_(_068741_, _068742_, _068743_);
  or g_125889_(_068729_, _068733_, _068744_);
  or g_125890_(_068737_, _068739_, _068745_);
  or g_125891_(_068744_, _068745_, _068746_);
  or g_125892_(_068743_, _068746_, _068747_);
  xor g_125893_(out[204], out[540], _068748_);
  or g_125894_(_068723_, _068748_, _068750_);
  or g_125895_(_068722_, _068734_, _068751_);
  or g_125896_(_068750_, _068751_, _068752_);
  or g_125897_(_068726_, _068732_, _068753_);
  or g_125898_(_068735_, _068753_, _068754_);
  or g_125899_(_068752_, _068754_, _068755_);
  or g_125900_(_068747_, _068755_, _068756_);
  or g_125901_(_068740_, _068756_, _068757_);
  xor g_125902_(out[179], out[531], _068758_);
  xor g_125903_(out[180], out[532], _068759_);
  xor g_125904_(out[190], out[542], _068761_);
  xor g_125905_(out[178], out[530], _068762_);
  xor g_125906_(out[181], out[533], _068763_);
  xor g_125907_(out[185], out[537], _068764_);
  xor g_125908_(out[184], out[536], _068765_);
  xor g_125909_(out[191], out[543], _068766_);
  xor g_125910_(out[186], out[538], _068767_);
  xor g_125911_(out[182], out[534], _068768_);
  xor g_125912_(out[176], out[528], _068769_);
  and g_125913_(_098195_, out[539], _068770_);
  and g_125914_(out[187], _049532_, _068772_);
  xor g_125915_(out[189], out[541], _068773_);
  or g_125916_(_068765_, _068773_, _068774_);
  xor g_125917_(out[177], out[529], _068775_);
  or g_125918_(_068762_, _068767_, _068776_);
  or g_125919_(_068774_, _068776_, _068777_);
  or g_125920_(_068758_, _068764_, _068778_);
  or g_125921_(_068763_, _068778_, _068779_);
  or g_125922_(_068777_, _068779_, _068780_);
  or g_125923_(_068759_, _068761_, _068781_);
  or g_125924_(_068780_, _068781_, _068783_);
  xor g_125925_(out[188], out[540], _068784_);
  or g_125926_(_068770_, _068784_, _068785_);
  xor g_125927_(out[183], out[535], _068786_);
  or g_125928_(_068768_, _068786_, _068787_);
  or g_125929_(_068785_, _068787_, _068788_);
  or g_125930_(_068772_, _068775_, _068789_);
  or g_125931_(_068766_, _068789_, _068790_);
  or g_125932_(_068788_, _068790_, _068791_);
  or g_125933_(_068769_, _068791_, _068792_);
  or g_125934_(_068783_, _068792_, _068794_);
  xor g_125935_(out[167], out[535], _068795_);
  and g_125936_(_098184_, out[539], _068796_);
  xor g_125937_(out[174], out[542], _068797_);
  xor g_125938_(out[168], out[536], _068798_);
  xor g_125939_(out[161], out[529], _068799_);
  xor g_125940_(out[173], out[541], _068800_);
  xor g_125941_(out[169], out[537], _068801_);
  xor g_125942_(out[164], out[532], _068802_);
  xor g_125943_(out[162], out[530], _068803_);
  and g_125944_(out[171], _049532_, _068805_);
  xor g_125945_(out[163], out[531], _068806_);
  xor g_125946_(out[166], out[534], _068807_);
  xor g_125947_(out[175], out[543], _068808_);
  xor g_125948_(out[170], out[538], _068809_);
  xor g_125949_(out[165], out[533], _068810_);
  xor g_125950_(out[160], out[528], _068811_);
  or g_125951_(_068797_, _068802_, _068812_);
  or g_125952_(_068798_, _068800_, _068813_);
  or g_125953_(_068803_, _068809_, _068814_);
  or g_125954_(_068813_, _068814_, _068816_);
  or g_125955_(_068801_, _068806_, _068817_);
  or g_125956_(_068810_, _068811_, _068818_);
  or g_125957_(_068817_, _068818_, _068819_);
  or g_125958_(_068816_, _068819_, _068820_);
  xor g_125959_(out[172], out[540], _068821_);
  or g_125960_(_068796_, _068821_, _068822_);
  or g_125961_(_068795_, _068807_, _068823_);
  or g_125962_(_068822_, _068823_, _068824_);
  or g_125963_(_068799_, _068805_, _068825_);
  or g_125964_(_068808_, _068825_, _068827_);
  or g_125965_(_068824_, _068827_, _068828_);
  or g_125966_(_068820_, _068828_, _068829_);
  or g_125967_(_068812_, _068829_, _068830_);
  not g_125968_(_068830_, _068831_);
  and g_125969_(_098173_, out[539], _068832_);
  xor g_125970_(out[154], out[538], _068833_);
  xor g_125971_(out[159], out[543], _068834_);
  xor g_125972_(out[144], out[528], _068835_);
  xor g_125973_(out[148], out[532], _068836_);
  xor g_125974_(out[146], out[530], _068838_);
  xor g_125975_(out[153], out[537], _068839_);
  xor g_125976_(out[149], out[533], _068840_);
  xor g_125977_(out[145], out[529], _068841_);
  xor g_125978_(out[152], out[536], _068842_);
  and g_125979_(out[155], _049532_, _068843_);
  xor g_125980_(out[150], out[534], _068844_);
  xor g_125981_(out[147], out[531], _068845_);
  xor g_125982_(out[157], out[541], _068846_);
  xor g_125983_(out[158], out[542], _068847_);
  or g_125984_(_068836_, _068847_, _068849_);
  or g_125985_(_068842_, _068846_, _068850_);
  or g_125986_(_068833_, _068838_, _068851_);
  or g_125987_(_068850_, _068851_, _068852_);
  or g_125988_(_068839_, _068845_, _068853_);
  or g_125989_(_068835_, _068840_, _068854_);
  or g_125990_(_068853_, _068854_, _068855_);
  or g_125991_(_068852_, _068855_, _068856_);
  xor g_125992_(out[156], out[540], _068857_);
  or g_125993_(_068832_, _068857_, _068858_);
  xor g_125994_(out[151], out[535], _068860_);
  or g_125995_(_068844_, _068860_, _068861_);
  or g_125996_(_068858_, _068861_, _068862_);
  or g_125997_(_068841_, _068843_, _068863_);
  or g_125998_(_068834_, _068863_, _068864_);
  or g_125999_(_068862_, _068864_, _068865_);
  or g_126000_(_068856_, _068865_, _068866_);
  or g_126001_(_068849_, _068866_, _068867_);
  xor g_126002_(out[135], out[535], _068868_);
  and g_126003_(_098162_, out[539], _068869_);
  xor g_126004_(out[142], out[542], _068871_);
  xor g_126005_(out[136], out[536], _068872_);
  xor g_126006_(out[129], out[529], _068873_);
  xor g_126007_(out[141], out[541], _068874_);
  xor g_126008_(out[137], out[537], _068875_);
  xor g_126009_(out[132], out[532], _068876_);
  xor g_126010_(out[130], out[530], _068877_);
  and g_126011_(out[139], _049532_, _068878_);
  xor g_126012_(out[131], out[531], _068879_);
  xor g_126013_(out[134], out[534], _068880_);
  xor g_126014_(out[143], out[543], _068882_);
  xor g_126015_(out[138], out[538], _068883_);
  xor g_126016_(out[133], out[533], _068884_);
  xor g_126017_(out[128], out[528], _068885_);
  or g_126018_(_068871_, _068876_, _068886_);
  or g_126019_(_068872_, _068874_, _068887_);
  or g_126020_(_068877_, _068883_, _068888_);
  or g_126021_(_068887_, _068888_, _068889_);
  or g_126022_(_068875_, _068879_, _068890_);
  or g_126023_(_068884_, _068885_, _068891_);
  or g_126024_(_068890_, _068891_, _068893_);
  or g_126025_(_068889_, _068893_, _068894_);
  xor g_126026_(out[140], out[540], _068895_);
  or g_126027_(_068869_, _068895_, _068896_);
  or g_126028_(_068868_, _068880_, _068897_);
  or g_126029_(_068896_, _068897_, _068898_);
  or g_126030_(_068873_, _068878_, _068899_);
  or g_126031_(_068882_, _068899_, _068900_);
  or g_126032_(_068898_, _068900_, _068901_);
  or g_126033_(_068894_, _068901_, _068902_);
  or g_126034_(_068886_, _068902_, _068904_);
  xor g_126035_(out[114], out[530], _068905_);
  xor g_126036_(out[112], out[528], _068906_);
  xor g_126037_(out[121], out[537], _068907_);
  xor g_126038_(out[120], out[536], _068908_);
  xor g_126039_(out[117], out[533], _068909_);
  xor g_126040_(out[126], out[542], _068910_);
  xor g_126041_(out[125], out[541], _068911_);
  xor g_126042_(out[127], out[543], _068912_);
  xor g_126043_(out[122], out[538], _068913_);
  xor g_126044_(out[118], out[534], _068915_);
  xor g_126045_(out[115], out[531], _068916_);
  and g_126046_(_098151_, out[539], _068917_);
  and g_126047_(out[123], _049532_, _068918_);
  xor g_126048_(out[116], out[532], _068919_);
  xor g_126049_(out[113], out[529], _068920_);
  or g_126050_(_068910_, _068919_, _068921_);
  or g_126051_(_068908_, _068911_, _068922_);
  or g_126052_(_068905_, _068913_, _068923_);
  or g_126053_(_068922_, _068923_, _068924_);
  or g_126054_(_068907_, _068916_, _068926_);
  or g_126055_(_068906_, _068909_, _068927_);
  or g_126056_(_068926_, _068927_, _068928_);
  or g_126057_(_068924_, _068928_, _068929_);
  xor g_126058_(out[124], out[540], _068930_);
  or g_126059_(_068917_, _068930_, _068931_);
  xor g_126060_(out[119], out[535], _068932_);
  or g_126061_(_068915_, _068932_, _068933_);
  or g_126062_(_068931_, _068933_, _068934_);
  or g_126063_(_068918_, _068920_, _068935_);
  or g_126064_(_068912_, _068935_, _068937_);
  or g_126065_(_068934_, _068937_, _068938_);
  or g_126066_(_068929_, _068938_, _068939_);
  or g_126067_(_068921_, _068939_, _068940_);
  not g_126068_(_068940_, _068941_);
  xor g_126069_(out[103], out[535], _068942_);
  and g_126070_(_098140_, out[539], _068943_);
  xor g_126071_(out[110], out[542], _068944_);
  xor g_126072_(out[104], out[536], _068945_);
  xor g_126073_(out[97], out[529], _068946_);
  xor g_126074_(out[109], out[541], _068948_);
  xor g_126075_(out[105], out[537], _068949_);
  xor g_126076_(out[100], out[532], _068950_);
  xor g_126077_(out[98], out[530], _068951_);
  and g_126078_(out[107], _049532_, _068952_);
  xor g_126079_(out[99], out[531], _068953_);
  xor g_126080_(out[102], out[534], _068954_);
  xor g_126081_(out[111], out[543], _068955_);
  xor g_126082_(out[106], out[538], _068956_);
  xor g_126083_(out[101], out[533], _068957_);
  xor g_126084_(out[96], out[528], _068959_);
  or g_126085_(_068944_, _068950_, _068960_);
  or g_126086_(_068945_, _068948_, _068961_);
  or g_126087_(_068951_, _068956_, _068962_);
  or g_126088_(_068961_, _068962_, _068963_);
  or g_126089_(_068949_, _068953_, _068964_);
  or g_126090_(_068957_, _068959_, _068965_);
  or g_126091_(_068964_, _068965_, _068966_);
  or g_126092_(_068963_, _068966_, _068967_);
  xor g_126093_(out[108], out[540], _068968_);
  or g_126094_(_068943_, _068968_, _068970_);
  or g_126095_(_068942_, _068954_, _068971_);
  or g_126096_(_068970_, _068971_, _068972_);
  or g_126097_(_068946_, _068952_, _068973_);
  or g_126098_(_068955_, _068973_, _068974_);
  or g_126099_(_068972_, _068974_, _068975_);
  or g_126100_(_068967_, _068975_, _068976_);
  or g_126101_(_068960_, _068976_, _068977_);
  not g_126102_(_068977_, _068978_);
  xor g_126103_(out[92], out[540], _068979_);
  and g_126104_(_098129_, out[539], _068981_);
  xor g_126105_(out[88], out[536], _068982_);
  xor g_126106_(out[86], out[534], _068983_);
  xor g_126107_(out[93], out[541], _068984_);
  xor g_126108_(out[94], out[542], _068985_);
  xor g_126109_(out[82], out[530], _068986_);
  xor g_126110_(out[89], out[537], _068987_);
  xor g_126111_(out[85], out[533], _068988_);
  xor g_126112_(out[81], out[529], _068989_);
  and g_126113_(out[91], _049532_, _068990_);
  or g_126114_(_068982_, _068984_, _068992_);
  xor g_126115_(out[95], out[543], _068993_);
  xor g_126116_(out[90], out[538], _068994_);
  xor g_126117_(out[84], out[532], _068995_);
  xor g_126118_(out[83], out[531], _068996_);
  xor g_126119_(out[80], out[528], _068997_);
  or g_126120_(_068986_, _068994_, _068998_);
  or g_126121_(_068992_, _068998_, _068999_);
  or g_126122_(_068987_, _068996_, _069000_);
  or g_126123_(_068988_, _069000_, _069001_);
  or g_126124_(_068999_, _069001_, _069003_);
  or g_126125_(_068985_, _068995_, _069004_);
  or g_126126_(_069003_, _069004_, _069005_);
  or g_126127_(_068979_, _068981_, _069006_);
  xor g_126128_(out[87], out[535], _069007_);
  or g_126129_(_068983_, _069007_, _069008_);
  or g_126130_(_069006_, _069008_, _069009_);
  or g_126131_(_068989_, _068990_, _069010_);
  or g_126132_(_068993_, _069010_, _069011_);
  or g_126133_(_069009_, _069011_, _069012_);
  or g_126134_(_068997_, _069012_, _069014_);
  or g_126135_(_069005_, _069014_, _069015_);
  not g_126136_(_069015_, _069016_);
  xor g_126137_(out[71], out[535], _069017_);
  and g_126138_(_098118_, out[539], _069018_);
  xor g_126139_(out[78], out[542], _069019_);
  xor g_126140_(out[72], out[536], _069020_);
  xor g_126141_(out[65], out[529], _069021_);
  xor g_126142_(out[77], out[541], _069022_);
  xor g_126143_(out[73], out[537], _069023_);
  xor g_126144_(out[68], out[532], _069025_);
  xor g_126145_(out[66], out[530], _069026_);
  and g_126146_(out[75], _049532_, _069027_);
  xor g_126147_(out[67], out[531], _069028_);
  xor g_126148_(out[70], out[534], _069029_);
  xor g_126149_(out[79], out[543], _069030_);
  xor g_126150_(out[74], out[538], _069031_);
  xor g_126151_(out[69], out[533], _069032_);
  xor g_126152_(out[64], out[528], _069033_);
  or g_126153_(_069019_, _069025_, _069034_);
  or g_126154_(_069020_, _069022_, _069036_);
  or g_126155_(_069026_, _069031_, _069037_);
  or g_126156_(_069036_, _069037_, _069038_);
  or g_126157_(_069023_, _069028_, _069039_);
  or g_126158_(_069032_, _069033_, _069040_);
  or g_126159_(_069039_, _069040_, _069041_);
  or g_126160_(_069038_, _069041_, _069042_);
  xor g_126161_(out[76], out[540], _069043_);
  or g_126162_(_069018_, _069043_, _069044_);
  or g_126163_(_069017_, _069029_, _069045_);
  or g_126164_(_069044_, _069045_, _069047_);
  or g_126165_(_069021_, _069027_, _069048_);
  or g_126166_(_069030_, _069048_, _069049_);
  or g_126167_(_069047_, _069049_, _069050_);
  or g_126168_(_069042_, _069050_, _069051_);
  or g_126169_(_069034_, _069051_, _069052_);
  not g_126170_(_069052_, _069053_);
  xor g_126171_(out[49], out[529], _069054_);
  and g_126172_(out[59], _049532_, _069055_);
  xor g_126173_(out[57], out[537], _069056_);
  xor g_126174_(out[48], out[528], _069058_);
  xor g_126175_(out[62], out[542], _069059_);
  xor g_126176_(out[52], out[532], _069060_);
  or g_126177_(_069059_, _069060_, _069061_);
  xor g_126178_(out[61], out[541], _069062_);
  xor g_126179_(out[51], out[531], _069063_);
  and g_126180_(_098107_, out[539], _069064_);
  xor g_126181_(out[54], out[534], _069065_);
  xor g_126182_(out[58], out[538], _069066_);
  xor g_126183_(out[53], out[533], _069067_);
  xor g_126184_(out[63], out[543], _069069_);
  xor g_126185_(out[56], out[536], _069070_);
  or g_126186_(_069062_, _069070_, _069071_);
  xor g_126187_(out[50], out[530], _069072_);
  or g_126188_(_069066_, _069072_, _069073_);
  or g_126189_(_069071_, _069073_, _069074_);
  or g_126190_(_069056_, _069063_, _069075_);
  or g_126191_(_069067_, _069075_, _069076_);
  or g_126192_(_069074_, _069076_, _069077_);
  or g_126193_(_069061_, _069077_, _069078_);
  xor g_126194_(out[60], out[540], _069080_);
  or g_126195_(_069064_, _069080_, _069081_);
  xor g_126196_(out[55], out[535], _069082_);
  or g_126197_(_069065_, _069082_, _069083_);
  or g_126198_(_069081_, _069083_, _069084_);
  or g_126199_(_069054_, _069055_, _069085_);
  or g_126200_(_069069_, _069085_, _069086_);
  or g_126201_(_069084_, _069086_, _069087_);
  or g_126202_(_069058_, _069087_, _069088_);
  or g_126203_(_069078_, _069088_, _069089_);
  xor g_126204_(out[39], out[535], _069091_);
  and g_126205_(_098096_, out[539], _069092_);
  xor g_126206_(out[46], out[542], _069093_);
  xor g_126207_(out[40], out[536], _069094_);
  xor g_126208_(out[33], out[529], _069095_);
  xor g_126209_(out[45], out[541], _069096_);
  xor g_126210_(out[41], out[537], _069097_);
  xor g_126211_(out[36], out[532], _069098_);
  xor g_126212_(out[34], out[530], _069099_);
  and g_126213_(out[43], _049532_, _069100_);
  xor g_126214_(out[35], out[531], _069102_);
  xor g_126215_(out[38], out[534], _069103_);
  xor g_126216_(out[47], out[543], _069104_);
  xor g_126217_(out[42], out[538], _069105_);
  xor g_126218_(out[37], out[533], _069106_);
  xor g_126219_(out[32], out[528], _069107_);
  or g_126220_(_069093_, _069098_, _069108_);
  or g_126221_(_069094_, _069096_, _069109_);
  or g_126222_(_069099_, _069105_, _069110_);
  or g_126223_(_069109_, _069110_, _069111_);
  or g_126224_(_069097_, _069102_, _069113_);
  or g_126225_(_069106_, _069107_, _069114_);
  or g_126226_(_069113_, _069114_, _069115_);
  or g_126227_(_069111_, _069115_, _069116_);
  xor g_126228_(out[44], out[540], _069117_);
  or g_126229_(_069092_, _069117_, _069118_);
  or g_126230_(_069091_, _069103_, _069119_);
  or g_126231_(_069118_, _069119_, _069120_);
  or g_126232_(_069095_, _069100_, _069121_);
  or g_126233_(_069104_, _069121_, _069122_);
  or g_126234_(_069120_, _069122_, _069124_);
  or g_126235_(_069116_, _069124_, _069125_);
  or g_126236_(_069108_, _069125_, _069126_);
  and g_126237_(out[27], _049532_, _069127_);
  xor g_126238_(out[20], out[532], _069128_);
  xor g_126239_(out[30], out[542], _069129_);
  or g_126240_(_069128_, _069129_, _069130_);
  xor g_126241_(out[29], out[541], _069131_);
  xor g_126242_(out[19], out[531], _069132_);
  xor g_126243_(out[16], out[528], _069133_);
  and g_126244_(_098063_, out[539], _069135_);
  xor g_126245_(out[26], out[538], _069136_);
  xor g_126246_(out[31], out[543], _069137_);
  xor g_126247_(out[22], out[534], _069138_);
  xor g_126248_(out[21], out[533], _069139_);
  xor g_126249_(out[24], out[536], _069140_);
  or g_126250_(_069131_, _069140_, _069141_);
  xor g_126251_(out[18], out[530], _069142_);
  xor g_126252_(out[25], out[537], _069143_);
  xor g_126253_(out[17], out[529], _069144_);
  or g_126254_(_069136_, _069142_, _069146_);
  or g_126255_(_069141_, _069146_, _069147_);
  or g_126256_(_069132_, _069143_, _069148_);
  or g_126257_(_069139_, _069148_, _069149_);
  or g_126258_(_069147_, _069149_, _069150_);
  or g_126259_(_069130_, _069150_, _069151_);
  xor g_126260_(out[28], out[540], _069152_);
  or g_126261_(_069135_, _069152_, _069153_);
  xor g_126262_(out[23], out[535], _069154_);
  or g_126263_(_069138_, _069154_, _069155_);
  or g_126264_(_069153_, _069155_, _069157_);
  or g_126265_(_069127_, _069144_, _069158_);
  or g_126266_(_069137_, _069158_, _069159_);
  or g_126267_(_069157_, _069159_, _069160_);
  or g_126268_(_069133_, _069160_, _069161_);
  or g_126269_(_069151_, _069161_, _069162_);
  not g_126270_(_069162_, _069163_);
  xor g_126271_(out[1], out[529], _069164_);
  and g_126272_(out[11], _049532_, _069165_);
  xor g_126273_(out[14], out[542], _069166_);
  xor g_126274_(out[3], out[531], _069168_);
  xor g_126275_(out[4], out[532], _069169_);
  xor g_126276_(out[2], out[530], _069170_);
  xor g_126277_(out[9], out[537], _069171_);
  xor g_126278_(out[0], out[528], _069172_);
  and g_126279_(_098041_, out[539], _069173_);
  xor g_126280_(out[6], out[534], _069174_);
  xor g_126281_(out[10], out[538], _069175_);
  xor g_126282_(out[5], out[533], _069176_);
  xor g_126283_(out[15], out[543], _069177_);
  xor g_126284_(out[13], out[541], _069179_);
  xor g_126285_(out[8], out[536], _069180_);
  or g_126286_(_069166_, _069169_, _069181_);
  or g_126287_(_069179_, _069180_, _069182_);
  or g_126288_(_069170_, _069175_, _069183_);
  or g_126289_(_069182_, _069183_, _069184_);
  or g_126290_(_069168_, _069171_, _069185_);
  or g_126291_(_069172_, _069176_, _069186_);
  or g_126292_(_069185_, _069186_, _069187_);
  or g_126293_(_069184_, _069187_, _069188_);
  xor g_126294_(out[12], out[540], _069190_);
  or g_126295_(_069173_, _069190_, _069191_);
  xor g_126296_(out[7], out[535], _069192_);
  or g_126297_(_069174_, _069192_, _069193_);
  or g_126298_(_069191_, _069193_, _069194_);
  or g_126299_(_069164_, _069165_, _069195_);
  or g_126300_(_069177_, _069195_, _069196_);
  or g_126301_(_069194_, _069196_, _069197_);
  or g_126302_(_069188_, _069197_, _069198_);
  or g_126303_(_069181_, _069198_, _069199_);
  xor g_126304_(out[471], out[519], _069201_);
  and g_126305_(_049499_, out[523], _069202_);
  xor g_126306_(out[478], out[526], _069203_);
  xor g_126307_(out[472], out[520], _069204_);
  xor g_126308_(out[465], out[513], _069205_);
  xor g_126309_(out[477], out[525], _069206_);
  xor g_126310_(out[473], out[521], _069207_);
  xor g_126311_(out[468], out[516], _069208_);
  xor g_126312_(out[466], out[514], _069209_);
  and g_126313_(out[475], _049521_, _069210_);
  xor g_126314_(out[467], out[515], _069212_);
  xor g_126315_(out[470], out[518], _069213_);
  xor g_126316_(out[479], out[527], _069214_);
  xor g_126317_(out[474], out[522], _069215_);
  xor g_126318_(out[469], out[517], _069216_);
  xor g_126319_(out[464], out[512], _069217_);
  or g_126320_(_069203_, _069208_, _069218_);
  or g_126321_(_069204_, _069206_, _069219_);
  or g_126322_(_069209_, _069215_, _069220_);
  or g_126323_(_069219_, _069220_, _069221_);
  or g_126324_(_069207_, _069212_, _069223_);
  or g_126325_(_069216_, _069217_, _069224_);
  or g_126326_(_069223_, _069224_, _069225_);
  or g_126327_(_069221_, _069225_, _069226_);
  xor g_126328_(out[476], out[524], _069227_);
  or g_126329_(_069202_, _069227_, _069228_);
  or g_126330_(_069201_, _069213_, _069229_);
  or g_126331_(_069228_, _069229_, _069230_);
  or g_126332_(_069205_, _069210_, _069231_);
  or g_126333_(_069214_, _069231_, _069232_);
  or g_126334_(_069230_, _069232_, _069234_);
  or g_126335_(_069226_, _069234_, _069235_);
  or g_126336_(_069218_, _069235_, _069236_);
  xor g_126337_(out[458], out[522], _069237_);
  xor g_126338_(out[450], out[514], _069238_);
  xor g_126339_(out[449], out[513], _069239_);
  and g_126340_(_049477_, out[523], _069240_);
  and g_126341_(out[459], _049521_, _069241_);
  xor g_126342_(out[461], out[525], _069242_);
  xor g_126343_(out[451], out[515], _069243_);
  xor g_126344_(out[462], out[526], _069245_);
  xor g_126345_(out[460], out[524], _069246_);
  xor g_126346_(out[456], out[520], _069247_);
  xor g_126347_(out[463], out[527], _069248_);
  xor g_126348_(out[453], out[517], _069249_);
  xor g_126349_(out[454], out[518], _069250_);
  xor g_126350_(out[448], out[512], _069251_);
  xor g_126351_(out[452], out[516], _069252_);
  or g_126352_(_069242_, _069247_, _069253_);
  xor g_126353_(out[457], out[521], _069254_);
  or g_126354_(_069237_, _069238_, _069256_);
  or g_126355_(_069253_, _069256_, _069257_);
  or g_126356_(_069243_, _069254_, _069258_);
  or g_126357_(_069249_, _069258_, _069259_);
  or g_126358_(_069257_, _069259_, _069260_);
  or g_126359_(_069245_, _069252_, _069261_);
  or g_126360_(_069260_, _069261_, _069262_);
  or g_126361_(_069240_, _069246_, _069263_);
  xor g_126362_(out[455], out[519], _069264_);
  or g_126363_(_069250_, _069264_, _069265_);
  or g_126364_(_069263_, _069265_, _069267_);
  or g_126365_(_069239_, _069241_, _069268_);
  or g_126366_(_069248_, _069268_, _069269_);
  or g_126367_(_069267_, _069269_, _069270_);
  or g_126368_(_069251_, _069270_, _069271_);
  or g_126369_(_069262_, _069271_, _069272_);
  not g_126370_(_069272_, _069273_);
  xor g_126371_(out[439], out[519], _069274_);
  and g_126372_(_049466_, out[523], _069275_);
  xor g_126373_(out[446], out[526], _069276_);
  xor g_126374_(out[440], out[520], _069278_);
  xor g_126375_(out[433], out[513], _069279_);
  xor g_126376_(out[445], out[525], _069280_);
  xor g_126377_(out[441], out[521], _069281_);
  xor g_126378_(out[436], out[516], _069282_);
  xor g_126379_(out[434], out[514], _069283_);
  and g_126380_(out[443], _049521_, _069284_);
  xor g_126381_(out[435], out[515], _069285_);
  xor g_126382_(out[438], out[518], _069286_);
  xor g_126383_(out[447], out[527], _069287_);
  xor g_126384_(out[442], out[522], _069289_);
  xor g_126385_(out[437], out[517], _069290_);
  xor g_126386_(out[432], out[512], _069291_);
  or g_126387_(_069276_, _069282_, _069292_);
  or g_126388_(_069278_, _069280_, _069293_);
  or g_126389_(_069283_, _069289_, _069294_);
  or g_126390_(_069293_, _069294_, _069295_);
  or g_126391_(_069281_, _069285_, _069296_);
  or g_126392_(_069290_, _069291_, _069297_);
  or g_126393_(_069296_, _069297_, _069298_);
  or g_126394_(_069295_, _069298_, _069300_);
  xor g_126395_(out[444], out[524], _069301_);
  or g_126396_(_069275_, _069301_, _069302_);
  or g_126397_(_069274_, _069286_, _069303_);
  or g_126398_(_069302_, _069303_, _069304_);
  or g_126399_(_069279_, _069284_, _069305_);
  or g_126400_(_069287_, _069305_, _069306_);
  or g_126401_(_069304_, _069306_, _069307_);
  or g_126402_(_069300_, _069307_, _069308_);
  or g_126403_(_069292_, _069308_, _069309_);
  not g_126404_(_069309_, _069311_);
  xor g_126405_(out[422], out[518], _069312_);
  xor g_126406_(out[417], out[513], _069313_);
  xor g_126407_(out[416], out[512], _069314_);
  xor g_126408_(out[418], out[514], _069315_);
  xor g_126409_(out[419], out[515], _069316_);
  xor g_126410_(out[425], out[521], _069317_);
  xor g_126411_(out[430], out[526], _069318_);
  and g_126412_(_049455_, out[523], _069319_);
  xor g_126413_(out[423], out[519], _069320_);
  and g_126414_(out[427], _049521_, _069322_);
  xor g_126415_(out[429], out[525], _069323_);
  xor g_126416_(out[424], out[520], _069324_);
  or g_126417_(_069323_, _069324_, _069325_);
  xor g_126418_(out[431], out[527], _069326_);
  xor g_126419_(out[426], out[522], _069327_);
  xor g_126420_(out[421], out[517], _069328_);
  xor g_126421_(out[420], out[516], _069329_);
  or g_126422_(_069315_, _069327_, _069330_);
  or g_126423_(_069325_, _069330_, _069331_);
  or g_126424_(_069316_, _069317_, _069333_);
  or g_126425_(_069328_, _069333_, _069334_);
  or g_126426_(_069331_, _069334_, _069335_);
  or g_126427_(_069318_, _069329_, _069336_);
  or g_126428_(_069335_, _069336_, _069337_);
  xor g_126429_(out[428], out[524], _069338_);
  or g_126430_(_069319_, _069338_, _069339_);
  or g_126431_(_069312_, _069320_, _069340_);
  or g_126432_(_069339_, _069340_, _069341_);
  or g_126433_(_069313_, _069322_, _069342_);
  or g_126434_(_069326_, _069342_, _069344_);
  or g_126435_(_069341_, _069344_, _069345_);
  or g_126436_(_069314_, _069345_, _069346_);
  or g_126437_(_069337_, _069346_, _069347_);
  not g_126438_(_069347_, _069348_);
  xor g_126439_(out[407], out[519], _069349_);
  and g_126440_(_049444_, out[523], _069350_);
  xor g_126441_(out[414], out[526], _069351_);
  xor g_126442_(out[408], out[520], _069352_);
  xor g_126443_(out[401], out[513], _069353_);
  xor g_126444_(out[413], out[525], _069355_);
  xor g_126445_(out[409], out[521], _069356_);
  xor g_126446_(out[404], out[516], _069357_);
  xor g_126447_(out[402], out[514], _069358_);
  and g_126448_(out[411], _049521_, _069359_);
  xor g_126449_(out[403], out[515], _069360_);
  xor g_126450_(out[406], out[518], _069361_);
  xor g_126451_(out[415], out[527], _069362_);
  xor g_126452_(out[410], out[522], _069363_);
  xor g_126453_(out[405], out[517], _069364_);
  xor g_126454_(out[400], out[512], _069366_);
  or g_126455_(_069351_, _069357_, _069367_);
  or g_126456_(_069352_, _069355_, _069368_);
  or g_126457_(_069358_, _069363_, _069369_);
  or g_126458_(_069368_, _069369_, _069370_);
  or g_126459_(_069356_, _069360_, _069371_);
  or g_126460_(_069364_, _069366_, _069372_);
  or g_126461_(_069371_, _069372_, _069373_);
  or g_126462_(_069370_, _069373_, _069374_);
  xor g_126463_(out[412], out[524], _069375_);
  or g_126464_(_069350_, _069375_, _069377_);
  or g_126465_(_069349_, _069361_, _069378_);
  or g_126466_(_069377_, _069378_, _069379_);
  or g_126467_(_069353_, _069359_, _069380_);
  or g_126468_(_069362_, _069380_, _069381_);
  or g_126469_(_069379_, _069381_, _069382_);
  or g_126470_(_069374_, _069382_, _069383_);
  or g_126471_(_069367_, _069383_, _069384_);
  xor g_126472_(out[385], out[513], _069385_);
  and g_126473_(out[395], _049521_, _069386_);
  xor g_126474_(out[393], out[521], _069388_);
  xor g_126475_(out[384], out[512], _069389_);
  xor g_126476_(out[398], out[526], _069390_);
  xor g_126477_(out[388], out[516], _069391_);
  or g_126478_(_069390_, _069391_, _069392_);
  xor g_126479_(out[397], out[525], _069393_);
  xor g_126480_(out[387], out[515], _069394_);
  and g_126481_(_049433_, out[523], _069395_);
  xor g_126482_(out[390], out[518], _069396_);
  xor g_126483_(out[394], out[522], _069397_);
  xor g_126484_(out[389], out[517], _069399_);
  xor g_126485_(out[399], out[527], _069400_);
  xor g_126486_(out[392], out[520], _069401_);
  or g_126487_(_069393_, _069401_, _069402_);
  xor g_126488_(out[386], out[514], _069403_);
  or g_126489_(_069397_, _069403_, _069404_);
  or g_126490_(_069402_, _069404_, _069405_);
  or g_126491_(_069388_, _069394_, _069406_);
  or g_126492_(_069399_, _069406_, _069407_);
  or g_126493_(_069405_, _069407_, _069408_);
  or g_126494_(_069392_, _069408_, _069410_);
  xor g_126495_(out[396], out[524], _069411_);
  or g_126496_(_069395_, _069411_, _069412_);
  xor g_126497_(out[391], out[519], _069413_);
  or g_126498_(_069396_, _069413_, _069414_);
  or g_126499_(_069412_, _069414_, _069415_);
  or g_126500_(_069385_, _069386_, _069416_);
  or g_126501_(_069400_, _069416_, _069417_);
  or g_126502_(_069415_, _069417_, _069418_);
  or g_126503_(_069389_, _069418_, _069419_);
  or g_126504_(_069410_, _069419_, _069421_);
  xor g_126505_(out[375], out[519], _069422_);
  and g_126506_(_049422_, out[523], _069423_);
  xor g_126507_(out[382], out[526], _069424_);
  xor g_126508_(out[376], out[520], _069425_);
  xor g_126509_(out[369], out[513], _069426_);
  xor g_126510_(out[381], out[525], _069427_);
  xor g_126511_(out[377], out[521], _069428_);
  xor g_126512_(out[372], out[516], _069429_);
  xor g_126513_(out[370], out[514], _069430_);
  and g_126514_(out[379], _049521_, _069432_);
  xor g_126515_(out[371], out[515], _069433_);
  xor g_126516_(out[374], out[518], _069434_);
  xor g_126517_(out[383], out[527], _069435_);
  xor g_126518_(out[378], out[522], _069436_);
  xor g_126519_(out[373], out[517], _069437_);
  xor g_126520_(out[368], out[512], _069438_);
  or g_126521_(_069424_, _069429_, _069439_);
  or g_126522_(_069425_, _069427_, _069440_);
  or g_126523_(_069430_, _069436_, _069441_);
  or g_126524_(_069440_, _069441_, _069443_);
  or g_126525_(_069428_, _069433_, _069444_);
  or g_126526_(_069437_, _069438_, _069445_);
  or g_126527_(_069444_, _069445_, _069446_);
  or g_126528_(_069443_, _069446_, _069447_);
  xor g_126529_(out[380], out[524], _069448_);
  or g_126530_(_069423_, _069448_, _069449_);
  or g_126531_(_069422_, _069434_, _069450_);
  or g_126532_(_069449_, _069450_, _069451_);
  or g_126533_(_069426_, _069432_, _069452_);
  or g_126534_(_069435_, _069452_, _069454_);
  or g_126535_(_069451_, _069454_, _069455_);
  or g_126536_(_069447_, _069455_, _069456_);
  or g_126537_(_069439_, _069456_, _069457_);
  xor g_126538_(out[353], out[513], _069458_);
  and g_126539_(_049411_, out[523], _069459_);
  and g_126540_(out[363], _049521_, _069460_);
  xor g_126541_(out[360], out[520], _069461_);
  xor g_126542_(out[362], out[522], _069462_);
  xor g_126543_(out[354], out[514], _069463_);
  xor g_126544_(out[356], out[516], _069465_);
  xor g_126545_(out[357], out[517], _069466_);
  xor g_126546_(out[361], out[521], _069467_);
  xor g_126547_(out[355], out[515], _069468_);
  xor g_126548_(out[366], out[526], _069469_);
  xor g_126549_(out[352], out[512], _069470_);
  xor g_126550_(out[367], out[527], _069471_);
  xor g_126551_(out[365], out[525], _069472_);
  or g_126552_(_069461_, _069472_, _069473_);
  xor g_126553_(out[358], out[518], _069474_);
  or g_126554_(_069462_, _069463_, _069476_);
  or g_126555_(_069473_, _069476_, _069477_);
  or g_126556_(_069467_, _069468_, _069478_);
  or g_126557_(_069466_, _069478_, _069479_);
  or g_126558_(_069477_, _069479_, _069480_);
  or g_126559_(_069465_, _069469_, _069481_);
  or g_126560_(_069480_, _069481_, _069482_);
  xor g_126561_(out[364], out[524], _069483_);
  or g_126562_(_069459_, _069483_, _069484_);
  xor g_126563_(out[359], out[519], _069485_);
  or g_126564_(_069474_, _069485_, _069487_);
  or g_126565_(_069484_, _069487_, _069488_);
  or g_126566_(_069458_, _069460_, _069489_);
  or g_126567_(_069471_, _069489_, _069490_);
  or g_126568_(_069488_, _069490_, _069491_);
  or g_126569_(_069470_, _069491_, _069492_);
  or g_126570_(_069482_, _069492_, _069493_);
  not g_126571_(_069493_, _069494_);
  xor g_126572_(out[343], out[519], _069495_);
  and g_126573_(_049400_, out[523], _069496_);
  xor g_126574_(out[350], out[526], _069498_);
  xor g_126575_(out[344], out[520], _069499_);
  xor g_126576_(out[337], out[513], _069500_);
  xor g_126577_(out[349], out[525], _069501_);
  xor g_126578_(out[345], out[521], _069502_);
  xor g_126579_(out[340], out[516], _069503_);
  xor g_126580_(out[338], out[514], _069504_);
  and g_126581_(out[347], _049521_, _069505_);
  xor g_126582_(out[339], out[515], _069506_);
  xor g_126583_(out[342], out[518], _069507_);
  xor g_126584_(out[351], out[527], _069509_);
  xor g_126585_(out[346], out[522], _069510_);
  xor g_126586_(out[341], out[517], _069511_);
  xor g_126587_(out[336], out[512], _069512_);
  or g_126588_(_069498_, _069503_, _069513_);
  or g_126589_(_069499_, _069501_, _069514_);
  or g_126590_(_069504_, _069510_, _069515_);
  or g_126591_(_069514_, _069515_, _069516_);
  or g_126592_(_069502_, _069506_, _069517_);
  or g_126593_(_069511_, _069512_, _069518_);
  or g_126594_(_069517_, _069518_, _069520_);
  or g_126595_(_069516_, _069520_, _069521_);
  xor g_126596_(out[348], out[524], _069522_);
  or g_126597_(_069496_, _069522_, _069523_);
  or g_126598_(_069495_, _069507_, _069524_);
  or g_126599_(_069523_, _069524_, _069525_);
  or g_126600_(_069500_, _069505_, _069526_);
  or g_126601_(_069509_, _069526_, _069527_);
  or g_126602_(_069525_, _069527_, _069528_);
  or g_126603_(_069521_, _069528_, _069529_);
  or g_126604_(_069513_, _069529_, _069531_);
  not g_126605_(_069531_, _069532_);
  and g_126606_(out[331], _049521_, _069533_);
  xor g_126607_(out[330], out[522], _069534_);
  xor g_126608_(out[335], out[527], _069535_);
  xor g_126609_(out[320], out[512], _069536_);
  xor g_126610_(out[321], out[513], _069537_);
  xor g_126611_(out[322], out[514], _069538_);
  xor g_126612_(out[323], out[515], _069539_);
  xor g_126613_(out[329], out[521], _069540_);
  xor g_126614_(out[334], out[526], _069542_);
  and g_126615_(_098294_, out[523], _069543_);
  xor g_126616_(out[325], out[517], _069544_);
  xor g_126617_(out[326], out[518], _069545_);
  xor g_126618_(out[324], out[516], _069546_);
  xor g_126619_(out[333], out[525], _069547_);
  xor g_126620_(out[328], out[520], _069548_);
  or g_126621_(_069547_, _069548_, _069549_);
  or g_126622_(_069534_, _069538_, _069550_);
  or g_126623_(_069549_, _069550_, _069551_);
  or g_126624_(_069539_, _069540_, _069553_);
  or g_126625_(_069544_, _069553_, _069554_);
  or g_126626_(_069551_, _069554_, _069555_);
  or g_126627_(_069542_, _069546_, _069556_);
  or g_126628_(_069555_, _069556_, _069557_);
  xor g_126629_(out[332], out[524], _069558_);
  or g_126630_(_069543_, _069558_, _069559_);
  xor g_126631_(out[327], out[519], _069560_);
  or g_126632_(_069545_, _069560_, _069561_);
  or g_126633_(_069559_, _069561_, _069562_);
  or g_126634_(_069533_, _069537_, _069564_);
  or g_126635_(_069535_, _069564_, _069565_);
  or g_126636_(_069562_, _069565_, _069566_);
  or g_126637_(_069536_, _069566_, _069567_);
  or g_126638_(_069557_, _069567_, _069568_);
  not g_126639_(_069568_, _069569_);
  xor g_126640_(out[311], out[519], _069570_);
  and g_126641_(_098283_, out[523], _069571_);
  xor g_126642_(out[318], out[526], _069572_);
  xor g_126643_(out[312], out[520], _069573_);
  xor g_126644_(out[305], out[513], _069575_);
  xor g_126645_(out[317], out[525], _069576_);
  xor g_126646_(out[313], out[521], _069577_);
  xor g_126647_(out[308], out[516], _069578_);
  xor g_126648_(out[306], out[514], _069579_);
  and g_126649_(out[315], _049521_, _069580_);
  xor g_126650_(out[307], out[515], _069581_);
  xor g_126651_(out[310], out[518], _069582_);
  xor g_126652_(out[319], out[527], _069583_);
  xor g_126653_(out[314], out[522], _069584_);
  xor g_126654_(out[309], out[517], _069586_);
  xor g_126655_(out[304], out[512], _069587_);
  or g_126656_(_069572_, _069578_, _069588_);
  or g_126657_(_069573_, _069576_, _069589_);
  or g_126658_(_069579_, _069584_, _069590_);
  or g_126659_(_069589_, _069590_, _069591_);
  or g_126660_(_069577_, _069581_, _069592_);
  or g_126661_(_069586_, _069587_, _069593_);
  or g_126662_(_069592_, _069593_, _069594_);
  or g_126663_(_069591_, _069594_, _069595_);
  xor g_126664_(out[316], out[524], _069597_);
  or g_126665_(_069571_, _069597_, _069598_);
  or g_126666_(_069570_, _069582_, _069599_);
  or g_126667_(_069598_, _069599_, _069600_);
  or g_126668_(_069575_, _069580_, _069601_);
  or g_126669_(_069583_, _069601_, _069602_);
  or g_126670_(_069600_, _069602_, _069603_);
  or g_126671_(_069595_, _069603_, _069604_);
  or g_126672_(_069588_, _069604_, _069605_);
  not g_126673_(_069605_, _069606_);
  xor g_126674_(out[289], out[513], _069608_);
  and g_126675_(_098272_, out[523], _069609_);
  and g_126676_(out[299], _049521_, _069610_);
  xor g_126677_(out[296], out[520], _069611_);
  xor g_126678_(out[298], out[522], _069612_);
  xor g_126679_(out[290], out[514], _069613_);
  xor g_126680_(out[292], out[516], _069614_);
  xor g_126681_(out[293], out[517], _069615_);
  xor g_126682_(out[297], out[521], _069616_);
  xor g_126683_(out[291], out[515], _069617_);
  xor g_126684_(out[302], out[526], _069619_);
  xor g_126685_(out[288], out[512], _069620_);
  xor g_126686_(out[303], out[527], _069621_);
  xor g_126687_(out[301], out[525], _069622_);
  or g_126688_(_069611_, _069622_, _069623_);
  xor g_126689_(out[294], out[518], _069624_);
  or g_126690_(_069612_, _069613_, _069625_);
  or g_126691_(_069623_, _069625_, _069626_);
  or g_126692_(_069616_, _069617_, _069627_);
  or g_126693_(_069615_, _069627_, _069628_);
  or g_126694_(_069626_, _069628_, _069630_);
  or g_126695_(_069614_, _069619_, _069631_);
  or g_126696_(_069630_, _069631_, _069632_);
  xor g_126697_(out[300], out[524], _069633_);
  or g_126698_(_069609_, _069633_, _069634_);
  xor g_126699_(out[295], out[519], _069635_);
  or g_126700_(_069624_, _069635_, _069636_);
  or g_126701_(_069634_, _069636_, _069637_);
  or g_126702_(_069608_, _069610_, _069638_);
  or g_126703_(_069621_, _069638_, _069639_);
  or g_126704_(_069637_, _069639_, _069641_);
  or g_126705_(_069620_, _069641_, _069642_);
  or g_126706_(_069632_, _069642_, _069643_);
  not g_126707_(_069643_, _069644_);
  xor g_126708_(out[279], out[519], _069645_);
  and g_126709_(_098261_, out[523], _069646_);
  xor g_126710_(out[286], out[526], _069647_);
  xor g_126711_(out[280], out[520], _069648_);
  xor g_126712_(out[273], out[513], _069649_);
  xor g_126713_(out[285], out[525], _069650_);
  xor g_126714_(out[281], out[521], _069652_);
  xor g_126715_(out[276], out[516], _069653_);
  xor g_126716_(out[274], out[514], _069654_);
  and g_126717_(out[283], _049521_, _069655_);
  xor g_126718_(out[275], out[515], _069656_);
  xor g_126719_(out[278], out[518], _069657_);
  xor g_126720_(out[287], out[527], _069658_);
  xor g_126721_(out[282], out[522], _069659_);
  xor g_126722_(out[277], out[517], _069660_);
  xor g_126723_(out[272], out[512], _069661_);
  or g_126724_(_069647_, _069653_, _069663_);
  or g_126725_(_069648_, _069650_, _069664_);
  or g_126726_(_069654_, _069659_, _069665_);
  or g_126727_(_069664_, _069665_, _069666_);
  or g_126728_(_069652_, _069656_, _069667_);
  or g_126729_(_069660_, _069661_, _069668_);
  or g_126730_(_069667_, _069668_, _069669_);
  or g_126731_(_069666_, _069669_, _069670_);
  xor g_126732_(out[284], out[524], _069671_);
  or g_126733_(_069646_, _069671_, _069672_);
  or g_126734_(_069645_, _069657_, _069674_);
  or g_126735_(_069672_, _069674_, _069675_);
  or g_126736_(_069649_, _069655_, _069676_);
  or g_126737_(_069658_, _069676_, _069677_);
  or g_126738_(_069675_, _069677_, _069678_);
  or g_126739_(_069670_, _069678_, _069679_);
  or g_126740_(_069663_, _069679_, _069680_);
  and g_126741_(out[267], _049521_, _069681_);
  xor g_126742_(out[260], out[516], _069682_);
  xor g_126743_(out[270], out[526], _069683_);
  or g_126744_(_069682_, _069683_, _069685_);
  xor g_126745_(out[269], out[525], _069686_);
  xor g_126746_(out[259], out[515], _069687_);
  xor g_126747_(out[256], out[512], _069688_);
  and g_126748_(_098250_, out[523], _069689_);
  xor g_126749_(out[266], out[522], _069690_);
  xor g_126750_(out[271], out[527], _069691_);
  xor g_126751_(out[262], out[518], _069692_);
  xor g_126752_(out[261], out[517], _069693_);
  xor g_126753_(out[264], out[520], _069694_);
  or g_126754_(_069686_, _069694_, _069696_);
  xor g_126755_(out[258], out[514], _069697_);
  xor g_126756_(out[265], out[521], _069698_);
  xor g_126757_(out[257], out[513], _069699_);
  or g_126758_(_069690_, _069697_, _069700_);
  or g_126759_(_069696_, _069700_, _069701_);
  or g_126760_(_069687_, _069698_, _069702_);
  or g_126761_(_069693_, _069702_, _069703_);
  or g_126762_(_069701_, _069703_, _069704_);
  or g_126763_(_069685_, _069704_, _069705_);
  xor g_126764_(out[268], out[524], _069707_);
  or g_126765_(_069689_, _069707_, _069708_);
  xor g_126766_(out[263], out[519], _069709_);
  or g_126767_(_069692_, _069709_, _069710_);
  or g_126768_(_069708_, _069710_, _069711_);
  or g_126769_(_069681_, _069699_, _069712_);
  or g_126770_(_069691_, _069712_, _069713_);
  or g_126771_(_069711_, _069713_, _069714_);
  or g_126772_(_069688_, _069714_, _069715_);
  or g_126773_(_069705_, _069715_, _069716_);
  not g_126774_(_069716_, _069718_);
  xor g_126775_(out[247], out[519], _069719_);
  and g_126776_(_098239_, out[523], _069720_);
  xor g_126777_(out[254], out[526], _069721_);
  xor g_126778_(out[248], out[520], _069722_);
  xor g_126779_(out[241], out[513], _069723_);
  xor g_126780_(out[253], out[525], _069724_);
  xor g_126781_(out[249], out[521], _069725_);
  xor g_126782_(out[244], out[516], _069726_);
  xor g_126783_(out[242], out[514], _069727_);
  and g_126784_(out[251], _049521_, _069729_);
  xor g_126785_(out[243], out[515], _069730_);
  xor g_126786_(out[246], out[518], _069731_);
  xor g_126787_(out[255], out[527], _069732_);
  xor g_126788_(out[250], out[522], _069733_);
  xor g_126789_(out[245], out[517], _069734_);
  xor g_126790_(out[240], out[512], _069735_);
  or g_126791_(_069721_, _069726_, _069736_);
  or g_126792_(_069722_, _069724_, _069737_);
  or g_126793_(_069727_, _069733_, _069738_);
  or g_126794_(_069737_, _069738_, _069740_);
  or g_126795_(_069725_, _069730_, _069741_);
  or g_126796_(_069734_, _069735_, _069742_);
  or g_126797_(_069741_, _069742_, _069743_);
  or g_126798_(_069740_, _069743_, _069744_);
  xor g_126799_(out[252], out[524], _069745_);
  or g_126800_(_069720_, _069745_, _069746_);
  or g_126801_(_069719_, _069731_, _069747_);
  or g_126802_(_069746_, _069747_, _069748_);
  or g_126803_(_069723_, _069729_, _069749_);
  or g_126804_(_069732_, _069749_, _069751_);
  or g_126805_(_069748_, _069751_, _069752_);
  or g_126806_(_069744_, _069752_, _069753_);
  or g_126807_(_069736_, _069753_, _069754_);
  not g_126808_(_069754_, _069755_);
  and g_126809_(out[235], _049521_, _069756_);
  xor g_126810_(out[228], out[516], _069757_);
  xor g_126811_(out[238], out[526], _069758_);
  or g_126812_(_069757_, _069758_, _069759_);
  xor g_126813_(out[237], out[525], _069760_);
  xor g_126814_(out[227], out[515], _069762_);
  xor g_126815_(out[224], out[512], _069763_);
  and g_126816_(_098228_, out[523], _069764_);
  xor g_126817_(out[234], out[522], _069765_);
  xor g_126818_(out[239], out[527], _069766_);
  xor g_126819_(out[230], out[518], _069767_);
  xor g_126820_(out[229], out[517], _069768_);
  xor g_126821_(out[232], out[520], _069769_);
  or g_126822_(_069760_, _069769_, _069770_);
  xor g_126823_(out[226], out[514], _069771_);
  xor g_126824_(out[233], out[521], _069773_);
  xor g_126825_(out[225], out[513], _069774_);
  or g_126826_(_069765_, _069771_, _069775_);
  or g_126827_(_069770_, _069775_, _069776_);
  or g_126828_(_069762_, _069773_, _069777_);
  or g_126829_(_069768_, _069777_, _069778_);
  or g_126830_(_069776_, _069778_, _069779_);
  or g_126831_(_069759_, _069779_, _069780_);
  xor g_126832_(out[236], out[524], _069781_);
  or g_126833_(_069764_, _069781_, _069782_);
  xor g_126834_(out[231], out[519], _069784_);
  or g_126835_(_069767_, _069784_, _069785_);
  or g_126836_(_069782_, _069785_, _069786_);
  or g_126837_(_069756_, _069774_, _069787_);
  or g_126838_(_069766_, _069787_, _069788_);
  or g_126839_(_069786_, _069788_, _069789_);
  or g_126840_(_069763_, _069789_, _069790_);
  or g_126841_(_069780_, _069790_, _069791_);
  xor g_126842_(out[215], out[519], _069792_);
  and g_126843_(_098217_, out[523], _069793_);
  xor g_126844_(out[222], out[526], _069795_);
  xor g_126845_(out[216], out[520], _069796_);
  xor g_126846_(out[209], out[513], _069797_);
  xor g_126847_(out[221], out[525], _069798_);
  xor g_126848_(out[217], out[521], _069799_);
  xor g_126849_(out[212], out[516], _069800_);
  xor g_126850_(out[210], out[514], _069801_);
  and g_126851_(out[219], _049521_, _069802_);
  xor g_126852_(out[211], out[515], _069803_);
  xor g_126853_(out[214], out[518], _069804_);
  xor g_126854_(out[223], out[527], _069806_);
  xor g_126855_(out[218], out[522], _069807_);
  xor g_126856_(out[213], out[517], _069808_);
  xor g_126857_(out[208], out[512], _069809_);
  or g_126858_(_069795_, _069800_, _069810_);
  or g_126859_(_069796_, _069798_, _069811_);
  or g_126860_(_069801_, _069807_, _069812_);
  or g_126861_(_069811_, _069812_, _069813_);
  or g_126862_(_069799_, _069803_, _069814_);
  or g_126863_(_069808_, _069809_, _069815_);
  or g_126864_(_069814_, _069815_, _069817_);
  or g_126865_(_069813_, _069817_, _069818_);
  xor g_126866_(out[220], out[524], _069819_);
  or g_126867_(_069793_, _069819_, _069820_);
  or g_126868_(_069792_, _069804_, _069821_);
  or g_126869_(_069820_, _069821_, _069822_);
  or g_126870_(_069797_, _069802_, _069823_);
  or g_126871_(_069806_, _069823_, _069824_);
  or g_126872_(_069822_, _069824_, _069825_);
  or g_126873_(_069818_, _069825_, _069826_);
  or g_126874_(_069810_, _069826_, _069828_);
  xor g_126875_(out[204], out[524], _069829_);
  and g_126876_(_098206_, out[523], _069830_);
  xor g_126877_(out[205], out[525], _069831_);
  xor g_126878_(out[198], out[518], _069832_);
  xor g_126879_(out[200], out[520], _069833_);
  xor g_126880_(out[201], out[521], _069834_);
  xor g_126881_(out[206], out[526], _069835_);
  xor g_126882_(out[196], out[516], _069836_);
  or g_126883_(_069835_, _069836_, _069837_);
  xor g_126884_(out[197], out[517], _069839_);
  xor g_126885_(out[193], out[513], _069840_);
  and g_126886_(out[203], _049521_, _069841_);
  xor g_126887_(out[207], out[527], _069842_);
  xor g_126888_(out[202], out[522], _069843_);
  xor g_126889_(out[192], out[512], _069844_);
  xor g_126890_(out[194], out[514], _069845_);
  xor g_126891_(out[195], out[515], _069846_);
  or g_126892_(_069831_, _069833_, _069847_);
  or g_126893_(_069843_, _069845_, _069848_);
  or g_126894_(_069847_, _069848_, _069850_);
  or g_126895_(_069834_, _069846_, _069851_);
  or g_126896_(_069839_, _069844_, _069852_);
  or g_126897_(_069851_, _069852_, _069853_);
  or g_126898_(_069850_, _069853_, _069854_);
  or g_126899_(_069829_, _069830_, _069855_);
  xor g_126900_(out[199], out[519], _069856_);
  or g_126901_(_069832_, _069856_, _069857_);
  or g_126902_(_069855_, _069857_, _069858_);
  or g_126903_(_069840_, _069841_, _069859_);
  or g_126904_(_069842_, _069859_, _069861_);
  or g_126905_(_069858_, _069861_, _069862_);
  or g_126906_(_069854_, _069862_, _069863_);
  or g_126907_(_069837_, _069863_, _069864_);
  not g_126908_(_069864_, _069865_);
  xor g_126909_(out[183], out[519], _069866_);
  and g_126910_(_098195_, out[523], _069867_);
  xor g_126911_(out[190], out[526], _069868_);
  xor g_126912_(out[184], out[520], _069869_);
  xor g_126913_(out[177], out[513], _069870_);
  xor g_126914_(out[189], out[525], _069872_);
  xor g_126915_(out[185], out[521], _069873_);
  xor g_126916_(out[180], out[516], _069874_);
  xor g_126917_(out[178], out[514], _069875_);
  and g_126918_(out[187], _049521_, _069876_);
  xor g_126919_(out[179], out[515], _069877_);
  xor g_126920_(out[182], out[518], _069878_);
  xor g_126921_(out[191], out[527], _069879_);
  xor g_126922_(out[186], out[522], _069880_);
  xor g_126923_(out[181], out[517], _069881_);
  xor g_126924_(out[176], out[512], _069883_);
  or g_126925_(_069868_, _069874_, _069884_);
  or g_126926_(_069869_, _069872_, _069885_);
  or g_126927_(_069875_, _069880_, _069886_);
  or g_126928_(_069885_, _069886_, _069887_);
  or g_126929_(_069873_, _069877_, _069888_);
  or g_126930_(_069881_, _069883_, _069889_);
  or g_126931_(_069888_, _069889_, _069890_);
  or g_126932_(_069887_, _069890_, _069891_);
  xor g_126933_(out[188], out[524], _069892_);
  or g_126934_(_069867_, _069892_, _069894_);
  or g_126935_(_069866_, _069878_, _069895_);
  or g_126936_(_069894_, _069895_, _069896_);
  or g_126937_(_069870_, _069876_, _069897_);
  or g_126938_(_069879_, _069897_, _069898_);
  or g_126939_(_069896_, _069898_, _069899_);
  or g_126940_(_069891_, _069899_, _069900_);
  or g_126941_(_069884_, _069900_, _069901_);
  xor g_126942_(out[172], out[524], _069902_);
  and g_126943_(_098184_, out[523], _069903_);
  xor g_126944_(out[168], out[520], _069905_);
  xor g_126945_(out[166], out[518], _069906_);
  xor g_126946_(out[173], out[525], _069907_);
  xor g_126947_(out[174], out[526], _069908_);
  xor g_126948_(out[162], out[514], _069909_);
  xor g_126949_(out[169], out[521], _069910_);
  xor g_126950_(out[165], out[517], _069911_);
  xor g_126951_(out[161], out[513], _069912_);
  and g_126952_(out[171], _049521_, _069913_);
  or g_126953_(_069905_, _069907_, _069914_);
  xor g_126954_(out[175], out[527], _069916_);
  xor g_126955_(out[170], out[522], _069917_);
  xor g_126956_(out[164], out[516], _069918_);
  xor g_126957_(out[163], out[515], _069919_);
  xor g_126958_(out[160], out[512], _069920_);
  or g_126959_(_069909_, _069917_, _069921_);
  or g_126960_(_069914_, _069921_, _069922_);
  or g_126961_(_069910_, _069919_, _069923_);
  or g_126962_(_069911_, _069923_, _069924_);
  or g_126963_(_069922_, _069924_, _069925_);
  or g_126964_(_069908_, _069918_, _069927_);
  or g_126965_(_069925_, _069927_, _069928_);
  or g_126966_(_069902_, _069903_, _069929_);
  xor g_126967_(out[167], out[519], _069930_);
  or g_126968_(_069906_, _069930_, _069931_);
  or g_126969_(_069929_, _069931_, _069932_);
  or g_126970_(_069912_, _069913_, _069933_);
  or g_126971_(_069916_, _069933_, _069934_);
  or g_126972_(_069932_, _069934_, _069935_);
  or g_126973_(_069920_, _069935_, _069936_);
  or g_126974_(_069928_, _069936_, _069938_);
  xor g_126975_(out[151], out[519], _069939_);
  and g_126976_(_098173_, out[523], _069940_);
  xor g_126977_(out[158], out[526], _069941_);
  xor g_126978_(out[152], out[520], _069942_);
  xor g_126979_(out[145], out[513], _069943_);
  xor g_126980_(out[157], out[525], _069944_);
  xor g_126981_(out[153], out[521], _069945_);
  xor g_126982_(out[148], out[516], _069946_);
  xor g_126983_(out[146], out[514], _069947_);
  and g_126984_(out[155], _049521_, _069949_);
  xor g_126985_(out[147], out[515], _069950_);
  xor g_126986_(out[150], out[518], _069951_);
  xor g_126987_(out[159], out[527], _069952_);
  xor g_126988_(out[154], out[522], _069953_);
  xor g_126989_(out[149], out[517], _069954_);
  xor g_126990_(out[144], out[512], _069955_);
  or g_126991_(_069941_, _069946_, _069956_);
  or g_126992_(_069942_, _069944_, _069957_);
  or g_126993_(_069947_, _069953_, _069958_);
  or g_126994_(_069957_, _069958_, _069960_);
  or g_126995_(_069945_, _069950_, _069961_);
  or g_126996_(_069954_, _069955_, _069962_);
  or g_126997_(_069961_, _069962_, _069963_);
  or g_126998_(_069960_, _069963_, _069964_);
  xor g_126999_(out[156], out[524], _069965_);
  or g_127000_(_069940_, _069965_, _069966_);
  or g_127001_(_069939_, _069951_, _069967_);
  or g_127002_(_069966_, _069967_, _069968_);
  or g_127003_(_069943_, _069949_, _069969_);
  or g_127004_(_069952_, _069969_, _069971_);
  or g_127005_(_069968_, _069971_, _069972_);
  or g_127006_(_069964_, _069972_, _069973_);
  or g_127007_(_069956_, _069973_, _069974_);
  not g_127008_(_069974_, _069975_);
  xor g_127009_(out[138], out[522], _069976_);
  xor g_127010_(out[130], out[514], _069977_);
  xor g_127011_(out[129], out[513], _069978_);
  and g_127012_(_098162_, out[523], _069979_);
  and g_127013_(out[139], _049521_, _069980_);
  xor g_127014_(out[141], out[525], _069982_);
  xor g_127015_(out[131], out[515], _069983_);
  xor g_127016_(out[142], out[526], _069984_);
  xor g_127017_(out[140], out[524], _069985_);
  xor g_127018_(out[136], out[520], _069986_);
  xor g_127019_(out[143], out[527], _069987_);
  xor g_127020_(out[133], out[517], _069988_);
  xor g_127021_(out[134], out[518], _069989_);
  xor g_127022_(out[128], out[512], _069990_);
  xor g_127023_(out[132], out[516], _069991_);
  or g_127024_(_069982_, _069986_, _069993_);
  xor g_127025_(out[137], out[521], _069994_);
  or g_127026_(_069976_, _069977_, _069995_);
  or g_127027_(_069993_, _069995_, _069996_);
  or g_127028_(_069983_, _069994_, _069997_);
  or g_127029_(_069988_, _069997_, _069998_);
  or g_127030_(_069996_, _069998_, _069999_);
  or g_127031_(_069984_, _069991_, _070000_);
  or g_127032_(_069999_, _070000_, _070001_);
  or g_127033_(_069979_, _069985_, _070002_);
  xor g_127034_(out[135], out[519], _070004_);
  or g_127035_(_069989_, _070004_, _070005_);
  or g_127036_(_070002_, _070005_, _070006_);
  or g_127037_(_069978_, _069980_, _070007_);
  or g_127038_(_069987_, _070007_, _070008_);
  or g_127039_(_070006_, _070008_, _070009_);
  or g_127040_(_069990_, _070009_, _070010_);
  or g_127041_(_070001_, _070010_, _070011_);
  not g_127042_(_070011_, _070012_);
  xor g_127043_(out[119], out[519], _070013_);
  and g_127044_(_098151_, out[523], _070015_);
  xor g_127045_(out[126], out[526], _070016_);
  xor g_127046_(out[120], out[520], _070017_);
  xor g_127047_(out[113], out[513], _070018_);
  xor g_127048_(out[125], out[525], _070019_);
  xor g_127049_(out[121], out[521], _070020_);
  xor g_127050_(out[116], out[516], _070021_);
  xor g_127051_(out[114], out[514], _070022_);
  and g_127052_(out[123], _049521_, _070023_);
  xor g_127053_(out[115], out[515], _070024_);
  xor g_127054_(out[118], out[518], _070026_);
  xor g_127055_(out[127], out[527], _070027_);
  xor g_127056_(out[122], out[522], _070028_);
  xor g_127057_(out[117], out[517], _070029_);
  xor g_127058_(out[112], out[512], _070030_);
  or g_127059_(_070016_, _070021_, _070031_);
  or g_127060_(_070017_, _070019_, _070032_);
  or g_127061_(_070022_, _070028_, _070033_);
  or g_127062_(_070032_, _070033_, _070034_);
  or g_127063_(_070020_, _070024_, _070035_);
  or g_127064_(_070029_, _070030_, _070037_);
  or g_127065_(_070035_, _070037_, _070038_);
  or g_127066_(_070034_, _070038_, _070039_);
  xor g_127067_(out[124], out[524], _070040_);
  or g_127068_(_070015_, _070040_, _070041_);
  or g_127069_(_070013_, _070026_, _070042_);
  or g_127070_(_070041_, _070042_, _070043_);
  or g_127071_(_070018_, _070023_, _070044_);
  or g_127072_(_070027_, _070044_, _070045_);
  or g_127073_(_070043_, _070045_, _070046_);
  or g_127074_(_070039_, _070046_, _070048_);
  or g_127075_(_070031_, _070048_, _070049_);
  and g_127076_(out[107], _049521_, _070050_);
  and g_127077_(_098140_, out[523], _070051_);
  xor g_127078_(out[104], out[520], _070052_);
  xor g_127079_(out[111], out[527], _070053_);
  xor g_127080_(out[97], out[513], _070054_);
  xor g_127081_(out[98], out[514], _070055_);
  xor g_127082_(out[100], out[516], _070056_);
  xor g_127083_(out[109], out[525], _070057_);
  xor g_127084_(out[105], out[521], _070059_);
  xor g_127085_(out[99], out[515], _070060_);
  xor g_127086_(out[101], out[517], _070061_);
  xor g_127087_(out[110], out[526], _070062_);
  xor g_127088_(out[96], out[512], _070063_);
  xor g_127089_(out[106], out[522], _070064_);
  or g_127090_(_070052_, _070057_, _070065_);
  xor g_127091_(out[102], out[518], _070066_);
  or g_127092_(_070055_, _070064_, _070067_);
  or g_127093_(_070065_, _070067_, _070068_);
  or g_127094_(_070059_, _070060_, _070070_);
  or g_127095_(_070061_, _070070_, _070071_);
  or g_127096_(_070068_, _070071_, _070072_);
  or g_127097_(_070056_, _070062_, _070073_);
  or g_127098_(_070072_, _070073_, _070074_);
  xor g_127099_(out[108], out[524], _070075_);
  or g_127100_(_070051_, _070075_, _070076_);
  xor g_127101_(out[103], out[519], _070077_);
  or g_127102_(_070066_, _070077_, _070078_);
  or g_127103_(_070076_, _070078_, _070079_);
  or g_127104_(_070050_, _070054_, _070081_);
  or g_127105_(_070053_, _070081_, _070082_);
  or g_127106_(_070079_, _070082_, _070083_);
  or g_127107_(_070063_, _070083_, _070084_);
  or g_127108_(_070074_, _070084_, _070085_);
  xor g_127109_(out[87], out[519], _070086_);
  and g_127110_(_098129_, out[523], _070087_);
  xor g_127111_(out[94], out[526], _070088_);
  xor g_127112_(out[88], out[520], _070089_);
  xor g_127113_(out[81], out[513], _070090_);
  xor g_127114_(out[93], out[525], _070092_);
  xor g_127115_(out[89], out[521], _070093_);
  xor g_127116_(out[84], out[516], _070094_);
  xor g_127117_(out[82], out[514], _070095_);
  and g_127118_(out[91], _049521_, _070096_);
  xor g_127119_(out[83], out[515], _070097_);
  xor g_127120_(out[86], out[518], _070098_);
  xor g_127121_(out[95], out[527], _070099_);
  xor g_127122_(out[90], out[522], _070100_);
  xor g_127123_(out[85], out[517], _070101_);
  xor g_127124_(out[80], out[512], _070103_);
  or g_127125_(_070088_, _070094_, _070104_);
  or g_127126_(_070089_, _070092_, _070105_);
  or g_127127_(_070095_, _070100_, _070106_);
  or g_127128_(_070105_, _070106_, _070107_);
  or g_127129_(_070093_, _070097_, _070108_);
  or g_127130_(_070101_, _070103_, _070109_);
  or g_127131_(_070108_, _070109_, _070110_);
  or g_127132_(_070107_, _070110_, _070111_);
  xor g_127133_(out[92], out[524], _070112_);
  or g_127134_(_070087_, _070112_, _070114_);
  or g_127135_(_070086_, _070098_, _070115_);
  or g_127136_(_070114_, _070115_, _070116_);
  or g_127137_(_070090_, _070096_, _070117_);
  or g_127138_(_070099_, _070117_, _070118_);
  or g_127139_(_070116_, _070118_, _070119_);
  or g_127140_(_070111_, _070119_, _070120_);
  or g_127141_(_070104_, _070120_, _070121_);
  not g_127142_(_070121_, _070122_);
  xor g_127143_(out[65], out[513], _070123_);
  and g_127144_(out[75], _049521_, _070125_);
  xor g_127145_(out[73], out[521], _070126_);
  xor g_127146_(out[64], out[512], _070127_);
  xor g_127147_(out[78], out[526], _070128_);
  xor g_127148_(out[68], out[516], _070129_);
  or g_127149_(_070128_, _070129_, _070130_);
  xor g_127150_(out[77], out[525], _070131_);
  xor g_127151_(out[67], out[515], _070132_);
  and g_127152_(_098118_, out[523], _070133_);
  xor g_127153_(out[70], out[518], _070134_);
  xor g_127154_(out[74], out[522], _070136_);
  xor g_127155_(out[69], out[517], _070137_);
  xor g_127156_(out[79], out[527], _070138_);
  xor g_127157_(out[72], out[520], _070139_);
  or g_127158_(_070131_, _070139_, _070140_);
  xor g_127159_(out[66], out[514], _070141_);
  or g_127160_(_070136_, _070141_, _070142_);
  or g_127161_(_070140_, _070142_, _070143_);
  or g_127162_(_070126_, _070132_, _070144_);
  or g_127163_(_070137_, _070144_, _070145_);
  or g_127164_(_070143_, _070145_, _070147_);
  or g_127165_(_070130_, _070147_, _070148_);
  xor g_127166_(out[76], out[524], _070149_);
  or g_127167_(_070133_, _070149_, _070150_);
  xor g_127168_(out[71], out[519], _070151_);
  or g_127169_(_070134_, _070151_, _070152_);
  or g_127170_(_070150_, _070152_, _070153_);
  or g_127171_(_070123_, _070125_, _070154_);
  or g_127172_(_070138_, _070154_, _070155_);
  or g_127173_(_070153_, _070155_, _070156_);
  or g_127174_(_070127_, _070156_, _070158_);
  or g_127175_(_070148_, _070158_, _070159_);
  xor g_127176_(out[55], out[519], _070160_);
  and g_127177_(_098107_, out[523], _070161_);
  xor g_127178_(out[62], out[526], _070162_);
  xor g_127179_(out[56], out[520], _070163_);
  xor g_127180_(out[49], out[513], _070164_);
  xor g_127181_(out[61], out[525], _070165_);
  xor g_127182_(out[57], out[521], _070166_);
  xor g_127183_(out[52], out[516], _070167_);
  xor g_127184_(out[50], out[514], _070169_);
  and g_127185_(out[59], _049521_, _070170_);
  xor g_127186_(out[51], out[515], _070171_);
  xor g_127187_(out[54], out[518], _070172_);
  xor g_127188_(out[63], out[527], _070173_);
  xor g_127189_(out[58], out[522], _070174_);
  xor g_127190_(out[53], out[517], _070175_);
  xor g_127191_(out[48], out[512], _070176_);
  or g_127192_(_070162_, _070167_, _070177_);
  or g_127193_(_070163_, _070165_, _070178_);
  or g_127194_(_070169_, _070174_, _070180_);
  or g_127195_(_070178_, _070180_, _070181_);
  or g_127196_(_070166_, _070171_, _070182_);
  or g_127197_(_070175_, _070176_, _070183_);
  or g_127198_(_070182_, _070183_, _070184_);
  or g_127199_(_070181_, _070184_, _070185_);
  xor g_127200_(out[60], out[524], _070186_);
  or g_127201_(_070161_, _070186_, _070187_);
  or g_127202_(_070160_, _070172_, _070188_);
  or g_127203_(_070187_, _070188_, _070189_);
  or g_127204_(_070164_, _070170_, _070191_);
  or g_127205_(_070173_, _070191_, _070192_);
  or g_127206_(_070189_, _070192_, _070193_);
  or g_127207_(_070185_, _070193_, _070194_);
  or g_127208_(_070177_, _070194_, _070195_);
  xor g_127209_(out[33], out[513], _070196_);
  and g_127210_(out[43], _049521_, _070197_);
  xor g_127211_(out[41], out[521], _070198_);
  xor g_127212_(out[32], out[512], _070199_);
  xor g_127213_(out[46], out[526], _070200_);
  xor g_127214_(out[36], out[516], _070202_);
  or g_127215_(_070200_, _070202_, _070203_);
  xor g_127216_(out[45], out[525], _070204_);
  xor g_127217_(out[35], out[515], _070205_);
  and g_127218_(_098096_, out[523], _070206_);
  xor g_127219_(out[38], out[518], _070207_);
  xor g_127220_(out[42], out[522], _070208_);
  xor g_127221_(out[37], out[517], _070209_);
  xor g_127222_(out[47], out[527], _070210_);
  xor g_127223_(out[40], out[520], _070211_);
  or g_127224_(_070204_, _070211_, _070213_);
  xor g_127225_(out[34], out[514], _070214_);
  or g_127226_(_070208_, _070214_, _070215_);
  or g_127227_(_070213_, _070215_, _070216_);
  or g_127228_(_070198_, _070205_, _070217_);
  or g_127229_(_070209_, _070217_, _070218_);
  or g_127230_(_070216_, _070218_, _070219_);
  or g_127231_(_070203_, _070219_, _070220_);
  xor g_127232_(out[44], out[524], _070221_);
  or g_127233_(_070206_, _070221_, _070222_);
  xor g_127234_(out[39], out[519], _070224_);
  or g_127235_(_070207_, _070224_, _070225_);
  or g_127236_(_070222_, _070225_, _070226_);
  or g_127237_(_070196_, _070197_, _070227_);
  or g_127238_(_070210_, _070227_, _070228_);
  or g_127239_(_070226_, _070228_, _070229_);
  or g_127240_(_070199_, _070229_, _070230_);
  or g_127241_(_070220_, _070230_, _070231_);
  xor g_127242_(out[23], out[519], _070232_);
  and g_127243_(_098063_, out[523], _070233_);
  xor g_127244_(out[30], out[526], _070235_);
  xor g_127245_(out[24], out[520], _070236_);
  xor g_127246_(out[17], out[513], _070237_);
  xor g_127247_(out[29], out[525], _070238_);
  xor g_127248_(out[25], out[521], _070239_);
  xor g_127249_(out[20], out[516], _070240_);
  xor g_127250_(out[18], out[514], _070241_);
  and g_127251_(out[27], _049521_, _070242_);
  xor g_127252_(out[19], out[515], _070243_);
  xor g_127253_(out[22], out[518], _070244_);
  xor g_127254_(out[31], out[527], _070246_);
  xor g_127255_(out[26], out[522], _070247_);
  xor g_127256_(out[21], out[517], _070248_);
  xor g_127257_(out[16], out[512], _070249_);
  or g_127258_(_070235_, _070240_, _070250_);
  or g_127259_(_070236_, _070238_, _070251_);
  or g_127260_(_070241_, _070247_, _070252_);
  or g_127261_(_070251_, _070252_, _070253_);
  or g_127262_(_070239_, _070243_, _070254_);
  or g_127263_(_070248_, _070249_, _070255_);
  or g_127264_(_070254_, _070255_, _070257_);
  or g_127265_(_070253_, _070257_, _070258_);
  xor g_127266_(out[28], out[524], _070259_);
  or g_127267_(_070233_, _070259_, _070260_);
  or g_127268_(_070232_, _070244_, _070261_);
  or g_127269_(_070260_, _070261_, _070262_);
  or g_127270_(_070237_, _070242_, _070263_);
  or g_127271_(_070246_, _070263_, _070264_);
  or g_127272_(_070262_, _070264_, _070265_);
  or g_127273_(_070258_, _070265_, _070266_);
  or g_127274_(_070250_, _070266_, _070268_);
  and g_127275_(out[11], _049521_, _070269_);
  xor g_127276_(out[4], out[516], _070270_);
  xor g_127277_(out[14], out[526], _070271_);
  or g_127278_(_070270_, _070271_, _070272_);
  xor g_127279_(out[13], out[525], _070273_);
  xor g_127280_(out[3], out[515], _070274_);
  xor g_127281_(out[0], out[512], _070275_);
  and g_127282_(_098041_, out[523], _070276_);
  xor g_127283_(out[10], out[522], _070277_);
  xor g_127284_(out[15], out[527], _070279_);
  xor g_127285_(out[6], out[518], _070280_);
  xor g_127286_(out[5], out[517], _070281_);
  xor g_127287_(out[8], out[520], _070282_);
  or g_127288_(_070273_, _070282_, _070283_);
  xor g_127289_(out[2], out[514], _070284_);
  xor g_127290_(out[9], out[521], _070285_);
  xor g_127291_(out[1], out[513], _070286_);
  or g_127292_(_070277_, _070284_, _070287_);
  or g_127293_(_070283_, _070287_, _070288_);
  or g_127294_(_070274_, _070285_, _070290_);
  or g_127295_(_070281_, _070290_, _070291_);
  or g_127296_(_070288_, _070291_, _070292_);
  or g_127297_(_070272_, _070292_, _070293_);
  not g_127298_(_070293_, _070294_);
  xor g_127299_(out[12], out[524], _070295_);
  or g_127300_(_070276_, _070295_, _070296_);
  xor g_127301_(out[7], out[519], _070297_);
  or g_127302_(_070280_, _070297_, _070298_);
  or g_127303_(_070296_, _070298_, _070299_);
  or g_127304_(_070269_, _070286_, _070301_);
  or g_127305_(_070279_, _070301_, _070302_);
  or g_127306_(_070299_, _070302_, _070303_);
  or g_127307_(_070275_, _070303_, _070304_);
  not g_127308_(_070304_, _070305_);
  and g_127309_(_070294_, _070305_, _070306_);
  not g_127310_(_070306_, _070307_);
  and g_127311_(out[475], _049510_, _070308_);
  xor g_127312_(out[468], out[500], _070309_);
  xor g_127313_(out[466], out[498], _070310_);
  xor g_127314_(out[473], out[505], _070312_);
  xor g_127315_(out[464], out[496], _070313_);
  xor g_127316_(out[467], out[499], _070314_);
  and g_127317_(_049499_, out[507], _070315_);
  xor g_127318_(out[474], out[506], _070316_);
  xor g_127319_(out[479], out[511], _070317_);
  xor g_127320_(out[470], out[502], _070318_);
  xor g_127321_(out[469], out[501], _070319_);
  xor g_127322_(out[477], out[509], _070320_);
  xor g_127323_(out[478], out[510], _070321_);
  xor g_127324_(out[472], out[504], _070323_);
  xor g_127325_(out[465], out[497], _070324_);
  or g_127326_(_070309_, _070321_, _070325_);
  or g_127327_(_070320_, _070323_, _070326_);
  or g_127328_(_070310_, _070316_, _070327_);
  or g_127329_(_070326_, _070327_, _070328_);
  or g_127330_(_070312_, _070314_, _070329_);
  or g_127331_(_070313_, _070319_, _070330_);
  or g_127332_(_070329_, _070330_, _070331_);
  or g_127333_(_070328_, _070331_, _070332_);
  xor g_127334_(out[476], out[508], _070334_);
  or g_127335_(_070315_, _070334_, _070335_);
  xor g_127336_(out[471], out[503], _070336_);
  or g_127337_(_070318_, _070336_, _070337_);
  or g_127338_(_070335_, _070337_, _070338_);
  or g_127339_(_070308_, _070324_, _070339_);
  or g_127340_(_070317_, _070339_, _070340_);
  or g_127341_(_070338_, _070340_, _070341_);
  or g_127342_(_070332_, _070341_, _070342_);
  or g_127343_(_070325_, _070342_, _070343_);
  xor g_127344_(out[455], out[503], _070345_);
  and g_127345_(_049477_, out[507], _070346_);
  xor g_127346_(out[462], out[510], _070347_);
  xor g_127347_(out[456], out[504], _070348_);
  xor g_127348_(out[449], out[497], _070349_);
  xor g_127349_(out[461], out[509], _070350_);
  xor g_127350_(out[457], out[505], _070351_);
  xor g_127351_(out[452], out[500], _070352_);
  xor g_127352_(out[450], out[498], _070353_);
  and g_127353_(out[459], _049510_, _070354_);
  xor g_127354_(out[451], out[499], _070356_);
  xor g_127355_(out[454], out[502], _070357_);
  xor g_127356_(out[463], out[511], _070358_);
  xor g_127357_(out[458], out[506], _070359_);
  xor g_127358_(out[453], out[501], _070360_);
  xor g_127359_(out[448], out[496], _070361_);
  or g_127360_(_070347_, _070352_, _070362_);
  or g_127361_(_070348_, _070350_, _070363_);
  or g_127362_(_070353_, _070359_, _070364_);
  or g_127363_(_070363_, _070364_, _070365_);
  or g_127364_(_070351_, _070356_, _070367_);
  or g_127365_(_070360_, _070361_, _070368_);
  or g_127366_(_070367_, _070368_, _070369_);
  or g_127367_(_070365_, _070369_, _070370_);
  xor g_127368_(out[460], out[508], _070371_);
  or g_127369_(_070346_, _070371_, _070372_);
  or g_127370_(_070345_, _070357_, _070373_);
  or g_127371_(_070372_, _070373_, _070374_);
  or g_127372_(_070349_, _070354_, _070375_);
  or g_127373_(_070358_, _070375_, _070376_);
  or g_127374_(_070374_, _070376_, _070378_);
  or g_127375_(_070370_, _070378_, _070379_);
  or g_127376_(_070362_, _070379_, _070380_);
  xor g_127377_(out[433], out[497], _070381_);
  and g_127378_(out[443], _049510_, _070382_);
  xor g_127379_(out[441], out[505], _070383_);
  xor g_127380_(out[432], out[496], _070384_);
  xor g_127381_(out[446], out[510], _070385_);
  xor g_127382_(out[436], out[500], _070386_);
  or g_127383_(_070385_, _070386_, _070387_);
  xor g_127384_(out[445], out[509], _070389_);
  xor g_127385_(out[435], out[499], _070390_);
  and g_127386_(_049466_, out[507], _070391_);
  xor g_127387_(out[438], out[502], _070392_);
  xor g_127388_(out[442], out[506], _070393_);
  xor g_127389_(out[437], out[501], _070394_);
  xor g_127390_(out[447], out[511], _070395_);
  xor g_127391_(out[440], out[504], _070396_);
  or g_127392_(_070389_, _070396_, _070397_);
  xor g_127393_(out[434], out[498], _070398_);
  or g_127394_(_070393_, _070398_, _070400_);
  or g_127395_(_070397_, _070400_, _070401_);
  or g_127396_(_070383_, _070390_, _070402_);
  or g_127397_(_070394_, _070402_, _070403_);
  or g_127398_(_070401_, _070403_, _070404_);
  or g_127399_(_070387_, _070404_, _070405_);
  xor g_127400_(out[444], out[508], _070406_);
  or g_127401_(_070391_, _070406_, _070407_);
  xor g_127402_(out[439], out[503], _070408_);
  or g_127403_(_070392_, _070408_, _070409_);
  or g_127404_(_070407_, _070409_, _070411_);
  or g_127405_(_070381_, _070382_, _070412_);
  or g_127406_(_070395_, _070412_, _070413_);
  or g_127407_(_070411_, _070413_, _070414_);
  or g_127408_(_070384_, _070414_, _070415_);
  or g_127409_(_070405_, _070415_, _070416_);
  xor g_127410_(out[423], out[503], _070417_);
  and g_127411_(_049455_, out[507], _070418_);
  xor g_127412_(out[430], out[510], _070419_);
  xor g_127413_(out[424], out[504], _070420_);
  xor g_127414_(out[417], out[497], _070422_);
  xor g_127415_(out[429], out[509], _070423_);
  xor g_127416_(out[425], out[505], _070424_);
  xor g_127417_(out[420], out[500], _070425_);
  xor g_127418_(out[418], out[498], _070426_);
  and g_127419_(out[427], _049510_, _070427_);
  xor g_127420_(out[419], out[499], _070428_);
  xor g_127421_(out[422], out[502], _070429_);
  xor g_127422_(out[431], out[511], _070430_);
  xor g_127423_(out[426], out[506], _070431_);
  xor g_127424_(out[421], out[501], _070433_);
  xor g_127425_(out[416], out[496], _070434_);
  or g_127426_(_070419_, _070425_, _070435_);
  or g_127427_(_070420_, _070423_, _070436_);
  or g_127428_(_070426_, _070431_, _070437_);
  or g_127429_(_070436_, _070437_, _070438_);
  or g_127430_(_070424_, _070428_, _070439_);
  or g_127431_(_070433_, _070434_, _070440_);
  or g_127432_(_070439_, _070440_, _070441_);
  or g_127433_(_070438_, _070441_, _070442_);
  xor g_127434_(out[428], out[508], _070444_);
  or g_127435_(_070418_, _070444_, _070445_);
  or g_127436_(_070417_, _070429_, _070446_);
  or g_127437_(_070445_, _070446_, _070447_);
  or g_127438_(_070422_, _070427_, _070448_);
  or g_127439_(_070430_, _070448_, _070449_);
  or g_127440_(_070447_, _070449_, _070450_);
  or g_127441_(_070442_, _070450_, _070451_);
  or g_127442_(_070435_, _070451_, _070452_);
  xor g_127443_(out[408], out[504], _070453_);
  xor g_127444_(out[405], out[501], _070455_);
  xor g_127445_(out[403], out[499], _070456_);
  xor g_127446_(out[414], out[510], _070457_);
  xor g_127447_(out[413], out[509], _070458_);
  xor g_127448_(out[402], out[498], _070459_);
  xor g_127449_(out[409], out[505], _070460_);
  xor g_127450_(out[406], out[502], _070461_);
  xor g_127451_(out[415], out[511], _070462_);
  xor g_127452_(out[410], out[506], _070463_);
  xor g_127453_(out[404], out[500], _070464_);
  xor g_127454_(out[400], out[496], _070466_);
  and g_127455_(_049444_, out[507], _070467_);
  and g_127456_(out[411], _049510_, _070468_);
  or g_127457_(_070453_, _070458_, _070469_);
  xor g_127458_(out[401], out[497], _070470_);
  or g_127459_(_070459_, _070463_, _070471_);
  or g_127460_(_070469_, _070471_, _070472_);
  or g_127461_(_070456_, _070460_, _070473_);
  or g_127462_(_070455_, _070473_, _070474_);
  or g_127463_(_070472_, _070474_, _070475_);
  or g_127464_(_070457_, _070464_, _070477_);
  or g_127465_(_070475_, _070477_, _070478_);
  xor g_127466_(out[412], out[508], _070479_);
  or g_127467_(_070467_, _070479_, _070480_);
  xor g_127468_(out[407], out[503], _070481_);
  or g_127469_(_070461_, _070481_, _070482_);
  or g_127470_(_070480_, _070482_, _070483_);
  or g_127471_(_070468_, _070470_, _070484_);
  or g_127472_(_070462_, _070484_, _070485_);
  or g_127473_(_070483_, _070485_, _070486_);
  or g_127474_(_070466_, _070486_, _070488_);
  or g_127475_(_070478_, _070488_, _070489_);
  not g_127476_(_070489_, _070490_);
  xor g_127477_(out[391], out[503], _070491_);
  and g_127478_(_049433_, out[507], _070492_);
  xor g_127479_(out[398], out[510], _070493_);
  xor g_127480_(out[392], out[504], _070494_);
  xor g_127481_(out[385], out[497], _070495_);
  xor g_127482_(out[397], out[509], _070496_);
  xor g_127483_(out[393], out[505], _070497_);
  xor g_127484_(out[388], out[500], _070499_);
  xor g_127485_(out[386], out[498], _070500_);
  and g_127486_(out[395], _049510_, _070501_);
  xor g_127487_(out[387], out[499], _070502_);
  xor g_127488_(out[390], out[502], _070503_);
  xor g_127489_(out[399], out[511], _070504_);
  xor g_127490_(out[394], out[506], _070505_);
  xor g_127491_(out[389], out[501], _070506_);
  xor g_127492_(out[384], out[496], _070507_);
  or g_127493_(_070493_, _070499_, _070508_);
  or g_127494_(_070494_, _070496_, _070510_);
  or g_127495_(_070500_, _070505_, _070511_);
  or g_127496_(_070510_, _070511_, _070512_);
  or g_127497_(_070497_, _070502_, _070513_);
  or g_127498_(_070506_, _070507_, _070514_);
  or g_127499_(_070513_, _070514_, _070515_);
  or g_127500_(_070512_, _070515_, _070516_);
  xor g_127501_(out[396], out[508], _070517_);
  or g_127502_(_070492_, _070517_, _070518_);
  or g_127503_(_070491_, _070503_, _070519_);
  or g_127504_(_070518_, _070519_, _070521_);
  or g_127505_(_070495_, _070501_, _070522_);
  or g_127506_(_070504_, _070522_, _070523_);
  or g_127507_(_070521_, _070523_, _070524_);
  or g_127508_(_070516_, _070524_, _070525_);
  or g_127509_(_070508_, _070525_, _070526_);
  xor g_127510_(out[378], out[506], _070527_);
  xor g_127511_(out[370], out[498], _070528_);
  xor g_127512_(out[369], out[497], _070529_);
  and g_127513_(_049422_, out[507], _070530_);
  and g_127514_(out[379], _049510_, _070532_);
  xor g_127515_(out[381], out[509], _070533_);
  xor g_127516_(out[371], out[499], _070534_);
  xor g_127517_(out[382], out[510], _070535_);
  xor g_127518_(out[380], out[508], _070536_);
  xor g_127519_(out[376], out[504], _070537_);
  xor g_127520_(out[383], out[511], _070538_);
  xor g_127521_(out[373], out[501], _070539_);
  xor g_127522_(out[374], out[502], _070540_);
  xor g_127523_(out[368], out[496], _070541_);
  xor g_127524_(out[372], out[500], _070543_);
  or g_127525_(_070533_, _070537_, _070544_);
  xor g_127526_(out[377], out[505], _070545_);
  or g_127527_(_070527_, _070528_, _070546_);
  or g_127528_(_070544_, _070546_, _070547_);
  or g_127529_(_070534_, _070545_, _070548_);
  or g_127530_(_070539_, _070548_, _070549_);
  or g_127531_(_070547_, _070549_, _070550_);
  or g_127532_(_070535_, _070543_, _070551_);
  or g_127533_(_070550_, _070551_, _070552_);
  or g_127534_(_070530_, _070536_, _070554_);
  xor g_127535_(out[375], out[503], _070555_);
  or g_127536_(_070540_, _070555_, _070556_);
  or g_127537_(_070554_, _070556_, _070557_);
  or g_127538_(_070529_, _070532_, _070558_);
  or g_127539_(_070538_, _070558_, _070559_);
  or g_127540_(_070557_, _070559_, _070560_);
  or g_127541_(_070541_, _070560_, _070561_);
  or g_127542_(_070552_, _070561_, _070562_);
  xor g_127543_(out[359], out[503], _070563_);
  and g_127544_(_049411_, out[507], _070565_);
  xor g_127545_(out[366], out[510], _070566_);
  xor g_127546_(out[360], out[504], _070567_);
  xor g_127547_(out[353], out[497], _070568_);
  xor g_127548_(out[365], out[509], _070569_);
  xor g_127549_(out[361], out[505], _070570_);
  xor g_127550_(out[356], out[500], _070571_);
  xor g_127551_(out[354], out[498], _070572_);
  and g_127552_(out[363], _049510_, _070573_);
  xor g_127553_(out[355], out[499], _070574_);
  xor g_127554_(out[358], out[502], _070576_);
  xor g_127555_(out[367], out[511], _070577_);
  xor g_127556_(out[362], out[506], _070578_);
  xor g_127557_(out[357], out[501], _070579_);
  xor g_127558_(out[352], out[496], _070580_);
  or g_127559_(_070566_, _070571_, _070581_);
  or g_127560_(_070567_, _070569_, _070582_);
  or g_127561_(_070572_, _070578_, _070583_);
  or g_127562_(_070582_, _070583_, _070584_);
  or g_127563_(_070570_, _070574_, _070585_);
  or g_127564_(_070579_, _070580_, _070587_);
  or g_127565_(_070585_, _070587_, _070588_);
  or g_127566_(_070584_, _070588_, _070589_);
  xor g_127567_(out[364], out[508], _070590_);
  or g_127568_(_070565_, _070590_, _070591_);
  or g_127569_(_070563_, _070576_, _070592_);
  or g_127570_(_070591_, _070592_, _070593_);
  or g_127571_(_070568_, _070573_, _070594_);
  or g_127572_(_070577_, _070594_, _070595_);
  or g_127573_(_070593_, _070595_, _070596_);
  or g_127574_(_070589_, _070596_, _070598_);
  or g_127575_(_070581_, _070598_, _070599_);
  and g_127576_(out[347], _049510_, _070600_);
  and g_127577_(_049400_, out[507], _070601_);
  xor g_127578_(out[344], out[504], _070602_);
  xor g_127579_(out[351], out[511], _070603_);
  xor g_127580_(out[337], out[497], _070604_);
  xor g_127581_(out[338], out[498], _070605_);
  xor g_127582_(out[340], out[500], _070606_);
  xor g_127583_(out[341], out[501], _070607_);
  xor g_127584_(out[345], out[505], _070609_);
  xor g_127585_(out[339], out[499], _070610_);
  xor g_127586_(out[350], out[510], _070611_);
  xor g_127587_(out[336], out[496], _070612_);
  xor g_127588_(out[346], out[506], _070613_);
  xor g_127589_(out[349], out[509], _070614_);
  or g_127590_(_070602_, _070614_, _070615_);
  xor g_127591_(out[342], out[502], _070616_);
  or g_127592_(_070605_, _070613_, _070617_);
  or g_127593_(_070615_, _070617_, _070618_);
  or g_127594_(_070609_, _070610_, _070620_);
  or g_127595_(_070607_, _070620_, _070621_);
  or g_127596_(_070618_, _070621_, _070622_);
  or g_127597_(_070606_, _070611_, _070623_);
  or g_127598_(_070622_, _070623_, _070624_);
  xor g_127599_(out[348], out[508], _070625_);
  or g_127600_(_070601_, _070625_, _070626_);
  xor g_127601_(out[343], out[503], _070627_);
  or g_127602_(_070616_, _070627_, _070628_);
  or g_127603_(_070626_, _070628_, _070629_);
  or g_127604_(_070600_, _070604_, _070631_);
  or g_127605_(_070603_, _070631_, _070632_);
  or g_127606_(_070629_, _070632_, _070633_);
  or g_127607_(_070612_, _070633_, _070634_);
  or g_127608_(_070624_, _070634_, _070635_);
  xor g_127609_(out[327], out[503], _070636_);
  and g_127610_(_098294_, out[507], _070637_);
  xor g_127611_(out[334], out[510], _070638_);
  xor g_127612_(out[328], out[504], _070639_);
  xor g_127613_(out[321], out[497], _070640_);
  xor g_127614_(out[333], out[509], _070642_);
  xor g_127615_(out[329], out[505], _070643_);
  xor g_127616_(out[324], out[500], _070644_);
  xor g_127617_(out[322], out[498], _070645_);
  and g_127618_(out[331], _049510_, _070646_);
  xor g_127619_(out[323], out[499], _070647_);
  xor g_127620_(out[326], out[502], _070648_);
  xor g_127621_(out[335], out[511], _070649_);
  xor g_127622_(out[330], out[506], _070650_);
  xor g_127623_(out[325], out[501], _070651_);
  xor g_127624_(out[320], out[496], _070653_);
  or g_127625_(_070638_, _070644_, _070654_);
  or g_127626_(_070639_, _070642_, _070655_);
  or g_127627_(_070645_, _070650_, _070656_);
  or g_127628_(_070655_, _070656_, _070657_);
  or g_127629_(_070643_, _070647_, _070658_);
  or g_127630_(_070651_, _070653_, _070659_);
  or g_127631_(_070658_, _070659_, _070660_);
  or g_127632_(_070657_, _070660_, _070661_);
  xor g_127633_(out[332], out[508], _070662_);
  or g_127634_(_070637_, _070662_, _070664_);
  or g_127635_(_070636_, _070648_, _070665_);
  or g_127636_(_070664_, _070665_, _070666_);
  or g_127637_(_070640_, _070646_, _070667_);
  or g_127638_(_070649_, _070667_, _070668_);
  or g_127639_(_070666_, _070668_, _070669_);
  or g_127640_(_070661_, _070669_, _070670_);
  or g_127641_(_070654_, _070670_, _070671_);
  not g_127642_(_070671_, _070672_);
  xor g_127643_(out[305], out[497], _070673_);
  and g_127644_(out[315], _049510_, _070675_);
  xor g_127645_(out[318], out[510], _070676_);
  xor g_127646_(out[307], out[499], _070677_);
  xor g_127647_(out[308], out[500], _070678_);
  xor g_127648_(out[306], out[498], _070679_);
  xor g_127649_(out[313], out[505], _070680_);
  xor g_127650_(out[304], out[496], _070681_);
  and g_127651_(_098283_, out[507], _070682_);
  xor g_127652_(out[310], out[502], _070683_);
  xor g_127653_(out[314], out[506], _070684_);
  xor g_127654_(out[309], out[501], _070686_);
  xor g_127655_(out[319], out[511], _070687_);
  xor g_127656_(out[317], out[509], _070688_);
  xor g_127657_(out[312], out[504], _070689_);
  or g_127658_(_070676_, _070678_, _070690_);
  or g_127659_(_070688_, _070689_, _070691_);
  or g_127660_(_070679_, _070684_, _070692_);
  or g_127661_(_070691_, _070692_, _070693_);
  or g_127662_(_070677_, _070680_, _070694_);
  or g_127663_(_070681_, _070686_, _070695_);
  or g_127664_(_070694_, _070695_, _070697_);
  or g_127665_(_070693_, _070697_, _070698_);
  xor g_127666_(out[316], out[508], _070699_);
  or g_127667_(_070682_, _070699_, _070700_);
  xor g_127668_(out[311], out[503], _070701_);
  or g_127669_(_070683_, _070701_, _070702_);
  or g_127670_(_070700_, _070702_, _070703_);
  or g_127671_(_070673_, _070675_, _070704_);
  or g_127672_(_070687_, _070704_, _070705_);
  or g_127673_(_070703_, _070705_, _070706_);
  or g_127674_(_070698_, _070706_, _070708_);
  or g_127675_(_070690_, _070708_, _070709_);
  xor g_127676_(out[295], out[503], _070710_);
  and g_127677_(_098272_, out[507], _070711_);
  xor g_127678_(out[302], out[510], _070712_);
  xor g_127679_(out[296], out[504], _070713_);
  xor g_127680_(out[289], out[497], _070714_);
  xor g_127681_(out[301], out[509], _070715_);
  xor g_127682_(out[297], out[505], _070716_);
  xor g_127683_(out[292], out[500], _070717_);
  xor g_127684_(out[290], out[498], _070719_);
  and g_127685_(out[299], _049510_, _070720_);
  xor g_127686_(out[291], out[499], _070721_);
  xor g_127687_(out[294], out[502], _070722_);
  xor g_127688_(out[303], out[511], _070723_);
  xor g_127689_(out[298], out[506], _070724_);
  xor g_127690_(out[293], out[501], _070725_);
  xor g_127691_(out[288], out[496], _070726_);
  or g_127692_(_070712_, _070717_, _070727_);
  or g_127693_(_070713_, _070715_, _070728_);
  or g_127694_(_070719_, _070724_, _070730_);
  or g_127695_(_070728_, _070730_, _070731_);
  or g_127696_(_070716_, _070721_, _070732_);
  or g_127697_(_070725_, _070726_, _070733_);
  or g_127698_(_070732_, _070733_, _070734_);
  or g_127699_(_070731_, _070734_, _070735_);
  xor g_127700_(out[300], out[508], _070736_);
  or g_127701_(_070711_, _070736_, _070737_);
  or g_127702_(_070710_, _070722_, _070738_);
  or g_127703_(_070737_, _070738_, _070739_);
  or g_127704_(_070714_, _070720_, _070741_);
  or g_127705_(_070723_, _070741_, _070742_);
  or g_127706_(_070739_, _070742_, _070743_);
  or g_127707_(_070735_, _070743_, _070744_);
  or g_127708_(_070727_, _070744_, _070745_);
  xor g_127709_(out[273], out[497], _070746_);
  and g_127710_(out[283], _049510_, _070747_);
  xor g_127711_(out[281], out[505], _070748_);
  xor g_127712_(out[272], out[496], _070749_);
  xor g_127713_(out[286], out[510], _070750_);
  xor g_127714_(out[276], out[500], _070752_);
  or g_127715_(_070750_, _070752_, _070753_);
  xor g_127716_(out[285], out[509], _070754_);
  xor g_127717_(out[275], out[499], _070755_);
  and g_127718_(_098261_, out[507], _070756_);
  xor g_127719_(out[278], out[502], _070757_);
  xor g_127720_(out[282], out[506], _070758_);
  xor g_127721_(out[277], out[501], _070759_);
  xor g_127722_(out[287], out[511], _070760_);
  xor g_127723_(out[280], out[504], _070761_);
  or g_127724_(_070754_, _070761_, _070763_);
  xor g_127725_(out[274], out[498], _070764_);
  or g_127726_(_070758_, _070764_, _070765_);
  or g_127727_(_070763_, _070765_, _070766_);
  or g_127728_(_070748_, _070755_, _070767_);
  or g_127729_(_070759_, _070767_, _070768_);
  or g_127730_(_070766_, _070768_, _070769_);
  or g_127731_(_070753_, _070769_, _070770_);
  xor g_127732_(out[284], out[508], _070771_);
  or g_127733_(_070756_, _070771_, _070772_);
  xor g_127734_(out[279], out[503], _070774_);
  or g_127735_(_070757_, _070774_, _070775_);
  or g_127736_(_070772_, _070775_, _070776_);
  or g_127737_(_070746_, _070747_, _070777_);
  or g_127738_(_070760_, _070777_, _070778_);
  or g_127739_(_070776_, _070778_, _070779_);
  or g_127740_(_070749_, _070779_, _070780_);
  or g_127741_(_070770_, _070780_, _070781_);
  xor g_127742_(out[263], out[503], _070782_);
  and g_127743_(_098250_, out[507], _070783_);
  xor g_127744_(out[270], out[510], _070785_);
  xor g_127745_(out[264], out[504], _070786_);
  xor g_127746_(out[257], out[497], _070787_);
  xor g_127747_(out[269], out[509], _070788_);
  xor g_127748_(out[265], out[505], _070789_);
  xor g_127749_(out[260], out[500], _070790_);
  xor g_127750_(out[258], out[498], _070791_);
  and g_127751_(out[267], _049510_, _070792_);
  xor g_127752_(out[259], out[499], _070793_);
  xor g_127753_(out[262], out[502], _070794_);
  xor g_127754_(out[271], out[511], _070796_);
  xor g_127755_(out[266], out[506], _070797_);
  xor g_127756_(out[261], out[501], _070798_);
  xor g_127757_(out[256], out[496], _070799_);
  or g_127758_(_070785_, _070790_, _070800_);
  or g_127759_(_070786_, _070788_, _070801_);
  or g_127760_(_070791_, _070797_, _070802_);
  or g_127761_(_070801_, _070802_, _070803_);
  or g_127762_(_070789_, _070793_, _070804_);
  or g_127763_(_070798_, _070799_, _070805_);
  or g_127764_(_070804_, _070805_, _070807_);
  or g_127765_(_070803_, _070807_, _070808_);
  xor g_127766_(out[268], out[508], _070809_);
  or g_127767_(_070783_, _070809_, _070810_);
  or g_127768_(_070782_, _070794_, _070811_);
  or g_127769_(_070810_, _070811_, _070812_);
  or g_127770_(_070787_, _070792_, _070813_);
  or g_127771_(_070796_, _070813_, _070814_);
  or g_127772_(_070812_, _070814_, _070815_);
  or g_127773_(_070808_, _070815_, _070816_);
  or g_127774_(_070800_, _070816_, _070818_);
  xor g_127775_(out[241], out[497], _070819_);
  and g_127776_(out[251], _049510_, _070820_);
  xor g_127777_(out[249], out[505], _070821_);
  xor g_127778_(out[240], out[496], _070822_);
  xor g_127779_(out[254], out[510], _070823_);
  xor g_127780_(out[244], out[500], _070824_);
  or g_127781_(_070823_, _070824_, _070825_);
  xor g_127782_(out[253], out[509], _070826_);
  xor g_127783_(out[243], out[499], _070827_);
  and g_127784_(_098239_, out[507], _070829_);
  xor g_127785_(out[246], out[502], _070830_);
  xor g_127786_(out[250], out[506], _070831_);
  xor g_127787_(out[245], out[501], _070832_);
  xor g_127788_(out[255], out[511], _070833_);
  xor g_127789_(out[248], out[504], _070834_);
  or g_127790_(_070826_, _070834_, _070835_);
  xor g_127791_(out[242], out[498], _070836_);
  or g_127792_(_070831_, _070836_, _070837_);
  or g_127793_(_070835_, _070837_, _070838_);
  or g_127794_(_070821_, _070827_, _070840_);
  or g_127795_(_070832_, _070840_, _070841_);
  or g_127796_(_070838_, _070841_, _070842_);
  or g_127797_(_070825_, _070842_, _070843_);
  xor g_127798_(out[252], out[508], _070844_);
  or g_127799_(_070829_, _070844_, _070845_);
  xor g_127800_(out[247], out[503], _070846_);
  or g_127801_(_070830_, _070846_, _070847_);
  or g_127802_(_070845_, _070847_, _070848_);
  or g_127803_(_070819_, _070820_, _070849_);
  or g_127804_(_070833_, _070849_, _070851_);
  or g_127805_(_070848_, _070851_, _070852_);
  or g_127806_(_070822_, _070852_, _070853_);
  or g_127807_(_070843_, _070853_, _070854_);
  xor g_127808_(out[231], out[503], _070855_);
  and g_127809_(_098228_, out[507], _070856_);
  xor g_127810_(out[238], out[510], _070857_);
  xor g_127811_(out[232], out[504], _070858_);
  xor g_127812_(out[225], out[497], _070859_);
  xor g_127813_(out[237], out[509], _070860_);
  xor g_127814_(out[233], out[505], _070862_);
  xor g_127815_(out[228], out[500], _070863_);
  xor g_127816_(out[226], out[498], _070864_);
  and g_127817_(out[235], _049510_, _070865_);
  xor g_127818_(out[227], out[499], _070866_);
  xor g_127819_(out[230], out[502], _070867_);
  xor g_127820_(out[239], out[511], _070868_);
  xor g_127821_(out[234], out[506], _070869_);
  xor g_127822_(out[229], out[501], _070870_);
  xor g_127823_(out[224], out[496], _070871_);
  or g_127824_(_070857_, _070863_, _070873_);
  or g_127825_(_070858_, _070860_, _070874_);
  or g_127826_(_070864_, _070869_, _070875_);
  or g_127827_(_070874_, _070875_, _070876_);
  or g_127828_(_070862_, _070866_, _070877_);
  or g_127829_(_070870_, _070871_, _070878_);
  or g_127830_(_070877_, _070878_, _070879_);
  or g_127831_(_070876_, _070879_, _070880_);
  xor g_127832_(out[236], out[508], _070881_);
  or g_127833_(_070856_, _070881_, _070882_);
  or g_127834_(_070855_, _070867_, _070884_);
  or g_127835_(_070882_, _070884_, _070885_);
  or g_127836_(_070859_, _070865_, _070886_);
  or g_127837_(_070868_, _070886_, _070887_);
  or g_127838_(_070885_, _070887_, _070888_);
  or g_127839_(_070880_, _070888_, _070889_);
  or g_127840_(_070873_, _070889_, _070890_);
  xor g_127841_(out[209], out[497], _070891_);
  and g_127842_(out[219], _049510_, _070892_);
  xor g_127843_(out[217], out[505], _070893_);
  xor g_127844_(out[208], out[496], _070895_);
  xor g_127845_(out[222], out[510], _070896_);
  xor g_127846_(out[212], out[500], _070897_);
  or g_127847_(_070896_, _070897_, _070898_);
  xor g_127848_(out[221], out[509], _070899_);
  xor g_127849_(out[211], out[499], _070900_);
  and g_127850_(_098217_, out[507], _070901_);
  xor g_127851_(out[214], out[502], _070902_);
  xor g_127852_(out[218], out[506], _070903_);
  xor g_127853_(out[213], out[501], _070904_);
  xor g_127854_(out[223], out[511], _070906_);
  xor g_127855_(out[216], out[504], _070907_);
  or g_127856_(_070899_, _070907_, _070908_);
  xor g_127857_(out[210], out[498], _070909_);
  or g_127858_(_070903_, _070909_, _070910_);
  or g_127859_(_070908_, _070910_, _070911_);
  or g_127860_(_070893_, _070900_, _070912_);
  or g_127861_(_070904_, _070912_, _070913_);
  or g_127862_(_070911_, _070913_, _070914_);
  or g_127863_(_070898_, _070914_, _070915_);
  xor g_127864_(out[220], out[508], _070917_);
  or g_127865_(_070901_, _070917_, _070918_);
  xor g_127866_(out[215], out[503], _070919_);
  or g_127867_(_070902_, _070919_, _070920_);
  or g_127868_(_070918_, _070920_, _070921_);
  or g_127869_(_070891_, _070892_, _070922_);
  or g_127870_(_070906_, _070922_, _070923_);
  or g_127871_(_070921_, _070923_, _070924_);
  or g_127872_(_070895_, _070924_, _070925_);
  or g_127873_(_070915_, _070925_, _070926_);
  xor g_127874_(out[199], out[503], _070928_);
  and g_127875_(_098206_, out[507], _070929_);
  xor g_127876_(out[206], out[510], _070930_);
  xor g_127877_(out[200], out[504], _070931_);
  xor g_127878_(out[193], out[497], _070932_);
  xor g_127879_(out[205], out[509], _070933_);
  xor g_127880_(out[201], out[505], _070934_);
  xor g_127881_(out[196], out[500], _070935_);
  xor g_127882_(out[194], out[498], _070936_);
  and g_127883_(out[203], _049510_, _070937_);
  xor g_127884_(out[195], out[499], _070939_);
  xor g_127885_(out[198], out[502], _070940_);
  xor g_127886_(out[207], out[511], _070941_);
  xor g_127887_(out[202], out[506], _070942_);
  xor g_127888_(out[197], out[501], _070943_);
  xor g_127889_(out[192], out[496], _070944_);
  or g_127890_(_070930_, _070935_, _070945_);
  or g_127891_(_070931_, _070933_, _070946_);
  or g_127892_(_070936_, _070942_, _070947_);
  or g_127893_(_070946_, _070947_, _070948_);
  or g_127894_(_070934_, _070939_, _070950_);
  or g_127895_(_070943_, _070944_, _070951_);
  or g_127896_(_070950_, _070951_, _070952_);
  or g_127897_(_070948_, _070952_, _070953_);
  xor g_127898_(out[204], out[508], _070954_);
  or g_127899_(_070929_, _070954_, _070955_);
  or g_127900_(_070928_, _070940_, _070956_);
  or g_127901_(_070955_, _070956_, _070957_);
  or g_127902_(_070932_, _070937_, _070958_);
  or g_127903_(_070941_, _070958_, _070959_);
  or g_127904_(_070957_, _070959_, _070961_);
  or g_127905_(_070953_, _070961_, _070962_);
  or g_127906_(_070945_, _070962_, _070963_);
  xor g_127907_(out[177], out[497], _070964_);
  and g_127908_(out[187], _049510_, _070965_);
  xor g_127909_(out[185], out[505], _070966_);
  xor g_127910_(out[176], out[496], _070967_);
  xor g_127911_(out[190], out[510], _070968_);
  xor g_127912_(out[180], out[500], _070969_);
  or g_127913_(_070968_, _070969_, _070970_);
  xor g_127914_(out[189], out[509], _070972_);
  xor g_127915_(out[179], out[499], _070973_);
  and g_127916_(_098195_, out[507], _070974_);
  xor g_127917_(out[182], out[502], _070975_);
  xor g_127918_(out[186], out[506], _070976_);
  xor g_127919_(out[181], out[501], _070977_);
  xor g_127920_(out[191], out[511], _070978_);
  xor g_127921_(out[184], out[504], _070979_);
  or g_127922_(_070972_, _070979_, _070980_);
  xor g_127923_(out[178], out[498], _070981_);
  or g_127924_(_070976_, _070981_, _070983_);
  or g_127925_(_070980_, _070983_, _070984_);
  or g_127926_(_070966_, _070973_, _070985_);
  or g_127927_(_070977_, _070985_, _070986_);
  or g_127928_(_070984_, _070986_, _070987_);
  or g_127929_(_070970_, _070987_, _070988_);
  xor g_127930_(out[188], out[508], _070989_);
  or g_127931_(_070974_, _070989_, _070990_);
  xor g_127932_(out[183], out[503], _070991_);
  or g_127933_(_070975_, _070991_, _070992_);
  or g_127934_(_070990_, _070992_, _070994_);
  or g_127935_(_070964_, _070965_, _070995_);
  or g_127936_(_070978_, _070995_, _070996_);
  or g_127937_(_070994_, _070996_, _070997_);
  or g_127938_(_070967_, _070997_, _070998_);
  or g_127939_(_070988_, _070998_, _070999_);
  xor g_127940_(out[167], out[503], _071000_);
  and g_127941_(_098184_, out[507], _071001_);
  xor g_127942_(out[174], out[510], _071002_);
  xor g_127943_(out[168], out[504], _071003_);
  xor g_127944_(out[161], out[497], _071005_);
  xor g_127945_(out[173], out[509], _071006_);
  xor g_127946_(out[169], out[505], _071007_);
  xor g_127947_(out[164], out[500], _071008_);
  xor g_127948_(out[162], out[498], _071009_);
  and g_127949_(out[171], _049510_, _071010_);
  xor g_127950_(out[163], out[499], _071011_);
  xor g_127951_(out[166], out[502], _071012_);
  xor g_127952_(out[175], out[511], _071013_);
  xor g_127953_(out[170], out[506], _071014_);
  xor g_127954_(out[165], out[501], _071016_);
  xor g_127955_(out[160], out[496], _071017_);
  or g_127956_(_071002_, _071008_, _071018_);
  or g_127957_(_071003_, _071006_, _071019_);
  or g_127958_(_071009_, _071014_, _071020_);
  or g_127959_(_071019_, _071020_, _071021_);
  or g_127960_(_071007_, _071011_, _071022_);
  or g_127961_(_071016_, _071017_, _071023_);
  or g_127962_(_071022_, _071023_, _071024_);
  or g_127963_(_071021_, _071024_, _071025_);
  xor g_127964_(out[172], out[508], _071027_);
  or g_127965_(_071001_, _071027_, _071028_);
  or g_127966_(_071000_, _071012_, _071029_);
  or g_127967_(_071028_, _071029_, _071030_);
  or g_127968_(_071005_, _071010_, _071031_);
  or g_127969_(_071013_, _071031_, _071032_);
  or g_127970_(_071030_, _071032_, _071033_);
  or g_127971_(_071025_, _071033_, _071034_);
  or g_127972_(_071018_, _071034_, _071035_);
  and g_127973_(out[155], _049510_, _071036_);
  xor g_127974_(out[148], out[500], _071038_);
  xor g_127975_(out[158], out[510], _071039_);
  or g_127976_(_071038_, _071039_, _071040_);
  xor g_127977_(out[157], out[509], _071041_);
  xor g_127978_(out[147], out[499], _071042_);
  xor g_127979_(out[144], out[496], _071043_);
  and g_127980_(_098173_, out[507], _071044_);
  xor g_127981_(out[154], out[506], _071045_);
  xor g_127982_(out[159], out[511], _071046_);
  xor g_127983_(out[150], out[502], _071047_);
  xor g_127984_(out[149], out[501], _071049_);
  xor g_127985_(out[152], out[504], _071050_);
  or g_127986_(_071041_, _071050_, _071051_);
  xor g_127987_(out[146], out[498], _071052_);
  xor g_127988_(out[153], out[505], _071053_);
  xor g_127989_(out[145], out[497], _071054_);
  or g_127990_(_071045_, _071052_, _071055_);
  or g_127991_(_071051_, _071055_, _071056_);
  or g_127992_(_071042_, _071053_, _071057_);
  or g_127993_(_071049_, _071057_, _071058_);
  or g_127994_(_071056_, _071058_, _071060_);
  or g_127995_(_071040_, _071060_, _071061_);
  xor g_127996_(out[156], out[508], _071062_);
  or g_127997_(_071044_, _071062_, _071063_);
  xor g_127998_(out[151], out[503], _071064_);
  or g_127999_(_071047_, _071064_, _071065_);
  or g_128000_(_071063_, _071065_, _071066_);
  or g_128001_(_071036_, _071054_, _071067_);
  or g_128002_(_071046_, _071067_, _071068_);
  or g_128003_(_071066_, _071068_, _071069_);
  or g_128004_(_071043_, _071069_, _071071_);
  or g_128005_(_071061_, _071071_, _071072_);
  xor g_128006_(out[135], out[503], _071073_);
  and g_128007_(_098162_, out[507], _071074_);
  xor g_128008_(out[142], out[510], _071075_);
  xor g_128009_(out[136], out[504], _071076_);
  xor g_128010_(out[129], out[497], _071077_);
  xor g_128011_(out[141], out[509], _071078_);
  xor g_128012_(out[137], out[505], _071079_);
  xor g_128013_(out[132], out[500], _071080_);
  xor g_128014_(out[130], out[498], _071082_);
  and g_128015_(out[139], _049510_, _071083_);
  xor g_128016_(out[131], out[499], _071084_);
  xor g_128017_(out[134], out[502], _071085_);
  xor g_128018_(out[143], out[511], _071086_);
  xor g_128019_(out[138], out[506], _071087_);
  xor g_128020_(out[133], out[501], _071088_);
  xor g_128021_(out[128], out[496], _071089_);
  or g_128022_(_071075_, _071080_, _071090_);
  or g_128023_(_071076_, _071078_, _071091_);
  or g_128024_(_071082_, _071087_, _071093_);
  or g_128025_(_071091_, _071093_, _071094_);
  or g_128026_(_071079_, _071084_, _071095_);
  or g_128027_(_071088_, _071089_, _071096_);
  or g_128028_(_071095_, _071096_, _071097_);
  or g_128029_(_071094_, _071097_, _071098_);
  xor g_128030_(out[140], out[508], _071099_);
  or g_128031_(_071074_, _071099_, _071100_);
  or g_128032_(_071073_, _071085_, _071101_);
  or g_128033_(_071100_, _071101_, _071102_);
  or g_128034_(_071077_, _071083_, _071104_);
  or g_128035_(_071086_, _071104_, _071105_);
  or g_128036_(_071102_, _071105_, _071106_);
  or g_128037_(_071098_, _071106_, _071107_);
  or g_128038_(_071090_, _071107_, _071108_);
  xor g_128039_(out[113], out[497], _071109_);
  and g_128040_(out[123], _049510_, _071110_);
  xor g_128041_(out[121], out[505], _071111_);
  xor g_128042_(out[112], out[496], _071112_);
  xor g_128043_(out[126], out[510], _071113_);
  xor g_128044_(out[116], out[500], _071115_);
  or g_128045_(_071113_, _071115_, _071116_);
  xor g_128046_(out[125], out[509], _071117_);
  xor g_128047_(out[115], out[499], _071118_);
  and g_128048_(_098151_, out[507], _071119_);
  xor g_128049_(out[118], out[502], _071120_);
  xor g_128050_(out[122], out[506], _071121_);
  xor g_128051_(out[117], out[501], _071122_);
  xor g_128052_(out[127], out[511], _071123_);
  xor g_128053_(out[120], out[504], _071124_);
  or g_128054_(_071117_, _071124_, _071126_);
  xor g_128055_(out[114], out[498], _071127_);
  or g_128056_(_071121_, _071127_, _071128_);
  or g_128057_(_071126_, _071128_, _071129_);
  or g_128058_(_071111_, _071118_, _071130_);
  or g_128059_(_071122_, _071130_, _071131_);
  or g_128060_(_071129_, _071131_, _071132_);
  or g_128061_(_071116_, _071132_, _071133_);
  xor g_128062_(out[124], out[508], _071134_);
  or g_128063_(_071119_, _071134_, _071135_);
  xor g_128064_(out[119], out[503], _071137_);
  or g_128065_(_071120_, _071137_, _071138_);
  or g_128066_(_071135_, _071138_, _071139_);
  or g_128067_(_071109_, _071110_, _071140_);
  or g_128068_(_071123_, _071140_, _071141_);
  or g_128069_(_071139_, _071141_, _071142_);
  or g_128070_(_071112_, _071142_, _071143_);
  or g_128071_(_071133_, _071143_, _071144_);
  xor g_128072_(out[103], out[503], _071145_);
  and g_128073_(_098140_, out[507], _071146_);
  xor g_128074_(out[110], out[510], _071148_);
  xor g_128075_(out[104], out[504], _071149_);
  xor g_128076_(out[97], out[497], _071150_);
  xor g_128077_(out[109], out[509], _071151_);
  xor g_128078_(out[105], out[505], _071152_);
  xor g_128079_(out[100], out[500], _071153_);
  xor g_128080_(out[98], out[498], _071154_);
  and g_128081_(out[107], _049510_, _071155_);
  xor g_128082_(out[99], out[499], _071156_);
  xor g_128083_(out[102], out[502], _071157_);
  xor g_128084_(out[111], out[511], _071159_);
  xor g_128085_(out[106], out[506], _071160_);
  xor g_128086_(out[101], out[501], _071161_);
  xor g_128087_(out[96], out[496], _071162_);
  or g_128088_(_071148_, _071153_, _071163_);
  or g_128089_(_071149_, _071151_, _071164_);
  or g_128090_(_071154_, _071160_, _071165_);
  or g_128091_(_071164_, _071165_, _071166_);
  or g_128092_(_071152_, _071156_, _071167_);
  or g_128093_(_071161_, _071162_, _071168_);
  or g_128094_(_071167_, _071168_, _071170_);
  or g_128095_(_071166_, _071170_, _071171_);
  xor g_128096_(out[108], out[508], _071172_);
  or g_128097_(_071146_, _071172_, _071173_);
  or g_128098_(_071145_, _071157_, _071174_);
  or g_128099_(_071173_, _071174_, _071175_);
  or g_128100_(_071150_, _071155_, _071176_);
  or g_128101_(_071159_, _071176_, _071177_);
  or g_128102_(_071175_, _071177_, _071178_);
  or g_128103_(_071171_, _071178_, _071179_);
  or g_128104_(_071163_, _071179_, _071181_);
  xor g_128105_(out[81], out[497], _071182_);
  and g_128106_(out[91], _049510_, _071183_);
  xor g_128107_(out[94], out[510], _071184_);
  xor g_128108_(out[83], out[499], _071185_);
  xor g_128109_(out[84], out[500], _071186_);
  xor g_128110_(out[82], out[498], _071187_);
  xor g_128111_(out[89], out[505], _071188_);
  xor g_128112_(out[80], out[496], _071189_);
  and g_128113_(_098129_, out[507], _071190_);
  xor g_128114_(out[86], out[502], _071192_);
  xor g_128115_(out[90], out[506], _071193_);
  xor g_128116_(out[85], out[501], _071194_);
  xor g_128117_(out[95], out[511], _071195_);
  xor g_128118_(out[93], out[509], _071196_);
  xor g_128119_(out[88], out[504], _071197_);
  or g_128120_(_071184_, _071186_, _071198_);
  or g_128121_(_071196_, _071197_, _071199_);
  or g_128122_(_071187_, _071193_, _071200_);
  or g_128123_(_071199_, _071200_, _071201_);
  or g_128124_(_071185_, _071188_, _071203_);
  or g_128125_(_071189_, _071194_, _071204_);
  or g_128126_(_071203_, _071204_, _071205_);
  or g_128127_(_071201_, _071205_, _071206_);
  xor g_128128_(out[92], out[508], _071207_);
  or g_128129_(_071190_, _071207_, _071208_);
  xor g_128130_(out[87], out[503], _071209_);
  or g_128131_(_071192_, _071209_, _071210_);
  or g_128132_(_071208_, _071210_, _071211_);
  or g_128133_(_071182_, _071183_, _071212_);
  or g_128134_(_071195_, _071212_, _071214_);
  or g_128135_(_071211_, _071214_, _071215_);
  or g_128136_(_071206_, _071215_, _071216_);
  or g_128137_(_071198_, _071216_, _071217_);
  xor g_128138_(out[71], out[503], _071218_);
  and g_128139_(_098118_, out[507], _071219_);
  xor g_128140_(out[78], out[510], _071220_);
  xor g_128141_(out[72], out[504], _071221_);
  xor g_128142_(out[65], out[497], _071222_);
  xor g_128143_(out[77], out[509], _071223_);
  xor g_128144_(out[73], out[505], _071225_);
  xor g_128145_(out[68], out[500], _071226_);
  xor g_128146_(out[66], out[498], _071227_);
  and g_128147_(out[75], _049510_, _071228_);
  xor g_128148_(out[67], out[499], _071229_);
  xor g_128149_(out[70], out[502], _071230_);
  xor g_128150_(out[79], out[511], _071231_);
  xor g_128151_(out[74], out[506], _071232_);
  xor g_128152_(out[69], out[501], _071233_);
  xor g_128153_(out[64], out[496], _071234_);
  or g_128154_(_071220_, _071226_, _071236_);
  or g_128155_(_071221_, _071223_, _071237_);
  or g_128156_(_071227_, _071232_, _071238_);
  or g_128157_(_071237_, _071238_, _071239_);
  or g_128158_(_071225_, _071229_, _071240_);
  or g_128159_(_071233_, _071234_, _071241_);
  or g_128160_(_071240_, _071241_, _071242_);
  or g_128161_(_071239_, _071242_, _071243_);
  xor g_128162_(out[76], out[508], _071244_);
  or g_128163_(_071219_, _071244_, _071245_);
  or g_128164_(_071218_, _071230_, _071247_);
  or g_128165_(_071245_, _071247_, _071248_);
  or g_128166_(_071222_, _071228_, _071249_);
  or g_128167_(_071231_, _071249_, _071250_);
  or g_128168_(_071248_, _071250_, _071251_);
  or g_128169_(_071243_, _071251_, _071252_);
  or g_128170_(_071236_, _071252_, _071253_);
  xor g_128171_(out[50], out[498], _071254_);
  xor g_128172_(out[48], out[496], _071255_);
  xor g_128173_(out[57], out[505], _071256_);
  xor g_128174_(out[56], out[504], _071258_);
  xor g_128175_(out[53], out[501], _071259_);
  xor g_128176_(out[62], out[510], _071260_);
  xor g_128177_(out[61], out[509], _071261_);
  xor g_128178_(out[63], out[511], _071262_);
  xor g_128179_(out[58], out[506], _071263_);
  xor g_128180_(out[54], out[502], _071264_);
  xor g_128181_(out[51], out[499], _071265_);
  and g_128182_(_098107_, out[507], _071266_);
  and g_128183_(out[59], _049510_, _071267_);
  xor g_128184_(out[52], out[500], _071269_);
  xor g_128185_(out[49], out[497], _071270_);
  or g_128186_(_071260_, _071269_, _071271_);
  or g_128187_(_071258_, _071261_, _071272_);
  or g_128188_(_071254_, _071263_, _071273_);
  or g_128189_(_071272_, _071273_, _071274_);
  or g_128190_(_071256_, _071265_, _071275_);
  or g_128191_(_071255_, _071259_, _071276_);
  or g_128192_(_071275_, _071276_, _071277_);
  or g_128193_(_071274_, _071277_, _071278_);
  xor g_128194_(out[60], out[508], _071280_);
  or g_128195_(_071266_, _071280_, _071281_);
  xor g_128196_(out[55], out[503], _071282_);
  or g_128197_(_071264_, _071282_, _071283_);
  or g_128198_(_071281_, _071283_, _071284_);
  or g_128199_(_071267_, _071270_, _071285_);
  or g_128200_(_071262_, _071285_, _071286_);
  or g_128201_(_071284_, _071286_, _071287_);
  or g_128202_(_071278_, _071287_, _071288_);
  or g_128203_(_071271_, _071288_, _071289_);
  xor g_128204_(out[39], out[503], _071291_);
  and g_128205_(_098096_, out[507], _071292_);
  xor g_128206_(out[46], out[510], _071293_);
  xor g_128207_(out[40], out[504], _071294_);
  xor g_128208_(out[33], out[497], _071295_);
  xor g_128209_(out[45], out[509], _071296_);
  xor g_128210_(out[41], out[505], _071297_);
  xor g_128211_(out[36], out[500], _071298_);
  xor g_128212_(out[34], out[498], _071299_);
  and g_128213_(out[43], _049510_, _071300_);
  xor g_128214_(out[35], out[499], _071302_);
  xor g_128215_(out[38], out[502], _071303_);
  xor g_128216_(out[47], out[511], _071304_);
  xor g_128217_(out[42], out[506], _071305_);
  xor g_128218_(out[37], out[501], _071306_);
  xor g_128219_(out[32], out[496], _071307_);
  or g_128220_(_071293_, _071298_, _071308_);
  or g_128221_(_071294_, _071296_, _071309_);
  or g_128222_(_071299_, _071305_, _071310_);
  or g_128223_(_071309_, _071310_, _071311_);
  or g_128224_(_071297_, _071302_, _071313_);
  or g_128225_(_071306_, _071307_, _071314_);
  or g_128226_(_071313_, _071314_, _071315_);
  or g_128227_(_071311_, _071315_, _071316_);
  xor g_128228_(out[44], out[508], _071317_);
  or g_128229_(_071292_, _071317_, _071318_);
  or g_128230_(_071291_, _071303_, _071319_);
  or g_128231_(_071318_, _071319_, _071320_);
  or g_128232_(_071295_, _071300_, _071321_);
  or g_128233_(_071304_, _071321_, _071322_);
  or g_128234_(_071320_, _071322_, _071324_);
  or g_128235_(_071316_, _071324_, _071325_);
  or g_128236_(_071308_, _071325_, _071326_);
  xor g_128237_(out[17], out[497], _071327_);
  and g_128238_(out[27], _049510_, _071328_);
  xor g_128239_(out[25], out[505], _071329_);
  xor g_128240_(out[16], out[496], _071330_);
  xor g_128241_(out[30], out[510], _071331_);
  xor g_128242_(out[20], out[500], _071332_);
  or g_128243_(_071331_, _071332_, _071333_);
  xor g_128244_(out[29], out[509], _071335_);
  xor g_128245_(out[19], out[499], _071336_);
  and g_128246_(_098063_, out[507], _071337_);
  xor g_128247_(out[22], out[502], _071338_);
  xor g_128248_(out[26], out[506], _071339_);
  xor g_128249_(out[21], out[501], _071340_);
  xor g_128250_(out[31], out[511], _071341_);
  xor g_128251_(out[24], out[504], _071342_);
  or g_128252_(_071335_, _071342_, _071343_);
  xor g_128253_(out[18], out[498], _071344_);
  or g_128254_(_071339_, _071344_, _071346_);
  or g_128255_(_071343_, _071346_, _071347_);
  or g_128256_(_071329_, _071336_, _071348_);
  or g_128257_(_071340_, _071348_, _071349_);
  or g_128258_(_071347_, _071349_, _071350_);
  or g_128259_(_071333_, _071350_, _071351_);
  xor g_128260_(out[28], out[508], _071352_);
  or g_128261_(_071337_, _071352_, _071353_);
  xor g_128262_(out[23], out[503], _071354_);
  or g_128263_(_071338_, _071354_, _071355_);
  or g_128264_(_071353_, _071355_, _071357_);
  or g_128265_(_071327_, _071328_, _071358_);
  or g_128266_(_071341_, _071358_, _071359_);
  or g_128267_(_071357_, _071359_, _071360_);
  or g_128268_(_071330_, _071360_, _071361_);
  or g_128269_(_071351_, _071361_, _071362_);
  not g_128270_(_071362_, _071363_);
  xor g_128271_(out[1], out[497], _071364_);
  and g_128272_(_098041_, out[507], _071365_);
  and g_128273_(out[11], _049510_, _071366_);
  xor g_128274_(out[8], out[504], _071368_);
  xor g_128275_(out[10], out[506], _071369_);
  xor g_128276_(out[2], out[498], _071370_);
  xor g_128277_(out[4], out[500], _071371_);
  xor g_128278_(out[5], out[501], _071372_);
  xor g_128279_(out[9], out[505], _071373_);
  xor g_128280_(out[3], out[499], _071374_);
  xor g_128281_(out[14], out[510], _071375_);
  xor g_128282_(out[0], out[496], _071376_);
  xor g_128283_(out[15], out[511], _071377_);
  xor g_128284_(out[13], out[509], _071379_);
  or g_128285_(_071368_, _071379_, _071380_);
  xor g_128286_(out[6], out[502], _071381_);
  or g_128287_(_071369_, _071370_, _071382_);
  or g_128288_(_071380_, _071382_, _071383_);
  or g_128289_(_071373_, _071374_, _071384_);
  or g_128290_(_071372_, _071384_, _071385_);
  or g_128291_(_071383_, _071385_, _071386_);
  or g_128292_(_071371_, _071375_, _071387_);
  or g_128293_(_071386_, _071387_, _071388_);
  xor g_128294_(out[12], out[508], _071390_);
  or g_128295_(_071365_, _071390_, _071391_);
  xor g_128296_(out[7], out[503], _071392_);
  or g_128297_(_071381_, _071392_, _071393_);
  or g_128298_(_071391_, _071393_, _071394_);
  or g_128299_(_071364_, _071366_, _071395_);
  or g_128300_(_071377_, _071395_, _071396_);
  or g_128301_(_071394_, _071396_, _071397_);
  or g_128302_(_071376_, _071397_, _071398_);
  or g_128303_(_071388_, _071398_, _071399_);
  xor g_128304_(out[481], out[465], _071401_);
  and g_128305_(_098030_, out[475], _071402_);
  and g_128306_(out[491], _049499_, _071403_);
  xor g_128307_(out[489], out[473], _071404_);
  xor g_128308_(out[480], out[464], _071405_);
  xor g_128309_(out[494], out[478], _071406_);
  xor g_128310_(out[484], out[468], _071407_);
  or g_128311_(_071406_, _071407_, _071408_);
  xor g_128312_(out[493], out[477], _071409_);
  xor g_128313_(out[483], out[467], _071410_);
  xor g_128314_(out[492], out[476], _071412_);
  xor g_128315_(out[486], out[470], _071413_);
  xor g_128316_(out[490], out[474], _071414_);
  xor g_128317_(out[485], out[469], _071415_);
  xor g_128318_(out[495], out[479], _071416_);
  xor g_128319_(out[488], out[472], _071417_);
  or g_128320_(_071409_, _071417_, _071418_);
  xor g_128321_(out[482], out[466], _071419_);
  or g_128322_(_071414_, _071419_, _071420_);
  or g_128323_(_071418_, _071420_, _071421_);
  or g_128324_(_071404_, _071410_, _071423_);
  or g_128325_(_071415_, _071423_, _071424_);
  or g_128326_(_071421_, _071424_, _071425_);
  or g_128327_(_071408_, _071425_, _071426_);
  or g_128328_(_071402_, _071412_, _071427_);
  xor g_128329_(out[487], out[471], _071428_);
  or g_128330_(_071413_, _071428_, _071429_);
  or g_128331_(_071427_, _071429_, _071430_);
  or g_128332_(_071401_, _071403_, _071431_);
  or g_128333_(_071416_, _071431_, _071432_);
  or g_128334_(_071430_, _071432_, _071434_);
  or g_128335_(_071405_, _071434_, _071435_);
  or g_128336_(_071426_, _071435_, _071436_);
  xor g_128337_(out[490], out[458], _071437_);
  xor g_128338_(out[488], out[456], _071438_);
  xor g_128339_(out[481], out[449], _071439_);
  and g_128340_(_098030_, out[459], _071440_);
  and g_128341_(out[491], _049477_, _071441_);
  xor g_128342_(out[482], out[450], _071442_);
  xor g_128343_(out[485], out[453], _071443_);
  xor g_128344_(out[489], out[457], _071445_);
  xor g_128345_(out[492], out[460], _071446_);
  xor g_128346_(out[493], out[461], _071447_);
  xor g_128347_(out[495], out[463], _071448_);
  xor g_128348_(out[484], out[452], _071449_);
  xor g_128349_(out[486], out[454], _071450_);
  xor g_128350_(out[483], out[451], _071451_);
  xor g_128351_(out[480], out[448], _071452_);
  xor g_128352_(out[494], out[462], _071453_);
  or g_128353_(_071449_, _071453_, _071454_);
  or g_128354_(_071438_, _071447_, _071456_);
  or g_128355_(_071437_, _071442_, _071457_);
  or g_128356_(_071456_, _071457_, _071458_);
  or g_128357_(_071445_, _071451_, _071459_);
  or g_128358_(_071443_, _071452_, _071460_);
  or g_128359_(_071459_, _071460_, _071461_);
  or g_128360_(_071458_, _071461_, _071462_);
  or g_128361_(_071440_, _071446_, _071463_);
  xor g_128362_(out[487], out[455], _071464_);
  or g_128363_(_071450_, _071464_, _071465_);
  or g_128364_(_071463_, _071465_, _071467_);
  or g_128365_(_071439_, _071441_, _071468_);
  or g_128366_(_071448_, _071468_, _071469_);
  or g_128367_(_071467_, _071469_, _071470_);
  or g_128368_(_071462_, _071470_, _071471_);
  or g_128369_(_071454_, _071471_, _071472_);
  not g_128370_(_071472_, _071473_);
  xor g_128371_(out[481], out[433], _071474_);
  and g_128372_(out[491], _049466_, _071475_);
  xor g_128373_(out[489], out[441], _071476_);
  xor g_128374_(out[480], out[432], _071478_);
  xor g_128375_(out[494], out[446], _071479_);
  xor g_128376_(out[484], out[436], _071480_);
  or g_128377_(_071479_, _071480_, _071481_);
  xor g_128378_(out[493], out[445], _071482_);
  xor g_128379_(out[483], out[435], _071483_);
  and g_128380_(_098030_, out[443], _071484_);
  xor g_128381_(out[486], out[438], _071485_);
  xor g_128382_(out[490], out[442], _071486_);
  xor g_128383_(out[485], out[437], _071487_);
  xor g_128384_(out[495], out[447], _071489_);
  xor g_128385_(out[488], out[440], _071490_);
  or g_128386_(_071482_, _071490_, _071491_);
  xor g_128387_(out[482], out[434], _071492_);
  or g_128388_(_071486_, _071492_, _071493_);
  or g_128389_(_071491_, _071493_, _071494_);
  or g_128390_(_071476_, _071483_, _071495_);
  or g_128391_(_071487_, _071495_, _071496_);
  or g_128392_(_071494_, _071496_, _071497_);
  or g_128393_(_071481_, _071497_, _071498_);
  not g_128394_(_071498_, _071500_);
  xor g_128395_(out[492], out[444], _071501_);
  or g_128396_(_071484_, _071501_, _071502_);
  xor g_128397_(out[487], out[439], _071503_);
  or g_128398_(_071485_, _071503_, _071504_);
  or g_128399_(_071502_, _071504_, _071505_);
  or g_128400_(_071474_, _071475_, _071506_);
  or g_128401_(_071489_, _071506_, _071507_);
  or g_128402_(_071505_, _071507_, _071508_);
  or g_128403_(_071478_, _071508_, _071509_);
  not g_128404_(_071509_, _071511_);
  and g_128405_(_071500_, _071511_, _071512_);
  not g_128406_(_071512_, _071513_);
  xor g_128407_(out[481], out[417], _071514_);
  and g_128408_(out[491], _049455_, _071515_);
  xor g_128409_(out[494], out[430], _071516_);
  xor g_128410_(out[483], out[419], _071517_);
  xor g_128411_(out[484], out[420], _071518_);
  xor g_128412_(out[482], out[418], _071519_);
  xor g_128413_(out[489], out[425], _071520_);
  xor g_128414_(out[480], out[416], _071522_);
  and g_128415_(_098030_, out[427], _071523_);
  xor g_128416_(out[486], out[422], _071524_);
  xor g_128417_(out[490], out[426], _071525_);
  xor g_128418_(out[485], out[421], _071526_);
  xor g_128419_(out[495], out[431], _071527_);
  xor g_128420_(out[493], out[429], _071528_);
  xor g_128421_(out[488], out[424], _071529_);
  or g_128422_(_071516_, _071518_, _071530_);
  or g_128423_(_071528_, _071529_, _071531_);
  or g_128424_(_071519_, _071525_, _071533_);
  or g_128425_(_071531_, _071533_, _071534_);
  or g_128426_(_071517_, _071520_, _071535_);
  or g_128427_(_071522_, _071526_, _071536_);
  or g_128428_(_071535_, _071536_, _071537_);
  or g_128429_(_071534_, _071537_, _071538_);
  xor g_128430_(out[492], out[428], _071539_);
  or g_128431_(_071523_, _071539_, _071540_);
  xor g_128432_(out[487], out[423], _071541_);
  or g_128433_(_071524_, _071541_, _071542_);
  or g_128434_(_071540_, _071542_, _071544_);
  or g_128435_(_071514_, _071515_, _071545_);
  or g_128436_(_071527_, _071545_, _071546_);
  or g_128437_(_071544_, _071546_, _071547_);
  or g_128438_(_071538_, _071547_, _071548_);
  or g_128439_(_071530_, _071548_, _071549_);
  not g_128440_(_071549_, _071550_);
  xor g_128441_(out[481], out[401], _071551_);
  and g_128442_(out[491], _049444_, _071552_);
  xor g_128443_(out[489], out[409], _071553_);
  xor g_128444_(out[480], out[400], _071555_);
  xor g_128445_(out[494], out[414], _071556_);
  xor g_128446_(out[484], out[404], _071557_);
  or g_128447_(_071556_, _071557_, _071558_);
  xor g_128448_(out[493], out[413], _071559_);
  xor g_128449_(out[483], out[403], _071560_);
  and g_128450_(_098030_, out[411], _071561_);
  xor g_128451_(out[486], out[406], _071562_);
  xor g_128452_(out[490], out[410], _071563_);
  xor g_128453_(out[485], out[405], _071564_);
  xor g_128454_(out[495], out[415], _071566_);
  xor g_128455_(out[488], out[408], _071567_);
  or g_128456_(_071559_, _071567_, _071568_);
  xor g_128457_(out[482], out[402], _071569_);
  or g_128458_(_071563_, _071569_, _071570_);
  or g_128459_(_071568_, _071570_, _071571_);
  or g_128460_(_071553_, _071560_, _071572_);
  or g_128461_(_071564_, _071572_, _071573_);
  or g_128462_(_071571_, _071573_, _071574_);
  or g_128463_(_071558_, _071574_, _071575_);
  xor g_128464_(out[492], out[412], _071577_);
  or g_128465_(_071561_, _071577_, _071578_);
  xor g_128466_(out[487], out[407], _071579_);
  or g_128467_(_071562_, _071579_, _071580_);
  or g_128468_(_071578_, _071580_, _071581_);
  or g_128469_(_071551_, _071552_, _071582_);
  or g_128470_(_071566_, _071582_, _071583_);
  or g_128471_(_071581_, _071583_, _071584_);
  or g_128472_(_071555_, _071584_, _071585_);
  or g_128473_(_071575_, _071585_, _071586_);
  not g_128474_(_071586_, _071588_);
  and g_128475_(out[491], _049433_, _071589_);
  and g_128476_(_098030_, out[395], _071590_);
  xor g_128477_(out[488], out[392], _071591_);
  xor g_128478_(out[495], out[399], _071592_);
  xor g_128479_(out[481], out[385], _071593_);
  xor g_128480_(out[482], out[386], _071594_);
  xor g_128481_(out[484], out[388], _071595_);
  xor g_128482_(out[493], out[397], _071596_);
  xor g_128483_(out[489], out[393], _071597_);
  xor g_128484_(out[483], out[387], _071599_);
  xor g_128485_(out[485], out[389], _071600_);
  xor g_128486_(out[494], out[398], _071601_);
  xor g_128487_(out[480], out[384], _071602_);
  xor g_128488_(out[490], out[394], _071603_);
  or g_128489_(_071591_, _071596_, _071604_);
  xor g_128490_(out[486], out[390], _071605_);
  or g_128491_(_071594_, _071603_, _071606_);
  or g_128492_(_071604_, _071606_, _071607_);
  or g_128493_(_071597_, _071599_, _071608_);
  or g_128494_(_071600_, _071608_, _071610_);
  or g_128495_(_071607_, _071610_, _071611_);
  or g_128496_(_071595_, _071601_, _071612_);
  or g_128497_(_071611_, _071612_, _071613_);
  xor g_128498_(out[492], out[396], _071614_);
  or g_128499_(_071590_, _071614_, _071615_);
  xor g_128500_(out[487], out[391], _071616_);
  or g_128501_(_071605_, _071616_, _071617_);
  or g_128502_(_071615_, _071617_, _071618_);
  or g_128503_(_071589_, _071593_, _071619_);
  or g_128504_(_071592_, _071619_, _071621_);
  or g_128505_(_071618_, _071621_, _071622_);
  or g_128506_(_071602_, _071622_, _071623_);
  or g_128507_(_071613_, _071623_, _071624_);
  not g_128508_(_071624_, _071625_);
  xor g_128509_(out[481], out[369], _071626_);
  and g_128510_(out[491], _049422_, _071627_);
  xor g_128511_(out[489], out[377], _071628_);
  xor g_128512_(out[480], out[368], _071629_);
  xor g_128513_(out[494], out[382], _071630_);
  xor g_128514_(out[484], out[372], _071632_);
  or g_128515_(_071630_, _071632_, _071633_);
  xor g_128516_(out[493], out[381], _071634_);
  xor g_128517_(out[483], out[371], _071635_);
  and g_128518_(_098030_, out[379], _071636_);
  xor g_128519_(out[486], out[374], _071637_);
  xor g_128520_(out[490], out[378], _071638_);
  xor g_128521_(out[485], out[373], _071639_);
  xor g_128522_(out[495], out[383], _071640_);
  xor g_128523_(out[488], out[376], _071641_);
  or g_128524_(_071634_, _071641_, _071643_);
  xor g_128525_(out[482], out[370], _071644_);
  or g_128526_(_071638_, _071644_, _071645_);
  or g_128527_(_071643_, _071645_, _071646_);
  or g_128528_(_071628_, _071635_, _071647_);
  or g_128529_(_071639_, _071647_, _071648_);
  or g_128530_(_071646_, _071648_, _071649_);
  or g_128531_(_071633_, _071649_, _071650_);
  xor g_128532_(out[492], out[380], _071651_);
  or g_128533_(_071636_, _071651_, _071652_);
  xor g_128534_(out[487], out[375], _071654_);
  or g_128535_(_071637_, _071654_, _071655_);
  or g_128536_(_071652_, _071655_, _071656_);
  or g_128537_(_071626_, _071627_, _071657_);
  or g_128538_(_071640_, _071657_, _071658_);
  or g_128539_(_071656_, _071658_, _071659_);
  or g_128540_(_071629_, _071659_, _071660_);
  or g_128541_(_071650_, _071660_, _071661_);
  not g_128542_(_071661_, _071662_);
  xor g_128543_(out[481], out[353], _071663_);
  and g_128544_(_098030_, out[363], _071665_);
  and g_128545_(out[491], _049411_, _071666_);
  xor g_128546_(out[494], out[366], _071667_);
  xor g_128547_(out[483], out[355], _071668_);
  xor g_128548_(out[484], out[356], _071669_);
  xor g_128549_(out[482], out[354], _071670_);
  xor g_128550_(out[489], out[361], _071671_);
  xor g_128551_(out[480], out[352], _071672_);
  xor g_128552_(out[492], out[364], _071673_);
  xor g_128553_(out[486], out[358], _071674_);
  xor g_128554_(out[490], out[362], _071676_);
  xor g_128555_(out[485], out[357], _071677_);
  xor g_128556_(out[495], out[367], _071678_);
  xor g_128557_(out[493], out[365], _071679_);
  xor g_128558_(out[488], out[360], _071680_);
  or g_128559_(_071667_, _071669_, _071681_);
  or g_128560_(_071679_, _071680_, _071682_);
  or g_128561_(_071670_, _071676_, _071683_);
  or g_128562_(_071682_, _071683_, _071684_);
  or g_128563_(_071668_, _071671_, _071685_);
  or g_128564_(_071672_, _071677_, _071687_);
  or g_128565_(_071685_, _071687_, _071688_);
  or g_128566_(_071684_, _071688_, _071689_);
  or g_128567_(_071665_, _071673_, _071690_);
  xor g_128568_(out[487], out[359], _071691_);
  or g_128569_(_071674_, _071691_, _071692_);
  or g_128570_(_071690_, _071692_, _071693_);
  or g_128571_(_071663_, _071666_, _071694_);
  or g_128572_(_071678_, _071694_, _071695_);
  or g_128573_(_071693_, _071695_, _071696_);
  or g_128574_(_071689_, _071696_, _071698_);
  or g_128575_(_071681_, _071698_, _071699_);
  xor g_128576_(out[482], out[338], _071700_);
  xor g_128577_(out[480], out[336], _071701_);
  xor g_128578_(out[489], out[345], _071702_);
  xor g_128579_(out[488], out[344], _071703_);
  xor g_128580_(out[485], out[341], _071704_);
  xor g_128581_(out[494], out[350], _071705_);
  xor g_128582_(out[493], out[349], _071706_);
  xor g_128583_(out[495], out[351], _071707_);
  xor g_128584_(out[490], out[346], _071709_);
  xor g_128585_(out[486], out[342], _071710_);
  xor g_128586_(out[483], out[339], _071711_);
  and g_128587_(_098030_, out[347], _071712_);
  and g_128588_(out[491], _049400_, _071713_);
  xor g_128589_(out[484], out[340], _071714_);
  xor g_128590_(out[481], out[337], _071715_);
  or g_128591_(_071705_, _071714_, _071716_);
  or g_128592_(_071703_, _071706_, _071717_);
  or g_128593_(_071700_, _071709_, _071718_);
  or g_128594_(_071717_, _071718_, _071720_);
  or g_128595_(_071702_, _071711_, _071721_);
  or g_128596_(_071701_, _071704_, _071722_);
  or g_128597_(_071721_, _071722_, _071723_);
  or g_128598_(_071720_, _071723_, _071724_);
  xor g_128599_(out[492], out[348], _071725_);
  or g_128600_(_071712_, _071725_, _071726_);
  xor g_128601_(out[487], out[343], _071727_);
  or g_128602_(_071710_, _071727_, _071728_);
  or g_128603_(_071726_, _071728_, _071729_);
  or g_128604_(_071713_, _071715_, _071731_);
  or g_128605_(_071707_, _071731_, _071732_);
  or g_128606_(_071729_, _071732_, _071733_);
  or g_128607_(_071724_, _071733_, _071734_);
  or g_128608_(_071716_, _071734_, _071735_);
  not g_128609_(_071735_, _071736_);
  and g_128610_(_098030_, out[331], _071737_);
  and g_128611_(out[491], _098294_, _071738_);
  xor g_128612_(out[484], out[324], _071739_);
  xor g_128613_(out[494], out[334], _071740_);
  or g_128614_(_071739_, _071740_, _071742_);
  xor g_128615_(out[493], out[333], _071743_);
  xor g_128616_(out[483], out[323], _071744_);
  xor g_128617_(out[480], out[320], _071745_);
  xor g_128618_(out[490], out[330], _071746_);
  xor g_128619_(out[495], out[335], _071747_);
  xor g_128620_(out[486], out[326], _071748_);
  xor g_128621_(out[485], out[325], _071749_);
  xor g_128622_(out[488], out[328], _071750_);
  or g_128623_(_071743_, _071750_, _071751_);
  xor g_128624_(out[482], out[322], _071753_);
  xor g_128625_(out[489], out[329], _071754_);
  xor g_128626_(out[481], out[321], _071755_);
  or g_128627_(_071746_, _071753_, _071756_);
  or g_128628_(_071751_, _071756_, _071757_);
  or g_128629_(_071744_, _071754_, _071758_);
  or g_128630_(_071749_, _071758_, _071759_);
  or g_128631_(_071757_, _071759_, _071760_);
  or g_128632_(_071742_, _071760_, _071761_);
  xor g_128633_(out[492], out[332], _071762_);
  or g_128634_(_071737_, _071762_, _071764_);
  xor g_128635_(out[487], out[327], _071765_);
  or g_128636_(_071748_, _071765_, _071766_);
  or g_128637_(_071764_, _071766_, _071767_);
  or g_128638_(_071738_, _071755_, _071768_);
  or g_128639_(_071747_, _071768_, _071769_);
  or g_128640_(_071767_, _071769_, _071770_);
  or g_128641_(_071745_, _071770_, _071771_);
  or g_128642_(_071761_, _071771_, _071772_);
  xor g_128643_(out[481], out[305], _071773_);
  and g_128644_(out[491], _098283_, _071775_);
  xor g_128645_(out[489], out[313], _071776_);
  xor g_128646_(out[480], out[304], _071777_);
  xor g_128647_(out[494], out[318], _071778_);
  xor g_128648_(out[484], out[308], _071779_);
  or g_128649_(_071778_, _071779_, _071780_);
  xor g_128650_(out[493], out[317], _071781_);
  xor g_128651_(out[483], out[307], _071782_);
  and g_128652_(_098030_, out[315], _071783_);
  xor g_128653_(out[486], out[310], _071784_);
  xor g_128654_(out[490], out[314], _071786_);
  xor g_128655_(out[485], out[309], _071787_);
  xor g_128656_(out[495], out[319], _071788_);
  xor g_128657_(out[488], out[312], _071789_);
  or g_128658_(_071781_, _071789_, _071790_);
  xor g_128659_(out[482], out[306], _071791_);
  or g_128660_(_071786_, _071791_, _071792_);
  or g_128661_(_071790_, _071792_, _071793_);
  or g_128662_(_071776_, _071782_, _071794_);
  or g_128663_(_071787_, _071794_, _071795_);
  or g_128664_(_071793_, _071795_, _071797_);
  or g_128665_(_071780_, _071797_, _071798_);
  xor g_128666_(out[492], out[316], _071799_);
  or g_128667_(_071783_, _071799_, _071800_);
  xor g_128668_(out[487], out[311], _071801_);
  or g_128669_(_071784_, _071801_, _071802_);
  or g_128670_(_071800_, _071802_, _071803_);
  or g_128671_(_071773_, _071775_, _071804_);
  or g_128672_(_071788_, _071804_, _071805_);
  or g_128673_(_071803_, _071805_, _071806_);
  or g_128674_(_071777_, _071806_, _071808_);
  or g_128675_(_071798_, _071808_, _071809_);
  xor g_128676_(out[481], out[289], _071810_);
  and g_128677_(out[491], _098272_, _071811_);
  xor g_128678_(out[489], out[297], _071812_);
  xor g_128679_(out[480], out[288], _071813_);
  xor g_128680_(out[494], out[302], _071814_);
  xor g_128681_(out[484], out[292], _071815_);
  or g_128682_(_071814_, _071815_, _071816_);
  xor g_128683_(out[493], out[301], _071817_);
  xor g_128684_(out[483], out[291], _071819_);
  and g_128685_(_098030_, out[299], _071820_);
  xor g_128686_(out[486], out[294], _071821_);
  xor g_128687_(out[490], out[298], _071822_);
  xor g_128688_(out[485], out[293], _071823_);
  xor g_128689_(out[495], out[303], _071824_);
  xor g_128690_(out[488], out[296], _071825_);
  or g_128691_(_071817_, _071825_, _071826_);
  xor g_128692_(out[482], out[290], _071827_);
  or g_128693_(_071822_, _071827_, _071828_);
  or g_128694_(_071826_, _071828_, _071830_);
  or g_128695_(_071812_, _071819_, _071831_);
  or g_128696_(_071823_, _071831_, _071832_);
  or g_128697_(_071830_, _071832_, _071833_);
  or g_128698_(_071816_, _071833_, _071834_);
  xor g_128699_(out[492], out[300], _071835_);
  or g_128700_(_071820_, _071835_, _071836_);
  xor g_128701_(out[487], out[295], _071837_);
  or g_128702_(_071821_, _071837_, _071838_);
  or g_128703_(_071836_, _071838_, _071839_);
  or g_128704_(_071810_, _071811_, _071841_);
  or g_128705_(_071824_, _071841_, _071842_);
  or g_128706_(_071839_, _071842_, _071843_);
  or g_128707_(_071813_, _071843_, _071844_);
  or g_128708_(_071834_, _071844_, _071845_);
  xor g_128709_(out[481], out[273], _071846_);
  and g_128710_(_098030_, out[283], _071847_);
  and g_128711_(out[491], _098261_, _071848_);
  xor g_128712_(out[494], out[286], _071849_);
  xor g_128713_(out[483], out[275], _071850_);
  xor g_128714_(out[484], out[276], _071852_);
  xor g_128715_(out[482], out[274], _071853_);
  xor g_128716_(out[489], out[281], _071854_);
  xor g_128717_(out[480], out[272], _071855_);
  xor g_128718_(out[492], out[284], _071856_);
  xor g_128719_(out[486], out[278], _071857_);
  xor g_128720_(out[490], out[282], _071858_);
  xor g_128721_(out[485], out[277], _071859_);
  xor g_128722_(out[495], out[287], _071860_);
  xor g_128723_(out[493], out[285], _071861_);
  xor g_128724_(out[488], out[280], _071863_);
  or g_128725_(_071849_, _071852_, _071864_);
  or g_128726_(_071861_, _071863_, _071865_);
  or g_128727_(_071853_, _071858_, _071866_);
  or g_128728_(_071865_, _071866_, _071867_);
  or g_128729_(_071850_, _071854_, _071868_);
  or g_128730_(_071855_, _071859_, _071869_);
  or g_128731_(_071868_, _071869_, _071870_);
  or g_128732_(_071867_, _071870_, _071871_);
  or g_128733_(_071847_, _071856_, _071872_);
  xor g_128734_(out[487], out[279], _071874_);
  or g_128735_(_071857_, _071874_, _071875_);
  or g_128736_(_071872_, _071875_, _071876_);
  or g_128737_(_071846_, _071848_, _071877_);
  or g_128738_(_071860_, _071877_, _071878_);
  or g_128739_(_071876_, _071878_, _071879_);
  or g_128740_(_071871_, _071879_, _071880_);
  or g_128741_(_071864_, _071880_, _071881_);
  and g_128742_(out[491], _098250_, _071882_);
  and g_128743_(_098030_, out[267], _071883_);
  xor g_128744_(out[484], out[260], _071885_);
  xor g_128745_(out[481], out[257], _071886_);
  xor g_128746_(out[485], out[261], _071887_);
  xor g_128747_(out[489], out[265], _071888_);
  xor g_128748_(out[493], out[269], _071889_);
  xor g_128749_(out[490], out[266], _071890_);
  xor g_128750_(out[486], out[262], _071891_);
  xor g_128751_(out[488], out[264], _071892_);
  or g_128752_(_071889_, _071892_, _071893_);
  xor g_128753_(out[482], out[258], _071894_);
  xor g_128754_(out[495], out[271], _071896_);
  xor g_128755_(out[483], out[259], _071897_);
  xor g_128756_(out[494], out[270], _071898_);
  xor g_128757_(out[480], out[256], _071899_);
  or g_128758_(_071890_, _071894_, _071900_);
  or g_128759_(_071893_, _071900_, _071901_);
  or g_128760_(_071888_, _071897_, _071902_);
  or g_128761_(_071887_, _071902_, _071903_);
  or g_128762_(_071901_, _071903_, _071904_);
  or g_128763_(_071885_, _071898_, _071905_);
  or g_128764_(_071904_, _071905_, _071907_);
  xor g_128765_(out[492], out[268], _071908_);
  or g_128766_(_071883_, _071908_, _071909_);
  xor g_128767_(out[487], out[263], _071910_);
  or g_128768_(_071891_, _071910_, _071911_);
  or g_128769_(_071909_, _071911_, _071912_);
  or g_128770_(_071882_, _071886_, _071913_);
  or g_128771_(_071896_, _071913_, _071914_);
  or g_128772_(_071912_, _071914_, _071915_);
  or g_128773_(_071899_, _071915_, _071916_);
  or g_128774_(_071907_, _071916_, _071918_);
  not g_128775_(_071918_, _071919_);
  xor g_128776_(out[488], out[248], _071920_);
  xor g_128777_(out[485], out[245], _071921_);
  xor g_128778_(out[483], out[243], _071922_);
  xor g_128779_(out[494], out[254], _071923_);
  xor g_128780_(out[493], out[253], _071924_);
  xor g_128781_(out[482], out[242], _071925_);
  xor g_128782_(out[489], out[249], _071926_);
  xor g_128783_(out[486], out[246], _071927_);
  xor g_128784_(out[495], out[255], _071929_);
  xor g_128785_(out[490], out[250], _071930_);
  xor g_128786_(out[484], out[244], _071931_);
  xor g_128787_(out[480], out[240], _071932_);
  and g_128788_(_098030_, out[251], _071933_);
  and g_128789_(out[491], _098239_, _071934_);
  or g_128790_(_071920_, _071924_, _071935_);
  xor g_128791_(out[481], out[241], _071936_);
  or g_128792_(_071925_, _071930_, _071937_);
  or g_128793_(_071935_, _071937_, _071938_);
  or g_128794_(_071922_, _071926_, _071940_);
  or g_128795_(_071921_, _071940_, _071941_);
  or g_128796_(_071938_, _071941_, _071942_);
  or g_128797_(_071923_, _071931_, _071943_);
  or g_128798_(_071942_, _071943_, _071944_);
  xor g_128799_(out[492], out[252], _071945_);
  or g_128800_(_071933_, _071945_, _071946_);
  xor g_128801_(out[487], out[247], _071947_);
  or g_128802_(_071927_, _071947_, _071948_);
  or g_128803_(_071946_, _071948_, _071949_);
  or g_128804_(_071934_, _071936_, _071951_);
  or g_128805_(_071929_, _071951_, _071952_);
  or g_128806_(_071949_, _071952_, _071953_);
  or g_128807_(_071932_, _071953_, _071954_);
  or g_128808_(_071944_, _071954_, _071955_);
  not g_128809_(_071955_, _071956_);
  and g_128810_(_098030_, out[235], _071957_);
  xor g_128811_(out[493], out[237], _071958_);
  xor g_128812_(out[480], out[224], _071959_);
  xor g_128813_(out[481], out[225], _071960_);
  and g_128814_(out[491], _098228_, _071962_);
  xor g_128815_(out[484], out[228], _071963_);
  xor g_128816_(out[488], out[232], _071964_);
  xor g_128817_(out[494], out[238], _071965_);
  xor g_128818_(out[485], out[229], _071966_);
  xor g_128819_(out[482], out[226], _071967_);
  xor g_128820_(out[489], out[233], _071968_);
  xor g_128821_(out[487], out[231], _071969_);
  xor g_128822_(out[483], out[227], _071970_);
  xor g_128823_(out[490], out[234], _071971_);
  xor g_128824_(out[495], out[239], _071973_);
  xor g_128825_(out[486], out[230], _071974_);
  or g_128826_(_071963_, _071965_, _071975_);
  or g_128827_(_071958_, _071964_, _071976_);
  or g_128828_(_071967_, _071971_, _071977_);
  or g_128829_(_071976_, _071977_, _071978_);
  or g_128830_(_071968_, _071970_, _071979_);
  or g_128831_(_071959_, _071966_, _071980_);
  or g_128832_(_071979_, _071980_, _071981_);
  or g_128833_(_071978_, _071981_, _071982_);
  xor g_128834_(out[492], out[236], _071984_);
  or g_128835_(_071957_, _071984_, _071985_);
  or g_128836_(_071969_, _071974_, _071986_);
  or g_128837_(_071985_, _071986_, _071987_);
  or g_128838_(_071960_, _071962_, _071988_);
  or g_128839_(_071973_, _071988_, _071989_);
  or g_128840_(_071987_, _071989_, _071990_);
  or g_128841_(_071982_, _071990_, _071991_);
  or g_128842_(_071975_, _071991_, _071992_);
  not g_128843_(_071992_, _071993_);
  xor g_128844_(out[481], out[209], _071995_);
  and g_128845_(out[491], _098217_, _071996_);
  xor g_128846_(out[489], out[217], _071997_);
  xor g_128847_(out[480], out[208], _071998_);
  xor g_128848_(out[494], out[222], _071999_);
  xor g_128849_(out[484], out[212], _072000_);
  or g_128850_(_071999_, _072000_, _072001_);
  xor g_128851_(out[493], out[221], _072002_);
  xor g_128852_(out[483], out[211], _072003_);
  and g_128853_(_098030_, out[219], _072004_);
  xor g_128854_(out[486], out[214], _072006_);
  xor g_128855_(out[490], out[218], _072007_);
  xor g_128856_(out[485], out[213], _072008_);
  xor g_128857_(out[495], out[223], _072009_);
  xor g_128858_(out[488], out[216], _072010_);
  or g_128859_(_072002_, _072010_, _072011_);
  xor g_128860_(out[482], out[210], _072012_);
  or g_128861_(_072007_, _072012_, _072013_);
  or g_128862_(_072011_, _072013_, _072014_);
  or g_128863_(_071997_, _072003_, _072015_);
  or g_128864_(_072008_, _072015_, _072017_);
  or g_128865_(_072014_, _072017_, _072018_);
  or g_128866_(_072001_, _072018_, _072019_);
  xor g_128867_(out[492], out[220], _072020_);
  or g_128868_(_072004_, _072020_, _072021_);
  xor g_128869_(out[487], out[215], _072022_);
  or g_128870_(_072006_, _072022_, _072023_);
  or g_128871_(_072021_, _072023_, _072024_);
  or g_128872_(_071995_, _071996_, _072025_);
  or g_128873_(_072009_, _072025_, _072026_);
  or g_128874_(_072024_, _072026_, _072028_);
  or g_128875_(_071998_, _072028_, _072029_);
  or g_128876_(_072019_, _072029_, _072030_);
  xor g_128877_(out[481], out[193], _072031_);
  and g_128878_(out[491], _098206_, _072032_);
  xor g_128879_(out[489], out[201], _072033_);
  xor g_128880_(out[480], out[192], _072034_);
  xor g_128881_(out[494], out[206], _072035_);
  xor g_128882_(out[484], out[196], _072036_);
  or g_128883_(_072035_, _072036_, _072037_);
  xor g_128884_(out[493], out[205], _072039_);
  xor g_128885_(out[483], out[195], _072040_);
  and g_128886_(_098030_, out[203], _072041_);
  xor g_128887_(out[486], out[198], _072042_);
  xor g_128888_(out[490], out[202], _072043_);
  xor g_128889_(out[485], out[197], _072044_);
  xor g_128890_(out[495], out[207], _072045_);
  xor g_128891_(out[488], out[200], _072046_);
  or g_128892_(_072039_, _072046_, _072047_);
  xor g_128893_(out[482], out[194], _072048_);
  or g_128894_(_072043_, _072048_, _072050_);
  or g_128895_(_072047_, _072050_, _072051_);
  or g_128896_(_072033_, _072040_, _072052_);
  or g_128897_(_072044_, _072052_, _072053_);
  or g_128898_(_072051_, _072053_, _072054_);
  or g_128899_(_072037_, _072054_, _072055_);
  xor g_128900_(out[492], out[204], _072056_);
  or g_128901_(_072041_, _072056_, _072057_);
  xor g_128902_(out[487], out[199], _072058_);
  or g_128903_(_072042_, _072058_, _072059_);
  or g_128904_(_072057_, _072059_, _072061_);
  or g_128905_(_072031_, _072032_, _072062_);
  or g_128906_(_072045_, _072062_, _072063_);
  or g_128907_(_072061_, _072063_, _072064_);
  or g_128908_(_072034_, _072064_, _072065_);
  or g_128909_(_072055_, _072065_, _072066_);
  and g_128910_(out[491], _098195_, _072067_);
  and g_128911_(_098030_, out[187], _072068_);
  xor g_128912_(out[481], out[177], _072069_);
  xor g_128913_(out[483], out[179], _072070_);
  xor g_128914_(out[487], out[183], _072072_);
  xor g_128915_(out[489], out[185], _072073_);
  xor g_128916_(out[495], out[191], _072074_);
  xor g_128917_(out[482], out[178], _072075_);
  xor g_128918_(out[494], out[190], _072076_);
  xor g_128919_(out[493], out[189], _072077_);
  xor g_128920_(out[488], out[184], _072078_);
  or g_128921_(_072077_, _072078_, _072079_);
  xor g_128922_(out[484], out[180], _072080_);
  xor g_128923_(out[486], out[182], _072081_);
  xor g_128924_(out[490], out[186], _072083_);
  xor g_128925_(out[485], out[181], _072084_);
  xor g_128926_(out[480], out[176], _072085_);
  or g_128927_(_072075_, _072083_, _072086_);
  or g_128928_(_072079_, _072086_, _072087_);
  or g_128929_(_072070_, _072073_, _072088_);
  or g_128930_(_072084_, _072088_, _072089_);
  or g_128931_(_072087_, _072089_, _072090_);
  or g_128932_(_072076_, _072080_, _072091_);
  or g_128933_(_072090_, _072091_, _072092_);
  xor g_128934_(out[492], out[188], _072094_);
  or g_128935_(_072068_, _072094_, _072095_);
  or g_128936_(_072072_, _072081_, _072096_);
  or g_128937_(_072095_, _072096_, _072097_);
  or g_128938_(_072067_, _072069_, _072098_);
  or g_128939_(_072074_, _072098_, _072099_);
  or g_128940_(_072097_, _072099_, _072100_);
  or g_128941_(_072085_, _072100_, _072101_);
  or g_128942_(_072092_, _072101_, _072102_);
  not g_128943_(_072102_, _072103_);
  xor g_128944_(out[490], out[170], _072105_);
  xor g_128945_(out[482], out[162], _072106_);
  xor g_128946_(out[481], out[161], _072107_);
  and g_128947_(_098030_, out[171], _072108_);
  and g_128948_(out[491], _098184_, _072109_);
  xor g_128949_(out[493], out[173], _072110_);
  xor g_128950_(out[483], out[163], _072111_);
  xor g_128951_(out[494], out[174], _072112_);
  xor g_128952_(out[492], out[172], _072113_);
  xor g_128953_(out[488], out[168], _072114_);
  xor g_128954_(out[495], out[175], _072116_);
  xor g_128955_(out[485], out[165], _072117_);
  xor g_128956_(out[486], out[166], _072118_);
  xor g_128957_(out[480], out[160], _072119_);
  xor g_128958_(out[484], out[164], _072120_);
  or g_128959_(_072110_, _072114_, _072121_);
  xor g_128960_(out[489], out[169], _072122_);
  or g_128961_(_072105_, _072106_, _072123_);
  or g_128962_(_072121_, _072123_, _072124_);
  or g_128963_(_072111_, _072122_, _072125_);
  or g_128964_(_072117_, _072125_, _072127_);
  or g_128965_(_072124_, _072127_, _072128_);
  or g_128966_(_072112_, _072120_, _072129_);
  or g_128967_(_072128_, _072129_, _072130_);
  or g_128968_(_072108_, _072113_, _072131_);
  xor g_128969_(out[487], out[167], _072132_);
  or g_128970_(_072118_, _072132_, _072133_);
  or g_128971_(_072131_, _072133_, _072134_);
  or g_128972_(_072107_, _072109_, _072135_);
  or g_128973_(_072116_, _072135_, _072136_);
  or g_128974_(_072134_, _072136_, _072138_);
  or g_128975_(_072119_, _072138_, _072139_);
  or g_128976_(_072130_, _072139_, _072140_);
  not g_128977_(_072140_, _072141_);
  xor g_128978_(out[490], out[154], _072142_);
  xor g_128979_(out[482], out[146], _072143_);
  xor g_128980_(out[481], out[145], _072144_);
  and g_128981_(_098030_, out[155], _072145_);
  and g_128982_(out[491], _098173_, _072146_);
  xor g_128983_(out[493], out[157], _072147_);
  xor g_128984_(out[483], out[147], _072149_);
  xor g_128985_(out[494], out[158], _072150_);
  xor g_128986_(out[492], out[156], _072151_);
  xor g_128987_(out[488], out[152], _072152_);
  xor g_128988_(out[495], out[159], _072153_);
  xor g_128989_(out[485], out[149], _072154_);
  xor g_128990_(out[486], out[150], _072155_);
  xor g_128991_(out[480], out[144], _072156_);
  xor g_128992_(out[484], out[148], _072157_);
  or g_128993_(_072147_, _072152_, _072158_);
  xor g_128994_(out[489], out[153], _072160_);
  or g_128995_(_072142_, _072143_, _072161_);
  or g_128996_(_072158_, _072161_, _072162_);
  or g_128997_(_072149_, _072160_, _072163_);
  or g_128998_(_072154_, _072163_, _072164_);
  or g_128999_(_072162_, _072164_, _072165_);
  or g_129000_(_072150_, _072157_, _072166_);
  or g_129001_(_072165_, _072166_, _072167_);
  or g_129002_(_072145_, _072151_, _072168_);
  xor g_129003_(out[487], out[151], _072169_);
  or g_129004_(_072155_, _072169_, _072171_);
  or g_129005_(_072168_, _072171_, _072172_);
  or g_129006_(_072144_, _072146_, _072173_);
  or g_129007_(_072153_, _072173_, _072174_);
  or g_129008_(_072172_, _072174_, _072175_);
  or g_129009_(_072156_, _072175_, _072176_);
  or g_129010_(_072167_, _072176_, _072177_);
  not g_129011_(_072177_, _072178_);
  xor g_129012_(out[481], out[129], _072179_);
  and g_129013_(out[491], _098162_, _072180_);
  xor g_129014_(out[494], out[142], _072182_);
  xor g_129015_(out[483], out[131], _072183_);
  xor g_129016_(out[484], out[132], _072184_);
  xor g_129017_(out[482], out[130], _072185_);
  xor g_129018_(out[489], out[137], _072186_);
  xor g_129019_(out[480], out[128], _072187_);
  and g_129020_(_098030_, out[139], _072188_);
  xor g_129021_(out[486], out[134], _072189_);
  xor g_129022_(out[490], out[138], _072190_);
  xor g_129023_(out[485], out[133], _072191_);
  xor g_129024_(out[495], out[143], _072193_);
  xor g_129025_(out[493], out[141], _072194_);
  xor g_129026_(out[488], out[136], _072195_);
  or g_129027_(_072182_, _072184_, _072196_);
  or g_129028_(_072194_, _072195_, _072197_);
  or g_129029_(_072185_, _072190_, _072198_);
  or g_129030_(_072197_, _072198_, _072199_);
  or g_129031_(_072183_, _072186_, _072200_);
  or g_129032_(_072187_, _072191_, _072201_);
  or g_129033_(_072200_, _072201_, _072202_);
  or g_129034_(_072199_, _072202_, _072204_);
  xor g_129035_(out[492], out[140], _072205_);
  or g_129036_(_072188_, _072205_, _072206_);
  xor g_129037_(out[487], out[135], _072207_);
  or g_129038_(_072189_, _072207_, _072208_);
  or g_129039_(_072206_, _072208_, _072209_);
  or g_129040_(_072179_, _072180_, _072210_);
  or g_129041_(_072193_, _072210_, _072211_);
  or g_129042_(_072209_, _072211_, _072212_);
  or g_129043_(_072204_, _072212_, _072213_);
  or g_129044_(_072196_, _072213_, _072215_);
  xor g_129045_(out[493], out[125], _072216_);
  xor g_129046_(out[482], out[114], _072217_);
  xor g_129047_(out[485], out[117], _072218_);
  xor g_129048_(out[489], out[121], _072219_);
  xor g_129049_(out[484], out[116], _072220_);
  xor g_129050_(out[488], out[120], _072221_);
  xor g_129051_(out[494], out[126], _072222_);
  xor g_129052_(out[486], out[118], _072223_);
  xor g_129053_(out[495], out[127], _072224_);
  xor g_129054_(out[490], out[122], _072226_);
  xor g_129055_(out[480], out[112], _072227_);
  xor g_129056_(out[483], out[115], _072228_);
  and g_129057_(_098030_, out[123], _072229_);
  and g_129058_(out[491], _098151_, _072230_);
  xor g_129059_(out[481], out[113], _072231_);
  or g_129060_(_072220_, _072222_, _072232_);
  or g_129061_(_072216_, _072221_, _072233_);
  or g_129062_(_072217_, _072226_, _072234_);
  or g_129063_(_072233_, _072234_, _072235_);
  or g_129064_(_072219_, _072228_, _072237_);
  or g_129065_(_072218_, _072227_, _072238_);
  or g_129066_(_072237_, _072238_, _072239_);
  or g_129067_(_072235_, _072239_, _072240_);
  xor g_129068_(out[492], out[124], _072241_);
  or g_129069_(_072229_, _072241_, _072242_);
  xor g_129070_(out[487], out[119], _072243_);
  or g_129071_(_072223_, _072243_, _072244_);
  or g_129072_(_072242_, _072244_, _072245_);
  or g_129073_(_072230_, _072231_, _072246_);
  or g_129074_(_072224_, _072246_, _072248_);
  or g_129075_(_072245_, _072248_, _072249_);
  or g_129076_(_072240_, _072249_, _072250_);
  or g_129077_(_072232_, _072250_, _072251_);
  xor g_129078_(out[481], out[97], _072252_);
  and g_129079_(out[491], _098140_, _072253_);
  xor g_129080_(out[489], out[105], _072254_);
  xor g_129081_(out[480], out[96], _072255_);
  xor g_129082_(out[494], out[110], _072256_);
  xor g_129083_(out[484], out[100], _072257_);
  or g_129084_(_072256_, _072257_, _072259_);
  xor g_129085_(out[493], out[109], _072260_);
  xor g_129086_(out[483], out[99], _072261_);
  and g_129087_(_098030_, out[107], _072262_);
  xor g_129088_(out[486], out[102], _072263_);
  xor g_129089_(out[490], out[106], _072264_);
  xor g_129090_(out[485], out[101], _072265_);
  xor g_129091_(out[495], out[111], _072266_);
  xor g_129092_(out[488], out[104], _072267_);
  or g_129093_(_072260_, _072267_, _072268_);
  xor g_129094_(out[482], out[98], _072270_);
  or g_129095_(_072264_, _072270_, _072271_);
  or g_129096_(_072268_, _072271_, _072272_);
  or g_129097_(_072254_, _072261_, _072273_);
  or g_129098_(_072265_, _072273_, _072274_);
  or g_129099_(_072272_, _072274_, _072275_);
  or g_129100_(_072259_, _072275_, _072276_);
  xor g_129101_(out[492], out[108], _072277_);
  or g_129102_(_072262_, _072277_, _072278_);
  xor g_129103_(out[487], out[103], _072279_);
  or g_129104_(_072263_, _072279_, _072281_);
  or g_129105_(_072278_, _072281_, _072282_);
  or g_129106_(_072252_, _072253_, _072283_);
  or g_129107_(_072266_, _072283_, _072284_);
  or g_129108_(_072282_, _072284_, _072285_);
  or g_129109_(_072255_, _072285_, _072286_);
  or g_129110_(_072276_, _072286_, _072287_);
  xor g_129111_(out[481], out[81], _072288_);
  and g_129112_(_098030_, out[91], _072289_);
  and g_129113_(out[491], _098129_, _072290_);
  xor g_129114_(out[489], out[89], _072292_);
  xor g_129115_(out[480], out[80], _072293_);
  xor g_129116_(out[494], out[94], _072294_);
  xor g_129117_(out[484], out[84], _072295_);
  or g_129118_(_072294_, _072295_, _072296_);
  xor g_129119_(out[493], out[93], _072297_);
  xor g_129120_(out[483], out[83], _072298_);
  xor g_129121_(out[492], out[92], _072299_);
  xor g_129122_(out[486], out[86], _072300_);
  xor g_129123_(out[490], out[90], _072301_);
  xor g_129124_(out[485], out[85], _072303_);
  xor g_129125_(out[495], out[95], _072304_);
  xor g_129126_(out[488], out[88], _072305_);
  or g_129127_(_072297_, _072305_, _072306_);
  xor g_129128_(out[482], out[82], _072307_);
  or g_129129_(_072301_, _072307_, _072308_);
  or g_129130_(_072306_, _072308_, _072309_);
  or g_129131_(_072292_, _072298_, _072310_);
  or g_129132_(_072303_, _072310_, _072311_);
  or g_129133_(_072309_, _072311_, _072312_);
  or g_129134_(_072296_, _072312_, _072314_);
  or g_129135_(_072289_, _072299_, _072315_);
  xor g_129136_(out[487], out[87], _072316_);
  or g_129137_(_072300_, _072316_, _072317_);
  or g_129138_(_072315_, _072317_, _072318_);
  or g_129139_(_072288_, _072290_, _072319_);
  or g_129140_(_072304_, _072319_, _072320_);
  or g_129141_(_072318_, _072320_, _072321_);
  or g_129142_(_072293_, _072321_, _072322_);
  or g_129143_(_072314_, _072322_, _072323_);
  xor g_129144_(out[492], out[76], _072325_);
  and g_129145_(_098030_, out[75], _072326_);
  xor g_129146_(out[488], out[72], _072327_);
  xor g_129147_(out[486], out[70], _072328_);
  xor g_129148_(out[493], out[77], _072329_);
  xor g_129149_(out[494], out[78], _072330_);
  xor g_129150_(out[482], out[66], _072331_);
  xor g_129151_(out[489], out[73], _072332_);
  xor g_129152_(out[485], out[69], _072333_);
  xor g_129153_(out[481], out[65], _072334_);
  and g_129154_(out[491], _098118_, _072336_);
  or g_129155_(_072327_, _072329_, _072337_);
  xor g_129156_(out[495], out[79], _072338_);
  xor g_129157_(out[490], out[74], _072339_);
  xor g_129158_(out[484], out[68], _072340_);
  xor g_129159_(out[483], out[67], _072341_);
  xor g_129160_(out[480], out[64], _072342_);
  or g_129161_(_072331_, _072339_, _072343_);
  or g_129162_(_072337_, _072343_, _072344_);
  or g_129163_(_072332_, _072341_, _072345_);
  or g_129164_(_072333_, _072345_, _072347_);
  or g_129165_(_072344_, _072347_, _072348_);
  or g_129166_(_072330_, _072340_, _072349_);
  or g_129167_(_072348_, _072349_, _072350_);
  or g_129168_(_072325_, _072326_, _072351_);
  xor g_129169_(out[487], out[71], _072352_);
  or g_129170_(_072328_, _072352_, _072353_);
  or g_129171_(_072351_, _072353_, _072354_);
  or g_129172_(_072334_, _072336_, _072355_);
  or g_129173_(_072338_, _072355_, _072356_);
  or g_129174_(_072354_, _072356_, _072358_);
  or g_129175_(_072342_, _072358_, _072359_);
  or g_129176_(_072350_, _072359_, _072360_);
  xor g_129177_(out[483], out[51], _072361_);
  xor g_129178_(out[484], out[52], _072362_);
  xor g_129179_(out[494], out[62], _072363_);
  xor g_129180_(out[482], out[50], _072364_);
  xor g_129181_(out[485], out[53], _072365_);
  xor g_129182_(out[489], out[57], _072366_);
  xor g_129183_(out[488], out[56], _072367_);
  xor g_129184_(out[495], out[63], _072369_);
  xor g_129185_(out[490], out[58], _072370_);
  xor g_129186_(out[486], out[54], _072371_);
  xor g_129187_(out[480], out[48], _072372_);
  and g_129188_(_098030_, out[59], _072373_);
  and g_129189_(out[491], _098107_, _072374_);
  xor g_129190_(out[493], out[61], _072375_);
  or g_129191_(_072367_, _072375_, _072376_);
  xor g_129192_(out[481], out[49], _072377_);
  or g_129193_(_072364_, _072370_, _072378_);
  or g_129194_(_072376_, _072378_, _072380_);
  or g_129195_(_072361_, _072366_, _072381_);
  or g_129196_(_072365_, _072381_, _072382_);
  or g_129197_(_072380_, _072382_, _072383_);
  or g_129198_(_072362_, _072363_, _072384_);
  or g_129199_(_072383_, _072384_, _072385_);
  xor g_129200_(out[492], out[60], _072386_);
  or g_129201_(_072373_, _072386_, _072387_);
  xor g_129202_(out[487], out[55], _072388_);
  or g_129203_(_072371_, _072388_, _072389_);
  or g_129204_(_072387_, _072389_, _072391_);
  or g_129205_(_072374_, _072377_, _072392_);
  or g_129206_(_072369_, _072392_, _072393_);
  or g_129207_(_072391_, _072393_, _072394_);
  or g_129208_(_072372_, _072394_, _072395_);
  or g_129209_(_072385_, _072395_, _072396_);
  xor g_129210_(out[482], out[34], _072397_);
  and g_129211_(_097986_, out[39], _072398_);
  xor g_129212_(out[485], out[37], _072399_);
  xor g_129213_(out[491], out[43], _072400_);
  or g_129214_(_072399_, _072400_, _072402_);
  xor g_129215_(out[483], out[35], _072403_);
  xor g_129216_(out[493], out[45], _072404_);
  xor g_129217_(out[484], out[36], _072405_);
  xor g_129218_(out[490], out[42], _072406_);
  xor g_129219_(out[486], out[38], _072407_);
  xor g_129220_(out[489], out[41], _072408_);
  and g_129221_(out[487], _098085_, _072409_);
  or g_129222_(_072403_, _072405_, _072410_);
  xor g_129223_(out[492], out[44], _072411_);
  xor g_129224_(out[481], out[33], _072413_);
  xor g_129225_(out[480], out[32], _072414_);
  xor g_129226_(out[494], out[46], _072415_);
  xor g_129227_(out[488], out[40], _072416_);
  or g_129228_(_072406_, _072407_, _072417_);
  or g_129229_(_072410_, _072417_, _072418_);
  or g_129230_(_072402_, _072404_, _072419_);
  or g_129231_(_072418_, _072419_, _072420_);
  or g_129232_(_072411_, _072414_, _072421_);
  or g_129233_(_072420_, _072421_, _072422_);
  or g_129234_(_072397_, _072398_, _072424_);
  xor g_129235_(out[495], out[47], _072425_);
  or g_129236_(_072415_, _072425_, _072426_);
  or g_129237_(_072424_, _072426_, _072427_);
  or g_129238_(_072408_, _072409_, _072428_);
  or g_129239_(_072413_, _072428_, _072429_);
  or g_129240_(_072427_, _072429_, _072430_);
  or g_129241_(_072416_, _072430_, _072431_);
  or g_129242_(_072422_, _072431_, _072432_);
  not g_129243_(_072432_, _072433_);
  xor g_129244_(out[486], out[22], _072435_);
  xor g_129245_(out[490], out[26], _072436_);
  xor g_129246_(out[485], out[21], _072437_);
  and g_129247_(out[492], _098074_, _072438_);
  xor g_129248_(out[481], out[17], _072439_);
  xor g_129249_(out[483], out[19], _072440_);
  xor g_129250_(out[495], out[31], _072441_);
  xor g_129251_(out[487], out[23], _072442_);
  xor g_129252_(out[480], out[16], _072443_);
  xor g_129253_(out[494], out[30], _072444_);
  xor g_129254_(out[484], out[20], _072446_);
  xor g_129255_(out[489], out[25], _072447_);
  xor g_129256_(out[491], out[27], _072448_);
  xor g_129257_(out[482], out[18], _072449_);
  and g_129258_(_098052_, out[28], _072450_);
  or g_129259_(_072444_, _072447_, _072451_);
  or g_129260_(_072435_, _072448_, _072452_);
  or g_129261_(_072451_, _072452_, _072453_);
  or g_129262_(_072436_, _072442_, _072454_);
  or g_129263_(_072446_, _072454_, _072455_);
  or g_129264_(_072453_, _072455_, _072457_);
  or g_129265_(_072443_, _072449_, _072458_);
  or g_129266_(_072457_, _072458_, _072459_);
  xor g_129267_(out[493], out[29], _072460_);
  or g_129268_(_072450_, _072460_, _072461_);
  xor g_129269_(out[488], out[24], _072462_);
  or g_129270_(_072439_, _072462_, _072463_);
  or g_129271_(_072461_, _072463_, _072464_);
  or g_129272_(_072437_, _072438_, _072465_);
  or g_129273_(_072441_, _072465_, _072466_);
  or g_129274_(_072464_, _072466_, _072468_);
  or g_129275_(_072440_, _072468_, _072469_);
  or g_129276_(_072459_, _072469_, _072470_);
  xor g_129277_(out[490], out[10], _072471_);
  xor g_129278_(out[485], out[5], _072472_);
  xor g_129279_(out[491], out[11], _072473_);
  xor g_129280_(out[480], out[0], _072474_);
  or g_129281_(out[487], _097997_, _072475_);
  or g_129282_(_097986_, out[7], _072476_);
  xor g_129283_(out[483], out[3], _072477_);
  xor g_129284_(out[493], out[13], _072479_);
  xor g_129285_(out[484], out[4], _072480_);
  xor g_129286_(out[486], out[6], _072481_);
  xor g_129287_(_097964_, out[1], _072482_);
  xor g_129288_(out[494], out[14], _072483_);
  xor g_129289_(_098019_, out[9], _072484_);
  xor g_129290_(out[492], out[12], _072485_);
  xor g_129291_(_098008_, out[8], _072486_);
  or g_129292_(_072477_, _072480_, _072487_);
  or g_129293_(_072471_, _072481_, _072488_);
  or g_129294_(_072487_, _072488_, _072490_);
  or g_129295_(_072472_, _072473_, _072491_);
  or g_129296_(_072479_, _072491_, _072492_);
  or g_129297_(_072490_, _072492_, _072493_);
  or g_129298_(_072474_, _072485_, _072494_);
  or g_129299_(_072493_, _072494_, _072495_);
  not g_129300_(_072495_, _072496_);
  xor g_129301_(_097975_, out[2], _072497_);
  and g_129302_(_072475_, _072497_, _072498_);
  xor g_129303_(out[495], out[15], _072499_);
  or g_129304_(_072483_, _072499_, _072501_);
  not g_129305_(_072501_, _072502_);
  and g_129306_(_072498_, _072502_, _072503_);
  and g_129307_(_072476_, _072484_, _072504_);
  and g_129308_(_072482_, _072504_, _072505_);
  and g_129309_(_072503_, _072505_, _072506_);
  and g_129310_(_072486_, _072506_, _072507_);
  and g_129311_(_072496_, _072507_, _072508_);
  not g_129312_(_072508_, _072509_);
  or g_129313_(_072470_, _072509_, _072510_);
  and g_129314_(_072470_, _072509_, _072512_);
  xor g_129315_(_072470_, _072508_, _072513_);
  xor g_129316_(_072433_, _072513_, _072514_);
  not g_129317_(_072514_, _072515_);
  or g_129318_(_072396_, _072514_, _072516_);
  xor g_129319_(_072396_, _072514_, _072517_);
  xor g_129320_(_072396_, _072515_, _072518_);
  or g_129321_(_072360_, _072518_, _072519_);
  xor g_129322_(_072360_, _072517_, _072520_);
  not g_129323_(_072520_, _072521_);
  or g_129324_(_072323_, _072520_, _072523_);
  xor g_129325_(_072323_, _072520_, _072524_);
  xor g_129326_(_072323_, _072521_, _072525_);
  or g_129327_(_072287_, _072525_, _072526_);
  xor g_129328_(_072287_, _072524_, _072527_);
  or g_129329_(_072251_, _072527_, _072528_);
  not g_129330_(_072528_, _072529_);
  and g_129331_(_072251_, _072527_, _072530_);
  xor g_129332_(_072251_, _072527_, _072531_);
  or g_129333_(_072529_, _072530_, _072532_);
  or g_129334_(_072215_, _072532_, _072534_);
  xor g_129335_(_072215_, _072531_, _072535_);
  or g_129336_(_072177_, _072535_, _072536_);
  xor g_129337_(_072178_, _072535_, _072537_);
  or g_129338_(_072140_, _072537_, _072538_);
  xor g_129339_(_072141_, _072537_, _072539_);
  or g_129340_(_072102_, _072539_, _072540_);
  xor g_129341_(_072103_, _072539_, _072541_);
  not g_129342_(_072541_, _072542_);
  or g_129343_(_072066_, _072541_, _072543_);
  xor g_129344_(_072066_, _072541_, _072545_);
  xor g_129345_(_072066_, _072542_, _072546_);
  or g_129346_(_072030_, _072546_, _072547_);
  xor g_129347_(_072030_, _072545_, _072548_);
  or g_129348_(_071992_, _072548_, _072549_);
  xor g_129349_(_071993_, _072548_, _072550_);
  or g_129350_(_071955_, _072550_, _072551_);
  xor g_129351_(_071956_, _072550_, _072552_);
  or g_129352_(_071918_, _072552_, _072553_);
  xor g_129353_(_071919_, _072552_, _072554_);
  or g_129354_(_071881_, _072554_, _072556_);
  not g_129355_(_072556_, _072557_);
  and g_129356_(_071881_, _072554_, _072558_);
  xor g_129357_(_071881_, _072554_, _072559_);
  or g_129358_(_072557_, _072558_, _072560_);
  or g_129359_(_071845_, _072560_, _072561_);
  xor g_129360_(_071845_, _072559_, _072562_);
  not g_129361_(_072562_, _072563_);
  or g_129362_(_071809_, _072562_, _072564_);
  xor g_129363_(_071809_, _072562_, _072565_);
  xor g_129364_(_071809_, _072563_, _072567_);
  or g_129365_(_071772_, _072567_, _072568_);
  xor g_129366_(_071772_, _072565_, _072569_);
  or g_129367_(_071735_, _072569_, _072570_);
  xor g_129368_(_071735_, _072569_, _072571_);
  xor g_129369_(_071736_, _072569_, _072572_);
  or g_129370_(_071699_, _072572_, _072573_);
  xor g_129371_(_071699_, _072571_, _072574_);
  or g_129372_(_071661_, _072574_, _072575_);
  xor g_129373_(_071662_, _072574_, _072576_);
  or g_129374_(_071624_, _072576_, _072578_);
  xor g_129375_(_071625_, _072576_, _072579_);
  or g_129376_(_071586_, _072579_, _072580_);
  xor g_129377_(_071588_, _072579_, _072581_);
  or g_129378_(_071549_, _072581_, _072582_);
  xor g_129379_(_071550_, _072581_, _072583_);
  or g_129380_(_071513_, _072583_, _072584_);
  xor g_129381_(_071512_, _072583_, _072585_);
  or g_129382_(_071472_, _072585_, _072586_);
  xor g_129383_(_071473_, _072585_, _072587_);
  not g_129384_(_072587_, _072589_);
  or g_129385_(_071436_, _072587_, _072590_);
  xor g_129386_(_071436_, _072587_, _072591_);
  xor g_129387_(_071436_, _072589_, _072592_);
  or g_129388_(_071399_, _072592_, _072593_);
  xor g_129389_(_071399_, _072591_, _072594_);
  or g_129390_(_071362_, _072594_, _072595_);
  xor g_129391_(_071363_, _072594_, _072596_);
  not g_129392_(_072596_, _072597_);
  or g_129393_(_071326_, _072596_, _072598_);
  xor g_129394_(_071326_, _072596_, _072600_);
  xor g_129395_(_071326_, _072597_, _072601_);
  or g_129396_(_071289_, _072601_, _072602_);
  xor g_129397_(_071289_, _072600_, _072603_);
  or g_129398_(_071253_, _072603_, _072604_);
  xor g_129399_(_071253_, _072603_, _072605_);
  not g_129400_(_072605_, _072606_);
  or g_129401_(_071217_, _072606_, _072607_);
  xor g_129402_(_071217_, _072605_, _072608_);
  not g_129403_(_072608_, _072609_);
  or g_129404_(_071181_, _072608_, _072611_);
  xor g_129405_(_071181_, _072608_, _072612_);
  xor g_129406_(_071181_, _072609_, _072613_);
  or g_129407_(_071144_, _072613_, _072614_);
  xor g_129408_(_071144_, _072612_, _072615_);
  not g_129409_(_072615_, _072616_);
  or g_129410_(_071108_, _072615_, _072617_);
  xor g_129411_(_071108_, _072615_, _072618_);
  xor g_129412_(_071108_, _072616_, _072619_);
  or g_129413_(_071072_, _072619_, _072620_);
  xor g_129414_(_071072_, _072618_, _072622_);
  not g_129415_(_072622_, _072623_);
  or g_129416_(_071035_, _072622_, _072624_);
  xor g_129417_(_071035_, _072622_, _072625_);
  xor g_129418_(_071035_, _072623_, _072626_);
  or g_129419_(_070999_, _072626_, _072627_);
  xor g_129420_(_070999_, _072625_, _072628_);
  or g_129421_(_070963_, _072628_, _072629_);
  not g_129422_(_072629_, _072630_);
  xor g_129423_(_070963_, _072628_, _072631_);
  not g_129424_(_072631_, _072633_);
  or g_129425_(_070926_, _072633_, _072634_);
  not g_129426_(_072634_, _072635_);
  xor g_129427_(_070926_, _072631_, _072636_);
  or g_129428_(_070890_, _072636_, _072637_);
  xor g_129429_(_070890_, _072636_, _072638_);
  not g_129430_(_072638_, _072639_);
  or g_129431_(_070854_, _072639_, _072640_);
  xor g_129432_(_070854_, _072638_, _072641_);
  not g_129433_(_072641_, _072642_);
  or g_129434_(_070818_, _072641_, _072644_);
  xor g_129435_(_070818_, _072641_, _072645_);
  xor g_129436_(_070818_, _072642_, _072646_);
  or g_129437_(_070781_, _072646_, _072647_);
  xor g_129438_(_070781_, _072645_, _072648_);
  not g_129439_(_072648_, _072649_);
  or g_129440_(_070745_, _072648_, _072650_);
  xor g_129441_(_070745_, _072648_, _072651_);
  xor g_129442_(_070745_, _072649_, _072652_);
  or g_129443_(_070709_, _072652_, _072653_);
  xor g_129444_(_070709_, _072651_, _072655_);
  or g_129445_(_070671_, _072655_, _072656_);
  xor g_129446_(_070672_, _072655_, _072657_);
  or g_129447_(_070635_, _072657_, _072658_);
  not g_129448_(_072658_, _072659_);
  xor g_129449_(_070635_, _072657_, _072660_);
  not g_129450_(_072660_, _072661_);
  or g_129451_(_070599_, _072661_, _072662_);
  not g_129452_(_072662_, _072663_);
  xor g_129453_(_070599_, _072660_, _072664_);
  not g_129454_(_072664_, _072666_);
  or g_129455_(_070562_, _072664_, _072667_);
  xor g_129456_(_070562_, _072664_, _072668_);
  xor g_129457_(_070562_, _072666_, _072669_);
  or g_129458_(_070526_, _072669_, _072670_);
  xor g_129459_(_070526_, _072668_, _072671_);
  or g_129460_(_070489_, _072671_, _072672_);
  not g_129461_(_072672_, _072673_);
  xor g_129462_(_070490_, _072671_, _072674_);
  not g_129463_(_072674_, _072675_);
  or g_129464_(_070452_, _072674_, _072677_);
  xor g_129465_(_070452_, _072674_, _072678_);
  xor g_129466_(_070452_, _072675_, _072679_);
  or g_129467_(_070416_, _072679_, _072680_);
  not g_129468_(_072680_, _072681_);
  xor g_129469_(_070416_, _072678_, _072682_);
  not g_129470_(_072682_, _072683_);
  or g_129471_(_070380_, _072682_, _072684_);
  xor g_129472_(_070380_, _072682_, _072685_);
  xor g_129473_(_070380_, _072683_, _072686_);
  or g_129474_(_070343_, _072686_, _072688_);
  xor g_129475_(_070343_, _072685_, _072689_);
  or g_129476_(_070307_, _072689_, _072690_);
  xor g_129477_(_070306_, _072689_, _072691_);
  not g_129478_(_072691_, _072692_);
  or g_129479_(_070268_, _072691_, _072693_);
  xor g_129480_(_070268_, _072691_, _072694_);
  xor g_129481_(_070268_, _072692_, _072695_);
  or g_129482_(_070231_, _072695_, _072696_);
  xor g_129483_(_070231_, _072694_, _072697_);
  not g_129484_(_072697_, _072699_);
  or g_129485_(_070195_, _072697_, _072700_);
  xor g_129486_(_070195_, _072697_, _072701_);
  xor g_129487_(_070195_, _072699_, _072702_);
  or g_129488_(_070159_, _072702_, _072703_);
  xor g_129489_(_070159_, _072701_, _072704_);
  or g_129490_(_070121_, _072704_, _072705_);
  xor g_129491_(_070122_, _072704_, _072706_);
  not g_129492_(_072706_, _072707_);
  or g_129493_(_070085_, _072706_, _072708_);
  xor g_129494_(_070085_, _072706_, _072710_);
  xor g_129495_(_070085_, _072707_, _072711_);
  or g_129496_(_070049_, _072711_, _072712_);
  xor g_129497_(_070049_, _072710_, _072713_);
  or g_129498_(_070011_, _072713_, _072714_);
  xor g_129499_(_070012_, _072713_, _072715_);
  or g_129500_(_069974_, _072715_, _072716_);
  xor g_129501_(_069975_, _072715_, _072717_);
  not g_129502_(_072717_, _072718_);
  or g_129503_(_069938_, _072717_, _072719_);
  xor g_129504_(_069938_, _072717_, _072721_);
  xor g_129505_(_069938_, _072718_, _072722_);
  or g_129506_(_069901_, _072722_, _072723_);
  xor g_129507_(_069901_, _072721_, _072724_);
  or g_129508_(_069864_, _072724_, _072725_);
  xor g_129509_(_069865_, _072724_, _072726_);
  or g_129510_(_069828_, _072726_, _072727_);
  not g_129511_(_072727_, _072728_);
  xor g_129512_(_069828_, _072726_, _072729_);
  not g_129513_(_072729_, _072730_);
  or g_129514_(_069791_, _072730_, _072732_);
  not g_129515_(_072732_, _072733_);
  xor g_129516_(_069791_, _072729_, _072734_);
  or g_129517_(_069754_, _072734_, _072735_);
  xor g_129518_(_069755_, _072734_, _072736_);
  or g_129519_(_069716_, _072736_, _072737_);
  xor g_129520_(_069718_, _072736_, _072738_);
  not g_129521_(_072738_, _072739_);
  or g_129522_(_069680_, _072738_, _072740_);
  xor g_129523_(_069680_, _072738_, _072741_);
  xor g_129524_(_069680_, _072739_, _072743_);
  and g_129525_(_069644_, _072741_, _072744_);
  or g_129526_(_069643_, _072743_, _072745_);
  xor g_129527_(_069643_, _072741_, _072746_);
  or g_129528_(_069605_, _072746_, _072747_);
  xor g_129529_(_069606_, _072746_, _072748_);
  or g_129530_(_069568_, _072748_, _072749_);
  xor g_129531_(_069569_, _072748_, _072750_);
  or g_129532_(_069531_, _072750_, _072751_);
  xor g_129533_(_069532_, _072750_, _072752_);
  or g_129534_(_069493_, _072752_, _072754_);
  xor g_129535_(_069494_, _072752_, _072755_);
  or g_129536_(_069457_, _072755_, _072756_);
  xor g_129537_(_069457_, _072755_, _072757_);
  not g_129538_(_072757_, _072758_);
  or g_129539_(_069421_, _072758_, _072759_);
  not g_129540_(_072759_, _072760_);
  xor g_129541_(_069421_, _072757_, _072761_);
  or g_129542_(_069384_, _072761_, _072762_);
  xor g_129543_(_069384_, _072761_, _072763_);
  not g_129544_(_072763_, _072765_);
  and g_129545_(_069348_, _072763_, _072766_);
  or g_129546_(_069347_, _072765_, _072767_);
  xor g_129547_(_069347_, _072763_, _072768_);
  or g_129548_(_069309_, _072768_, _072769_);
  not g_129549_(_072769_, _072770_);
  xor g_129550_(_069311_, _072768_, _072771_);
  or g_129551_(_069272_, _072771_, _072772_);
  not g_129552_(_072772_, _072773_);
  xor g_129553_(_069273_, _072771_, _072774_);
  or g_129554_(_069236_, _072774_, _072776_);
  not g_129555_(_072776_, _072777_);
  xor g_129556_(_069236_, _072774_, _072778_);
  not g_129557_(_072778_, _072779_);
  or g_129558_(_069199_, _072779_, _072780_);
  xor g_129559_(_069199_, _072778_, _072781_);
  or g_129560_(_069162_, _072781_, _072782_);
  not g_129561_(_072782_, _072783_);
  xor g_129562_(_069163_, _072781_, _072784_);
  or g_129563_(_069126_, _072784_, _072785_);
  not g_129564_(_072785_, _072787_);
  and g_129565_(_069126_, _072784_, _072788_);
  xor g_129566_(_069126_, _072784_, _072789_);
  or g_129567_(_072787_, _072788_, _072790_);
  or g_129568_(_069089_, _072790_, _072791_);
  xor g_129569_(_069089_, _072789_, _072792_);
  or g_129570_(_069052_, _072792_, _072793_);
  xor g_129571_(_069053_, _072792_, _072794_);
  or g_129572_(_069015_, _072794_, _072795_);
  xor g_129573_(_069016_, _072794_, _072796_);
  or g_129574_(_068977_, _072796_, _072798_);
  xor g_129575_(_068978_, _072796_, _072799_);
  or g_129576_(_068940_, _072799_, _072800_);
  xor g_129577_(_068941_, _072799_, _072801_);
  or g_129578_(_068904_, _072801_, _072802_);
  xor g_129579_(_068904_, _072801_, _072803_);
  not g_129580_(_072803_, _072804_);
  or g_129581_(_068867_, _072804_, _072805_);
  not g_129582_(_072805_, _072806_);
  xor g_129583_(_068867_, _072803_, _072807_);
  or g_129584_(_068830_, _072807_, _072809_);
  not g_129585_(_072809_, _072810_);
  xor g_129586_(_068831_, _072807_, _072811_);
  or g_129587_(_068794_, _072811_, _072812_);
  not g_129588_(_072812_, _072813_);
  xor g_129589_(_068794_, _072811_, _072814_);
  not g_129590_(_072814_, _072815_);
  or g_129591_(_068757_, _072815_, _072816_);
  not g_129592_(_072816_, _072817_);
  xor g_129593_(_068757_, _072814_, _072818_);
  not g_129594_(_072818_, _072820_);
  or g_129595_(_068721_, _072818_, _072821_);
  xor g_129596_(_068721_, _072818_, _072822_);
  xor g_129597_(_068721_, _072820_, _072823_);
  or g_129598_(_068685_, _072823_, _072824_);
  xor g_129599_(_068685_, _072822_, _072825_);
  or g_129600_(_068647_, _072825_, _072826_);
  xor g_129601_(_068648_, _072825_, _072827_);
  or g_129602_(_068610_, _072827_, _072828_);
  xor g_129603_(_068611_, _072827_, _072829_);
  not g_129604_(_072829_, _072831_);
  or g_129605_(_068574_, _072829_, _072832_);
  xor g_129606_(_068574_, _072829_, _072833_);
  xor g_129607_(_068574_, _072831_, _072834_);
  or g_129608_(_068537_, _072834_, _072835_);
  xor g_129609_(_068537_, _072833_, _072836_);
  not g_129610_(_072836_, _072837_);
  or g_129611_(_068501_, _072836_, _072838_);
  xor g_129612_(_068501_, _072836_, _072839_);
  xor g_129613_(_068501_, _072837_, _072840_);
  or g_129614_(_068465_, _072840_, _072842_);
  xor g_129615_(_068465_, _072839_, _072843_);
  not g_129616_(_072843_, _072844_);
  or g_129617_(_068428_, _072843_, _072845_);
  xor g_129618_(_068428_, _072843_, _072846_);
  xor g_129619_(_068428_, _072844_, _072847_);
  or g_129620_(_068392_, _072847_, _072848_);
  xor g_129621_(_068392_, _072846_, _072849_);
  or g_129622_(_068355_, _072849_, _072850_);
  xor g_129623_(_068356_, _072849_, _072851_);
  not g_129624_(_072851_, _072853_);
  or g_129625_(_068318_, _072851_, _072854_);
  xor g_129626_(_068318_, _072851_, _072855_);
  xor g_129627_(_068318_, _072853_, _072856_);
  or g_129628_(_068282_, _072856_, _072857_);
  xor g_129629_(_068282_, _072855_, _072858_);
  or g_129630_(_068246_, _072858_, _072859_);
  not g_129631_(_072859_, _072860_);
  and g_129632_(_068246_, _072858_, _072861_);
  xor g_129633_(_068246_, _072858_, _072862_);
  or g_129634_(_072860_, _072861_, _072864_);
  or g_129635_(_068209_, _072864_, _072865_);
  xor g_129636_(_068209_, _072862_, _072866_);
  or g_129637_(_068172_, _072866_, _072867_);
  xor g_129638_(_068173_, _072866_, _072868_);
  or g_129639_(_068135_, _072868_, _072869_);
  xor g_129640_(_068136_, _072868_, _072870_);
  or g_129641_(_068098_, _072870_, _072871_);
  not g_129642_(_072871_, _072872_);
  xor g_129643_(_068098_, _072870_, _072873_);
  not g_129644_(_072873_, _072875_);
  or g_129645_(_068062_, _072875_, _072876_);
  and g_129646_(_068062_, _072875_, _072877_);
  xor g_129647_(_068062_, _072873_, _072878_);
  not g_129648_(_072878_, _072879_);
  and g_129649_(_068026_, _072879_, _072880_);
  not g_129650_(_072880_, _072881_);
  xor g_129651_(_068025_, _072878_, _072882_);
  not g_129652_(_072882_, _072883_);
  or g_129653_(_067988_, _072883_, _072884_);
  xor g_129654_(_067988_, _072882_, _072886_);
  or g_129655_(_067951_, _072886_, _072887_);
  not g_129656_(_072887_, _072888_);
  xor g_129657_(_067952_, _072886_, _072889_);
  or g_129658_(_067914_, _072889_, _072890_);
  xor g_129659_(_067915_, _072889_, _072891_);
  or g_129660_(_067876_, _072891_, _072892_);
  xor g_129661_(_067877_, _072891_, _072893_);
  not g_129662_(_072893_, _072894_);
  or g_129663_(_067840_, _072893_, _072895_);
  xor g_129664_(_067840_, _072893_, _072897_);
  xor g_129665_(_067840_, _072894_, _072898_);
  or g_129666_(_067804_, _072898_, _072899_);
  xor g_129667_(_067804_, _072897_, _072900_);
  or g_129668_(_067767_, _072900_, _072901_);
  not g_129669_(_072901_, _072902_);
  xor g_129670_(_067767_, _072900_, _072903_);
  not g_129671_(_072903_, _072904_);
  or g_129672_(_067731_, _072904_, _072905_);
  xor g_129673_(_067731_, _072903_, _072906_);
  not g_129674_(_072906_, _072908_);
  or g_129675_(_067695_, _072906_, _072909_);
  xor g_129676_(_067695_, _072906_, _072910_);
  xor g_129677_(_067695_, _072908_, _072911_);
  or g_129678_(_067658_, _072911_, _072912_);
  not g_129679_(_072912_, _072913_);
  xor g_129680_(_067658_, _072910_, _072914_);
  not g_129681_(_072914_, _072915_);
  or g_129682_(_067622_, _072914_, _072916_);
  xor g_129683_(_067622_, _072914_, _072917_);
  xor g_129684_(_067622_, _072915_, _072919_);
  or g_129685_(_067586_, _072919_, _072920_);
  xor g_129686_(_067586_, _072917_, _072921_);
  not g_129687_(_072921_, _072922_);
  or g_129688_(_067549_, _072921_, _072923_);
  xor g_129689_(_067549_, _072921_, _072924_);
  xor g_129690_(_067549_, _072922_, _072925_);
  or g_129691_(_067513_, _072925_, _072926_);
  xor g_129692_(_067513_, _072924_, _072927_);
  or g_129693_(_067477_, _072927_, _072928_);
  xor g_129694_(_067477_, _072927_, _072930_);
  not g_129695_(_072930_, _072931_);
  or g_129696_(_067441_, _072931_, _072932_);
  not g_129697_(_072932_, _072933_);
  xor g_129698_(_067441_, _072930_, _072934_);
  not g_129699_(_072934_, _072935_);
  or g_129700_(_067404_, _072934_, _072936_);
  xor g_129701_(_067404_, _072934_, _072937_);
  xor g_129702_(_067404_, _072935_, _072938_);
  or g_129703_(_067368_, _072938_, _072939_);
  xor g_129704_(_067368_, _072937_, _072941_);
  not g_129705_(_072941_, _072942_);
  or g_129706_(_067332_, _072941_, _072943_);
  xor g_129707_(_067332_, _072941_, _072944_);
  xor g_129708_(_067332_, _072942_, _072945_);
  or g_129709_(_067295_, _072945_, _072946_);
  xor g_129710_(_067295_, _072944_, _072947_);
  or g_129711_(_067258_, _072947_, _072948_);
  not g_129712_(_072948_, _072949_);
  xor g_129713_(_067259_, _072947_, _072950_);
  not g_129714_(_072950_, _072952_);
  and g_129715_(_067222_, _072952_, _072953_);
  or g_129716_(_067221_, _072950_, _072954_);
  xor g_129717_(_067222_, _072950_, _072955_);
  or g_129718_(_067184_, _072955_, _072956_);
  xor g_129719_(_067184_, _072955_, _072957_);
  not g_129720_(_072957_, _072958_);
  or g_129721_(_067148_, _072958_, _072959_);
  xor g_129722_(_067148_, _072957_, _072960_);
  not g_129723_(_072960_, _072961_);
  or g_129724_(_067112_, _072960_, _072963_);
  xor g_129725_(_067112_, _072960_, _072964_);
  xor g_129726_(_067112_, _072961_, _072965_);
  and g_129727_(_067075_, _072964_, _072966_);
  or g_129728_(_067074_, _072965_, _072967_);
  xor g_129729_(_067074_, _072964_, _072968_);
  or g_129730_(_067037_, _072968_, _072969_);
  xor g_129731_(_067038_, _072968_, _072970_);
  or g_129732_(_066999_, _072970_, _072971_);
  xor g_129733_(_067001_, _072970_, _072972_);
  or g_129734_(_066962_, _072972_, _072974_);
  xor g_129735_(_066963_, _072972_, _072975_);
  or g_129736_(_066926_, _072975_, _072976_);
  not g_129737_(_072976_, _072977_);
  xor g_129738_(_066926_, _072975_, _072978_);
  not g_129739_(_072978_, _072979_);
  or g_129740_(_066889_, _072979_, _072980_);
  not g_129741_(_072980_, _072981_);
  xor g_129742_(_066889_, _072978_, _072982_);
  or g_129743_(_066853_, _072982_, _072983_);
  xor g_129744_(_066853_, _072982_, _072985_);
  not g_129745_(_072985_, _072986_);
  or g_129746_(_066817_, _072986_, _072987_);
  xor g_129747_(_066817_, _072985_, _072988_);
  not g_129748_(_072988_, _072989_);
  or g_129749_(_066781_, _072988_, _072990_);
  xor g_129750_(_066781_, _072988_, _072991_);
  xor g_129751_(_066781_, _072989_, _072992_);
  or g_129752_(_066744_, _072992_, _072993_);
  xor g_129753_(_066744_, _072991_, _072994_);
  not g_129754_(_072994_, _072996_);
  or g_129755_(_066708_, _072994_, _072997_);
  xor g_129756_(_066708_, _072994_, _072998_);
  xor g_129757_(_066708_, _072996_, _072999_);
  or g_129758_(_066672_, _072999_, _073000_);
  xor g_129759_(_066672_, _072998_, _073001_);
  or g_129760_(_066634_, _073001_, _073002_);
  xor g_129761_(_066635_, _073001_, _073003_);
  not g_129762_(_073003_, _073004_);
  or g_129763_(_066598_, _073003_, _073005_);
  xor g_129764_(_066598_, _073003_, _073007_);
  xor g_129765_(_066598_, _073004_, _073008_);
  or g_129766_(_066562_, _073008_, _073009_);
  xor g_129767_(_066562_, _073007_, _073010_);
  not g_129768_(_073010_, _073011_);
  or g_129769_(_066525_, _073010_, _073012_);
  xor g_129770_(_066525_, _073010_, _073013_);
  xor g_129771_(_066525_, _073011_, _073014_);
  or g_129772_(_066489_, _073014_, _073015_);
  xor g_129773_(_066489_, _073013_, _073016_);
  or g_129774_(_066453_, _073016_, _073018_);
  not g_129775_(_073018_, _073019_);
  and g_129776_(_066453_, _073016_, _073020_);
  xor g_129777_(_066453_, _073016_, _073021_);
  or g_129778_(_073019_, _073020_, _073022_);
  or g_129779_(_066416_, _073022_, _073023_);
  and g_129780_(_066416_, _073022_, _073024_);
  xor g_129781_(_066416_, _073021_, _073025_);
  or g_129782_(_066379_, _073024_, _073026_);
  or g_129783_(_066379_, _073025_, _073027_);
  xor g_129784_(_066380_, _073025_, _073029_);
  or g_129785_(_066343_, _073029_, _073030_);
  not g_129786_(_073030_, _073031_);
  and g_129787_(_066343_, _073029_, _073032_);
  xor g_129788_(_066343_, _073029_, _073033_);
  or g_129789_(_073031_, _073032_, _073034_);
  or g_129790_(_066306_, _073034_, _073035_);
  not g_129791_(_073035_, _073036_);
  xor g_129792_(_066306_, _073033_, _073037_);
  not g_129793_(_073037_, _073038_);
  or g_129794_(_066270_, _073037_, _073040_);
  xor g_129795_(_066270_, _073037_, _073041_);
  xor g_129796_(_066270_, _073038_, _073042_);
  or g_129797_(_066234_, _073042_, _073043_);
  xor g_129798_(_066234_, _073041_, _073044_);
  or g_129799_(_066196_, _073044_, _073045_);
  xor g_129800_(_066198_, _073044_, _073046_);
  or g_129801_(_066159_, _073046_, _073047_);
  xor g_129802_(_066160_, _073046_, _073048_);
  not g_129803_(_073048_, _073049_);
  or g_129804_(_066123_, _073048_, _073051_);
  xor g_129805_(_066123_, _073048_, _073052_);
  xor g_129806_(_066123_, _073049_, _073053_);
  or g_129807_(_066086_, _073053_, _073054_);
  xor g_129808_(_066086_, _073052_, _073055_);
  or g_129809_(_066049_, _073055_, _073056_);
  xor g_129810_(_066050_, _073055_, _073057_);
  or g_129811_(_066012_, _073057_, _073058_);
  not g_129812_(_073058_, _073059_);
  xor g_129813_(_066013_, _073057_, _073060_);
  not g_129814_(_073060_, _073062_);
  or g_129815_(_065975_, _073060_, _073063_);
  xor g_129816_(_065975_, _073060_, _073064_);
  xor g_129817_(_065975_, _073062_, _073065_);
  or g_129818_(_065939_, _073065_, _073066_);
  xor g_129819_(_065939_, _073064_, _073067_);
  not g_129820_(_073067_, _073068_);
  or g_129821_(_065903_, _073067_, _073069_);
  xor g_129822_(_065903_, _073067_, _073070_);
  xor g_129823_(_065903_, _073068_, _073071_);
  or g_129824_(_065866_, _073071_, _073073_);
  xor g_129825_(_065866_, _073070_, _073074_);
  or g_129826_(_065829_, _073074_, _073075_);
  xor g_129827_(_065830_, _073074_, _073076_);
  not g_129828_(_073076_, _073077_);
  or g_129829_(_065793_, _073076_, _073078_);
  xor g_129830_(_065793_, _073076_, _073079_);
  xor g_129831_(_065793_, _073077_, _073080_);
  or g_129832_(_065756_, _073080_, _073081_);
  xor g_129833_(_065756_, _073079_, _073082_);
  or g_129834_(_065719_, _073082_, _073084_);
  xor g_129835_(_065720_, _073082_, _073085_);
  not g_129836_(_073085_, _073086_);
  or g_129837_(_065683_, _073085_, _073087_);
  xor g_129838_(_065683_, _073085_, _073088_);
  xor g_129839_(_065683_, _073086_, _073089_);
  or g_129840_(_065646_, _073089_, _073090_);
  xor g_129841_(_065646_, _073088_, _073091_);
  or g_129842_(_065610_, _073091_, _073092_);
  not g_129843_(_073092_, _073093_);
  xor g_129844_(_065610_, _073091_, _073095_);
  not g_129845_(_073095_, _073096_);
  or g_129846_(_065574_, _073096_, _073097_);
  xor g_129847_(_065574_, _073095_, _073098_);
  not g_129848_(_073098_, _073099_);
  or g_129849_(_065538_, _073098_, _073100_);
  xor g_129850_(_065538_, _073098_, _073101_);
  xor g_129851_(_065538_, _073099_, _073102_);
  or g_129852_(_065501_, _073102_, _073103_);
  xor g_129853_(_065501_, _073101_, _073104_);
  or g_129854_(_065464_, _073104_, _073106_);
  not g_129855_(_073106_, _073107_);
  xor g_129856_(_065465_, _073104_, _073108_);
  or g_129857_(_065428_, _073108_, _073109_);
  xor g_129858_(_065428_, _073108_, _073110_);
  not g_129859_(_073110_, _073111_);
  and g_129860_(_065391_, _073110_, _073112_);
  or g_129861_(_065390_, _073111_, _073113_);
  xor g_129862_(_065390_, _073110_, _073114_);
  or g_129863_(_065353_, _073114_, _073115_);
  not g_129864_(_073115_, _073117_);
  xor g_129865_(_065354_, _073114_, _073118_);
  or g_129866_(_065316_, _073118_, _073119_);
  xor g_129867_(_065316_, _073118_, _073120_);
  not g_129868_(_073120_, _073121_);
  or g_129869_(_065280_, _073121_, _073122_);
  xor g_129870_(_065280_, _073120_, _073123_);
  or g_129871_(_065243_, _073123_, _073124_);
  xor g_129872_(_065244_, _073123_, _073125_);
  not g_129873_(_073125_, _073126_);
  or g_129874_(_065206_, _073125_, _073128_);
  xor g_129875_(_065206_, _073125_, _073129_);
  xor g_129876_(_065206_, _073126_, _073130_);
  or g_129877_(_065170_, _073130_, _073131_);
  not g_129878_(_073131_, _073132_);
  xor g_129879_(_065170_, _073129_, _073133_);
  or g_129880_(_065134_, _073133_, _073134_);
  not g_129881_(_073134_, _073135_);
  xor g_129882_(_065134_, _073133_, _073136_);
  not g_129883_(_073136_, _073137_);
  or g_129884_(_065098_, _073137_, _073139_);
  not g_129885_(_073139_, _073140_);
  xor g_129886_(_065098_, _073136_, _073141_);
  not g_129887_(_073141_, _073142_);
  or g_129888_(_065061_, _073141_, _073143_);
  xor g_129889_(_065061_, _073141_, _073144_);
  xor g_129890_(_065061_, _073142_, _073145_);
  or g_129891_(_065025_, _073145_, _073146_);
  xor g_129892_(_065025_, _073144_, _073147_);
  or g_129893_(_064989_, _073147_, _073148_);
  xor g_129894_(_064989_, _073147_, _073150_);
  not g_129895_(_073150_, _073151_);
  or g_129896_(_064952_, _073151_, _073152_);
  xor g_129897_(_064952_, _073150_, _073153_);
  or g_129898_(_064915_, _073153_, _073154_);
  xor g_129899_(_064916_, _073153_, _073155_);
  or g_129900_(_064878_, _073155_, _073156_);
  xor g_129901_(_064879_, _073155_, _073157_);
  or g_129902_(_064840_, _073157_, _073158_);
  xor g_129903_(_064841_, _073157_, _073159_);
  not g_129904_(_073159_, _073161_);
  or g_129905_(_064804_, _073159_, _073162_);
  xor g_129906_(_064804_, _073159_, _073163_);
  xor g_129907_(_064804_, _073161_, _073164_);
  or g_129908_(_064768_, _073164_, _073165_);
  xor g_129909_(_064768_, _073163_, _073166_);
  or g_129910_(_064731_, _073166_, _073167_);
  xor g_129911_(_064731_, _073166_, _073168_);
  not g_129912_(_073168_, _073169_);
  or g_129913_(_064695_, _073169_, _073170_);
  not g_129914_(_073170_, _073172_);
  xor g_129915_(_064695_, _073168_, _073173_);
  or g_129916_(_064659_, _073173_, _073174_);
  not g_129917_(_073174_, _073175_);
  and g_129918_(_064659_, _073173_, _073176_);
  xor g_129919_(_064659_, _073173_, _073177_);
  or g_129920_(_073175_, _073176_, _073178_);
  or g_129921_(_064622_, _073178_, _073179_);
  xor g_129922_(_064622_, _073177_, _073180_);
  or g_129923_(_064586_, _073180_, _073181_);
  not g_129924_(_073181_, _073183_);
  xor g_129925_(_064585_, _073180_, _073184_);
  or g_129926_(_064545_, _073184_, _073185_);
  xor g_129927_(_064546_, _073184_, _073186_);
  not g_129928_(_073186_, _073187_);
  or g_129929_(_064509_, _073186_, _073188_);
  xor g_129930_(_064509_, _073186_, _073189_);
  xor g_129931_(_064509_, _073187_, _073190_);
  or g_129932_(_064473_, _073190_, _073191_);
  xor g_129933_(_064473_, _073189_, _073192_);
  or g_129934_(_064436_, _073192_, _073194_);
  xor g_129935_(_064436_, _073192_, _073195_);
  not g_129936_(_073195_, _073196_);
  or g_129937_(_064400_, _073196_, _073197_);
  not g_129938_(_073197_, _073198_);
  xor g_129939_(_064400_, _073195_, _073199_);
  or g_129940_(_064363_, _073199_, _073200_);
  not g_129941_(_073200_, _073201_);
  xor g_129942_(_064364_, _073199_, _073202_);
  or g_129943_(_064326_, _073202_, _073203_);
  not g_129944_(_073203_, _073205_);
  and g_129945_(_064326_, _073202_, _073206_);
  xor g_129946_(_064326_, _073202_, _073207_);
  or g_129947_(_073205_, _073206_, _073208_);
  or g_129948_(_064290_, _073208_, _073209_);
  xor g_129949_(_064290_, _073207_, _073210_);
  or g_129950_(_064254_, _073210_, _073211_);
  not g_129951_(_073211_, _073212_);
  xor g_129952_(_064254_, _073210_, _073213_);
  not g_129953_(_073213_, _073214_);
  or g_129954_(_064218_, _073214_, _073216_);
  not g_129955_(_073216_, _073217_);
  xor g_129956_(_064218_, _073213_, _073218_);
  or g_129957_(_064181_, _073218_, _073219_);
  not g_129958_(_073219_, _073220_);
  and g_129959_(_064181_, _073218_, _073221_);
  xor g_129960_(_064181_, _073218_, _073222_);
  or g_129961_(_073220_, _073221_, _073223_);
  or g_129962_(_064144_, _073223_, _073224_);
  xor g_129963_(_064145_, _073222_, _073225_);
  xor g_129964_(_064144_, _073222_, _073227_);
  or g_129965_(_064108_, _073227_, _073228_);
  xor g_129966_(_064108_, _073225_, _073229_);
  not g_129967_(_073229_, _073230_);
  or g_129968_(_064071_, _073229_, _073231_);
  xor g_129969_(_064071_, _073229_, _073232_);
  xor g_129970_(_064071_, _073230_, _073233_);
  or g_129971_(_064035_, _073233_, _073234_);
  xor g_129972_(_064035_, _073232_, _073235_);
  not g_129973_(_073235_, _073236_);
  or g_129974_(_063999_, _073235_, _073238_);
  xor g_129975_(_063999_, _073235_, _073239_);
  xor g_129976_(_063999_, _073236_, _073240_);
  or g_129977_(_063962_, _073240_, _073241_);
  xor g_129978_(_063962_, _073239_, _073242_);
  or g_129979_(_063926_, _073242_, _073243_);
  not g_129980_(_073243_, _073244_);
  and g_129981_(_063926_, _073242_, _073245_);
  xor g_129982_(_063926_, _073242_, _073246_);
  or g_129983_(_073244_, _073245_, _073247_);
  or g_129984_(_063890_, _073247_, _073249_);
  xor g_129985_(_063890_, _073246_, _073250_);
  not g_129986_(_073250_, _073251_);
  or g_129987_(_063853_, _073250_, _073252_);
  xor g_129988_(_063853_, _073250_, _073253_);
  xor g_129989_(_063853_, _073251_, _073254_);
  or g_129990_(_063817_, _073254_, _073255_);
  xor g_129991_(_063817_, _073253_, _073256_);
  or g_129992_(_063780_, _073256_, _073257_);
  xor g_129993_(_063781_, _073256_, _073258_);
  not g_129994_(_073258_, _073260_);
  or g_129995_(_063743_, _073258_, _073261_);
  xor g_129996_(_063743_, _073258_, _073262_);
  xor g_129997_(_063743_, _073260_, _073263_);
  or g_129998_(_063707_, _073263_, _073264_);
  xor g_129999_(_063707_, _073262_, _073265_);
  or g_130000_(_063670_, _073265_, _073266_);
  xor g_130001_(_063671_, _073265_, _073267_);
  or g_130002_(_063632_, _073267_, _073268_);
  xor g_130003_(_063633_, _073267_, _073269_);
  or g_130004_(_063596_, _073269_, _073271_);
  not g_130005_(_073271_, _073272_);
  and g_130006_(_063596_, _073269_, _073273_);
  xor g_130007_(_063596_, _073269_, _073274_);
  or g_130008_(_073272_, _073273_, _073275_);
  or g_130009_(_063560_, _073275_, _073276_);
  xor g_130010_(_063560_, _073274_, _073277_);
  or g_130011_(_063522_, _073277_, _073278_);
  not g_130012_(_073278_, _073279_);
  xor g_130013_(_063523_, _073277_, _073280_);
  or g_130014_(_063485_, _073280_, _073282_);
  xor g_130015_(_063486_, _073280_, _073283_);
  not g_130016_(_073283_, _073284_);
  or g_130017_(_063449_, _073283_, _073285_);
  xor g_130018_(_063449_, _073283_, _073286_);
  xor g_130019_(_063449_, _073284_, _073287_);
  or g_130020_(_063412_, _073287_, _073288_);
  xor g_130021_(_063412_, _073286_, _073289_);
  or g_130022_(_063376_, _073289_, _073290_);
  not g_130023_(_073290_, _073291_);
  and g_130024_(_063376_, _073289_, _073293_);
  xor g_130025_(_063376_, _073289_, _073294_);
  or g_130026_(_073291_, _073293_, _073295_);
  or g_130027_(_063340_, _073295_, _073296_);
  xor g_130028_(_063340_, _073294_, _073297_);
  or g_130029_(_063302_, _073297_, _073298_);
  not g_130030_(_073298_, _073299_);
  xor g_130031_(_063303_, _073297_, _073300_);
  not g_130032_(_073300_, _073301_);
  or g_130033_(_063266_, _073300_, _073302_);
  xor g_130034_(_063266_, _073300_, _073304_);
  xor g_130035_(_063266_, _073301_, _073305_);
  or g_130036_(_063230_, _073305_, _073306_);
  xor g_130037_(_063230_, _073304_, _073307_);
  or g_130038_(_063193_, _073307_, _073308_);
  not g_130039_(_073308_, _073309_);
  xor g_130040_(_063192_, _073307_, _073310_);
  or g_130041_(_063153_, _073310_, _073311_);
  xor g_130042_(_063154_, _073310_, _073312_);
  or g_130043_(_063115_, _073312_, _073313_);
  and g_130044_(_063115_, _073312_, _073315_);
  xor g_130045_(_063116_, _073312_, _073316_);
  not g_130046_(_073316_, _073317_);
  or g_130047_(_063079_, _073315_, _073318_);
  or g_130048_(_063079_, _073316_, _073319_);
  xor g_130049_(_063079_, _073316_, _073320_);
  xor g_130050_(_063079_, _073317_, _073321_);
  or g_130051_(_063043_, _073321_, _073322_);
  xor g_130052_(_063043_, _073320_, _073323_);
  or g_130053_(_063005_, _073323_, _073324_);
  xor g_130054_(_063006_, _073323_, _073326_);
  or g_130055_(_062969_, _073326_, _073327_);
  not g_130056_(_073327_, _073328_);
  and g_130057_(_062969_, _073326_, _073329_);
  xor g_130058_(_062969_, _073326_, _073330_);
  or g_130059_(_073328_, _073329_, _073331_);
  or g_130060_(_062933_, _073331_, _073332_);
  xor g_130061_(_062933_, _073330_, _073333_);
  not g_130062_(_073333_, _073334_);
  or g_130063_(_062896_, _073333_, _073335_);
  xor g_130064_(_062896_, _073333_, _073337_);
  xor g_130065_(_062896_, _073334_, _073338_);
  or g_130066_(_062860_, _073338_, _073339_);
  xor g_130067_(_062860_, _073337_, _073340_);
  or g_130068_(_062823_, _073340_, _073341_);
  not g_130069_(_073341_, _073342_);
  xor g_130070_(_062824_, _073340_, _073343_);
  or g_130071_(_062786_, _073343_, _073344_);
  and g_130072_(_062786_, _073343_, _073345_);
  xor g_130073_(_062786_, _073343_, _073346_);
  and g_130074_(_062750_, _073346_, _073348_);
  not g_130075_(_073348_, _073349_);
  or g_130076_(_062749_, _073345_, _073350_);
  xor g_130077_(_062749_, _073346_, _073351_);
  or g_130078_(_062713_, _073351_, _073352_);
  not g_130079_(_073352_, _073353_);
  and g_130080_(_062713_, _073351_, _073354_);
  xor g_130081_(_062713_, _073351_, _073355_);
  or g_130082_(_073353_, _073354_, _073356_);
  or g_130083_(_062676_, _073356_, _073357_);
  xor g_130084_(_062676_, _073355_, _073359_);
  or g_130085_(_062640_, _073359_, _073360_);
  xor g_130086_(_062640_, _073359_, _073361_);
  not g_130087_(_073361_, _073362_);
  and g_130088_(_062604_, _073361_, _073363_);
  or g_130089_(_062603_, _073362_, _073364_);
  xor g_130090_(_062603_, _073361_, _073365_);
  not g_130091_(_073365_, _073366_);
  or g_130092_(_062566_, _073365_, _073367_);
  xor g_130093_(_062566_, _073365_, _073368_);
  xor g_130094_(_062566_, _073366_, _073370_);
  or g_130095_(_062530_, _073370_, _073371_);
  not g_130096_(_073371_, _073372_);
  xor g_130097_(_062530_, _073368_, _073373_);
  not g_130098_(_073373_, _073374_);
  or g_130099_(_062494_, _073373_, _073375_);
  xor g_130100_(_062494_, _073374_, _073376_);
  not g_130101_(_073376_, _073377_);
  or g_130102_(_062458_, _073376_, _073378_);
  xor g_130103_(_062458_, _073376_, _073379_);
  xor g_130104_(_062458_, _073377_, _073381_);
  or g_130105_(_062421_, _073381_, _073382_);
  xor g_130106_(_062421_, _073379_, _073383_);
  not g_130107_(_073383_, _073384_);
  or g_130108_(_062385_, _073383_, _073385_);
  xor g_130109_(_062385_, _073383_, _073386_);
  xor g_130110_(_062385_, _073384_, _073387_);
  or g_130111_(_062349_, _073387_, _073388_);
  xor g_130112_(_062349_, _073387_, _073389_);
  xor g_130113_(_062349_, _073386_, _073390_);
  or g_130114_(_062312_, _073390_, _073392_);
  not g_130115_(_073392_, _073393_);
  xor g_130116_(_062312_, _073389_, _073394_);
  or g_130117_(_062275_, _073394_, _073395_);
  xor g_130118_(_062276_, _073394_, _073396_);
  not g_130119_(_073396_, _073397_);
  or g_130120_(_062239_, _073396_, _073398_);
  xor g_130121_(_062239_, _073396_, _073399_);
  xor g_130122_(_062239_, _073397_, _073400_);
  or g_130123_(_062202_, _073400_, _073401_);
  xor g_130124_(_062202_, _073399_, _073403_);
  or g_130125_(_062166_, _073403_, _073404_);
  not g_130126_(_073404_, _073405_);
  and g_130127_(_062166_, _073403_, _073406_);
  xor g_130128_(_062166_, _073403_, _073407_);
  or g_130129_(_073405_, _073406_, _073408_);
  or g_130130_(_062130_, _073408_, _073409_);
  xor g_130131_(_062130_, _073407_, _073410_);
  or g_130132_(_062093_, _073410_, _073411_);
  xor g_130133_(_062093_, _073410_, _073412_);
  not g_130134_(_073412_, _073414_);
  and g_130135_(_062057_, _073412_, _073415_);
  or g_130136_(_062056_, _073414_, _073416_);
  xor g_130137_(_062056_, _073412_, _073417_);
  not g_130138_(_073417_, _073418_);
  or g_130139_(_062020_, _073417_, _073419_);
  xor g_130140_(_062020_, _073417_, _073420_);
  xor g_130141_(_062020_, _073418_, _073421_);
  or g_130142_(_061983_, _073421_, _073422_);
  not g_130143_(_073422_, _073423_);
  xor g_130144_(_061983_, _073420_, _073425_);
  or g_130145_(_061946_, _073425_, _073426_);
  xor g_130146_(_061947_, _073425_, _073427_);
  not g_130147_(_073427_, _073428_);
  or g_130148_(_061910_, _073427_, _073429_);
  xor g_130149_(_061910_, _073427_, _073430_);
  xor g_130150_(_061910_, _073428_, _073431_);
  or g_130151_(_061873_, _073431_, _073432_);
  xor g_130152_(_061873_, _073430_, _073433_);
  not g_130153_(_073433_, _073434_);
  or g_130154_(_061837_, _073433_, _073436_);
  xor g_130155_(_061837_, _073433_, _073437_);
  xor g_130156_(_061837_, _073434_, _073438_);
  or g_130157_(_061801_, _073438_, _073439_);
  xor g_130158_(_061801_, _073437_, _073440_);
  or g_130159_(_061763_, _073440_, _073441_);
  xor g_130160_(_061765_, _073440_, _073442_);
  or g_130161_(_061726_, _073442_, _073443_);
  xor g_130162_(_061727_, _073442_, _073444_);
  not g_130163_(_073444_, _073445_);
  or g_130164_(_061690_, _073444_, _073447_);
  xor g_130165_(_061690_, _073444_, _073448_);
  xor g_130166_(_061690_, _073445_, _073449_);
  or g_130167_(_061653_, _073449_, _073450_);
  xor g_130168_(_061653_, _073448_, _073451_);
  or g_130169_(_061616_, _073451_, _073452_);
  xor g_130170_(_061617_, _073451_, _073453_);
  or g_130171_(_061579_, _073453_, _073454_);
  xor g_130172_(_061580_, _073453_, _073455_);
  not g_130173_(_073455_, _073456_);
  or g_130174_(_061542_, _073455_, _073458_);
  xor g_130175_(_061542_, _073455_, _073459_);
  xor g_130176_(_061542_, _073456_, _073460_);
  or g_130177_(_061506_, _073460_, _073461_);
  xor g_130178_(_061506_, _073459_, _073462_);
  not g_130179_(_073462_, _073463_);
  or g_130180_(_061470_, _073462_, _073464_);
  xor g_130181_(_061470_, _073462_, _073465_);
  xor g_130182_(_061470_, _073463_, _073466_);
  or g_130183_(_061433_, _073466_, _073467_);
  xor g_130184_(_061433_, _073465_, _073469_);
  or g_130185_(_061397_, _073469_, _073470_);
  not g_130186_(_073470_, _073471_);
  xor g_130187_(_061397_, _073469_, _073472_);
  not g_130188_(_073472_, _073473_);
  or g_130189_(_061361_, _073473_, _073474_);
  xor g_130190_(_061361_, _073472_, _073475_);
  not g_130191_(_073475_, _073476_);
  or g_130192_(_061325_, _073475_, _073477_);
  xor g_130193_(_061325_, _073475_, _073478_);
  xor g_130194_(_061325_, _073476_, _073480_);
  or g_130195_(_061288_, _073480_, _073481_);
  xor g_130196_(_061288_, _073478_, _073482_);
  or g_130197_(_061252_, _073482_, _073483_);
  xor g_130198_(_061252_, _073482_, _073484_);
  not g_130199_(_073484_, _073485_);
  or g_130200_(_061216_, _073485_, _073486_);
  not g_130201_(_073486_, _073487_);
  xor g_130202_(_061216_, _073484_, _073488_);
  or g_130203_(_061178_, _073488_, _073489_);
  xor g_130204_(_061179_, _073488_, _073491_);
  or g_130205_(_061141_, _073491_, _073492_);
  xor g_130206_(_061142_, _073491_, _073493_);
  not g_130207_(_073493_, _073494_);
  or g_130208_(_061105_, _073493_, _073495_);
  xor g_130209_(_061105_, _073493_, _073496_);
  xor g_130210_(_061105_, _073494_, _073497_);
  or g_130211_(_061068_, _073497_, _073498_);
  xor g_130212_(_061068_, _073496_, _073499_);
  or g_130213_(_061032_, _073499_, _073500_);
  xor g_130214_(_061032_, _073499_, _073502_);
  not g_130215_(_073502_, _073503_);
  or g_130216_(_060996_, _073503_, _073504_);
  xor g_130217_(_060996_, _073502_, _073505_);
  not g_130218_(_073505_, _073506_);
  or g_130219_(_060959_, _073505_, _073507_);
  xor g_130220_(_060959_, _073505_, _073508_);
  xor g_130221_(_060959_, _073506_, _073509_);
  or g_130222_(_060923_, _073509_, _073510_);
  xor g_130223_(_060923_, _073508_, _073511_);
  or g_130224_(_060887_, _073511_, _073513_);
  not g_130225_(_073513_, _073514_);
  xor g_130226_(_060887_, _073511_, _073515_);
  not g_130227_(_073515_, _073516_);
  or g_130228_(_060850_, _073516_, _073517_);
  xor g_130229_(_060850_, _073515_, _073518_);
  or g_130230_(_060814_, _073518_, _073519_);
  xor g_130231_(_060814_, _073518_, _073520_);
  not g_130232_(_073520_, _073521_);
  or g_130233_(_060778_, _073521_, _073522_);
  xor g_130234_(_060778_, _073520_, _073524_);
  or g_130235_(_060740_, _073524_, _073525_);
  xor g_130236_(_060742_, _073524_, _073526_);
  or g_130237_(_060704_, _073526_, _073527_);
  xor g_130238_(_060704_, _073526_, _073528_);
  not g_130239_(_073528_, _073529_);
  or g_130240_(_060668_, _073529_, _073530_);
  xor g_130241_(_060668_, _073528_, _073531_);
  or g_130242_(_060630_, _073531_, _073532_);
  xor g_130243_(_060632_, _073531_, _073533_);
  not g_130244_(_073533_, _073535_);
  or g_130245_(_060594_, _073533_, _073536_);
  xor g_130246_(_060594_, _073533_, _073537_);
  xor g_130247_(_060594_, _073535_, _073538_);
  or g_130248_(_060558_, _073538_, _073539_);
  xor g_130249_(_060558_, _073537_, _073540_);
  or g_130250_(_060520_, _073540_, _073541_);
  xor g_130251_(_060522_, _073540_, _073542_);
  not g_130252_(_073542_, _073543_);
  or g_130253_(_060484_, _073542_, _073544_);
  xor g_130254_(_060484_, _073542_, _073546_);
  xor g_130255_(_060484_, _073543_, _073547_);
  or g_130256_(_060448_, _073547_, _073548_);
  xor g_130257_(_060448_, _073546_, _073549_);
  or g_130258_(_060410_, _073549_, _073550_);
  not g_130259_(_073550_, _073551_);
  xor g_130260_(_060412_, _073549_, _073552_);
  or g_130261_(_060373_, _073552_, _073553_);
  xor g_130262_(_060374_, _073552_, _073554_);
  or g_130263_(_060336_, _073554_, _073555_);
  xor g_130264_(_060337_, _073554_, _073557_);
  or g_130265_(_060299_, _073557_, _073558_);
  not g_130266_(_073558_, _073559_);
  and g_130267_(_060299_, _073557_, _073560_);
  xor g_130268_(_060299_, _073557_, _073561_);
  or g_130269_(_073559_, _073560_, _073562_);
  or g_130270_(_060263_, _073562_, _073563_);
  xor g_130271_(_060263_, _073561_, _073564_);
  or g_130272_(_060226_, _073564_, _073565_);
  xor g_130273_(_060227_, _073564_, _073566_);
  or g_130274_(_060189_, _073566_, _073568_);
  xor g_130275_(_060189_, _073566_, _073569_);
  not g_130276_(_073569_, _073570_);
  or g_130277_(_060153_, _073570_, _073571_);
  xor g_130278_(_060153_, _073569_, _073572_);
  or g_130279_(_060117_, _073572_, _073573_);
  not g_130280_(_073573_, _073574_);
  and g_130281_(_060117_, _073572_, _073575_);
  xor g_130282_(_060117_, _073572_, _073576_);
  or g_130283_(_073574_, _073575_, _073577_);
  or g_130284_(_060080_, _073577_, _073579_);
  xor g_130285_(_060080_, _073576_, _073580_);
  or g_130286_(_060043_, _073580_, _073581_);
  xor g_130287_(_060044_, _073580_, _073582_);
  or g_130288_(_060007_, _073582_, _073583_);
  xor g_130289_(_060007_, _073582_, _073584_);
  not g_130290_(_073584_, _073585_);
  or g_130291_(_059970_, _073585_, _073586_);
  xor g_130292_(_059970_, _073584_, _073587_);
  or g_130293_(_059934_, _073587_, _073588_);
  not g_130294_(_073588_, _073590_);
  xor g_130295_(_059934_, _073587_, _073591_);
  not g_130296_(_073591_, _073592_);
  or g_130297_(_059898_, _073592_, _073593_);
  not g_130298_(_073593_, _073594_);
  xor g_130299_(_059898_, _073591_, _073595_);
  or g_130300_(_059860_, _073595_, _073596_);
  xor g_130301_(_059862_, _073595_, _073597_);
  or g_130302_(_059824_, _073597_, _073598_);
  not g_130303_(_073598_, _073599_);
  xor g_130304_(_059824_, _073597_, _073601_);
  not g_130305_(_073601_, _073602_);
  or g_130306_(_059788_, _073602_, _073603_);
  xor g_130307_(_059788_, _073601_, _073604_);
  or g_130308_(_059750_, _073604_, _073605_);
  xor g_130309_(_059752_, _073604_, _073606_);
  not g_130310_(_073606_, _073607_);
  or g_130311_(_059714_, _073606_, _073608_);
  xor g_130312_(_059714_, _073606_, _073609_);
  xor g_130313_(_059714_, _073607_, _073610_);
  or g_130314_(_059678_, _073610_, _073612_);
  not g_130315_(_073612_, _073613_);
  xor g_130316_(_059678_, _073609_, _073614_);
  or g_130317_(_059640_, _073614_, _073615_);
  xor g_130318_(_059640_, _073614_, _073616_);
  xor g_130319_(_059642_, _073614_, _073617_);
  and g_130320_(_059604_, _073616_, _073618_);
  or g_130321_(_059603_, _073617_, _073619_);
  and g_130322_(_059603_, _073617_, _073620_);
  xor g_130323_(_059604_, _073616_, _073621_);
  or g_130324_(_059567_, _073620_, _073623_);
  or g_130325_(_073618_, _073623_, _073624_);
  xor g_130326_(_059567_, _073621_, _073625_);
  or g_130327_(_059530_, _073625_, _073626_);
  xor g_130328_(_059530_, _073625_, _073627_);
  not g_130329_(_073627_, _073628_);
  or g_130330_(_059494_, _073628_, _073629_);
  xor g_130331_(_059494_, _073627_, _073630_);
  or g_130332_(_059458_, _073630_, _073631_);
  xor g_130333_(_059458_, _073630_, _073632_);
  not g_130334_(_073632_, _073634_);
  or g_130335_(_059422_, _073634_, _073635_);
  not g_130336_(_073635_, _073636_);
  xor g_130337_(_059422_, _073632_, _073637_);
  not g_130338_(_073637_, _073638_);
  or g_130339_(_059385_, _073637_, _073639_);
  not g_130340_(_073639_, _073640_);
  xor g_130341_(_059385_, _073638_, _073641_);
  not g_130342_(_073641_, _073642_);
  or g_130343_(_059349_, _073641_, _073643_);
  xor g_130344_(_059349_, _073641_, _073645_);
  xor g_130345_(_059349_, _073642_, _073646_);
  or g_130346_(_059313_, _073646_, _073647_);
  xor g_130347_(_059313_, _073645_, _073648_);
  not g_130348_(_073648_, _073649_);
  or g_130349_(_059276_, _073648_, _073650_);
  xor g_130350_(_059276_, _073648_, _073651_);
  xor g_130351_(_059276_, _073649_, _073652_);
  or g_130352_(_059240_, _073652_, _073653_);
  xor g_130353_(_059240_, _073651_, _073654_);
  or g_130354_(_059203_, _073654_, _073656_);
  xor g_130355_(_059204_, _073654_, _073657_);
  or g_130356_(_059165_, _073657_, _073658_);
  xor g_130357_(_059166_, _073657_, _073659_);
  or g_130358_(_059129_, _073659_, _073660_);
  not g_130359_(_073660_, _073661_);
  and g_130360_(_059129_, _073659_, _073662_);
  xor g_130361_(_059129_, _073659_, _073663_);
  or g_130362_(_073661_, _073662_, _073664_);
  or g_130363_(_059093_, _073664_, _073665_);
  xor g_130364_(_059093_, _073663_, _073667_);
  not g_130365_(_073667_, _073668_);
  or g_130366_(_059056_, _073667_, _073669_);
  xor g_130367_(_059056_, _073667_, _073670_);
  xor g_130368_(_059056_, _073668_, _073671_);
  or g_130369_(_059020_, _073671_, _073672_);
  xor g_130370_(_059020_, _073670_, _073673_);
  or g_130371_(_058983_, _073673_, _073674_);
  xor g_130372_(_058984_, _073673_, _073675_);
  not g_130373_(_073675_, _073676_);
  or g_130374_(_058946_, _073675_, _073678_);
  not g_130375_(_073678_, _073679_);
  xor g_130376_(_058946_, _073676_, _073680_);
  or g_130377_(_058909_, _073680_, _073681_);
  xor g_130378_(_058909_, _073680_, _073682_);
  xor g_130379_(_058910_, _073680_, _073683_);
  and g_130380_(_058873_, _073682_, _073684_);
  or g_130381_(_058872_, _073683_, _073685_);
  xor g_130382_(_058872_, _073682_, _073686_);
  or g_130383_(_058834_, _073686_, _073687_);
  not g_130384_(_073687_, _073689_);
  xor g_130385_(_058835_, _073686_, _073690_);
  or g_130386_(_058798_, _073690_, _073691_);
  xor g_130387_(_058798_, _073690_, _073692_);
  not g_130388_(_073692_, _073693_);
  or g_130389_(_058762_, _073693_, _073694_);
  not g_130390_(_073694_, _073695_);
  xor g_130391_(_058762_, _073692_, _073696_);
  not g_130392_(_073696_, _073697_);
  or g_130393_(_058725_, _073696_, _073698_);
  xor g_130394_(_058725_, _073696_, _073700_);
  xor g_130395_(_058725_, _073697_, _073701_);
  or g_130396_(_058689_, _073701_, _073702_);
  xor g_130397_(_058689_, _073700_, _073703_);
  or g_130398_(_058652_, _073703_, _073704_);
  xor g_130399_(_058653_, _073703_, _073705_);
  not g_130400_(_073705_, _073706_);
  or g_130401_(_058615_, _073705_, _073707_);
  xor g_130402_(_058615_, _073705_, _073708_);
  xor g_130403_(_058615_, _073706_, _073709_);
  or g_130404_(_058579_, _073709_, _073711_);
  xor g_130405_(_058579_, _073708_, _073712_);
  or g_130406_(_058542_, _073712_, _073713_);
  xor g_130407_(_058542_, _073712_, _073714_);
  xor g_130408_(_058543_, _073712_, _073715_);
  or g_130409_(_058505_, _073715_, _073716_);
  xor g_130410_(_058505_, _073714_, _073717_);
  or g_130411_(_058469_, _073717_, _073718_);
  not g_130412_(_073718_, _073719_);
  and g_130413_(_058469_, _073717_, _073720_);
  xor g_130414_(_058469_, _073717_, _073722_);
  or g_130415_(_073719_, _073720_, _073723_);
  or g_130416_(_058433_, _073723_, _073724_);
  not g_130417_(_073724_, _073725_);
  xor g_130418_(_058433_, _073722_, _073726_);
  not g_130419_(_073726_, _073727_);
  or g_130420_(_058396_, _073726_, _073728_);
  xor g_130421_(_058396_, _073726_, _073729_);
  xor g_130422_(_058396_, _073727_, _073730_);
  or g_130423_(_058360_, _073730_, _073731_);
  xor g_130424_(_058360_, _073729_, _073733_);
  not g_130425_(_073733_, _073734_);
  or g_130426_(_058324_, _073733_, _073735_);
  xor g_130427_(_058324_, _073734_, _073736_);
  or g_130428_(_058286_, _073736_, _073737_);
  xor g_130429_(_058287_, _073736_, _073738_);
  or g_130430_(_058250_, _073738_, _073739_);
  xor g_130431_(_058250_, _073738_, _073740_);
  not g_130432_(_073740_, _073741_);
  or g_130433_(_058214_, _073741_, _073742_);
  not g_130434_(_073742_, _073744_);
  xor g_130435_(_058214_, _073740_, _073745_);
  or g_130436_(_058176_, _073745_, _073746_);
  xor g_130437_(_058177_, _073745_, _073747_);
  not g_130438_(_073747_, _073748_);
  or g_130439_(_058140_, _073747_, _073749_);
  xor g_130440_(_058140_, _073747_, _073750_);
  xor g_130441_(_058140_, _073748_, _073751_);
  or g_130442_(_058104_, _073751_, _073752_);
  xor g_130443_(_058104_, _073750_, _073753_);
  or g_130444_(_058066_, _073753_, _073755_);
  xor g_130445_(_058066_, _073753_, _073756_);
  xor g_130446_(_058067_, _073753_, _073757_);
  or g_130447_(_058030_, _073757_, _073758_);
  xor g_130448_(_058030_, _073756_, _073759_);
  not g_130449_(_073759_, _073760_);
  or g_130450_(_057994_, _073759_, _073761_);
  xor g_130451_(_057994_, _073759_, _073762_);
  xor g_130452_(_057994_, _073760_, _073763_);
  or g_130453_(_057957_, _073763_, _073764_);
  xor g_130454_(_057957_, _073762_, _073766_);
  not g_130455_(_073766_, _073767_);
  or g_130456_(_057921_, _073766_, _073768_);
  xor g_130457_(_057921_, _073766_, _073769_);
  xor g_130458_(_057921_, _073767_, _073770_);
  or g_130459_(_057885_, _073770_, _073771_);
  not g_130460_(_073771_, _073772_);
  xor g_130461_(_057885_, _073769_, _073773_);
  or g_130462_(_057849_, _073773_, _073774_);
  xor g_130463_(_057847_, _073773_, _073775_);
  or g_130464_(_057808_, _073775_, _073777_);
  xor g_130465_(_057809_, _073775_, _073778_);
  or g_130466_(_057772_, _073778_, _073779_);
  xor g_130467_(_057772_, _073778_, _073780_);
  not g_130468_(_073780_, _073781_);
  or g_130469_(_057735_, _073781_, _073782_);
  xor g_130470_(_057735_, _073780_, _073783_);
  not g_130471_(_073783_, _073784_);
  or g_130472_(_057699_, _073783_, _073785_);
  xor g_130473_(_057699_, _073783_, _073786_);
  xor g_130474_(_057699_, _073784_, _073788_);
  or g_130475_(_057663_, _073788_, _073789_);
  xor g_130476_(_057663_, _073786_, _073790_);
  or g_130477_(_057625_, _073790_, _073791_);
  xor g_130478_(_057626_, _073790_, _073792_);
  or g_130479_(_057589_, _073792_, _073793_);
  not g_130480_(_073793_, _073794_);
  and g_130481_(_057589_, _073792_, _073795_);
  xor g_130482_(_057589_, _073792_, _073796_);
  or g_130483_(_073794_, _073795_, _073797_);
  or g_130484_(_057553_, _073797_, _073799_);
  xor g_130485_(_057553_, _073796_, _073800_);
  not g_130486_(_073800_, _073801_);
  or g_130487_(_057516_, _073800_, _073802_);
  xor g_130488_(_057516_, _073800_, _073803_);
  xor g_130489_(_057516_, _073801_, _073804_);
  or g_130490_(_057480_, _073804_, _073805_);
  xor g_130491_(_057480_, _073803_, _073806_);
  or g_130492_(_057444_, _073806_, _073807_);
  not g_130493_(_073807_, _073808_);
  and g_130494_(_057444_, _073806_, _073810_);
  xor g_130495_(_057444_, _073806_, _073811_);
  or g_130496_(_073808_, _073810_, _073812_);
  or g_130497_(_057407_, _073812_, _073813_);
  xor g_130498_(_057407_, _073811_, _073814_);
  not g_130499_(_073814_, _073815_);
  or g_130500_(_057371_, _073814_, _073816_);
  xor g_130501_(_057371_, _073814_, _073817_);
  xor g_130502_(_057371_, _073815_, _073818_);
  or g_130503_(_057335_, _073818_, _073819_);
  not g_130504_(_073819_, _073821_);
  xor g_130505_(_057335_, _073817_, _073822_);
  or g_130506_(_057299_, _073822_, _073823_);
  not g_130507_(_073823_, _073824_);
  and g_130508_(_057299_, _073822_, _073825_);
  xor g_130509_(_057299_, _073822_, _073826_);
  or g_130510_(_073824_, _073825_, _073827_);
  or g_130511_(_057262_, _073827_, _073828_);
  xor g_130512_(_057262_, _073826_, _073829_);
  or g_130513_(_057225_, _073829_, _073830_);
  xor g_130514_(_057226_, _073829_, _073832_);
  or g_130515_(_057187_, _073832_, _073833_);
  xor g_130516_(_057189_, _073832_, _073834_);
  not g_130517_(_073834_, _073835_);
  or g_130518_(_057151_, _073834_, _073836_);
  xor g_130519_(_057151_, _073834_, _073837_);
  xor g_130520_(_057151_, _073835_, _073838_);
  or g_130521_(_057115_, _073838_, _073839_);
  xor g_130522_(_057115_, _073837_, _073840_);
  not g_130523_(_073840_, _073841_);
  or g_130524_(_057079_, _073840_, _073843_);
  xor g_130525_(_057079_, _073841_, _073844_);
  or g_130526_(_057042_, _073844_, _073845_);
  xor g_130527_(_057042_, _073844_, _073846_);
  not g_130528_(_073846_, _073847_);
  or g_130529_(_057006_, _073847_, _073848_);
  xor g_130530_(_057006_, _073846_, _073849_);
  or g_130531_(_056969_, _073849_, _073850_);
  xor g_130532_(_056970_, _073849_, _073851_);
  or g_130533_(_056932_, _073851_, _073852_);
  not g_130534_(_073852_, _073854_);
  xor g_130535_(_056932_, _073851_, _073855_);
  not g_130536_(_073855_, _073856_);
  or g_130537_(_056896_, _073856_, _073857_);
  xor g_130538_(_056896_, _073855_, _073858_);
  or g_130539_(_056859_, _073858_, _073859_);
  xor g_130540_(_056860_, _073858_, _073860_);
  or g_130541_(_056821_, _073860_, _073861_);
  xor g_130542_(_056822_, _073860_, _073862_);
  or g_130543_(_056784_, _073862_, _073863_);
  xor g_130544_(_056785_, _073862_, _073865_);
  or g_130545_(_056746_, _073865_, _073866_);
  xor g_130546_(_056746_, _073865_, _073867_);
  xor g_130547_(_056747_, _073865_, _073868_);
  and g_130548_(_056710_, _073867_, _073869_);
  or g_130549_(_056709_, _073868_, _073870_);
  xor g_130550_(_056709_, _073867_, _073871_);
  or g_130551_(_056672_, _073871_, _073872_);
  not g_130552_(_073872_, _073873_);
  xor g_130553_(_056673_, _073871_, _073874_);
  not g_130554_(_073874_, _073876_);
  or g_130555_(_056635_, _073874_, _073877_);
  xor g_130556_(_056635_, _073874_, _073878_);
  xor g_130557_(_056635_, _073876_, _073879_);
  and g_130558_(_056599_, _073878_, _073880_);
  or g_130559_(_056598_, _073879_, _073881_);
  xor g_130560_(_056598_, _073878_, _073882_);
  or g_130561_(_056562_, _073882_, _073883_);
  not g_130562_(_073883_, _073884_);
  xor g_130563_(_056562_, _073882_, _073885_);
  not g_130564_(_073885_, _073887_);
  or g_130565_(_056525_, _073887_, _073888_);
  xor g_130566_(_056525_, _073885_, _073889_);
  not g_130567_(_073889_, _073890_);
  or g_130568_(_056489_, _073889_, _073891_);
  xor g_130569_(_056489_, _073890_, _073892_);
  not g_130570_(_073892_, _073893_);
  or g_130571_(_056453_, _073892_, _073894_);
  xor g_130572_(_056453_, _073893_, _073895_);
  or g_130573_(_056415_, _073895_, _073896_);
  xor g_130574_(_056416_, _073895_, _073898_);
  or g_130575_(_056378_, _073898_, _073899_);
  not g_130576_(_073899_, _073900_);
  xor g_130577_(_056379_, _073898_, _073901_);
  or g_130578_(_056342_, _073901_, _073902_);
  not g_130579_(_073902_, _073903_);
  and g_130580_(_056342_, _073901_, _073904_);
  xor g_130581_(_056342_, _073901_, _073905_);
  or g_130582_(_073903_, _073904_, _073906_);
  or g_130583_(_056305_, _073906_, _073907_);
  xor g_130584_(_056305_, _073905_, _073909_);
  or g_130585_(_056269_, _073909_, _073910_);
  not g_130586_(_073910_, _073911_);
  xor g_130587_(_056269_, _073909_, _073912_);
  not g_130588_(_073912_, _073913_);
  or g_130589_(_056233_, _073913_, _073914_);
  xor g_130590_(_056233_, _073912_, _073915_);
  not g_130591_(_073915_, _073916_);
  or g_130592_(_056196_, _073915_, _073917_);
  xor g_130593_(_056196_, _073916_, _073918_);
  not g_130594_(_073918_, _073920_);
  or g_130595_(_056160_, _073918_, _073921_);
  xor g_130596_(_056160_, _073918_, _073922_);
  xor g_130597_(_056160_, _073920_, _073923_);
  or g_130598_(_056124_, _073923_, _073924_);
  xor g_130599_(_056124_, _073922_, _073925_);
  not g_130600_(_073925_, _073926_);
  or g_130601_(_056087_, _073925_, _073927_);
  xor g_130602_(_056087_, _073925_, _073928_);
  xor g_130603_(_056087_, _073926_, _073929_);
  or g_130604_(_056051_, _073929_, _073931_);
  xor g_130605_(_056051_, _073928_, _073932_);
  not g_130606_(_073932_, _073933_);
  or g_130607_(_056015_, _073932_, _073934_);
  xor g_130608_(_056015_, _073932_, _073935_);
  xor g_130609_(_056015_, _073933_, _073936_);
  or g_130610_(_055979_, _073936_, _073937_);
  xor g_130611_(_055979_, _073935_, _073938_);
  not g_130612_(_073938_, _073939_);
  or g_130613_(_055942_, _073938_, _073940_);
  xor g_130614_(_055942_, _073938_, _073942_);
  xor g_130615_(_055942_, _073939_, _073943_);
  or g_130616_(_055906_, _073943_, _073944_);
  xor g_130617_(_055906_, _073942_, _073945_);
  not g_130618_(_073945_, _073946_);
  or g_130619_(_055870_, _073945_, _073947_);
  xor g_130620_(_055870_, _073946_, _073948_);
  not g_130621_(_073948_, _073949_);
  or g_130622_(_055833_, _073948_, _073950_);
  not g_130623_(_073950_, _073951_);
  xor g_130624_(_055833_, _073949_, _073953_);
  not g_130625_(_073953_, _073954_);
  or g_130626_(_055797_, _073953_, _073955_);
  xor g_130627_(_055797_, _073953_, _073956_);
  xor g_130628_(_055797_, _073954_, _073957_);
  or g_130629_(_055761_, _073957_, _073958_);
  xor g_130630_(_055761_, _073956_, _073959_);
  not g_130631_(_073959_, _073960_);
  or g_130632_(_055724_, _073959_, _073961_);
  xor g_130633_(_055724_, _073959_, _073962_);
  xor g_130634_(_055724_, _073960_, _073964_);
  or g_130635_(_055688_, _073964_, _073965_);
  xor g_130636_(_055688_, _073962_, _073966_);
  not g_130637_(_073966_, _073967_);
  or g_130638_(_055652_, _073966_, _073968_);
  xor g_130639_(_055652_, _073966_, _073969_);
  xor g_130640_(_055652_, _073967_, _073970_);
  or g_130641_(_055616_, _073970_, _073971_);
  not g_130642_(_073971_, _073972_);
  xor g_130643_(_055616_, _073969_, _073973_);
  or g_130644_(_055579_, _073973_, _073975_);
  not g_130645_(_073975_, _073976_);
  and g_130646_(_055579_, _073973_, _073977_);
  xor g_130647_(_055579_, _073973_, _073978_);
  or g_130648_(_073976_, _073977_, _073979_);
  or g_130649_(_055543_, _073979_, _073980_);
  not g_130650_(_073980_, _073981_);
  xor g_130651_(_055543_, _073978_, _073982_);
  or g_130652_(_055506_, _073982_, _073983_);
  not g_130653_(_073983_, _073984_);
  xor g_130654_(_055507_, _073982_, _073986_);
  or g_130655_(_055468_, _073986_, _073987_);
  xor g_130656_(_055469_, _073986_, _073988_);
  or g_130657_(_055432_, _073988_, _073989_);
  not g_130658_(_073989_, _073990_);
  and g_130659_(_055432_, _073988_, _073991_);
  xor g_130660_(_055432_, _073988_, _073992_);
  or g_130661_(_073990_, _073991_, _073993_);
  or g_130662_(_055396_, _073993_, _073994_);
  xor g_130663_(_055396_, _073992_, _073995_);
  or g_130664_(_055358_, _073995_, _073997_);
  xor g_130665_(_055359_, _073995_, _073998_);
  or g_130666_(_055321_, _073998_, _073999_);
  xor g_130667_(_055322_, _073998_, _074000_);
  not g_130668_(_074000_, _074001_);
  or g_130669_(_055284_, _074000_, _074002_);
  xor g_130670_(_055284_, _074000_, _074003_);
  xor g_130671_(_055284_, _074001_, _074004_);
  or g_130672_(_055248_, _074004_, _074005_);
  xor g_130673_(_055248_, _074003_, _074006_);
  or g_130674_(_055212_, _074006_, _074008_);
  xor g_130675_(_055212_, _074006_, _074009_);
  not g_130676_(_074009_, _074010_);
  or g_130677_(_055176_, _074010_, _074011_);
  not g_130678_(_074011_, _074012_);
  xor g_130679_(_055176_, _074009_, _074013_);
  not g_130680_(_074013_, _074014_);
  or g_130681_(_055139_, _074013_, _074015_);
  not g_130682_(_074015_, _074016_);
  xor g_130683_(_055139_, _074013_, _074017_);
  xor g_130684_(_055139_, _074014_, _074019_);
  or g_130685_(_055103_, _074019_, _074020_);
  xor g_130686_(_055103_, _074017_, _074021_);
  or g_130687_(_055067_, _074021_, _074022_);
  xor g_130688_(_055067_, _074021_, _074023_);
  not g_130689_(_074023_, _074024_);
  or g_130690_(_055030_, _074024_, _074025_);
  xor g_130691_(_055030_, _074023_, _074026_);
  or g_130692_(_054994_, _074026_, _074027_);
  not g_130693_(_074027_, _074028_);
  and g_130694_(_054994_, _074026_, _074030_);
  xor g_130695_(_054994_, _074026_, _074031_);
  or g_130696_(_074028_, _074030_, _074032_);
  or g_130697_(_054958_, _074032_, _074033_);
  not g_130698_(_074033_, _074034_);
  xor g_130699_(_054958_, _074031_, _074035_);
  or g_130700_(_054921_, _074035_, _074036_);
  not g_130701_(_074036_, _074037_);
  and g_130702_(_054921_, _074035_, _074038_);
  xor g_130703_(_054921_, _074035_, _074039_);
  or g_130704_(_074037_, _074038_, _074041_);
  and g_130705_(_054885_, _074039_, _074042_);
  or g_130706_(_054884_, _074041_, _074043_);
  xor g_130707_(_054885_, _074039_, _074044_);
  xor g_130708_(_054884_, _074039_, _074045_);
  or g_130709_(_054848_, _074045_, _074046_);
  xor g_130710_(_054848_, _074044_, _074047_);
  or g_130711_(_054810_, _074047_, _074048_);
  xor g_130712_(_054811_, _074047_, _074049_);
  not g_130713_(_074049_, _074050_);
  or g_130714_(_054774_, _074049_, _074052_);
  xor g_130715_(_054774_, _074049_, _074053_);
  xor g_130716_(_054774_, _074050_, _074054_);
  or g_130717_(_054738_, _074054_, _074055_);
  xor g_130718_(_054738_, _074053_, _074056_);
  not g_130719_(_074056_, _074057_);
  or g_130720_(_054701_, _074056_, _074058_);
  xor g_130721_(_054701_, _074056_, _074059_);
  xor g_130722_(_054701_, _074057_, _074060_);
  or g_130723_(_054665_, _074060_, _074061_);
  xor g_130724_(_054665_, _074059_, _074063_);
  not g_130725_(_074063_, _074064_);
  or g_130726_(_054629_, _074063_, _074065_);
  xor g_130727_(_054629_, _074063_, _074066_);
  xor g_130728_(_054629_, _074064_, _074067_);
  or g_130729_(_054593_, _074067_, _074068_);
  xor g_130730_(_054593_, _074066_, _074069_);
  not g_130731_(_074069_, _074070_);
  or g_130732_(_054556_, _074069_, _074071_);
  xor g_130733_(_054556_, _074069_, _074072_);
  xor g_130734_(_054556_, _074070_, _074074_);
  or g_130735_(_054520_, _074074_, _074075_);
  xor g_130736_(_054520_, _074072_, _074076_);
  or g_130737_(_054484_, _074076_, _074077_);
  not g_130738_(_074077_, _074078_);
  and g_130739_(_054484_, _074076_, _074079_);
  xor g_130740_(_054484_, _074076_, _074080_);
  or g_130741_(_074078_, _074079_, _074081_);
  or g_130742_(_054447_, _074081_, _074082_);
  xor g_130743_(_054447_, _074080_, _074083_);
  or g_130744_(_054411_, _074083_, _074085_);
  xor g_130745_(_054411_, _074083_, _074086_);
  not g_130746_(_074086_, _074087_);
  or g_130747_(_054375_, _074087_, _074088_);
  xor g_130748_(_054375_, _074086_, _074089_);
  or g_130749_(_054337_, _074089_, _074090_);
  xor g_130750_(_054338_, _074089_, _074091_);
  or g_130751_(_054301_, _074091_, _074092_);
  xor g_130752_(_054301_, _074091_, _074093_);
  not g_130753_(_074093_, _074094_);
  or g_130754_(_054265_, _074094_, _074096_);
  xor g_130755_(_054265_, _074093_, _074097_);
  or g_130756_(_054227_, _074097_, _074098_);
  xor g_130757_(_054228_, _074097_, _074099_);
  or g_130758_(_054190_, _074099_, _074100_);
  xor g_130759_(_054191_, _074099_, _074101_);
  not g_130760_(_074101_, _074102_);
  or g_130761_(_054154_, _074101_, _074103_);
  xor g_130762_(_054154_, _074101_, _074104_);
  xor g_130763_(_054154_, _074102_, _074105_);
  or g_130764_(_054117_, _074105_, _074107_);
  xor g_130765_(_054117_, _074104_, _074108_);
  or g_130766_(_054080_, _074108_, _074109_);
  xor g_130767_(_054081_, _074108_, _074110_);
  or g_130768_(_054044_, _074110_, _074111_);
  not g_130769_(_074111_, _074112_);
  and g_130770_(_054044_, _074110_, _074113_);
  xor g_130771_(_054044_, _074110_, _074114_);
  or g_130772_(_074112_, _074113_, _074115_);
  or g_130773_(_054007_, _074115_, _074116_);
  xor g_130774_(_054007_, _074114_, _074118_);
  or g_130775_(_053970_, _074118_, _074119_);
  xor g_130776_(_053971_, _074118_, _074120_);
  or g_130777_(_053933_, _074120_, _074121_);
  not g_130778_(_074121_, _074122_);
  xor g_130779_(_053934_, _074120_, _074123_);
  not g_130780_(_074123_, _074124_);
  or g_130781_(_053896_, _074123_, _074125_);
  xor g_130782_(_053896_, _074123_, _074126_);
  xor g_130783_(_053896_, _074124_, _074127_);
  or g_130784_(_053860_, _074127_, _074129_);
  xor g_130785_(_053860_, _074126_, _074130_);
  not g_130786_(_074130_, _074131_);
  or g_130787_(_053824_, _074130_, _074132_);
  xor g_130788_(_053824_, _074130_, _074133_);
  xor g_130789_(_053824_, _074131_, _074134_);
  or g_130790_(_053787_, _074134_, _074135_);
  xor g_130791_(_053787_, _074133_, _074136_);
  or g_130792_(_053750_, _074136_, _074137_);
  xor g_130793_(_053751_, _074136_, _074138_);
  or g_130794_(_053713_, _074138_, _074140_);
  xor g_130795_(_053713_, _074138_, _074141_);
  xor g_130796_(_053714_, _074138_, _074142_);
  or g_130797_(_053676_, _074142_, _074143_);
  xor g_130798_(_053676_, _074141_, _074144_);
  or g_130799_(_053640_, _074144_, _074145_);
  not g_130800_(_074145_, _074146_);
  xor g_130801_(_053640_, _074144_, _074147_);
  not g_130802_(_074147_, _074148_);
  or g_130803_(_053604_, _074148_, _074149_);
  xor g_130804_(_053604_, _074147_, _074151_);
  or g_130805_(_053567_, _074151_, _074152_);
  xor g_130806_(_053567_, _074151_, _074153_);
  not g_130807_(_074153_, _074154_);
  or g_130808_(_053531_, _074154_, _074155_);
  xor g_130809_(_053531_, _074153_, _074156_);
  or g_130810_(_053494_, _074156_, _074157_);
  xor g_130811_(_053495_, _074156_, _074158_);
  or g_130812_(_053456_, _074158_, _074159_);
  xor g_130813_(_053457_, _074158_, _074160_);
  not g_130814_(_074160_, _074162_);
  or g_130815_(_053420_, _074160_, _074163_);
  xor g_130816_(_053420_, _074160_, _074164_);
  xor g_130817_(_053420_, _074162_, _074165_);
  or g_130818_(_053384_, _074165_, _074166_);
  xor g_130819_(_053384_, _074164_, _074167_);
  or g_130820_(_053346_, _074167_, _074168_);
  xor g_130821_(_053347_, _074167_, _074169_);
  or g_130822_(_053310_, _074169_, _074170_);
  xor g_130823_(_053310_, _074169_, _074171_);
  not g_130824_(_074171_, _074173_);
  or g_130825_(_053274_, _074173_, _074174_);
  not g_130826_(_074174_, _074175_);
  xor g_130827_(_053274_, _074171_, _074176_);
  or g_130828_(_053236_, _074176_, _074177_);
  xor g_130829_(_053237_, _074176_, _074178_);
  or g_130830_(_053199_, _074178_, _074179_);
  xor g_130831_(_053200_, _074178_, _074180_);
  or g_130832_(_053163_, _074180_, _074181_);
  not g_130833_(_074181_, _074182_);
  and g_130834_(_053163_, _074180_, _074184_);
  xor g_130835_(_053163_, _074180_, _074185_);
  or g_130836_(_074182_, _074184_, _074186_);
  or g_130837_(_053126_, _074186_, _074187_);
  not g_130838_(_074187_, _074188_);
  xor g_130839_(_053126_, _074185_, _074189_);
  not g_130840_(_074189_, _074190_);
  and g_130841_(_053090_, _074190_, _074191_);
  or g_130842_(_053089_, _074189_, _074192_);
  xor g_130843_(_053089_, _074189_, _074193_);
  not g_130844_(_074193_, _074195_);
  or g_130845_(_053053_, _074195_, _074196_);
  not g_130846_(_074196_, _074197_);
  xor g_130847_(_053053_, _074193_, _074198_);
  not g_130848_(_074198_, _074199_);
  or g_130849_(_053016_, _074198_, _074200_);
  xor g_130850_(_053016_, _074199_, _074201_);
  or g_130851_(_052980_, _074201_, _074202_);
  not g_130852_(_074202_, _074203_);
  xor g_130853_(_052980_, _074201_, _074204_);
  not g_130854_(_074204_, _074206_);
  or g_130855_(_052944_, _074206_, _074207_);
  xor g_130856_(_052944_, _074204_, _074208_);
  not g_130857_(_074208_, _074209_);
  or g_130858_(_052907_, _074208_, _074210_);
  xor g_130859_(_052907_, _074208_, _074211_);
  xor g_130860_(_052907_, _074209_, _074212_);
  or g_130861_(_052871_, _074212_, _074213_);
  xor g_130862_(_052871_, _074211_, _074214_);
  not g_130863_(_074214_, _074215_);
  or g_130864_(_052835_, _074214_, _074217_);
  xor g_130865_(_052835_, _074214_, _074218_);
  xor g_130866_(_052835_, _074215_, _074219_);
  or g_130867_(_052798_, _074219_, _074220_);
  xor g_130868_(_052798_, _074218_, _074221_);
  or g_130869_(_052762_, _074221_, _074222_);
  not g_130870_(_074222_, _074223_);
  xor g_130871_(_052762_, _074221_, _074224_);
  not g_130872_(_074224_, _074225_);
  or g_130873_(_052726_, _074225_, _074226_);
  xor g_130874_(_052726_, _074224_, _074228_);
  or g_130875_(_052688_, _074228_, _074229_);
  xor g_130876_(_052690_, _074228_, _074230_);
  not g_130877_(_074230_, _074231_);
  or g_130878_(_052652_, _074230_, _074232_);
  xor g_130879_(_052652_, _074230_, _074233_);
  xor g_130880_(_052652_, _074231_, _074234_);
  or g_130881_(_052616_, _074234_, _074235_);
  xor g_130882_(_052616_, _074233_, _074236_);
  not g_130883_(_074236_, _074237_);
  or g_130884_(_052580_, _074236_, _074239_);
  xor g_130885_(_052580_, _074236_, _074240_);
  xor g_130886_(_052580_, _074237_, _074241_);
  or g_130887_(_052543_, _074241_, _074242_);
  xor g_130888_(_052543_, _074240_, _074243_);
  or g_130889_(_052506_, _074243_, _074244_);
  not g_130890_(_074244_, _074245_);
  xor g_130891_(_052507_, _074243_, _074246_);
  not g_130892_(_074246_, _074247_);
  or g_130893_(_052470_, _074246_, _074248_);
  xor g_130894_(_052470_, _074246_, _074250_);
  xor g_130895_(_052470_, _074247_, _074251_);
  or g_130896_(_052433_, _074251_, _074252_);
  xor g_130897_(_052433_, _074250_, _074253_);
  or g_130898_(_052397_, _074253_, _074254_);
  xor g_130899_(_052397_, _074253_, _074255_);
  not g_130900_(_074255_, _074256_);
  or g_130901_(_052361_, _074256_, _074257_);
  xor g_130902_(_052361_, _074255_, _074258_);
  or g_130903_(_052323_, _074258_, _074259_);
  xor g_130904_(_052324_, _074258_, _074261_);
  or g_130905_(_052287_, _074261_, _074262_);
  not g_130906_(_074262_, _074263_);
  and g_130907_(_052287_, _074261_, _074264_);
  xor g_130908_(_052287_, _074261_, _074265_);
  or g_130909_(_074263_, _074264_, _074266_);
  or g_130910_(_052251_, _074266_, _074267_);
  xor g_130911_(_052251_, _074265_, _074268_);
  or g_130912_(_052213_, _074268_, _074269_);
  xor g_130913_(_052214_, _074268_, _074270_);
  not g_130914_(_074270_, _074272_);
  or g_130915_(_052177_, _074270_, _074273_);
  xor g_130916_(_052177_, _074270_, _074274_);
  xor g_130917_(_052177_, _074272_, _074275_);
  or g_130918_(_052141_, _074275_, _074276_);
  xor g_130919_(_052141_, _074274_, _074277_);
  or g_130920_(_052103_, _074277_, _074278_);
  xor g_130921_(_052104_, _074277_, _074279_);
  or g_130922_(_052066_, _074279_, _074280_);
  not g_130923_(_074280_, _074281_);
  xor g_130924_(_052067_, _074279_, _074283_);
  not g_130925_(_074283_, _074284_);
  or g_130926_(_052030_, _074283_, _074285_);
  xor g_130927_(_052030_, _074283_, _074286_);
  xor g_130928_(_052030_, _074284_, _074287_);
  or g_130929_(_051993_, _074287_, _074288_);
  xor g_130930_(_051993_, _074286_, _074289_);
  or g_130931_(_051956_, _074289_, _074290_);
  xor g_130932_(_051957_, _074289_, _074291_);
  or g_130933_(_051918_, _074291_, _074292_);
  xor g_130934_(_051920_, _074291_, _074294_);
  or g_130935_(_051881_, _074294_, _074295_);
  xor g_130936_(_051881_, _074294_, _074296_);
  xor g_130937_(_051882_, _074294_, _074297_);
  or g_130938_(_051845_, _074297_, _074298_);
  xor g_130939_(_051845_, _074296_, _074299_);
  not g_130940_(_074299_, _074300_);
  or g_130941_(_051808_, _074299_, _074301_);
  xor g_130942_(_051808_, _074299_, _074302_);
  xor g_130943_(_051808_, _074300_, _074303_);
  or g_130944_(_051772_, _074303_, _074305_);
  xor g_130945_(_051772_, _074302_, _074306_);
  or g_130946_(_051736_, _074306_, _074307_);
  not g_130947_(_074307_, _074308_);
  xor g_130948_(_051736_, _074306_, _074309_);
  not g_130949_(_074309_, _074310_);
  or g_130950_(_051700_, _074310_, _074311_);
  xor g_130951_(_051700_, _074309_, _074312_);
  or g_130952_(_051663_, _074312_, _074313_);
  xor g_130953_(_051663_, _074312_, _074314_);
  not g_130954_(_074314_, _074316_);
  or g_130955_(_051627_, _074316_, _074317_);
  not g_130956_(_074317_, _074318_);
  xor g_130957_(_051627_, _074314_, _074319_);
  or g_130958_(_051590_, _074319_, _074320_);
  xor g_130959_(_051591_, _074319_, _074321_);
  or g_130960_(_051552_, _074321_, _074322_);
  xor g_130961_(_051553_, _074321_, _074323_);
  or g_130962_(_051515_, _074323_, _074324_);
  xor g_130963_(_051516_, _074323_, _074325_);
  or g_130964_(_051478_, _074325_, _074327_);
  not g_130965_(_074327_, _074328_);
  and g_130966_(_051478_, _074325_, _074329_);
  xor g_130967_(_051478_, _074325_, _074330_);
  or g_130968_(_074328_, _074329_, _074331_);
  or g_130969_(_051442_, _074331_, _074332_);
  not g_130970_(_074332_, _074333_);
  xor g_130971_(_051442_, _074330_, _074334_);
  not g_130972_(_074334_, _074335_);
  or g_130973_(_051406_, _074334_, _074336_);
  xor g_130974_(_051406_, _074334_, _074338_);
  xor g_130975_(_051406_, _074335_, _074339_);
  or g_130976_(_051370_, _074339_, _074340_);
  xor g_130977_(_051370_, _074338_, _074341_);
  or g_130978_(_051332_, _074341_, _074342_);
  xor g_130979_(_051333_, _074341_, _074343_);
  or g_130980_(_051296_, _074343_, _074344_);
  xor g_130981_(_051296_, _074343_, _074345_);
  and g_130982_(_051260_, _074345_, _074346_);
  not g_130983_(_074346_, _074347_);
  xor g_130984_(_051258_, _074345_, _074349_);
  or g_130985_(_051222_, _074349_, _074350_);
  xor g_130986_(_051222_, _074349_, _074351_);
  not g_130987_(_074351_, _074352_);
  or g_130988_(_051186_, _074352_, _074353_);
  not g_130989_(_074353_, _074354_);
  xor g_130990_(_051186_, _074351_, _074355_);
  or g_130991_(_051148_, _074355_, _074356_);
  xor g_130992_(_051150_, _074355_, _074357_);
  or g_130993_(_051111_, _074357_, _074358_);
  xor g_130994_(_051112_, _074357_, _074360_);
  not g_130995_(_074360_, _074361_);
  or g_130996_(_051075_, _074360_, _074362_);
  xor g_130997_(_051075_, _074360_, _074363_);
  xor g_130998_(_051075_, _074361_, _074364_);
  or g_130999_(_051038_, _074364_, _074365_);
  xor g_131000_(_051038_, _074363_, _074366_);
  not g_131001_(_074366_, _074367_);
  or g_131002_(_051002_, _074366_, _074368_);
  xor g_131003_(_051002_, _074366_, _074369_);
  xor g_131004_(_051002_, _074367_, _074371_);
  and g_131005_(_050966_, _074369_, _074372_);
  or g_131006_(_050965_, _074371_, _074373_);
  xor g_131007_(_050966_, _074369_, _074374_);
  xor g_131008_(_050965_, _074369_, _074375_);
  and g_131009_(_050928_, _074374_, _074376_);
  or g_131010_(_050927_, _074375_, _074377_);
  xor g_131011_(_050928_, _074374_, _074378_);
  xor g_131012_(_050927_, _074374_, _074379_);
  or g_131013_(_050891_, _074379_, _074380_);
  xor g_131014_(_050891_, _074378_, _074382_);
  or g_131015_(_050854_, _074382_, _074383_);
  not g_131016_(_074383_, _074384_);
  xor g_131017_(_050855_, _074382_, _074385_);
  or g_131018_(_050816_, _074385_, _074386_);
  xor g_131019_(_050817_, _074385_, _074387_);
  or g_131020_(_050779_, _074387_, _074388_);
  xor g_131021_(_050780_, _074387_, _074389_);
  or g_131022_(_050741_, _074389_, _074390_);
  xor g_131023_(_050741_, _074389_, _074391_);
  xor g_131024_(_050743_, _074389_, _074393_);
  or g_131025_(_050705_, _074393_, _074394_);
  xor g_131026_(_050705_, _074391_, _074395_);
  or g_131027_(_050669_, _074395_, _074396_);
  xor g_131028_(_050669_, _074395_, _074397_);
  not g_131029_(_074397_, _074398_);
  and g_131030_(_050633_, _074397_, _074399_);
  or g_131031_(_050631_, _074398_, _074400_);
  xor g_131032_(_050631_, _074397_, _074401_);
  not g_131033_(_074401_, _074402_);
  or g_131034_(_050595_, _074401_, _074404_);
  not g_131035_(_074404_, _074405_);
  xor g_131036_(_050595_, _074402_, _074406_);
  or g_131037_(_050559_, _074406_, _074407_);
  xor g_131038_(_050559_, _074406_, _074408_);
  not g_131039_(_074408_, _074409_);
  or g_131040_(_050523_, _074409_, _074410_);
  not g_131041_(_074410_, _074411_);
  xor g_131042_(_050523_, _074408_, _074412_);
  or g_131043_(_050486_, _074412_, _074413_);
  not g_131044_(_074413_, _074415_);
  and g_131045_(_050486_, _074412_, _074416_);
  xor g_131046_(_050486_, _074412_, _074417_);
  or g_131047_(_074415_, _074416_, _074418_);
  or g_131048_(_050450_, _074418_, _074419_);
  xor g_131049_(_050450_, _074417_, _074420_);
  not g_131050_(_074420_, _074421_);
  or g_131051_(_050414_, _074420_, _074422_);
  xor g_131052_(_050414_, _074420_, _074423_);
  xor g_131053_(_050414_, _074421_, _074424_);
  or g_131054_(_050377_, _074424_, _074426_);
  xor g_131055_(_050377_, _074423_, _074427_);
  not g_131056_(_074427_, _074428_);
  or g_131057_(_050341_, _074427_, _074429_);
  xor g_131058_(_050341_, _074428_, _074430_);
  or g_131059_(_050304_, _074430_, _074431_);
  xor g_131060_(_050305_, _074430_, _074432_);
  not g_131061_(_074432_, _074433_);
  or g_131062_(_050267_, _074432_, _074434_);
  xor g_131063_(_050267_, _074432_, _074435_);
  xor g_131064_(_050267_, _074433_, _074437_);
  or g_131065_(_050231_, _074437_, _074438_);
  xor g_131066_(_050231_, _074435_, _074439_);
  not g_131067_(_074439_, _074440_);
  or g_131068_(_050195_, _074439_, _074441_);
  xor g_131069_(_050195_, _074439_, _074442_);
  xor g_131070_(_050195_, _074440_, _074443_);
  or g_131071_(_050158_, _074443_, _074444_);
  xor g_131072_(_050158_, _074442_, _074445_);
  or g_131073_(_050122_, _074445_, _074446_);
  xor g_131074_(_050122_, _074445_, _074448_);
  not g_131075_(_074448_, _074449_);
  or g_131076_(_050086_, _074449_, _074450_);
  not g_131077_(_074450_, _074451_);
  xor g_131078_(_050086_, _074448_, _074452_);
  not g_131079_(_074452_, _074453_);
  or g_131080_(_050050_, _074452_, _074454_);
  xor g_131081_(_050050_, _074452_, _074455_);
  xor g_131082_(_050050_, _074453_, _074456_);
  or g_131083_(_050013_, _074456_, _074457_);
  xor g_131084_(_050013_, _074455_, _074459_);
  not g_131085_(_074459_, _074460_);
  or g_131086_(_049977_, _074459_, _074461_);
  xor g_131087_(_049977_, _074460_, _074462_);
  not g_131088_(_074462_, _074463_);
  or g_131089_(_049941_, _074462_, _074464_);
  xor g_131090_(_049941_, _074463_, _074465_);
  or g_131091_(_049904_, _074465_, _074466_);
  not g_131092_(_074466_, _074467_);
  xor g_131093_(_049904_, _074465_, _074468_);
  not g_131094_(_074468_, _074470_);
  or g_131095_(_049868_, _074470_, _074471_);
  xor g_131096_(_049868_, _074468_, _074472_);
  not g_131097_(_074472_, _074473_);
  or g_131098_(_049832_, _074472_, _074474_);
  xor g_131099_(_049832_, _074472_, _074475_);
  xor g_131100_(_049832_, _074473_, _074476_);
  or g_131101_(_049795_, _074476_, _074477_);
  xor g_131102_(_049795_, _074475_, _074478_);
  or g_131103_(_049758_, _074478_, _074479_);
  not g_131104_(_074479_, _074481_);
  xor g_131105_(_049759_, _074478_, _074482_);
  not g_131106_(_074482_, _074483_);
  or g_131107_(_049722_, _074482_, _074484_);
  not g_131108_(_074484_, _074485_);
  xor g_131109_(_049722_, _074483_, _074486_);
  or g_131110_(_049684_, _074486_, _074487_);
  xor g_131111_(_049684_, _074486_, _074488_);
  xor g_131112_(_049685_, _074486_, _074489_);
  and g_131113_(_049648_, _074488_, _074490_);
  or g_131114_(_049647_, _074489_, _074492_);
  xor g_131115_(_049647_, _074488_, _074493_);
  not g_131116_(_074493_, _074494_);
  or g_131117_(_049611_, _074493_, _074495_);
  xor g_131118_(_049611_, _074494_, _074496_);
  or g_131119_(_049574_, _074496_, _074497_);
  xor g_131120_(_049574_, _074496_, _074498_);
  not g_131121_(_074498_, _074499_);
  or g_131122_(_049538_, _074499_, _074500_);
  xor g_131123_(_049538_, _074498_, _074501_);
  or g_131124_(_049501_, _074501_, _074503_);
  xor g_131125_(_049502_, _074501_, _074504_);
  not g_131126_(_074504_, _074505_);
  or g_131127_(_049464_, _074504_, _074506_);
  xor g_131128_(_049464_, _074504_, _074507_);
  xor g_131129_(_049464_, _074505_, _074508_);
  or g_131130_(_049428_, _074508_, _074509_);
  not g_131131_(_074509_, _074510_);
  xor g_131132_(_049428_, _074507_, _074511_);
  or g_131133_(_049391_, _074511_, _074512_);
  xor g_131134_(_049392_, _074511_, _074514_);
  or g_131135_(_098259_, _074514_, _074515_);
  xor g_131136_(_098259_, _074514_, _074516_);
  not g_131137_(_074516_, _074517_);
  and g_131138_(_098223_, _074516_, _074518_);
  or g_131139_(_098222_, _074517_, _074519_);
  xor g_131140_(_098222_, _074516_, _074520_);
  or g_131141_(_098185_, _074520_, _074521_);
  xor g_131142_(_098186_, _074520_, _074522_);
  or g_131143_(_098147_, _074522_, _074523_);
  xor g_131144_(_098148_, _074522_, _074525_);
  not g_131145_(_074525_, _074526_);
  or g_131146_(_098111_, _074525_, _074527_);
  xor g_131147_(_098111_, _074525_, _074528_);
  xor g_131148_(_098111_, _074526_, _074529_);
  or g_131149_(_098075_, _074529_, _074530_);
  xor g_131150_(_098075_, _074528_, _074531_);
  or g_131151_(_098037_, _074531_, _074532_);
  xor g_131152_(_098038_, _074531_, _074533_);
  or g_131153_(_098000_, _074533_, _074534_);
  xor g_131154_(_098001_, _074533_, _074536_);
  not g_131155_(_074536_, _074537_);
  or g_131156_(_097963_, _074536_, _074538_);
  xor g_131157_(_097963_, _074536_, _074539_);
  xor g_131158_(_097963_, _074537_, _074540_);
  or g_131159_(_097930_, _074540_, _074541_);
  xor g_131160_(_097930_, _074539_, _074542_);
  or g_131161_(_097896_, _074542_, _074543_);
  xor g_131162_(_097897_, _074542_, _074544_);
  not g_131163_(_074544_, _074545_);
  or g_131164_(_097863_, _074544_, _074547_);
  xor g_131165_(_097863_, _074544_, _074548_);
  xor g_131166_(_097863_, _074545_, _074549_);
  or g_131167_(_097830_, _074549_, _074550_);
  xor g_131168_(_097830_, _074548_, _074551_);
  not g_131169_(_074551_, _074552_);
  or g_131170_(_097797_, _074551_, _074553_);
  xor g_131171_(_097797_, _074551_, _074554_);
  xor g_131172_(_097797_, _074552_, _074555_);
  or g_131173_(_097764_, _074555_, _074556_);
  xor g_131174_(_097764_, _074554_, _074558_);
  or g_131175_(_097730_, _074558_, _074559_);
  xor g_131176_(_097731_, _074558_, _074560_);
  or g_131177_(_097696_, _074560_, _074561_);
  xor g_131178_(_097697_, _074560_, _074562_);
  or g_131179_(_097662_, _074562_, _074563_);
  xor g_131180_(_097663_, _074562_, _074564_);
  not g_131181_(_074564_, _074565_);
  or g_131182_(_097629_, _074564_, _074566_);
  xor g_131183_(_097629_, _074564_, _074567_);
  xor g_131184_(_097629_, _074565_, _074569_);
  or g_131185_(_097596_, _074569_, _074570_);
  xor g_131186_(_097596_, _074567_, _074571_);
  not g_131187_(_074571_, _074572_);
  or g_131188_(_097563_, _074571_, _074573_);
  xor g_131189_(_097563_, _074571_, _074574_);
  xor g_131190_(_097563_, _074572_, _074575_);
  or g_131191_(_097530_, _074575_, _074576_);
  xor g_131192_(_097530_, _074574_, _074577_);
  or g_131193_(_097497_, _074577_, _074578_);
  not g_131194_(_074578_, _074580_);
  xor g_131195_(_097497_, _074577_, _074581_);
  not g_131196_(_074581_, _074582_);
  or g_131197_(_097464_, _074582_, _074583_);
  not g_131198_(_074583_, _074584_);
  xor g_131199_(_097464_, _074581_, _074585_);
  or g_131200_(_097430_, _074585_, _074586_);
  not g_131201_(_074586_, _074587_);
  xor g_131202_(_097431_, _074585_, _074588_);
  or g_131203_(_097396_, _074588_, _074589_);
  xor g_131204_(_097397_, _074588_, _074591_);
  not g_131205_(_074591_, _074592_);
  or g_131206_(_097363_, _074591_, _074593_);
  xor g_131207_(_097363_, _074591_, _074594_);
  xor g_131208_(_097363_, _074592_, _074595_);
  or g_131209_(_097330_, _074595_, _074596_);
  xor g_131210_(_097330_, _074594_, _074597_);
  or g_131211_(_097296_, _074597_, _074598_);
  xor g_131212_(_097297_, _074597_, _074599_);
  or g_131213_(_097263_, _074599_, _074600_);
  xor g_131214_(_097263_, _074599_, _074602_);
  not g_131215_(_074602_, _074603_);
  or g_131216_(_097230_, _074603_, _074604_);
  xor g_131217_(_097230_, _074602_, _074605_);
  or g_131218_(_097196_, _074605_, _074606_);
  xor g_131219_(_097197_, _074605_, _074607_);
  or g_131220_(_097163_, _074607_, _074608_);
  not g_131221_(_074608_, _074609_);
  and g_131222_(_097163_, _074607_, _074610_);
  xor g_131223_(_097163_, _074607_, _074611_);
  or g_131224_(_074609_, _074610_, _074613_);
  or g_131225_(_097130_, _074613_, _074614_);
  xor g_131226_(_097130_, _074611_, _074615_);
  or g_131227_(_097096_, _074615_, _074616_);
  xor g_131228_(_097097_, _074615_, _074617_);
  not g_131229_(_074617_, _074618_);
  or g_131230_(_097063_, _074617_, _074619_);
  xor g_131231_(_097063_, _074617_, _074620_);
  xor g_131232_(_097063_, _074618_, _074621_);
  or g_131233_(_097030_, _074621_, _074622_);
  xor g_131234_(_097030_, _074620_, _074624_);
  or g_131235_(_096997_, _074624_, _074625_);
  xor g_131236_(_096997_, _074624_, _074626_);
  not g_131237_(_074626_, _074627_);
  or g_131238_(_096964_, _074627_, _074628_);
  xor g_131239_(_096964_, _074626_, _074629_);
  not g_131240_(_074629_, _074630_);
  or g_131241_(_096931_, _074629_, _074631_);
  xor g_131242_(_096931_, _074629_, _074632_);
  xor g_131243_(_096931_, _074630_, _074633_);
  or g_131244_(_096898_, _074633_, _074635_);
  xor g_131245_(_096898_, _074632_, _074636_);
  or g_131246_(_096864_, _074636_, _074637_);
  xor g_131247_(_096865_, _074636_, _074638_);
  or g_131248_(_096831_, _074638_, _074639_);
  xor g_131249_(_096831_, _074638_, _074640_);
  not g_131250_(_074640_, _074641_);
  or g_131251_(_096798_, _074641_, _074642_);
  not g_131252_(_074642_, _074643_);
  xor g_131253_(_096798_, _074640_, _074644_);
  or g_131254_(_096764_, _074644_, _074646_);
  not g_131255_(_074646_, _074647_);
  xor g_131256_(_096765_, _074644_, _074648_);
  not g_131257_(_074648_, _074649_);
  or g_131258_(_096731_, _074648_, _074650_);
  xor g_131259_(_096731_, _074648_, _074651_);
  xor g_131260_(_096731_, _074649_, _074652_);
  or g_131261_(_096698_, _074652_, _074653_);
  xor g_131262_(_096698_, _074651_, _074654_);
  or g_131263_(_096664_, _074654_, _074655_);
  not g_131264_(_074655_, _074657_);
  xor g_131265_(_096665_, _074654_, _074658_);
  not g_131266_(_074658_, _074659_);
  or g_131267_(_096631_, _074658_, _074660_);
  xor g_131268_(_096631_, _074658_, _074661_);
  xor g_131269_(_096631_, _074659_, _074662_);
  or g_131270_(_096598_, _074662_, _074663_);
  xor g_131271_(_096598_, _074661_, _074664_);
  or g_131272_(_096564_, _074664_, _074665_);
  xor g_131273_(_096565_, _074664_, _074666_);
  or g_131274_(_096531_, _074666_, _074668_);
  not g_131275_(_074668_, _074669_);
  and g_131276_(_096531_, _074666_, _074670_);
  xor g_131277_(_096531_, _074666_, _074671_);
  or g_131278_(_074669_, _074670_, _074672_);
  or g_131279_(_096498_, _074672_, _074673_);
  xor g_131280_(_096498_, _074671_, _074674_);
  not g_131281_(_074674_, _074675_);
  or g_131282_(_096465_, _074674_, _074676_);
  xor g_131283_(_096465_, _074674_, _074677_);
  xor g_131284_(_096465_, _074675_, _074679_);
  or g_131285_(_096432_, _074679_, _074680_);
  xor g_131286_(_096432_, _074677_, _074681_);
  or g_131287_(_096398_, _074681_, _074682_);
  not g_131288_(_074682_, _074683_);
  xor g_131289_(_096399_, _074681_, _074684_);
  or g_131290_(_096364_, _074684_, _074685_);
  xor g_131291_(_096365_, _074684_, _074686_);
  or g_131292_(_096330_, _074686_, _074687_);
  xor g_131293_(_096331_, _074686_, _074688_);
  or g_131294_(_096296_, _074688_, _074690_);
  xor g_131295_(_096297_, _074688_, _074691_);
  not g_131296_(_074691_, _074692_);
  or g_131297_(_096263_, _074691_, _074693_);
  xor g_131298_(_096263_, _074691_, _074694_);
  xor g_131299_(_096263_, _074692_, _074695_);
  or g_131300_(_096230_, _074695_, _074696_);
  xor g_131301_(_096230_, _074694_, _074697_);
  or g_131302_(_096196_, _074697_, _074698_);
  xor g_131303_(_096197_, _074697_, _074699_);
  not g_131304_(_074699_, _074701_);
  or g_131305_(_096163_, _074699_, _074702_);
  xor g_131306_(_096163_, _074699_, _074703_);
  xor g_131307_(_096163_, _074701_, _074704_);
  or g_131308_(_096130_, _074704_, _074705_);
  xor g_131309_(_096130_, _074703_, _074706_);
  or g_131310_(_096096_, _074706_, _074707_);
  xor g_131311_(_096097_, _074706_, _074708_);
  or g_131312_(_096063_, _074708_, _074709_);
  not g_131313_(_074709_, _074710_);
  and g_131314_(_096063_, _074708_, _074712_);
  or g_131315_(_074710_, _074712_, _074713_);
  not g_131316_(_074713_, _074714_);
  or g_131317_(_096030_, _074713_, _074715_);
  or g_131318_(_096030_, _074712_, _074716_);
  xor g_131319_(_096030_, _074713_, _074717_);
  xor g_131320_(_096030_, _074714_, _074718_);
  or g_131321_(_095997_, _074718_, _074719_);
  xor g_131322_(_095997_, _074717_, _074720_);
  or g_131323_(_095964_, _074720_, _074721_);
  xor g_131324_(_095964_, _074720_, _074723_);
  not g_131325_(_074723_, _074724_);
  or g_131326_(_095931_, _074724_, _074725_);
  not g_131327_(_074725_, _074726_);
  xor g_131328_(_095931_, _074723_, _074727_);
  not g_131329_(_074727_, _074728_);
  or g_131330_(_095898_, _074727_, _074729_);
  xor g_131331_(_095898_, _074727_, _074730_);
  xor g_131332_(_095898_, _074728_, _074731_);
  or g_131333_(_095865_, _074731_, _074732_);
  xor g_131334_(_095865_, _074730_, _074734_);
  or g_131335_(_095831_, _074734_, _074735_);
  xor g_131336_(_095832_, _074734_, _074736_);
  not g_131337_(_074736_, _074737_);
  or g_131338_(_095798_, _074736_, _074738_);
  xor g_131339_(_095798_, _074736_, _074739_);
  xor g_131340_(_095798_, _074737_, _074740_);
  or g_131341_(_095765_, _074740_, _074741_);
  xor g_131342_(_095765_, _074739_, _074742_);
  or g_131343_(_095732_, _074742_, _074743_);
  not g_131344_(_074743_, _074745_);
  and g_131345_(_095732_, _074742_, _074746_);
  xor g_131346_(_095732_, _074742_, _074747_);
  or g_131347_(_074745_, _074746_, _074748_);
  or g_131348_(_095699_, _074748_, _074749_);
  xor g_131349_(_095699_, _074747_, _074750_);
  or g_131350_(_095665_, _074750_, _074751_);
  xor g_131351_(_095666_, _074750_, _074752_);
  not g_131352_(_074752_, _074753_);
  or g_131353_(_095632_, _074752_, _074754_);
  xor g_131354_(_095632_, _074752_, _074756_);
  xor g_131355_(_095632_, _074753_, _074757_);
  or g_131356_(_095599_, _074757_, _074758_);
  not g_131357_(_074758_, _074759_);
  xor g_131358_(_095599_, _074756_, _074760_);
  or g_131359_(_095565_, _074760_, _074761_);
  xor g_131360_(_095566_, _074760_, _074762_);
  or g_131361_(_095531_, _074762_, _074763_);
  xor g_131362_(_095532_, _074762_, _074764_);
  not g_131363_(_074764_, _074765_);
  or g_131364_(_095498_, _074764_, _074767_);
  xor g_131365_(_095498_, _074764_, _074768_);
  xor g_131366_(_095498_, _074765_, _074769_);
  or g_131367_(_095465_, _074769_, _074770_);
  xor g_131368_(_095465_, _074768_, _074771_);
  or g_131369_(_095432_, _074771_, _074772_);
  not g_131370_(_074772_, _074773_);
  and g_131371_(_095432_, _074771_, _074774_);
  xor g_131372_(_095432_, _074771_, _074775_);
  or g_131373_(_074773_, _074774_, _074776_);
  or g_131374_(_095399_, _074776_, _074778_);
  xor g_131375_(_095399_, _074775_, _074779_);
  or g_131376_(_095365_, _074779_, _074780_);
  xor g_131377_(_095366_, _074779_, _074781_);
  or g_131378_(_095331_, _074781_, _074782_);
  xor g_131379_(_095332_, _074781_, _074783_);
  or g_131380_(_095297_, _074783_, _074784_);
  xor g_131381_(_095298_, _074783_, _074785_);
  not g_131382_(_074785_, _074786_);
  or g_131383_(_095264_, _074785_, _074787_);
  xor g_131384_(_095264_, _074785_, _074789_);
  xor g_131385_(_095264_, _074786_, _074790_);
  or g_131386_(_095231_, _074790_, _074791_);
  xor g_131387_(_095231_, _074789_, _074792_);
  or g_131388_(_095197_, _074792_, _074793_);
  xor g_131389_(_095198_, _074792_, _074794_);
  or g_131390_(_095163_, _074794_, _074795_);
  not g_131391_(_074795_, _074796_);
  xor g_131392_(_095164_, _074794_, _074797_);
  or g_131393_(_095129_, _074797_, _074798_);
  xor g_131394_(_095130_, _074797_, _074800_);
  not g_131395_(_074800_, _074801_);
  or g_131396_(_095096_, _074800_, _074802_);
  xor g_131397_(_095096_, _074800_, _074803_);
  xor g_131398_(_095096_, _074801_, _074804_);
  or g_131399_(_095063_, _074804_, _074805_);
  not g_131400_(_074805_, _074806_);
  xor g_131401_(_095063_, _074803_, _074807_);
  or g_131402_(_095030_, _074807_, _074808_);
  xor g_131403_(_095030_, _074807_, _074809_);
  not g_131404_(_074809_, _074811_);
  or g_131405_(_094997_, _074811_, _074812_);
  xor g_131406_(_094997_, _074809_, _074813_);
  or g_131407_(_094963_, _074813_, _074814_);
  xor g_131408_(_094964_, _074813_, _074815_);
  or g_131409_(_094929_, _074815_, _074816_);
  xor g_131410_(_094930_, _074815_, _074817_);
  not g_131411_(_074817_, _074818_);
  or g_131412_(_094896_, _074817_, _074819_);
  xor g_131413_(_094896_, _074817_, _074820_);
  xor g_131414_(_094896_, _074818_, _074822_);
  or g_131415_(_094863_, _074822_, _074823_);
  xor g_131416_(_094863_, _074820_, _074824_);
  or g_131417_(_094829_, _074824_, _074825_);
  xor g_131418_(_094830_, _074824_, _074826_);
  or g_131419_(_094796_, _074826_, _074827_);
  not g_131420_(_074827_, _074828_);
  and g_131421_(_094796_, _074826_, _074829_);
  xor g_131422_(_094796_, _074826_, _074830_);
  or g_131423_(_074828_, _074829_, _074831_);
  or g_131424_(_094763_, _074831_, _074833_);
  xor g_131425_(_094763_, _074830_, _074834_);
  or g_131426_(_094729_, _074834_, _074835_);
  xor g_131427_(_094730_, _074834_, _074836_);
  or g_131428_(_094695_, _074836_, _074837_);
  xor g_131429_(_094696_, _074836_, _074838_);
  or g_131430_(_094662_, _074838_, _074839_);
  xor g_131431_(_094662_, _074838_, _074840_);
  not g_131432_(_074840_, _074841_);
  and g_131433_(_094629_, _074840_, _074842_);
  or g_131434_(_094628_, _074841_, _074844_);
  xor g_131435_(_094628_, _074840_, _074845_);
  or g_131436_(_094595_, _074845_, _074846_);
  xor g_131437_(_094594_, _074845_, _074847_);
  not g_131438_(_074847_, _074848_);
  or g_131439_(_094559_, _074847_, _074849_);
  xor g_131440_(_094559_, _074847_, _074850_);
  xor g_131441_(_094559_, _074848_, _074851_);
  or g_131442_(_094526_, _074851_, _074852_);
  xor g_131443_(_094526_, _074850_, _074853_);
  or g_131444_(_094493_, _074853_, _074855_);
  not g_131445_(_074855_, _074856_);
  and g_131446_(_094493_, _074853_, _074857_);
  xor g_131447_(_094493_, _074853_, _074858_);
  or g_131448_(_074856_, _074857_, _074859_);
  or g_131449_(_094460_, _074859_, _074860_);
  xor g_131450_(_094460_, _074858_, _074861_);
  not g_131451_(_074861_, _074862_);
  or g_131452_(_094427_, _074861_, _074863_);
  not g_131453_(_074863_, _074864_);
  xor g_131454_(_094427_, _074862_, _074866_);
  or g_131455_(_094394_, _074866_, _074867_);
  not g_131456_(_074867_, _074868_);
  xor g_131457_(_094394_, _074866_, _074869_);
  not g_131458_(_074869_, _074870_);
  or g_131459_(_094361_, _074870_, _074871_);
  xor g_131460_(_094361_, _074869_, _074872_);
  or g_131461_(_094327_, _074872_, _074873_);
  xor g_131462_(_094328_, _074872_, _074874_);
  or g_131463_(_094293_, _074874_, _074875_);
  xor g_131464_(_094294_, _074874_, _074877_);
  or g_131465_(_094259_, _074877_, _074878_);
  xor g_131466_(_094260_, _074877_, _074879_);
  or g_131467_(_094225_, _074879_, _074880_);
  xor g_131468_(_094226_, _074879_, _074881_);
  or g_131469_(_094191_, _074881_, _074882_);
  xor g_131470_(_094191_, _074881_, _074883_);
  xor g_131471_(_094192_, _074881_, _074884_);
  or g_131472_(_094158_, _074884_, _074885_);
  xor g_131473_(_094158_, _074883_, _074886_);
  not g_131474_(_074886_, _074888_);
  or g_131475_(_094125_, _074886_, _074889_);
  xor g_131476_(_094125_, _074886_, _074890_);
  xor g_131477_(_094125_, _074888_, _074891_);
  and g_131478_(_094092_, _074890_, _074892_);
  or g_131479_(_094091_, _074891_, _074893_);
  xor g_131480_(_094092_, _074890_, _074894_);
  not g_131481_(_074894_, _074895_);
  and g_131482_(_094058_, _074894_, _074896_);
  or g_131483_(_094057_, _074895_, _074897_);
  xor g_131484_(_094057_, _074894_, _074899_);
  or g_131485_(_094024_, _074899_, _074900_);
  xor g_131486_(_094024_, _074899_, _074901_);
  and g_131487_(_093991_, _074901_, _074902_);
  not g_131488_(_074902_, _074903_);
  xor g_131489_(_093990_, _074901_, _074904_);
  not g_131490_(_074904_, _074905_);
  and g_131491_(_093957_, _074905_, _074906_);
  or g_131492_(_093956_, _074904_, _074907_);
  xor g_131493_(_093956_, _074904_, _074908_);
  xor g_131494_(_093957_, _074904_, _074910_);
  and g_131495_(_093923_, _074908_, _074911_);
  or g_131496_(_093922_, _074910_, _074912_);
  xor g_131497_(_093922_, _074908_, _074913_);
  not g_131498_(_074913_, _074914_);
  or g_131499_(_093889_, _074913_, _074915_);
  xor g_131500_(_093889_, _074913_, _074916_);
  xor g_131501_(_093889_, _074914_, _074917_);
  or g_131502_(_093856_, _074917_, _074918_);
  xor g_131503_(_093856_, _074916_, _074919_);
  or g_131504_(_093823_, _074919_, _074921_);
  xor g_131505_(_093823_, _074919_, _074922_);
  not g_131506_(_074922_, _074923_);
  or g_131507_(_093790_, _074923_, _074924_);
  xor g_131508_(_093790_, _074922_, _074925_);
  not g_131509_(_074925_, _074926_);
  or g_131510_(_093757_, _074925_, _074927_);
  xor g_131511_(_093757_, _074925_, _074928_);
  xor g_131512_(_093757_, _074926_, _074929_);
  or g_131513_(_093724_, _074929_, _074930_);
  xor g_131514_(_093724_, _074928_, _074932_);
  not g_131515_(_074932_, _074933_);
  or g_131516_(_093691_, _074932_, _074934_);
  xor g_131517_(_093691_, _074933_, _074935_);
  or g_131518_(_093657_, _074935_, _074936_);
  xor g_131519_(_093658_, _074935_, _074937_);
  or g_131520_(_093624_, _074937_, _074938_);
  xor g_131521_(_093624_, _074937_, _074939_);
  not g_131522_(_074939_, _074940_);
  or g_131523_(_093591_, _074940_, _074941_);
  xor g_131524_(_093591_, _074939_, _074943_);
  not g_131525_(_074943_, _074944_);
  or g_131526_(_093558_, _074943_, _074945_);
  xor g_131527_(_093558_, _074943_, _074946_);
  xor g_131528_(_093558_, _074944_, _074947_);
  or g_131529_(_093525_, _074947_, _074948_);
  xor g_131530_(_093525_, _074946_, _074949_);
  or g_131531_(_093491_, _074949_, _074950_);
  xor g_131532_(_093492_, _074949_, _074951_);
  or g_131533_(_093458_, _074951_, _074952_);
  not g_131534_(_074952_, _074954_);
  xor g_131535_(_093458_, _074951_, _074955_);
  not g_131536_(_074955_, _074956_);
  or g_131537_(_093425_, _074956_, _074957_);
  xor g_131538_(_093425_, _074955_, _074958_);
  or g_131539_(_093391_, _074958_, _074959_);
  xor g_131540_(_093392_, _074958_, _074960_);
  or g_131541_(_093357_, _074960_, _074961_);
  xor g_131542_(_093358_, _074960_, _074962_);
  or g_131543_(_093323_, _074962_, _074963_);
  not g_131544_(_074963_, _074965_);
  xor g_131545_(_093324_, _074962_, _074966_);
  or g_131546_(_093289_, _074966_, _074967_);
  xor g_131547_(_093290_, _074966_, _074968_);
  not g_131548_(_074968_, _074969_);
  or g_131549_(_093256_, _074968_, _074970_);
  xor g_131550_(_093256_, _074968_, _074971_);
  xor g_131551_(_093256_, _074969_, _074972_);
  or g_131552_(_092942_, _074972_, _074973_);
  not g_131553_(_074973_, _074974_);
  xor g_131554_(_092942_, _074971_, _074976_);
  not g_131555_(_074976_, _074977_);
  or g_131556_(_092579_, _074976_, _074978_);
  xor g_131557_(_092579_, _074976_, _074979_);
  xor g_131558_(_092579_, _074977_, _074980_);
  or g_131559_(_092216_, _074980_, _074981_);
  not g_131560_(_074981_, _074982_);
  xor g_131561_(_092216_, _074979_, _074983_);
  or g_131562_(_091854_, _074983_, _074984_);
  not g_131563_(_074984_, _074985_);
  and g_131564_(_091854_, _074983_, _074987_);
  xor g_131565_(_091854_, _074983_, _074988_);
  or g_131566_(_074985_, _074987_, _074989_);
  or g_131567_(_091491_, _074989_, _074990_);
  xor g_131568_(_091491_, _074988_, _074991_);
  not g_131569_(_074991_, _074992_);
  or g_131570_(_091128_, _074991_, _074993_);
  xor g_131571_(_091128_, _074991_, _074994_);
  xor g_131572_(_091128_, _074992_, _074995_);
  or g_131573_(_090765_, _074995_, _074996_);
  not g_131574_(_074996_, _074998_);
  xor g_131575_(_090765_, _074994_, _074999_);
  or g_131576_(_090391_, _074999_, _075000_);
  xor g_131577_(_090402_, _074999_, _075001_);
  not g_131578_(_075001_, _075002_);
  or g_131579_(_090028_, _075001_, _075003_);
  xor g_131580_(_090028_, _075001_, _075004_);
  xor g_131581_(_090028_, _075002_, _075005_);
  or g_131582_(_089665_, _075005_, _075006_);
  xor g_131583_(_089665_, _075004_, _075007_);
  or g_131584_(_089292_, _075007_, _075009_);
  not g_131585_(_075009_, _075010_);
  xor g_131586_(_089303_, _075007_, _075011_);
  not g_131587_(_075011_, _075012_);
  or g_131588_(_088929_, _075011_, _075013_);
  xor g_131589_(_088929_, _075012_, _075014_);
  or g_131590_(_088555_, _075014_, _075015_);
  xor g_131591_(_088566_, _075014_, _075016_);
  or g_131592_(_088192_, _075016_, _075017_);
  not g_131593_(_075017_, _075018_);
  xor g_131594_(_088192_, _075016_, _075020_);
  and g_131595_(_087829_, _075020_, _075021_);
  not g_131596_(_075021_, _075022_);
  xor g_131597_(_087818_, _075020_, _075023_);
  or g_131598_(_087444_, _075023_, _075024_);
  xor g_131599_(_087455_, _075023_, _075025_);
  or g_131600_(_087070_, _075025_, _075026_);
  xor g_131601_(_087081_, _075025_, _075027_);
  not g_131602_(_075027_, _075028_);
  or g_131603_(_086708_, _075027_, _075029_);
  xor g_131604_(_086708_, _075027_, _075031_);
  xor g_131605_(_086708_, _075028_, _075032_);
  or g_131606_(_086345_, _075032_, _075033_);
  xor g_131607_(_086345_, _075031_, _075034_);
  or g_131608_(_085971_, _075034_, _075035_);
  xor g_131609_(_085982_, _075034_, _075036_);
  not g_131610_(_075036_, _075037_);
  or g_131611_(_085608_, _075036_, _075038_);
  xor g_131612_(_085608_, _075036_, _075039_);
  xor g_131613_(_085608_, _075037_, _075040_);
  or g_131614_(_085245_, _075040_, _075042_);
  not g_131615_(_075042_, _075043_);
  xor g_131616_(_085245_, _075039_, _075044_);
  not g_131617_(_075044_, _075045_);
  or g_131618_(_084882_, _075044_, _075046_);
  xor g_131619_(_084882_, _075044_, _075047_);
  xor g_131620_(_084882_, _075045_, _075048_);
  or g_131621_(_084519_, _075048_, _075049_);
  xor g_131622_(_084519_, _075047_, _075050_);
  not g_131623_(_075050_, _075051_);
  or g_131624_(_084156_, _075050_, _075053_);
  xor g_131625_(_084156_, _075050_, _075054_);
  xor g_131626_(_084156_, _075051_, _075055_);
  or g_131627_(_083794_, _075055_, _075056_);
  xor g_131628_(_083794_, _075054_, _075057_);
  or g_131629_(_083420_, _075057_, _075058_);
  xor g_131630_(_083431_, _075057_, _075059_);
  or g_131631_(_083057_, _075059_, _075060_);
  not g_131632_(_075060_, _075061_);
  xor g_131633_(_083057_, _075059_, _075062_);
  not g_131634_(_075062_, _075064_);
  or g_131635_(_082694_, _075064_, _075065_);
  xor g_131636_(_082694_, _075062_, _075066_);
  or g_131637_(_082320_, _075066_, _075067_);
  xor g_131638_(_082331_, _075066_, _075068_);
  not g_131639_(_075068_, _075069_);
  or g_131640_(_081957_, _075068_, _075070_);
  xor g_131641_(_081957_, _075068_, _075071_);
  xor g_131642_(_081957_, _075069_, _075072_);
  or g_131643_(_081594_, _075072_, _075073_);
  xor g_131644_(_081594_, _075071_, _075075_);
  or g_131645_(_081220_, _075075_, _075076_);
  xor g_131646_(_081231_, _075075_, _075077_);
  or g_131647_(_080847_, _075077_, _075078_);
  xor g_131648_(_080858_, _075077_, _075079_);
  not g_131649_(_075079_, _075080_);
  or g_131650_(_080484_, _075079_, _075081_);
  xor g_131651_(_080484_, _075079_, _075082_);
  xor g_131652_(_080484_, _075080_, _075083_);
  or g_131653_(_080121_, _075083_, _075084_);
  xor g_131654_(_080121_, _075082_, _075086_);
  or g_131655_(_079758_, _075086_, _075087_);
  not g_131656_(_075087_, _075088_);
  and g_131657_(_079758_, _075086_, _075089_);
  xor g_131658_(_079758_, _075086_, _075090_);
  or g_131659_(_075088_, _075089_, _075091_);
  or g_131660_(_079395_, _075091_, _075092_);
  xor g_131661_(_079395_, _075090_, _075093_);
  or g_131662_(_079021_, _075093_, _075094_);
  xor g_131663_(_079032_, _075093_, _075095_);
  or g_131664_(_078647_, _075095_, _075097_);
  not g_131665_(_075097_, _075098_);
  xor g_131666_(_078658_, _075095_, _075099_);
  or g_131667_(_078284_, _075099_, _075100_);
  xor g_131668_(_078284_, _075099_, _075101_);
  not g_131669_(_075101_, _075102_);
  or g_131670_(_077922_, _075102_, _075103_);
  xor g_131671_(_077922_, _075101_, _075104_);
  or g_131672_(_077548_, _075104_, _075105_);
  not g_131673_(_075105_, _075106_);
  xor g_131674_(_077559_, _075104_, _075108_);
  or g_131675_(_077174_, _075108_, _075109_);
  xor g_131676_(_077185_, _075108_, _075110_);
  not g_131677_(_075110_, _075111_);
  or g_131678_(_076811_, _075110_, _075112_);
  xor g_131679_(_076811_, _075110_, _075113_);
  xor g_131680_(_076811_, _075111_, _075114_);
  or g_131681_(_076448_, _075114_, _075115_);
  not g_131682_(_075115_, _075116_);
  xor g_131683_(_076448_, _075113_, _075117_);
  not g_131684_(_075117_, _075119_);
  and g_131685_(_076085_, _075119_, _075120_);
  xor g_131686_(_076074_, _075117_, _075121_);
  xor g_131687_(_076085_, _075117_, _075122_);
  or g_131688_(_075711_, _075122_, _075123_);
  xor g_131689_(_075711_, _075121_, _075124_);
  not g_131690_(_075124_, _075125_);
  or g_131691_(_075349_, _075124_, _075126_);
  xor g_131692_(_075349_, _075124_, _075127_);
  xor g_131693_(_075349_, _075125_, _075128_);
  or g_131694_(_074986_, _075128_, _075130_);
  not g_131695_(_075130_, _075131_);
  xor g_131696_(_074986_, _075127_, _075132_);
  or g_131697_(_074623_, _075132_, _075133_);
  not g_131698_(_075133_, _075134_);
  and g_131699_(_074623_, _075132_, _075135_);
  xor g_131700_(_074623_, _075132_, _075136_);
  or g_131701_(_075134_, _075135_, _075137_);
  or g_131702_(_074260_, _075137_, _075138_);
  xor g_131703_(_074260_, _075136_, _075139_);
  or g_131704_(_073886_, _075139_, _075141_);
  xor g_131705_(_073897_, _075139_, _075142_);
  not g_131706_(_075142_, _075143_);
  or g_131707_(_073523_, _075142_, _075144_);
  not g_131708_(_075144_, _075145_);
  xor g_131709_(_073523_, _075143_, _075146_);
  or g_131710_(_073160_, _075146_, _075147_);
  not g_131711_(_075147_, _075148_);
  xor g_131712_(_073160_, _075146_, _075149_);
  not g_131713_(_075149_, _075150_);
  or g_131714_(_072797_, _075150_, _075152_);
  xor g_131715_(_072797_, _075149_, _075153_);
  or g_131716_(_072423_, _075153_, _075154_);
  xor g_131717_(_072423_, _075153_, _075155_);
  xor g_131718_(_072434_, _075153_, _075156_);
  and g_131719_(_072060_, _075155_, _075157_);
  or g_131720_(_072049_, _075156_, _075158_);
  xor g_131721_(_072049_, _075155_, _075159_);
  or g_131722_(_071675_, _075159_, _075160_);
  xor g_131723_(_071686_, _075159_, _075161_);
  or g_131724_(_071312_, _075161_, _075163_);
  xor g_131725_(_071312_, _075161_, _075164_);
  not g_131726_(_075164_, _075165_);
  or g_131727_(_070949_, _075165_, _075166_);
  xor g_131728_(_070949_, _075164_, _075167_);
  not g_131729_(_075167_, _075168_);
  or g_131730_(_070586_, _075167_, _075169_);
  xor g_131731_(_070586_, _075167_, _075170_);
  xor g_131732_(_070586_, _075168_, _075171_);
  or g_131733_(_070223_, _075171_, _075172_);
  xor g_131734_(_070223_, _075170_, _075174_);
  or g_131735_(_069849_, _075174_, _075175_);
  not g_131736_(_075175_, _075176_);
  xor g_131737_(_069860_, _075174_, _075177_);
  or g_131738_(_069475_, _075177_, _075178_);
  not g_131739_(_075178_, _075179_);
  xor g_131740_(_069486_, _075177_, _075180_);
  not g_131741_(_075180_, _075181_);
  or g_131742_(_069112_, _075180_, _075182_);
  xor g_131743_(_069112_, _075180_, _075183_);
  xor g_131744_(_069112_, _075181_, _075185_);
  or g_131745_(_068749_, _075185_, _075186_);
  not g_131746_(_075186_, _075187_);
  xor g_131747_(_068749_, _075183_, _075188_);
  not g_131748_(_075188_, _075189_);
  or g_131749_(_068386_, _075188_, _075190_);
  xor g_131750_(_068386_, _075188_, _075191_);
  xor g_131751_(_068386_, _075189_, _075192_);
  or g_131752_(_068023_, _075192_, _075193_);
  xor g_131753_(_068023_, _075191_, _075194_);
  not g_131754_(_075194_, _075196_);
  or g_131755_(_067660_, _075194_, _075197_);
  xor g_131756_(_067660_, _075194_, _075198_);
  xor g_131757_(_067660_, _075196_, _075199_);
  or g_131758_(_067297_, _075199_, _075200_);
  xor g_131759_(_067297_, _075198_, _075201_);
  not g_131760_(_075201_, _075202_);
  or g_131761_(_066934_, _075201_, _075203_);
  xor g_131762_(_066934_, _075202_, _075204_);
  not g_131763_(_075204_, _075205_);
  or g_131764_(_066571_, _075204_, _075207_);
  xor g_131765_(_066571_, _075204_, _075208_);
  xor g_131766_(_066571_, _075205_, _075209_);
  or g_131767_(_066208_, _075209_, _075210_);
  not g_131768_(_075210_, _075211_);
  xor g_131769_(_066208_, _075208_, _075212_);
  or g_131770_(_065834_, _075212_, _075213_);
  xor g_131771_(_065845_, _075212_, _075214_);
  not g_131772_(_075214_, _075215_);
  or g_131773_(_065471_, _075214_, _075216_);
  xor g_131774_(_065471_, _075214_, _075218_);
  xor g_131775_(_065471_, _075215_, _075219_);
  or g_131776_(_065108_, _075219_, _075220_);
  xor g_131777_(_065108_, _075218_, _075221_);
  not g_131778_(_075221_, _075222_);
  or g_131779_(_064745_, _075221_, _075223_);
  xor g_131780_(_064745_, _075221_, _075224_);
  xor g_131781_(_064745_, _075222_, _075225_);
  or g_131782_(_064382_, _075225_, _075226_);
  xor g_131783_(_064382_, _075224_, _075227_);
  not g_131784_(_075227_, _075229_);
  or g_131785_(_064019_, _075227_, _075230_);
  xor g_131786_(_064019_, _075227_, _075231_);
  xor g_131787_(_064019_, _075229_, _075232_);
  or g_131788_(_063656_, _075232_, _075233_);
  xor g_131789_(_063656_, _075231_, _075234_);
  or g_131790_(_063282_, _075234_, _075235_);
  xor g_131791_(_063293_, _075234_, _075236_);
  or g_131792_(_062908_, _075236_, _075237_);
  xor g_131793_(_062908_, _075236_, _075238_);
  xor g_131794_(_062919_, _075236_, _075240_);
  or g_131795_(_062545_, _075240_, _075241_);
  xor g_131796_(_062545_, _075238_, _075242_);
  not g_131797_(_075242_, _075243_);
  or g_131798_(_062182_, _075242_, _075244_);
  xor g_131799_(_062182_, _075242_, _075245_);
  xor g_131800_(_062182_, _075243_, _075246_);
  and g_131801_(_061819_, _075245_, _075247_);
  or g_131802_(_061808_, _075246_, _075248_);
  xor g_131803_(_061808_, _075245_, _075249_);
  not g_131804_(_075249_, _075251_);
  or g_131805_(_061445_, _075249_, _075252_);
  not g_131806_(_075252_, _075253_);
  xor g_131807_(_061445_, _075251_, _075254_);
  not g_131808_(_075254_, _075255_);
  or g_131809_(_061082_, _075254_, _075256_);
  xor g_131810_(_061082_, _075254_, _075257_);
  xor g_131811_(_061082_, _075255_, _075258_);
  or g_131812_(_060719_, _075258_, _075259_);
  not g_131813_(_075259_, _075260_);
  xor g_131814_(_060719_, _075257_, _075262_);
  or g_131815_(_060356_, _075262_, _075263_);
  not g_131816_(_075263_, _075264_);
  and g_131817_(_060356_, _075262_, _075265_);
  or g_131818_(_075264_, _075265_, _075266_);
  not g_131819_(_075266_, _075267_);
  or g_131820_(_059993_, _075266_, _075268_);
  xor g_131821_(_059993_, _075267_, _075269_);
  or g_131822_(_059630_, _075269_, _075270_);
  xor g_131823_(_059630_, _075269_, _075271_);
  not g_131824_(_075271_, _075273_);
  or g_131825_(_059267_, _075273_, _075274_);
  not g_131826_(_075274_, _075275_);
  xor g_131827_(_059267_, _075271_, _075276_);
  not g_131828_(_075276_, _075277_);
  or g_131829_(_058904_, _075276_, _075278_);
  xor g_131830_(_058904_, _075277_, _075279_);
  not g_131831_(_075279_, _075280_);
  or g_131832_(_058541_, _075279_, _075281_);
  xor g_131833_(_058541_, _075279_, _075282_);
  xor g_131834_(_058541_, _075280_, _075284_);
  or g_131835_(_058178_, _075284_, _075285_);
  xor g_131836_(_058178_, _075282_, _075286_);
  not g_131837_(_075286_, _075287_);
  or g_131838_(_057815_, _075286_, _075288_);
  xor g_131839_(_057815_, _075286_, _075289_);
  xor g_131840_(_057815_, _075287_, _075290_);
  or g_131841_(_057452_, _075290_, _075291_);
  xor g_131842_(_057452_, _075289_, _075292_);
  not g_131843_(_075292_, _075293_);
  or g_131844_(_057089_, _075292_, _075295_);
  xor g_131845_(_057089_, _075293_, _075296_);
  not g_131846_(_075296_, _075297_);
  or g_131847_(_056726_, _075296_, _075298_);
  xor g_131848_(_056726_, _075297_, _075299_);
  not g_131849_(_075299_, _075300_);
  or g_131850_(_056363_, _075299_, _075301_);
  xor g_131851_(_056363_, _075299_, _075302_);
  xor g_131852_(_056363_, _075300_, _075303_);
  or g_131853_(_056000_, _075303_, _075304_);
  xor g_131854_(_056000_, _075302_, _075306_);
  not g_131855_(_075306_, _075307_);
  or g_131856_(_055637_, _075306_, _075308_);
  xor g_131857_(_055637_, _075307_, _075309_);
  not g_131858_(_075309_, _075310_);
  or g_131859_(_055274_, _075309_, _075311_);
  xor g_131860_(_055274_, _075310_, _075312_);
  or g_131861_(_054911_, _075312_, _075313_);
  xor g_131862_(_054911_, _075312_, _075314_);
  not g_131863_(_075314_, _075315_);
  or g_131864_(_054548_, _075315_, _075317_);
  xor g_131865_(_054548_, _075314_, _075318_);
  not g_131866_(_075318_, _075319_);
  or g_131867_(_054185_, _075318_, _075320_);
  xor g_131868_(_054185_, _075319_, _075321_);
  not g_131869_(_075321_, _075322_);
  or g_131870_(_053822_, _075321_, _075323_);
  xor g_131871_(_053822_, _075322_, _075324_);
  not g_131872_(_075324_, _075325_);
  or g_131873_(_053459_, _075324_, _075326_);
  xor g_131874_(_053459_, _075324_, _075328_);
  xor g_131875_(_053459_, _075325_, _075329_);
  or g_131876_(_053096_, _075329_, _075330_);
  xor g_131877_(_053096_, _075328_, _075331_);
  not g_131878_(_075331_, _075332_);
  or g_131879_(_052733_, _075331_, _075333_);
  xor g_131880_(_052733_, _075331_, _075334_);
  xor g_131881_(_052733_, _075332_, _075335_);
  or g_131882_(_052370_, _075335_, _075336_);
  xor g_131883_(_052370_, _075334_, _075337_);
  not g_131884_(_075337_, _075339_);
  or g_131885_(_052007_, _075337_, _075340_);
  xor g_131886_(_052007_, _075339_, _075341_);
  not g_131887_(_075341_, _075342_);
  or g_131888_(_051644_, _075341_, _075343_);
  xor g_131889_(_051644_, _075342_, _075344_);
  or g_131890_(_051281_, _075344_, _075345_);
  xor g_131891_(_051281_, _075344_, _075346_);
  not g_131892_(_075346_, _075347_);
  or g_131893_(_050918_, _075347_, _075348_);
  xor g_131894_(_050918_, _075346_, _075350_);
  not g_131895_(_075350_, _075351_);
  or g_131896_(_050555_, _075350_, _075352_);
  xor g_131897_(_050555_, _075351_, _075353_);
  or g_131898_(_050192_, _075353_, _075354_);
  not g_131899_(_075354_, _075355_);
  xor g_131900_(_050192_, _075353_, out[960]);
  and g_131901_(_075330_, _075333_, _075356_);
  and g_131902_(_075323_, _075326_, _075357_);
  and g_131903_(_075311_, _075313_, _075358_);
  and g_131904_(_075237_, _075241_, _075360_);
  and g_131905_(_075220_, _075223_, _075361_);
  and g_131906_(_075130_, _075133_, _075362_);
  not g_131907_(_075362_, _075363_);
  and g_131908_(_075123_, _075126_, _075364_);
  and g_131909_(_075049_, _075053_, _075365_);
  not g_131910_(_075365_, _075366_);
  and g_131911_(_075035_, _075038_, _075367_);
  not g_131912_(_075367_, _075368_);
  and g_131913_(_075000_, _075003_, _075369_);
  and g_131914_(_074978_, _074981_, _075371_);
  not g_131915_(_075371_, _075372_);
  and g_131916_(_074959_, _074961_, _075373_);
  and g_131917_(_074948_, _074950_, _075374_);
  and g_131918_(_074882_, _074885_, _075375_);
  and g_131919_(_074823_, _074825_, _075376_);
  and g_131920_(_074751_, _074754_, _075377_);
  and g_131921_(_074709_, _074716_, _075378_);
  and g_131922_(_074702_, _074705_, _075379_);
  and g_131923_(_074655_, _074660_, _075380_);
  and g_131924_(_074563_, _074566_, _075382_);
  and g_131925_(_074556_, _074559_, _075383_);
  and g_131926_(_074550_, _074553_, _075384_);
  and g_131927_(_074386_, _074388_, _075385_);
  and g_131928_(_074380_, _074383_, _075386_);
  and g_131929_(_074362_, _074365_, _075387_);
  and g_131930_(_074342_, _074344_, _075388_);
  and g_131931_(_074327_, _074332_, _075389_);
  and g_131932_(_074290_, _074292_, _075390_);
  and g_131933_(_074267_, _074269_, _075391_);
  and g_131934_(_074252_, _074254_, _075393_);
  and g_131935_(_074168_, _074170_, _075394_);
  not g_131936_(_075394_, _075395_);
  and g_131937_(_074103_, _074107_, _075396_);
  and g_131938_(_074075_, _074077_, _075397_);
  and g_131939_(_073999_, _074002_, _075398_);
  and g_131940_(_073975_, _073980_, _075399_);
  and g_131941_(_073934_, _073937_, _075400_);
  and g_131942_(_073863_, _073866_, _075401_);
  and g_131943_(_073764_, _073768_, _075402_);
  and g_131944_(_073724_, _073728_, _075404_);
  and g_131945_(_073541_, _073544_, _075405_);
  not g_131946_(_075405_, _075406_);
  and g_131947_(_073477_, _073481_, _075407_);
  and g_131948_(_073452_, _073454_, _075408_);
  not g_131949_(_075408_, _075409_);
  and g_131950_(_073447_, _073450_, _075410_);
  and g_131951_(_073441_, _073443_, _075411_);
  and g_131952_(_073426_, _073429_, _075412_);
  not g_131953_(_075412_, _075413_);
  and g_131954_(_073382_, _073385_, _075415_);
  and g_131955_(_073375_, _073378_, _075416_);
  and g_131956_(_073344_, _073350_, _075417_);
  not g_131957_(_075417_, _075418_);
  and g_131958_(_073255_, _073257_, _075419_);
  and g_131959_(_073234_, _073238_, _075420_);
  not g_131960_(_075420_, _075421_);
  and g_131961_(_073185_, _073188_, _075422_);
  and g_131962_(_073154_, _073156_, _075423_);
  and g_131963_(_073148_, _073152_, _075424_);
  not g_131964_(_075424_, _075426_);
  and g_131965_(_073143_, _073146_, _075427_);
  and g_131966_(_073087_, _073090_, _075428_);
  and g_131967_(_073058_, _073063_, _075429_);
  not g_131968_(_075429_, _075430_);
  and g_131969_(_073040_, _073043_, _075431_);
  not g_131970_(_075431_, _075432_);
  and g_131971_(_072865_, _072867_, _075433_);
  not g_131972_(_075433_, _075434_);
  and g_131973_(_072751_, _072754_, _075435_);
  and g_131974_(_072700_, _072703_, _075437_);
  and g_131975_(_072580_, _072582_, _075438_);
  not g_131976_(_075438_, _075439_);
  and g_131977_(_072570_, _072573_, _075440_);
  and g_131978_(_072564_, _072568_, _075441_);
  and g_131979_(_072556_, _072561_, _075442_);
  and g_131980_(_072551_, _072553_, _075443_);
  not g_131981_(_075443_, _075444_);
  and g_131982_(_072547_, _072549_, _075445_);
  not g_131983_(_075445_, _075446_);
  and g_131984_(_072540_, _072543_, _075448_);
  not g_131985_(_075448_, _075449_);
  and g_131986_(_072536_, _072538_, _075450_);
  not g_131987_(_075450_, _075451_);
  and g_131988_(_072432_, _072510_, _075452_);
  or g_131989_(_072512_, _075452_, _075453_);
  not g_131990_(_075453_, _075454_);
  or g_131991_(_072516_, _075453_, _075455_);
  not g_131992_(_075455_, _075456_);
  or g_131993_(_072519_, _075453_, _075457_);
  xor g_131994_(_072519_, _075454_, _075459_);
  and g_131995_(_072516_, _075459_, _075460_);
  or g_131996_(_075456_, _075460_, _075461_);
  and g_131997_(_072523_, _072526_, _075462_);
  or g_131998_(_075461_, _075462_, _075463_);
  xor g_131999_(_075461_, _075462_, _075464_);
  not g_132000_(_075464_, _075465_);
  or g_132001_(_072534_, _075465_, _075466_);
  and g_132002_(_072528_, _072534_, _075467_);
  and g_132003_(_072529_, _075464_, _075468_);
  or g_132004_(_072528_, _075465_, _075470_);
  xor g_132005_(_075464_, _075467_, _075471_);
  xor g_132006_(_075451_, _075471_, _075472_);
  xor g_132007_(_075449_, _075472_, _075473_);
  xor g_132008_(_075446_, _075473_, _075474_);
  xor g_132009_(_075444_, _075474_, _075475_);
  xor g_132010_(_075444_, _075474_, _075476_);
  xor g_132011_(_075443_, _075474_, _075477_);
  xor g_132012_(_075442_, _075477_, _075478_);
  not g_132013_(_075478_, _075479_);
  xor g_132014_(_075441_, _075479_, _075481_);
  not g_132015_(_075481_, _075482_);
  xor g_132016_(_075440_, _075482_, _075483_);
  not g_132017_(_075483_, _075484_);
  or g_132018_(_072578_, _075483_, _075485_);
  and g_132019_(_072575_, _072578_, _075486_);
  or g_132020_(_072575_, _075483_, _075487_);
  xor g_132021_(_075484_, _075486_, _075488_);
  xor g_132022_(_075439_, _075488_, _075489_);
  not g_132023_(_075489_, _075490_);
  or g_132024_(_072586_, _075489_, _075492_);
  and g_132025_(_072584_, _072586_, _075493_);
  or g_132026_(_072584_, _075489_, _075494_);
  not g_132027_(_075494_, _075495_);
  xor g_132028_(_075490_, _075493_, _075496_);
  xor g_132029_(_075489_, _075493_, _075497_);
  or g_132030_(_072590_, _075496_, _075498_);
  xor g_132031_(_072590_, _075497_, _075499_);
  not g_132032_(_075499_, _075500_);
  or g_132033_(_072593_, _075499_, _075501_);
  xor g_132034_(_072593_, _075499_, _075503_);
  xor g_132035_(_072593_, _075500_, _075504_);
  or g_132036_(_072595_, _075504_, _075505_);
  xor g_132037_(_072595_, _075503_, _075506_);
  not g_132038_(_075506_, _075507_);
  or g_132039_(_072598_, _075506_, _075508_);
  xor g_132040_(_072598_, _075507_, _075509_);
  not g_132041_(_075509_, _075510_);
  and g_132042_(_072602_, _072604_, _075511_);
  or g_132043_(_072602_, _075509_, _075512_);
  or g_132044_(_072604_, _075509_, _075514_);
  xor g_132045_(_075510_, _075511_, _075515_);
  not g_132046_(_075515_, _075516_);
  and g_132047_(_072607_, _072611_, _075517_);
  xor g_132048_(_075516_, _075517_, _075518_);
  and g_132049_(_072614_, _072617_, _075519_);
  or g_132050_(_072607_, _075515_, _075520_);
  not g_132051_(_075520_, _075521_);
  or g_132052_(_072611_, _075515_, _075522_);
  xor g_132053_(_075518_, _075519_, _075523_);
  not g_132054_(_075523_, _075525_);
  and g_132055_(_072620_, _072624_, _075526_);
  xor g_132056_(_075523_, _075526_, _075527_);
  xor g_132057_(_075523_, _075526_, _075528_);
  not g_132058_(_075528_, _075529_);
  or g_132059_(_072620_, _075525_, _075530_);
  or g_132060_(_072624_, _075525_, _075531_);
  or g_132061_(_072627_, _075527_, _075532_);
  xor g_132062_(_072627_, _075528_, _075533_);
  xor g_132063_(_072627_, _075529_, _075534_);
  and g_132064_(_072629_, _075534_, _075536_);
  or g_132065_(_072630_, _075533_, _075537_);
  or g_132066_(_072629_, _075527_, _075538_);
  not g_132067_(_075538_, _075539_);
  and g_132068_(_075537_, _075538_, _075540_);
  or g_132069_(_075536_, _075539_, _075541_);
  and g_132070_(_072634_, _075541_, _075542_);
  or g_132071_(_072635_, _075540_, _075543_);
  or g_132072_(_072634_, _075534_, _075544_);
  not g_132073_(_075544_, _075545_);
  and g_132074_(_075543_, _075544_, _075547_);
  or g_132075_(_075542_, _075545_, _075548_);
  or g_132076_(_072637_, _075548_, _075549_);
  xor g_132077_(_072637_, _075547_, _075550_);
  not g_132078_(_075550_, _075551_);
  or g_132079_(_072640_, _075550_, _075552_);
  xor g_132080_(_072640_, _075550_, _075553_);
  xor g_132081_(_072640_, _075551_, _075554_);
  or g_132082_(_072644_, _075554_, _075555_);
  xor g_132083_(_072644_, _075553_, _075556_);
  not g_132084_(_075556_, _075558_);
  or g_132085_(_072647_, _075556_, _075559_);
  xor g_132086_(_072647_, _075556_, _075560_);
  xor g_132087_(_072647_, _075558_, _075561_);
  or g_132088_(_072650_, _075561_, _075562_);
  or g_132089_(_072653_, _075561_, _075563_);
  and g_132090_(_072650_, _072653_, _075564_);
  xor g_132091_(_075560_, _075564_, _075565_);
  not g_132092_(_075565_, _075566_);
  or g_132093_(_072656_, _075565_, _075567_);
  xor g_132094_(_072656_, _075565_, _075569_);
  xor g_132095_(_072656_, _075566_, _075570_);
  and g_132096_(_072658_, _075570_, _075571_);
  or g_132097_(_072659_, _075569_, _075572_);
  or g_132098_(_072658_, _075565_, _075573_);
  not g_132099_(_075573_, _075574_);
  and g_132100_(_075572_, _075573_, _075575_);
  or g_132101_(_075571_, _075574_, _075576_);
  and g_132102_(_072662_, _075576_, _075577_);
  or g_132103_(_072663_, _075575_, _075578_);
  or g_132104_(_072662_, _075571_, _075580_);
  not g_132105_(_075580_, _075581_);
  and g_132106_(_075578_, _075580_, _075582_);
  or g_132107_(_075577_, _075581_, _075583_);
  and g_132108_(_072667_, _072670_, _075584_);
  not g_132109_(_075584_, _075585_);
  or g_132110_(_072667_, _075583_, _075586_);
  or g_132111_(_072670_, _075583_, _075587_);
  xor g_132112_(_075582_, _075585_, _075588_);
  not g_132113_(_075588_, _075589_);
  and g_132114_(_072672_, _072677_, _075591_);
  not g_132115_(_075591_, _075592_);
  and g_132116_(_072673_, _075588_, _075593_);
  or g_132117_(_072677_, _075589_, _075594_);
  or g_132118_(_075589_, _075591_, _075595_);
  xor g_132119_(_075588_, _075592_, _075596_);
  not g_132120_(_075596_, _075597_);
  and g_132121_(_072681_, _075596_, _075598_);
  or g_132122_(_072680_, _075597_, _075599_);
  xor g_132123_(_072681_, _075596_, _075600_);
  xor g_132124_(_072680_, _075596_, _075602_);
  or g_132125_(_072688_, _075602_, _075603_);
  not g_132126_(_075603_, _075604_);
  or g_132127_(_072684_, _075597_, _075605_);
  xor g_132128_(_072684_, _075600_, _075606_);
  and g_132129_(_072688_, _075606_, _075607_);
  or g_132130_(_075604_, _075607_, _075608_);
  and g_132131_(_072690_, _075608_, _075609_);
  or g_132132_(_072690_, _075606_, _075610_);
  not g_132133_(_075610_, _075611_);
  or g_132134_(_075609_, _075611_, _075613_);
  and g_132135_(_072693_, _072696_, _075614_);
  not g_132136_(_075614_, _075615_);
  xor g_132137_(_075613_, _075615_, _075616_);
  not g_132138_(_075616_, _075617_);
  or g_132139_(_072700_, _075616_, _075618_);
  or g_132140_(_072703_, _075616_, _075619_);
  xor g_132141_(_075437_, _075617_, _075620_);
  xor g_132142_(_075437_, _075616_, _075621_);
  or g_132143_(_072705_, _075620_, _075622_);
  xor g_132144_(_072705_, _075621_, _075624_);
  or g_132145_(_072708_, _075624_, _075625_);
  xor g_132146_(_072708_, _075624_, _075626_);
  not g_132147_(_075626_, _075627_);
  or g_132148_(_072712_, _075627_, _075628_);
  not g_132149_(_075628_, _075629_);
  xor g_132150_(_072712_, _075626_, _075630_);
  not g_132151_(_075630_, _075631_);
  or g_132152_(_072714_, _075630_, _075632_);
  not g_132153_(_075632_, _075633_);
  xor g_132154_(_072714_, _075631_, _075635_);
  or g_132155_(_072716_, _075635_, _075636_);
  xor g_132156_(_072716_, _075635_, _075637_);
  not g_132157_(_075637_, _075638_);
  and g_132158_(_072719_, _072723_, _075639_);
  xor g_132159_(_075637_, _075639_, _075640_);
  not g_132160_(_075640_, _075641_);
  or g_132161_(_072725_, _075640_, _075642_);
  xor g_132162_(_072725_, _075640_, _075643_);
  xor g_132163_(_072725_, _075641_, _075644_);
  and g_132164_(_072727_, _075644_, _075646_);
  or g_132165_(_072728_, _075643_, _075647_);
  or g_132166_(_072727_, _075640_, _075648_);
  not g_132167_(_075648_, _075649_);
  and g_132168_(_075647_, _075648_, _075650_);
  or g_132169_(_075646_, _075649_, _075651_);
  and g_132170_(_072732_, _075651_, _075652_);
  or g_132171_(_072733_, _075650_, _075653_);
  or g_132172_(_072732_, _075644_, _075654_);
  not g_132173_(_075654_, _075655_);
  and g_132174_(_075653_, _075654_, _075657_);
  or g_132175_(_075652_, _075655_, _075658_);
  or g_132176_(_072735_, _075658_, _075659_);
  xor g_132177_(_072735_, _075657_, _075660_);
  and g_132178_(_072737_, _072740_, _075661_);
  not g_132179_(_075661_, _075662_);
  xor g_132180_(_075660_, _075662_, _075663_);
  or g_132181_(_072745_, _075663_, _075664_);
  xor g_132182_(_072744_, _075663_, _075665_);
  not g_132183_(_075665_, _075666_);
  and g_132184_(_072747_, _072749_, _075668_);
  xor g_132185_(_075665_, _075668_, _075669_);
  xor g_132186_(_075666_, _075668_, _075670_);
  or g_132187_(_075435_, _075670_, _075671_);
  xor g_132188_(_075435_, _075669_, _075672_);
  not g_132189_(_075672_, _075673_);
  or g_132190_(_072756_, _075672_, _075674_);
  xor g_132191_(_072756_, _075672_, _075675_);
  xor g_132192_(_072756_, _075673_, _075676_);
  and g_132193_(_072760_, _075675_, _075677_);
  or g_132194_(_072759_, _075676_, _075679_);
  or g_132195_(_072762_, _075676_, _075680_);
  xor g_132196_(_072762_, _075675_, _075681_);
  and g_132197_(_072759_, _075681_, _075682_);
  or g_132198_(_075677_, _075682_, _075683_);
  or g_132199_(_072767_, _075683_, _075684_);
  xor g_132200_(_072766_, _075683_, _075685_);
  or g_132201_(_072769_, _075685_, _075686_);
  xor g_132202_(_072770_, _075685_, _075687_);
  or g_132203_(_072772_, _075687_, _075688_);
  xor g_132204_(_072773_, _075687_, _075690_);
  or g_132205_(_072776_, _075690_, _075691_);
  xor g_132206_(_072777_, _075690_, _075692_);
  and g_132207_(_072780_, _075692_, _075693_);
  not g_132208_(_075693_, _075694_);
  or g_132209_(_072780_, _075690_, _075695_);
  not g_132210_(_075695_, _075696_);
  or g_132211_(_075693_, _075696_, _075697_);
  and g_132212_(_072782_, _075697_, _075698_);
  and g_132213_(_072783_, _075694_, _075699_);
  not g_132214_(_075699_, _075701_);
  or g_132215_(_075698_, _075699_, _075702_);
  or g_132216_(_072785_, _075702_, _075703_);
  xor g_132217_(_072787_, _075702_, _075704_);
  and g_132218_(_072791_, _075704_, _075705_);
  or g_132219_(_072791_, _075702_, _075706_);
  not g_132220_(_075706_, _075707_);
  or g_132221_(_075705_, _075707_, _075708_);
  or g_132222_(_072795_, _075708_, _075709_);
  not g_132223_(_075709_, _075710_);
  and g_132224_(_072793_, _075708_, _075712_);
  or g_132225_(_072793_, _075704_, _075713_);
  not g_132226_(_075713_, _075714_);
  or g_132227_(_075712_, _075714_, _075715_);
  and g_132228_(_072795_, _075715_, _075716_);
  or g_132229_(_075710_, _075716_, _075717_);
  and g_132230_(_072798_, _072800_, _075718_);
  not g_132231_(_075718_, _075719_);
  or g_132232_(_075717_, _075718_, _075720_);
  xor g_132233_(_075717_, _075719_, _075721_);
  not g_132234_(_075721_, _075723_);
  or g_132235_(_072802_, _075721_, _075724_);
  xor g_132236_(_072802_, _075721_, _075725_);
  xor g_132237_(_072802_, _075723_, _075726_);
  and g_132238_(_072805_, _075726_, _075727_);
  or g_132239_(_072806_, _075725_, _075728_);
  or g_132240_(_072805_, _075721_, _075729_);
  not g_132241_(_075729_, _075730_);
  and g_132242_(_075728_, _075729_, _075731_);
  or g_132243_(_075727_, _075730_, _075732_);
  or g_132244_(_072812_, _075732_, _075734_);
  not g_132245_(_075734_, _075735_);
  and g_132246_(_072809_, _075732_, _075736_);
  or g_132247_(_072810_, _075731_, _075737_);
  or g_132248_(_072809_, _075727_, _075738_);
  not g_132249_(_075738_, _075739_);
  and g_132250_(_075737_, _075738_, _075740_);
  or g_132251_(_075736_, _075739_, _075741_);
  and g_132252_(_072812_, _075741_, _075742_);
  or g_132253_(_072813_, _075740_, _075743_);
  and g_132254_(_075734_, _075743_, _075745_);
  or g_132255_(_075735_, _075742_, _075746_);
  and g_132256_(_072816_, _075746_, _075747_);
  or g_132257_(_072817_, _075745_, _075748_);
  or g_132258_(_072816_, _075741_, _075749_);
  not g_132259_(_075749_, _075750_);
  and g_132260_(_075748_, _075749_, _075751_);
  or g_132261_(_075747_, _075750_, _075752_);
  and g_132262_(_072821_, _072824_, _075753_);
  not g_132263_(_075753_, _075754_);
  xor g_132264_(_075751_, _075753_, _075756_);
  xor g_132265_(_075751_, _075754_, _075757_);
  or g_132266_(_072826_, _075756_, _075758_);
  not g_132267_(_075758_, _075759_);
  xor g_132268_(_072826_, _075757_, _075760_);
  and g_132269_(_072828_, _072832_, _075761_);
  not g_132270_(_075761_, _075762_);
  xor g_132271_(_075760_, _075762_, _075763_);
  not g_132272_(_075763_, _075764_);
  or g_132273_(_072838_, _075763_, _075765_);
  or g_132274_(_072835_, _075763_, _075767_);
  and g_132275_(_075765_, _075767_, _075768_);
  and g_132276_(_072835_, _072838_, _075769_);
  xor g_132277_(_075763_, _075769_, _075770_);
  xor g_132278_(_075764_, _075769_, _075771_);
  or g_132279_(_072842_, _075771_, _075772_);
  xor g_132280_(_072842_, _075770_, _075773_);
  not g_132281_(_075773_, _075774_);
  or g_132282_(_072845_, _075773_, _075775_);
  xor g_132283_(_072845_, _075773_, _075776_);
  xor g_132284_(_072845_, _075774_, _075778_);
  and g_132285_(_072848_, _072850_, _075779_);
  xor g_132286_(_075776_, _075779_, _075780_);
  and g_132287_(_072854_, _072857_, _075781_);
  not g_132288_(_075781_, _075782_);
  or g_132289_(_075780_, _075781_, _075783_);
  xor g_132290_(_075780_, _075782_, _075784_);
  or g_132291_(_072859_, _075784_, _075785_);
  not g_132292_(_075785_, _075786_);
  xor g_132293_(_072860_, _075784_, _075787_);
  or g_132294_(_072865_, _075787_, _075789_);
  or g_132295_(_072867_, _075787_, _075790_);
  not g_132296_(_075790_, _075791_);
  xor g_132297_(_075434_, _075787_, _075792_);
  or g_132298_(_072869_, _075792_, _075793_);
  xor g_132299_(_072869_, _075792_, _075794_);
  not g_132300_(_075794_, _075795_);
  or g_132301_(_072872_, _075794_, _075796_);
  or g_132302_(_072871_, _075792_, _075797_);
  and g_132303_(_075796_, _075797_, _075798_);
  and g_132304_(_072876_, _075798_, _075800_);
  not g_132305_(_075800_, _075801_);
  xor g_132306_(_072876_, _075798_, _075802_);
  and g_132307_(_072881_, _075802_, _075803_);
  and g_132308_(_072880_, _075798_, _075804_);
  or g_132309_(_072877_, _075801_, _075805_);
  or g_132310_(_075803_, _075804_, _075806_);
  not g_132311_(_075806_, _075807_);
  and g_132312_(_072888_, _075807_, _075808_);
  not g_132313_(_075808_, _075809_);
  and g_132314_(_072884_, _075806_, _075811_);
  or g_132315_(_072884_, _075802_, _075812_);
  not g_132316_(_075812_, _075813_);
  or g_132317_(_075811_, _075813_, _075814_);
  and g_132318_(_072887_, _075814_, _075815_);
  or g_132319_(_075808_, _075815_, _075816_);
  and g_132320_(_072890_, _075816_, _075817_);
  or g_132321_(_072890_, _075814_, _075818_);
  not g_132322_(_075818_, _075819_);
  or g_132323_(_072889_, _075814_, _075820_);
  or g_132324_(_075817_, _075819_, _075822_);
  not g_132325_(_075822_, _075823_);
  and g_132326_(_072892_, _072895_, _075824_);
  or g_132327_(_075822_, _075824_, _075825_);
  xor g_132328_(_075822_, _075824_, _075826_);
  xor g_132329_(_075823_, _075824_, _075827_);
  or g_132330_(_072899_, _075827_, _075828_);
  xor g_132331_(_072899_, _075826_, _075829_);
  and g_132332_(_072901_, _075829_, _075830_);
  and g_132333_(_072902_, _075826_, _075831_);
  or g_132334_(_072901_, _075827_, _075833_);
  or g_132335_(_075830_, _075831_, _075834_);
  or g_132336_(_072909_, _075834_, _075835_);
  not g_132337_(_075835_, _075836_);
  and g_132338_(_072905_, _075834_, _075837_);
  or g_132339_(_072905_, _075830_, _075838_);
  not g_132340_(_075838_, _075839_);
  or g_132341_(_075837_, _075839_, _075840_);
  and g_132342_(_072909_, _075840_, _075841_);
  or g_132343_(_075836_, _075841_, _075842_);
  or g_132344_(_072912_, _075840_, _075844_);
  xor g_132345_(_072913_, _075842_, _075845_);
  and g_132346_(_072916_, _072920_, _075846_);
  not g_132347_(_075846_, _075847_);
  or g_132348_(_072920_, _075845_, _075848_);
  or g_132349_(_072916_, _075845_, _075849_);
  xor g_132350_(_075845_, _075847_, _075850_);
  not g_132351_(_075850_, _075851_);
  and g_132352_(_072923_, _072926_, _075852_);
  or g_132353_(_075850_, _075852_, _075853_);
  xor g_132354_(_075850_, _075852_, _075855_);
  xor g_132355_(_075851_, _075852_, _075856_);
  or g_132356_(_072928_, _075856_, _075857_);
  xor g_132357_(_072928_, _075855_, _075858_);
  and g_132358_(_072932_, _075858_, _075859_);
  and g_132359_(_072933_, _075855_, _075860_);
  or g_132360_(_072932_, _075856_, _075861_);
  or g_132361_(_075859_, _075860_, _075862_);
  and g_132362_(_072936_, _072939_, _075863_);
  not g_132363_(_075863_, _075864_);
  xor g_132364_(_075862_, _075864_, _075866_);
  and g_132365_(_072943_, _072946_, _075867_);
  not g_132366_(_075867_, _075868_);
  or g_132367_(_072946_, _075866_, _075869_);
  or g_132368_(_072943_, _075866_, _075870_);
  xor g_132369_(_075866_, _075867_, _075871_);
  xor g_132370_(_075866_, _075868_, _075872_);
  and g_132371_(_072949_, _075871_, _075873_);
  or g_132372_(_072948_, _075872_, _075874_);
  xor g_132373_(_072948_, _075871_, _075875_);
  and g_132374_(_072954_, _075875_, _075877_);
  and g_132375_(_072953_, _075871_, _075878_);
  or g_132376_(_072954_, _075872_, _075879_);
  or g_132377_(_075877_, _075878_, _075880_);
  or g_132378_(_072959_, _075880_, _075881_);
  not g_132379_(_075881_, _075882_);
  and g_132380_(_072956_, _075880_, _075883_);
  or g_132381_(_072956_, _075875_, _075884_);
  not g_132382_(_075884_, _075885_);
  or g_132383_(_075883_, _075885_, _075886_);
  and g_132384_(_072959_, _075886_, _075888_);
  or g_132385_(_075882_, _075888_, _075889_);
  and g_132386_(_072963_, _075889_, _075890_);
  or g_132387_(_072963_, _075886_, _075891_);
  not g_132388_(_075891_, _075892_);
  or g_132389_(_075890_, _075892_, _075893_);
  or g_132390_(_072969_, _075893_, _075894_);
  not g_132391_(_075894_, _075895_);
  or g_132392_(_072967_, _075893_, _075896_);
  xor g_132393_(_072966_, _075893_, _075897_);
  and g_132394_(_072969_, _075897_, _075899_);
  or g_132395_(_075895_, _075899_, _075900_);
  and g_132396_(_072971_, _075900_, _075901_);
  not g_132397_(_075901_, _075902_);
  or g_132398_(_072971_, _075897_, _075903_);
  not g_132399_(_075903_, _075904_);
  and g_132400_(_075902_, _075903_, _075905_);
  or g_132401_(_075901_, _075904_, _075906_);
  and g_132402_(_072977_, _075905_, _075907_);
  not g_132403_(_075907_, _075908_);
  and g_132404_(_072974_, _075906_, _075910_);
  or g_132405_(_072974_, _075900_, _075911_);
  not g_132406_(_075911_, _075912_);
  or g_132407_(_075910_, _075912_, _075913_);
  not g_132408_(_075913_, _075914_);
  and g_132409_(_072976_, _075913_, _075915_);
  or g_132410_(_075907_, _075915_, _075916_);
  and g_132411_(_072980_, _075916_, _075917_);
  and g_132412_(_072981_, _075914_, _075918_);
  not g_132413_(_075918_, _075919_);
  or g_132414_(_075917_, _075918_, _075921_);
  and g_132415_(_072983_, _072987_, _075922_);
  not g_132416_(_075922_, _075923_);
  xor g_132417_(_075921_, _075923_, _075924_);
  and g_132418_(_072990_, _072993_, _075925_);
  not g_132419_(_075925_, _075926_);
  or g_132420_(_075924_, _075925_, _075927_);
  xor g_132421_(_075924_, _075926_, _075928_);
  not g_132422_(_075928_, _075929_);
  or g_132423_(_072997_, _075928_, _075930_);
  xor g_132424_(_072997_, _075928_, _075932_);
  xor g_132425_(_072997_, _075929_, _075933_);
  or g_132426_(_073000_, _075928_, _075934_);
  xor g_132427_(_073000_, _075932_, _075935_);
  and g_132428_(_073002_, _073005_, _075936_);
  xor g_132429_(_075935_, _075936_, _075937_);
  not g_132430_(_075937_, _075938_);
  or g_132431_(_073009_, _075938_, _075939_);
  not g_132432_(_075939_, _075940_);
  or g_132433_(_073012_, _075938_, _075941_);
  xor g_132434_(_073012_, _075937_, _075943_);
  and g_132435_(_073009_, _075943_, _075944_);
  or g_132436_(_075940_, _075944_, _075945_);
  not g_132437_(_075945_, _075946_);
  or g_132438_(_073015_, _075945_, _075947_);
  xor g_132439_(_073015_, _075946_, _075948_);
  and g_132440_(_073009_, _073012_, _075949_);
  xor g_132441_(_075937_, _075949_, _075950_);
  xor g_132442_(_073015_, _075950_, _075951_);
  and g_132443_(_073018_, _075948_, _075952_);
  or g_132444_(_073019_, _075951_, _075954_);
  or g_132445_(_073018_, _075945_, _075955_);
  not g_132446_(_075955_, _075956_);
  or g_132447_(_073018_, _075950_, _075957_);
  and g_132448_(_075954_, _075957_, _075958_);
  or g_132449_(_075952_, _075956_, _075959_);
  and g_132450_(_073023_, _073026_, _075960_);
  xor g_132451_(_075959_, _075960_, _075961_);
  xor g_132452_(_075958_, _075960_, _075962_);
  or g_132453_(_073031_, _073036_, _075963_);
  and g_132454_(_075961_, _075963_, _075965_);
  not g_132455_(_075965_, _075966_);
  xor g_132456_(_075962_, _075963_, _075967_);
  xor g_132457_(_075431_, _075967_, _075968_);
  xor g_132458_(_075432_, _075967_, _075969_);
  or g_132459_(_073045_, _075969_, _075970_);
  xor g_132460_(_073045_, _075969_, _075971_);
  xor g_132461_(_073045_, _075968_, _075972_);
  or g_132462_(_073047_, _075972_, _075973_);
  xor g_132463_(_073047_, _075971_, _075974_);
  not g_132464_(_075974_, _075976_);
  or g_132465_(_073051_, _075974_, _075977_);
  xor g_132466_(_073051_, _075974_, _075978_);
  xor g_132467_(_073051_, _075976_, _075979_);
  and g_132468_(_073054_, _073056_, _075980_);
  xor g_132469_(_075978_, _075980_, _075981_);
  not g_132470_(_075981_, _075982_);
  xor g_132471_(_075430_, _075981_, _075983_);
  or g_132472_(_073066_, _075983_, _075984_);
  not g_132473_(_075984_, _075985_);
  xor g_132474_(_073066_, _075983_, _075987_);
  not g_132475_(_075987_, _075988_);
  and g_132476_(_073069_, _073073_, _075989_);
  not g_132477_(_075989_, _075990_);
  or g_132478_(_073073_, _075988_, _075991_);
  or g_132479_(_073069_, _075983_, _075992_);
  and g_132480_(_075987_, _075990_, _075993_);
  xor g_132481_(_075987_, _075990_, _075994_);
  xor g_132482_(_075987_, _075989_, _075995_);
  or g_132483_(_073075_, _075995_, _075996_);
  xor g_132484_(_073075_, _075994_, _075998_);
  and g_132485_(_073078_, _075998_, _075999_);
  or g_132486_(_073078_, _075995_, _076000_);
  not g_132487_(_076000_, _076001_);
  or g_132488_(_075999_, _076001_, _076002_);
  and g_132489_(_073081_, _073084_, _076003_);
  xor g_132490_(_076002_, _076003_, _076004_);
  not g_132491_(_076004_, _076005_);
  xor g_132492_(_075428_, _076004_, _076006_);
  or g_132493_(_073092_, _076006_, _076007_);
  xor g_132494_(_073092_, _076006_, _076009_);
  xor g_132495_(_073093_, _076006_, _076010_);
  or g_132496_(_073097_, _076010_, _076011_);
  not g_132497_(_076011_, _076012_);
  xor g_132498_(_073097_, _076009_, _076013_);
  not g_132499_(_076013_, _076014_);
  or g_132500_(_073100_, _076013_, _076015_);
  xor g_132501_(_073100_, _076013_, _076016_);
  xor g_132502_(_073100_, _076014_, _076017_);
  or g_132503_(_073103_, _076017_, _076018_);
  not g_132504_(_076018_, _076020_);
  xor g_132505_(_073103_, _076016_, _076021_);
  and g_132506_(_073106_, _076021_, _076022_);
  not g_132507_(_076022_, _076023_);
  and g_132508_(_073107_, _076016_, _076024_);
  or g_132509_(_073106_, _076017_, _076025_);
  and g_132510_(_076023_, _076025_, _076026_);
  or g_132511_(_076022_, _076024_, _076027_);
  and g_132512_(_073112_, _076026_, _076028_);
  not g_132513_(_076028_, _076029_);
  and g_132514_(_073109_, _076027_, _076031_);
  or g_132515_(_073109_, _076021_, _076032_);
  not g_132516_(_076032_, _076033_);
  or g_132517_(_076031_, _076033_, _076034_);
  not g_132518_(_076034_, _076035_);
  and g_132519_(_073113_, _076034_, _076036_);
  or g_132520_(_076028_, _076036_, _076037_);
  and g_132521_(_073115_, _076037_, _076038_);
  and g_132522_(_073117_, _076035_, _076039_);
  not g_132523_(_076039_, _076040_);
  or g_132524_(_076038_, _076039_, _076042_);
  or g_132525_(_073122_, _076042_, _076043_);
  not g_132526_(_076043_, _076044_);
  and g_132527_(_073119_, _076042_, _076045_);
  or g_132528_(_073119_, _076037_, _076046_);
  not g_132529_(_076046_, _076047_);
  or g_132530_(_076045_, _076047_, _076048_);
  and g_132531_(_073122_, _076048_, _076049_);
  or g_132532_(_076044_, _076049_, _076050_);
  and g_132533_(_073124_, _076050_, _076051_);
  or g_132534_(_073124_, _076048_, _076053_);
  not g_132535_(_076053_, _076054_);
  or g_132536_(_076051_, _076054_, _076055_);
  not g_132537_(_076055_, _076056_);
  or g_132538_(_073131_, _076055_, _076057_);
  not g_132539_(_076057_, _076058_);
  xor g_132540_(_073128_, _076056_, _076059_);
  xor g_132541_(_073128_, _076055_, _076060_);
  and g_132542_(_073131_, _076059_, _076061_);
  or g_132543_(_073132_, _076060_, _076062_);
  and g_132544_(_076057_, _076062_, _076064_);
  or g_132545_(_076058_, _076061_, _076065_);
  or g_132546_(_073128_, _076050_, _076066_);
  or g_132547_(_073135_, _076064_, _076067_);
  or g_132548_(_073139_, _076065_, _076068_);
  or g_132549_(_073134_, _076059_, _076069_);
  and g_132550_(_076068_, _076069_, _076070_);
  and g_132551_(_076067_, _076069_, _076071_);
  or g_132552_(_073140_, _076071_, _076072_);
  and g_132553_(_076068_, _076072_, _076073_);
  not g_132554_(_076073_, _076075_);
  xor g_132555_(_075427_, _076073_, _076076_);
  xor g_132556_(_075426_, _076076_, _076077_);
  not g_132557_(_076077_, _076078_);
  xor g_132558_(_075423_, _076078_, _076079_);
  xor g_132559_(_075423_, _076077_, _076080_);
  or g_132560_(_073158_, _076079_, _076081_);
  not g_132561_(_076081_, _076082_);
  xor g_132562_(_073158_, _076080_, _076083_);
  and g_132563_(_073162_, _073165_, _076084_);
  not g_132564_(_076084_, _076086_);
  xor g_132565_(_076083_, _076086_, _076087_);
  not g_132566_(_076087_, _076088_);
  or g_132567_(_073167_, _076087_, _076089_);
  xor g_132568_(_073167_, _076087_, _076090_);
  xor g_132569_(_073167_, _076088_, _076091_);
  or g_132570_(_073172_, _076090_, _076092_);
  or g_132571_(_073170_, _076087_, _076093_);
  and g_132572_(_076092_, _076093_, _076094_);
  or g_132573_(_073175_, _076094_, _076095_);
  or g_132574_(_073174_, _076091_, _076097_);
  and g_132575_(_076095_, _076097_, _076098_);
  not g_132576_(_076098_, _076099_);
  and g_132577_(_073179_, _073181_, _076100_);
  and g_132578_(_073183_, _076098_, _076101_);
  not g_132579_(_076101_, _076102_);
  or g_132580_(_073179_, _076099_, _076103_);
  xor g_132581_(_076098_, _076100_, _076104_);
  not g_132582_(_076104_, _076105_);
  xor g_132583_(_075422_, _076104_, _076106_);
  xor g_132584_(_075422_, _076105_, _076108_);
  and g_132585_(_073191_, _076108_, _076109_);
  or g_132586_(_073191_, _076108_, _076110_);
  xor g_132587_(_073191_, _076106_, _076111_);
  not g_132588_(_076111_, _076112_);
  xor g_132589_(_073194_, _076112_, _076113_);
  xor g_132590_(_073194_, _076111_, _076114_);
  and g_132591_(_073197_, _076113_, _076115_);
  or g_132592_(_073198_, _076114_, _076116_);
  or g_132593_(_073197_, _076111_, _076117_);
  not g_132594_(_076117_, _076119_);
  and g_132595_(_076116_, _076117_, _076120_);
  or g_132596_(_076115_, _076119_, _076121_);
  or g_132597_(_073203_, _076121_, _076122_);
  not g_132598_(_076122_, _076123_);
  and g_132599_(_073200_, _076121_, _076124_);
  or g_132600_(_073201_, _076120_, _076125_);
  or g_132601_(_073200_, _076113_, _076126_);
  not g_132602_(_076126_, _076127_);
  and g_132603_(_076125_, _076126_, _076128_);
  or g_132604_(_076124_, _076127_, _076130_);
  and g_132605_(_073203_, _076130_, _076131_);
  or g_132606_(_073205_, _076128_, _076132_);
  and g_132607_(_076122_, _076132_, _076133_);
  or g_132608_(_076123_, _076131_, _076134_);
  or g_132609_(_073209_, _076134_, _076135_);
  xor g_132610_(_073209_, _076133_, _076136_);
  and g_132611_(_076122_, _076126_, _076137_);
  and g_132612_(_073211_, _076136_, _076138_);
  not g_132613_(_076138_, _076139_);
  and g_132614_(_073212_, _076133_, _076141_);
  or g_132615_(_073211_, _076134_, _076142_);
  and g_132616_(_076139_, _076142_, _076143_);
  or g_132617_(_076138_, _076141_, _076144_);
  and g_132618_(_073220_, _076143_, _076145_);
  not g_132619_(_076145_, _076146_);
  and g_132620_(_073216_, _076144_, _076147_);
  or g_132621_(_073217_, _076143_, _076148_);
  or g_132622_(_073216_, _076138_, _076149_);
  not g_132623_(_076149_, _076150_);
  and g_132624_(_076148_, _076149_, _076152_);
  or g_132625_(_076147_, _076150_, _076153_);
  and g_132626_(_073219_, _076153_, _076154_);
  or g_132627_(_076145_, _076154_, _076155_);
  and g_132628_(_073224_, _076155_, _076156_);
  or g_132629_(_073224_, _076153_, _076157_);
  not g_132630_(_076157_, _076158_);
  or g_132631_(_076156_, _076158_, _076159_);
  or g_132632_(_073231_, _076159_, _076160_);
  and g_132633_(_073222_, _076152_, _076161_);
  and g_132634_(_064145_, _076161_, _076163_);
  or g_132635_(_076156_, _076163_, _076164_);
  and g_132636_(_073228_, _073231_, _076165_);
  not g_132637_(_076165_, _076166_);
  or g_132638_(_073228_, _076159_, _076167_);
  xor g_132639_(_076164_, _076166_, _076168_);
  or g_132640_(_075420_, _076168_, _076169_);
  xor g_132641_(_075421_, _076168_, _076170_);
  or g_132642_(_073241_, _076170_, _076171_);
  not g_132643_(_076171_, _076172_);
  and g_132644_(_073241_, _076170_, _076174_);
  xor g_132645_(_073241_, _076170_, _076175_);
  or g_132646_(_076172_, _076174_, _076176_);
  and g_132647_(_073243_, _076176_, _076177_);
  or g_132648_(_073244_, _076175_, _076178_);
  or g_132649_(_073243_, _076170_, _076179_);
  not g_132650_(_076179_, _076180_);
  and g_132651_(_076178_, _076179_, _076181_);
  not g_132652_(_076181_, _076182_);
  and g_132653_(_073249_, _073252_, _076183_);
  xor g_132654_(_076181_, _076183_, _076185_);
  not g_132655_(_076185_, _076186_);
  or g_132656_(_075419_, _076185_, _076187_);
  xor g_132657_(_075419_, _076185_, _076188_);
  xor g_132658_(_075419_, _076186_, _076189_);
  or g_132659_(_073261_, _076189_, _076190_);
  xor g_132660_(_073261_, _076188_, _076191_);
  and g_132661_(_073264_, _073266_, _076192_);
  or g_132662_(_073266_, _076191_, _076193_);
  or g_132663_(_073264_, _076189_, _076194_);
  and g_132664_(_076193_, _076194_, _076196_);
  xor g_132665_(_076191_, _076192_, _076197_);
  not g_132666_(_076197_, _076198_);
  and g_132667_(_073268_, _073271_, _076199_);
  and g_132668_(_073272_, _076197_, _076200_);
  or g_132669_(_073271_, _076198_, _076201_);
  or g_132670_(_073268_, _076198_, _076202_);
  xor g_132671_(_076197_, _076199_, _076203_);
  and g_132672_(_073276_, _076203_, _076204_);
  or g_132673_(_073276_, _076203_, _076205_);
  not g_132674_(_076205_, _076207_);
  xor g_132675_(_073276_, _076203_, _076208_);
  or g_132676_(_076204_, _076207_, _076209_);
  and g_132677_(_073278_, _076209_, _076210_);
  or g_132678_(_073279_, _076208_, _076211_);
  or g_132679_(_073278_, _076203_, _076212_);
  not g_132680_(_076212_, _076213_);
  and g_132681_(_076211_, _076212_, _076214_);
  or g_132682_(_076210_, _076213_, _076215_);
  and g_132683_(_073282_, _073285_, _076216_);
  or g_132684_(_073285_, _076215_, _076218_);
  or g_132685_(_073282_, _076209_, _076219_);
  or g_132686_(_076215_, _076216_, _076220_);
  xor g_132687_(_076214_, _076216_, _076221_);
  not g_132688_(_076221_, _076222_);
  or g_132689_(_073288_, _076221_, _076223_);
  xor g_132690_(_073288_, _076221_, _076224_);
  xor g_132691_(_073288_, _076222_, _076225_);
  or g_132692_(_073291_, _076224_, _076226_);
  and g_132693_(_073291_, _076222_, _076227_);
  or g_132694_(_073290_, _076221_, _076229_);
  and g_132695_(_076226_, _076229_, _076230_);
  not g_132696_(_076230_, _076231_);
  and g_132697_(_073299_, _076230_, _076232_);
  or g_132698_(_073298_, _076231_, _076233_);
  xor g_132699_(_073296_, _076230_, _076234_);
  and g_132700_(_073298_, _076234_, _076235_);
  or g_132701_(_076232_, _076235_, _076236_);
  or g_132702_(_073306_, _076236_, _076237_);
  not g_132703_(_076237_, _076238_);
  and g_132704_(_073302_, _076236_, _076240_);
  or g_132705_(_073302_, _076234_, _076241_);
  not g_132706_(_076241_, _076242_);
  or g_132707_(_076238_, _076242_, _076243_);
  or g_132708_(_076240_, _076242_, _076244_);
  and g_132709_(_073306_, _076244_, _076245_);
  or g_132710_(_076238_, _076245_, _076246_);
  or g_132711_(_073308_, _076246_, _076247_);
  xor g_132712_(_073309_, _076246_, _076248_);
  and g_132713_(_073311_, _076248_, _076249_);
  or g_132714_(_073311_, _076246_, _076251_);
  not g_132715_(_076251_, _076252_);
  or g_132716_(_076249_, _076252_, _076253_);
  and g_132717_(_073313_, _073318_, _076254_);
  not g_132718_(_076254_, _076255_);
  xor g_132719_(_076253_, _076255_, _076256_);
  xor g_132720_(_076253_, _076254_, _076257_);
  or g_132721_(_073322_, _076256_, _076258_);
  xor g_132722_(_073322_, _076257_, _076259_);
  or g_132723_(_073324_, _076259_, _076260_);
  not g_132724_(_076260_, _076262_);
  or g_132725_(_073327_, _076259_, _076263_);
  xor g_132726_(_073328_, _076259_, _076264_);
  and g_132727_(_073324_, _076264_, _076265_);
  or g_132728_(_076262_, _076265_, _076266_);
  not g_132729_(_076266_, _076267_);
  or g_132730_(_073332_, _076266_, _076268_);
  xor g_132731_(_073332_, _076267_, _076269_);
  and g_132732_(_073335_, _073339_, _076270_);
  not g_132733_(_076270_, _076271_);
  xor g_132734_(_076269_, _076271_, _076273_);
  or g_132735_(_073341_, _076273_, _076274_);
  not g_132736_(_076274_, _076275_);
  xor g_132737_(_073342_, _076273_, _076276_);
  xor g_132738_(_075418_, _076276_, _076277_);
  or g_132739_(_073352_, _076277_, _076278_);
  not g_132740_(_076278_, _076279_);
  xor g_132741_(_073353_, _076277_, _076280_);
  and g_132742_(_073357_, _073360_, _076281_);
  xor g_132743_(_076280_, _076281_, _076282_);
  not g_132744_(_076282_, _076284_);
  or g_132745_(_073367_, _076284_, _076285_);
  not g_132746_(_076285_, _076286_);
  and g_132747_(_073364_, _073367_, _076287_);
  not g_132748_(_076287_, _076288_);
  or g_132749_(_076282_, _076288_, _076289_);
  and g_132750_(_073363_, _076282_, _076290_);
  not g_132751_(_076290_, _076291_);
  and g_132752_(_076289_, _076291_, _076292_);
  and g_132753_(_076285_, _076292_, _076293_);
  and g_132754_(_073372_, _076293_, _076295_);
  not g_132755_(_076295_, _076296_);
  xor g_132756_(_073371_, _076293_, _076297_);
  xor g_132757_(_076282_, _076287_, _076298_);
  xor g_132758_(_073371_, _076298_, _076299_);
  xor g_132759_(_075416_, _076299_, _076300_);
  xor g_132760_(_075415_, _076300_, _076301_);
  not g_132761_(_076301_, _076302_);
  or g_132762_(_073388_, _076302_, _076303_);
  not g_132763_(_076303_, _076304_);
  xor g_132764_(_073388_, _076301_, _076306_);
  or g_132765_(_073392_, _076306_, _076307_);
  xor g_132766_(_073393_, _076306_, _076308_);
  and g_132767_(_073395_, _076308_, _076309_);
  or g_132768_(_073395_, _076306_, _076310_);
  not g_132769_(_076310_, _076311_);
  or g_132770_(_076309_, _076311_, _076312_);
  and g_132771_(_073398_, _073401_, _076313_);
  xor g_132772_(_076312_, _076313_, _076314_);
  not g_132773_(_076314_, _076315_);
  and g_132774_(_073405_, _076314_, _076317_);
  or g_132775_(_073404_, _076315_, _076318_);
  or g_132776_(_073409_, _076315_, _076319_);
  xor g_132777_(_073409_, _076314_, _076320_);
  and g_132778_(_073404_, _076320_, _076321_);
  or g_132779_(_076317_, _076321_, _076322_);
  or g_132780_(_073411_, _076322_, _076323_);
  not g_132781_(_076323_, _076324_);
  and g_132782_(_073411_, _076322_, _076325_);
  xor g_132783_(_073411_, _076322_, _076326_);
  or g_132784_(_076324_, _076325_, _076328_);
  or g_132785_(_073415_, _076326_, _076329_);
  or g_132786_(_073416_, _076322_, _076330_);
  not g_132787_(_076330_, _076331_);
  and g_132788_(_076329_, _076330_, _076332_);
  and g_132789_(_073419_, _073422_, _076333_);
  xor g_132790_(_076332_, _076333_, _076334_);
  xor g_132791_(_075413_, _076334_, _076335_);
  not g_132792_(_076335_, _076336_);
  or g_132793_(_073432_, _076335_, _076337_);
  xor g_132794_(_073432_, _076335_, _076339_);
  xor g_132795_(_073432_, _076336_, _076340_);
  or g_132796_(_073436_, _076340_, _076341_);
  not g_132797_(_076341_, _076342_);
  or g_132798_(_073439_, _076340_, _076343_);
  not g_132799_(_076343_, _076344_);
  xor g_132800_(_073439_, _076339_, _076345_);
  and g_132801_(_073436_, _076345_, _076346_);
  or g_132802_(_076342_, _076346_, _076347_);
  and g_132803_(_073436_, _073439_, _076348_);
  xor g_132804_(_076339_, _076348_, _076350_);
  xor g_132805_(_076340_, _076348_, _076351_);
  xor g_132806_(_075411_, _076350_, _076352_);
  xor g_132807_(_075411_, _076351_, _076353_);
  xor g_132808_(_075410_, _076352_, _076354_);
  xor g_132809_(_075408_, _076354_, _076355_);
  xor g_132810_(_075409_, _076354_, _076356_);
  or g_132811_(_073458_, _076356_, _076357_);
  not g_132812_(_076357_, _076358_);
  xor g_132813_(_073458_, _076355_, _076359_);
  not g_132814_(_076359_, _076361_);
  or g_132815_(_073461_, _076359_, _076362_);
  xor g_132816_(_073461_, _076361_, _076363_);
  and g_132817_(_073464_, _073467_, _076364_);
  not g_132818_(_076364_, _076365_);
  or g_132819_(_073464_, _076363_, _076366_);
  or g_132820_(_073467_, _076363_, _076367_);
  not g_132821_(_076367_, _076368_);
  xor g_132822_(_076363_, _076365_, _076369_);
  not g_132823_(_076369_, _076370_);
  or g_132824_(_073474_, _076369_, _076372_);
  not g_132825_(_076372_, _076373_);
  and g_132826_(_073470_, _073474_, _076374_);
  and g_132827_(_076369_, _076374_, _076375_);
  and g_132828_(_073471_, _076370_, _076376_);
  not g_132829_(_076376_, _076377_);
  or g_132830_(_076375_, _076376_, _076378_);
  or g_132831_(_076373_, _076378_, _076379_);
  or g_132832_(_075407_, _076379_, _076380_);
  xor g_132833_(_076369_, _076374_, _076381_);
  xor g_132834_(_075407_, _076381_, _076383_);
  not g_132835_(_076383_, _076384_);
  or g_132836_(_073486_, _076383_, _076385_);
  not g_132837_(_076385_, _076386_);
  or g_132838_(_073483_, _076383_, _076387_);
  xor g_132839_(_073483_, _076383_, _076388_);
  xor g_132840_(_073483_, _076384_, _076389_);
  and g_132841_(_073486_, _076389_, _076390_);
  or g_132842_(_073487_, _076388_, _076391_);
  and g_132843_(_076385_, _076391_, _076392_);
  or g_132844_(_076386_, _076390_, _076394_);
  and g_132845_(_073489_, _073492_, _076395_);
  or g_132846_(_073492_, _076394_, _076396_);
  or g_132847_(_073489_, _076389_, _076397_);
  or g_132848_(_076394_, _076395_, _076398_);
  xor g_132849_(_076392_, _076395_, _076399_);
  not g_132850_(_076399_, _076400_);
  or g_132851_(_073495_, _076399_, _076401_);
  or g_132852_(_073498_, _076399_, _076402_);
  and g_132853_(_073495_, _073498_, _076403_);
  or g_132854_(_076399_, _076403_, _076405_);
  xor g_132855_(_076400_, _076403_, _076406_);
  and g_132856_(_073500_, _073504_, _076407_);
  xor g_132857_(_076399_, _076403_, _076408_);
  or g_132858_(_073500_, _076406_, _076409_);
  or g_132859_(_073504_, _076406_, _076410_);
  not g_132860_(_076410_, _076411_);
  and g_132861_(_076409_, _076410_, _076412_);
  xor g_132862_(_076407_, _076408_, _076413_);
  and g_132863_(_073507_, _073510_, _076414_);
  not g_132864_(_076414_, _076416_);
  or g_132865_(_073507_, _076413_, _076417_);
  or g_132866_(_073510_, _076413_, _076418_);
  xor g_132867_(_076413_, _076416_, _076419_);
  or g_132868_(_073513_, _076419_, _076420_);
  xor g_132869_(_073513_, _076419_, _076421_);
  xor g_132870_(_073514_, _076419_, _076422_);
  or g_132871_(_073517_, _076422_, _076423_);
  not g_132872_(_076423_, _076424_);
  or g_132873_(_073519_, _076422_, _076425_);
  xor g_132874_(_073519_, _076421_, _076427_);
  and g_132875_(_073517_, _076427_, _076428_);
  or g_132876_(_076424_, _076428_, _076429_);
  or g_132877_(_073522_, _076429_, _076430_);
  or g_132878_(_073525_, _076429_, _076431_);
  not g_132879_(_076431_, _076432_);
  and g_132880_(_073522_, _073525_, _076433_);
  xor g_132881_(_076429_, _076433_, _076434_);
  not g_132882_(_076434_, _076435_);
  or g_132883_(_073530_, _076435_, _076436_);
  not g_132884_(_076436_, _076438_);
  or g_132885_(_073527_, _076435_, _076439_);
  xor g_132886_(_073527_, _076434_, _076440_);
  and g_132887_(_073530_, _076440_, _076441_);
  or g_132888_(_076438_, _076441_, _076442_);
  and g_132889_(_073532_, _076442_, _076443_);
  or g_132890_(_073532_, _076440_, _076444_);
  not g_132891_(_076444_, _076445_);
  or g_132892_(_076443_, _076445_, _076446_);
  and g_132893_(_073536_, _073539_, _076447_);
  not g_132894_(_076447_, _076449_);
  xor g_132895_(_076446_, _076449_, _076450_);
  xor g_132896_(_075406_, _076450_, _076451_);
  xor g_132897_(_075405_, _076450_, _076452_);
  or g_132898_(_073548_, _076451_, _076453_);
  xor g_132899_(_073548_, _076452_, _076454_);
  or g_132900_(_073550_, _076454_, _076455_);
  xor g_132901_(_073550_, _076454_, _076456_);
  xor g_132902_(_073551_, _076454_, _076457_);
  and g_132903_(_073553_, _073555_, _076458_);
  xor g_132904_(_076457_, _076458_, _076460_);
  xor g_132905_(_076456_, _076458_, _076461_);
  and g_132906_(_073558_, _073563_, _076462_);
  and g_132907_(_073559_, _076460_, _076463_);
  not g_132908_(_076463_, _076464_);
  or g_132909_(_073563_, _076461_, _076465_);
  xor g_132910_(_076461_, _076462_, _076466_);
  xor g_132911_(_076460_, _076462_, _076467_);
  or g_132912_(_073565_, _076467_, _076468_);
  xor g_132913_(_073565_, _076466_, _076469_);
  and g_132914_(_073568_, _076469_, _076471_);
  or g_132915_(_073568_, _076467_, _076472_);
  not g_132916_(_076472_, _076473_);
  or g_132917_(_076471_, _076473_, _076474_);
  and g_132918_(_073571_, _076474_, _076475_);
  or g_132919_(_073571_, _076471_, _076476_);
  not g_132920_(_076476_, _076477_);
  or g_132921_(_076475_, _076477_, _076478_);
  or g_132922_(_073573_, _076478_, _076479_);
  xor g_132923_(_073574_, _076478_, _076480_);
  and g_132924_(_073579_, _073581_, _076482_);
  not g_132925_(_076482_, _076483_);
  xor g_132926_(_076480_, _076483_, _076484_);
  or g_132927_(_073579_, _076480_, _076485_);
  or g_132928_(_073581_, _076480_, _076486_);
  xor g_132929_(_076480_, _076482_, _076487_);
  or g_132930_(_073583_, _076484_, _076488_);
  xor g_132931_(_073583_, _076487_, _076489_);
  or g_132932_(_073586_, _076489_, _076490_);
  not g_132933_(_076490_, _076491_);
  or g_132934_(_073588_, _076489_, _076493_);
  not g_132935_(_076493_, _076494_);
  xor g_132936_(_073590_, _076489_, _076495_);
  and g_132937_(_073586_, _076495_, _076496_);
  or g_132938_(_076491_, _076496_, _076497_);
  or g_132939_(_073593_, _076497_, _076498_);
  or g_132940_(_073596_, _076497_, _076499_);
  xor g_132941_(_073596_, _076497_, _076500_);
  or g_132942_(_073594_, _076500_, _076501_);
  and g_132943_(_076498_, _076501_, _076502_);
  not g_132944_(_076502_, _076504_);
  and g_132945_(_073599_, _076502_, _076505_);
  not g_132946_(_076505_, _076506_);
  or g_132947_(_073603_, _076504_, _076507_);
  xor g_132948_(_073603_, _076502_, _076508_);
  and g_132949_(_073598_, _076508_, _076509_);
  or g_132950_(_076505_, _076509_, _076510_);
  not g_132951_(_076510_, _076511_);
  or g_132952_(_073605_, _076510_, _076512_);
  xor g_132953_(_073605_, _076510_, _076513_);
  xor g_132954_(_073605_, _076511_, _076515_);
  and g_132955_(_073608_, _073612_, _076516_);
  xor g_132956_(_076513_, _076516_, _076517_);
  and g_132957_(_073615_, _076517_, _076518_);
  or g_132958_(_073615_, _076517_, _076519_);
  not g_132959_(_076519_, _076520_);
  xor g_132960_(_073615_, _076517_, _076521_);
  or g_132961_(_076518_, _076520_, _076522_);
  and g_132962_(_073619_, _073623_, _076523_);
  xor g_132963_(_076521_, _076523_, _076524_);
  not g_132964_(_076524_, _076526_);
  and g_132965_(_073626_, _073629_, _076527_);
  xor g_132966_(_076526_, _076527_, _076528_);
  or g_132967_(_073631_, _076528_, _076529_);
  xor g_132968_(_073631_, _076528_, _076530_);
  not g_132969_(_076530_, _076531_);
  or g_132970_(_073626_, _076524_, _076532_);
  or g_132971_(_073629_, _076524_, _076533_);
  and g_132972_(_073635_, _076531_, _076534_);
  or g_132973_(_073636_, _076530_, _076535_);
  or g_132974_(_073635_, _076528_, _076537_);
  not g_132975_(_076537_, _076538_);
  and g_132976_(_076535_, _076537_, _076539_);
  or g_132977_(_076534_, _076538_, _076540_);
  and g_132978_(_073639_, _073643_, _076541_);
  xor g_132979_(_076539_, _076541_, _076542_);
  not g_132980_(_076542_, _076543_);
  and g_132981_(_073647_, _073650_, _076544_);
  or g_132982_(_076542_, _076544_, _076545_);
  xor g_132983_(_076543_, _076544_, _076546_);
  and g_132984_(_073653_, _073656_, _076548_);
  not g_132985_(_076548_, _076549_);
  xor g_132986_(_076546_, _076549_, _076550_);
  or g_132987_(_073658_, _076550_, _076551_);
  xor g_132988_(_073658_, _076550_, _076552_);
  not g_132989_(_076552_, _076553_);
  or g_132990_(_073656_, _076546_, _076554_);
  or g_132991_(_073653_, _076546_, _076555_);
  or g_132992_(_073660_, _076553_, _076556_);
  xor g_132993_(_073661_, _076552_, _076557_);
  xor g_132994_(_073660_, _076552_, _076559_);
  or g_132995_(_073665_, _076559_, _076560_);
  xor g_132996_(_073665_, _076557_, _076561_);
  not g_132997_(_076561_, _076562_);
  and g_132998_(_073669_, _073672_, _076563_);
  xor g_132999_(_076561_, _076563_, _076564_);
  xor g_133000_(_076562_, _076563_, _076565_);
  and g_133001_(_073679_, _076564_, _076566_);
  or g_133002_(_073678_, _076565_, _076567_);
  and g_133003_(_073674_, _073678_, _076568_);
  or g_133004_(_073674_, _076565_, _076570_);
  not g_133005_(_076570_, _076571_);
  xor g_133006_(_076564_, _076568_, _076572_);
  not g_133007_(_076572_, _076573_);
  or g_133008_(_073681_, _076572_, _076574_);
  xor g_133009_(_073681_, _076572_, _076575_);
  xor g_133010_(_073681_, _076573_, _076576_);
  and g_133011_(_073685_, _076576_, _076577_);
  or g_133012_(_073684_, _076575_, _076578_);
  or g_133013_(_073685_, _076572_, _076579_);
  not g_133014_(_076579_, _076581_);
  and g_133015_(_076578_, _076579_, _076582_);
  or g_133016_(_076577_, _076581_, _076583_);
  and g_133017_(_073687_, _076583_, _076584_);
  or g_133018_(_073689_, _076582_, _076585_);
  or g_133019_(_073687_, _076576_, _076586_);
  not g_133020_(_076586_, _076587_);
  and g_133021_(_076585_, _076586_, _076588_);
  or g_133022_(_076584_, _076587_, _076589_);
  or g_133023_(_073691_, _076589_, _076590_);
  xor g_133024_(_073691_, _076588_, _076592_);
  and g_133025_(_073694_, _076592_, _076593_);
  and g_133026_(_073695_, _076588_, _076594_);
  or g_133027_(_073694_, _076589_, _076595_);
  or g_133028_(_076593_, _076594_, _076596_);
  and g_133029_(_073698_, _076596_, _076597_);
  or g_133030_(_073698_, _076592_, _076598_);
  not g_133031_(_076598_, _076599_);
  or g_133032_(_076597_, _076599_, _076600_);
  not g_133033_(_076600_, _076601_);
  and g_133034_(_073702_, _073704_, _076603_);
  or g_133035_(_073702_, _076600_, _076604_);
  xor g_133036_(_076600_, _076603_, _076605_);
  xor g_133037_(_076601_, _076603_, _076606_);
  or g_133038_(_073707_, _076606_, _076607_);
  xor g_133039_(_073707_, _076605_, _076608_);
  not g_133040_(_076608_, _076609_);
  or g_133041_(_073711_, _076608_, _076610_);
  xor g_133042_(_073711_, _076609_, _076611_);
  or g_133043_(_073713_, _076611_, _076612_);
  xor g_133044_(_073713_, _076611_, _076614_);
  and g_133045_(_073716_, _073718_, _076615_);
  not g_133046_(_076615_, _076616_);
  xor g_133047_(_076614_, _076616_, _076617_);
  xor g_133048_(_076614_, _076615_, _076618_);
  xor g_133049_(_075404_, _076617_, _076619_);
  xor g_133050_(_075404_, _076618_, _076620_);
  or g_133051_(_073731_, _076619_, _076621_);
  xor g_133052_(_073731_, _076620_, _076622_);
  and g_133053_(_073735_, _076622_, _076623_);
  or g_133054_(_073735_, _076619_, _076625_);
  not g_133055_(_076625_, _076626_);
  or g_133056_(_076623_, _076626_, _076627_);
  and g_133057_(_073737_, _076627_, _076628_);
  or g_133058_(_073737_, _076623_, _076629_);
  not g_133059_(_076629_, _076630_);
  or g_133060_(_076628_, _076630_, _076631_);
  not g_133061_(_076631_, _076632_);
  or g_133062_(_073739_, _076631_, _076633_);
  xor g_133063_(_073739_, _076631_, _076634_);
  xor g_133064_(_073739_, _076632_, _076636_);
  and g_133065_(_073742_, _076636_, _076637_);
  or g_133066_(_073744_, _076634_, _076638_);
  or g_133067_(_073742_, _076631_, _076639_);
  not g_133068_(_076639_, _076640_);
  and g_133069_(_076638_, _076639_, _076641_);
  or g_133070_(_076637_, _076640_, _076642_);
  and g_133071_(_073746_, _073749_, _076643_);
  xor g_133072_(_076641_, _076643_, _076644_);
  and g_133073_(_073752_, _073755_, _076645_);
  or g_133074_(_073755_, _076644_, _076647_);
  or g_133075_(_073752_, _076644_, _076648_);
  or g_133076_(_076644_, _076645_, _076649_);
  xor g_133077_(_076644_, _076645_, _076650_);
  not g_133078_(_076650_, _076651_);
  or g_133079_(_073758_, _076651_, _076652_);
  xor g_133080_(_073758_, _076650_, _076653_);
  and g_133081_(_073761_, _076653_, _076654_);
  or g_133082_(_073761_, _076651_, _076655_);
  not g_133083_(_076655_, _076656_);
  or g_133084_(_076654_, _076656_, _076658_);
  xor g_133085_(_073761_, _076653_, _076659_);
  xor g_133086_(_075402_, _076658_, _076660_);
  xor g_133087_(_075402_, _076659_, _076661_);
  and g_133088_(_073772_, _076660_, _076662_);
  or g_133089_(_073771_, _076661_, _076663_);
  or g_133090_(_073774_, _076661_, _076664_);
  xor g_133091_(_073774_, _076661_, _076665_);
  not g_133092_(_076665_, _076666_);
  and g_133093_(_073771_, _076666_, _076667_);
  or g_133094_(_073772_, _076665_, _076669_);
  and g_133095_(_076663_, _076669_, _076670_);
  or g_133096_(_076662_, _076667_, _076671_);
  or g_133097_(_073777_, _076671_, _076672_);
  xor g_133098_(_073777_, _076670_, _076673_);
  and g_133099_(_073779_, _076673_, _076674_);
  or g_133100_(_073779_, _076671_, _076675_);
  not g_133101_(_076675_, _076676_);
  or g_133102_(_076674_, _076676_, _076677_);
  and g_133103_(_073782_, _076677_, _076678_);
  or g_133104_(_073782_, _076673_, _076680_);
  not g_133105_(_076680_, _076681_);
  or g_133106_(_076678_, _076681_, _076682_);
  not g_133107_(_076682_, _076683_);
  and g_133108_(_073785_, _073789_, _076684_);
  xor g_133109_(_076683_, _076684_, _076685_);
  xor g_133110_(_076682_, _076684_, _076686_);
  or g_133111_(_073791_, _076685_, _076687_);
  xor g_133112_(_073791_, _076686_, _076688_);
  or g_133113_(_073793_, _076688_, _076689_);
  xor g_133114_(_073794_, _076688_, _076691_);
  and g_133115_(_073799_, _076691_, _076692_);
  or g_133116_(_073799_, _076688_, _076693_);
  not g_133117_(_076693_, _076694_);
  or g_133118_(_076692_, _076694_, _076695_);
  and g_133119_(_073802_, _073805_, _076696_);
  not g_133120_(_076696_, _076697_);
  xor g_133121_(_076695_, _076697_, _076698_);
  or g_133122_(_073807_, _076698_, _076699_);
  xor g_133123_(_073808_, _076698_, _076700_);
  and g_133124_(_073813_, _073816_, _076702_);
  xor g_133125_(_076700_, _076702_, _076703_);
  and g_133126_(_073819_, _073823_, _076704_);
  not g_133127_(_076704_, _076705_);
  and g_133128_(_073824_, _076703_, _076706_);
  not g_133129_(_076706_, _076707_);
  and g_133130_(_073821_, _076703_, _076708_);
  not g_133131_(_076708_, _076709_);
  xor g_133132_(_076703_, _076705_, _076710_);
  xor g_133133_(_076703_, _076704_, _076711_);
  or g_133134_(_073828_, _076711_, _076713_);
  xor g_133135_(_073828_, _076710_, _076714_);
  or g_133136_(_073833_, _076714_, _076715_);
  or g_133137_(_073830_, _076714_, _076716_);
  and g_133138_(_073830_, _073833_, _076717_);
  not g_133139_(_076717_, _076718_);
  xor g_133140_(_076714_, _076717_, _076719_);
  xor g_133141_(_076714_, _076718_, _076720_);
  or g_133142_(_073836_, _076720_, _076721_);
  xor g_133143_(_073836_, _076719_, _076722_);
  not g_133144_(_076722_, _076724_);
  or g_133145_(_073839_, _076722_, _076725_);
  xor g_133146_(_073839_, _076724_, _076726_);
  or g_133147_(_073845_, _076726_, _076727_);
  not g_133148_(_076727_, _076728_);
  or g_133149_(_073843_, _076722_, _076729_);
  not g_133150_(_076729_, _076730_);
  and g_133151_(_073843_, _076726_, _076731_);
  or g_133152_(_076730_, _076731_, _076732_);
  and g_133153_(_073845_, _076732_, _076733_);
  or g_133154_(_076728_, _076733_, _076735_);
  and g_133155_(_073848_, _073850_, _076736_);
  not g_133156_(_076736_, _076737_);
  xor g_133157_(_076735_, _076737_, _076738_);
  or g_133158_(_073852_, _076738_, _076739_);
  not g_133159_(_076739_, _076740_);
  xor g_133160_(_073854_, _076738_, _076741_);
  and g_133161_(_073857_, _076741_, _076742_);
  or g_133162_(_073857_, _076738_, _076743_);
  not g_133163_(_076743_, _076744_);
  or g_133164_(_076742_, _076744_, _076746_);
  and g_133165_(_073859_, _073861_, _076747_);
  xor g_133166_(_076746_, _076747_, _076748_);
  not g_133167_(_076748_, _076749_);
  or g_133168_(_075401_, _076749_, _076750_);
  xor g_133169_(_075401_, _076748_, _076751_);
  or g_133170_(_073870_, _076751_, _076752_);
  not g_133171_(_076752_, _076753_);
  xor g_133172_(_073870_, _076751_, _076754_);
  xor g_133173_(_073869_, _076751_, _076755_);
  and g_133174_(_073872_, _076755_, _076757_);
  or g_133175_(_073873_, _076754_, _076758_);
  or g_133176_(_073872_, _076751_, _076759_);
  not g_133177_(_076759_, _076760_);
  and g_133178_(_076758_, _076759_, _076761_);
  or g_133179_(_076757_, _076760_, _076762_);
  and g_133180_(_073880_, _076761_, _076763_);
  not g_133181_(_076763_, _076764_);
  and g_133182_(_073877_, _076762_, _076765_);
  or g_133183_(_073877_, _076755_, _076766_);
  not g_133184_(_076766_, _076768_);
  or g_133185_(_076765_, _076768_, _076769_);
  not g_133186_(_076769_, _076770_);
  and g_133187_(_073881_, _076769_, _076771_);
  or g_133188_(_076763_, _076771_, _076772_);
  and g_133189_(_073883_, _076772_, _076773_);
  and g_133190_(_073884_, _076770_, _076774_);
  not g_133191_(_076774_, _076775_);
  or g_133192_(_076773_, _076774_, _076776_);
  or g_133193_(_073891_, _076776_, _076777_);
  not g_133194_(_076777_, _076779_);
  and g_133195_(_073888_, _076776_, _076780_);
  or g_133196_(_073888_, _076772_, _076781_);
  not g_133197_(_076781_, _076782_);
  or g_133198_(_076780_, _076782_, _076783_);
  and g_133199_(_073891_, _076783_, _076784_);
  or g_133200_(_076779_, _076784_, _076785_);
  and g_133201_(_073894_, _076785_, _076786_);
  or g_133202_(_073894_, _076783_, _076787_);
  not g_133203_(_076787_, _076788_);
  or g_133204_(_076786_, _076788_, _076790_);
  not g_133205_(_076790_, _076791_);
  or g_133206_(_073899_, _076790_, _076792_);
  not g_133207_(_076792_, _076793_);
  or g_133208_(_073896_, _076790_, _076794_);
  xor g_133209_(_073896_, _076790_, _076795_);
  xor g_133210_(_073896_, _076791_, _076796_);
  and g_133211_(_073899_, _076796_, _076797_);
  or g_133212_(_073900_, _076795_, _076798_);
  and g_133213_(_076792_, _076798_, _076799_);
  or g_133214_(_076793_, _076797_, _076801_);
  or g_133215_(_073903_, _076799_, _076802_);
  or g_133216_(_073902_, _076796_, _076803_);
  and g_133217_(_076802_, _076803_, _076804_);
  and g_133218_(_073911_, _076804_, _076805_);
  not g_133219_(_076805_, _076806_);
  xor g_133220_(_073907_, _076804_, _076807_);
  and g_133221_(_073910_, _076807_, _076808_);
  or g_133222_(_076805_, _076808_, _076809_);
  or g_133223_(_073917_, _076809_, _076810_);
  not g_133224_(_076810_, _076812_);
  or g_133225_(_073917_, _076812_, _076813_);
  and g_133226_(_073914_, _076809_, _076814_);
  or g_133227_(_073914_, _076807_, _076815_);
  and g_133228_(_076810_, _076815_, _076816_);
  not g_133229_(_076816_, _076817_);
  or g_133230_(_076814_, _076817_, _076818_);
  and g_133231_(_076813_, _076818_, _076819_);
  or g_133232_(_073924_, _076819_, _076820_);
  not g_133233_(_076820_, _076821_);
  or g_133234_(_073921_, _076819_, _076823_);
  not g_133235_(_076823_, _076824_);
  and g_133236_(_073921_, _073924_, _076825_);
  not g_133237_(_076825_, _076826_);
  or g_133238_(_076819_, _076825_, _076827_);
  xor g_133239_(_076819_, _076826_, _076828_);
  not g_133240_(_076828_, _076829_);
  and g_133241_(_073927_, _073931_, _076830_);
  or g_133242_(_073931_, _076828_, _076831_);
  or g_133243_(_073927_, _076828_, _076832_);
  xor g_133244_(_076829_, _076830_, _076834_);
  xor g_133245_(_075400_, _076834_, _076835_);
  not g_133246_(_076835_, _076836_);
  or g_133247_(_073940_, _076836_, _076837_);
  not g_133248_(_076837_, _076838_);
  xor g_133249_(_073940_, _076835_, _076839_);
  or g_133250_(_073944_, _076839_, _076840_);
  not g_133251_(_076840_, _076841_);
  xor g_133252_(_073944_, _076839_, _076842_);
  not g_133253_(_076842_, _076843_);
  and g_133254_(_073947_, _073950_, _076845_);
  xor g_133255_(_076842_, _076845_, _076846_);
  or g_133256_(_073958_, _076846_, _076847_);
  not g_133257_(_076847_, _076848_);
  and g_133258_(_073955_, _073958_, _076849_);
  not g_133259_(_076849_, _076850_);
  or g_133260_(_073955_, _076846_, _076851_);
  not g_133261_(_076851_, _076852_);
  xor g_133262_(_076846_, _076850_, _076853_);
  or g_133263_(_073961_, _076853_, _076854_);
  not g_133264_(_076854_, _076856_);
  and g_133265_(_073961_, _076853_, _076857_);
  xor g_133266_(_073961_, _076853_, _076858_);
  or g_133267_(_076856_, _076857_, _076859_);
  or g_133268_(_073965_, _076859_, _076860_);
  xor g_133269_(_073965_, _076859_, _076861_);
  xor g_133270_(_073965_, _076858_, _076862_);
  and g_133271_(_073968_, _073971_, _076863_);
  xor g_133272_(_076862_, _076863_, _076864_);
  not g_133273_(_076864_, _076865_);
  xor g_133274_(_075399_, _076864_, _076867_);
  or g_133275_(_073983_, _076867_, _076868_);
  xor g_133276_(_073984_, _076867_, _076869_);
  or g_133277_(_073989_, _076869_, _076870_);
  not g_133278_(_076870_, _076871_);
  xor g_133279_(_073990_, _076869_, _076872_);
  and g_133280_(_073987_, _076872_, _076873_);
  or g_133281_(_073987_, _076869_, _076874_);
  not g_133282_(_076874_, _076875_);
  or g_133283_(_076873_, _076875_, _076876_);
  or g_133284_(_073994_, _076876_, _076878_);
  not g_133285_(_076878_, _076879_);
  or g_133286_(_073997_, _076876_, _076880_);
  xor g_133287_(_073997_, _076876_, _076881_);
  not g_133288_(_076881_, _076882_);
  and g_133289_(_073994_, _076882_, _076883_);
  or g_133290_(_076879_, _076883_, _076884_);
  and g_133291_(_073994_, _073997_, _076885_);
  xor g_133292_(_076876_, _076885_, _076886_);
  xor g_133293_(_075398_, _076886_, _076887_);
  and g_133294_(_074005_, _074008_, _076889_);
  xor g_133295_(_076887_, _076889_, _076890_);
  or g_133296_(_074005_, _076887_, _076891_);
  not g_133297_(_076891_, _076892_);
  or g_133298_(_074008_, _076887_, _076893_);
  not g_133299_(_076893_, _076894_);
  and g_133300_(_074012_, _076890_, _076895_);
  not g_133301_(_076895_, _076896_);
  xor g_133302_(_074011_, _076890_, _076897_);
  and g_133303_(_074015_, _076897_, _076898_);
  and g_133304_(_074016_, _076890_, _076900_);
  not g_133305_(_076900_, _076901_);
  or g_133306_(_076898_, _076900_, _076902_);
  and g_133307_(_074020_, _076902_, _076903_);
  or g_133308_(_074020_, _076897_, _076904_);
  not g_133309_(_076904_, _076905_);
  or g_133310_(_076903_, _076905_, _076906_);
  not g_133311_(_076906_, _076907_);
  or g_133312_(_074022_, _076906_, _076908_);
  xor g_133313_(_074022_, _076907_, _076909_);
  or g_133314_(_074027_, _076909_, _076911_);
  and g_133315_(_074028_, _076909_, _076912_);
  and g_133316_(_074025_, _076909_, _076913_);
  not g_133317_(_076913_, _076914_);
  or g_133318_(_074025_, _076906_, _076915_);
  and g_133319_(_076911_, _076915_, _076916_);
  and g_133320_(_076914_, _076916_, _076917_);
  or g_133321_(_076912_, _076917_, _076918_);
  not g_133322_(_076918_, _076919_);
  or g_133323_(_074033_, _076919_, _076920_);
  xor g_133324_(_074034_, _076918_, _076922_);
  xor g_133325_(_074033_, _076918_, _076923_);
  or g_133326_(_074037_, _076922_, _076924_);
  or g_133327_(_074036_, _076919_, _076925_);
  and g_133328_(_076924_, _076925_, _076926_);
  or g_133329_(_074042_, _076926_, _076927_);
  or g_133330_(_074043_, _076923_, _076928_);
  not g_133331_(_076928_, _076929_);
  and g_133332_(_076927_, _076928_, _076930_);
  not g_133333_(_076930_, _076931_);
  or g_133334_(_074046_, _076931_, _076933_);
  xor g_133335_(_074046_, _076930_, _076934_);
  not g_133336_(_076934_, _076935_);
  and g_133337_(_074048_, _074052_, _076936_);
  or g_133338_(_076934_, _076936_, _076937_);
  xor g_133339_(_076934_, _076936_, _076938_);
  xor g_133340_(_076935_, _076936_, _076939_);
  or g_133341_(_074055_, _076939_, _076940_);
  xor g_133342_(_074055_, _076938_, _076941_);
  not g_133343_(_076941_, _076942_);
  or g_133344_(_074058_, _076941_, _076944_);
  xor g_133345_(_074058_, _076942_, _076945_);
  and g_133346_(_074061_, _074065_, _076946_);
  not g_133347_(_076946_, _076947_);
  xor g_133348_(_076945_, _076947_, _076948_);
  or g_133349_(_074071_, _076948_, _076949_);
  and g_133350_(_074068_, _074071_, _076950_);
  not g_133351_(_076950_, _076951_);
  or g_133352_(_074068_, _076948_, _076952_);
  not g_133353_(_076952_, _076953_);
  xor g_133354_(_076948_, _076950_, _076955_);
  xor g_133355_(_076948_, _076951_, _076956_);
  xor g_133356_(_075397_, _076955_, _076957_);
  xor g_133357_(_075397_, _076956_, _076958_);
  or g_133358_(_074082_, _076957_, _076959_);
  xor g_133359_(_074082_, _076957_, _076960_);
  xor g_133360_(_074082_, _076958_, _076961_);
  or g_133361_(_074085_, _076961_, _076962_);
  xor g_133362_(_074085_, _076960_, _076963_);
  and g_133363_(_074088_, _076963_, _076964_);
  or g_133364_(_074088_, _076961_, _076966_);
  not g_133365_(_076966_, _076967_);
  or g_133366_(_076964_, _076967_, _076968_);
  and g_133367_(_074090_, _074092_, _076969_);
  not g_133368_(_076969_, _076970_);
  xor g_133369_(_076968_, _076969_, _076971_);
  xor g_133370_(_076968_, _076970_, _076972_);
  or g_133371_(_074098_, _076972_, _076973_);
  not g_133372_(_076973_, _076974_);
  and g_133373_(_074096_, _074098_, _076975_);
  not g_133374_(_076975_, _076977_);
  and g_133375_(_076972_, _076975_, _076978_);
  or g_133376_(_076971_, _076977_, _076979_);
  or g_133377_(_074096_, _076972_, _076980_);
  not g_133378_(_076980_, _076981_);
  and g_133379_(_076979_, _076980_, _076982_);
  or g_133380_(_076978_, _076981_, _076983_);
  and g_133381_(_076973_, _076982_, _076984_);
  or g_133382_(_076974_, _076983_, _076985_);
  or g_133383_(_074100_, _076985_, _076986_);
  xor g_133384_(_074100_, _076984_, _076988_);
  xor g_133385_(_075396_, _076988_, _076989_);
  not g_133386_(_076989_, _076990_);
  or g_133387_(_074109_, _076990_, _076991_);
  xor g_133388_(_074109_, _076989_, _076992_);
  and g_133389_(_074111_, _076992_, _076993_);
  and g_133390_(_074112_, _076989_, _076994_);
  not g_133391_(_076994_, _076995_);
  or g_133392_(_076993_, _076994_, _076996_);
  and g_133393_(_074116_, _074119_, _076997_);
  not g_133394_(_076997_, _076999_);
  xor g_133395_(_076996_, _076999_, _077000_);
  or g_133396_(_074121_, _077000_, _077001_);
  xor g_133397_(_074122_, _077000_, _077002_);
  and g_133398_(_074125_, _074129_, _077003_);
  xor g_133399_(_077002_, _077003_, _077004_);
  not g_133400_(_077004_, _077005_);
  or g_133401_(_074132_, _077005_, _077006_);
  not g_133402_(_077006_, _077007_);
  xor g_133403_(_074132_, _077004_, _077008_);
  not g_133404_(_077008_, _077010_);
  or g_133405_(_074135_, _077008_, _077011_);
  xor g_133406_(_074135_, _077008_, _077012_);
  xor g_133407_(_074135_, _077010_, _077013_);
  or g_133408_(_074137_, _077013_, _077014_);
  xor g_133409_(_074137_, _077012_, _077015_);
  and g_133410_(_074140_, _074143_, _077016_);
  not g_133411_(_077016_, _077017_);
  or g_133412_(_074140_, _077015_, _077018_);
  or g_133413_(_074143_, _077015_, _077019_);
  or g_133414_(_077015_, _077016_, _077021_);
  xor g_133415_(_077015_, _077017_, _077022_);
  or g_133416_(_074145_, _077022_, _077023_);
  xor g_133417_(_074146_, _077022_, _077024_);
  or g_133418_(_074152_, _077024_, _077025_);
  not g_133419_(_077025_, _077026_);
  and g_133420_(_074149_, _077024_, _077027_);
  or g_133421_(_074149_, _077022_, _077028_);
  not g_133422_(_077028_, _077029_);
  or g_133423_(_077027_, _077029_, _077030_);
  and g_133424_(_074152_, _077030_, _077032_);
  or g_133425_(_077026_, _077032_, _077033_);
  and g_133426_(_074155_, _077033_, _077034_);
  or g_133427_(_074155_, _077030_, _077035_);
  not g_133428_(_077035_, _077036_);
  or g_133429_(_077034_, _077036_, _077037_);
  and g_133430_(_074157_, _074159_, _077038_);
  xor g_133431_(_077037_, _077038_, _077039_);
  not g_133432_(_077039_, _077040_);
  and g_133433_(_074163_, _074166_, _077041_);
  or g_133434_(_074166_, _077040_, _077043_);
  or g_133435_(_074163_, _077040_, _077044_);
  and g_133436_(_077043_, _077044_, _077045_);
  xor g_133437_(_077039_, _077041_, _077046_);
  or g_133438_(_075394_, _077046_, _077047_);
  xor g_133439_(_075395_, _077046_, _077048_);
  or g_133440_(_074174_, _077048_, _077049_);
  xor g_133441_(_074175_, _077048_, _077050_);
  not g_133442_(_077050_, _077051_);
  or g_133443_(_074177_, _077050_, _077052_);
  xor g_133444_(_074177_, _077050_, _077054_);
  xor g_133445_(_074177_, _077051_, _077055_);
  and g_133446_(_074179_, _074181_, _077056_);
  xor g_133447_(_077055_, _077056_, _077057_);
  xor g_133448_(_077054_, _077056_, _077058_);
  and g_133449_(_074188_, _077057_, _077059_);
  not g_133450_(_077059_, _077060_);
  xor g_133451_(_074187_, _077058_, _077061_);
  xor g_133452_(_074188_, _077058_, _077062_);
  and g_133453_(_074192_, _077062_, _077063_);
  or g_133454_(_074191_, _077061_, _077065_);
  and g_133455_(_074191_, _077057_, _077066_);
  or g_133456_(_074192_, _077058_, _077067_);
  and g_133457_(_077065_, _077067_, _077068_);
  or g_133458_(_077063_, _077066_, _077069_);
  and g_133459_(_074196_, _077069_, _077070_);
  or g_133460_(_074197_, _077068_, _077071_);
  or g_133461_(_074196_, _077062_, _077072_);
  not g_133462_(_077072_, _077073_);
  and g_133463_(_077071_, _077072_, _077074_);
  or g_133464_(_077070_, _077073_, _077076_);
  and g_133465_(_074203_, _077074_, _077077_);
  or g_133466_(_074202_, _077076_, _077078_);
  or g_133467_(_074200_, _077076_, _077079_);
  xor g_133468_(_074200_, _077074_, _077080_);
  and g_133469_(_074202_, _077080_, _077081_);
  or g_133470_(_077077_, _077081_, _077082_);
  and g_133471_(_074207_, _077082_, _077083_);
  or g_133472_(_074207_, _077080_, _077084_);
  not g_133473_(_077084_, _077085_);
  or g_133474_(_077083_, _077085_, _077087_);
  and g_133475_(_074210_, _077087_, _077088_);
  or g_133476_(_074210_, _077082_, _077089_);
  not g_133477_(_077089_, _077090_);
  or g_133478_(_077088_, _077090_, _077091_);
  and g_133479_(_074213_, _077091_, _077092_);
  or g_133480_(_074213_, _077087_, _077093_);
  not g_133481_(_077093_, _077094_);
  or g_133482_(_077092_, _077094_, _077095_);
  not g_133483_(_077095_, _077096_);
  and g_133484_(_074217_, _074220_, _077098_);
  xor g_133485_(_077096_, _077098_, _077099_);
  or g_133486_(_074222_, _077099_, _077100_);
  not g_133487_(_077100_, _077101_);
  xor g_133488_(_074223_, _077099_, _077102_);
  and g_133489_(_074226_, _077102_, _077103_);
  or g_133490_(_074226_, _077099_, _077104_);
  not g_133491_(_077104_, _077105_);
  or g_133492_(_077103_, _077105_, _077106_);
  and g_133493_(_074229_, _074232_, _077107_);
  not g_133494_(_077107_, _077109_);
  xor g_133495_(_077106_, _077107_, _077110_);
  xor g_133496_(_077106_, _077109_, _077111_);
  or g_133497_(_074235_, _077111_, _077112_);
  xor g_133498_(_074235_, _077110_, _077113_);
  or g_133499_(_074239_, _077113_, _077114_);
  or g_133500_(_074242_, _077113_, _077115_);
  and g_133501_(_074239_, _074242_, _077116_);
  not g_133502_(_077116_, _077117_);
  xor g_133503_(_077113_, _077116_, _077118_);
  xor g_133504_(_077113_, _077117_, _077120_);
  and g_133505_(_074245_, _077118_, _077121_);
  not g_133506_(_077121_, _077122_);
  or g_133507_(_074248_, _077120_, _077123_);
  not g_133508_(_077123_, _077124_);
  xor g_133509_(_074248_, _077118_, _077125_);
  and g_133510_(_074244_, _077125_, _077126_);
  or g_133511_(_077121_, _077126_, _077127_);
  and g_133512_(_074244_, _074248_, _077128_);
  xor g_133513_(_077120_, _077128_, _077129_);
  xor g_133514_(_075393_, _077129_, _077131_);
  or g_133515_(_074259_, _077131_, _077132_);
  not g_133516_(_077132_, _077133_);
  and g_133517_(_074257_, _074259_, _077134_);
  and g_133518_(_077131_, _077134_, _077135_);
  or g_133519_(_074257_, _077131_, _077136_);
  not g_133520_(_077136_, _077137_);
  or g_133521_(_077135_, _077137_, _077138_);
  or g_133522_(_077133_, _077138_, _077139_);
  or g_133523_(_074262_, _077139_, _077140_);
  xor g_133524_(_074262_, _077139_, _077142_);
  xor g_133525_(_074263_, _077139_, _077143_);
  xor g_133526_(_075391_, _077142_, _077144_);
  and g_133527_(_074273_, _077144_, _077145_);
  or g_133528_(_074273_, _077144_, _077146_);
  not g_133529_(_077146_, _077147_);
  xor g_133530_(_074273_, _077144_, _077148_);
  or g_133531_(_077145_, _077147_, _077149_);
  and g_133532_(_074276_, _074278_, _077150_);
  xor g_133533_(_077148_, _077150_, _077151_);
  or g_133534_(_074280_, _077151_, _077153_);
  not g_133535_(_077153_, _077154_);
  xor g_133536_(_074280_, _077151_, _077155_);
  xor g_133537_(_074281_, _077151_, _077156_);
  and g_133538_(_074285_, _074288_, _077157_);
  xor g_133539_(_077156_, _077157_, _077158_);
  xor g_133540_(_077155_, _077157_, _077159_);
  xor g_133541_(_075390_, _077158_, _077160_);
  xor g_133542_(_075390_, _077159_, _077161_);
  or g_133543_(_074295_, _077160_, _077162_);
  xor g_133544_(_074295_, _077161_, _077164_);
  and g_133545_(_074298_, _077164_, _077165_);
  or g_133546_(_074298_, _077160_, _077166_);
  not g_133547_(_077166_, _077167_);
  or g_133548_(_077165_, _077167_, _077168_);
  and g_133549_(_074301_, _077168_, _077169_);
  or g_133550_(_074301_, _077164_, _077170_);
  not g_133551_(_077170_, _077171_);
  or g_133552_(_077169_, _077171_, _077172_);
  and g_133553_(_074305_, _077172_, _077173_);
  or g_133554_(_074305_, _077168_, _077175_);
  not g_133555_(_077175_, _077176_);
  or g_133556_(_077173_, _077176_, _077177_);
  or g_133557_(_074307_, _077177_, _077178_);
  xor g_133558_(_074308_, _077177_, _077179_);
  or g_133559_(_074313_, _077179_, _077180_);
  not g_133560_(_077180_, _077181_);
  or g_133561_(_074311_, _077177_, _077182_);
  not g_133562_(_077182_, _077183_);
  and g_133563_(_074311_, _077179_, _077184_);
  or g_133564_(_077183_, _077184_, _077186_);
  and g_133565_(_074313_, _077186_, _077187_);
  or g_133566_(_077181_, _077187_, _077188_);
  or g_133567_(_074317_, _077188_, _077189_);
  xor g_133568_(_074318_, _077188_, _077190_);
  and g_133569_(_074320_, _077190_, _077191_);
  or g_133570_(_074320_, _077188_, _077192_);
  not g_133571_(_077192_, _077193_);
  or g_133572_(_077191_, _077193_, _077194_);
  not g_133573_(_077194_, _077195_);
  and g_133574_(_074322_, _074324_, _077197_);
  xor g_133575_(_077194_, _077197_, _077198_);
  xor g_133576_(_077195_, _077197_, _077199_);
  xor g_133577_(_075389_, _077198_, _077200_);
  xor g_133578_(_075389_, _077199_, _077201_);
  and g_133579_(_074336_, _074340_, _077202_);
  xor g_133580_(_077201_, _077202_, _077203_);
  xor g_133581_(_075388_, _077203_, _077204_);
  not g_133582_(_077204_, _077205_);
  and g_133583_(_074346_, _077204_, _077206_);
  or g_133584_(_074347_, _077205_, _077208_);
  xor g_133585_(_074346_, _077204_, _077209_);
  xor g_133586_(_074347_, _077204_, _077210_);
  or g_133587_(_074350_, _077210_, _077211_);
  xor g_133588_(_074350_, _077209_, _077212_);
  or g_133589_(_074353_, _077212_, _077213_);
  xor g_133590_(_074354_, _077212_, _077214_);
  not g_133591_(_077214_, _077215_);
  and g_133592_(_074356_, _074358_, _077216_);
  xor g_133593_(_077214_, _077216_, _077217_);
  xor g_133594_(_077215_, _077216_, _077219_);
  xor g_133595_(_075387_, _077217_, _077220_);
  or g_133596_(_074368_, _077220_, _077221_);
  xor g_133597_(_074368_, _077220_, _077222_);
  not g_133598_(_077222_, _077223_);
  or g_133599_(_074377_, _077223_, _077224_);
  not g_133600_(_077224_, _077225_);
  or g_133601_(_074372_, _077222_, _077226_);
  or g_133602_(_074373_, _077220_, _077227_);
  and g_133603_(_077226_, _077227_, _077228_);
  not g_133604_(_077228_, _077230_);
  and g_133605_(_074377_, _077230_, _077231_);
  or g_133606_(_074376_, _077228_, _077232_);
  and g_133607_(_077224_, _077227_, _077233_);
  not g_133608_(_077233_, _077234_);
  and g_133609_(_077224_, _077232_, _077235_);
  or g_133610_(_077225_, _077231_, _077236_);
  xor g_133611_(_075386_, _077235_, _077237_);
  not g_133612_(_077237_, _077238_);
  xor g_133613_(_075385_, _077238_, _077239_);
  xor g_133614_(_075385_, _077237_, _077241_);
  or g_133615_(_074394_, _077239_, _077242_);
  or g_133616_(_074390_, _077239_, _077243_);
  and g_133617_(_074390_, _074394_, _077244_);
  or g_133618_(_077239_, _077244_, _077245_);
  xor g_133619_(_077241_, _077244_, _077246_);
  not g_133620_(_077246_, _077247_);
  or g_133621_(_074396_, _077246_, _077248_);
  xor g_133622_(_074396_, _077246_, _077249_);
  xor g_133623_(_074396_, _077247_, _077250_);
  and g_133624_(_074400_, _077250_, _077252_);
  or g_133625_(_074399_, _077249_, _077253_);
  or g_133626_(_074400_, _077246_, _077254_);
  not g_133627_(_077254_, _077255_);
  and g_133628_(_077253_, _077254_, _077256_);
  or g_133629_(_077252_, _077255_, _077257_);
  and g_133630_(_074404_, _077257_, _077258_);
  or g_133631_(_074405_, _077256_, _077259_);
  or g_133632_(_074404_, _077250_, _077260_);
  not g_133633_(_077260_, _077261_);
  and g_133634_(_077259_, _077260_, _077263_);
  or g_133635_(_077258_, _077261_, _077264_);
  or g_133636_(_074407_, _077264_, _077265_);
  xor g_133637_(_074407_, _077264_, _077266_);
  xor g_133638_(_074407_, _077263_, _077267_);
  and g_133639_(_074410_, _077267_, _077268_);
  and g_133640_(_074411_, _077263_, _077269_);
  or g_133641_(_074410_, _077264_, _077270_);
  or g_133642_(_077268_, _077269_, _077271_);
  or g_133643_(_074419_, _077271_, _077272_);
  not g_133644_(_077272_, _077274_);
  and g_133645_(_074413_, _077271_, _077275_);
  and g_133646_(_074415_, _077266_, _077276_);
  not g_133647_(_077276_, _077277_);
  or g_133648_(_077275_, _077276_, _077278_);
  and g_133649_(_074419_, _077278_, _077279_);
  or g_133650_(_077274_, _077279_, _077280_);
  not g_133651_(_077280_, _077281_);
  or g_133652_(_074422_, _077280_, _077282_);
  xor g_133653_(_074422_, _077281_, _077283_);
  and g_133654_(_074426_, _074429_, _077285_);
  not g_133655_(_077285_, _077286_);
  or g_133656_(_074426_, _077283_, _077287_);
  or g_133657_(_074429_, _077283_, _077288_);
  not g_133658_(_077288_, _077289_);
  xor g_133659_(_077283_, _077286_, _077290_);
  and g_133660_(_074431_, _074434_, _077291_);
  not g_133661_(_077291_, _077292_);
  xor g_133662_(_077290_, _077292_, _077293_);
  or g_133663_(_074438_, _077293_, _077294_);
  not g_133664_(_077294_, _077296_);
  and g_133665_(_074438_, _077293_, _077297_);
  xor g_133666_(_074438_, _077293_, _077298_);
  or g_133667_(_077296_, _077297_, _077299_);
  or g_133668_(_074434_, _077290_, _077300_);
  or g_133669_(_074431_, _077290_, _077301_);
  or g_133670_(_074441_, _077299_, _077302_);
  xor g_133671_(_074441_, _077298_, _077303_);
  not g_133672_(_077303_, _077304_);
  or g_133673_(_074444_, _077303_, _077305_);
  xor g_133674_(_074444_, _077304_, _077307_);
  not g_133675_(_077307_, _077308_);
  or g_133676_(_074446_, _077307_, _077309_);
  xor g_133677_(_074446_, _077307_, _077310_);
  xor g_133678_(_074446_, _077308_, _077311_);
  and g_133679_(_074450_, _077311_, _077312_);
  or g_133680_(_074451_, _077310_, _077313_);
  or g_133681_(_074450_, _077307_, _077314_);
  not g_133682_(_077314_, _077315_);
  and g_133683_(_077313_, _077314_, _077316_);
  or g_133684_(_077312_, _077315_, _077318_);
  and g_133685_(_074454_, _074457_, _077319_);
  xor g_133686_(_077316_, _077319_, _077320_);
  not g_133687_(_077320_, _077321_);
  or g_133688_(_074464_, _077320_, _077322_);
  or g_133689_(_074461_, _077320_, _077323_);
  not g_133690_(_077323_, _077324_);
  and g_133691_(_074461_, _074464_, _077325_);
  or g_133692_(_077320_, _077325_, _077326_);
  xor g_133693_(_077321_, _077325_, _077327_);
  or g_133694_(_074466_, _077327_, _077329_);
  xor g_133695_(_074467_, _077327_, _077330_);
  and g_133696_(_074471_, _077330_, _077331_);
  or g_133697_(_074471_, _077327_, _077332_);
  not g_133698_(_077332_, _077333_);
  or g_133699_(_077331_, _077333_, _077334_);
  and g_133700_(_074474_, _074477_, _077335_);
  xor g_133701_(_077334_, _077335_, _077336_);
  and g_133702_(_074479_, _074484_, _077337_);
  or g_133703_(_074481_, _074485_, _077338_);
  xor g_133704_(_077336_, _077337_, _077340_);
  xor g_133705_(_077336_, _077338_, _077341_);
  or g_133706_(_074487_, _077340_, _077342_);
  xor g_133707_(_074487_, _077341_, _077343_);
  and g_133708_(_074492_, _077343_, _077344_);
  and g_133709_(_074490_, _077341_, _077345_);
  or g_133710_(_074492_, _077340_, _077346_);
  or g_133711_(_077344_, _077345_, _077347_);
  or g_133712_(_074497_, _077347_, _077348_);
  not g_133713_(_077348_, _077349_);
  and g_133714_(_074495_, _077347_, _077351_);
  or g_133715_(_074495_, _077343_, _077352_);
  not g_133716_(_077352_, _077353_);
  or g_133717_(_077351_, _077353_, _077354_);
  and g_133718_(_074497_, _077354_, _077355_);
  or g_133719_(_077349_, _077355_, _077356_);
  and g_133720_(_074500_, _077356_, _077357_);
  or g_133721_(_074500_, _077354_, _077358_);
  not g_133722_(_077358_, _077359_);
  or g_133723_(_077357_, _077359_, _077360_);
  and g_133724_(_074503_, _074506_, _077362_);
  not g_133725_(_077362_, _077363_);
  xor g_133726_(_077360_, _077363_, _077364_);
  not g_133727_(_077364_, _077365_);
  and g_133728_(_074509_, _074512_, _077366_);
  xor g_133729_(_077365_, _077366_, _077367_);
  or g_133730_(_074515_, _077367_, _077368_);
  xor g_133731_(_074515_, _077367_, _077369_);
  not g_133732_(_077369_, _077370_);
  and g_133733_(_074510_, _077365_, _077371_);
  not g_133734_(_077371_, _077373_);
  or g_133735_(_074512_, _077364_, _077374_);
  or g_133736_(_074519_, _077370_, _077375_);
  xor g_133737_(_074518_, _077369_, _077376_);
  not g_133738_(_077376_, _077377_);
  and g_133739_(_074521_, _074523_, _077378_);
  xor g_133740_(_077376_, _077378_, _077379_);
  not g_133741_(_077379_, _077380_);
  or g_133742_(_074527_, _077379_, _077381_);
  xor g_133743_(_074527_, _077380_, _077382_);
  not g_133744_(_077382_, _077384_);
  and g_133745_(_074530_, _074532_, _077385_);
  or g_133746_(_074532_, _077382_, _077386_);
  or g_133747_(_074530_, _077379_, _077387_);
  and g_133748_(_077386_, _077387_, _077388_);
  xor g_133749_(_077382_, _077385_, _077389_);
  xor g_133750_(_077384_, _077385_, _077390_);
  and g_133751_(_074534_, _074538_, _077391_);
  xor g_133752_(_077389_, _077391_, _077392_);
  xor g_133753_(_077390_, _077391_, _077393_);
  or g_133754_(_074541_, _077392_, _077395_);
  xor g_133755_(_074541_, _077392_, _077396_);
  xor g_133756_(_074541_, _077393_, _077397_);
  or g_133757_(_074543_, _077397_, _077398_);
  not g_133758_(_077398_, _077399_);
  or g_133759_(_074547_, _077397_, _077400_);
  not g_133760_(_077400_, _077401_);
  xor g_133761_(_074547_, _077396_, _077402_);
  and g_133762_(_074543_, _077402_, _077403_);
  or g_133763_(_077399_, _077403_, _077404_);
  and g_133764_(_074543_, _074547_, _077406_);
  xor g_133765_(_077397_, _077406_, _077407_);
  xor g_133766_(_075384_, _077407_, _077408_);
  not g_133767_(_077408_, _077409_);
  xor g_133768_(_075383_, _077409_, _077410_);
  not g_133769_(_077410_, _077411_);
  or g_133770_(_074561_, _077410_, _077412_);
  not g_133771_(_077412_, _077413_);
  xor g_133772_(_074561_, _077411_, _077414_);
  not g_133773_(_077414_, _077415_);
  xor g_133774_(_075382_, _077415_, _077417_);
  not g_133775_(_077417_, _077418_);
  or g_133776_(_074570_, _077417_, _077419_);
  xor g_133777_(_074570_, _077418_, _077420_);
  not g_133778_(_077420_, _077421_);
  and g_133779_(_074573_, _074576_, _077422_);
  xor g_133780_(_077421_, _077422_, _077423_);
  not g_133781_(_077423_, _077424_);
  and g_133782_(_074584_, _077424_, _077425_);
  and g_133783_(_074578_, _074583_, _077426_);
  and g_133784_(_077423_, _077426_, _077428_);
  and g_133785_(_074580_, _077424_, _077429_);
  not g_133786_(_077429_, _077430_);
  or g_133787_(_077428_, _077429_, _077431_);
  or g_133788_(_077425_, _077431_, _077432_);
  or g_133789_(_074589_, _077432_, _077433_);
  or g_133790_(_074586_, _077432_, _077434_);
  xor g_133791_(_074587_, _077432_, _077435_);
  or g_133792_(_074593_, _077435_, _077436_);
  and g_133793_(_074589_, _074593_, _077437_);
  xor g_133794_(_077423_, _077426_, _077439_);
  xor g_133795_(_074587_, _077439_, _077440_);
  xor g_133796_(_074586_, _077439_, _077441_);
  xor g_133797_(_077437_, _077441_, _077442_);
  xor g_133798_(_077437_, _077440_, _077443_);
  or g_133799_(_074596_, _077443_, _077444_);
  xor g_133800_(_074596_, _077442_, _077445_);
  and g_133801_(_074598_, _077445_, _077446_);
  or g_133802_(_074598_, _077443_, _077447_);
  not g_133803_(_077447_, _077448_);
  or g_133804_(_077446_, _077448_, _077450_);
  or g_133805_(_074604_, _077450_, _077451_);
  not g_133806_(_077451_, _077452_);
  and g_133807_(_074600_, _077450_, _077453_);
  or g_133808_(_074600_, _077445_, _077454_);
  not g_133809_(_077454_, _077455_);
  or g_133810_(_077453_, _077455_, _077456_);
  and g_133811_(_074604_, _077456_, _077457_);
  or g_133812_(_077452_, _077457_, _077458_);
  and g_133813_(_074606_, _077458_, _077459_);
  or g_133814_(_074606_, _077456_, _077461_);
  not g_133815_(_077461_, _077462_);
  or g_133816_(_077459_, _077462_, _077463_);
  or g_133817_(_074608_, _077463_, _077464_);
  xor g_133818_(_074608_, _077463_, _077465_);
  xor g_133819_(_074609_, _077463_, _077466_);
  or g_133820_(_074614_, _077463_, _077467_);
  xor g_133821_(_074614_, _077465_, _077468_);
  and g_133822_(_074616_, _077468_, _077469_);
  or g_133823_(_074616_, _077466_, _077470_);
  not g_133824_(_077470_, _077472_);
  or g_133825_(_077469_, _077472_, _077473_);
  and g_133826_(_074619_, _077473_, _077474_);
  or g_133827_(_074619_, _077469_, _077475_);
  not g_133828_(_077475_, _077476_);
  or g_133829_(_077474_, _077476_, _077477_);
  and g_133830_(_074622_, _074625_, _077478_);
  not g_133831_(_077478_, _077479_);
  xor g_133832_(_077477_, _077478_, _077480_);
  xor g_133833_(_077477_, _077479_, _077481_);
  or g_133834_(_074631_, _077481_, _077483_);
  not g_133835_(_077483_, _077484_);
  and g_133836_(_074628_, _074631_, _077485_);
  not g_133837_(_077485_, _077486_);
  and g_133838_(_077481_, _077485_, _077487_);
  or g_133839_(_077480_, _077486_, _077488_);
  or g_133840_(_074628_, _077481_, _077489_);
  not g_133841_(_077489_, _077490_);
  and g_133842_(_077488_, _077489_, _077491_);
  or g_133843_(_077487_, _077490_, _077492_);
  and g_133844_(_077483_, _077491_, _077494_);
  or g_133845_(_077484_, _077492_, _077495_);
  or g_133846_(_074635_, _077495_, _077496_);
  xor g_133847_(_074635_, _077494_, _077497_);
  xor g_133848_(_077480_, _077485_, _077498_);
  xor g_133849_(_074635_, _077498_, _077499_);
  or g_133850_(_074637_, _077497_, _077500_);
  xor g_133851_(_074637_, _077499_, _077501_);
  or g_133852_(_074639_, _077501_, _077502_);
  xor g_133853_(_074639_, _077501_, _077503_);
  not g_133854_(_077503_, _077505_);
  and g_133855_(_074643_, _077503_, _077506_);
  not g_133856_(_077506_, _077507_);
  and g_133857_(_074647_, _077503_, _077508_);
  or g_133858_(_074646_, _077505_, _077509_);
  xor g_133859_(_074646_, _077503_, _077510_);
  and g_133860_(_074642_, _077510_, _077511_);
  or g_133861_(_077506_, _077511_, _077512_);
  and g_133862_(_074650_, _074653_, _077513_);
  xor g_133863_(_077512_, _077513_, _077514_);
  not g_133864_(_077514_, _077516_);
  xor g_133865_(_075380_, _077514_, _077517_);
  not g_133866_(_077517_, _077518_);
  and g_133867_(_074663_, _074665_, _077519_);
  xor g_133868_(_077518_, _077519_, _077520_);
  or g_133869_(_074668_, _077520_, _077521_);
  not g_133870_(_077521_, _077522_);
  xor g_133871_(_074669_, _077520_, _077523_);
  not g_133872_(_077523_, _077524_);
  or g_133873_(_074673_, _077523_, _077525_);
  not g_133874_(_077525_, _077527_);
  xor g_133875_(_074673_, _077524_, _077528_);
  not g_133876_(_077528_, _077529_);
  and g_133877_(_074676_, _074680_, _077530_);
  xor g_133878_(_077528_, _077530_, _077531_);
  xor g_133879_(_077529_, _077530_, _077532_);
  and g_133880_(_074682_, _074685_, _077533_);
  and g_133881_(_074683_, _077531_, _077534_);
  or g_133882_(_074682_, _077532_, _077535_);
  or g_133883_(_074685_, _077532_, _077536_);
  not g_133884_(_077536_, _077538_);
  xor g_133885_(_077531_, _077533_, _077539_);
  not g_133886_(_077539_, _077540_);
  or g_133887_(_074687_, _077539_, _077541_);
  xor g_133888_(_074687_, _077540_, _077542_);
  not g_133889_(_077542_, _077543_);
  and g_133890_(_074690_, _074693_, _077544_);
  or g_133891_(_074693_, _077542_, _077545_);
  or g_133892_(_074690_, _077542_, _077546_);
  xor g_133893_(_077543_, _077544_, _077547_);
  not g_133894_(_077547_, _077549_);
  and g_133895_(_074696_, _074698_, _077550_);
  or g_133896_(_074698_, _077547_, _077551_);
  or g_133897_(_074696_, _077547_, _077552_);
  and g_133898_(_077551_, _077552_, _077553_);
  xor g_133899_(_077549_, _077550_, _077554_);
  not g_133900_(_077554_, _077555_);
  xor g_133901_(_075379_, _077555_, _077556_);
  not g_133902_(_077556_, _077557_);
  or g_133903_(_074707_, _077556_, _077558_);
  xor g_133904_(_074707_, _077557_, _077560_);
  not g_133905_(_077560_, _077561_);
  xor g_133906_(_075378_, _077561_, _077562_);
  not g_133907_(_077562_, _077563_);
  or g_133908_(_074719_, _077562_, _077564_);
  xor g_133909_(_074719_, _077563_, _077565_);
  not g_133910_(_077565_, _077566_);
  and g_133911_(_074726_, _077566_, _077567_);
  not g_133912_(_077567_, _077568_);
  and g_133913_(_074721_, _077565_, _077569_);
  or g_133914_(_074721_, _077562_, _077571_);
  not g_133915_(_077571_, _077572_);
  or g_133916_(_077569_, _077572_, _077573_);
  and g_133917_(_074725_, _077573_, _077574_);
  or g_133918_(_077567_, _077574_, _077575_);
  and g_133919_(_074729_, _074732_, _077576_);
  xor g_133920_(_077575_, _077576_, _077577_);
  not g_133921_(_077577_, _077578_);
  or g_133922_(_074735_, _077578_, _077579_);
  not g_133923_(_077579_, _077580_);
  xor g_133924_(_074735_, _077577_, _077582_);
  not g_133925_(_077582_, _077583_);
  and g_133926_(_074738_, _074741_, _077584_);
  xor g_133927_(_077583_, _077584_, _077585_);
  or g_133928_(_074743_, _077585_, _077586_);
  not g_133929_(_077586_, _077587_);
  xor g_133930_(_074745_, _077585_, _077588_);
  and g_133931_(_074749_, _077588_, _077589_);
  or g_133932_(_074749_, _077585_, _077590_);
  not g_133933_(_077590_, _077591_);
  or g_133934_(_077589_, _077591_, _077593_);
  not g_133935_(_077593_, _077594_);
  xor g_133936_(_075377_, _077594_, _077595_);
  not g_133937_(_077595_, _077596_);
  and g_133938_(_074759_, _077596_, _077597_);
  or g_133939_(_074758_, _077595_, _077598_);
  or g_133940_(_074761_, _077595_, _077599_);
  xor g_133941_(_074761_, _077596_, _077600_);
  and g_133942_(_074758_, _077600_, _077601_);
  or g_133943_(_077597_, _077601_, _077602_);
  and g_133944_(_074758_, _074761_, _077604_);
  xor g_133945_(_077595_, _077604_, _077605_);
  or g_133946_(_074763_, _077602_, _077606_);
  xor g_133947_(_074763_, _077605_, _077607_);
  and g_133948_(_074767_, _077607_, _077608_);
  not g_133949_(_077608_, _077609_);
  or g_133950_(_074767_, _077602_, _077610_);
  not g_133951_(_077610_, _077611_);
  and g_133952_(_077609_, _077610_, _077612_);
  not g_133953_(_077612_, _077613_);
  and g_133954_(_074770_, _074772_, _077615_);
  xor g_133955_(_077612_, _077615_, _077616_);
  not g_133956_(_077616_, _077617_);
  or g_133957_(_074780_, _077616_, _077618_);
  not g_133958_(_077618_, _077619_);
  and g_133959_(_074778_, _074780_, _077620_);
  or g_133960_(_074778_, _077616_, _077621_);
  not g_133961_(_077621_, _077622_);
  xor g_133962_(_077617_, _077620_, _077623_);
  or g_133963_(_074782_, _077623_, _077624_);
  xor g_133964_(_074782_, _077623_, _077626_);
  not g_133965_(_077626_, _077627_);
  and g_133966_(_074784_, _074787_, _077628_);
  not g_133967_(_077628_, _077629_);
  or g_133968_(_074787_, _077627_, _077630_);
  or g_133969_(_074784_, _077623_, _077631_);
  or g_133970_(_077627_, _077628_, _077632_);
  not g_133971_(_077632_, _077633_);
  xor g_133972_(_077626_, _077629_, _077634_);
  xor g_133973_(_077626_, _077628_, _077635_);
  or g_133974_(_074791_, _077635_, _077637_);
  not g_133975_(_077637_, _077638_);
  xor g_133976_(_074791_, _077634_, _077639_);
  or g_133977_(_074793_, _077639_, _077640_);
  not g_133978_(_077640_, _077641_);
  or g_133979_(_074795_, _077639_, _077642_);
  xor g_133980_(_074796_, _077639_, _077643_);
  and g_133981_(_074793_, _077643_, _077644_);
  or g_133982_(_077641_, _077644_, _077645_);
  and g_133983_(_074798_, _074802_, _077646_);
  not g_133984_(_077646_, _077648_);
  or g_133985_(_074798_, _077645_, _077649_);
  or g_133986_(_074802_, _077645_, _077650_);
  and g_133987_(_077649_, _077650_, _077651_);
  xor g_133988_(_077645_, _077648_, _077652_);
  not g_133989_(_077652_, _077653_);
  and g_133990_(_074806_, _077653_, _077654_);
  not g_133991_(_077654_, _077655_);
  or g_133992_(_074808_, _077652_, _077656_);
  and g_133993_(_074805_, _074808_, _077657_);
  not g_133994_(_077657_, _077659_);
  and g_133995_(_074805_, _077652_, _077660_);
  and g_133996_(_077653_, _077659_, _077661_);
  and g_133997_(_074808_, _077660_, _077662_);
  or g_133998_(_077661_, _077662_, _077663_);
  xor g_133999_(_077652_, _077659_, _077664_);
  xor g_134000_(_077652_, _077657_, _077665_);
  or g_134001_(_074812_, _077663_, _077666_);
  xor g_134002_(_074812_, _077664_, _077667_);
  xor g_134003_(_074812_, _077665_, _077668_);
  and g_134004_(_074814_, _074816_, _077670_);
  xor g_134005_(_077667_, _077670_, _077671_);
  not g_134006_(_077671_, _077672_);
  or g_134007_(_074819_, _077671_, _077673_);
  xor g_134008_(_074819_, _077672_, _077674_);
  xor g_134009_(_075376_, _077674_, _077675_);
  not g_134010_(_077675_, _077676_);
  and g_134011_(_074828_, _077675_, _077677_);
  not g_134012_(_077677_, _077678_);
  xor g_134013_(_074827_, _077675_, _077679_);
  not g_134014_(_077679_, _077681_);
  and g_134015_(_074833_, _074835_, _077682_);
  xor g_134016_(_077679_, _077682_, _077683_);
  xor g_134017_(_077681_, _077682_, _077684_);
  or g_134018_(_074839_, _077684_, _077685_);
  or g_134019_(_074837_, _077684_, _077686_);
  and g_134020_(_074837_, _074839_, _077687_);
  not g_134021_(_077687_, _077688_);
  and g_134022_(_077683_, _077688_, _077689_);
  xor g_134023_(_077683_, _077687_, _077690_);
  or g_134024_(_074844_, _077690_, _077692_);
  xor g_134025_(_074842_, _077690_, _077693_);
  and g_134026_(_074846_, _077693_, _077694_);
  or g_134027_(_074846_, _077690_, _077695_);
  not g_134028_(_077695_, _077696_);
  or g_134029_(_077694_, _077696_, _077697_);
  and g_134030_(_074849_, _074852_, _077698_);
  xor g_134031_(_077697_, _077698_, _077699_);
  not g_134032_(_077699_, _077700_);
  or g_134033_(_074855_, _077700_, _077701_);
  not g_134034_(_077701_, _077703_);
  xor g_134035_(_074856_, _077699_, _077704_);
  xor g_134036_(_074855_, _077699_, _077705_);
  or g_134037_(_074860_, _077700_, _077706_);
  xor g_134038_(_074860_, _077705_, _077707_);
  xor g_134039_(_074860_, _077704_, _077708_);
  and g_134040_(_074863_, _077708_, _077709_);
  or g_134041_(_074864_, _077707_, _077710_);
  or g_134042_(_074863_, _077705_, _077711_);
  not g_134043_(_077711_, _077712_);
  and g_134044_(_077710_, _077711_, _077714_);
  or g_134045_(_077709_, _077712_, _077715_);
  or g_134046_(_074871_, _077715_, _077716_);
  or g_134047_(_074871_, _077714_, _077717_);
  not g_134048_(_077717_, _077718_);
  or g_134049_(_074868_, _077714_, _077719_);
  or g_134050_(_074867_, _077708_, _077720_);
  and g_134051_(_077716_, _077720_, _077721_);
  not g_134052_(_077721_, _077722_);
  and g_134053_(_077719_, _077721_, _077723_);
  or g_134054_(_077718_, _077723_, _077725_);
  not g_134055_(_077725_, _077726_);
  and g_134056_(_074873_, _074875_, _077727_);
  xor g_134057_(_077725_, _077727_, _077728_);
  not g_134058_(_077728_, _077729_);
  and g_134059_(_074878_, _074880_, _077730_);
  or g_134060_(_074880_, _077728_, _077731_);
  not g_134061_(_077731_, _077732_);
  or g_134062_(_074878_, _077728_, _077733_);
  not g_134063_(_077733_, _077734_);
  xor g_134064_(_077728_, _077730_, _077736_);
  xor g_134065_(_077729_, _077730_, _077737_);
  xor g_134066_(_075375_, _077736_, _077738_);
  not g_134067_(_077738_, _077739_);
  or g_134068_(_074889_, _077738_, _077740_);
  xor g_134069_(_074889_, _077738_, _077741_);
  xor g_134070_(_074889_, _077739_, _077742_);
  and g_134071_(_074893_, _077742_, _077743_);
  or g_134072_(_074892_, _077741_, _077744_);
  or g_134073_(_074893_, _077738_, _077745_);
  and g_134074_(_077744_, _077745_, _077747_);
  or g_134075_(_074896_, _077747_, _077748_);
  or g_134076_(_074897_, _077743_, _077749_);
  and g_134077_(_077748_, _077749_, _077750_);
  not g_134078_(_077750_, _077751_);
  or g_134079_(_074900_, _077751_, _077752_);
  xor g_134080_(_074900_, _077751_, _077753_);
  xor g_134081_(_074900_, _077750_, _077754_);
  or g_134082_(_074907_, _077754_, _077755_);
  or g_134083_(_074902_, _077753_, _077756_);
  or g_134084_(_074903_, _077751_, _077758_);
  and g_134085_(_077756_, _077758_, _077759_);
  or g_134086_(_074906_, _077759_, _077760_);
  and g_134087_(_077755_, _077760_, _077761_);
  not g_134088_(_077761_, _077762_);
  and g_134089_(_074906_, _077754_, _077763_);
  and g_134090_(_077755_, _077758_, _077764_);
  and g_134091_(_077756_, _077764_, _077765_);
  or g_134092_(_077763_, _077765_, _077766_);
  and g_134093_(_074911_, _077761_, _077767_);
  or g_134094_(_074912_, _077762_, _077769_);
  xor g_134095_(_074911_, _077766_, _077770_);
  xor g_134096_(_074912_, _077766_, _077771_);
  or g_134097_(_074915_, _077771_, _077772_);
  not g_134098_(_077772_, _077773_);
  or g_134099_(_074918_, _077771_, _077774_);
  not g_134100_(_077774_, _077775_);
  xor g_134101_(_074918_, _077770_, _077776_);
  and g_134102_(_074915_, _077776_, _077777_);
  or g_134103_(_077773_, _077777_, _077778_);
  not g_134104_(_077778_, _077780_);
  or g_134105_(_074921_, _077778_, _077781_);
  not g_134106_(_077781_, _077782_);
  xor g_134107_(_074921_, _077780_, _077783_);
  and g_134108_(_074924_, _077783_, _077784_);
  or g_134109_(_074924_, _077778_, _077785_);
  not g_134110_(_077785_, _077786_);
  or g_134111_(_077784_, _077786_, _077787_);
  not g_134112_(_077787_, _077788_);
  and g_134113_(_074927_, _074930_, _077789_);
  xor g_134114_(_077787_, _077789_, _077791_);
  xor g_134115_(_077788_, _077789_, _077792_);
  and g_134116_(_074934_, _074936_, _077793_);
  or g_134117_(_074936_, _077792_, _077794_);
  or g_134118_(_074934_, _077792_, _077795_);
  and g_134119_(_077794_, _077795_, _077796_);
  xor g_134120_(_077791_, _077793_, _077797_);
  not g_134121_(_077797_, _077798_);
  or g_134122_(_074938_, _077797_, _077799_);
  xor g_134123_(_074938_, _077798_, _077800_);
  and g_134124_(_074941_, _077800_, _077802_);
  or g_134125_(_074941_, _077797_, _077803_);
  not g_134126_(_077803_, _077804_);
  or g_134127_(_077802_, _077804_, _077805_);
  and g_134128_(_074945_, _077805_, _077806_);
  or g_134129_(_074945_, _077800_, _077807_);
  not g_134130_(_077807_, _077808_);
  or g_134131_(_077806_, _077808_, _077809_);
  xor g_134132_(_075374_, _077809_, _077810_);
  not g_134133_(_077810_, _077811_);
  and g_134134_(_074954_, _077810_, _077813_);
  or g_134135_(_074952_, _077811_, _077814_);
  xor g_134136_(_074952_, _077810_, _077815_);
  and g_134137_(_074957_, _077815_, _077816_);
  or g_134138_(_074957_, _077811_, _077817_);
  not g_134139_(_077817_, _077818_);
  or g_134140_(_077816_, _077818_, _077819_);
  not g_134141_(_077819_, _077820_);
  or g_134142_(_074959_, _077815_, _077821_);
  or g_134143_(_074961_, _077819_, _077822_);
  or g_134144_(_075373_, _077819_, _077824_);
  xor g_134145_(_075373_, _077820_, _077825_);
  or g_134146_(_074963_, _077825_, _077826_);
  xor g_134147_(_074965_, _077825_, _077827_);
  or g_134148_(_074967_, _077827_, _077828_);
  xor g_134149_(_074967_, _077827_, _077829_);
  and g_134150_(_074970_, _074973_, _077830_);
  xor g_134151_(_077829_, _077830_, _077831_);
  not g_134152_(_077831_, _077832_);
  xor g_134153_(_075372_, _077831_, _077833_);
  or g_134154_(_074984_, _077833_, _077835_);
  xor g_134155_(_074985_, _077833_, _077836_);
  not g_134156_(_077836_, _077837_);
  and g_134157_(_074990_, _074993_, _077838_);
  xor g_134158_(_077837_, _077838_, _077839_);
  or g_134159_(_074996_, _077839_, _077840_);
  xor g_134160_(_074998_, _077839_, _077841_);
  xor g_134161_(_075369_, _077841_, _077842_);
  not g_134162_(_077842_, _077843_);
  or g_134163_(_075006_, _077843_, _077844_);
  xor g_134164_(_075006_, _077842_, _077846_);
  and g_134165_(_075009_, _077846_, _077847_);
  and g_134166_(_075010_, _077842_, _077848_);
  not g_134167_(_077848_, _077849_);
  or g_134168_(_077847_, _077848_, _077850_);
  and g_134169_(_075013_, _075015_, _077851_);
  xor g_134170_(_077850_, _077851_, _077852_);
  and g_134171_(_075018_, _077852_, _077853_);
  not g_134172_(_077853_, _077854_);
  xor g_134173_(_075017_, _077852_, _077855_);
  and g_134174_(_075022_, _077855_, _077857_);
  and g_134175_(_075021_, _077852_, _077858_);
  not g_134176_(_077858_, _077859_);
  or g_134177_(_077857_, _077858_, _077860_);
  and g_134178_(_075024_, _077860_, _077861_);
  or g_134179_(_075024_, _077855_, _077862_);
  not g_134180_(_077862_, _077863_);
  or g_134181_(_077861_, _077863_, _077864_);
  not g_134182_(_077864_, _077865_);
  and g_134183_(_075026_, _075029_, _077866_);
  xor g_134184_(_077864_, _077866_, _077868_);
  xor g_134185_(_077865_, _077866_, _077869_);
  or g_134186_(_075033_, _077869_, _077870_);
  not g_134187_(_077870_, _077871_);
  xor g_134188_(_075033_, _077868_, _077872_);
  xor g_134189_(_075368_, _077872_, _077873_);
  or g_134190_(_075042_, _077873_, _077874_);
  not g_134191_(_077874_, _077875_);
  xor g_134192_(_075043_, _077873_, _077876_);
  and g_134193_(_075046_, _077876_, _077877_);
  or g_134194_(_075046_, _077873_, _077879_);
  not g_134195_(_077879_, _077880_);
  or g_134196_(_077877_, _077880_, _077881_);
  xor g_134197_(_075365_, _077881_, _077882_);
  xor g_134198_(_075366_, _077881_, _077883_);
  and g_134199_(_075056_, _075058_, _077884_);
  or g_134200_(_075058_, _077883_, _077885_);
  or g_134201_(_075056_, _077883_, _077886_);
  or g_134202_(_077883_, _077884_, _077887_);
  xor g_134203_(_077882_, _077884_, _077888_);
  or g_134204_(_075060_, _077888_, _077890_);
  xor g_134205_(_075061_, _077888_, _077891_);
  and g_134206_(_075065_, _077891_, _077892_);
  or g_134207_(_075065_, _077888_, _077893_);
  not g_134208_(_077893_, _077894_);
  or g_134209_(_077892_, _077894_, _077895_);
  and g_134210_(_075067_, _075070_, _077896_);
  not g_134211_(_077896_, _077897_);
  xor g_134212_(_077895_, _077896_, _077898_);
  xor g_134213_(_077895_, _077897_, _077899_);
  and g_134214_(_075073_, _075076_, _077901_);
  or g_134215_(_075076_, _077899_, _077902_);
  or g_134216_(_075073_, _077899_, _077903_);
  xor g_134217_(_077899_, _077901_, _077904_);
  xor g_134218_(_077898_, _077901_, _077905_);
  or g_134219_(_075078_, _077905_, _077906_);
  xor g_134220_(_075078_, _077904_, _077907_);
  and g_134221_(_075081_, _077907_, _077908_);
  or g_134222_(_075081_, _077905_, _077909_);
  not g_134223_(_077909_, _077910_);
  or g_134224_(_077908_, _077910_, _077912_);
  and g_134225_(_075084_, _077912_, _077913_);
  or g_134226_(_075084_, _077908_, _077914_);
  not g_134227_(_077914_, _077915_);
  or g_134228_(_077913_, _077915_, _077916_);
  or g_134229_(_075087_, _077916_, _077917_);
  xor g_134230_(_075088_, _077916_, _077918_);
  and g_134231_(_075092_, _075094_, _077919_);
  not g_134232_(_077919_, _077920_);
  xor g_134233_(_077918_, _077920_, _077921_);
  or g_134234_(_075097_, _077921_, _077923_);
  not g_134235_(_077923_, _077924_);
  xor g_134236_(_075098_, _077921_, _077925_);
  and g_134237_(_075100_, _077925_, _077926_);
  or g_134238_(_075100_, _077921_, _077927_);
  not g_134239_(_077927_, _077928_);
  or g_134240_(_077926_, _077928_, _077929_);
  and g_134241_(_075103_, _077929_, _077930_);
  or g_134242_(_075103_, _077926_, _077931_);
  not g_134243_(_077931_, _077932_);
  or g_134244_(_077930_, _077932_, _077934_);
  or g_134245_(_075105_, _077934_, _077935_);
  xor g_134246_(_075106_, _077934_, _077936_);
  or g_134247_(_075109_, _077936_, _077937_);
  not g_134248_(_077937_, _077938_);
  xor g_134249_(_075109_, _077936_, _077939_);
  and g_134250_(_075112_, _075115_, _077940_);
  xor g_134251_(_077939_, _077940_, _077941_);
  not g_134252_(_077941_, _077942_);
  and g_134253_(_075120_, _077942_, _077943_);
  xor g_134254_(_075120_, _077941_, _077945_);
  xor g_134255_(_075364_, _077945_, _077946_);
  xor g_134256_(_075362_, _077946_, _077947_);
  xor g_134257_(_075363_, _077946_, _077948_);
  or g_134258_(_075138_, _077947_, _077949_);
  not g_134259_(_077949_, _077950_);
  xor g_134260_(_075138_, _077948_, _077951_);
  or g_134261_(_075141_, _077951_, _077952_);
  not g_134262_(_077952_, _077953_);
  or g_134263_(_075144_, _077951_, _077954_);
  xor g_134264_(_075145_, _077951_, _077956_);
  and g_134265_(_075141_, _077956_, _077957_);
  or g_134266_(_077953_, _077957_, _077958_);
  or g_134267_(_075147_, _077958_, _077959_);
  xor g_134268_(_075148_, _077958_, _077960_);
  or g_134269_(_075154_, _077960_, _077961_);
  not g_134270_(_077961_, _077962_);
  and g_134271_(_075152_, _077960_, _077963_);
  or g_134272_(_075152_, _077958_, _077964_);
  not g_134273_(_077964_, _077965_);
  or g_134274_(_077963_, _077965_, _077967_);
  and g_134275_(_075154_, _077967_, _077968_);
  and g_134276_(_077961_, _077964_, _077969_);
  or g_134277_(_077962_, _077968_, _077970_);
  or g_134278_(_075158_, _077970_, _077971_);
  not g_134279_(_077971_, _077972_);
  xor g_134280_(_075157_, _077970_, _077973_);
  and g_134281_(_075160_, _077973_, _077974_);
  or g_134282_(_075160_, _077970_, _077975_);
  not g_134283_(_077975_, _077976_);
  or g_134284_(_077974_, _077976_, _077978_);
  and g_134285_(_075163_, _075166_, _077979_);
  not g_134286_(_077979_, _077980_);
  xor g_134287_(_077978_, _077980_, _077981_);
  or g_134288_(_075169_, _077981_, _077982_);
  xor g_134289_(_075169_, _077981_, _077983_);
  and g_134290_(_075172_, _075175_, _077984_);
  not g_134291_(_077984_, _077985_);
  xor g_134292_(_077983_, _077985_, _077986_);
  xor g_134293_(_077983_, _077984_, _077987_);
  or g_134294_(_075182_, _077987_, _077989_);
  not g_134295_(_077989_, _077990_);
  and g_134296_(_075178_, _075182_, _077991_);
  and g_134297_(_077987_, _077991_, _077992_);
  and g_134298_(_075179_, _077986_, _077993_);
  or g_134299_(_075178_, _077987_, _077994_);
  or g_134300_(_077992_, _077993_, _077995_);
  or g_134301_(_077990_, _077995_, _077996_);
  or g_134302_(_075186_, _077996_, _077997_);
  not g_134303_(_077997_, _077998_);
  xor g_134304_(_075187_, _077996_, _078000_);
  and g_134305_(_075190_, _078000_, _078001_);
  or g_134306_(_075190_, _077996_, _078002_);
  not g_134307_(_078002_, _078003_);
  or g_134308_(_078001_, _078003_, _078004_);
  and g_134309_(_075193_, _078004_, _078005_);
  or g_134310_(_075193_, _078000_, _078006_);
  not g_134311_(_078006_, _078007_);
  or g_134312_(_078005_, _078007_, _078008_);
  and g_134313_(_075197_, _075200_, _078009_);
  not g_134314_(_078009_, _078011_);
  xor g_134315_(_078008_, _078011_, _078012_);
  and g_134316_(_075203_, _075207_, _078013_);
  not g_134317_(_078013_, _078014_);
  or g_134318_(_075203_, _078012_, _078015_);
  or g_134319_(_075207_, _078012_, _078016_);
  xor g_134320_(_078012_, _078014_, _078017_);
  or g_134321_(_075210_, _078017_, _078018_);
  xor g_134322_(_075211_, _078017_, _078019_);
  or g_134323_(_075216_, _078019_, _078020_);
  not g_134324_(_078020_, _078022_);
  or g_134325_(_075213_, _078017_, _078023_);
  not g_134326_(_078023_, _078024_);
  and g_134327_(_075213_, _075216_, _078025_);
  not g_134328_(_078025_, _078026_);
  xor g_134329_(_078019_, _078026_, _078027_);
  not g_134330_(_078027_, _078028_);
  xor g_134331_(_075361_, _078028_, _078029_);
  xor g_134332_(_075361_, _078027_, _078030_);
  or g_134333_(_075226_, _078029_, _078031_);
  xor g_134334_(_075226_, _078030_, _078033_);
  and g_134335_(_075230_, _078033_, _078034_);
  or g_134336_(_075230_, _078029_, _078035_);
  not g_134337_(_078035_, _078036_);
  or g_134338_(_078034_, _078036_, _078037_);
  not g_134339_(_078037_, _078038_);
  and g_134340_(_075233_, _075235_, _078039_);
  xor g_134341_(_078037_, _078039_, _078040_);
  xor g_134342_(_078038_, _078039_, _078041_);
  or g_134343_(_075360_, _078041_, _078042_);
  xor g_134344_(_075360_, _078040_, _078044_);
  not g_134345_(_078044_, _078045_);
  or g_134346_(_075244_, _078044_, _078046_);
  xor g_134347_(_075244_, _078044_, _078047_);
  xor g_134348_(_075244_, _078045_, _078048_);
  or g_134349_(_075247_, _078047_, _078049_);
  or g_134350_(_075248_, _078044_, _078050_);
  not g_134351_(_078050_, _078051_);
  and g_134352_(_078049_, _078050_, _078052_);
  or g_134353_(_075253_, _078052_, _078053_);
  or g_134354_(_075252_, _078048_, _078055_);
  and g_134355_(_078053_, _078055_, _078056_);
  not g_134356_(_078056_, _078057_);
  or g_134357_(_075256_, _078057_, _078058_);
  not g_134358_(_078058_, _078059_);
  xor g_134359_(_075256_, _078056_, _078060_);
  or g_134360_(_075259_, _078060_, _078061_);
  xor g_134361_(_075260_, _078060_, _078062_);
  or g_134362_(_075268_, _078062_, _078063_);
  not g_134363_(_078063_, _078064_);
  or g_134364_(_075263_, _078062_, _078066_);
  xor g_134365_(_075264_, _078062_, _078067_);
  and g_134366_(_075268_, _078067_, _078068_);
  or g_134367_(_078064_, _078068_, _078069_);
  and g_134368_(_075270_, _078069_, _078070_);
  not g_134369_(_078070_, _078071_);
  or g_134370_(_075270_, _078067_, _078072_);
  not g_134371_(_078072_, _078073_);
  and g_134372_(_078071_, _078072_, _078074_);
  or g_134373_(_078070_, _078073_, _078075_);
  and g_134374_(_075274_, _078075_, _078077_);
  or g_134375_(_075275_, _078074_, _078078_);
  or g_134376_(_075274_, _078069_, _078079_);
  not g_134377_(_078079_, _078080_);
  and g_134378_(_078078_, _078079_, _078081_);
  or g_134379_(_078077_, _078080_, _078082_);
  or g_134380_(_075278_, _078082_, _078083_);
  xor g_134381_(_075278_, _078081_, _078084_);
  not g_134382_(_078084_, _078085_);
  or g_134383_(_075281_, _078084_, _078086_);
  xor g_134384_(_075281_, _078085_, _078088_);
  not g_134385_(_078088_, _078089_);
  and g_134386_(_075285_, _075288_, _078090_);
  xor g_134387_(_078089_, _078090_, _078091_);
  not g_134388_(_078091_, _078092_);
  or g_134389_(_075291_, _078091_, _078093_);
  xor g_134390_(_075291_, _078092_, _078094_);
  not g_134391_(_078094_, _078095_);
  and g_134392_(_075295_, _075298_, _078096_);
  xor g_134393_(_078095_, _078096_, _078097_);
  not g_134394_(_078097_, _078099_);
  or g_134395_(_075304_, _078097_, _078100_);
  or g_134396_(_075301_, _078097_, _078101_);
  and g_134397_(_075301_, _075304_, _078102_);
  or g_134398_(_078097_, _078102_, _078103_);
  xor g_134399_(_078097_, _078102_, _078104_);
  xor g_134400_(_078099_, _078102_, _078105_);
  or g_134401_(_075308_, _078105_, _078106_);
  xor g_134402_(_075308_, _078104_, _078107_);
  not g_134403_(_078107_, _078108_);
  or g_134404_(_075358_, _078107_, _078110_);
  xor g_134405_(_075358_, _078108_, _078111_);
  or g_134406_(_075317_, _078111_, _078112_);
  xor g_134407_(_075317_, _078111_, _078113_);
  not g_134408_(_078113_, _078114_);
  and g_134409_(_075320_, _078114_, _078115_);
  or g_134410_(_075320_, _078111_, _078116_);
  not g_134411_(_078116_, _078117_);
  or g_134412_(_078115_, _078117_, _078118_);
  not g_134413_(_078118_, _078119_);
  xor g_134414_(_075357_, _078119_, _078121_);
  not g_134415_(_078121_, _078122_);
  xor g_134416_(_075356_, _078122_, _078123_);
  xor g_134417_(_075356_, _078121_, _078124_);
  or g_134418_(_075336_, _078123_, _078125_);
  xor g_134419_(_075336_, _078124_, _078126_);
  not g_134420_(_078126_, _078127_);
  or g_134421_(_075340_, _078126_, _078128_);
  not g_134422_(_078128_, _078129_);
  or g_134423_(_075343_, _078126_, _078130_);
  xor g_134424_(_075343_, _078127_, _078132_);
  and g_134425_(_075340_, _078132_, _078133_);
  or g_134426_(_078129_, _078133_, _078134_);
  not g_134427_(_078134_, _078135_);
  or g_134428_(_075345_, _078134_, _078136_);
  xor g_134429_(_075345_, _078135_, _078137_);
  and g_134430_(_075348_, _078137_, _078138_);
  or g_134431_(_075348_, _078134_, _078139_);
  not g_134432_(_078139_, _078140_);
  or g_134433_(_078138_, _078140_, _078141_);
  and g_134434_(_075352_, _078141_, _078143_);
  not g_134435_(_078143_, _078144_);
  or g_134436_(_075352_, _078137_, _078145_);
  and g_134437_(_078144_, _078145_, _078146_);
  or g_134438_(_075355_, _078146_, _078147_);
  or g_134439_(_075354_, _078143_, _078148_);
  and g_134440_(_078147_, _078148_, out[961]);
  or g_134441_(_075330_, _078121_, _078149_);
  not g_134442_(_078149_, _078150_);
  or g_134443_(_075298_, _078094_, _078151_);
  or g_134444_(_075200_, _078008_, _078153_);
  not g_134445_(_078153_, _078154_);
  or g_134446_(_075197_, _078004_, _078155_);
  not g_134447_(_078155_, _078156_);
  and g_134448_(_075176_, _077983_, _078157_);
  not g_134449_(_078157_, _078158_);
  or g_134450_(_075166_, _077978_, _078159_);
  or g_134451_(_075163_, _077973_, _078160_);
  and g_134452_(_075131_, _077946_, _078161_);
  not g_134453_(_078161_, _078162_);
  or g_134454_(_075126_, _077945_, _078164_);
  and g_134455_(_075116_, _077939_, _078165_);
  not g_134456_(_078165_, _078166_);
  or g_134457_(_075112_, _077936_, _078167_);
  or g_134458_(_075092_, _077918_, _078168_);
  not g_134459_(_078168_, _078169_);
  or g_134460_(_075070_, _077895_, _078170_);
  or g_134461_(_075053_, _077881_, _078171_);
  not g_134462_(_078171_, _078172_);
  or g_134463_(_075049_, _077876_, _078173_);
  or g_134464_(_075035_, _077872_, _078175_);
  or g_134465_(_075029_, _077864_, _078176_);
  or g_134466_(_075003_, _077841_, _078177_);
  or g_134467_(_075000_, _077839_, _078178_);
  or g_134468_(_074993_, _077836_, _078179_);
  or g_134469_(_074978_, _077831_, _078180_);
  and g_134470_(_074974_, _077829_, _078181_);
  not g_134471_(_078181_, _078182_);
  or g_134472_(_074970_, _077827_, _078183_);
  and g_134473_(_077826_, _077828_, _078184_);
  or g_134474_(_074950_, _077809_, _078186_);
  not g_134475_(_078186_, _078187_);
  or g_134476_(_074930_, _077787_, _078188_);
  not g_134477_(_078188_, _078189_);
  or g_134478_(_074882_, _077737_, _078190_);
  or g_134479_(_074875_, _077726_, _078191_);
  or g_134480_(_074873_, _077726_, _078192_);
  or g_134481_(_074852_, _077697_, _078193_);
  or g_134482_(_074825_, _077674_, _078194_);
  or g_134483_(_074816_, _077668_, _078195_);
  and g_134484_(_074773_, _077612_, _078197_);
  or g_134485_(_074772_, _077613_, _078198_);
  or g_134486_(_074754_, _077593_, _078199_);
  or g_134487_(_074741_, _077582_, _078200_);
  or g_134488_(_074738_, _077582_, _078201_);
  not g_134489_(_078201_, _078202_);
  or g_134490_(_074729_, _077573_, _078203_);
  not g_134491_(_078203_, _078204_);
  or g_134492_(_074705_, _077554_, _078205_);
  or g_134493_(_074680_, _077528_, _078206_);
  or g_134494_(_074676_, _077523_, _078208_);
  not g_134495_(_078208_, _078209_);
  or g_134496_(_074665_, _077517_, _078210_);
  or g_134497_(_074663_, _077517_, _078211_);
  not g_134498_(_078211_, _078212_);
  or g_134499_(_074660_, _077516_, _078213_);
  or g_134500_(_074653_, _077512_, _078214_);
  or g_134501_(_074625_, _077477_, _078215_);
  or g_134502_(_074622_, _077473_, _078216_);
  not g_134503_(_078216_, _078217_);
  or g_134504_(_074576_, _077420_, _078219_);
  or g_134505_(_074566_, _077414_, _078220_);
  or g_134506_(_074559_, _077408_, _078221_);
  or g_134507_(_074553_, _077404_, _078222_);
  or g_134508_(_074550_, _077404_, _078223_);
  or g_134509_(_074538_, _077390_, _078224_);
  or g_134510_(_074534_, _077390_, _078225_);
  and g_134511_(_077388_, _078225_, _078226_);
  or g_134512_(_074521_, _077370_, _078227_);
  not g_134513_(_078227_, _078228_);
  or g_134514_(_074506_, _077360_, _078230_);
  and g_134515_(_074485_, _077336_, _078231_);
  not g_134516_(_078231_, _078232_);
  and g_134517_(_074481_, _077336_, _078233_);
  not g_134518_(_078233_, _078234_);
  or g_134519_(_074477_, _077334_, _078235_);
  or g_134520_(_074457_, _077318_, _078236_);
  not g_134521_(_078236_, _078237_);
  or g_134522_(_074388_, _077237_, _078238_);
  not g_134523_(_078238_, _078239_);
  or g_134524_(_074386_, _077237_, _078241_);
  and g_134525_(_074384_, _077235_, _078242_);
  or g_134526_(_074383_, _077236_, _078243_);
  or g_134527_(_074380_, _077236_, _078244_);
  or g_134528_(_074362_, _077219_, _078245_);
  or g_134529_(_074358_, _077214_, _078246_);
  or g_134530_(_074344_, _077203_, _078247_);
  or g_134531_(_074342_, _077203_, _078248_);
  or g_134532_(_074340_, _077200_, _078249_);
  or g_134533_(_074336_, _077200_, _078250_);
  not g_134534_(_078250_, _078252_);
  and g_134535_(_074333_, _077198_, _078253_);
  or g_134536_(_074332_, _077199_, _078254_);
  or g_134537_(_074324_, _077194_, _078255_);
  or g_134538_(_074292_, _077159_, _078256_);
  not g_134539_(_078256_, _078257_);
  or g_134540_(_074290_, _077159_, _078258_);
  or g_134541_(_074278_, _077149_, _078259_);
  or g_134542_(_074269_, _077143_, _078260_);
  or g_134543_(_074267_, _077139_, _078261_);
  or g_134544_(_074252_, _077127_, _078263_);
  not g_134545_(_078263_, _078264_);
  or g_134546_(_074220_, _077095_, _078265_);
  and g_134547_(_074182_, _077054_, _078266_);
  or g_134548_(_074181_, _077055_, _078267_);
  or g_134549_(_074179_, _077050_, _078268_);
  and g_134550_(_077049_, _077052_, _078269_);
  or g_134551_(_074159_, _077037_, _078270_);
  and g_134552_(_077021_, _077023_, _078271_);
  not g_134553_(_078271_, _078272_);
  or g_134554_(_074129_, _077002_, _078274_);
  or g_134555_(_074119_, _076996_, _078275_);
  or g_134556_(_074107_, _076988_, _078276_);
  or g_134557_(_074092_, _076968_, _078277_);
  and g_134558_(_074078_, _076955_, _078278_);
  or g_134559_(_074077_, _076956_, _078279_);
  or g_134560_(_074075_, _076956_, _078280_);
  and g_134561_(_076920_, _076925_, _078281_);
  and g_134562_(_076904_, _076908_, _078282_);
  or g_134563_(_074002_, _076884_, _078283_);
  and g_134564_(_073976_, _076864_, _078285_);
  not g_134565_(_078285_, _078286_);
  and g_134566_(_073972_, _076861_, _078287_);
  not g_134567_(_078287_, _078288_);
  or g_134568_(_073968_, _076859_, _078289_);
  and g_134569_(_073951_, _076842_, _078290_);
  or g_134570_(_073950_, _076843_, _078291_);
  or g_134571_(_073947_, _076839_, _078292_);
  or g_134572_(_073937_, _076834_, _078293_);
  not g_134573_(_078293_, _078294_);
  or g_134574_(_073934_, _076834_, _078296_);
  not g_134575_(_078296_, _078297_);
  and g_134576_(_076827_, _076832_, _078298_);
  or g_134577_(_073861_, _076746_, _078299_);
  or g_134578_(_073850_, _076735_, _078300_);
  or g_134579_(_073805_, _076695_, _078301_);
  or g_134580_(_073789_, _076682_, _078302_);
  or g_134581_(_073785_, _076682_, _078303_);
  not g_134582_(_078303_, _078304_);
  or g_134583_(_073768_, _076658_, _078305_);
  not g_134584_(_078305_, _078307_);
  or g_134585_(_073749_, _076642_, _078308_);
  not g_134586_(_078308_, _078309_);
  or g_134587_(_073728_, _076618_, _078310_);
  and g_134588_(_073725_, _076617_, _078311_);
  not g_134589_(_078311_, _078312_);
  and g_134590_(_073719_, _076614_, _078313_);
  not g_134591_(_078313_, _078314_);
  or g_134592_(_073716_, _076611_, _078315_);
  and g_134593_(_076610_, _076612_, _078316_);
  and g_134594_(_076586_, _076590_, _078318_);
  or g_134595_(_073643_, _076540_, _078319_);
  or g_134596_(_073624_, _076522_, _078320_);
  and g_134597_(_073613_, _076513_, _078321_);
  or g_134598_(_073612_, _076515_, _078322_);
  or g_134599_(_073608_, _076510_, _078323_);
  and g_134600_(_076476_, _076479_, _078324_);
  or g_134601_(_073553_, _076454_, _078325_);
  or g_134602_(_073544_, _076450_, _078326_);
  and g_134603_(_076418_, _076420_, _078327_);
  and g_134604_(_076412_, _076417_, _078329_);
  or g_134605_(_073452_, _076354_, _078330_);
  or g_134606_(_073450_, _076353_, _078331_);
  or g_134607_(_073447_, _076353_, _078332_);
  not g_134608_(_078332_, _078333_);
  or g_134609_(_073443_, _076347_, _078334_);
  not g_134610_(_078334_, _078335_);
  or g_134611_(_073441_, _076347_, _078336_);
  or g_134612_(_073429_, _076334_, _078337_);
  not g_134613_(_078337_, _078338_);
  or g_134614_(_073426_, _076334_, _078340_);
  and g_134615_(_073423_, _076332_, _078341_);
  not g_134616_(_078341_, _078342_);
  or g_134617_(_073401_, _076312_, _078343_);
  or g_134618_(_073385_, _076300_, _078344_);
  or g_134619_(_073382_, _076300_, _078345_);
  or g_134620_(_073378_, _076297_, _078346_);
  or g_134621_(_073375_, _076297_, _078347_);
  not g_134622_(_078347_, _078348_);
  or g_134623_(_073360_, _076280_, _078349_);
  or g_134624_(_073349_, _076276_, _078351_);
  or g_134625_(_073339_, _076269_, _078352_);
  not g_134626_(_078352_, _078353_);
  or g_134627_(_073335_, _076266_, _078354_);
  and g_134628_(_076263_, _076268_, _078355_);
  or g_134629_(_073319_, _076253_, _078356_);
  or g_134630_(_073313_, _076248_, _078357_);
  and g_134631_(_076196_, _076202_, _078358_);
  or g_134632_(_073252_, _076182_, _078359_);
  and g_134633_(_076169_, _076171_, _078360_);
  or g_134634_(_073188_, _076104_, _078362_);
  or g_134635_(_073185_, _076104_, _078363_);
  or g_134636_(_073165_, _076083_, _078364_);
  or g_134637_(_073162_, _076083_, _078365_);
  or g_134638_(_073156_, _076077_, _078366_);
  or g_134639_(_073154_, _076077_, _078367_);
  or g_134640_(_073152_, _076076_, _078368_);
  not g_134641_(_078368_, _078369_);
  or g_134642_(_073146_, _076075_, _078370_);
  or g_134643_(_073143_, _076075_, _078371_);
  or g_134644_(_073087_, _076005_, _078373_);
  or g_134645_(_073084_, _076002_, _078374_);
  or g_134646_(_073063_, _075981_, _078375_);
  not g_134647_(_078375_, _078376_);
  and g_134648_(_073059_, _075982_, _078377_);
  not g_134649_(_078377_, _078378_);
  or g_134650_(_073056_, _075979_, _078379_);
  or g_134651_(_073043_, _075967_, _078380_);
  or g_134652_(_073027_, _075959_, _078381_);
  or g_134653_(_073023_, _075948_, _078382_);
  or g_134654_(_072987_, _075921_, _078384_);
  or g_134655_(_075904_, _075912_, _078385_);
  or g_134656_(_072939_, _075862_, _078386_);
  or g_134657_(_072828_, _075760_, _078387_);
  or g_134658_(_072824_, _075752_, _078388_);
  and g_134659_(_075758_, _078388_, _078389_);
  and g_134660_(_075688_, _075691_, _078390_);
  or g_134661_(_072737_, _075658_, _078391_);
  and g_134662_(_075654_, _075659_, _078392_);
  or g_134663_(_072696_, _075613_, _078393_);
  and g_134664_(_075552_, _075555_, _078395_);
  not g_134665_(_078395_, _078396_);
  and g_134666_(_075544_, _075549_, _078397_);
  not g_134667_(_078397_, _078398_);
  or g_134668_(_072568_, _075478_, _078399_);
  or g_134669_(_072564_, _075478_, _078400_);
  or g_134670_(_072553_, _075474_, _078401_);
  or g_134671_(_072551_, _075474_, _078402_);
  or g_134672_(_072543_, _075472_, _078403_);
  or g_134673_(_072540_, _075472_, _078404_);
  and g_134674_(_075455_, _075457_, _078406_);
  and g_134675_(_075463_, _078406_, _078407_);
  or g_134676_(_075470_, _078407_, _078408_);
  xor g_134677_(_075468_, _078407_, _078409_);
  not g_134678_(_078409_, _078410_);
  or g_134679_(_075466_, _078409_, _078411_);
  xor g_134680_(_075466_, _078409_, _078412_);
  xor g_134681_(_075466_, _078410_, _078413_);
  or g_134682_(_072538_, _075471_, _078414_);
  or g_134683_(_072536_, _075471_, _078415_);
  or g_134684_(_078413_, _078415_, _078417_);
  xor g_134685_(_078412_, _078415_, _078418_);
  not g_134686_(_078418_, _078419_);
  or g_134687_(_078414_, _078418_, _078420_);
  xor g_134688_(_078414_, _078418_, _078421_);
  xor g_134689_(_078414_, _078419_, _078422_);
  or g_134690_(_078404_, _078422_, _078423_);
  xor g_134691_(_078404_, _078421_, _078424_);
  not g_134692_(_078424_, _078425_);
  or g_134693_(_078403_, _078424_, _078426_);
  xor g_134694_(_078403_, _078424_, _078428_);
  xor g_134695_(_078403_, _078425_, _078429_);
  or g_134696_(_072547_, _075473_, _078430_);
  or g_134697_(_078429_, _078430_, _078431_);
  xor g_134698_(_078428_, _078430_, _078432_);
  or g_134699_(_072549_, _075473_, _078433_);
  not g_134700_(_078433_, _078434_);
  or g_134701_(_078432_, _078433_, _078435_);
  xor g_134702_(_078432_, _078434_, _078436_);
  not g_134703_(_078436_, _078437_);
  or g_134704_(_078402_, _078436_, _078439_);
  xor g_134705_(_078402_, _078436_, _078440_);
  xor g_134706_(_078402_, _078437_, _078441_);
  or g_134707_(_078401_, _078441_, _078442_);
  xor g_134708_(_078401_, _078440_, _078443_);
  or g_134709_(_072556_, _075475_, _078444_);
  or g_134710_(_078443_, _078444_, _078445_);
  or g_134711_(_072561_, _075476_, _078446_);
  and g_134712_(_072557_, _075477_, _078447_);
  or g_134713_(_072556_, _075476_, _078448_);
  or g_134714_(_078443_, _078448_, _078450_);
  xor g_134715_(_078443_, _078447_, _078451_);
  not g_134716_(_078451_, _078452_);
  or g_134717_(_078446_, _078451_, _078453_);
  xor g_134718_(_078446_, _078452_, _078454_);
  not g_134719_(_078454_, _078455_);
  or g_134720_(_078400_, _078454_, _078456_);
  xor g_134721_(_078400_, _078455_, _078457_);
  not g_134722_(_078457_, _078458_);
  or g_134723_(_078399_, _078457_, _078459_);
  xor g_134724_(_078399_, _078458_, _078461_);
  or g_134725_(_072570_, _075481_, _078462_);
  not g_134726_(_078462_, _078463_);
  or g_134727_(_078461_, _078462_, _078464_);
  xor g_134728_(_078461_, _078463_, _078465_);
  or g_134729_(_072573_, _075481_, _078466_);
  not g_134730_(_078466_, _078467_);
  or g_134731_(_078465_, _078466_, _078468_);
  xor g_134732_(_078465_, _078466_, _078469_);
  xor g_134733_(_078465_, _078467_, _078470_);
  or g_134734_(_075487_, _078470_, _078472_);
  xor g_134735_(_075487_, _078469_, _078473_);
  not g_134736_(_078473_, _078474_);
  or g_134737_(_075485_, _078473_, _078475_);
  xor g_134738_(_075485_, _078474_, _078476_);
  or g_134739_(_072582_, _075488_, _078477_);
  or g_134740_(_072580_, _075488_, _078478_);
  not g_134741_(_078478_, _078479_);
  or g_134742_(_078476_, _078478_, _078480_);
  xor g_134743_(_078476_, _078479_, _078481_);
  not g_134744_(_078481_, _078483_);
  or g_134745_(_078477_, _078481_, _078484_);
  xor g_134746_(_078477_, _078483_, _078485_);
  or g_134747_(_075494_, _078485_, _078486_);
  xor g_134748_(_075495_, _078485_, _078487_);
  not g_134749_(_078487_, _078488_);
  or g_134750_(_075492_, _078487_, _078489_);
  xor g_134751_(_075492_, _078488_, _078490_);
  not g_134752_(_078490_, _078491_);
  or g_134753_(_075498_, _078490_, _078492_);
  xor g_134754_(_075498_, _078491_, _078494_);
  not g_134755_(_078494_, _078495_);
  or g_134756_(_075505_, _078494_, _078496_);
  not g_134757_(_078496_, _078497_);
  or g_134758_(_075501_, _078494_, _078498_);
  xor g_134759_(_075501_, _078495_, _078499_);
  and g_134760_(_075505_, _078499_, _078500_);
  or g_134761_(_078497_, _078500_, _078501_);
  and g_134762_(_075508_, _078501_, _078502_);
  or g_134763_(_075508_, _078499_, _078503_);
  not g_134764_(_078503_, _078505_);
  or g_134765_(_078502_, _078505_, _078506_);
  not g_134766_(_078506_, _078507_);
  or g_134767_(_075512_, _078506_, _078508_);
  xor g_134768_(_075512_, _078506_, _078509_);
  xor g_134769_(_075512_, _078507_, _078510_);
  or g_134770_(_075514_, _078510_, _078511_);
  xor g_134771_(_075514_, _078509_, _078512_);
  or g_134772_(_075520_, _078512_, _078513_);
  xor g_134773_(_075521_, _078512_, _078514_);
  not g_134774_(_078514_, _078516_);
  or g_134775_(_075522_, _078514_, _078517_);
  xor g_134776_(_075522_, _078516_, _078518_);
  or g_134777_(_072614_, _075518_, _078519_);
  not g_134778_(_078519_, _078520_);
  or g_134779_(_078518_, _078519_, _078521_);
  xor g_134780_(_078518_, _078520_, _078522_);
  not g_134781_(_078522_, _078523_);
  or g_134782_(_072617_, _075518_, _078524_);
  or g_134783_(_078522_, _078524_, _078525_);
  xor g_134784_(_078523_, _078524_, _078527_);
  not g_134785_(_078527_, _078528_);
  or g_134786_(_075530_, _078527_, _078529_);
  xor g_134787_(_075530_, _078527_, _078530_);
  xor g_134788_(_075530_, _078528_, _078531_);
  or g_134789_(_075531_, _078531_, _078532_);
  xor g_134790_(_075531_, _078530_, _078533_);
  not g_134791_(_078533_, _078534_);
  or g_134792_(_075532_, _078533_, _078535_);
  xor g_134793_(_075532_, _078534_, _078536_);
  or g_134794_(_075538_, _078536_, _078538_);
  xor g_134795_(_075539_, _078536_, _078539_);
  xor g_134796_(_078398_, _078539_, _078540_);
  xor g_134797_(_078395_, _078540_, _078541_);
  xor g_134798_(_078396_, _078540_, _078542_);
  or g_134799_(_075559_, _078542_, _078543_);
  xor g_134800_(_075559_, _078541_, _078544_);
  or g_134801_(_075562_, _078544_, _078545_);
  xor g_134802_(_075562_, _078544_, _078546_);
  not g_134803_(_078546_, _078547_);
  or g_134804_(_075563_, _078547_, _078549_);
  not g_134805_(_078549_, _078550_);
  xor g_134806_(_075563_, _078546_, _078551_);
  or g_134807_(_075567_, _078551_, _078552_);
  xor g_134808_(_075567_, _078551_, _078553_);
  not g_134809_(_078553_, _078554_);
  or g_134810_(_075573_, _078554_, _078555_);
  xor g_134811_(_075573_, _078553_, _078556_);
  not g_134812_(_078556_, _078557_);
  and g_134813_(_075580_, _075586_, _078558_);
  xor g_134814_(_078556_, _078558_, _078560_);
  xor g_134815_(_078557_, _078558_, _078561_);
  or g_134816_(_075587_, _078561_, _078562_);
  not g_134817_(_078562_, _078563_);
  xor g_134818_(_075587_, _078560_, _078564_);
  not g_134819_(_078564_, _078565_);
  or g_134820_(_075595_, _078564_, _078566_);
  xor g_134821_(_075595_, _078565_, _078567_);
  or g_134822_(_075599_, _078567_, _078568_);
  xor g_134823_(_075598_, _078567_, _078569_);
  or g_134824_(_075605_, _078569_, _078571_);
  xor g_134825_(_075605_, _078569_, _078572_);
  not g_134826_(_078572_, _078573_);
  and g_134827_(_075604_, _078572_, _078574_);
  or g_134828_(_075603_, _078573_, _078575_);
  xor g_134829_(_075603_, _078572_, _078576_);
  or g_134830_(_075610_, _078576_, _078577_);
  xor g_134831_(_075611_, _078576_, _078578_);
  or g_134832_(_072693_, _075608_, _078579_);
  not g_134833_(_078579_, _078580_);
  or g_134834_(_078578_, _078579_, _078582_);
  xor g_134835_(_078578_, _078579_, _078583_);
  xor g_134836_(_078578_, _078580_, _078584_);
  or g_134837_(_078393_, _078584_, _078585_);
  xor g_134838_(_078393_, _078583_, _078586_);
  not g_134839_(_078586_, _078587_);
  or g_134840_(_075618_, _078586_, _078588_);
  xor g_134841_(_075618_, _078586_, _078589_);
  xor g_134842_(_075618_, _078587_, _078590_);
  or g_134843_(_075619_, _078590_, _078591_);
  xor g_134844_(_075619_, _078589_, _078593_);
  not g_134845_(_078593_, _078594_);
  and g_134846_(_075622_, _075625_, _078595_);
  xor g_134847_(_078594_, _078595_, _078596_);
  not g_134848_(_078596_, _078597_);
  and g_134849_(_075633_, _078597_, _078598_);
  not g_134850_(_078598_, _078599_);
  and g_134851_(_075629_, _078597_, _078600_);
  not g_134852_(_078600_, _078601_);
  or g_134853_(_078598_, _078600_, _078602_);
  and g_134854_(_075628_, _078596_, _078604_);
  and g_134855_(_075632_, _078604_, _078605_);
  or g_134856_(_078602_, _078605_, _078606_);
  or g_134857_(_075636_, _078606_, _078607_);
  not g_134858_(_078607_, _078608_);
  xor g_134859_(_075636_, _078606_, _078609_);
  not g_134860_(_078609_, _078610_);
  or g_134861_(_072719_, _075635_, _078611_);
  or g_134862_(_078610_, _078611_, _078612_);
  not g_134863_(_078612_, _078613_);
  xor g_134864_(_078609_, _078611_, _078615_);
  not g_134865_(_078615_, _078616_);
  or g_134866_(_072723_, _075638_, _078617_);
  and g_134867_(_075642_, _078617_, _078618_);
  and g_134868_(_075648_, _078618_, _078619_);
  xor g_134869_(_078616_, _078619_, _078620_);
  not g_134870_(_078620_, _078621_);
  xor g_134871_(_078392_, _078621_, _078622_);
  not g_134872_(_078622_, _078623_);
  or g_134873_(_078391_, _078622_, _078624_);
  xor g_134874_(_078391_, _078622_, _078626_);
  xor g_134875_(_078391_, _078623_, _078627_);
  or g_134876_(_072740_, _075660_, _078628_);
  or g_134877_(_078627_, _078628_, _078629_);
  xor g_134878_(_078626_, _078628_, _078630_);
  and g_134879_(_075664_, _078630_, _078631_);
  or g_134880_(_075664_, _078630_, _078632_);
  not g_134881_(_078632_, _078633_);
  xor g_134882_(_075664_, _078630_, _078634_);
  or g_134883_(_078631_, _078633_, _078635_);
  or g_134884_(_072747_, _075663_, _078637_);
  or g_134885_(_078635_, _078637_, _078638_);
  xor g_134886_(_078634_, _078637_, _078639_);
  or g_134887_(_072749_, _075665_, _078640_);
  not g_134888_(_078640_, _078641_);
  or g_134889_(_078639_, _078640_, _078642_);
  xor g_134890_(_078639_, _078641_, _078643_);
  not g_134891_(_078643_, _078644_);
  and g_134892_(_075671_, _075674_, _078645_);
  xor g_134893_(_078644_, _078645_, _078646_);
  or g_134894_(_075679_, _078646_, _078648_);
  xor g_134895_(_075679_, _078646_, _078649_);
  not g_134896_(_078649_, _078650_);
  or g_134897_(_075680_, _078650_, _078651_);
  not g_134898_(_078651_, _078652_);
  xor g_134899_(_075680_, _078649_, _078653_);
  not g_134900_(_078653_, _078654_);
  and g_134901_(_075684_, _075686_, _078655_);
  xor g_134902_(_078654_, _078655_, _078656_);
  not g_134903_(_078656_, _078657_);
  xor g_134904_(_078390_, _078657_, _078659_);
  or g_134905_(_075695_, _078659_, _078660_);
  not g_134906_(_078660_, _078661_);
  xor g_134907_(_075695_, _078659_, _078662_);
  not g_134908_(_078662_, _078663_);
  and g_134909_(_075699_, _078662_, _078664_);
  not g_134910_(_078664_, _078665_);
  or g_134911_(_075703_, _078663_, _078666_);
  not g_134912_(_078666_, _078667_);
  xor g_134913_(_075703_, _078662_, _078668_);
  and g_134914_(_075701_, _078668_, _078670_);
  or g_134915_(_078664_, _078670_, _078671_);
  or g_134916_(_075707_, _075714_, _078672_);
  xor g_134917_(_078671_, _078672_, _078673_);
  not g_134918_(_078673_, _078674_);
  and g_134919_(_075709_, _075720_, _078675_);
  xor g_134920_(_078674_, _078675_, _078676_);
  or g_134921_(_075724_, _078676_, _078677_);
  not g_134922_(_078677_, _078678_);
  xor g_134923_(_075724_, _078676_, _078679_);
  not g_134924_(_078679_, _078681_);
  and g_134925_(_075730_, _078679_, _078682_);
  or g_134926_(_075729_, _078681_, _078683_);
  xor g_134927_(_075729_, _078679_, _078684_);
  or g_134928_(_075738_, _078684_, _078685_);
  xor g_134929_(_075739_, _078684_, _078686_);
  or g_134930_(_075734_, _078686_, _078687_);
  xor g_134931_(_075735_, _078686_, _078688_);
  or g_134932_(_072821_, _075752_, _078689_);
  and g_134933_(_075749_, _078689_, _078690_);
  xor g_134934_(_078688_, _078690_, _078692_);
  not g_134935_(_078692_, _078693_);
  xor g_134936_(_078389_, _078692_, _078694_);
  and g_134937_(_078387_, _078694_, _078695_);
  or g_134938_(_078387_, _078694_, _078696_);
  not g_134939_(_078696_, _078697_);
  xor g_134940_(_078387_, _078694_, _078698_);
  or g_134941_(_078695_, _078697_, _078699_);
  or g_134942_(_072832_, _075760_, _078700_);
  or g_134943_(_078699_, _078700_, _078701_);
  not g_134944_(_078701_, _078703_);
  xor g_134945_(_078698_, _078700_, _078704_);
  not g_134946_(_078704_, _078705_);
  and g_134947_(_075768_, _075772_, _078706_);
  and g_134948_(_075775_, _078706_, _078707_);
  xor g_134949_(_078705_, _078707_, _078708_);
  or g_134950_(_072848_, _075773_, _078709_);
  not g_134951_(_078709_, _078710_);
  or g_134952_(_078708_, _078709_, _078711_);
  xor g_134953_(_078708_, _078710_, _078712_);
  or g_134954_(_072850_, _075778_, _078714_);
  or g_134955_(_078712_, _078714_, _078715_);
  not g_134956_(_078715_, _078716_);
  and g_134957_(_078712_, _078714_, _078717_);
  xor g_134958_(_078712_, _078714_, _078718_);
  or g_134959_(_078716_, _078717_, _078719_);
  and g_134960_(_075783_, _075785_, _078720_);
  xor g_134961_(_078718_, _078720_, _078721_);
  or g_134962_(_075789_, _078721_, _078722_);
  xor g_134963_(_075789_, _078721_, _078723_);
  not g_134964_(_078723_, _078725_);
  and g_134965_(_075791_, _078723_, _078726_);
  or g_134966_(_075790_, _078725_, _078727_);
  xor g_134967_(_075790_, _078723_, _078728_);
  not g_134968_(_078728_, _078729_);
  or g_134969_(_075793_, _078728_, _078730_);
  xor g_134970_(_075793_, _078728_, _078731_);
  xor g_134971_(_075793_, _078729_, _078732_);
  or g_134972_(_075797_, _078732_, _078733_);
  xor g_134973_(_075797_, _078731_, _078734_);
  or g_134974_(_072876_, _075795_, _078736_);
  and g_134975_(_078734_, _078736_, _078737_);
  or g_134976_(_078734_, _078736_, _078738_);
  not g_134977_(_078738_, _078739_);
  xor g_134978_(_078734_, _078736_, _078740_);
  or g_134979_(_078737_, _078739_, _078741_);
  or g_134980_(_075805_, _078741_, _078742_);
  or g_134981_(_068025_, _078742_, _078743_);
  or g_134982_(_075804_, _078740_, _078744_);
  and g_134983_(_078743_, _078744_, _078745_);
  not g_134984_(_078745_, _078747_);
  or g_134985_(_075812_, _078747_, _078748_);
  xor g_134986_(_075812_, _078745_, _078749_);
  or g_134987_(_075809_, _078749_, _078750_);
  xor g_134988_(_075808_, _078749_, _078751_);
  or g_134989_(_075818_, _078751_, _078752_);
  xor g_134990_(_075819_, _078751_, _078753_);
  not g_134991_(_078753_, _078754_);
  and g_134992_(_075825_, _075828_, _078755_);
  xor g_134993_(_078754_, _078755_, _078756_);
  or g_134994_(_075833_, _078756_, _078758_);
  xor g_134995_(_075831_, _078756_, _078759_);
  or g_134996_(_075838_, _078759_, _078760_);
  xor g_134997_(_075839_, _078759_, _078761_);
  or g_134998_(_075835_, _078761_, _078762_);
  not g_134999_(_078762_, _078763_);
  xor g_135000_(_075836_, _078761_, _078764_);
  not g_135001_(_078764_, _078765_);
  or g_135002_(_075844_, _078764_, _078766_);
  xor g_135003_(_075844_, _078765_, _078767_);
  and g_135004_(_075849_, _078767_, _078769_);
  or g_135005_(_075849_, _078767_, _078770_);
  not g_135006_(_078770_, _078771_);
  or g_135007_(_078769_, _078771_, _078772_);
  not g_135008_(_078772_, _078773_);
  or g_135009_(_075848_, _078772_, _078774_);
  xor g_135010_(_075848_, _078773_, _078775_);
  not g_135011_(_078775_, _078776_);
  and g_135012_(_075853_, _075857_, _078777_);
  xor g_135013_(_078776_, _078777_, _078778_);
  or g_135014_(_075861_, _078778_, _078780_);
  xor g_135015_(_075860_, _078778_, _078781_);
  or g_135016_(_072936_, _075858_, _078782_);
  or g_135017_(_078781_, _078782_, _078783_);
  xor g_135018_(_078781_, _078782_, _078784_);
  not g_135019_(_078784_, _078785_);
  or g_135020_(_078386_, _078785_, _078786_);
  xor g_135021_(_078386_, _078784_, _078787_);
  not g_135022_(_078787_, _078788_);
  or g_135023_(_075870_, _078787_, _078789_);
  xor g_135024_(_075870_, _078788_, _078791_);
  or g_135025_(_075869_, _078791_, _078792_);
  not g_135026_(_078792_, _078793_);
  and g_135027_(_075869_, _078791_, _078794_);
  xor g_135028_(_075869_, _078791_, _078795_);
  or g_135029_(_078793_, _078794_, _078796_);
  and g_135030_(_075874_, _075879_, _078797_);
  and g_135031_(_078796_, _078797_, _078798_);
  and g_135032_(_075878_, _078795_, _078799_);
  or g_135033_(_075879_, _078796_, _078800_);
  and g_135034_(_075873_, _078795_, _078802_);
  or g_135035_(_075874_, _078796_, _078803_);
  or g_135036_(_078799_, _078802_, _078804_);
  or g_135037_(_078798_, _078804_, _078805_);
  or g_135038_(_075884_, _078805_, _078806_);
  xor g_135039_(_075885_, _078805_, _078807_);
  or g_135040_(_075881_, _078807_, _078808_);
  not g_135041_(_078808_, _078809_);
  xor g_135042_(_075882_, _078807_, _078810_);
  or g_135043_(_075891_, _078810_, _078811_);
  not g_135044_(_078811_, _078813_);
  or g_135045_(_075896_, _078810_, _078814_);
  not g_135046_(_078814_, _078815_);
  and g_135047_(_075896_, _078810_, _078816_);
  or g_135048_(_078815_, _078816_, _078817_);
  and g_135049_(_075891_, _078817_, _078818_);
  or g_135050_(_078813_, _078818_, _078819_);
  xor g_135051_(_075895_, _078819_, _078820_);
  xor g_135052_(_078385_, _078820_, _078821_);
  or g_135053_(_075908_, _078821_, _078822_);
  not g_135054_(_078822_, _078824_);
  xor g_135055_(_075907_, _078821_, _078825_);
  or g_135056_(_075919_, _078825_, _078826_);
  xor g_135057_(_075918_, _078825_, _078827_);
  or g_135058_(_072983_, _075916_, _078828_);
  not g_135059_(_078828_, _078829_);
  or g_135060_(_078827_, _078828_, _078830_);
  xor g_135061_(_078827_, _078828_, _078831_);
  xor g_135062_(_078827_, _078829_, _078832_);
  or g_135063_(_078384_, _078832_, _078833_);
  xor g_135064_(_078384_, _078831_, _078835_);
  not g_135065_(_078835_, _078836_);
  and g_135066_(_075927_, _075930_, _078837_);
  xor g_135067_(_078836_, _078837_, _078838_);
  and g_135068_(_075934_, _078838_, _078839_);
  or g_135069_(_075934_, _078838_, _078840_);
  not g_135070_(_078840_, _078841_);
  xor g_135071_(_075934_, _078838_, _078842_);
  or g_135072_(_078839_, _078841_, _078843_);
  or g_135073_(_073002_, _075933_, _078844_);
  or g_135074_(_078843_, _078844_, _078846_);
  not g_135075_(_078846_, _078847_);
  xor g_135076_(_078842_, _078844_, _078848_);
  or g_135077_(_073005_, _075935_, _078849_);
  or g_135078_(_078848_, _078849_, _078850_);
  xor g_135079_(_078848_, _078849_, _078851_);
  not g_135080_(_078851_, _078852_);
  or g_135081_(_075939_, _078852_, _078853_);
  xor g_135082_(_075939_, _078851_, _078854_);
  or g_135083_(_075941_, _078854_, _078855_);
  not g_135084_(_078855_, _078857_);
  and g_135085_(_075941_, _078854_, _078858_);
  or g_135086_(_078857_, _078858_, _078859_);
  and g_135087_(_075947_, _075955_, _078860_);
  xor g_135088_(_078859_, _078860_, _078861_);
  not g_135089_(_078861_, _078862_);
  or g_135090_(_078382_, _078862_, _078863_);
  not g_135091_(_078863_, _078864_);
  xor g_135092_(_078382_, _078861_, _078865_);
  not g_135093_(_078865_, _078866_);
  or g_135094_(_078381_, _078865_, _078868_);
  xor g_135095_(_078381_, _078866_, _078869_);
  not g_135096_(_078869_, _078870_);
  or g_135097_(_073040_, _075967_, _078871_);
  and g_135098_(_075966_, _078871_, _078872_);
  xor g_135099_(_078870_, _078872_, _078873_);
  xor g_135100_(_078869_, _078872_, _078874_);
  or g_135101_(_078380_, _078873_, _078875_);
  not g_135102_(_078875_, _078876_);
  xor g_135103_(_078380_, _078874_, _078877_);
  not g_135104_(_078877_, _078879_);
  and g_135105_(_075970_, _075973_, _078880_);
  or g_135106_(_078877_, _078880_, _078881_);
  xor g_135107_(_078877_, _078880_, _078882_);
  xor g_135108_(_078879_, _078880_, _078883_);
  or g_135109_(_075977_, _078883_, _078884_);
  xor g_135110_(_075977_, _078882_, _078885_);
  or g_135111_(_073054_, _075974_, _078886_);
  not g_135112_(_078886_, _078887_);
  or g_135113_(_078885_, _078886_, _078888_);
  not g_135114_(_078888_, _078890_);
  xor g_135115_(_078885_, _078887_, _078891_);
  or g_135116_(_078379_, _078891_, _078892_);
  not g_135117_(_078892_, _078893_);
  and g_135118_(_078379_, _078891_, _078894_);
  or g_135119_(_078893_, _078894_, _078895_);
  or g_135120_(_078378_, _078895_, _078896_);
  not g_135121_(_078896_, _078897_);
  xor g_135122_(_078377_, _078895_, _078898_);
  or g_135123_(_078375_, _078898_, _078899_);
  xor g_135124_(_078376_, _078898_, _078901_);
  or g_135125_(_075984_, _078901_, _078902_);
  xor g_135126_(_075985_, _078901_, _078903_);
  xor g_135127_(_075993_, _078903_, _078904_);
  or g_135128_(_075996_, _078904_, _078905_);
  xor g_135129_(_075996_, _078904_, _078906_);
  not g_135130_(_078906_, _078907_);
  or g_135131_(_076000_, _078907_, _078908_);
  not g_135132_(_078908_, _078909_);
  xor g_135133_(_076000_, _078906_, _078910_);
  not g_135134_(_078910_, _078912_);
  or g_135135_(_073081_, _075998_, _078913_);
  or g_135136_(_078910_, _078913_, _078914_);
  xor g_135137_(_078910_, _078913_, _078915_);
  xor g_135138_(_078912_, _078913_, _078916_);
  or g_135139_(_078374_, _078916_, _078917_);
  not g_135140_(_078917_, _078918_);
  xor g_135141_(_078374_, _078915_, _078919_);
  and g_135142_(_078373_, _078919_, _078920_);
  or g_135143_(_078373_, _078919_, _078921_);
  not g_135144_(_078921_, _078923_);
  or g_135145_(_078920_, _078923_, _078924_);
  or g_135146_(_073090_, _076005_, _078925_);
  not g_135147_(_078925_, _078926_);
  or g_135148_(_078924_, _078925_, _078927_);
  xor g_135149_(_078924_, _078925_, _078928_);
  xor g_135150_(_078924_, _078926_, _078929_);
  or g_135151_(_076007_, _078929_, _078930_);
  xor g_135152_(_076007_, _078928_, _078931_);
  not g_135153_(_078931_, _078932_);
  and g_135154_(_076011_, _076015_, _078934_);
  xor g_135155_(_078931_, _078934_, _078935_);
  xor g_135156_(_078932_, _078934_, _078936_);
  and g_135157_(_076020_, _078935_, _078937_);
  or g_135158_(_076018_, _078936_, _078938_);
  xor g_135159_(_076018_, _078935_, _078939_);
  or g_135160_(_076025_, _078939_, _078940_);
  xor g_135161_(_076024_, _078939_, _078941_);
  or g_135162_(_076032_, _078941_, _078942_);
  xor g_135163_(_076033_, _078941_, _078943_);
  or g_135164_(_076029_, _078943_, _078945_);
  not g_135165_(_078945_, _078946_);
  xor g_135166_(_076028_, _078943_, _078947_);
  not g_135167_(_078947_, _078948_);
  and g_135168_(_076039_, _078948_, _078949_);
  xor g_135169_(_076039_, _078947_, _078950_);
  or g_135170_(_076046_, _078950_, _078951_);
  not g_135171_(_078951_, _078952_);
  xor g_135172_(_076047_, _078950_, _078953_);
  or g_135173_(_076043_, _078953_, _078954_);
  not g_135174_(_078954_, _078956_);
  xor g_135175_(_076044_, _078953_, _078957_);
  or g_135176_(_076053_, _078957_, _078958_);
  xor g_135177_(_076054_, _078957_, _078959_);
  not g_135178_(_078959_, _078960_);
  or g_135179_(_076066_, _078959_, _078961_);
  xor g_135180_(_076066_, _078960_, _078962_);
  or g_135181_(_076057_, _078962_, _078963_);
  not g_135182_(_078963_, _078964_);
  xor g_135183_(_076057_, _078962_, _078965_);
  not g_135184_(_078965_, _078967_);
  xor g_135185_(_076070_, _078965_, _078968_);
  or g_135186_(_078371_, _078968_, _078969_);
  xor g_135187_(_078371_, _078968_, _078970_);
  not g_135188_(_078970_, _078971_);
  or g_135189_(_078370_, _078971_, _078972_);
  xor g_135190_(_078370_, _078970_, _078973_);
  or g_135191_(_073148_, _076076_, _078974_);
  not g_135192_(_078974_, _078975_);
  or g_135193_(_078973_, _078974_, _078976_);
  xor g_135194_(_078973_, _078975_, _078978_);
  or g_135195_(_078368_, _078978_, _078979_);
  xor g_135196_(_078369_, _078978_, _078980_);
  not g_135197_(_078980_, _078981_);
  or g_135198_(_078367_, _078980_, _078982_);
  xor g_135199_(_078367_, _078981_, _078983_);
  not g_135200_(_078983_, _078984_);
  or g_135201_(_078366_, _078983_, _078985_);
  not g_135202_(_078985_, _078986_);
  xor g_135203_(_078366_, _078984_, _078987_);
  or g_135204_(_076081_, _078987_, _078989_);
  xor g_135205_(_076082_, _078987_, _078990_);
  and g_135206_(_078365_, _078990_, _078991_);
  or g_135207_(_078365_, _078990_, _078992_);
  not g_135208_(_078992_, _078993_);
  xor g_135209_(_078365_, _078990_, _078994_);
  or g_135210_(_078991_, _078993_, _078995_);
  or g_135211_(_078364_, _078995_, _078996_);
  xor g_135212_(_078364_, _078994_, _078997_);
  or g_135213_(_076089_, _078997_, _078998_);
  not g_135214_(_078998_, _079000_);
  xor g_135215_(_076089_, _078997_, _079001_);
  not g_135216_(_079001_, _079002_);
  or g_135217_(_076093_, _079002_, _079003_);
  not g_135218_(_079003_, _079004_);
  xor g_135219_(_076093_, _079001_, _079005_);
  not g_135220_(_079005_, _079006_);
  or g_135221_(_076097_, _079005_, _079007_);
  xor g_135222_(_076097_, _079006_, _079008_);
  or g_135223_(_076102_, _079008_, _079009_);
  xor g_135224_(_076102_, _079008_, _079011_);
  xor g_135225_(_076103_, _079011_, _079012_);
  or g_135226_(_078363_, _079012_, _079013_);
  xor g_135227_(_078363_, _079012_, _079014_);
  not g_135228_(_079014_, _079015_);
  or g_135229_(_078362_, _079015_, _079016_);
  xor g_135230_(_078362_, _079014_, _079017_);
  or g_135231_(_076110_, _079017_, _079018_);
  not g_135232_(_079018_, _079019_);
  xor g_135233_(_076110_, _079017_, _079020_);
  not g_135234_(_079020_, _079022_);
  or g_135235_(_073194_, _076109_, _079023_);
  not g_135236_(_079023_, _079024_);
  and g_135237_(_079020_, _079024_, _079025_);
  or g_135238_(_079022_, _079023_, _079026_);
  xor g_135239_(_079020_, _079023_, _079027_);
  not g_135240_(_079027_, _079028_);
  and g_135241_(_076119_, _079028_, _079029_);
  or g_135242_(_076117_, _079027_, _079030_);
  xor g_135243_(_076119_, _079027_, _079031_);
  not g_135244_(_079031_, _079033_);
  xor g_135245_(_076137_, _079033_, _079034_);
  xor g_135246_(_076137_, _079031_, _079035_);
  or g_135247_(_076135_, _079034_, _079036_);
  xor g_135248_(_076135_, _079035_, _079037_);
  or g_135249_(_076142_, _079037_, _079038_);
  xor g_135250_(_076141_, _079037_, _079039_);
  or g_135251_(_076149_, _079039_, _079040_);
  xor g_135252_(_076150_, _079039_, _079041_);
  or g_135253_(_076146_, _079041_, _079042_);
  xor g_135254_(_076145_, _079041_, _079044_);
  and g_135255_(_076157_, _076167_, _079045_);
  and g_135256_(_076160_, _079045_, _079046_);
  xor g_135257_(_079044_, _079046_, _079047_);
  not g_135258_(_079047_, _079048_);
  xor g_135259_(_078360_, _079047_, _079049_);
  or g_135260_(_076179_, _079049_, _079050_);
  xor g_135261_(_076180_, _079049_, _079051_);
  or g_135262_(_073249_, _076177_, _079052_);
  or g_135263_(_079051_, _079052_, _079053_);
  xor g_135264_(_079051_, _079052_, _079055_);
  not g_135265_(_079055_, _079056_);
  or g_135266_(_078359_, _079056_, _079057_);
  xor g_135267_(_078359_, _079055_, _079058_);
  not g_135268_(_079058_, _079059_);
  and g_135269_(_076187_, _076190_, _079060_);
  xor g_135270_(_079059_, _079060_, _079061_);
  not g_135271_(_079061_, _079062_);
  xor g_135272_(_078358_, _079061_, _079063_);
  not g_135273_(_079063_, _079064_);
  and g_135274_(_076200_, _079063_, _079066_);
  or g_135275_(_076201_, _079064_, _079067_);
  xor g_135276_(_076200_, _079063_, _079068_);
  not g_135277_(_079068_, _079069_);
  and g_135278_(_076207_, _079068_, _079070_);
  or g_135279_(_076205_, _079069_, _079071_);
  xor g_135280_(_076205_, _079068_, _079072_);
  not g_135281_(_079072_, _079073_);
  and g_135282_(_076213_, _079073_, _079074_);
  not g_135283_(_079074_, _079075_);
  xor g_135284_(_076213_, _079072_, _079077_);
  and g_135285_(_076220_, _079077_, _079078_);
  not g_135286_(_079078_, _079079_);
  or g_135287_(_076218_, _079072_, _079080_);
  not g_135288_(_079080_, _079081_);
  or g_135289_(_076219_, _079077_, _079082_);
  and g_135290_(_079080_, _079082_, _079083_);
  not g_135291_(_079083_, _079084_);
  and g_135292_(_079079_, _079083_, _079085_);
  or g_135293_(_079078_, _079084_, _079086_);
  or g_135294_(_076223_, _079086_, _079088_);
  xor g_135295_(_076223_, _079085_, _079089_);
  or g_135296_(_076229_, _079089_, _079090_);
  xor g_135297_(_076227_, _079089_, _079091_);
  or g_135298_(_073296_, _076225_, _079092_);
  and g_135299_(_079091_, _079092_, _079093_);
  or g_135300_(_079091_, _079092_, _079094_);
  not g_135301_(_079094_, _079095_);
  or g_135302_(_079093_, _079095_, _079096_);
  or g_135303_(_076233_, _079096_, _079097_);
  not g_135304_(_079097_, _079099_);
  xor g_135305_(_076232_, _079096_, _079100_);
  xor g_135306_(_076243_, _079100_, _079101_);
  and g_135307_(_076247_, _079101_, _079102_);
  and g_135308_(_076251_, _079102_, _079103_);
  or g_135309_(_076251_, _079101_, _079104_);
  or g_135310_(_076247_, _079101_, _079105_);
  not g_135311_(_079105_, _079106_);
  and g_135312_(_079104_, _079105_, _079107_);
  not g_135313_(_079107_, _079108_);
  or g_135314_(_079103_, _079108_, _079110_);
  not g_135315_(_079110_, _079111_);
  or g_135316_(_078357_, _079110_, _079112_);
  xor g_135317_(_078357_, _079111_, _079113_);
  not g_135318_(_079113_, _079114_);
  or g_135319_(_078356_, _079113_, _079115_);
  xor g_135320_(_078356_, _079113_, _079116_);
  xor g_135321_(_078356_, _079114_, _079117_);
  and g_135322_(_076258_, _076260_, _079118_);
  xor g_135323_(_079116_, _079118_, _079119_);
  xor g_135324_(_078355_, _079119_, _079121_);
  not g_135325_(_079121_, _079122_);
  or g_135326_(_078354_, _079122_, _079123_);
  xor g_135327_(_078354_, _079121_, _079124_);
  or g_135328_(_078352_, _079124_, _079125_);
  xor g_135329_(_078353_, _079124_, _079126_);
  or g_135330_(_076274_, _079126_, _079127_);
  not g_135331_(_079127_, _079128_);
  xor g_135332_(_076275_, _079126_, _079129_);
  or g_135333_(_073344_, _076273_, _079130_);
  and g_135334_(_079129_, _079130_, _079132_);
  or g_135335_(_079129_, _079130_, _079133_);
  not g_135336_(_079133_, _079134_);
  xor g_135337_(_079129_, _079130_, _079135_);
  or g_135338_(_079132_, _079134_, _079136_);
  or g_135339_(_078351_, _079136_, _079137_);
  not g_135340_(_079137_, _079138_);
  xor g_135341_(_078351_, _079135_, _079139_);
  or g_135342_(_076278_, _079139_, _079140_);
  xor g_135343_(_076279_, _079139_, _079141_);
  not g_135344_(_079141_, _079143_);
  or g_135345_(_073357_, _076277_, _079144_);
  or g_135346_(_079141_, _079144_, _079145_);
  xor g_135347_(_079141_, _079144_, _079146_);
  xor g_135348_(_079143_, _079144_, _079147_);
  or g_135349_(_078349_, _079147_, _079148_);
  xor g_135350_(_078349_, _079146_, _079149_);
  or g_135351_(_076291_, _079149_, _079150_);
  not g_135352_(_079150_, _079151_);
  xor g_135353_(_076290_, _079149_, _079152_);
  or g_135354_(_076285_, _079152_, _079154_);
  xor g_135355_(_076285_, _079152_, _079155_);
  xor g_135356_(_076286_, _079152_, _079156_);
  or g_135357_(_076295_, _079155_, _079157_);
  or g_135358_(_078348_, _079157_, _079158_);
  or g_135359_(_076296_, _079156_, _079159_);
  not g_135360_(_079159_, _079160_);
  or g_135361_(_078347_, _079156_, _079161_);
  and g_135362_(_079159_, _079161_, _079162_);
  and g_135363_(_079158_, _079162_, _079163_);
  not g_135364_(_079163_, _079165_);
  or g_135365_(_078346_, _079165_, _079166_);
  xor g_135366_(_078346_, _079163_, _079167_);
  not g_135367_(_079167_, _079168_);
  or g_135368_(_078345_, _079167_, _079169_);
  xor g_135369_(_078345_, _079167_, _079170_);
  xor g_135370_(_078345_, _079168_, _079171_);
  or g_135371_(_078344_, _079171_, _079172_);
  not g_135372_(_079172_, _079173_);
  xor g_135373_(_078344_, _079170_, _079174_);
  or g_135374_(_076303_, _079174_, _079176_);
  xor g_135375_(_076303_, _079174_, _079177_);
  xor g_135376_(_076304_, _079174_, _079178_);
  or g_135377_(_076307_, _079178_, _079179_);
  xor g_135378_(_076307_, _079177_, _079180_);
  and g_135379_(_076310_, _079180_, _079181_);
  or g_135380_(_076310_, _079174_, _079182_);
  not g_135381_(_079182_, _079183_);
  or g_135382_(_079181_, _079183_, _079184_);
  or g_135383_(_073398_, _076308_, _079185_);
  not g_135384_(_079185_, _079187_);
  or g_135385_(_079184_, _079185_, _079188_);
  xor g_135386_(_079184_, _079185_, _079189_);
  xor g_135387_(_079184_, _079187_, _079190_);
  or g_135388_(_078343_, _079190_, _079191_);
  xor g_135389_(_078343_, _079189_, _079192_);
  or g_135390_(_076318_, _079192_, _079193_);
  xor g_135391_(_076318_, _079192_, _079194_);
  xor g_135392_(_076317_, _079192_, _079195_);
  or g_135393_(_076319_, _079195_, _079196_);
  xor g_135394_(_076319_, _079194_, _079198_);
  or g_135395_(_076323_, _079198_, _079199_);
  xor g_135396_(_076324_, _079198_, _079200_);
  or g_135397_(_076330_, _079200_, _079201_);
  not g_135398_(_079201_, _079202_);
  xor g_135399_(_076330_, _079200_, _079203_);
  xor g_135400_(_076331_, _079200_, _079204_);
  or g_135401_(_073419_, _076328_, _079205_);
  or g_135402_(_079204_, _079205_, _079206_);
  xor g_135403_(_079203_, _079205_, _079207_);
  or g_135404_(_078342_, _079207_, _079209_);
  xor g_135405_(_078342_, _079207_, _079210_);
  xor g_135406_(_078341_, _079207_, _079211_);
  or g_135407_(_078340_, _079211_, _079212_);
  xor g_135408_(_078340_, _079210_, _079213_);
  or g_135409_(_078337_, _079213_, _079214_);
  xor g_135410_(_078338_, _079213_, _079215_);
  and g_135411_(_076337_, _076341_, _079216_);
  not g_135412_(_079216_, _079217_);
  xor g_135413_(_079215_, _079217_, _079218_);
  or g_135414_(_076343_, _079218_, _079220_);
  xor g_135415_(_076343_, _079218_, _079221_);
  xor g_135416_(_076344_, _079218_, _079222_);
  or g_135417_(_078336_, _079222_, _079223_);
  xor g_135418_(_078336_, _079221_, _079224_);
  or g_135419_(_078334_, _079224_, _079225_);
  xor g_135420_(_078335_, _079224_, _079226_);
  or g_135421_(_078332_, _079226_, _079227_);
  not g_135422_(_079227_, _079228_);
  xor g_135423_(_078333_, _079226_, _079229_);
  not g_135424_(_079229_, _079231_);
  or g_135425_(_078331_, _079229_, _079232_);
  not g_135426_(_079232_, _079233_);
  xor g_135427_(_078331_, _079229_, _079234_);
  xor g_135428_(_078331_, _079231_, _079235_);
  or g_135429_(_078330_, _079235_, _079236_);
  xor g_135430_(_078330_, _079234_, _079237_);
  or g_135431_(_073454_, _076354_, _079238_);
  not g_135432_(_079238_, _079239_);
  or g_135433_(_079237_, _079238_, _079240_);
  xor g_135434_(_079237_, _079239_, _079242_);
  or g_135435_(_076357_, _079242_, _079243_);
  xor g_135436_(_076358_, _079242_, _079244_);
  and g_135437_(_076362_, _076366_, _079245_);
  xor g_135438_(_079244_, _079245_, _079246_);
  not g_135439_(_079246_, _079247_);
  and g_135440_(_076368_, _079246_, _079248_);
  or g_135441_(_076367_, _079247_, _079249_);
  xor g_135442_(_076367_, _079246_, _079250_);
  or g_135443_(_076377_, _079250_, _079251_);
  not g_135444_(_079251_, _079253_);
  xor g_135445_(_076376_, _079250_, _079254_);
  or g_135446_(_076372_, _079254_, _079255_);
  not g_135447_(_079255_, _079256_);
  xor g_135448_(_076372_, _079254_, _079257_);
  xor g_135449_(_076373_, _079254_, _079258_);
  xor g_135450_(_076380_, _079257_, _079259_);
  or g_135451_(_076387_, _079259_, _079260_);
  xor g_135452_(_076387_, _079259_, _079261_);
  not g_135453_(_079261_, _079262_);
  or g_135454_(_076385_, _079262_, _079264_);
  xor g_135455_(_076385_, _079261_, _079265_);
  not g_135456_(_079265_, _079266_);
  xor g_135457_(_076398_, _079266_, _079267_);
  xor g_135458_(_076405_, _079267_, _079268_);
  not g_135459_(_079268_, _079269_);
  xor g_135460_(_078329_, _079268_, _079270_);
  xor g_135461_(_078327_, _079270_, _079271_);
  not g_135462_(_079271_, _079272_);
  or g_135463_(_076423_, _079272_, _079273_);
  xor g_135464_(_076423_, _079271_, _079275_);
  not g_135465_(_079275_, _079276_);
  or g_135466_(_076425_, _079275_, _079277_);
  xor g_135467_(_076425_, _079275_, _079278_);
  xor g_135468_(_076425_, _079276_, _079279_);
  or g_135469_(_076430_, _079279_, _079280_);
  xor g_135470_(_076430_, _079278_, _079281_);
  or g_135471_(_076431_, _079281_, _079282_);
  xor g_135472_(_076432_, _079281_, _079283_);
  or g_135473_(_076436_, _079283_, _079284_);
  xor g_135474_(_076438_, _079283_, _079286_);
  not g_135475_(_079286_, _079287_);
  xor g_135476_(_076439_, _079287_, _079288_);
  or g_135477_(_076444_, _079288_, _079289_);
  not g_135478_(_079289_, _079290_);
  xor g_135479_(_076445_, _079288_, _079291_);
  not g_135480_(_079291_, _079292_);
  or g_135481_(_073536_, _076442_, _079293_);
  or g_135482_(_079291_, _079293_, _079294_);
  not g_135483_(_079294_, _079295_);
  xor g_135484_(_079292_, _079293_, _079297_);
  not g_135485_(_079297_, _079298_);
  or g_135486_(_073539_, _076446_, _079299_);
  or g_135487_(_079297_, _079299_, _079300_);
  not g_135488_(_079300_, _079301_);
  xor g_135489_(_079298_, _079299_, _079302_);
  or g_135490_(_073541_, _076450_, _079303_);
  or g_135491_(_079302_, _079303_, _079304_);
  not g_135492_(_079304_, _079305_);
  xor g_135493_(_079302_, _079303_, _079306_);
  not g_135494_(_079306_, _079308_);
  or g_135495_(_078326_, _079308_, _079309_);
  xor g_135496_(_078326_, _079306_, _079310_);
  not g_135497_(_079310_, _079311_);
  and g_135498_(_076453_, _076455_, _079312_);
  xor g_135499_(_079311_, _079312_, _079313_);
  xor g_135500_(_079310_, _079312_, _079314_);
  or g_135501_(_078325_, _079313_, _079315_);
  xor g_135502_(_078325_, _079314_, _079316_);
  or g_135503_(_073555_, _076457_, _079317_);
  or g_135504_(_079316_, _079317_, _079319_);
  not g_135505_(_079319_, _079320_);
  xor g_135506_(_079316_, _079317_, _079321_);
  and g_135507_(_076463_, _079321_, _079322_);
  xor g_135508_(_076463_, _079321_, _079323_);
  xor g_135509_(_076464_, _079321_, _079324_);
  or g_135510_(_076465_, _079324_, _079325_);
  not g_135511_(_079325_, _079326_);
  xor g_135512_(_076465_, _079323_, _079327_);
  and g_135513_(_076468_, _076472_, _079328_);
  and g_135514_(_079327_, _079328_, _079330_);
  not g_135515_(_079330_, _079331_);
  or g_135516_(_076472_, _079327_, _079332_);
  or g_135517_(_076468_, _079327_, _079333_);
  not g_135518_(_079333_, _079334_);
  and g_135519_(_079332_, _079333_, _079335_);
  not g_135520_(_079335_, _079336_);
  and g_135521_(_079331_, _079335_, _079337_);
  or g_135522_(_079330_, _079336_, _079338_);
  xor g_135523_(_078324_, _079337_, _079339_);
  or g_135524_(_076485_, _079339_, _079341_);
  xor g_135525_(_076485_, _079339_, _079342_);
  not g_135526_(_079342_, _079343_);
  or g_135527_(_076486_, _079343_, _079344_);
  xor g_135528_(_076486_, _079342_, _079345_);
  or g_135529_(_076488_, _079345_, _079346_);
  not g_135530_(_079346_, _079347_);
  xor g_135531_(_076488_, _079345_, _079348_);
  not g_135532_(_079348_, _079349_);
  or g_135533_(_076490_, _079349_, _079350_);
  not g_135534_(_079350_, _079352_);
  xor g_135535_(_076490_, _079348_, _079353_);
  or g_135536_(_076493_, _079353_, _079354_);
  xor g_135537_(_076494_, _079353_, _079355_);
  not g_135538_(_079355_, _079356_);
  or g_135539_(_076498_, _079355_, _079357_);
  xor g_135540_(_076498_, _079355_, _079358_);
  xor g_135541_(_076498_, _079356_, _079359_);
  or g_135542_(_076499_, _079359_, _079360_);
  xor g_135543_(_076499_, _079358_, _079361_);
  or g_135544_(_076506_, _079361_, _079363_);
  xor g_135545_(_076505_, _079361_, _079364_);
  and g_135546_(_076507_, _076512_, _079365_);
  xor g_135547_(_079364_, _079365_, _079366_);
  not g_135548_(_079366_, _079367_);
  or g_135549_(_078323_, _079367_, _079368_);
  not g_135550_(_079368_, _079369_);
  xor g_135551_(_078323_, _079366_, _079370_);
  or g_135552_(_078322_, _079370_, _079371_);
  xor g_135553_(_078321_, _079370_, _079372_);
  or g_135554_(_076519_, _079372_, _079374_);
  not g_135555_(_079374_, _079375_);
  xor g_135556_(_076520_, _079372_, _079376_);
  or g_135557_(_073619_, _076517_, _079377_);
  not g_135558_(_079377_, _079378_);
  or g_135559_(_079376_, _079377_, _079379_);
  xor g_135560_(_079376_, _079377_, _079380_);
  xor g_135561_(_079376_, _079378_, _079381_);
  or g_135562_(_078320_, _079381_, _079382_);
  xor g_135563_(_078320_, _079380_, _079383_);
  not g_135564_(_079383_, _079385_);
  or g_135565_(_076532_, _079383_, _079386_);
  xor g_135566_(_076532_, _079383_, _079387_);
  xor g_135567_(_076532_, _079385_, _079388_);
  or g_135568_(_076533_, _079388_, _079389_);
  xor g_135569_(_076533_, _079387_, _079390_);
  or g_135570_(_076529_, _079390_, _079391_);
  not g_135571_(_079391_, _079392_);
  xor g_135572_(_076529_, _079390_, _079393_);
  not g_135573_(_079393_, _079394_);
  and g_135574_(_076538_, _079393_, _079396_);
  or g_135575_(_076537_, _079394_, _079397_);
  xor g_135576_(_076537_, _079393_, _079398_);
  not g_135577_(_079398_, _079399_);
  and g_135578_(_073640_, _076530_, _079400_);
  or g_135579_(_073639_, _076531_, _079401_);
  and g_135580_(_079399_, _079400_, _079402_);
  or g_135581_(_079398_, _079401_, _079403_);
  xor g_135582_(_079398_, _079401_, _079404_);
  xor g_135583_(_079398_, _079400_, _079405_);
  or g_135584_(_078319_, _079405_, _079407_);
  not g_135585_(_079407_, _079408_);
  xor g_135586_(_078319_, _079404_, _079409_);
  and g_135587_(_076545_, _076555_, _079410_);
  xor g_135588_(_079409_, _079410_, _079411_);
  not g_135589_(_079411_, _079412_);
  or g_135590_(_076554_, _079412_, _079413_);
  xor g_135591_(_076554_, _079411_, _079414_);
  not g_135592_(_079414_, _079415_);
  and g_135593_(_076551_, _076556_, _079416_);
  xor g_135594_(_079415_, _079416_, _079418_);
  or g_135595_(_076560_, _079418_, _079419_);
  not g_135596_(_079419_, _079420_);
  xor g_135597_(_076560_, _079418_, _079421_);
  not g_135598_(_079421_, _079422_);
  or g_135599_(_073669_, _076559_, _079423_);
  or g_135600_(_079422_, _079423_, _079424_);
  not g_135601_(_079424_, _079425_);
  xor g_135602_(_079421_, _079423_, _079426_);
  or g_135603_(_073672_, _076561_, _079427_);
  or g_135604_(_079426_, _079427_, _079429_);
  not g_135605_(_079429_, _079430_);
  xor g_135606_(_079426_, _079427_, _079431_);
  and g_135607_(_076571_, _079431_, _079432_);
  not g_135608_(_079432_, _079433_);
  xor g_135609_(_076570_, _079431_, _079434_);
  or g_135610_(_076567_, _079434_, _079435_);
  xor g_135611_(_076566_, _079434_, _079436_);
  and g_135612_(_076574_, _076579_, _079437_);
  and g_135613_(_079436_, _079437_, _079438_);
  or g_135614_(_076579_, _079436_, _079440_);
  not g_135615_(_079440_, _079441_);
  or g_135616_(_076574_, _079436_, _079442_);
  and g_135617_(_079440_, _079442_, _079443_);
  not g_135618_(_079443_, _079444_);
  or g_135619_(_079438_, _079444_, _079445_);
  not g_135620_(_079445_, _079446_);
  xor g_135621_(_078318_, _079446_, _079447_);
  or g_135622_(_076595_, _079447_, _079448_);
  xor g_135623_(_076595_, _079447_, _079449_);
  xor g_135624_(_076594_, _079447_, _079451_);
  and g_135625_(_076598_, _076604_, _079452_);
  xor g_135626_(_079449_, _079452_, _079453_);
  or g_135627_(_076607_, _079453_, _079454_);
  not g_135628_(_079454_, _079455_);
  or g_135629_(_073704_, _076600_, _079456_);
  and g_135630_(_079453_, _079456_, _079457_);
  and g_135631_(_076607_, _079457_, _079458_);
  or g_135632_(_079453_, _079456_, _079459_);
  not g_135633_(_079459_, _079460_);
  or g_135634_(_079458_, _079460_, _079462_);
  or g_135635_(_079455_, _079462_, _079463_);
  not g_135636_(_079463_, _079464_);
  xor g_135637_(_078316_, _079463_, _079465_);
  xor g_135638_(_078316_, _079464_, _079466_);
  or g_135639_(_078315_, _079466_, _079467_);
  xor g_135640_(_078315_, _079465_, _079468_);
  not g_135641_(_079468_, _079469_);
  and g_135642_(_078313_, _079469_, _079470_);
  or g_135643_(_078314_, _079468_, _079471_);
  xor g_135644_(_078313_, _079468_, _079473_);
  not g_135645_(_079473_, _079474_);
  and g_135646_(_078311_, _079474_, _079475_);
  or g_135647_(_078312_, _079473_, _079476_);
  xor g_135648_(_078311_, _079473_, _079477_);
  not g_135649_(_079477_, _079478_);
  or g_135650_(_078310_, _079477_, _079479_);
  xor g_135651_(_078310_, _079477_, _079480_);
  xor g_135652_(_078310_, _079478_, _079481_);
  or g_135653_(_076621_, _079481_, _079482_);
  xor g_135654_(_076621_, _079480_, _079484_);
  or g_135655_(_076625_, _079484_, _079485_);
  xor g_135656_(_076626_, _079484_, _079486_);
  not g_135657_(_079486_, _079487_);
  and g_135658_(_076629_, _076633_, _079488_);
  xor g_135659_(_079487_, _079488_, _079489_);
  or g_135660_(_076639_, _079489_, _079490_);
  xor g_135661_(_076640_, _079489_, _079491_);
  or g_135662_(_073746_, _076636_, _079492_);
  or g_135663_(_079491_, _079492_, _079493_);
  xor g_135664_(_079491_, _079492_, _079495_);
  and g_135665_(_078309_, _079495_, _079496_);
  not g_135666_(_079496_, _079497_);
  xor g_135667_(_078308_, _079495_, _079498_);
  not g_135668_(_079498_, _079499_);
  and g_135669_(_076649_, _076652_, _079500_);
  xor g_135670_(_079499_, _079500_, _079501_);
  xor g_135671_(_079498_, _079500_, _079502_);
  or g_135672_(_076655_, _079501_, _079503_);
  xor g_135673_(_076655_, _079502_, _079504_);
  or g_135674_(_073764_, _076653_, _079506_);
  or g_135675_(_079504_, _079506_, _079507_);
  xor g_135676_(_079504_, _079506_, _079508_);
  and g_135677_(_078307_, _079508_, _079509_);
  not g_135678_(_079509_, _079510_);
  xor g_135679_(_078305_, _079508_, _079511_);
  or g_135680_(_076663_, _079511_, _079512_);
  xor g_135681_(_076663_, _079511_, _079513_);
  xor g_135682_(_076662_, _079511_, _079514_);
  or g_135683_(_076664_, _079514_, _079515_);
  xor g_135684_(_076664_, _079513_, _079517_);
  not g_135685_(_079517_, _079518_);
  or g_135686_(_076672_, _079517_, _079519_);
  xor g_135687_(_076672_, _079517_, _079520_);
  xor g_135688_(_076672_, _079518_, _079521_);
  or g_135689_(_076675_, _079521_, _079522_);
  xor g_135690_(_076675_, _079520_, _079523_);
  or g_135691_(_076680_, _079523_, _079524_);
  xor g_135692_(_076680_, _079523_, _079525_);
  not g_135693_(_079525_, _079526_);
  and g_135694_(_078304_, _079525_, _079528_);
  or g_135695_(_078303_, _079526_, _079529_);
  xor g_135696_(_078303_, _079525_, _079530_);
  not g_135697_(_079530_, _079531_);
  or g_135698_(_078302_, _079530_, _079532_);
  xor g_135699_(_078302_, _079531_, _079533_);
  and g_135700_(_076687_, _076689_, _079534_);
  xor g_135701_(_079533_, _079534_, _079535_);
  not g_135702_(_079535_, _079536_);
  or g_135703_(_076693_, _079536_, _079537_);
  not g_135704_(_079537_, _079539_);
  xor g_135705_(_076693_, _079535_, _079540_);
  or g_135706_(_073802_, _076691_, _079541_);
  or g_135707_(_079540_, _079541_, _079542_);
  not g_135708_(_079542_, _079543_);
  xor g_135709_(_079540_, _079541_, _079544_);
  not g_135710_(_079544_, _079545_);
  or g_135711_(_078301_, _079545_, _079546_);
  not g_135712_(_079546_, _079547_);
  xor g_135713_(_078301_, _079544_, _079548_);
  not g_135714_(_079548_, _079550_);
  or g_135715_(_076699_, _079548_, _079551_);
  not g_135716_(_079551_, _079552_);
  xor g_135717_(_076699_, _079550_, _079553_);
  or g_135718_(_073813_, _076698_, _079554_);
  or g_135719_(_079553_, _079554_, _079555_);
  not g_135720_(_079555_, _079556_);
  xor g_135721_(_079553_, _079554_, _079557_);
  not g_135722_(_079557_, _079558_);
  or g_135723_(_073816_, _076700_, _079559_);
  or g_135724_(_079558_, _079559_, _079561_);
  not g_135725_(_079561_, _079562_);
  xor g_135726_(_079557_, _079559_, _079563_);
  or g_135727_(_076709_, _079563_, _079564_);
  not g_135728_(_079564_, _079565_);
  xor g_135729_(_076708_, _079563_, _079566_);
  not g_135730_(_079566_, _079567_);
  and g_135731_(_076706_, _079567_, _079568_);
  or g_135732_(_076707_, _079566_, _079569_);
  xor g_135733_(_076706_, _079566_, _079570_);
  and g_135734_(_076713_, _076716_, _079572_);
  not g_135735_(_079572_, _079573_);
  xor g_135736_(_079570_, _079573_, _079574_);
  not g_135737_(_079574_, _079575_);
  or g_135738_(_076715_, _079574_, _079576_);
  xor g_135739_(_076715_, _079575_, _079577_);
  or g_135740_(_076725_, _079577_, _079578_);
  not g_135741_(_079578_, _079579_);
  and g_135742_(_076721_, _079577_, _079580_);
  and g_135743_(_076725_, _079580_, _079581_);
  or g_135744_(_076721_, _079577_, _079583_);
  not g_135745_(_079583_, _079584_);
  or g_135746_(_079581_, _079584_, _079585_);
  or g_135747_(_079579_, _079585_, _079586_);
  or g_135748_(_076729_, _079586_, _079587_);
  xor g_135749_(_076730_, _079586_, _079588_);
  or g_135750_(_076727_, _079588_, _079589_);
  or g_135751_(_073848_, _076735_, _079590_);
  or g_135752_(_079588_, _079590_, _079591_);
  and g_135753_(_079589_, _079591_, _079592_);
  not g_135754_(_079592_, _079594_);
  and g_135755_(_076727_, _079588_, _079595_);
  and g_135756_(_079590_, _079595_, _079596_);
  or g_135757_(_079594_, _079596_, _079597_);
  not g_135758_(_079597_, _079598_);
  or g_135759_(_078300_, _079597_, _079599_);
  xor g_135760_(_078300_, _079598_, _079600_);
  or g_135761_(_076739_, _079600_, _079601_);
  xor g_135762_(_076740_, _079600_, _079602_);
  or g_135763_(_076743_, _079602_, _079603_);
  xor g_135764_(_076743_, _079602_, _079605_);
  not g_135765_(_079605_, _079606_);
  or g_135766_(_073859_, _076742_, _079607_);
  or g_135767_(_079606_, _079607_, _079608_);
  xor g_135768_(_079605_, _079607_, _079609_);
  or g_135769_(_078299_, _079609_, _079610_);
  xor g_135770_(_078299_, _079609_, _079611_);
  not g_135771_(_079611_, _079612_);
  and g_135772_(_076750_, _076752_, _079613_);
  xor g_135773_(_079612_, _079613_, _079614_);
  and g_135774_(_076760_, _079614_, _079616_);
  not g_135775_(_079616_, _079617_);
  xor g_135776_(_076759_, _079614_, _079618_);
  or g_135777_(_076766_, _079618_, _079619_);
  xor g_135778_(_076768_, _079618_, _079620_);
  or g_135779_(_076764_, _079620_, _079621_);
  xor g_135780_(_076763_, _079620_, _079622_);
  not g_135781_(_079622_, _079623_);
  and g_135782_(_076774_, _079623_, _079624_);
  or g_135783_(_076775_, _079622_, _079625_);
  xor g_135784_(_076774_, _079622_, _079627_);
  or g_135785_(_076781_, _079627_, _079628_);
  xor g_135786_(_076782_, _079627_, _079629_);
  or g_135787_(_076777_, _079629_, _079630_);
  xor g_135788_(_076779_, _079629_, _079631_);
  and g_135789_(_076787_, _076794_, _079632_);
  not g_135790_(_079632_, _079633_);
  xor g_135791_(_079631_, _079633_, _079634_);
  or g_135792_(_076792_, _079634_, _079635_);
  xor g_135793_(_076793_, _079634_, _079636_);
  not g_135794_(_079636_, _079638_);
  or g_135795_(_076803_, _079636_, _079639_);
  xor g_135796_(_076803_, _079636_, _079640_);
  xor g_135797_(_076803_, _079638_, _079641_);
  or g_135798_(_073907_, _076801_, _079642_);
  or g_135799_(_079641_, _079642_, _079643_);
  xor g_135800_(_079640_, _079642_, _079644_);
  or g_135801_(_076806_, _079644_, _079645_);
  xor g_135802_(_076805_, _079644_, _079646_);
  xor g_135803_(_076817_, _079646_, _079647_);
  not g_135804_(_079647_, _079649_);
  xor g_135805_(_078298_, _079647_, _079650_);
  not g_135806_(_079650_, _079651_);
  or g_135807_(_076831_, _079651_, _079652_);
  not g_135808_(_079652_, _079653_);
  xor g_135809_(_076831_, _079650_, _079654_);
  or g_135810_(_078296_, _079654_, _079655_);
  not g_135811_(_079655_, _079656_);
  xor g_135812_(_078297_, _079654_, _079657_);
  or g_135813_(_078293_, _079657_, _079658_);
  xor g_135814_(_078294_, _079657_, _079660_);
  or g_135815_(_076837_, _079660_, _079661_);
  not g_135816_(_079661_, _079662_);
  or g_135817_(_076840_, _079660_, _079663_);
  xor g_135818_(_076840_, _079660_, _079664_);
  xor g_135819_(_076841_, _079660_, _079665_);
  and g_135820_(_076837_, _079665_, _079666_);
  or g_135821_(_076838_, _079664_, _079667_);
  and g_135822_(_079661_, _079667_, _079668_);
  or g_135823_(_079662_, _079666_, _079669_);
  or g_135824_(_078292_, _079669_, _079671_);
  not g_135825_(_079671_, _079672_);
  xor g_135826_(_078292_, _079669_, _079673_);
  xor g_135827_(_078292_, _079668_, _079674_);
  and g_135828_(_078290_, _079673_, _079675_);
  or g_135829_(_078291_, _079674_, _079676_);
  xor g_135830_(_078291_, _079673_, _079677_);
  or g_135831_(_076851_, _079677_, _079678_);
  xor g_135832_(_076851_, _079677_, _079679_);
  xor g_135833_(_076852_, _079677_, _079680_);
  and g_135834_(_076848_, _079679_, _079682_);
  or g_135835_(_076847_, _079680_, _079683_);
  xor g_135836_(_076847_, _079679_, _079684_);
  not g_135837_(_079684_, _079685_);
  and g_135838_(_076854_, _076860_, _079686_);
  or g_135839_(_079684_, _079686_, _079687_);
  xor g_135840_(_079684_, _079686_, _079688_);
  xor g_135841_(_079685_, _079686_, _079689_);
  or g_135842_(_078289_, _079689_, _079690_);
  not g_135843_(_079690_, _079691_);
  xor g_135844_(_078289_, _079688_, _079693_);
  or g_135845_(_078288_, _079693_, _079694_);
  not g_135846_(_079694_, _079695_);
  xor g_135847_(_078287_, _079693_, _079696_);
  not g_135848_(_079696_, _079697_);
  and g_135849_(_078285_, _079697_, _079698_);
  or g_135850_(_078286_, _079696_, _079699_);
  xor g_135851_(_078285_, _079696_, _079700_);
  and g_135852_(_073981_, _076864_, _079701_);
  or g_135853_(_073980_, _076865_, _079702_);
  or g_135854_(_079700_, _079702_, _079704_);
  xor g_135855_(_079700_, _079701_, _079705_);
  and g_135856_(_076868_, _076874_, _079706_);
  xor g_135857_(_079705_, _079706_, _079707_);
  not g_135858_(_079707_, _079708_);
  and g_135859_(_076871_, _079707_, _079709_);
  or g_135860_(_076870_, _079708_, _079710_);
  xor g_135861_(_076871_, _079707_, _079711_);
  not g_135862_(_079711_, _079712_);
  and g_135863_(_076879_, _079711_, _079713_);
  or g_135864_(_076878_, _079712_, _079715_);
  xor g_135865_(_076878_, _079711_, _079716_);
  and g_135866_(_076880_, _079716_, _079717_);
  or g_135867_(_076880_, _079716_, _079718_);
  not g_135868_(_079718_, _079719_);
  xor g_135869_(_076880_, _079716_, _079720_);
  or g_135870_(_079717_, _079719_, _079721_);
  or g_135871_(_073999_, _076884_, _079722_);
  or g_135872_(_079721_, _079722_, _079723_);
  xor g_135873_(_079720_, _079722_, _079724_);
  not g_135874_(_079724_, _079726_);
  or g_135875_(_078283_, _079724_, _079727_);
  xor g_135876_(_078283_, _079726_, _079728_);
  or g_135877_(_076891_, _079728_, _079729_);
  xor g_135878_(_076891_, _079728_, _079730_);
  xor g_135879_(_076892_, _079728_, _079731_);
  and g_135880_(_076894_, _079730_, _079732_);
  or g_135881_(_076893_, _079731_, _079733_);
  xor g_135882_(_076893_, _079730_, _079734_);
  not g_135883_(_079734_, _079735_);
  or g_135884_(_076895_, _076900_, _079737_);
  not g_135885_(_079737_, _079738_);
  and g_135886_(_079734_, _079738_, _079739_);
  or g_135887_(_076901_, _079734_, _079740_);
  not g_135888_(_079740_, _079741_);
  and g_135889_(_076895_, _079735_, _079742_);
  or g_135890_(_076896_, _079734_, _079743_);
  or g_135891_(_079741_, _079742_, _079744_);
  or g_135892_(_079739_, _079744_, _079745_);
  not g_135893_(_079745_, _079746_);
  xor g_135894_(_078282_, _079746_, _079748_);
  not g_135895_(_079748_, _079749_);
  xor g_135896_(_076916_, _079749_, _079750_);
  not g_135897_(_079750_, _079751_);
  xor g_135898_(_078281_, _079751_, _079752_);
  or g_135899_(_076933_, _079752_, _079753_);
  not g_135900_(_079753_, _079754_);
  or g_135901_(_076928_, _079752_, _079755_);
  xor g_135902_(_076929_, _079752_, _079756_);
  and g_135903_(_076933_, _079756_, _079757_);
  or g_135904_(_079754_, _079757_, _079759_);
  not g_135905_(_079759_, _079760_);
  and g_135906_(_076937_, _076940_, _079761_);
  xor g_135907_(_079759_, _079761_, _079762_);
  xor g_135908_(_079760_, _079761_, _079763_);
  or g_135909_(_076944_, _079763_, _079764_);
  xor g_135910_(_076944_, _079762_, _079765_);
  or g_135911_(_074061_, _076941_, _079766_);
  not g_135912_(_079766_, _079767_);
  or g_135913_(_079765_, _079766_, _079768_);
  xor g_135914_(_079765_, _079766_, _079770_);
  xor g_135915_(_079765_, _079767_, _079771_);
  or g_135916_(_074065_, _076945_, _079772_);
  or g_135917_(_079771_, _079772_, _079773_);
  xor g_135918_(_079770_, _079772_, _079774_);
  or g_135919_(_076952_, _079774_, _079775_);
  xor g_135920_(_076953_, _079774_, _079776_);
  or g_135921_(_076949_, _079776_, _079777_);
  xor g_135922_(_076949_, _079776_, _079778_);
  not g_135923_(_079778_, _079779_);
  or g_135924_(_078280_, _079779_, _079781_);
  not g_135925_(_079781_, _079782_);
  xor g_135926_(_078280_, _079778_, _079783_);
  or g_135927_(_078279_, _079783_, _079784_);
  xor g_135928_(_078278_, _079783_, _079785_);
  not g_135929_(_079785_, _079786_);
  and g_135930_(_076959_, _076962_, _079787_);
  xor g_135931_(_079786_, _079787_, _079788_);
  or g_135932_(_076966_, _079788_, _079789_);
  xor g_135933_(_076967_, _079788_, _079790_);
  or g_135934_(_074090_, _076963_, _079792_);
  not g_135935_(_079792_, _079793_);
  or g_135936_(_079790_, _079792_, _079794_);
  xor g_135937_(_079790_, _079792_, _079795_);
  xor g_135938_(_079790_, _079793_, _079796_);
  or g_135939_(_078277_, _079796_, _079797_);
  not g_135940_(_079797_, _079798_);
  xor g_135941_(_078277_, _079795_, _079799_);
  or g_135942_(_076980_, _079799_, _079800_);
  not g_135943_(_079800_, _079801_);
  xor g_135944_(_076981_, _079799_, _079803_);
  or g_135945_(_076973_, _079803_, _079804_);
  not g_135946_(_079804_, _079805_);
  xor g_135947_(_076974_, _079803_, _079806_);
  or g_135948_(_074103_, _076988_, _079807_);
  and g_135949_(_076986_, _079807_, _079808_);
  not g_135950_(_079808_, _079809_);
  xor g_135951_(_079806_, _079809_, _079810_);
  or g_135952_(_078276_, _079810_, _079811_);
  xor g_135953_(_078276_, _079810_, _079812_);
  not g_135954_(_079812_, _079814_);
  or g_135955_(_076991_, _079814_, _079815_);
  not g_135956_(_079815_, _079816_);
  xor g_135957_(_076991_, _079812_, _079817_);
  or g_135958_(_076995_, _079817_, _079818_);
  xor g_135959_(_076994_, _079817_, _079819_);
  or g_135960_(_074116_, _076992_, _079820_);
  not g_135961_(_079820_, _079821_);
  or g_135962_(_079819_, _079820_, _079822_);
  xor g_135963_(_079819_, _079821_, _079823_);
  not g_135964_(_079823_, _079825_);
  or g_135965_(_078275_, _079823_, _079826_);
  xor g_135966_(_078275_, _079825_, _079827_);
  not g_135967_(_079827_, _079828_);
  or g_135968_(_074125_, _077000_, _079829_);
  and g_135969_(_077001_, _079829_, _079830_);
  xor g_135970_(_079827_, _079830_, _079831_);
  xor g_135971_(_079828_, _079830_, _079832_);
  or g_135972_(_078274_, _079832_, _079833_);
  xor g_135973_(_078274_, _079831_, _079834_);
  or g_135974_(_077006_, _079834_, _079836_);
  not g_135975_(_079836_, _079837_);
  xor g_135976_(_077007_, _079834_, _079838_);
  and g_135977_(_077011_, _077014_, _079839_);
  not g_135978_(_079839_, _079840_);
  xor g_135979_(_079838_, _079840_, _079841_);
  xor g_135980_(_078272_, _079841_, _079842_);
  or g_135981_(_077026_, _077029_, _079843_);
  xor g_135982_(_079842_, _079843_, _079844_);
  not g_135983_(_079844_, _079845_);
  or g_135984_(_074157_, _077037_, _079847_);
  and g_135985_(_077035_, _079847_, _079848_);
  xor g_135986_(_079844_, _079848_, _079849_);
  xor g_135987_(_079845_, _079848_, _079850_);
  or g_135988_(_078270_, _079850_, _079851_);
  not g_135989_(_079851_, _079852_);
  xor g_135990_(_078270_, _079849_, _079853_);
  and g_135991_(_077045_, _079853_, _079854_);
  or g_135992_(_077044_, _079853_, _079855_);
  not g_135993_(_079855_, _079856_);
  or g_135994_(_077043_, _079853_, _079858_);
  not g_135995_(_079858_, _079859_);
  and g_135996_(_079855_, _079858_, _079860_);
  not g_135997_(_079860_, _079861_);
  or g_135998_(_079854_, _079861_, _079862_);
  not g_135999_(_079862_, _079863_);
  xor g_136000_(_077047_, _079863_, _079864_);
  xor g_136001_(_078269_, _079864_, _079865_);
  not g_136002_(_079865_, _079866_);
  or g_136003_(_078268_, _079866_, _079867_);
  xor g_136004_(_078268_, _079865_, _079869_);
  or g_136005_(_078267_, _079869_, _079870_);
  xor g_136006_(_078266_, _079869_, _079871_);
  or g_136007_(_077060_, _079871_, _079872_);
  xor g_136008_(_077059_, _079871_, _079873_);
  or g_136009_(_077067_, _079873_, _079874_);
  not g_136010_(_079874_, _079875_);
  xor g_136011_(_077066_, _079873_, _079876_);
  or g_136012_(_077072_, _079876_, _079877_);
  xor g_136013_(_077072_, _079876_, _079878_);
  xor g_136014_(_077073_, _079876_, _079880_);
  or g_136015_(_077079_, _079880_, _079881_);
  xor g_136016_(_077079_, _079878_, _079882_);
  xor g_136017_(_077077_, _079882_, _079883_);
  or g_136018_(_077084_, _079883_, _079884_);
  xor g_136019_(_077085_, _079883_, _079885_);
  or g_136020_(_077089_, _079885_, _079886_);
  xor g_136021_(_077089_, _079885_, _079887_);
  xor g_136022_(_077090_, _079885_, _079888_);
  or g_136023_(_074217_, _077095_, _079889_);
  and g_136024_(_077093_, _079889_, _079891_);
  xor g_136025_(_079887_, _079891_, _079892_);
  or g_136026_(_078265_, _079892_, _079893_);
  not g_136027_(_079893_, _079894_);
  xor g_136028_(_078265_, _079892_, _079895_);
  not g_136029_(_079895_, _079896_);
  and g_136030_(_077101_, _079895_, _079897_);
  or g_136031_(_077100_, _079896_, _079898_);
  xor g_136032_(_077100_, _079895_, _079899_);
  or g_136033_(_077104_, _079899_, _079900_);
  xor g_136034_(_077105_, _079899_, _079902_);
  or g_136035_(_074229_, _077102_, _079903_);
  not g_136036_(_079903_, _079904_);
  or g_136037_(_079902_, _079903_, _079905_);
  xor g_136038_(_079902_, _079903_, _079906_);
  xor g_136039_(_079902_, _079904_, _079907_);
  or g_136040_(_074232_, _077106_, _079908_);
  or g_136041_(_079907_, _079908_, _079909_);
  xor g_136042_(_079906_, _079908_, _079910_);
  not g_136043_(_079910_, _079911_);
  and g_136044_(_077112_, _077114_, _079913_);
  xor g_136045_(_079911_, _079913_, _079914_);
  or g_136046_(_077115_, _079914_, _079915_);
  not g_136047_(_079915_, _079916_);
  xor g_136048_(_077115_, _079914_, _079917_);
  and g_136049_(_077121_, _079917_, _079918_);
  not g_136050_(_079918_, _079919_);
  xor g_136051_(_077122_, _079917_, _079920_);
  or g_136052_(_077123_, _079920_, _079921_);
  xor g_136053_(_077124_, _079920_, _079922_);
  or g_136054_(_078263_, _079922_, _079924_);
  not g_136055_(_079924_, _079925_);
  xor g_136056_(_078264_, _079922_, _079926_);
  not g_136057_(_079926_, _079927_);
  or g_136058_(_074254_, _077127_, _079928_);
  and g_136059_(_077136_, _079928_, _079929_);
  xor g_136060_(_079927_, _079929_, _079930_);
  xor g_136061_(_079926_, _079929_, _079931_);
  and g_136062_(_077132_, _077140_, _079932_);
  or g_136063_(_079930_, _079932_, _079933_);
  xor g_136064_(_079931_, _079932_, _079935_);
  not g_136065_(_079935_, _079936_);
  or g_136066_(_078261_, _079935_, _079937_);
  xor g_136067_(_078261_, _079935_, _079938_);
  xor g_136068_(_078261_, _079936_, _079939_);
  or g_136069_(_078260_, _079939_, _079940_);
  xor g_136070_(_078260_, _079938_, _079941_);
  or g_136071_(_077146_, _079941_, _079942_);
  xor g_136072_(_077147_, _079941_, _079943_);
  or g_136073_(_074276_, _077144_, _079944_);
  or g_136074_(_079943_, _079944_, _079946_);
  xor g_136075_(_079943_, _079944_, _079947_);
  not g_136076_(_079947_, _079948_);
  or g_136077_(_078259_, _079948_, _079949_);
  xor g_136078_(_078259_, _079947_, _079950_);
  or g_136079_(_077153_, _079950_, _079951_);
  xor g_136080_(_077154_, _079950_, _079952_);
  or g_136081_(_074285_, _077151_, _079953_);
  not g_136082_(_079953_, _079954_);
  or g_136083_(_079952_, _079953_, _079955_);
  xor g_136084_(_079952_, _079954_, _079957_);
  or g_136085_(_074288_, _077156_, _079958_);
  or g_136086_(_079957_, _079958_, _079959_);
  xor g_136087_(_079957_, _079958_, _079960_);
  not g_136088_(_079960_, _079961_);
  or g_136089_(_078258_, _079961_, _079962_);
  xor g_136090_(_078258_, _079960_, _079963_);
  or g_136091_(_078256_, _079963_, _079964_);
  not g_136092_(_079964_, _079965_);
  xor g_136093_(_078257_, _079963_, _079966_);
  or g_136094_(_077162_, _079966_, _079968_);
  xor g_136095_(_077162_, _079966_, _079969_);
  not g_136096_(_079969_, _079970_);
  or g_136097_(_077166_, _079970_, _079971_);
  xor g_136098_(_077166_, _079969_, _079972_);
  or g_136099_(_077170_, _079972_, _079973_);
  xor g_136100_(_077171_, _079972_, _079974_);
  not g_136101_(_079974_, _079975_);
  and g_136102_(_077175_, _077178_, _079976_);
  xor g_136103_(_079975_, _079976_, _079977_);
  or g_136104_(_077182_, _079977_, _079979_);
  xor g_136105_(_077183_, _079977_, _079980_);
  not g_136106_(_079980_, _079981_);
  and g_136107_(_077180_, _077189_, _079982_);
  xor g_136108_(_079981_, _079982_, _079983_);
  or g_136109_(_077192_, _079983_, _079984_);
  not g_136110_(_079984_, _079985_);
  xor g_136111_(_077193_, _079983_, _079986_);
  or g_136112_(_074322_, _077194_, _079987_);
  not g_136113_(_079987_, _079988_);
  xor g_136114_(_079986_, _079987_, _079990_);
  xor g_136115_(_079986_, _079988_, _079991_);
  or g_136116_(_078255_, _079991_, _079992_);
  xor g_136117_(_078255_, _079990_, _079993_);
  and g_136118_(_074328_, _077198_, _079994_);
  or g_136119_(_074327_, _077199_, _079995_);
  or g_136120_(_079993_, _079995_, _079996_);
  not g_136121_(_079996_, _079997_);
  xor g_136122_(_079993_, _079994_, _079998_);
  or g_136123_(_078254_, _079998_, _079999_);
  not g_136124_(_079999_, _080001_);
  xor g_136125_(_078253_, _079998_, _080002_);
  or g_136126_(_078250_, _080002_, _080003_);
  not g_136127_(_080003_, _080004_);
  xor g_136128_(_078252_, _080002_, _080005_);
  not g_136129_(_080005_, _080006_);
  or g_136130_(_078249_, _080005_, _080007_);
  xor g_136131_(_078249_, _080005_, _080008_);
  xor g_136132_(_078249_, _080006_, _080009_);
  or g_136133_(_078248_, _080009_, _080010_);
  xor g_136134_(_078248_, _080008_, _080012_);
  not g_136135_(_080012_, _080013_);
  or g_136136_(_078247_, _080012_, _080014_);
  xor g_136137_(_078247_, _080013_, _080015_);
  not g_136138_(_080015_, _080016_);
  and g_136139_(_077208_, _077211_, _080017_);
  xor g_136140_(_080015_, _080017_, _080018_);
  xor g_136141_(_080016_, _080017_, _080019_);
  or g_136142_(_077213_, _080019_, _080020_);
  xor g_136143_(_077213_, _080018_, _080021_);
  or g_136144_(_074356_, _077212_, _080023_);
  not g_136145_(_080023_, _080024_);
  or g_136146_(_080021_, _080023_, _080025_);
  xor g_136147_(_080021_, _080023_, _080026_);
  xor g_136148_(_080021_, _080024_, _080027_);
  or g_136149_(_078246_, _080027_, _080028_);
  not g_136150_(_080028_, _080029_);
  xor g_136151_(_078246_, _080026_, _080030_);
  not g_136152_(_080030_, _080031_);
  or g_136153_(_078245_, _080030_, _080032_);
  xor g_136154_(_078245_, _080031_, _080034_);
  not g_136155_(_080034_, _080035_);
  or g_136156_(_074365_, _077219_, _080036_);
  or g_136157_(_080034_, _080036_, _080037_);
  xor g_136158_(_080034_, _080036_, _080038_);
  xor g_136159_(_080035_, _080036_, _080039_);
  or g_136160_(_077221_, _080039_, _080040_);
  xor g_136161_(_077221_, _080038_, _080041_);
  xor g_136162_(_077233_, _080041_, _080042_);
  xor g_136163_(_077234_, _080041_, _080043_);
  or g_136164_(_078244_, _080043_, _080045_);
  not g_136165_(_080045_, _080046_);
  xor g_136166_(_078244_, _080042_, _080047_);
  or g_136167_(_078243_, _080047_, _080048_);
  xor g_136168_(_078242_, _080047_, _080049_);
  not g_136169_(_080049_, _080050_);
  or g_136170_(_078241_, _080049_, _080051_);
  xor g_136171_(_078241_, _080050_, _080052_);
  or g_136172_(_078238_, _080052_, _080053_);
  xor g_136173_(_078239_, _080052_, _080054_);
  not g_136174_(_080054_, _080056_);
  and g_136175_(_077245_, _077248_, _080057_);
  xor g_136176_(_080056_, _080057_, _080058_);
  or g_136177_(_077254_, _080058_, _080059_);
  xor g_136178_(_077255_, _080058_, _080060_);
  and g_136179_(_077260_, _077265_, _080061_);
  not g_136180_(_080061_, _080062_);
  xor g_136181_(_080060_, _080062_, _080063_);
  and g_136182_(_077270_, _077277_, _080064_);
  and g_136183_(_080063_, _080064_, _080065_);
  or g_136184_(_077277_, _080063_, _080067_);
  or g_136185_(_077270_, _080063_, _080068_);
  and g_136186_(_080067_, _080068_, _080069_);
  not g_136187_(_080069_, _080070_);
  or g_136188_(_080065_, _080070_, _080071_);
  and g_136189_(_077272_, _077282_, _080072_);
  not g_136190_(_080072_, _080073_);
  or g_136191_(_080071_, _080072_, _080074_);
  xor g_136192_(_080071_, _080072_, _080075_);
  xor g_136193_(_080071_, _080073_, _080076_);
  or g_136194_(_077287_, _080076_, _080078_);
  xor g_136195_(_077287_, _080075_, _080079_);
  xor g_136196_(_077289_, _080079_, _080080_);
  or g_136197_(_077301_, _080080_, _080081_);
  xor g_136198_(_077301_, _080080_, _080082_);
  not g_136199_(_080082_, _080083_);
  or g_136200_(_077300_, _080083_, _080084_);
  not g_136201_(_080084_, _080085_);
  xor g_136202_(_077300_, _080082_, _080086_);
  not g_136203_(_080086_, _080087_);
  and g_136204_(_077294_, _077302_, _080089_);
  or g_136205_(_080086_, _080089_, _080090_);
  xor g_136206_(_080087_, _080089_, _080091_);
  not g_136207_(_080091_, _080092_);
  or g_136208_(_077305_, _080091_, _080093_);
  xor g_136209_(_077305_, _080091_, _080094_);
  xor g_136210_(_077305_, _080092_, _080095_);
  or g_136211_(_077309_, _080095_, _080096_);
  xor g_136212_(_077309_, _080094_, _080097_);
  or g_136213_(_077314_, _080097_, _080098_);
  not g_136214_(_080098_, _080100_);
  xor g_136215_(_077315_, _080097_, _080101_);
  or g_136216_(_074454_, _077311_, _080102_);
  or g_136217_(_080101_, _080102_, _080103_);
  xor g_136218_(_080101_, _080102_, _080104_);
  not g_136219_(_080104_, _080105_);
  and g_136220_(_078237_, _080104_, _080106_);
  or g_136221_(_078236_, _080105_, _080107_);
  xor g_136222_(_078236_, _080104_, _080108_);
  not g_136223_(_080108_, _080109_);
  and g_136224_(_077326_, _077329_, _080111_);
  xor g_136225_(_080109_, _080111_, _080112_);
  or g_136226_(_077332_, _080112_, _080113_);
  xor g_136227_(_077333_, _080112_, _080114_);
  or g_136228_(_074474_, _077330_, _080115_);
  or g_136229_(_080114_, _080115_, _080116_);
  xor g_136230_(_080114_, _080115_, _080117_);
  not g_136231_(_080117_, _080118_);
  or g_136232_(_078235_, _080118_, _080119_);
  xor g_136233_(_078235_, _080117_, _080120_);
  or g_136234_(_078234_, _080120_, _080122_);
  xor g_136235_(_078233_, _080120_, _080123_);
  or g_136236_(_078232_, _080123_, _080124_);
  xor g_136237_(_078231_, _080123_, _080125_);
  not g_136238_(_080125_, _080126_);
  or g_136239_(_077342_, _080125_, _080127_);
  xor g_136240_(_077342_, _080126_, _080128_);
  or g_136241_(_077346_, _080128_, _080129_);
  xor g_136242_(_077345_, _080128_, _080130_);
  or g_136243_(_077352_, _080130_, _080131_);
  xor g_136244_(_077353_, _080130_, _080133_);
  or g_136245_(_077348_, _080133_, _080134_);
  xor g_136246_(_077349_, _080133_, _080135_);
  not g_136247_(_080135_, _080136_);
  or g_136248_(_074503_, _077360_, _080137_);
  and g_136249_(_077358_, _080137_, _080138_);
  xor g_136250_(_080136_, _080138_, _080139_);
  or g_136251_(_078230_, _080139_, _080140_);
  xor g_136252_(_078230_, _080139_, _080141_);
  and g_136253_(_077371_, _080141_, _080142_);
  not g_136254_(_080142_, _080144_);
  xor g_136255_(_077371_, _080141_, _080145_);
  xor g_136256_(_077373_, _080141_, _080146_);
  or g_136257_(_077374_, _080146_, _080147_);
  xor g_136258_(_077374_, _080145_, _080148_);
  not g_136259_(_080148_, _080149_);
  and g_136260_(_077368_, _077375_, _080150_);
  xor g_136261_(_080149_, _080150_, _080151_);
  or g_136262_(_078227_, _080151_, _080152_);
  xor g_136263_(_078228_, _080151_, _080153_);
  not g_136264_(_080153_, _080155_);
  or g_136265_(_074523_, _077377_, _080156_);
  and g_136266_(_077381_, _080156_, _080157_);
  xor g_136267_(_080155_, _080157_, _080158_);
  not g_136268_(_080158_, _080159_);
  xor g_136269_(_078226_, _080159_, _080160_);
  not g_136270_(_080160_, _080161_);
  or g_136271_(_078224_, _080160_, _080162_);
  xor g_136272_(_078224_, _080160_, _080163_);
  xor g_136273_(_078224_, _080161_, _080164_);
  and g_136274_(_077395_, _077398_, _080166_);
  xor g_136275_(_080163_, _080166_, _080167_);
  or g_136276_(_077400_, _080167_, _080168_);
  not g_136277_(_080168_, _080169_);
  xor g_136278_(_077400_, _080167_, _080170_);
  xor g_136279_(_077401_, _080167_, _080171_);
  or g_136280_(_078223_, _080171_, _080172_);
  not g_136281_(_080172_, _080173_);
  xor g_136282_(_078223_, _080170_, _080174_);
  not g_136283_(_080174_, _080175_);
  or g_136284_(_078222_, _080174_, _080177_);
  xor g_136285_(_078222_, _080175_, _080178_);
  or g_136286_(_074556_, _077408_, _080179_);
  not g_136287_(_080179_, _080180_);
  or g_136288_(_080178_, _080179_, _080181_);
  xor g_136289_(_080178_, _080179_, _080182_);
  xor g_136290_(_080178_, _080180_, _080183_);
  or g_136291_(_078221_, _080183_, _080184_);
  not g_136292_(_080184_, _080185_);
  xor g_136293_(_078221_, _080182_, _080186_);
  or g_136294_(_077412_, _080186_, _080188_);
  not g_136295_(_080188_, _080189_);
  xor g_136296_(_077413_, _080186_, _080190_);
  or g_136297_(_074563_, _077410_, _080191_);
  or g_136298_(_080190_, _080191_, _080192_);
  not g_136299_(_080192_, _080193_);
  xor g_136300_(_080190_, _080191_, _080194_);
  not g_136301_(_080194_, _080195_);
  or g_136302_(_078220_, _080195_, _080196_);
  xor g_136303_(_078220_, _080194_, _080197_);
  not g_136304_(_080197_, _080199_);
  or g_136305_(_077419_, _080197_, _080200_);
  not g_136306_(_080200_, _080201_);
  xor g_136307_(_077419_, _080199_, _080202_);
  or g_136308_(_074573_, _077417_, _080203_);
  not g_136309_(_080203_, _080204_);
  or g_136310_(_080202_, _080203_, _080205_);
  xor g_136311_(_080202_, _080203_, _080206_);
  xor g_136312_(_080202_, _080204_, _080207_);
  or g_136313_(_078219_, _080207_, _080208_);
  xor g_136314_(_078219_, _080206_, _080210_);
  not g_136315_(_080210_, _080211_);
  and g_136316_(_077429_, _080211_, _080212_);
  or g_136317_(_077430_, _080210_, _080213_);
  xor g_136318_(_077429_, _080210_, _080214_);
  not g_136319_(_080214_, _080215_);
  and g_136320_(_077425_, _080215_, _080216_);
  xor g_136321_(_077425_, _080214_, _080217_);
  not g_136322_(_080217_, _080218_);
  and g_136323_(_077433_, _077434_, _080219_);
  xor g_136324_(_080218_, _080219_, _080221_);
  or g_136325_(_077436_, _080221_, _080222_);
  xor g_136326_(_077436_, _080221_, _080223_);
  not g_136327_(_080223_, _080224_);
  or g_136328_(_077444_, _080224_, _080225_);
  xor g_136329_(_077444_, _080223_, _080226_);
  or g_136330_(_077447_, _080226_, _080227_);
  xor g_136331_(_077448_, _080226_, _080228_);
  or g_136332_(_077454_, _080228_, _080229_);
  xor g_136333_(_077455_, _080228_, _080230_);
  or g_136334_(_077451_, _080230_, _080232_);
  xor g_136335_(_077451_, _080230_, _080233_);
  xor g_136336_(_077452_, _080230_, _080234_);
  and g_136337_(_077461_, _077464_, _080235_);
  xor g_136338_(_080233_, _080235_, _080236_);
  or g_136339_(_077467_, _080236_, _080237_);
  xor g_136340_(_077467_, _080236_, _080238_);
  not g_136341_(_080238_, _080239_);
  or g_136342_(_077470_, _080239_, _080240_);
  xor g_136343_(_077470_, _080238_, _080241_);
  or g_136344_(_077475_, _080241_, _080243_);
  xor g_136345_(_077476_, _080241_, _080244_);
  or g_136346_(_078216_, _080244_, _080245_);
  xor g_136347_(_078217_, _080244_, _080246_);
  not g_136348_(_080246_, _080247_);
  or g_136349_(_078215_, _080246_, _080248_);
  xor g_136350_(_078215_, _080247_, _080249_);
  or g_136351_(_077489_, _080249_, _080250_);
  xor g_136352_(_077489_, _080249_, _080251_);
  not g_136353_(_080251_, _080252_);
  and g_136354_(_077484_, _080251_, _080254_);
  or g_136355_(_077483_, _080252_, _080255_);
  xor g_136356_(_077483_, _080251_, _080256_);
  and g_136357_(_077496_, _077500_, _080257_);
  and g_136358_(_080256_, _080257_, _080258_);
  not g_136359_(_080258_, _080259_);
  or g_136360_(_077500_, _080256_, _080260_);
  or g_136361_(_077496_, _080256_, _080261_);
  and g_136362_(_080260_, _080261_, _080262_);
  not g_136363_(_080262_, _080263_);
  and g_136364_(_080259_, _080262_, _080265_);
  or g_136365_(_080258_, _080263_, _080266_);
  or g_136366_(_077502_, _080266_, _080267_);
  xor g_136367_(_077502_, _080265_, _080268_);
  or g_136368_(_077507_, _080268_, _080269_);
  xor g_136369_(_077506_, _080268_, _080270_);
  or g_136370_(_077509_, _080270_, _080271_);
  xor g_136371_(_077508_, _080270_, _080272_);
  or g_136372_(_074650_, _077512_, _080273_);
  not g_136373_(_080273_, _080274_);
  or g_136374_(_080272_, _080273_, _080276_);
  xor g_136375_(_080272_, _080273_, _080277_);
  xor g_136376_(_080272_, _080274_, _080278_);
  or g_136377_(_078214_, _080278_, _080279_);
  xor g_136378_(_078214_, _080277_, _080280_);
  not g_136379_(_080280_, _080281_);
  and g_136380_(_074657_, _077514_, _080282_);
  not g_136381_(_080282_, _080283_);
  and g_136382_(_080281_, _080282_, _080284_);
  or g_136383_(_080280_, _080283_, _080285_);
  xor g_136384_(_080280_, _080282_, _080287_);
  not g_136385_(_080287_, _080288_);
  or g_136386_(_078213_, _080287_, _080289_);
  xor g_136387_(_078213_, _080287_, _080290_);
  xor g_136388_(_078213_, _080288_, _080291_);
  and g_136389_(_078212_, _080290_, _080292_);
  or g_136390_(_078211_, _080291_, _080293_);
  xor g_136391_(_078211_, _080290_, _080294_);
  not g_136392_(_080294_, _080295_);
  or g_136393_(_078210_, _080294_, _080296_);
  xor g_136394_(_078210_, _080294_, _080298_);
  xor g_136395_(_078210_, _080295_, _080299_);
  and g_136396_(_077527_, _080298_, _080300_);
  or g_136397_(_077525_, _080299_, _080301_);
  and g_136398_(_077522_, _080298_, _080302_);
  or g_136399_(_077521_, _080299_, _080303_);
  and g_136400_(_080301_, _080303_, _080304_);
  or g_136401_(_080300_, _080302_, _080305_);
  and g_136402_(_077521_, _080299_, _080306_);
  and g_136403_(_077525_, _080306_, _080307_);
  or g_136404_(_080305_, _080307_, _080309_);
  or g_136405_(_078208_, _080309_, _080310_);
  xor g_136406_(_078208_, _080309_, _080311_);
  xor g_136407_(_078209_, _080309_, _080312_);
  or g_136408_(_078206_, _080312_, _080313_);
  xor g_136409_(_078206_, _080311_, _080314_);
  or g_136410_(_077535_, _080314_, _080315_);
  xor g_136411_(_077534_, _080314_, _080316_);
  or g_136412_(_077536_, _080316_, _080317_);
  xor g_136413_(_077538_, _080316_, _080318_);
  and g_136414_(_077541_, _077546_, _080320_);
  xor g_136415_(_080318_, _080320_, _080321_);
  not g_136416_(_080321_, _080322_);
  or g_136417_(_077545_, _080322_, _080323_);
  not g_136418_(_080323_, _080324_);
  xor g_136419_(_077545_, _080321_, _080325_);
  not g_136420_(_080325_, _080326_);
  or g_136421_(_074702_, _077554_, _080327_);
  and g_136422_(_077553_, _080327_, _080328_);
  xor g_136423_(_080326_, _080328_, _080329_);
  or g_136424_(_078205_, _080329_, _080331_);
  xor g_136425_(_078205_, _080329_, _080332_);
  not g_136426_(_080332_, _080333_);
  or g_136427_(_077558_, _080333_, _080334_);
  xor g_136428_(_077558_, _080332_, _080335_);
  or g_136429_(_074709_, _077556_, _080336_);
  not g_136430_(_080336_, _080337_);
  or g_136431_(_080335_, _080336_, _080338_);
  xor g_136432_(_080335_, _080337_, _080339_);
  not g_136433_(_080339_, _080340_);
  or g_136434_(_074715_, _077560_, _080342_);
  and g_136435_(_077564_, _080342_, _080343_);
  xor g_136436_(_080340_, _080343_, _080344_);
  or g_136437_(_077571_, _080344_, _080345_);
  xor g_136438_(_077571_, _080344_, _080346_);
  not g_136439_(_080346_, _080347_);
  and g_136440_(_077567_, _080346_, _080348_);
  or g_136441_(_077568_, _080347_, _080349_);
  xor g_136442_(_077568_, _080346_, _080350_);
  or g_136443_(_078203_, _080350_, _080351_);
  xor g_136444_(_078204_, _080350_, _080353_);
  or g_136445_(_074732_, _077575_, _080354_);
  not g_136446_(_080354_, _080355_);
  or g_136447_(_080353_, _080354_, _080356_);
  xor g_136448_(_080353_, _080354_, _080357_);
  xor g_136449_(_080353_, _080355_, _080358_);
  and g_136450_(_077579_, _080358_, _080359_);
  or g_136451_(_077580_, _080357_, _080360_);
  and g_136452_(_078201_, _080359_, _080361_);
  or g_136453_(_078202_, _080360_, _080362_);
  or g_136454_(_078201_, _080358_, _080364_);
  or g_136455_(_077579_, _080358_, _080365_);
  not g_136456_(_080365_, _080366_);
  and g_136457_(_080364_, _080365_, _080367_);
  not g_136458_(_080367_, _080368_);
  and g_136459_(_080362_, _080367_, _080369_);
  or g_136460_(_080361_, _080368_, _080370_);
  or g_136461_(_078200_, _080370_, _080371_);
  xor g_136462_(_078200_, _080369_, _080372_);
  or g_136463_(_077586_, _080372_, _080373_);
  not g_136464_(_080373_, _080375_);
  xor g_136465_(_077587_, _080372_, _080376_);
  or g_136466_(_077590_, _080376_, _080377_);
  xor g_136467_(_077591_, _080376_, _080378_);
  or g_136468_(_074751_, _077588_, _080379_);
  not g_136469_(_080379_, _080380_);
  or g_136470_(_080378_, _080379_, _080381_);
  xor g_136471_(_080378_, _080379_, _080382_);
  xor g_136472_(_080378_, _080380_, _080383_);
  or g_136473_(_078199_, _080383_, _080384_);
  xor g_136474_(_078199_, _080382_, _080386_);
  or g_136475_(_077598_, _080386_, _080387_);
  xor g_136476_(_077598_, _080386_, _080388_);
  xor g_136477_(_077597_, _080386_, _080389_);
  or g_136478_(_077599_, _080389_, _080390_);
  not g_136479_(_080390_, _080391_);
  xor g_136480_(_077599_, _080388_, _080392_);
  not g_136481_(_080392_, _080393_);
  or g_136482_(_077606_, _080392_, _080394_);
  xor g_136483_(_077606_, _080393_, _080395_);
  or g_136484_(_077610_, _080395_, _080397_);
  not g_136485_(_080397_, _080398_);
  xor g_136486_(_077610_, _080395_, _080399_);
  xor g_136487_(_077611_, _080395_, _080400_);
  or g_136488_(_074770_, _077608_, _080401_);
  or g_136489_(_080400_, _080401_, _080402_);
  xor g_136490_(_080399_, _080401_, _080403_);
  or g_136491_(_078198_, _080403_, _080404_);
  xor g_136492_(_078197_, _080403_, _080405_);
  or g_136493_(_077621_, _080405_, _080406_);
  not g_136494_(_080406_, _080408_);
  xor g_136495_(_077622_, _080405_, _080409_);
  or g_136496_(_077618_, _080409_, _080410_);
  xor g_136497_(_077619_, _080409_, _080411_);
  not g_136498_(_080411_, _080412_);
  or g_136499_(_077624_, _080411_, _080413_);
  xor g_136500_(_077624_, _080412_, _080414_);
  xor g_136501_(_077632_, _080414_, _080415_);
  xor g_136502_(_077633_, _080414_, _080416_);
  and g_136503_(_077638_, _080415_, _080417_);
  or g_136504_(_077637_, _080416_, _080419_);
  xor g_136505_(_077637_, _080415_, _080420_);
  or g_136506_(_077640_, _080420_, _080421_);
  xor g_136507_(_077641_, _080420_, _080422_);
  not g_136508_(_080422_, _080423_);
  or g_136509_(_077642_, _080422_, _080424_);
  xor g_136510_(_077642_, _080422_, _080425_);
  xor g_136511_(_077642_, _080423_, _080426_);
  xor g_136512_(_077651_, _080425_, _080427_);
  xor g_136513_(_077661_, _080427_, _080428_);
  not g_136514_(_080428_, _080430_);
  or g_136515_(_077666_, _080428_, _080431_);
  xor g_136516_(_077666_, _080430_, _080432_);
  or g_136517_(_074814_, _077663_, _080433_);
  not g_136518_(_080433_, _080434_);
  or g_136519_(_080432_, _080433_, _080435_);
  xor g_136520_(_080432_, _080433_, _080436_);
  xor g_136521_(_080432_, _080434_, _080437_);
  or g_136522_(_078195_, _080437_, _080438_);
  xor g_136523_(_078195_, _080436_, _080439_);
  not g_136524_(_080439_, _080441_);
  or g_136525_(_077673_, _080439_, _080442_);
  xor g_136526_(_077673_, _080441_, _080443_);
  or g_136527_(_074823_, _077671_, _080444_);
  not g_136528_(_080444_, _080445_);
  or g_136529_(_080443_, _080444_, _080446_);
  xor g_136530_(_080443_, _080445_, _080447_);
  not g_136531_(_080447_, _080448_);
  or g_136532_(_078194_, _080447_, _080449_);
  not g_136533_(_080449_, _080450_);
  xor g_136534_(_078194_, _080448_, _080452_);
  or g_136535_(_077678_, _080452_, _080453_);
  xor g_136536_(_077677_, _080452_, _080454_);
  not g_136537_(_080454_, _080455_);
  or g_136538_(_074833_, _077676_, _080456_);
  or g_136539_(_080454_, _080456_, _080457_);
  xor g_136540_(_080454_, _080456_, _080458_);
  xor g_136541_(_080455_, _080456_, _080459_);
  or g_136542_(_074835_, _077679_, _080460_);
  or g_136543_(_080459_, _080460_, _080461_);
  xor g_136544_(_080458_, _080460_, _080463_);
  or g_136545_(_077692_, _080463_, _080464_);
  not g_136546_(_080464_, _080465_);
  xor g_136547_(_077689_, _080463_, _080466_);
  and g_136548_(_077692_, _080466_, _080467_);
  or g_136549_(_080465_, _080467_, _080468_);
  or g_136550_(_077695_, _080468_, _080469_);
  xor g_136551_(_077696_, _080468_, _080470_);
  or g_136552_(_074849_, _077693_, _080471_);
  not g_136553_(_080471_, _080472_);
  or g_136554_(_080470_, _080471_, _080474_);
  xor g_136555_(_080470_, _080471_, _080475_);
  xor g_136556_(_080470_, _080472_, _080476_);
  or g_136557_(_078193_, _080476_, _080477_);
  xor g_136558_(_078193_, _080475_, _080478_);
  or g_136559_(_077701_, _080478_, _080479_);
  xor g_136560_(_077701_, _080478_, _080480_);
  xor g_136561_(_077703_, _080478_, _080481_);
  or g_136562_(_077706_, _080481_, _080482_);
  xor g_136563_(_077706_, _080480_, _080483_);
  or g_136564_(_077711_, _080483_, _080485_);
  xor g_136565_(_077712_, _080483_, _080486_);
  xor g_136566_(_077722_, _080486_, _080487_);
  or g_136567_(_078192_, _080487_, _080488_);
  xor g_136568_(_078192_, _080487_, _080489_);
  not g_136569_(_080489_, _080490_);
  or g_136570_(_078191_, _080490_, _080491_);
  xor g_136571_(_078191_, _080489_, _080492_);
  or g_136572_(_077733_, _080492_, _080493_);
  xor g_136573_(_077733_, _080492_, _080494_);
  xor g_136574_(_077734_, _080492_, _080496_);
  and g_136575_(_077732_, _080494_, _080497_);
  or g_136576_(_077731_, _080496_, _080498_);
  xor g_136577_(_077732_, _080494_, _080499_);
  xor g_136578_(_077731_, _080494_, _080500_);
  or g_136579_(_078190_, _080500_, _080501_);
  xor g_136580_(_078190_, _080499_, _080502_);
  or g_136581_(_074885_, _077737_, _080503_);
  not g_136582_(_080503_, _080504_);
  or g_136583_(_080502_, _080503_, _080505_);
  xor g_136584_(_080502_, _080504_, _080507_);
  not g_136585_(_080507_, _080508_);
  or g_136586_(_077740_, _080507_, _080509_);
  xor g_136587_(_077740_, _080507_, _080510_);
  xor g_136588_(_077740_, _080508_, _080511_);
  or g_136589_(_077745_, _080511_, _080512_);
  xor g_136590_(_077745_, _080510_, _080513_);
  not g_136591_(_080513_, _080514_);
  or g_136592_(_077749_, _080513_, _080515_);
  xor g_136593_(_077749_, _080514_, _080516_);
  not g_136594_(_080516_, _080518_);
  or g_136595_(_077752_, _080516_, _080519_);
  xor g_136596_(_077752_, _080516_, _080520_);
  xor g_136597_(_077752_, _080518_, _080521_);
  xor g_136598_(_077764_, _080520_, _080522_);
  not g_136599_(_080522_, _080523_);
  and g_136600_(_077769_, _080522_, _080524_);
  and g_136601_(_077772_, _080524_, _080525_);
  or g_136602_(_077772_, _080522_, _080526_);
  not g_136603_(_080526_, _080527_);
  and g_136604_(_077767_, _080523_, _080529_);
  not g_136605_(_080529_, _080530_);
  or g_136606_(_080527_, _080529_, _080531_);
  or g_136607_(_080525_, _080531_, _080532_);
  or g_136608_(_077774_, _080532_, _080533_);
  xor g_136609_(_077775_, _080532_, _080534_);
  or g_136610_(_077781_, _080534_, _080535_);
  xor g_136611_(_077782_, _080534_, _080536_);
  or g_136612_(_077785_, _080536_, _080537_);
  xor g_136613_(_077786_, _080536_, _080538_);
  or g_136614_(_074927_, _077783_, _080540_);
  or g_136615_(_080538_, _080540_, _080541_);
  xor g_136616_(_080538_, _080540_, _080542_);
  not g_136617_(_080542_, _080543_);
  and g_136618_(_078189_, _080542_, _080544_);
  or g_136619_(_078188_, _080543_, _080545_);
  xor g_136620_(_078188_, _080542_, _080546_);
  not g_136621_(_080546_, _080547_);
  and g_136622_(_077796_, _077799_, _080548_);
  xor g_136623_(_080547_, _080548_, _080549_);
  or g_136624_(_077803_, _080549_, _080551_);
  xor g_136625_(_077804_, _080549_, _080552_);
  not g_136626_(_080552_, _080553_);
  or g_136627_(_074948_, _077809_, _080554_);
  and g_136628_(_077807_, _080554_, _080555_);
  xor g_136629_(_080553_, _080555_, _080556_);
  or g_136630_(_078186_, _080556_, _080557_);
  xor g_136631_(_078187_, _080556_, _080558_);
  not g_136632_(_080558_, _080559_);
  and g_136633_(_077814_, _077817_, _080560_);
  and g_136634_(_080558_, _080560_, _080562_);
  or g_136635_(_077817_, _080558_, _080563_);
  not g_136636_(_080563_, _080564_);
  and g_136637_(_077813_, _080559_, _080565_);
  not g_136638_(_080565_, _080566_);
  or g_136639_(_080564_, _080565_, _080567_);
  or g_136640_(_080562_, _080567_, _080568_);
  not g_136641_(_080568_, _080569_);
  xor g_136642_(_077824_, _080569_, _080570_);
  or g_136643_(_078184_, _080570_, _080571_);
  not g_136644_(_080571_, _080573_);
  xor g_136645_(_078184_, _080570_, _080574_);
  not g_136646_(_080574_, _080575_);
  or g_136647_(_078183_, _080575_, _080576_);
  not g_136648_(_080576_, _080577_);
  xor g_136649_(_078183_, _080574_, _080578_);
  or g_136650_(_078182_, _080578_, _080579_);
  xor g_136651_(_078181_, _080578_, _080580_);
  not g_136652_(_080580_, _080581_);
  or g_136653_(_078180_, _080580_, _080582_);
  xor g_136654_(_078180_, _080581_, _080584_);
  not g_136655_(_080584_, _080585_);
  and g_136656_(_074982_, _077832_, _080586_);
  not g_136657_(_080586_, _080587_);
  and g_136658_(_080585_, _080586_, _080588_);
  or g_136659_(_080584_, _080587_, _080589_);
  xor g_136660_(_080584_, _080586_, _080590_);
  not g_136661_(_080590_, _080591_);
  or g_136662_(_077835_, _080590_, _080592_);
  not g_136663_(_080592_, _080593_);
  xor g_136664_(_077835_, _080590_, _080595_);
  xor g_136665_(_077835_, _080591_, _080596_);
  or g_136666_(_074990_, _077836_, _080597_);
  not g_136667_(_080597_, _080598_);
  or g_136668_(_080595_, _080598_, _080599_);
  or g_136669_(_074990_, _077833_, _080600_);
  or g_136670_(_080596_, _080600_, _080601_);
  not g_136671_(_080601_, _080602_);
  and g_136672_(_080599_, _080601_, _080603_);
  not g_136673_(_080603_, _080604_);
  or g_136674_(_078179_, _080604_, _080606_);
  xor g_136675_(_078179_, _080603_, _080607_);
  not g_136676_(_080607_, _080608_);
  or g_136677_(_077840_, _080607_, _080609_);
  xor g_136678_(_077840_, _080607_, _080610_);
  xor g_136679_(_077840_, _080608_, _080611_);
  or g_136680_(_078178_, _080611_, _080612_);
  xor g_136681_(_078178_, _080610_, _080613_);
  and g_136682_(_078177_, _080613_, _080614_);
  or g_136683_(_078177_, _080613_, _080615_);
  not g_136684_(_080615_, _080617_);
  xor g_136685_(_078177_, _080613_, _080618_);
  or g_136686_(_080614_, _080617_, _080619_);
  or g_136687_(_077844_, _080619_, _080620_);
  xor g_136688_(_077844_, _080618_, _080621_);
  or g_136689_(_077849_, _080621_, _080622_);
  xor g_136690_(_077848_, _080621_, _080623_);
  not g_136691_(_080623_, _080624_);
  or g_136692_(_075013_, _077846_, _080625_);
  or g_136693_(_080623_, _080625_, _080626_);
  xor g_136694_(_080623_, _080625_, _080628_);
  xor g_136695_(_080624_, _080625_, _080629_);
  or g_136696_(_075015_, _077850_, _080630_);
  or g_136697_(_080629_, _080630_, _080631_);
  xor g_136698_(_080628_, _080630_, _080632_);
  or g_136699_(_077854_, _080632_, _080633_);
  xor g_136700_(_077853_, _080632_, _080634_);
  or g_136701_(_077859_, _080634_, _080635_);
  xor g_136702_(_077858_, _080634_, _080636_);
  or g_136703_(_077862_, _080636_, _080637_);
  xor g_136704_(_077863_, _080636_, _080639_);
  or g_136705_(_075026_, _077860_, _080640_);
  not g_136706_(_080640_, _080641_);
  or g_136707_(_080639_, _080640_, _080642_);
  xor g_136708_(_080639_, _080640_, _080643_);
  xor g_136709_(_080639_, _080641_, _080644_);
  or g_136710_(_078176_, _080644_, _080645_);
  xor g_136711_(_078176_, _080643_, _080646_);
  or g_136712_(_077870_, _080646_, _080647_);
  xor g_136713_(_077870_, _080646_, _080648_);
  xor g_136714_(_077871_, _080646_, _080650_);
  or g_136715_(_078175_, _080650_, _080651_);
  xor g_136716_(_078175_, _080648_, _080652_);
  or g_136717_(_075038_, _077872_, _080653_);
  not g_136718_(_080653_, _080654_);
  or g_136719_(_080652_, _080653_, _080655_);
  xor g_136720_(_080652_, _080654_, _080656_);
  or g_136721_(_077874_, _080656_, _080657_);
  not g_136722_(_080657_, _080658_);
  or g_136723_(_077879_, _080656_, _080659_);
  xor g_136724_(_077879_, _080656_, _080661_);
  xor g_136725_(_077880_, _080656_, _080662_);
  and g_136726_(_077874_, _080662_, _080663_);
  or g_136727_(_077875_, _080661_, _080664_);
  and g_136728_(_080657_, _080664_, _080665_);
  or g_136729_(_080658_, _080663_, _080666_);
  or g_136730_(_078173_, _080666_, _080667_);
  xor g_136731_(_078173_, _080665_, _080668_);
  or g_136732_(_078171_, _080668_, _080669_);
  not g_136733_(_080669_, _080670_);
  xor g_136734_(_078172_, _080668_, _080672_);
  not g_136735_(_080672_, _080673_);
  and g_136736_(_077887_, _077890_, _080674_);
  xor g_136737_(_080673_, _080674_, _080675_);
  xor g_136738_(_080672_, _080674_, _080676_);
  or g_136739_(_077893_, _080675_, _080677_);
  xor g_136740_(_077893_, _080676_, _080678_);
  or g_136741_(_075067_, _077892_, _080679_);
  or g_136742_(_080678_, _080679_, _080680_);
  xor g_136743_(_080678_, _080679_, _080681_);
  not g_136744_(_080681_, _080683_);
  or g_136745_(_078170_, _080683_, _080684_);
  xor g_136746_(_078170_, _080681_, _080685_);
  or g_136747_(_077903_, _080685_, _080686_);
  xor g_136748_(_077903_, _080685_, _080687_);
  not g_136749_(_080687_, _080688_);
  or g_136750_(_077902_, _080688_, _080689_);
  xor g_136751_(_077902_, _080687_, _080690_);
  and g_136752_(_077906_, _077909_, _080691_);
  xor g_136753_(_080690_, _080691_, _080692_);
  not g_136754_(_080692_, _080694_);
  or g_136755_(_077914_, _080694_, _080695_);
  not g_136756_(_080695_, _080696_);
  or g_136757_(_077917_, _080694_, _080697_);
  xor g_136758_(_077917_, _080692_, _080698_);
  and g_136759_(_077914_, _080698_, _080699_);
  or g_136760_(_080696_, _080699_, _080700_);
  or g_136761_(_078168_, _080700_, _080701_);
  xor g_136762_(_078169_, _080700_, _080702_);
  or g_136763_(_075094_, _077918_, _080703_);
  not g_136764_(_080703_, _080705_);
  or g_136765_(_080702_, _080703_, _080706_);
  not g_136766_(_080706_, _080707_);
  xor g_136767_(_080702_, _080705_, _080708_);
  or g_136768_(_077923_, _080708_, _080709_);
  not g_136769_(_080709_, _080710_);
  xor g_136770_(_077924_, _080708_, _080711_);
  or g_136771_(_077927_, _080711_, _080712_);
  xor g_136772_(_077928_, _080711_, _080713_);
  or g_136773_(_077931_, _080713_, _080714_);
  xor g_136774_(_077931_, _080713_, _080716_);
  not g_136775_(_080716_, _080717_);
  and g_136776_(_077935_, _077937_, _080718_);
  not g_136777_(_080718_, _080719_);
  xor g_136778_(_080716_, _080719_, _080720_);
  xor g_136779_(_080716_, _080718_, _080721_);
  or g_136780_(_078167_, _080721_, _080722_);
  xor g_136781_(_078167_, _080720_, _080723_);
  or g_136782_(_078166_, _080723_, _080724_);
  not g_136783_(_080724_, _080725_);
  xor g_136784_(_078165_, _080723_, _080727_);
  not g_136785_(_080727_, _080728_);
  and g_136786_(_077943_, _080728_, _080729_);
  not g_136787_(_080729_, _080730_);
  xor g_136788_(_077943_, _080727_, _080731_);
  or g_136789_(_075123_, _077941_, _080732_);
  and g_136790_(_080731_, _080732_, _080733_);
  or g_136791_(_080731_, _080732_, _080734_);
  not g_136792_(_080734_, _080735_);
  xor g_136793_(_080731_, _080732_, _080736_);
  or g_136794_(_080733_, _080735_, _080738_);
  or g_136795_(_078164_, _080738_, _080739_);
  xor g_136796_(_078164_, _080736_, _080740_);
  or g_136797_(_078162_, _080740_, _080741_);
  xor g_136798_(_078161_, _080740_, _080742_);
  and g_136799_(_075134_, _077946_, _080743_);
  not g_136800_(_080743_, _080744_);
  or g_136801_(_080742_, _080744_, _080745_);
  xor g_136802_(_080742_, _080743_, _080746_);
  or g_136803_(_077949_, _080746_, _080747_);
  xor g_136804_(_077950_, _080746_, _080749_);
  or g_136805_(_077952_, _080749_, _080750_);
  xor g_136806_(_077953_, _080749_, _080751_);
  or g_136807_(_077954_, _080751_, _080752_);
  not g_136808_(_080752_, _080753_);
  xor g_136809_(_077954_, _080751_, _080754_);
  not g_136810_(_080754_, _080755_);
  or g_136811_(_077959_, _080755_, _080756_);
  not g_136812_(_080756_, _080757_);
  xor g_136813_(_077959_, _080754_, _080758_);
  xor g_136814_(_077969_, _080758_, _080760_);
  not g_136815_(_080760_, _080761_);
  and g_136816_(_077971_, _077975_, _080762_);
  xor g_136817_(_080760_, _080762_, _080763_);
  or g_136818_(_078160_, _080763_, _080764_);
  not g_136819_(_080764_, _080765_);
  xor g_136820_(_078160_, _080763_, _080766_);
  not g_136821_(_080766_, _080767_);
  or g_136822_(_078159_, _080767_, _080768_);
  xor g_136823_(_078159_, _080766_, _080769_);
  not g_136824_(_080769_, _080771_);
  or g_136825_(_077982_, _080769_, _080772_);
  xor g_136826_(_077982_, _080769_, _080773_);
  xor g_136827_(_077982_, _080771_, _080774_);
  or g_136828_(_075172_, _077981_, _080775_);
  or g_136829_(_080774_, _080775_, _080776_);
  xor g_136830_(_080773_, _080775_, _080777_);
  not g_136831_(_080777_, _080778_);
  and g_136832_(_078157_, _080778_, _080779_);
  or g_136833_(_078158_, _080777_, _080780_);
  xor g_136834_(_078157_, _080777_, _080782_);
  or g_136835_(_077994_, _080782_, _080783_);
  not g_136836_(_080783_, _080784_);
  xor g_136837_(_077993_, _080782_, _080785_);
  or g_136838_(_077989_, _080785_, _080786_);
  xor g_136839_(_077990_, _080785_, _080787_);
  or g_136840_(_077997_, _080787_, _080788_);
  xor g_136841_(_077998_, _080787_, _080789_);
  or g_136842_(_078002_, _080789_, _080790_);
  not g_136843_(_080790_, _080791_);
  xor g_136844_(_078002_, _080789_, _080793_);
  not g_136845_(_080793_, _080794_);
  and g_136846_(_078007_, _080793_, _080795_);
  or g_136847_(_078006_, _080794_, _080796_);
  xor g_136848_(_078006_, _080793_, _080797_);
  or g_136849_(_078155_, _080797_, _080798_);
  xor g_136850_(_078156_, _080797_, _080799_);
  not g_136851_(_080799_, _080800_);
  and g_136852_(_078154_, _080800_, _080801_);
  not g_136853_(_080801_, _080802_);
  xor g_136854_(_078154_, _080799_, _080804_);
  or g_136855_(_078015_, _080804_, _080805_);
  not g_136856_(_080805_, _080806_);
  xor g_136857_(_078015_, _080804_, _080807_);
  xor g_136858_(_078016_, _080807_, _080808_);
  and g_136859_(_078018_, _080808_, _080809_);
  or g_136860_(_078018_, _080804_, _080810_);
  not g_136861_(_080810_, _080811_);
  or g_136862_(_080809_, _080811_, _080812_);
  or g_136863_(_078023_, _080812_, _080813_);
  xor g_136864_(_078024_, _080812_, _080815_);
  or g_136865_(_078020_, _080815_, _080816_);
  not g_136866_(_080816_, _080817_);
  xor g_136867_(_078022_, _080815_, _080818_);
  or g_136868_(_075220_, _078027_, _080819_);
  not g_136869_(_080819_, _080820_);
  or g_136870_(_080818_, _080819_, _080821_);
  not g_136871_(_080821_, _080822_);
  xor g_136872_(_080818_, _080820_, _080823_);
  or g_136873_(_075223_, _078027_, _080824_);
  not g_136874_(_080824_, _080826_);
  or g_136875_(_080823_, _080824_, _080827_);
  xor g_136876_(_080823_, _080826_, _080828_);
  not g_136877_(_080828_, _080829_);
  or g_136878_(_078031_, _080828_, _080830_);
  not g_136879_(_080830_, _080831_);
  xor g_136880_(_078031_, _080828_, _080832_);
  xor g_136881_(_078031_, _080829_, _080833_);
  or g_136882_(_078035_, _080833_, _080834_);
  xor g_136883_(_078035_, _080832_, _080835_);
  or g_136884_(_075233_, _078033_, _080837_);
  not g_136885_(_080837_, _080838_);
  or g_136886_(_080835_, _080837_, _080839_);
  xor g_136887_(_080835_, _080838_, _080840_);
  or g_136888_(_075235_, _078037_, _080841_);
  not g_136889_(_080841_, _080842_);
  or g_136890_(_080840_, _080841_, _080843_);
  not g_136891_(_080843_, _080844_);
  xor g_136892_(_080840_, _080842_, _080845_);
  not g_136893_(_080845_, _080846_);
  and g_136894_(_078042_, _078046_, _080848_);
  xor g_136895_(_080846_, _080848_, _080849_);
  or g_136896_(_078050_, _080849_, _080850_);
  not g_136897_(_080850_, _080851_);
  xor g_136898_(_078050_, _080849_, _080852_);
  xor g_136899_(_078051_, _080849_, _080853_);
  and g_136900_(_078055_, _078058_, _080854_);
  xor g_136901_(_080852_, _080854_, _080855_);
  not g_136902_(_080855_, _080856_);
  and g_136903_(_078061_, _078066_, _080857_);
  xor g_136904_(_080856_, _080857_, _080859_);
  or g_136905_(_078063_, _080859_, _080860_);
  xor g_136906_(_078063_, _080859_, _080861_);
  not g_136907_(_080861_, _080862_);
  or g_136908_(_078072_, _080862_, _080863_);
  xor g_136909_(_078072_, _080861_, _080864_);
  and g_136910_(_078079_, _080864_, _080865_);
  and g_136911_(_078083_, _080865_, _080866_);
  not g_136912_(_080866_, _080867_);
  or g_136913_(_078083_, _080864_, _080868_);
  not g_136914_(_080868_, _080870_);
  or g_136915_(_078079_, _080864_, _080871_);
  not g_136916_(_080871_, _080872_);
  and g_136917_(_080868_, _080871_, _080873_);
  not g_136918_(_080873_, _080874_);
  and g_136919_(_080867_, _080873_, _080875_);
  or g_136920_(_080866_, _080874_, _080876_);
  or g_136921_(_078086_, _080876_, _080877_);
  xor g_136922_(_078086_, _080876_, _080878_);
  xor g_136923_(_078086_, _080875_, _080879_);
  or g_136924_(_075285_, _078084_, _080881_);
  or g_136925_(_080879_, _080881_, _080882_);
  xor g_136926_(_080878_, _080881_, _080883_);
  or g_136927_(_075288_, _078088_, _080884_);
  not g_136928_(_080884_, _080885_);
  or g_136929_(_080883_, _080884_, _080886_);
  xor g_136930_(_080883_, _080885_, _080887_);
  not g_136931_(_080887_, _080888_);
  or g_136932_(_075295_, _078091_, _080889_);
  and g_136933_(_078093_, _080889_, _080890_);
  xor g_136934_(_080888_, _080890_, _080892_);
  or g_136935_(_078151_, _080892_, _080893_);
  xor g_136936_(_078151_, _080892_, _080894_);
  not g_136937_(_080894_, _080895_);
  xor g_136938_(_078103_, _080894_, _080896_);
  not g_136939_(_080896_, _080897_);
  or g_136940_(_078106_, _080896_, _080898_);
  xor g_136941_(_078106_, _080897_, _080899_);
  not g_136942_(_080899_, _080900_);
  and g_136943_(_078110_, _078112_, _080901_);
  xor g_136944_(_080900_, _080901_, _080903_);
  or g_136945_(_078116_, _080903_, _080904_);
  xor g_136946_(_078117_, _080903_, _080905_);
  or g_136947_(_075323_, _078115_, _080906_);
  and g_136948_(_080905_, _080906_, _080907_);
  or g_136949_(_080905_, _080906_, _080908_);
  not g_136950_(_080908_, _080909_);
  or g_136951_(_080907_, _080909_, _080910_);
  or g_136952_(_075326_, _078118_, _080911_);
  or g_136953_(_080910_, _080911_, _080912_);
  not g_136954_(_080912_, _080914_);
  xor g_136955_(_080910_, _080911_, _080915_);
  not g_136956_(_080915_, _080916_);
  and g_136957_(_078150_, _080915_, _080917_);
  or g_136958_(_078149_, _080916_, _080918_);
  xor g_136959_(_078149_, _080915_, _080919_);
  or g_136960_(_075333_, _078121_, _080920_);
  and g_136961_(_078125_, _080920_, _080921_);
  xor g_136962_(_080919_, _080921_, _080922_);
  not g_136963_(_080922_, _080923_);
  or g_136964_(_078128_, _080923_, _080925_);
  xor g_136965_(_078128_, _080922_, _080926_);
  not g_136966_(_080926_, _080927_);
  or g_136967_(_078130_, _080926_, _080928_);
  xor g_136968_(_078130_, _080927_, _080929_);
  not g_136969_(_080929_, _080930_);
  or g_136970_(_078136_, _080929_, _080931_);
  xor g_136971_(_078136_, _080930_, _080932_);
  or g_136972_(_078139_, _080932_, _080933_);
  xor g_136973_(_078139_, _080932_, _080934_);
  not g_136974_(_080934_, _080936_);
  or g_136975_(_078145_, _080936_, _080937_);
  not g_136976_(_080937_, _080938_);
  xor g_136977_(_078145_, _080934_, _080939_);
  or g_136978_(_078148_, _080939_, _080940_);
  xor g_136979_(_078148_, _080939_, out[962]);
  or g_136980_(_078125_, _080919_, _080941_);
  or g_136981_(_080919_, _080920_, _080942_);
  or g_136982_(_078107_, _080896_, _080943_);
  or g_136983_(_075313_, _080943_, _080944_);
  or g_136984_(_075311_, _080943_, _080946_);
  or g_136985_(_078101_, _080895_, _080947_);
  not g_136986_(_080947_, _080948_);
  or g_136987_(_080887_, _080889_, _080949_);
  not g_136988_(_080949_, _080950_);
  or g_136989_(_078093_, _080887_, _080951_);
  and g_136990_(_080886_, _080951_, _080952_);
  or g_136991_(_078066_, _080855_, _080953_);
  or g_136992_(_078061_, _080855_, _080954_);
  not g_136993_(_080954_, _080955_);
  and g_136994_(_078059_, _080852_, _080957_);
  not g_136995_(_080957_, _080958_);
  or g_136996_(_078055_, _080853_, _080959_);
  not g_136997_(_080959_, _080960_);
  or g_136998_(_078046_, _080845_, _080961_);
  not g_136999_(_080961_, _080962_);
  or g_137000_(_078041_, _080845_, _080963_);
  or g_137001_(_075241_, _080963_, _080964_);
  or g_137002_(_075237_, _080963_, _080965_);
  and g_137003_(_080790_, _080796_, _080966_);
  not g_137004_(_080966_, _080968_);
  and g_137005_(_077976_, _080760_, _080969_);
  not g_137006_(_080969_, _080970_);
  and g_137007_(_077972_, _080760_, _080971_);
  or g_137008_(_077971_, _080761_, _080972_);
  and g_137009_(_077962_, _080754_, _080973_);
  or g_137010_(_077961_, _080755_, _080974_);
  or g_137011_(_077964_, _080758_, _080975_);
  and g_137012_(_077938_, _080716_, _080976_);
  not g_137013_(_080976_, _080977_);
  or g_137014_(_077935_, _080717_, _080979_);
  not g_137015_(_080979_, _080980_);
  or g_137016_(_077909_, _080690_, _080981_);
  or g_137017_(_077906_, _080690_, _080982_);
  or g_137018_(_077890_, _080672_, _080983_);
  or g_137019_(_077885_, _080672_, _080984_);
  or g_137020_(_077886_, _080672_, _080985_);
  not g_137021_(_080985_, _080986_);
  or g_137022_(_080552_, _080554_, _080987_);
  or g_137023_(_077799_, _080546_, _080988_);
  or g_137024_(_077794_, _080546_, _080990_);
  not g_137025_(_080990_, _080991_);
  or g_137026_(_077755_, _080516_, _080992_);
  or g_137027_(_077716_, _080486_, _080993_);
  or g_137028_(_077720_, _080486_, _080994_);
  or g_137029_(_077685_, _080463_, _080995_);
  or g_137030_(_077686_, _080463_, _080996_);
  not g_137031_(_080996_, _080997_);
  or g_137032_(_077656_, _080427_, _080998_);
  or g_137033_(_077655_, _080426_, _080999_);
  or g_137034_(_077649_, _080426_, _081001_);
  or g_137035_(_077630_, _080411_, _081002_);
  not g_137036_(_081002_, _081003_);
  or g_137037_(_077631_, _080414_, _081004_);
  or g_137038_(_077564_, _080339_, _081005_);
  or g_137039_(_080325_, _080327_, _081006_);
  or g_137040_(_077551_, _080325_, _081007_);
  or g_137041_(_077552_, _080325_, _081008_);
  or g_137042_(_077546_, _080318_, _081009_);
  or g_137043_(_077541_, _080318_, _081010_);
  and g_137044_(_080248_, _080250_, _081012_);
  and g_137045_(_080243_, _080245_, _081013_);
  or g_137046_(_077464_, _080234_, _081014_);
  or g_137047_(_077433_, _080217_, _081015_);
  or g_137048_(_077434_, _080217_, _081016_);
  or g_137049_(_077398_, _080164_, _081017_);
  or g_137050_(_077395_, _080164_, _081018_);
  or g_137051_(_077386_, _080158_, _081019_);
  not g_137052_(_081019_, _081020_);
  or g_137053_(_077387_, _080158_, _081021_);
  or g_137054_(_077381_, _080153_, _081023_);
  or g_137055_(_077375_, _080148_, _081024_);
  not g_137056_(_081024_, _081025_);
  or g_137057_(_077358_, _080135_, _081026_);
  or g_137058_(_077329_, _080108_, _081027_);
  or g_137059_(_077322_, _080108_, _081028_);
  and g_137060_(_077324_, _080109_, _081029_);
  and g_137061_(_080098_, _080103_, _081030_);
  and g_137062_(_080093_, _080096_, _081031_);
  and g_137063_(_077289_, _080075_, _081032_);
  or g_137064_(_077288_, _080076_, _081034_);
  or g_137065_(_077265_, _080060_, _081035_);
  and g_137066_(_080068_, _081035_, _081036_);
  not g_137067_(_081036_, _081037_);
  or g_137068_(_077248_, _080054_, _081038_);
  or g_137069_(_077242_, _080054_, _081039_);
  or g_137070_(_077243_, _080054_, _081040_);
  and g_137071_(_080053_, _081040_, _081041_);
  or g_137072_(_077224_, _080039_, _081042_);
  or g_137073_(_077227_, _080041_, _081043_);
  or g_137074_(_077211_, _080015_, _081045_);
  or g_137075_(_077189_, _079980_, _081046_);
  or g_137076_(_077180_, _079980_, _081047_);
  or g_137077_(_077178_, _079974_, _081048_);
  or g_137078_(_077136_, _079926_, _081049_);
  or g_137079_(_079926_, _079928_, _081050_);
  or g_137080_(_077114_, _079910_, _081051_);
  or g_137081_(_079888_, _079889_, _081052_);
  or g_137082_(_077093_, _079888_, _081053_);
  and g_137083_(_077077_, _079878_, _081054_);
  or g_137084_(_077078_, _079880_, _081056_);
  or g_137085_(_077052_, _079864_, _081057_);
  or g_137086_(_077046_, _079862_, _081058_);
  or g_137087_(_074168_, _081058_, _081059_);
  or g_137088_(_079844_, _079847_, _081060_);
  or g_137089_(_077035_, _079844_, _081061_);
  or g_137090_(_077025_, _079842_, _081062_);
  or g_137091_(_077028_, _079842_, _081063_);
  not g_137092_(_081063_, _081064_);
  or g_137093_(_077023_, _079841_, _081065_);
  not g_137094_(_081065_, _081067_);
  or g_137095_(_079827_, _079829_, _081068_);
  and g_137096_(_079833_, _081068_, _081069_);
  or g_137097_(_079806_, _079807_, _081070_);
  not g_137098_(_081070_, _081071_);
  or g_137099_(_076962_, _079785_, _081072_);
  not g_137100_(_081072_, _081073_);
  or g_137101_(_076959_, _079785_, _081074_);
  not g_137102_(_081074_, _081075_);
  and g_137103_(_079775_, _079777_, _081076_);
  or g_137104_(_076940_, _079759_, _081078_);
  not g_137105_(_081078_, _081079_);
  or g_137106_(_076934_, _079756_, _081080_);
  or g_137107_(_074052_, _081080_, _081081_);
  not g_137108_(_081081_, _081082_);
  or g_137109_(_074048_, _081080_, _081083_);
  or g_137110_(_076925_, _079750_, _081084_);
  or g_137111_(_076920_, _079750_, _081085_);
  or g_137112_(_076911_, _079748_, _081086_);
  or g_137113_(_076915_, _079748_, _081087_);
  or g_137114_(_076908_, _079745_, _081089_);
  or g_137115_(_076904_, _079745_, _081090_);
  not g_137116_(_081090_, _081091_);
  or g_137117_(_076874_, _079705_, _081092_);
  not g_137118_(_081092_, _081093_);
  or g_137119_(_076868_, _079705_, _081094_);
  or g_137120_(_076832_, _079647_, _081095_);
  and g_137121_(_076821_, _079649_, _081096_);
  not g_137122_(_081096_, _081097_);
  and g_137123_(_076824_, _079649_, _081098_);
  not g_137124_(_081098_, _081100_);
  or g_137125_(_076810_, _079646_, _081101_);
  not g_137126_(_081101_, _081102_);
  or g_137127_(_076815_, _079646_, _081103_);
  or g_137128_(_076787_, _079631_, _081104_);
  and g_137129_(_076753_, _079611_, _081105_);
  or g_137130_(_076752_, _079612_, _081106_);
  or g_137131_(_076749_, _079612_, _081107_);
  or g_137132_(_073866_, _081107_, _081108_);
  not g_137133_(_081108_, _081109_);
  and g_137134_(_079599_, _079601_, _081111_);
  not g_137135_(_081111_, _081112_);
  or g_137136_(_076716_, _079570_, _081113_);
  not g_137137_(_081113_, _081114_);
  or g_137138_(_076713_, _079570_, _081115_);
  not g_137139_(_081115_, _081116_);
  and g_137140_(_079522_, _079524_, _081117_);
  or g_137141_(_076652_, _079498_, _081118_);
  or g_137142_(_076647_, _079498_, _081119_);
  or g_137143_(_076648_, _079498_, _081120_);
  or g_137144_(_076633_, _079486_, _081122_);
  and g_137145_(_079490_, _081122_, _081123_);
  or g_137146_(_076612_, _079463_, _081124_);
  not g_137147_(_081124_, _081125_);
  or g_137148_(_076610_, _079463_, _081126_);
  and g_137149_(_079454_, _081126_, _081127_);
  or g_137150_(_076598_, _079451_, _081128_);
  not g_137151_(_081128_, _081129_);
  or g_137152_(_076586_, _079445_, _081130_);
  not g_137153_(_081130_, _081131_);
  or g_137154_(_079430_, _079432_, _081133_);
  or g_137155_(_076556_, _079414_, _081134_);
  not g_137156_(_081134_, _081135_);
  or g_137157_(_076551_, _079414_, _081136_);
  or g_137158_(_076542_, _079409_, _081137_);
  or g_137159_(_073650_, _081137_, _081138_);
  or g_137160_(_073647_, _081137_, _081139_);
  not g_137161_(_081139_, _081140_);
  or g_137162_(_076512_, _079364_, _081141_);
  not g_137163_(_081141_, _081142_);
  or g_137164_(_076507_, _079364_, _081144_);
  and g_137165_(_079360_, _079363_, _081145_);
  or g_137166_(_076479_, _079338_, _081146_);
  or g_137167_(_076455_, _079310_, _081147_);
  not g_137168_(_081147_, _081148_);
  or g_137169_(_076420_, _079270_, _081149_);
  or g_137170_(_076418_, _079270_, _081150_);
  not g_137171_(_081150_, _081151_);
  or g_137172_(_076409_, _079267_, _081152_);
  not g_137173_(_081152_, _081153_);
  or g_137174_(_076401_, _079267_, _081155_);
  not g_137175_(_081155_, _081156_);
  or g_137176_(_076396_, _079265_, _081157_);
  or g_137177_(_076379_, _079258_, _081158_);
  or g_137178_(_073481_, _081158_, _081159_);
  not g_137179_(_081159_, _081160_);
  or g_137180_(_073477_, _081158_, _081161_);
  or g_137181_(_076366_, _079244_, _081162_);
  or g_137182_(_076362_, _079242_, _081163_);
  or g_137183_(_076341_, _079215_, _081164_);
  not g_137184_(_081164_, _081166_);
  or g_137185_(_076337_, _079215_, _081167_);
  and g_137186_(_079201_, _079206_, _081168_);
  and g_137187_(_079182_, _079188_, _081169_);
  or g_137188_(_076268_, _079119_, _081170_);
  not g_137189_(_081170_, _081171_);
  and g_137190_(_076262_, _079116_, _081172_);
  or g_137191_(_076260_, _079117_, _081173_);
  or g_137192_(_076258_, _079117_, _081174_);
  or g_137193_(_076237_, _079096_, _081175_);
  or g_137194_(_076202_, _079061_, _081177_);
  not g_137195_(_081177_, _081178_);
  or g_137196_(_076193_, _079061_, _081179_);
  or g_137197_(_076194_, _079061_, _081180_);
  not g_137198_(_081180_, _081181_);
  or g_137199_(_073255_, _076185_, _081182_);
  or g_137200_(_079058_, _081182_, _081183_);
  not g_137201_(_081183_, _081184_);
  and g_137202_(_076172_, _079047_, _081185_);
  or g_137203_(_076171_, _079048_, _081186_);
  or g_137204_(_076168_, _079048_, _081188_);
  or g_137205_(_073238_, _081188_, _081189_);
  not g_137206_(_081189_, _081190_);
  or g_137207_(_076160_, _079044_, _081191_);
  not g_137208_(_081191_, _081192_);
  or g_137209_(_076167_, _079044_, _081193_);
  or g_137210_(_076157_, _079044_, _081194_);
  not g_137211_(_081194_, _081195_);
  and g_137212_(_079040_, _079042_, _081196_);
  or g_137213_(_076126_, _079031_, _081197_);
  or g_137214_(_076068_, _078962_, _081199_);
  or g_137215_(_076069_, _078967_, _081200_);
  not g_137216_(_081200_, _081201_);
  or g_137217_(_076015_, _078931_, _081202_);
  not g_137218_(_081202_, _081203_);
  and g_137219_(_076012_, _078928_, _081204_);
  or g_137220_(_076011_, _078929_, _081205_);
  or g_137221_(_075991_, _078901_, _081206_);
  not g_137222_(_081206_, _081207_);
  or g_137223_(_075992_, _078903_, _081208_);
  not g_137224_(_081208_, _081210_);
  and g_137225_(_073031_, _075961_, _081211_);
  not g_137226_(_081211_, _081212_);
  or g_137227_(_078869_, _081212_, _081213_);
  not g_137228_(_081213_, _081214_);
  or g_137229_(_075955_, _078859_, _081215_);
  or g_137230_(_075947_, _078859_, _081216_);
  or g_137231_(_072993_, _075924_, _081217_);
  or g_137232_(_078835_, _081217_, _081218_);
  not g_137233_(_081218_, _081219_);
  or g_137234_(_072990_, _075924_, _081221_);
  or g_137235_(_078835_, _081221_, _081222_);
  not g_137236_(_081222_, _081223_);
  or g_137237_(_075911_, _078819_, _081224_);
  not g_137238_(_081224_, _081225_);
  or g_137239_(_075857_, _078775_, _081226_);
  or g_137240_(_075850_, _078772_, _081227_);
  or g_137241_(_072926_, _081227_, _081228_);
  not g_137242_(_081228_, _081229_);
  or g_137243_(_075828_, _078753_, _081230_);
  not g_137244_(_081230_, _081232_);
  or g_137245_(_075822_, _078751_, _081233_);
  or g_137246_(_072895_, _081233_, _081234_);
  or g_137247_(_075780_, _078719_, _081235_);
  or g_137248_(_072857_, _081235_, _081236_);
  or g_137249_(_072854_, _081235_, _081237_);
  or g_137250_(_075775_, _078704_, _081238_);
  or g_137251_(_075767_, _078704_, _081239_);
  not g_137252_(_081239_, _081240_);
  and g_137253_(_075759_, _078692_, _081241_);
  or g_137254_(_075758_, _078693_, _081243_);
  or g_137255_(_078688_, _078689_, _081244_);
  or g_137256_(_075717_, _078673_, _081245_);
  or g_137257_(_072798_, _081245_, _081246_);
  or g_137258_(_075709_, _078673_, _081247_);
  or g_137259_(_075713_, _078671_, _081248_);
  or g_137260_(_075691_, _078656_, _081249_);
  or g_137261_(_075688_, _078656_, _081250_);
  not g_137262_(_081250_, _081251_);
  or g_137263_(_075686_, _078653_, _081252_);
  or g_137264_(_075684_, _078653_, _081254_);
  not g_137265_(_081254_, _081255_);
  or g_137266_(_075674_, _078643_, _081256_);
  not g_137267_(_081256_, _081257_);
  or g_137268_(_075670_, _078643_, _081258_);
  or g_137269_(_072754_, _081258_, _081259_);
  not g_137270_(_081259_, _081260_);
  or g_137271_(_075659_, _078620_, _081261_);
  not g_137272_(_081261_, _081262_);
  or g_137273_(_075648_, _078615_, _081263_);
  or g_137274_(_075625_, _078593_, _081265_);
  not g_137275_(_081265_, _081266_);
  or g_137276_(_075622_, _078593_, _081267_);
  and g_137277_(_078566_, _078568_, _081268_);
  not g_137278_(_081268_, _081269_);
  or g_137279_(_075580_, _078556_, _081270_);
  or g_137280_(_075555_, _078540_, _081271_);
  or g_137281_(_075552_, _078540_, _081272_);
  and g_137282_(_078525_, _078529_, _081273_);
  and g_137283_(_078511_, _078513_, _081274_);
  and g_137284_(_078411_, _078417_, _081276_);
  and g_137285_(_078408_, _081276_, _081277_);
  and g_137286_(_078420_, _078423_, _081278_);
  and g_137287_(_081277_, _081278_, _081279_);
  and g_137288_(_078426_, _078431_, _081280_);
  and g_137289_(_081279_, _081280_, _081281_);
  and g_137290_(_078435_, _081281_, _081282_);
  and g_137291_(_078442_, _078445_, _081283_);
  or g_137292_(_081282_, _081283_, _081284_);
  and g_137293_(_078459_, _078464_, _081285_);
  and g_137294_(_078453_, _078456_, _081287_);
  or g_137295_(_078439_, _081282_, _081288_);
  xor g_137296_(_078439_, _081282_, _081289_);
  and g_137297_(_078442_, _078450_, _081290_);
  xor g_137298_(_081289_, _081290_, _081291_);
  not g_137299_(_081291_, _081292_);
  or g_137300_(_081287_, _081291_, _081293_);
  xor g_137301_(_081287_, _081291_, _081294_);
  xor g_137302_(_081287_, _081292_, _081295_);
  or g_137303_(_081285_, _081295_, _081296_);
  xor g_137304_(_081285_, _081294_, _081298_);
  not g_137305_(_081298_, _081299_);
  or g_137306_(_078468_, _081298_, _081300_);
  xor g_137307_(_078468_, _081299_, _081301_);
  not g_137308_(_081301_, _081302_);
  or g_137309_(_078472_, _081301_, _081303_);
  xor g_137310_(_078472_, _081302_, _081304_);
  not g_137311_(_081304_, _081305_);
  and g_137312_(_078475_, _078480_, _081306_);
  or g_137313_(_081304_, _081306_, _081307_);
  xor g_137314_(_081305_, _081306_, _081309_);
  not g_137315_(_081309_, _081310_);
  and g_137316_(_078484_, _078486_, _081311_);
  xor g_137317_(_081310_, _081311_, _081312_);
  not g_137318_(_081312_, _081313_);
  or g_137319_(_078489_, _081312_, _081314_);
  xor g_137320_(_078489_, _081313_, _081315_);
  and g_137321_(_078492_, _081315_, _081316_);
  or g_137322_(_078492_, _081312_, _081317_);
  not g_137323_(_081317_, _081318_);
  or g_137324_(_081316_, _081318_, _081320_);
  not g_137325_(_081320_, _081321_);
  and g_137326_(_078496_, _078498_, _081322_);
  xor g_137327_(_081321_, _081322_, _081323_);
  not g_137328_(_081323_, _081324_);
  or g_137329_(_078503_, _081323_, _081325_);
  not g_137330_(_081325_, _081326_);
  or g_137331_(_078508_, _081323_, _081327_);
  xor g_137332_(_078508_, _081324_, _081328_);
  and g_137333_(_078503_, _081328_, _081329_);
  or g_137334_(_081326_, _081329_, _081331_);
  not g_137335_(_081331_, _081332_);
  or g_137336_(_081274_, _081331_, _081333_);
  xor g_137337_(_081274_, _081332_, _081334_);
  not g_137338_(_081334_, _081335_);
  or g_137339_(_078521_, _081334_, _081336_);
  not g_137340_(_081336_, _081337_);
  or g_137341_(_078517_, _081334_, _081338_);
  xor g_137342_(_078517_, _081335_, _081339_);
  and g_137343_(_078521_, _081339_, _081340_);
  not g_137344_(_081340_, _081342_);
  and g_137345_(_081336_, _081342_, _081343_);
  or g_137346_(_081337_, _081340_, _081344_);
  xor g_137347_(_081273_, _081343_, _081345_);
  or g_137348_(_078532_, _081345_, _081346_);
  xor g_137349_(_078532_, _081345_, _081347_);
  not g_137350_(_081347_, _081348_);
  or g_137351_(_078535_, _081348_, _081349_);
  xor g_137352_(_078535_, _081347_, _081350_);
  not g_137353_(_081350_, _081351_);
  or g_137354_(_075544_, _078539_, _081353_);
  and g_137355_(_078538_, _081353_, _081354_);
  xor g_137356_(_081351_, _081354_, _081355_);
  or g_137357_(_075549_, _078539_, _081356_);
  not g_137358_(_081356_, _081357_);
  or g_137359_(_081355_, _081356_, _081358_);
  xor g_137360_(_081355_, _081356_, _081359_);
  xor g_137361_(_081355_, _081357_, _081360_);
  or g_137362_(_081272_, _081360_, _081361_);
  xor g_137363_(_081272_, _081359_, _081362_);
  not g_137364_(_081362_, _081364_);
  or g_137365_(_081271_, _081362_, _081365_);
  xor g_137366_(_081271_, _081364_, _081366_);
  not g_137367_(_081366_, _081367_);
  and g_137368_(_078543_, _078545_, _081368_);
  xor g_137369_(_081367_, _081368_, _081369_);
  or g_137370_(_078549_, _081369_, _081370_);
  xor g_137371_(_078549_, _081369_, _081371_);
  xor g_137372_(_078550_, _081369_, _081372_);
  and g_137373_(_078552_, _078555_, _081373_);
  xor g_137374_(_081371_, _081373_, _081375_);
  or g_137375_(_081270_, _081375_, _081376_);
  xor g_137376_(_081270_, _081375_, _081377_);
  or g_137377_(_075586_, _078556_, _081378_);
  not g_137378_(_081378_, _081379_);
  and g_137379_(_078562_, _081378_, _081380_);
  xor g_137380_(_081377_, _081380_, _081381_);
  xor g_137381_(_081268_, _081381_, _081382_);
  xor g_137382_(_081269_, _081381_, _081383_);
  or g_137383_(_078575_, _081383_, _081384_);
  or g_137384_(_078571_, _081383_, _081386_);
  xor g_137385_(_078571_, _081382_, _081387_);
  or g_137386_(_078577_, _081387_, _081388_);
  xor g_137387_(_078577_, _081387_, _081389_);
  or g_137388_(_078574_, _081389_, _081390_);
  and g_137389_(_081384_, _081390_, _081391_);
  not g_137390_(_081391_, _081392_);
  or g_137391_(_078582_, _081392_, _081393_);
  xor g_137392_(_078582_, _081391_, _081394_);
  not g_137393_(_081394_, _081395_);
  or g_137394_(_078585_, _081394_, _081397_);
  xor g_137395_(_078585_, _081395_, _081398_);
  and g_137396_(_078588_, _078591_, _081399_);
  and g_137397_(_081398_, _081399_, _081400_);
  not g_137398_(_081400_, _081401_);
  or g_137399_(_078591_, _081398_, _081402_);
  or g_137400_(_078588_, _081398_, _081403_);
  and g_137401_(_081402_, _081403_, _081404_);
  not g_137402_(_081404_, _081405_);
  and g_137403_(_081401_, _081404_, _081406_);
  or g_137404_(_081400_, _081405_, _081408_);
  or g_137405_(_081267_, _081408_, _081409_);
  xor g_137406_(_081267_, _081406_, _081410_);
  or g_137407_(_081265_, _081410_, _081411_);
  not g_137408_(_081411_, _081412_);
  xor g_137409_(_081265_, _081410_, _081413_);
  xor g_137410_(_081266_, _081410_, _081414_);
  or g_137411_(_078602_, _081413_, _081415_);
  not g_137412_(_081415_, _081416_);
  and g_137413_(_078600_, _081413_, _081417_);
  or g_137414_(_078601_, _081414_, _081419_);
  and g_137415_(_078598_, _081413_, _081420_);
  or g_137416_(_078599_, _081414_, _081421_);
  and g_137417_(_081419_, _081421_, _081422_);
  or g_137418_(_081417_, _081420_, _081423_);
  and g_137419_(_081415_, _081422_, _081424_);
  or g_137420_(_081416_, _081423_, _081425_);
  or g_137421_(_078608_, _081424_, _081426_);
  not g_137422_(_081426_, _081427_);
  and g_137423_(_078612_, _081427_, _081428_);
  or g_137424_(_078613_, _081426_, _081430_);
  or g_137425_(_078607_, _081425_, _081431_);
  or g_137426_(_078612_, _081425_, _081432_);
  not g_137427_(_081432_, _081433_);
  and g_137428_(_081431_, _081432_, _081434_);
  not g_137429_(_081434_, _081435_);
  and g_137430_(_081430_, _081434_, _081436_);
  or g_137431_(_081428_, _081435_, _081437_);
  or g_137432_(_078615_, _078618_, _081438_);
  xor g_137433_(_081436_, _081438_, _081439_);
  or g_137434_(_081263_, _081439_, _081441_);
  not g_137435_(_081441_, _081442_);
  xor g_137436_(_081263_, _081439_, _081443_);
  not g_137437_(_081443_, _081444_);
  or g_137438_(_075654_, _078620_, _081445_);
  or g_137439_(_081444_, _081445_, _081446_);
  not g_137440_(_081446_, _081447_);
  xor g_137441_(_081443_, _081445_, _081448_);
  or g_137442_(_081261_, _081448_, _081449_);
  xor g_137443_(_081262_, _081448_, _081450_);
  not g_137444_(_081450_, _081452_);
  or g_137445_(_078624_, _081450_, _081453_);
  xor g_137446_(_078624_, _081450_, _081454_);
  xor g_137447_(_078624_, _081452_, _081455_);
  or g_137448_(_078629_, _081455_, _081456_);
  not g_137449_(_081456_, _081457_);
  xor g_137450_(_078629_, _081454_, _081458_);
  or g_137451_(_078632_, _081458_, _081459_);
  xor g_137452_(_078633_, _081458_, _081460_);
  and g_137453_(_078638_, _078642_, _081461_);
  not g_137454_(_081461_, _081463_);
  xor g_137455_(_081460_, _081463_, _081464_);
  or g_137456_(_072751_, _081258_, _081465_);
  not g_137457_(_081465_, _081466_);
  or g_137458_(_081464_, _081465_, _081467_);
  xor g_137459_(_081464_, _081466_, _081468_);
  or g_137460_(_081259_, _081468_, _081469_);
  xor g_137461_(_081260_, _081468_, _081470_);
  or g_137462_(_081256_, _081470_, _081471_);
  xor g_137463_(_081257_, _081470_, _081472_);
  not g_137464_(_081472_, _081474_);
  or g_137465_(_078648_, _081472_, _081475_);
  xor g_137466_(_078648_, _081472_, _081476_);
  xor g_137467_(_078648_, _081474_, _081477_);
  or g_137468_(_081254_, _081477_, _081478_);
  not g_137469_(_081478_, _081479_);
  and g_137470_(_078651_, _081477_, _081480_);
  or g_137471_(_078652_, _081476_, _081481_);
  and g_137472_(_081254_, _081480_, _081482_);
  or g_137473_(_081255_, _081481_, _081483_);
  or g_137474_(_078651_, _081477_, _081485_);
  not g_137475_(_081485_, _081486_);
  and g_137476_(_081483_, _081485_, _081487_);
  or g_137477_(_081482_, _081486_, _081488_);
  and g_137478_(_081478_, _081487_, _081489_);
  or g_137479_(_081479_, _081488_, _081490_);
  or g_137480_(_081252_, _081490_, _081491_);
  xor g_137481_(_081252_, _081489_, _081492_);
  or g_137482_(_081250_, _081492_, _081493_);
  xor g_137483_(_081251_, _081492_, _081494_);
  or g_137484_(_081249_, _081494_, _081496_);
  xor g_137485_(_081249_, _081494_, _081497_);
  not g_137486_(_081497_, _081498_);
  and g_137487_(_078661_, _081497_, _081499_);
  or g_137488_(_078660_, _081498_, _081500_);
  xor g_137489_(_078660_, _081497_, _081501_);
  not g_137490_(_081501_, _081502_);
  and g_137491_(_078664_, _081502_, _081503_);
  or g_137492_(_078665_, _081501_, _081504_);
  xor g_137493_(_078664_, _081501_, _081505_);
  or g_137494_(_078666_, _081505_, _081507_);
  xor g_137495_(_078667_, _081505_, _081508_);
  or g_137496_(_075706_, _078671_, _081509_);
  or g_137497_(_081508_, _081509_, _081510_);
  xor g_137498_(_081508_, _081509_, _081511_);
  not g_137499_(_081511_, _081512_);
  or g_137500_(_081248_, _081512_, _081513_);
  xor g_137501_(_081248_, _081511_, _081514_);
  not g_137502_(_081514_, _081515_);
  or g_137503_(_081247_, _081514_, _081516_);
  xor g_137504_(_081247_, _081514_, _081518_);
  xor g_137505_(_081247_, _081515_, _081519_);
  or g_137506_(_081246_, _081519_, _081520_);
  xor g_137507_(_081246_, _081518_, _081521_);
  or g_137508_(_072800_, _081245_, _081522_);
  not g_137509_(_081522_, _081523_);
  or g_137510_(_081521_, _081522_, _081524_);
  xor g_137511_(_081521_, _081523_, _081525_);
  or g_137512_(_078678_, _078682_, _081526_);
  xor g_137513_(_081525_, _081526_, _081527_);
  not g_137514_(_081527_, _081529_);
  or g_137515_(_078685_, _081527_, _081530_);
  xor g_137516_(_078685_, _081527_, _081531_);
  xor g_137517_(_078685_, _081529_, _081532_);
  or g_137518_(_078687_, _081532_, _081533_);
  xor g_137519_(_078687_, _081531_, _081534_);
  or g_137520_(_075749_, _078684_, _081535_);
  not g_137521_(_081535_, _081536_);
  or g_137522_(_081534_, _081535_, _081537_);
  xor g_137523_(_081534_, _081536_, _081538_);
  or g_137524_(_081244_, _081538_, _081540_);
  xor g_137525_(_081244_, _081538_, _081541_);
  not g_137526_(_081541_, _081542_);
  or g_137527_(_078388_, _078688_, _081543_);
  not g_137528_(_081543_, _081544_);
  and g_137529_(_081541_, _081544_, _081545_);
  or g_137530_(_081542_, _081543_, _081546_);
  xor g_137531_(_081541_, _081543_, _081547_);
  or g_137532_(_081243_, _081547_, _081548_);
  not g_137533_(_081548_, _081549_);
  xor g_137534_(_081241_, _081547_, _081551_);
  or g_137535_(_078696_, _081551_, _081552_);
  xor g_137536_(_078696_, _081551_, _081553_);
  xor g_137537_(_078697_, _081551_, _081554_);
  and g_137538_(_078701_, _081554_, _081555_);
  or g_137539_(_078703_, _081553_, _081556_);
  and g_137540_(_081239_, _081555_, _081557_);
  or g_137541_(_081240_, _081556_, _081558_);
  or g_137542_(_081239_, _081554_, _081559_);
  or g_137543_(_078701_, _081554_, _081560_);
  and g_137544_(_081559_, _081560_, _081562_);
  not g_137545_(_081562_, _081563_);
  and g_137546_(_081558_, _081562_, _081564_);
  or g_137547_(_081557_, _081563_, _081565_);
  or g_137548_(_075765_, _078704_, _081566_);
  or g_137549_(_075772_, _078704_, _081567_);
  and g_137550_(_081566_, _081567_, _081568_);
  xor g_137551_(_081564_, _081568_, _081569_);
  or g_137552_(_081238_, _081569_, _081570_);
  xor g_137553_(_081238_, _081569_, _081571_);
  not g_137554_(_081571_, _081573_);
  or g_137555_(_078711_, _081573_, _081574_);
  xor g_137556_(_078711_, _081571_, _081575_);
  or g_137557_(_078715_, _081575_, _081576_);
  xor g_137558_(_078716_, _081575_, _081577_);
  not g_137559_(_081577_, _081578_);
  or g_137560_(_081237_, _081577_, _081579_);
  xor g_137561_(_081237_, _081577_, _081580_);
  xor g_137562_(_081237_, _081578_, _081581_);
  or g_137563_(_081236_, _081581_, _081582_);
  xor g_137564_(_081236_, _081580_, _081584_);
  or g_137565_(_078722_, _081584_, _081585_);
  not g_137566_(_081585_, _081586_);
  and g_137567_(_075786_, _078718_, _081587_);
  or g_137568_(_075785_, _078719_, _081588_);
  or g_137569_(_081584_, _081588_, _081589_);
  xor g_137570_(_081584_, _081587_, _081590_);
  and g_137571_(_078722_, _081590_, _081591_);
  or g_137572_(_081586_, _081591_, _081592_);
  or g_137573_(_078727_, _081592_, _081593_);
  xor g_137574_(_078726_, _081592_, _081595_);
  and g_137575_(_078730_, _078733_, _081596_);
  not g_137576_(_081596_, _081597_);
  xor g_137577_(_081595_, _081597_, _081598_);
  or g_137578_(_078738_, _081598_, _081599_);
  xor g_137579_(_078739_, _081598_, _081600_);
  or g_137580_(_078748_, _081600_, _081601_);
  not g_137581_(_081601_, _081602_);
  and g_137582_(_078743_, _081600_, _081603_);
  and g_137583_(_078748_, _081603_, _081604_);
  or g_137584_(_078743_, _081598_, _081606_);
  not g_137585_(_081606_, _081607_);
  or g_137586_(_081604_, _081607_, _081608_);
  or g_137587_(_081602_, _081608_, _081609_);
  not g_137588_(_081609_, _081610_);
  or g_137589_(_078750_, _081609_, _081611_);
  xor g_137590_(_078750_, _081609_, _081612_);
  xor g_137591_(_078750_, _081610_, _081613_);
  and g_137592_(_078752_, _081613_, _081614_);
  or g_137593_(_075820_, _078751_, _081615_);
  not g_137594_(_081615_, _081617_);
  and g_137595_(_081612_, _081617_, _081618_);
  or g_137596_(_081613_, _081615_, _081619_);
  and g_137597_(_067915_, _081618_, _081620_);
  or g_137598_(_067914_, _081619_, _081621_);
  or g_137599_(_081614_, _081620_, _081622_);
  or g_137600_(_072891_, _081233_, _081623_);
  or g_137601_(_067876_, _081623_, _081624_);
  and g_137602_(_081622_, _081624_, _081625_);
  not g_137603_(_081625_, _081626_);
  or g_137604_(_081622_, _081623_, _081628_);
  not g_137605_(_081628_, _081629_);
  or g_137606_(_067876_, _081628_, _081630_);
  and g_137607_(_081626_, _081630_, _081631_);
  not g_137608_(_081631_, _081632_);
  or g_137609_(_081234_, _081632_, _081633_);
  xor g_137610_(_081234_, _081631_, _081634_);
  or g_137611_(_081230_, _081634_, _081635_);
  xor g_137612_(_081232_, _081634_, _081636_);
  and g_137613_(_078758_, _078760_, _081637_);
  not g_137614_(_081637_, _081639_);
  xor g_137615_(_081636_, _081639_, _081640_);
  or g_137616_(_078766_, _081640_, _081641_);
  not g_137617_(_081641_, _081642_);
  or g_137618_(_078762_, _081640_, _081643_);
  xor g_137619_(_078763_, _081640_, _081644_);
  and g_137620_(_078766_, _081644_, _081645_);
  or g_137621_(_081642_, _081645_, _081646_);
  or g_137622_(_078770_, _081646_, _081647_);
  not g_137623_(_081647_, _081648_);
  xor g_137624_(_078771_, _081646_, _081650_);
  or g_137625_(_072923_, _081227_, _081651_);
  and g_137626_(_078774_, _081651_, _081652_);
  not g_137627_(_081652_, _081653_);
  xor g_137628_(_081650_, _081653_, _081654_);
  not g_137629_(_081654_, _081655_);
  and g_137630_(_081229_, _081655_, _081656_);
  not g_137631_(_081656_, _081657_);
  xor g_137632_(_081228_, _081654_, _081658_);
  not g_137633_(_081658_, _081659_);
  or g_137634_(_081226_, _081659_, _081661_);
  xor g_137635_(_081226_, _081658_, _081662_);
  and g_137636_(_078780_, _078783_, _081663_);
  or g_137637_(_081662_, _081663_, _081664_);
  xor g_137638_(_081662_, _081663_, _081665_);
  not g_137639_(_081665_, _081666_);
  or g_137640_(_078786_, _081666_, _081667_);
  xor g_137641_(_078786_, _081665_, _081668_);
  or g_137642_(_078789_, _081668_, _081669_);
  not g_137643_(_081669_, _081670_);
  or g_137644_(_078792_, _081668_, _081672_);
  xor g_137645_(_078793_, _081668_, _081673_);
  and g_137646_(_078789_, _081673_, _081674_);
  or g_137647_(_081670_, _081674_, _081675_);
  or g_137648_(_078806_, _081675_, _081676_);
  not g_137649_(_081676_, _081677_);
  or g_137650_(_078803_, _081675_, _081678_);
  xor g_137651_(_078802_, _081675_, _081679_);
  or g_137652_(_078800_, _081679_, _081680_);
  not g_137653_(_081680_, _081681_);
  xor g_137654_(_078799_, _081679_, _081683_);
  and g_137655_(_078806_, _081683_, _081684_);
  or g_137656_(_081677_, _081684_, _081685_);
  or g_137657_(_078808_, _081685_, _081686_);
  xor g_137658_(_078808_, _081685_, _081687_);
  xor g_137659_(_078809_, _081685_, _081688_);
  and g_137660_(_078811_, _081688_, _081689_);
  or g_137661_(_075891_, _078805_, _081690_);
  not g_137662_(_081690_, _081691_);
  and g_137663_(_081687_, _081691_, _081692_);
  or g_137664_(_081688_, _081690_, _081694_);
  or g_137665_(_081689_, _081692_, _081695_);
  or g_137666_(_078814_, _081695_, _081696_);
  xor g_137667_(_078815_, _081695_, _081697_);
  or g_137668_(_075894_, _078810_, _081698_);
  not g_137669_(_081698_, _081699_);
  or g_137670_(_081697_, _081698_, _081700_);
  xor g_137671_(_081697_, _081699_, _081701_);
  or g_137672_(_075903_, _078820_, _081702_);
  not g_137673_(_081702_, _081703_);
  or g_137674_(_081701_, _081702_, _081705_);
  xor g_137675_(_081701_, _081703_, _081706_);
  or g_137676_(_081224_, _081706_, _081707_);
  xor g_137677_(_081225_, _081706_, _081708_);
  or g_137678_(_078822_, _081708_, _081709_);
  xor g_137679_(_078824_, _081708_, _081710_);
  not g_137680_(_081710_, _081711_);
  and g_137681_(_078826_, _078830_, _081712_);
  xor g_137682_(_081710_, _081712_, _081713_);
  xor g_137683_(_081711_, _081712_, _081714_);
  or g_137684_(_078833_, _081714_, _081716_);
  xor g_137685_(_078833_, _081713_, _081717_);
  or g_137686_(_081222_, _081717_, _081718_);
  not g_137687_(_081718_, _081719_);
  xor g_137688_(_081223_, _081717_, _081720_);
  not g_137689_(_081720_, _081721_);
  or g_137690_(_081218_, _081720_, _081722_);
  not g_137691_(_081722_, _081723_);
  xor g_137692_(_081218_, _081720_, _081724_);
  xor g_137693_(_081219_, _081720_, _081725_);
  and g_137694_(_078841_, _081724_, _081727_);
  or g_137695_(_078840_, _081725_, _081728_);
  or g_137696_(_075930_, _078835_, _081729_);
  not g_137697_(_081729_, _081730_);
  and g_137698_(_081721_, _081730_, _081731_);
  not g_137699_(_081731_, _081732_);
  or g_137700_(_081727_, _081731_, _081733_);
  not g_137701_(_081733_, _081734_);
  and g_137702_(_081725_, _081729_, _081735_);
  and g_137703_(_078840_, _081735_, _081736_);
  or g_137704_(_081733_, _081736_, _081738_);
  or g_137705_(_078846_, _081738_, _081739_);
  xor g_137706_(_078847_, _081738_, _081740_);
  and g_137707_(_078850_, _078853_, _081741_);
  not g_137708_(_081741_, _081742_);
  xor g_137709_(_081740_, _081742_, _081743_);
  or g_137710_(_078855_, _081743_, _081744_);
  xor g_137711_(_078857_, _081743_, _081745_);
  not g_137712_(_081745_, _081746_);
  or g_137713_(_081216_, _081745_, _081747_);
  xor g_137714_(_081216_, _081745_, _081749_);
  xor g_137715_(_081216_, _081746_, _081750_);
  or g_137716_(_081215_, _081750_, _081751_);
  xor g_137717_(_081215_, _081749_, _081752_);
  or g_137718_(_078863_, _081752_, _081753_);
  xor g_137719_(_078863_, _081752_, _081754_);
  xor g_137720_(_078864_, _081752_, _081755_);
  or g_137721_(_078868_, _081755_, _081756_);
  xor g_137722_(_078868_, _081754_, _081757_);
  or g_137723_(_081213_, _081757_, _081758_);
  xor g_137724_(_081214_, _081757_, _081760_);
  and g_137725_(_073036_, _075961_, _081761_);
  not g_137726_(_081761_, _081762_);
  or g_137727_(_078869_, _081762_, _081763_);
  or g_137728_(_078869_, _078871_, _081764_);
  and g_137729_(_081763_, _081764_, _081765_);
  not g_137730_(_081765_, _081766_);
  xor g_137731_(_081760_, _081766_, _081767_);
  or g_137732_(_078875_, _081767_, _081768_);
  xor g_137733_(_078875_, _081767_, _081769_);
  xor g_137734_(_078876_, _081767_, _081771_);
  and g_137735_(_078881_, _078884_, _081772_);
  xor g_137736_(_081769_, _081772_, _081773_);
  or g_137737_(_078888_, _081773_, _081774_);
  xor g_137738_(_078890_, _081773_, _081775_);
  or g_137739_(_078892_, _081775_, _081776_);
  xor g_137740_(_078893_, _081775_, _081777_);
  or g_137741_(_078896_, _081777_, _081778_);
  xor g_137742_(_078897_, _081777_, _081779_);
  and g_137743_(_078899_, _078902_, _081780_);
  not g_137744_(_081780_, _081782_);
  xor g_137745_(_081779_, _081782_, _081783_);
  not g_137746_(_081783_, _081784_);
  and g_137747_(_081210_, _081784_, _081785_);
  not g_137748_(_081785_, _081786_);
  xor g_137749_(_081208_, _081783_, _081787_);
  not g_137750_(_081787_, _081788_);
  and g_137751_(_081207_, _081787_, _081789_);
  or g_137752_(_081206_, _081788_, _081790_);
  xor g_137753_(_081206_, _081787_, _081791_);
  or g_137754_(_078905_, _081791_, _081793_);
  xor g_137755_(_078905_, _081791_, _081794_);
  not g_137756_(_081794_, _081795_);
  and g_137757_(_078909_, _081794_, _081796_);
  not g_137758_(_081796_, _081797_);
  or g_137759_(_078914_, _081795_, _081798_);
  xor g_137760_(_078914_, _081794_, _081799_);
  and g_137761_(_078908_, _081799_, _081800_);
  or g_137762_(_081796_, _081800_, _081801_);
  or g_137763_(_078917_, _081801_, _081802_);
  xor g_137764_(_078918_, _081801_, _081804_);
  and g_137765_(_078921_, _081804_, _081805_);
  or g_137766_(_078921_, _081804_, _081806_);
  xor g_137767_(_078923_, _081804_, _081807_);
  not g_137768_(_081807_, _081808_);
  or g_137769_(_078927_, _081807_, _081809_);
  xor g_137770_(_078927_, _081808_, _081810_);
  and g_137771_(_078930_, _081810_, _081811_);
  or g_137772_(_078930_, _081807_, _081812_);
  not g_137773_(_081812_, _081813_);
  or g_137774_(_081811_, _081813_, _081815_);
  or g_137775_(_081205_, _081815_, _081816_);
  xor g_137776_(_081204_, _081815_, _081817_);
  or g_137777_(_081202_, _081817_, _081818_);
  xor g_137778_(_081203_, _081817_, _081819_);
  or g_137779_(_078938_, _081819_, _081820_);
  xor g_137780_(_078937_, _081819_, _081821_);
  and g_137781_(_078940_, _078942_, _081822_);
  not g_137782_(_081822_, _081823_);
  xor g_137783_(_081821_, _081823_, _081824_);
  xor g_137784_(_081821_, _081822_, _081826_);
  and g_137785_(_078946_, _081826_, _081827_);
  or g_137786_(_078945_, _081824_, _081828_);
  xor g_137787_(_078945_, _081824_, _081829_);
  xor g_137788_(_078946_, _081824_, _081830_);
  or g_137789_(_078949_, _081829_, _081831_);
  or g_137790_(_076040_, _078941_, _081832_);
  or g_137791_(_081830_, _081832_, _081833_);
  and g_137792_(_081831_, _081833_, _081834_);
  and g_137793_(_078952_, _081834_, _081835_);
  xor g_137794_(_078951_, _081834_, _081837_);
  and g_137795_(_078954_, _081837_, _081838_);
  and g_137796_(_078956_, _081834_, _081839_);
  or g_137797_(_081838_, _081839_, _081840_);
  and g_137798_(_078958_, _078961_, _081841_);
  not g_137799_(_081841_, _081842_);
  xor g_137800_(_081840_, _081841_, _081843_);
  xor g_137801_(_081840_, _081842_, _081844_);
  and g_137802_(_081201_, _081843_, _081845_);
  or g_137803_(_081200_, _081844_, _081846_);
  and g_137804_(_078964_, _081843_, _081848_);
  or g_137805_(_078963_, _081844_, _081849_);
  and g_137806_(_081846_, _081849_, _081850_);
  or g_137807_(_081845_, _081848_, _081851_);
  and g_137808_(_078963_, _081844_, _081852_);
  and g_137809_(_081200_, _081852_, _081853_);
  or g_137810_(_081851_, _081853_, _081854_);
  not g_137811_(_081854_, _081855_);
  or g_137812_(_081199_, _081854_, _081856_);
  xor g_137813_(_081199_, _081854_, _081857_);
  xor g_137814_(_081199_, _081855_, _081859_);
  or g_137815_(_078969_, _081859_, _081860_);
  xor g_137816_(_078969_, _081857_, _081861_);
  and g_137817_(_078972_, _081861_, _081862_);
  or g_137818_(_078972_, _081861_, _081863_);
  not g_137819_(_081863_, _081864_);
  xor g_137820_(_078972_, _081861_, _081865_);
  or g_137821_(_081862_, _081864_, _081866_);
  and g_137822_(_078976_, _078979_, _081867_);
  xor g_137823_(_081865_, _081867_, _081868_);
  or g_137824_(_078982_, _081868_, _081870_);
  xor g_137825_(_078982_, _081868_, _081871_);
  not g_137826_(_081871_, _081872_);
  and g_137827_(_078986_, _081871_, _081873_);
  or g_137828_(_078985_, _081872_, _081874_);
  or g_137829_(_078989_, _081872_, _081875_);
  xor g_137830_(_078989_, _081871_, _081876_);
  and g_137831_(_078985_, _081876_, _081877_);
  or g_137832_(_081873_, _081877_, _081878_);
  or g_137833_(_078992_, _081878_, _081879_);
  xor g_137834_(_078993_, _081878_, _081881_);
  not g_137835_(_081881_, _081882_);
  or g_137836_(_078996_, _081881_, _081883_);
  xor g_137837_(_078996_, _081881_, _081884_);
  xor g_137838_(_078996_, _081882_, _081885_);
  and g_137839_(_078998_, _079003_, _081886_);
  and g_137840_(_081885_, _081886_, _081887_);
  and g_137841_(_079000_, _081884_, _081888_);
  or g_137842_(_078998_, _081885_, _081889_);
  and g_137843_(_079004_, _081884_, _081890_);
  or g_137844_(_079003_, _081885_, _081892_);
  or g_137845_(_081888_, _081890_, _081893_);
  or g_137846_(_081887_, _081893_, _081894_);
  not g_137847_(_081894_, _081895_);
  or g_137848_(_076103_, _079008_, _081896_);
  and g_137849_(_079007_, _081896_, _081897_);
  xor g_137850_(_081895_, _081897_, _081898_);
  xor g_137851_(_081894_, _081897_, _081899_);
  or g_137852_(_079009_, _081898_, _081900_);
  not g_137853_(_081900_, _081901_);
  xor g_137854_(_079009_, _081899_, _081903_);
  and g_137855_(_079013_, _079016_, _081904_);
  xor g_137856_(_081903_, _081904_, _081905_);
  not g_137857_(_081905_, _081906_);
  or g_137858_(_079018_, _081906_, _081907_);
  xor g_137859_(_079019_, _081905_, _081908_);
  xor g_137860_(_079018_, _081905_, _081909_);
  or g_137861_(_079025_, _081908_, _081910_);
  or g_137862_(_079029_, _081910_, _081911_);
  or g_137863_(_079030_, _081909_, _081912_);
  not g_137864_(_081912_, _081914_);
  and g_137865_(_079025_, _081908_, _081915_);
  or g_137866_(_079026_, _081909_, _081916_);
  and g_137867_(_081912_, _081916_, _081917_);
  and g_137868_(_081911_, _081917_, _081918_);
  not g_137869_(_081918_, _081919_);
  or g_137870_(_081197_, _081919_, _081920_);
  xor g_137871_(_081197_, _081918_, _081921_);
  or g_137872_(_076122_, _079027_, _081922_);
  not g_137873_(_081922_, _081923_);
  or g_137874_(_081921_, _081922_, _081925_);
  xor g_137875_(_081921_, _081923_, _081926_);
  and g_137876_(_079036_, _079038_, _081927_);
  not g_137877_(_081927_, _081928_);
  xor g_137878_(_081926_, _081928_, _081929_);
  xor g_137879_(_081926_, _081927_, _081930_);
  xor g_137880_(_081196_, _081929_, _081931_);
  xor g_137881_(_081196_, _081930_, _081932_);
  or g_137882_(_081195_, _081931_, _081933_);
  or g_137883_(_076157_, _079039_, _081934_);
  or g_137884_(_081932_, _081934_, _081936_);
  not g_137885_(_081936_, _081937_);
  and g_137886_(_081933_, _081936_, _081938_);
  not g_137887_(_081938_, _081939_);
  or g_137888_(_081193_, _081939_, _081940_);
  xor g_137889_(_081193_, _081938_, _081941_);
  or g_137890_(_081191_, _081941_, _081942_);
  xor g_137891_(_081192_, _081941_, _081943_);
  or g_137892_(_073234_, _081188_, _081944_);
  or g_137893_(_081943_, _081944_, _081945_);
  xor g_137894_(_081943_, _081944_, _081947_);
  not g_137895_(_081947_, _081948_);
  and g_137896_(_081190_, _081947_, _081949_);
  or g_137897_(_081189_, _081948_, _081950_);
  xor g_137898_(_081189_, _081947_, _081951_);
  or g_137899_(_081186_, _081951_, _081952_);
  xor g_137900_(_081185_, _081951_, _081953_);
  and g_137901_(_079050_, _079053_, _081954_);
  or g_137902_(_081953_, _081954_, _081955_);
  xor g_137903_(_081953_, _081954_, _081956_);
  not g_137904_(_081956_, _081958_);
  or g_137905_(_079057_, _081958_, _081959_);
  xor g_137906_(_079057_, _081956_, _081960_);
  or g_137907_(_081183_, _081960_, _081961_);
  xor g_137908_(_081184_, _081960_, _081962_);
  or g_137909_(_073257_, _076185_, _081963_);
  or g_137910_(_079058_, _081963_, _081964_);
  not g_137911_(_081964_, _081965_);
  or g_137912_(_081962_, _081964_, _081966_);
  xor g_137913_(_081962_, _081964_, _081967_);
  xor g_137914_(_081962_, _081965_, _081969_);
  or g_137915_(_076190_, _079058_, _081970_);
  not g_137916_(_081970_, _081971_);
  and g_137917_(_081969_, _081970_, _081972_);
  or g_137918_(_081967_, _081971_, _081973_);
  and g_137919_(_081180_, _081972_, _081974_);
  or g_137920_(_081181_, _081973_, _081975_);
  or g_137921_(_081180_, _081969_, _081976_);
  or g_137922_(_081969_, _081970_, _081977_);
  and g_137923_(_081976_, _081977_, _081978_);
  not g_137924_(_081978_, _081980_);
  and g_137925_(_081975_, _081978_, _081981_);
  or g_137926_(_081974_, _081980_, _081982_);
  or g_137927_(_081179_, _081982_, _081983_);
  xor g_137928_(_081179_, _081981_, _081984_);
  or g_137929_(_081177_, _081984_, _081985_);
  xor g_137930_(_081177_, _081984_, _081986_);
  xor g_137931_(_081178_, _081984_, _081987_);
  and g_137932_(_079067_, _081987_, _081988_);
  or g_137933_(_079066_, _081986_, _081989_);
  and g_137934_(_076200_, _079062_, _081991_);
  or g_137935_(_076201_, _079061_, _081992_);
  and g_137936_(_081986_, _081991_, _081993_);
  or g_137937_(_081987_, _081992_, _081994_);
  and g_137938_(_081989_, _081994_, _081995_);
  or g_137939_(_081988_, _081993_, _081996_);
  or g_137940_(_079070_, _081995_, _081997_);
  or g_137941_(_079074_, _081997_, _081998_);
  or g_137942_(_079075_, _081996_, _081999_);
  not g_137943_(_081999_, _082000_);
  or g_137944_(_079071_, _081996_, _082002_);
  and g_137945_(_081999_, _082002_, _082003_);
  and g_137946_(_081998_, _082003_, _082004_);
  not g_137947_(_082004_, _082005_);
  or g_137948_(_079082_, _082005_, _082006_);
  xor g_137949_(_079082_, _082004_, _082007_);
  or g_137950_(_079080_, _082007_, _082008_);
  xor g_137951_(_079081_, _082007_, _082009_);
  and g_137952_(_079088_, _079090_, _082010_);
  and g_137953_(_082009_, _082010_, _082011_);
  not g_137954_(_082011_, _082013_);
  or g_137955_(_079088_, _082009_, _082014_);
  or g_137956_(_079090_, _082009_, _082015_);
  and g_137957_(_082014_, _082015_, _082016_);
  and g_137958_(_082013_, _082016_, _082017_);
  not g_137959_(_082017_, _082018_);
  or g_137960_(_079094_, _082018_, _082019_);
  xor g_137961_(_079095_, _082017_, _082020_);
  xor g_137962_(_079094_, _082017_, _082021_);
  or g_137963_(_076241_, _079100_, _082022_);
  not g_137964_(_082022_, _082024_);
  or g_137965_(_082021_, _082022_, _082025_);
  or g_137966_(_079097_, _082021_, _082026_);
  and g_137967_(_082025_, _082026_, _082027_);
  not g_137968_(_082027_, _082028_);
  and g_137969_(_079097_, _082021_, _082029_);
  or g_137970_(_079099_, _082020_, _082030_);
  and g_137971_(_082022_, _082029_, _082031_);
  or g_137972_(_082024_, _082030_, _082032_);
  and g_137973_(_082027_, _082032_, _082033_);
  or g_137974_(_082028_, _082031_, _082035_);
  or g_137975_(_081175_, _082035_, _082036_);
  xor g_137976_(_081175_, _082033_, _082037_);
  or g_137977_(_079105_, _082037_, _082038_);
  xor g_137978_(_079106_, _082037_, _082039_);
  not g_137979_(_082039_, _082040_);
  or g_137980_(_079104_, _082039_, _082041_);
  xor g_137981_(_079104_, _082039_, _082042_);
  xor g_137982_(_079104_, _082040_, _082043_);
  or g_137983_(_079112_, _082043_, _082044_);
  xor g_137984_(_079112_, _082042_, _082046_);
  or g_137985_(_079115_, _082046_, _082047_);
  xor g_137986_(_079115_, _082046_, _082048_);
  not g_137987_(_082048_, _082049_);
  or g_137988_(_081174_, _082049_, _082050_);
  xor g_137989_(_081174_, _082048_, _082051_);
  or g_137990_(_081173_, _082051_, _082052_);
  xor g_137991_(_081172_, _082051_, _082053_);
  or g_137992_(_076263_, _079119_, _082054_);
  not g_137993_(_082054_, _082055_);
  or g_137994_(_082053_, _082054_, _082057_);
  xor g_137995_(_082053_, _082055_, _082058_);
  or g_137996_(_081170_, _082058_, _082059_);
  xor g_137997_(_081170_, _082058_, _082060_);
  xor g_137998_(_081171_, _082058_, _082061_);
  or g_137999_(_079123_, _082061_, _082062_);
  xor g_138000_(_079123_, _082061_, _082063_);
  xor g_138001_(_079123_, _082060_, _082064_);
  or g_138002_(_079125_, _082064_, _082065_);
  not g_138003_(_082065_, _082066_);
  xor g_138004_(_079125_, _082063_, _082068_);
  or g_138005_(_079127_, _082068_, _082069_);
  xor g_138006_(_079128_, _082068_, _082070_);
  or g_138007_(_079133_, _082070_, _082071_);
  not g_138008_(_082071_, _082072_);
  xor g_138009_(_079134_, _082070_, _082073_);
  or g_138010_(_079137_, _082073_, _082074_);
  xor g_138011_(_079138_, _082073_, _082075_);
  not g_138012_(_082075_, _082076_);
  and g_138013_(_079140_, _079145_, _082077_);
  xor g_138014_(_082075_, _082077_, _082079_);
  xor g_138015_(_082076_, _082077_, _082080_);
  or g_138016_(_079148_, _082080_, _082081_);
  xor g_138017_(_079148_, _082079_, _082082_);
  and g_138018_(_079150_, _079154_, _082083_);
  or g_138019_(_082082_, _082083_, _082084_);
  not g_138020_(_082084_, _082085_);
  xor g_138021_(_082082_, _082083_, _082086_);
  not g_138022_(_082086_, _082087_);
  and g_138023_(_079160_, _082086_, _082088_);
  or g_138024_(_079159_, _082087_, _082090_);
  xor g_138025_(_079159_, _082086_, _082091_);
  not g_138026_(_082091_, _082092_);
  or g_138027_(_079161_, _082091_, _082093_);
  not g_138028_(_082093_, _082094_);
  xor g_138029_(_079161_, _082091_, _082095_);
  xor g_138030_(_079161_, _082092_, _082096_);
  or g_138031_(_079166_, _082096_, _082097_);
  not g_138032_(_082097_, _082098_);
  xor g_138033_(_079166_, _082096_, _082099_);
  xor g_138034_(_079166_, _082095_, _082101_);
  or g_138035_(_079169_, _082101_, _082102_);
  not g_138036_(_082102_, _082103_);
  xor g_138037_(_079169_, _082099_, _082104_);
  or g_138038_(_079172_, _082104_, _082105_);
  xor g_138039_(_079173_, _082104_, _082106_);
  and g_138040_(_079176_, _079179_, _082107_);
  not g_138041_(_082107_, _082108_);
  xor g_138042_(_082106_, _082108_, _082109_);
  not g_138043_(_082109_, _082110_);
  xor g_138044_(_081169_, _082110_, _082112_);
  or g_138045_(_079191_, _082112_, _082113_);
  xor g_138046_(_079191_, _082112_, _082114_);
  not g_138047_(_082114_, _082115_);
  or g_138048_(_079193_, _082115_, _082116_);
  xor g_138049_(_079193_, _082114_, _082117_);
  not g_138050_(_082117_, _082118_);
  and g_138051_(_079196_, _079199_, _082119_);
  or g_138052_(_082117_, _082119_, _082120_);
  xor g_138053_(_082117_, _082119_, _082121_);
  xor g_138054_(_082118_, _082119_, _082123_);
  xor g_138055_(_081168_, _082121_, _082124_);
  or g_138056_(_079209_, _082124_, _082125_);
  not g_138057_(_082125_, _082126_);
  and g_138058_(_079209_, _082124_, _082127_);
  xor g_138059_(_079209_, _082124_, _082128_);
  or g_138060_(_082126_, _082127_, _082129_);
  or g_138061_(_079212_, _082129_, _082130_);
  xor g_138062_(_079212_, _082128_, _082131_);
  not g_138063_(_082131_, _082132_);
  or g_138064_(_079214_, _082131_, _082134_);
  xor g_138065_(_079214_, _082131_, _082135_);
  xor g_138066_(_079214_, _082132_, _082136_);
  or g_138067_(_081167_, _082136_, _082137_);
  not g_138068_(_082137_, _082138_);
  xor g_138069_(_081167_, _082135_, _082139_);
  or g_138070_(_081164_, _082139_, _082140_);
  xor g_138071_(_081164_, _082139_, _082141_);
  xor g_138072_(_081166_, _082139_, _082142_);
  or g_138073_(_079220_, _082142_, _082143_);
  not g_138074_(_082143_, _082145_);
  xor g_138075_(_079220_, _082141_, _082146_);
  not g_138076_(_082146_, _082147_);
  or g_138077_(_079223_, _082146_, _082148_);
  xor g_138078_(_079223_, _082146_, _082149_);
  xor g_138079_(_079223_, _082147_, _082150_);
  or g_138080_(_079225_, _082150_, _082151_);
  xor g_138081_(_079225_, _082149_, _082152_);
  or g_138082_(_079227_, _082152_, _082153_);
  not g_138083_(_082153_, _082154_);
  xor g_138084_(_079228_, _082152_, _082156_);
  or g_138085_(_079232_, _082156_, _082157_);
  xor g_138086_(_079232_, _082156_, _082158_);
  xor g_138087_(_079233_, _082156_, _082159_);
  and g_138088_(_079236_, _079240_, _082160_);
  xor g_138089_(_082158_, _082160_, _082161_);
  or g_138090_(_079243_, _082161_, _082162_);
  not g_138091_(_082162_, _082163_);
  xor g_138092_(_079243_, _082161_, _082164_);
  xor g_138093_(_081163_, _082164_, _082165_);
  or g_138094_(_081162_, _082165_, _082167_);
  not g_138095_(_082167_, _082168_);
  xor g_138096_(_081162_, _082165_, _082169_);
  not g_138097_(_082169_, _082170_);
  and g_138098_(_079248_, _082169_, _082171_);
  or g_138099_(_079249_, _082170_, _082172_);
  xor g_138100_(_079248_, _082169_, _082173_);
  xor g_138101_(_079249_, _082169_, _082174_);
  or g_138102_(_079255_, _082174_, _082175_);
  or g_138103_(_079251_, _082174_, _082176_);
  and g_138104_(_082175_, _082176_, _082178_);
  not g_138105_(_082178_, _082179_);
  and g_138106_(_079251_, _082174_, _082180_);
  or g_138107_(_079253_, _082173_, _082181_);
  and g_138108_(_079255_, _082180_, _082182_);
  or g_138109_(_079256_, _082181_, _082183_);
  and g_138110_(_082178_, _082183_, _082184_);
  or g_138111_(_082179_, _082182_, _082185_);
  or g_138112_(_081161_, _082185_, _082186_);
  xor g_138113_(_081161_, _082184_, _082187_);
  or g_138114_(_081159_, _082187_, _082189_);
  not g_138115_(_082189_, _082190_);
  xor g_138116_(_081160_, _082187_, _082191_);
  not g_138117_(_082191_, _082192_);
  or g_138118_(_079260_, _082191_, _082193_);
  xor g_138119_(_079260_, _082191_, _082194_);
  xor g_138120_(_079260_, _082192_, _082195_);
  or g_138121_(_076397_, _079265_, _082196_);
  and g_138122_(_079264_, _082196_, _082197_);
  xor g_138123_(_082194_, _082197_, _082198_);
  or g_138124_(_081157_, _082198_, _082200_);
  not g_138125_(_082200_, _082201_);
  xor g_138126_(_081157_, _082198_, _082202_);
  not g_138127_(_082202_, _082203_);
  or g_138128_(_081155_, _082203_, _082204_);
  not g_138129_(_082204_, _082205_);
  xor g_138130_(_081156_, _082202_, _082206_);
  xor g_138131_(_081155_, _082202_, _082207_);
  or g_138132_(_076402_, _079267_, _082208_);
  or g_138133_(_082207_, _082208_, _082209_);
  xor g_138134_(_082206_, _082208_, _082211_);
  or g_138135_(_081152_, _082211_, _082212_);
  xor g_138136_(_081153_, _082211_, _082213_);
  and g_138137_(_076411_, _079268_, _082214_);
  or g_138138_(_076410_, _079269_, _082215_);
  or g_138139_(_082213_, _082215_, _082216_);
  not g_138140_(_082216_, _082217_);
  or g_138141_(_076417_, _079269_, _082218_);
  or g_138142_(_082213_, _082218_, _082219_);
  not g_138143_(_082219_, _082220_);
  xor g_138144_(_082213_, _082218_, _082222_);
  or g_138145_(_082214_, _082222_, _082223_);
  and g_138146_(_082216_, _082223_, _082224_);
  not g_138147_(_082224_, _082225_);
  and g_138148_(_081151_, _082224_, _082226_);
  or g_138149_(_081150_, _082225_, _082227_);
  xor g_138150_(_081151_, _082224_, _082228_);
  xor g_138151_(_081150_, _082224_, _082229_);
  or g_138152_(_081149_, _082229_, _082230_);
  not g_138153_(_082230_, _082231_);
  xor g_138154_(_081149_, _082228_, _082233_);
  and g_138155_(_079273_, _079277_, _082234_);
  xor g_138156_(_082233_, _082234_, _082235_);
  not g_138157_(_082235_, _082236_);
  or g_138158_(_079280_, _082236_, _082237_);
  not g_138159_(_082237_, _082238_);
  xor g_138160_(_079280_, _082235_, _082239_);
  not g_138161_(_082239_, _082240_);
  or g_138162_(_076439_, _079283_, _082241_);
  not g_138163_(_082241_, _082242_);
  and g_138164_(_079282_, _082241_, _082244_);
  not g_138165_(_082244_, _082245_);
  xor g_138166_(_082239_, _082245_, _082246_);
  or g_138167_(_079284_, _082246_, _082247_);
  xor g_138168_(_079284_, _082246_, _082248_);
  not g_138169_(_082248_, _082249_);
  and g_138170_(_079290_, _082248_, _082250_);
  or g_138171_(_079289_, _082249_, _082251_);
  and g_138172_(_079295_, _082248_, _082252_);
  or g_138173_(_079294_, _082249_, _082253_);
  xor g_138174_(_079294_, _082248_, _082255_);
  and g_138175_(_079289_, _082255_, _082256_);
  or g_138176_(_082250_, _082256_, _082257_);
  or g_138177_(_079300_, _082257_, _082258_);
  xor g_138178_(_079301_, _082257_, _082259_);
  or g_138179_(_079304_, _082259_, _082260_);
  xor g_138180_(_079305_, _082259_, _082261_);
  or g_138181_(_076453_, _079310_, _082262_);
  and g_138182_(_079309_, _082262_, _082263_);
  xor g_138183_(_082261_, _082263_, _082264_);
  and g_138184_(_081148_, _082264_, _082266_);
  not g_138185_(_082266_, _082267_);
  xor g_138186_(_081147_, _082264_, _082268_);
  not g_138187_(_082268_, _082269_);
  and g_138188_(_079315_, _079319_, _082270_);
  xor g_138189_(_082268_, _082270_, _082271_);
  and g_138190_(_079322_, _082271_, _082272_);
  not g_138191_(_082272_, _082273_);
  xor g_138192_(_079322_, _082271_, _082274_);
  and g_138193_(_079326_, _082274_, _082275_);
  not g_138194_(_082275_, _082277_);
  xor g_138195_(_079325_, _082274_, _082278_);
  or g_138196_(_079333_, _082278_, _082279_);
  xor g_138197_(_079334_, _082278_, _082280_);
  not g_138198_(_082280_, _082281_);
  or g_138199_(_079332_, _082280_, _082282_);
  xor g_138200_(_079332_, _082280_, _082283_);
  xor g_138201_(_079332_, _082281_, _082284_);
  or g_138202_(_076476_, _079338_, _082285_);
  or g_138203_(_082284_, _082285_, _082286_);
  xor g_138204_(_082283_, _082285_, _082288_);
  not g_138205_(_082288_, _082289_);
  or g_138206_(_081146_, _082288_, _082290_);
  xor g_138207_(_081146_, _082288_, _082291_);
  xor g_138208_(_081146_, _082289_, _082292_);
  or g_138209_(_079344_, _082292_, _082293_);
  not g_138210_(_082293_, _082294_);
  or g_138211_(_079341_, _082292_, _082295_);
  xor g_138212_(_079341_, _082291_, _082296_);
  or g_138213_(_079346_, _082296_, _082297_);
  not g_138214_(_082297_, _082299_);
  xor g_138215_(_079347_, _082296_, _082300_);
  and g_138216_(_079344_, _082300_, _082301_);
  or g_138217_(_082294_, _082301_, _082302_);
  or g_138218_(_079350_, _082302_, _082303_);
  xor g_138219_(_079352_, _082302_, _082304_);
  and g_138220_(_079354_, _079357_, _082305_);
  not g_138221_(_082305_, _082306_);
  xor g_138222_(_082304_, _082306_, _082307_);
  xor g_138223_(_081145_, _082307_, _082308_);
  not g_138224_(_082308_, _082310_);
  or g_138225_(_081144_, _082310_, _082311_);
  xor g_138226_(_081144_, _082308_, _082312_);
  or g_138227_(_081141_, _082312_, _082313_);
  xor g_138228_(_081142_, _082312_, _082314_);
  or g_138229_(_079368_, _082314_, _082315_);
  xor g_138230_(_079369_, _082314_, _082316_);
  not g_138231_(_082316_, _082317_);
  and g_138232_(_079371_, _079374_, _082318_);
  xor g_138233_(_082317_, _082318_, _082319_);
  xor g_138234_(_082316_, _082318_, _082321_);
  and g_138235_(_079379_, _079382_, _082322_);
  xor g_138236_(_082321_, _082322_, _082323_);
  or g_138237_(_079386_, _082323_, _082324_);
  xor g_138238_(_079386_, _082323_, _082325_);
  not g_138239_(_082325_, _082326_);
  or g_138240_(_079389_, _082326_, _082327_);
  xor g_138241_(_079389_, _082325_, _082328_);
  or g_138242_(_079391_, _082328_, _082329_);
  xor g_138243_(_079391_, _082328_, _082330_);
  xor g_138244_(_079392_, _082328_, _082332_);
  or g_138245_(_079403_, _082332_, _082333_);
  not g_138246_(_082333_, _082334_);
  or g_138247_(_079397_, _082332_, _082335_);
  not g_138248_(_082335_, _082336_);
  and g_138249_(_082333_, _082335_, _082337_);
  or g_138250_(_082334_, _082336_, _082338_);
  and g_138251_(_079397_, _082332_, _082339_);
  or g_138252_(_079396_, _082330_, _082340_);
  and g_138253_(_079403_, _082339_, _082341_);
  or g_138254_(_079402_, _082340_, _082343_);
  and g_138255_(_082337_, _082343_, _082344_);
  or g_138256_(_082338_, _082341_, _082345_);
  or g_138257_(_081139_, _082345_, _082346_);
  not g_138258_(_082346_, _082347_);
  and g_138259_(_079407_, _082345_, _082348_);
  or g_138260_(_079408_, _082344_, _082349_);
  and g_138261_(_081139_, _082348_, _082350_);
  or g_138262_(_081140_, _082349_, _082351_);
  or g_138263_(_079407_, _082345_, _082352_);
  not g_138264_(_082352_, _082354_);
  and g_138265_(_082351_, _082352_, _082355_);
  or g_138266_(_082350_, _082354_, _082356_);
  and g_138267_(_082346_, _082355_, _082357_);
  or g_138268_(_082347_, _082356_, _082358_);
  or g_138269_(_081138_, _082358_, _082359_);
  xor g_138270_(_081138_, _082357_, _082360_);
  or g_138271_(_076555_, _079409_, _082361_);
  and g_138272_(_079413_, _082361_, _082362_);
  xor g_138273_(_082360_, _082362_, _082363_);
  not g_138274_(_082363_, _082365_);
  or g_138275_(_081136_, _082365_, _082366_);
  xor g_138276_(_081136_, _082363_, _082367_);
  or g_138277_(_081134_, _082367_, _082368_);
  xor g_138278_(_081134_, _082367_, _082369_);
  xor g_138279_(_081135_, _082367_, _082370_);
  and g_138280_(_079425_, _082369_, _082371_);
  or g_138281_(_079424_, _082370_, _082372_);
  and g_138282_(_079420_, _082369_, _082373_);
  or g_138283_(_079419_, _082370_, _082374_);
  and g_138284_(_082372_, _082374_, _082376_);
  or g_138285_(_082371_, _082373_, _082377_);
  and g_138286_(_079419_, _082370_, _082378_);
  and g_138287_(_079424_, _082378_, _082379_);
  or g_138288_(_082377_, _082379_, _082380_);
  not g_138289_(_082380_, _082381_);
  xor g_138290_(_081133_, _082380_, _082382_);
  or g_138291_(_079435_, _082382_, _082383_);
  xor g_138292_(_079435_, _082382_, _082384_);
  not g_138293_(_082384_, _082385_);
  or g_138294_(_079442_, _082385_, _082387_);
  xor g_138295_(_079442_, _082384_, _082388_);
  or g_138296_(_079440_, _082388_, _082389_);
  not g_138297_(_082389_, _082390_);
  xor g_138298_(_079441_, _082388_, _082391_);
  or g_138299_(_081130_, _082391_, _082392_);
  xor g_138300_(_081131_, _082391_, _082393_);
  or g_138301_(_079448_, _082393_, _082394_);
  not g_138302_(_082394_, _082395_);
  or g_138303_(_076590_, _079445_, _082396_);
  and g_138304_(_082393_, _082396_, _082398_);
  and g_138305_(_079448_, _082398_, _082399_);
  or g_138306_(_082393_, _082396_, _082400_);
  not g_138307_(_082400_, _082401_);
  or g_138308_(_082399_, _082401_, _082402_);
  or g_138309_(_082395_, _082402_, _082403_);
  or g_138310_(_081128_, _082403_, _082404_);
  xor g_138311_(_081128_, _082403_, _082405_);
  xor g_138312_(_081129_, _082403_, _082406_);
  or g_138313_(_076604_, _079451_, _082407_);
  not g_138314_(_082407_, _082409_);
  and g_138315_(_079459_, _082407_, _082410_);
  xor g_138316_(_082405_, _082410_, _082411_);
  not g_138317_(_082411_, _082412_);
  xor g_138318_(_081127_, _082412_, _082413_);
  or g_138319_(_081124_, _082413_, _082414_);
  not g_138320_(_082414_, _082415_);
  xor g_138321_(_081124_, _082413_, _082416_);
  xor g_138322_(_081125_, _082413_, _082417_);
  or g_138323_(_079467_, _082417_, _082418_);
  not g_138324_(_082418_, _082420_);
  xor g_138325_(_079467_, _082416_, _082421_);
  or g_138326_(_079471_, _082421_, _082422_);
  xor g_138327_(_079470_, _082421_, _082423_);
  or g_138328_(_079476_, _082423_, _082424_);
  xor g_138329_(_079475_, _082423_, _082425_);
  not g_138330_(_082425_, _082426_);
  or g_138331_(_079479_, _082425_, _082427_);
  not g_138332_(_082427_, _082428_);
  xor g_138333_(_079479_, _082425_, _082429_);
  xor g_138334_(_079479_, _082426_, _082431_);
  or g_138335_(_079482_, _082431_, _082432_);
  xor g_138336_(_079482_, _082429_, _082433_);
  not g_138337_(_082433_, _082434_);
  or g_138338_(_076629_, _079486_, _082435_);
  and g_138339_(_079485_, _082435_, _082436_);
  xor g_138340_(_082434_, _082436_, _082437_);
  xor g_138341_(_081123_, _082437_, _082438_);
  not g_138342_(_082438_, _082439_);
  or g_138343_(_079493_, _082439_, _082440_);
  not g_138344_(_082440_, _082442_);
  xor g_138345_(_079493_, _082438_, _082443_);
  or g_138346_(_079497_, _082443_, _082444_);
  not g_138347_(_082444_, _082445_);
  xor g_138348_(_079496_, _082443_, _082446_);
  not g_138349_(_082446_, _082447_);
  or g_138350_(_081120_, _082446_, _082448_);
  not g_138351_(_082448_, _082449_);
  xor g_138352_(_081120_, _082447_, _082450_);
  and g_138353_(_081119_, _082450_, _082451_);
  or g_138354_(_081119_, _082450_, _082453_);
  not g_138355_(_082453_, _082454_);
  xor g_138356_(_081119_, _082450_, _082455_);
  or g_138357_(_082451_, _082454_, _082456_);
  or g_138358_(_081118_, _082456_, _082457_);
  xor g_138359_(_081118_, _082455_, _082458_);
  or g_138360_(_079503_, _082458_, _082459_);
  xor g_138361_(_079503_, _082458_, _082460_);
  not g_138362_(_082460_, _082461_);
  or g_138363_(_079507_, _082461_, _082462_);
  not g_138364_(_082462_, _082464_);
  xor g_138365_(_079507_, _082460_, _082465_);
  not g_138366_(_082465_, _082466_);
  or g_138367_(_079512_, _082465_, _082467_);
  not g_138368_(_082467_, _082468_);
  and g_138369_(_079509_, _082466_, _082469_);
  or g_138370_(_079510_, _082465_, _082470_);
  xor g_138371_(_079509_, _082465_, _082471_);
  and g_138372_(_079512_, _082471_, _082472_);
  or g_138373_(_082468_, _082472_, _082473_);
  not g_138374_(_082473_, _082475_);
  and g_138375_(_079515_, _079519_, _082476_);
  or g_138376_(_082473_, _082476_, _082477_);
  not g_138377_(_082477_, _082478_);
  xor g_138378_(_082475_, _082476_, _082479_);
  not g_138379_(_082479_, _082480_);
  or g_138380_(_081117_, _082479_, _082481_);
  not g_138381_(_082481_, _082482_);
  xor g_138382_(_081117_, _082480_, _082483_);
  or g_138383_(_079529_, _082483_, _082484_);
  not g_138384_(_082484_, _082486_);
  xor g_138385_(_079528_, _082483_, _082487_);
  or g_138386_(_076687_, _079533_, _082488_);
  and g_138387_(_079532_, _082488_, _082489_);
  not g_138388_(_082489_, _082490_);
  xor g_138389_(_082487_, _082489_, _082491_);
  xor g_138390_(_082487_, _082490_, _082492_);
  or g_138391_(_076689_, _079533_, _082493_);
  not g_138392_(_082493_, _082494_);
  and g_138393_(_082492_, _082493_, _082495_);
  and g_138394_(_079537_, _082495_, _082497_);
  and g_138395_(_079539_, _082491_, _082498_);
  or g_138396_(_079537_, _082492_, _082499_);
  and g_138397_(_082491_, _082494_, _082500_);
  not g_138398_(_082500_, _082501_);
  or g_138399_(_082498_, _082500_, _082502_);
  or g_138400_(_082497_, _082502_, _082503_);
  or g_138401_(_079542_, _082503_, _082504_);
  xor g_138402_(_079543_, _082503_, _082505_);
  or g_138403_(_079546_, _082505_, _082506_);
  xor g_138404_(_079546_, _082505_, _082508_);
  xor g_138405_(_079547_, _082505_, _082509_);
  and g_138406_(_079552_, _082508_, _082510_);
  or g_138407_(_079551_, _082509_, _082511_);
  xor g_138408_(_079552_, _082508_, _082512_);
  and g_138409_(_079556_, _082512_, _082513_);
  not g_138410_(_082513_, _082514_);
  xor g_138411_(_079556_, _082512_, _082515_);
  xor g_138412_(_079555_, _082512_, _082516_);
  and g_138413_(_079561_, _082516_, _082517_);
  and g_138414_(_079564_, _082517_, _082519_);
  and g_138415_(_079562_, _082512_, _082520_);
  not g_138416_(_082520_, _082521_);
  and g_138417_(_079565_, _082515_, _082522_);
  not g_138418_(_082522_, _082523_);
  or g_138419_(_082520_, _082522_, _082524_);
  or g_138420_(_082519_, _082524_, _082525_);
  not g_138421_(_082525_, _082526_);
  and g_138422_(_079568_, _082526_, _082527_);
  or g_138423_(_079569_, _082525_, _082528_);
  xor g_138424_(_079569_, _082525_, _082530_);
  xor g_138425_(_079568_, _082525_, _082531_);
  and g_138426_(_081116_, _082530_, _082532_);
  or g_138427_(_081115_, _082531_, _082533_);
  xor g_138428_(_081115_, _082530_, _082534_);
  or g_138429_(_081113_, _082534_, _082535_);
  not g_138430_(_082535_, _082536_);
  xor g_138431_(_081113_, _082534_, _082537_);
  xor g_138432_(_081114_, _082534_, _082538_);
  and g_138433_(_079576_, _079583_, _082539_);
  xor g_138434_(_082537_, _082539_, _082541_);
  or g_138435_(_079578_, _082541_, _082542_);
  not g_138436_(_082542_, _082543_);
  xor g_138437_(_079578_, _082541_, _082544_);
  not g_138438_(_082544_, _082545_);
  or g_138439_(_079587_, _082545_, _082546_);
  not g_138440_(_082546_, _082547_);
  xor g_138441_(_079587_, _082544_, _082548_);
  xor g_138442_(_079594_, _082548_, _082549_);
  xor g_138443_(_081112_, _082549_, _082550_);
  and g_138444_(_079603_, _082550_, _082552_);
  and g_138445_(_079608_, _082552_, _082553_);
  or g_138446_(_079608_, _082550_, _082554_);
  not g_138447_(_082554_, _082555_);
  or g_138448_(_079603_, _082550_, _082556_);
  not g_138449_(_082556_, _082557_);
  or g_138450_(_082555_, _082557_, _082558_);
  or g_138451_(_082553_, _082558_, _082559_);
  or g_138452_(_073863_, _081107_, _082560_);
  and g_138453_(_079610_, _082560_, _082561_);
  or g_138454_(_082559_, _082561_, _082563_);
  xor g_138455_(_082559_, _082561_, _082564_);
  not g_138456_(_082564_, _082565_);
  and g_138457_(_081109_, _082564_, _082566_);
  or g_138458_(_081108_, _082565_, _082567_);
  xor g_138459_(_081108_, _082564_, _082568_);
  or g_138460_(_081106_, _082568_, _082569_);
  not g_138461_(_082569_, _082570_);
  xor g_138462_(_081105_, _082568_, _082571_);
  not g_138463_(_082571_, _082572_);
  and g_138464_(_079616_, _082572_, _082574_);
  or g_138465_(_079617_, _082571_, _082575_);
  xor g_138466_(_079616_, _082571_, _082576_);
  and g_138467_(_079619_, _079621_, _082577_);
  not g_138468_(_082577_, _082578_);
  xor g_138469_(_082576_, _082578_, _082579_);
  xor g_138470_(_082576_, _082577_, _082580_);
  and g_138471_(_079625_, _082579_, _082581_);
  or g_138472_(_079624_, _082580_, _082582_);
  or g_138473_(_076775_, _079618_, _082583_);
  or g_138474_(_082579_, _082583_, _082585_);
  not g_138475_(_082585_, _082586_);
  and g_138476_(_082582_, _082585_, _082587_);
  or g_138477_(_082581_, _082586_, _082588_);
  and g_138478_(_079628_, _079630_, _082589_);
  xor g_138479_(_082588_, _082589_, _082590_);
  xor g_138480_(_082587_, _082589_, _082591_);
  or g_138481_(_081104_, _082591_, _082592_);
  xor g_138482_(_081104_, _082591_, _082593_);
  xor g_138483_(_081104_, _082590_, _082594_);
  or g_138484_(_076794_, _079631_, _082596_);
  and g_138485_(_079635_, _082596_, _082597_);
  xor g_138486_(_082593_, _082597_, _082598_);
  and g_138487_(_079639_, _082598_, _082599_);
  or g_138488_(_079639_, _082598_, _082600_);
  not g_138489_(_082600_, _082601_);
  xor g_138490_(_079639_, _082598_, _082602_);
  or g_138491_(_082599_, _082601_, _082603_);
  and g_138492_(_079643_, _079645_, _082604_);
  xor g_138493_(_082602_, _082604_, _082605_);
  or g_138494_(_081103_, _082605_, _082607_);
  xor g_138495_(_081103_, _082605_, _082608_);
  not g_138496_(_082608_, _082609_);
  and g_138497_(_081102_, _082608_, _082610_);
  or g_138498_(_081101_, _082609_, _082611_);
  xor g_138499_(_081101_, _082608_, _082612_);
  or g_138500_(_081100_, _082612_, _082613_);
  not g_138501_(_082613_, _082614_);
  xor g_138502_(_081098_, _082612_, _082615_);
  or g_138503_(_081097_, _082615_, _082616_);
  not g_138504_(_082616_, _082618_);
  xor g_138505_(_081096_, _082615_, _082619_);
  not g_138506_(_082619_, _082620_);
  or g_138507_(_081095_, _082619_, _082621_);
  xor g_138508_(_081095_, _082620_, _082622_);
  or g_138509_(_079652_, _082622_, _082623_);
  xor g_138510_(_079653_, _082622_, _082624_);
  or g_138511_(_079655_, _082624_, _082625_);
  not g_138512_(_082625_, _082626_);
  xor g_138513_(_079655_, _082624_, _082627_);
  xor g_138514_(_079656_, _082624_, _082629_);
  and g_138515_(_079658_, _079661_, _082630_);
  xor g_138516_(_082627_, _082630_, _082631_);
  or g_138517_(_079663_, _082631_, _082632_);
  xor g_138518_(_079663_, _082631_, _082633_);
  and g_138519_(_079672_, _082633_, _082634_);
  not g_138520_(_082634_, _082635_);
  xor g_138521_(_079671_, _082633_, _082636_);
  or g_138522_(_079676_, _082636_, _082637_);
  not g_138523_(_082637_, _082638_);
  xor g_138524_(_079675_, _082636_, _082640_);
  not g_138525_(_082640_, _082641_);
  or g_138526_(_079683_, _082640_, _082642_);
  not g_138527_(_082642_, _082643_);
  or g_138528_(_079678_, _082640_, _082644_);
  xor g_138529_(_079678_, _082640_, _082645_);
  xor g_138530_(_079678_, _082641_, _082646_);
  and g_138531_(_079683_, _082646_, _082647_);
  or g_138532_(_079682_, _082645_, _082648_);
  and g_138533_(_082642_, _082648_, _082649_);
  or g_138534_(_082643_, _082647_, _082651_);
  xor g_138535_(_079687_, _082649_, _082652_);
  xor g_138536_(_079687_, _082651_, _082653_);
  and g_138537_(_079691_, _082653_, _082654_);
  not g_138538_(_082654_, _082655_);
  xor g_138539_(_079690_, _082652_, _082656_);
  not g_138540_(_082656_, _082657_);
  and g_138541_(_079695_, _082656_, _082658_);
  or g_138542_(_079694_, _082657_, _082659_);
  xor g_138543_(_079694_, _082656_, _082660_);
  or g_138544_(_079699_, _082660_, _082662_);
  xor g_138545_(_079698_, _082660_, _082663_);
  not g_138546_(_082663_, _082664_);
  or g_138547_(_079704_, _082663_, _082665_);
  xor g_138548_(_079704_, _082663_, _082666_);
  xor g_138549_(_079704_, _082664_, _082667_);
  or g_138550_(_081094_, _082667_, _082668_);
  not g_138551_(_082668_, _082669_);
  xor g_138552_(_081094_, _082666_, _082670_);
  or g_138553_(_081092_, _082670_, _082671_);
  not g_138554_(_082671_, _082673_);
  xor g_138555_(_081092_, _082670_, _082674_);
  xor g_138556_(_081093_, _082670_, _082675_);
  and g_138557_(_079713_, _082674_, _082676_);
  or g_138558_(_079715_, _082675_, _082677_);
  or g_138559_(_079710_, _082675_, _082678_);
  not g_138560_(_082678_, _082679_);
  and g_138561_(_082677_, _082678_, _082680_);
  or g_138562_(_082676_, _082679_, _082681_);
  and g_138563_(_079710_, _082675_, _082682_);
  or g_138564_(_079709_, _082674_, _082684_);
  and g_138565_(_079715_, _082682_, _082685_);
  or g_138566_(_079713_, _082684_, _082686_);
  and g_138567_(_082680_, _082686_, _082687_);
  or g_138568_(_082681_, _082685_, _082688_);
  and g_138569_(_079719_, _082687_, _082689_);
  or g_138570_(_079718_, _082688_, _082690_);
  xor g_138571_(_079719_, _082687_, _082691_);
  xor g_138572_(_079718_, _082687_, _082692_);
  or g_138573_(_079723_, _082692_, _082693_);
  not g_138574_(_082693_, _082695_);
  xor g_138575_(_079723_, _082692_, _082696_);
  xor g_138576_(_079723_, _082691_, _082697_);
  and g_138577_(_079727_, _079729_, _082698_);
  xor g_138578_(_082696_, _082698_, _082699_);
  xor g_138579_(_082697_, _082698_, _082700_);
  and g_138580_(_079742_, _082700_, _082701_);
  not g_138581_(_082701_, _082702_);
  and g_138582_(_079733_, _082699_, _082703_);
  and g_138583_(_079743_, _082703_, _082704_);
  and g_138584_(_079732_, _082700_, _082706_);
  not g_138585_(_082706_, _082707_);
  or g_138586_(_082704_, _082706_, _082708_);
  or g_138587_(_082701_, _082708_, _082709_);
  or g_138588_(_079740_, _082709_, _082710_);
  xor g_138589_(_079741_, _082709_, _082711_);
  or g_138590_(_081090_, _082711_, _082712_);
  xor g_138591_(_081091_, _082711_, _082713_);
  not g_138592_(_082713_, _082714_);
  or g_138593_(_081089_, _082713_, _082715_);
  xor g_138594_(_081089_, _082713_, _082717_);
  xor g_138595_(_081089_, _082714_, _082718_);
  or g_138596_(_081087_, _082718_, _082719_);
  xor g_138597_(_081087_, _082717_, _082720_);
  or g_138598_(_081086_, _082720_, _082721_);
  xor g_138599_(_081086_, _082720_, _082722_);
  not g_138600_(_082722_, _082723_);
  or g_138601_(_081085_, _082723_, _082724_);
  not g_138602_(_082724_, _082725_);
  xor g_138603_(_081085_, _082722_, _082726_);
  not g_138604_(_082726_, _082728_);
  or g_138605_(_081084_, _082726_, _082729_);
  xor g_138606_(_081084_, _082726_, _082730_);
  xor g_138607_(_081084_, _082728_, _082731_);
  and g_138608_(_079753_, _079755_, _082732_);
  xor g_138609_(_082730_, _082732_, _082733_);
  or g_138610_(_081083_, _082733_, _082734_);
  not g_138611_(_082734_, _082735_);
  xor g_138612_(_081083_, _082733_, _082736_);
  not g_138613_(_082736_, _082737_);
  and g_138614_(_081082_, _082736_, _082739_);
  or g_138615_(_081081_, _082737_, _082740_);
  xor g_138616_(_081081_, _082736_, _082741_);
  or g_138617_(_081078_, _082741_, _082742_);
  xor g_138618_(_081079_, _082741_, _082743_);
  or g_138619_(_079768_, _082743_, _082744_);
  not g_138620_(_082744_, _082745_);
  and g_138621_(_079764_, _082743_, _082746_);
  and g_138622_(_079768_, _082746_, _082747_);
  or g_138623_(_079764_, _082743_, _082748_);
  not g_138624_(_082748_, _082750_);
  or g_138625_(_082747_, _082750_, _082751_);
  or g_138626_(_082745_, _082751_, _082752_);
  and g_138627_(_079773_, _082752_, _082753_);
  or g_138628_(_079773_, _082752_, _082754_);
  not g_138629_(_082754_, _082755_);
  xor g_138630_(_079773_, _082752_, _082756_);
  or g_138631_(_082753_, _082755_, _082757_);
  xor g_138632_(_081076_, _082756_, _082758_);
  or g_138633_(_079781_, _082758_, _082759_);
  not g_138634_(_082759_, _082761_);
  xor g_138635_(_079781_, _082758_, _082762_);
  xor g_138636_(_079782_, _082758_, _082763_);
  and g_138637_(_078278_, _079778_, _082764_);
  and g_138638_(_082762_, _082764_, _082765_);
  not g_138639_(_082765_, _082766_);
  and g_138640_(_079784_, _082763_, _082767_);
  or g_138641_(_082765_, _082767_, _082768_);
  or g_138642_(_081074_, _082768_, _082769_);
  xor g_138643_(_081075_, _082768_, _082770_);
  or g_138644_(_081072_, _082770_, _082772_);
  xor g_138645_(_081073_, _082770_, _082773_);
  and g_138646_(_079789_, _079794_, _082774_);
  not g_138647_(_082774_, _082775_);
  or g_138648_(_082773_, _082774_, _082776_);
  not g_138649_(_082776_, _082777_);
  xor g_138650_(_082773_, _082775_, _082778_);
  or g_138651_(_079797_, _082778_, _082779_);
  xor g_138652_(_079797_, _082778_, _082780_);
  xor g_138653_(_079798_, _082778_, _082781_);
  and g_138654_(_079801_, _082780_, _082783_);
  or g_138655_(_079800_, _082781_, _082784_);
  xor g_138656_(_079801_, _082780_, _082785_);
  or g_138657_(_076986_, _079806_, _082786_);
  not g_138658_(_082786_, _082787_);
  and g_138659_(_079804_, _082786_, _082788_);
  xor g_138660_(_082785_, _082788_, _082789_);
  or g_138661_(_081070_, _082789_, _082790_);
  xor g_138662_(_081071_, _082789_, _082791_);
  not g_138663_(_082791_, _082792_);
  or g_138664_(_079815_, _082791_, _082794_);
  not g_138665_(_082794_, _082795_);
  or g_138666_(_079811_, _082791_, _082796_);
  xor g_138667_(_079811_, _082791_, _082797_);
  xor g_138668_(_079811_, _082792_, _082798_);
  and g_138669_(_079815_, _082798_, _082799_);
  or g_138670_(_079816_, _082797_, _082800_);
  and g_138671_(_082794_, _082800_, _082801_);
  or g_138672_(_082795_, _082799_, _082802_);
  and g_138673_(_079818_, _079822_, _082803_);
  xor g_138674_(_082801_, _082803_, _082805_);
  not g_138675_(_082805_, _082806_);
  or g_138676_(_077001_, _079827_, _082807_);
  and g_138677_(_079826_, _082807_, _082808_);
  or g_138678_(_082805_, _082808_, _082809_);
  not g_138679_(_082809_, _082810_);
  xor g_138680_(_082806_, _082808_, _082811_);
  not g_138681_(_082811_, _082812_);
  xor g_138682_(_081069_, _082812_, _082813_);
  not g_138683_(_082813_, _082814_);
  or g_138684_(_077011_, _079834_, _082816_);
  and g_138685_(_079836_, _082816_, _082817_);
  xor g_138686_(_082813_, _082817_, _082818_);
  not g_138687_(_082818_, _082819_);
  or g_138688_(_077018_, _079841_, _082820_);
  not g_138689_(_082820_, _082821_);
  or g_138690_(_077014_, _079838_, _082822_);
  not g_138691_(_082822_, _082823_);
  and g_138692_(_082820_, _082822_, _082824_);
  xor g_138693_(_082818_, _082824_, _082825_);
  or g_138694_(_081065_, _082825_, _082827_);
  or g_138695_(_077019_, _079841_, _082828_);
  or g_138696_(_082825_, _082828_, _082829_);
  xor g_138697_(_082825_, _082828_, _082830_);
  not g_138698_(_082830_, _082831_);
  or g_138699_(_081067_, _082830_, _082832_);
  and g_138700_(_082827_, _082832_, _082833_);
  not g_138701_(_082833_, _082834_);
  xor g_138702_(_081063_, _082833_, _082835_);
  or g_138703_(_081062_, _082835_, _082836_);
  xor g_138704_(_081062_, _082835_, _082838_);
  xor g_138705_(_081061_, _082838_, _082839_);
  or g_138706_(_081060_, _082839_, _082840_);
  not g_138707_(_082840_, _082841_);
  xor g_138708_(_081060_, _082839_, _082842_);
  not g_138709_(_082842_, _082843_);
  and g_138710_(_079852_, _082842_, _082844_);
  or g_138711_(_079851_, _082843_, _082845_);
  xor g_138712_(_079851_, _082842_, _082846_);
  or g_138713_(_079855_, _082846_, _082847_);
  not g_138714_(_082847_, _082849_);
  xor g_138715_(_079856_, _082846_, _082850_);
  or g_138716_(_079858_, _082850_, _082851_);
  not g_138717_(_082851_, _082852_);
  xor g_138718_(_079859_, _082850_, _082853_);
  and g_138719_(_081059_, _082853_, _082854_);
  or g_138720_(_081059_, _082853_, _082855_);
  not g_138721_(_082855_, _082856_);
  xor g_138722_(_081059_, _082853_, _082857_);
  or g_138723_(_082854_, _082856_, _082858_);
  or g_138724_(_077049_, _079862_, _082860_);
  or g_138725_(_074170_, _081058_, _082861_);
  and g_138726_(_082860_, _082861_, _082862_);
  xor g_138727_(_082857_, _082862_, _082863_);
  or g_138728_(_081057_, _082863_, _082864_);
  xor g_138729_(_081057_, _082863_, _082865_);
  not g_138730_(_082865_, _082866_);
  or g_138731_(_079867_, _082866_, _082867_);
  xor g_138732_(_079867_, _082865_, _082868_);
  and g_138733_(_079870_, _082868_, _082869_);
  and g_138734_(_079872_, _082869_, _082871_);
  or g_138735_(_079872_, _082868_, _082872_);
  not g_138736_(_082872_, _082873_);
  or g_138737_(_079870_, _082868_, _082874_);
  and g_138738_(_082872_, _082874_, _082875_);
  not g_138739_(_082875_, _082876_);
  or g_138740_(_082871_, _082876_, _082877_);
  or g_138741_(_079877_, _082877_, _082878_);
  not g_138742_(_082878_, _082879_);
  or g_138743_(_079874_, _082877_, _082880_);
  xor g_138744_(_079874_, _082877_, _082882_);
  xor g_138745_(_079875_, _082877_, _082883_);
  or g_138746_(_079881_, _082883_, _082884_);
  xor g_138747_(_079881_, _082882_, _082885_);
  and g_138748_(_079877_, _082885_, _082886_);
  or g_138749_(_082879_, _082886_, _082887_);
  not g_138750_(_082887_, _082888_);
  and g_138751_(_081054_, _082888_, _082889_);
  or g_138752_(_081056_, _082887_, _082890_);
  xor g_138753_(_081056_, _082887_, _082891_);
  xor g_138754_(_081054_, _082887_, _082893_);
  and g_138755_(_079884_, _079886_, _082894_);
  xor g_138756_(_082891_, _082894_, _082895_);
  not g_138757_(_082895_, _082896_);
  or g_138758_(_081053_, _082895_, _082897_);
  xor g_138759_(_081053_, _082895_, _082898_);
  xor g_138760_(_081053_, _082896_, _082899_);
  or g_138761_(_081052_, _082899_, _082900_);
  xor g_138762_(_081052_, _082898_, _082901_);
  or g_138763_(_079893_, _082901_, _082902_);
  not g_138764_(_082902_, _082904_);
  xor g_138765_(_079894_, _082901_, _082905_);
  or g_138766_(_079898_, _082905_, _082906_);
  xor g_138767_(_079897_, _082905_, _082907_);
  not g_138768_(_082907_, _082908_);
  and g_138769_(_079900_, _079905_, _082909_);
  or g_138770_(_082907_, _082909_, _082910_);
  not g_138771_(_082910_, _082911_);
  xor g_138772_(_082908_, _082909_, _082912_);
  not g_138773_(_082912_, _082913_);
  or g_138774_(_077112_, _079910_, _082915_);
  and g_138775_(_079909_, _082915_, _082916_);
  xor g_138776_(_082912_, _082916_, _082917_);
  xor g_138777_(_082913_, _082916_, _082918_);
  or g_138778_(_081051_, _082918_, _082919_);
  xor g_138779_(_081051_, _082917_, _082920_);
  or g_138780_(_079916_, _079918_, _082921_);
  xor g_138781_(_082920_, _082921_, _082922_);
  not g_138782_(_082922_, _082923_);
  or g_138783_(_079921_, _082922_, _082924_);
  not g_138784_(_082924_, _082926_);
  xor g_138785_(_079921_, _082922_, _082927_);
  xor g_138786_(_079921_, _082923_, _082928_);
  and g_138787_(_079925_, _082927_, _082929_);
  or g_138788_(_079924_, _082928_, _082930_);
  xor g_138789_(_079925_, _082927_, _082931_);
  xor g_138790_(_081050_, _082931_, _082932_);
  or g_138791_(_081049_, _082932_, _082933_);
  not g_138792_(_082933_, _082934_);
  xor g_138793_(_081049_, _082932_, _082935_);
  not g_138794_(_082935_, _082937_);
  xor g_138795_(_079933_, _082935_, _082938_);
  or g_138796_(_079937_, _082938_, _082939_);
  not g_138797_(_082939_, _082940_);
  and g_138798_(_079937_, _082938_, _082941_);
  xor g_138799_(_079937_, _082938_, _082942_);
  or g_138800_(_082940_, _082941_, _082943_);
  or g_138801_(_079940_, _082943_, _082944_);
  xor g_138802_(_079940_, _082942_, _082945_);
  not g_138803_(_082945_, _082946_);
  or g_138804_(_079942_, _082945_, _082948_);
  xor g_138805_(_079942_, _082946_, _082949_);
  or g_138806_(_079949_, _082949_, _082950_);
  not g_138807_(_082950_, _082951_);
  and g_138808_(_079946_, _082949_, _082952_);
  and g_138809_(_079949_, _082952_, _082953_);
  or g_138810_(_079946_, _082949_, _082954_);
  not g_138811_(_082954_, _082955_);
  or g_138812_(_082953_, _082955_, _082956_);
  or g_138813_(_082951_, _082956_, _082957_);
  and g_138814_(_079951_, _079955_, _082959_);
  not g_138815_(_082959_, _082960_);
  xor g_138816_(_082957_, _082960_, _082961_);
  or g_138817_(_079959_, _082961_, _082962_);
  not g_138818_(_082962_, _082963_);
  xor g_138819_(_079959_, _082961_, _082964_);
  not g_138820_(_082964_, _082965_);
  or g_138821_(_079962_, _082965_, _082966_);
  not g_138822_(_082966_, _082967_);
  xor g_138823_(_079962_, _082964_, _082968_);
  or g_138824_(_079964_, _082968_, _082970_);
  xor g_138825_(_079965_, _082968_, _082971_);
  not g_138826_(_082971_, _082972_);
  or g_138827_(_079968_, _082971_, _082973_);
  xor g_138828_(_079968_, _082971_, _082974_);
  xor g_138829_(_079968_, _082972_, _082975_);
  or g_138830_(_079971_, _082975_, _082976_);
  xor g_138831_(_079971_, _082974_, _082977_);
  or g_138832_(_077175_, _079974_, _082978_);
  and g_138833_(_079973_, _082978_, _082979_);
  and g_138834_(_082977_, _082979_, _082981_);
  or g_138835_(_082977_, _082979_, _082982_);
  not g_138836_(_082982_, _082983_);
  xor g_138837_(_082977_, _082979_, _082984_);
  or g_138838_(_082981_, _082983_, _082985_);
  or g_138839_(_081048_, _082985_, _082986_);
  xor g_138840_(_081048_, _082984_, _082987_);
  and g_138841_(_079979_, _082987_, _082988_);
  and g_138842_(_081047_, _082988_, _082989_);
  not g_138843_(_082989_, _082990_);
  or g_138844_(_079979_, _082987_, _082992_);
  or g_138845_(_081047_, _082987_, _082993_);
  not g_138846_(_082993_, _082994_);
  and g_138847_(_082992_, _082993_, _082995_);
  not g_138848_(_082995_, _082996_);
  and g_138849_(_082990_, _082995_, _082997_);
  or g_138850_(_082989_, _082996_, _082998_);
  or g_138851_(_081046_, _082998_, _082999_);
  xor g_138852_(_081046_, _082997_, _083000_);
  or g_138853_(_079984_, _083000_, _083001_);
  xor g_138854_(_079985_, _083000_, _083003_);
  or g_138855_(_074322_, _077190_, _083004_);
  or g_138856_(_079986_, _083004_, _083005_);
  not g_138857_(_083005_, _083006_);
  or g_138858_(_083003_, _083005_, _083007_);
  xor g_138859_(_083003_, _083006_, _083008_);
  not g_138860_(_083008_, _083009_);
  or g_138861_(_079992_, _083008_, _083010_);
  not g_138862_(_083010_, _083011_);
  xor g_138863_(_079992_, _083008_, _083012_);
  xor g_138864_(_079992_, _083009_, _083014_);
  or g_138865_(_079996_, _083014_, _083015_);
  not g_138866_(_083015_, _083016_);
  xor g_138867_(_079997_, _083012_, _083017_);
  not g_138868_(_083017_, _083018_);
  and g_138869_(_080001_, _083017_, _083019_);
  or g_138870_(_079999_, _083018_, _083020_);
  xor g_138871_(_079999_, _083017_, _083021_);
  or g_138872_(_080003_, _083021_, _083022_);
  xor g_138873_(_080004_, _083021_, _083023_);
  and g_138874_(_080007_, _080010_, _083025_);
  xor g_138875_(_083023_, _083025_, _083026_);
  not g_138876_(_083026_, _083027_);
  or g_138877_(_080014_, _083027_, _083028_);
  not g_138878_(_083028_, _083029_);
  xor g_138879_(_080014_, _083026_, _083030_);
  and g_138880_(_077206_, _080016_, _083031_);
  or g_138881_(_077208_, _080015_, _083032_);
  or g_138882_(_083030_, _083032_, _083033_);
  not g_138883_(_083033_, _083034_);
  xor g_138884_(_083030_, _083031_, _083036_);
  not g_138885_(_083036_, _083037_);
  or g_138886_(_081045_, _083036_, _083038_);
  not g_138887_(_083038_, _083039_);
  xor g_138888_(_081045_, _083037_, _083040_);
  not g_138889_(_083040_, _083041_);
  and g_138890_(_080020_, _080025_, _083042_);
  xor g_138891_(_083041_, _083042_, _083043_);
  or g_138892_(_080028_, _083043_, _083044_);
  xor g_138893_(_080029_, _083043_, _083045_);
  not g_138894_(_083045_, _083047_);
  and g_138895_(_080032_, _080037_, _083048_);
  xor g_138896_(_083047_, _083048_, _083049_);
  xor g_138897_(_083045_, _083048_, _083050_);
  or g_138898_(_080040_, _083049_, _083051_);
  xor g_138899_(_080040_, _083049_, _083052_);
  xor g_138900_(_080040_, _083050_, _083053_);
  or g_138901_(_081043_, _083053_, _083054_);
  xor g_138902_(_081043_, _083052_, _083055_);
  or g_138903_(_081042_, _083055_, _083056_);
  not g_138904_(_083056_, _083058_);
  xor g_138905_(_081042_, _083055_, _083059_);
  not g_138906_(_083059_, _083060_);
  and g_138907_(_080046_, _083059_, _083061_);
  or g_138908_(_080045_, _083060_, _083062_);
  xor g_138909_(_080045_, _083059_, _083063_);
  not g_138910_(_083063_, _083064_);
  and g_138911_(_080048_, _080051_, _083065_);
  xor g_138912_(_083063_, _083065_, _083066_);
  xor g_138913_(_083064_, _083065_, _083067_);
  xor g_138914_(_081041_, _083066_, _083069_);
  or g_138915_(_081039_, _083069_, _083070_);
  xor g_138916_(_081039_, _083069_, _083071_);
  not g_138917_(_083071_, _083072_);
  or g_138918_(_081038_, _083072_, _083073_);
  xor g_138919_(_081038_, _083071_, _083074_);
  not g_138920_(_083074_, _083075_);
  or g_138921_(_077260_, _080060_, _083076_);
  and g_138922_(_080059_, _083076_, _083077_);
  xor g_138923_(_083075_, _083077_, _083078_);
  xor g_138924_(_081037_, _083078_, _083080_);
  or g_138925_(_080067_, _083080_, _083081_);
  not g_138926_(_083081_, _083082_);
  xor g_138927_(_080067_, _083080_, _083083_);
  xor g_138928_(_080074_, _083083_, _083084_);
  not g_138929_(_083084_, _083085_);
  or g_138930_(_080078_, _083084_, _083086_);
  not g_138931_(_083086_, _083087_);
  xor g_138932_(_080078_, _083085_, _083088_);
  or g_138933_(_081034_, _083088_, _083089_);
  xor g_138934_(_081032_, _083088_, _083091_);
  or g_138935_(_080081_, _083091_, _083092_);
  xor g_138936_(_080081_, _083091_, _083093_);
  not g_138937_(_083093_, _083094_);
  and g_138938_(_080084_, _080090_, _083095_);
  xor g_138939_(_083093_, _083095_, _083096_);
  or g_138940_(_081031_, _083096_, _083097_);
  xor g_138941_(_081031_, _083096_, _083098_);
  not g_138942_(_083098_, _083099_);
  xor g_138943_(_081030_, _083098_, _083100_);
  or g_138944_(_080107_, _083100_, _083102_);
  xor g_138945_(_080106_, _083100_, _083103_);
  not g_138946_(_083103_, _083104_);
  and g_138947_(_081029_, _083104_, _083105_);
  not g_138948_(_083105_, _083106_);
  xor g_138949_(_081029_, _083103_, _083107_);
  not g_138950_(_083107_, _083108_);
  or g_138951_(_081028_, _083107_, _083109_);
  xor g_138952_(_081028_, _083107_, _083110_);
  xor g_138953_(_081028_, _083108_, _083111_);
  or g_138954_(_081027_, _083111_, _083113_);
  xor g_138955_(_081027_, _083110_, _083114_);
  or g_138956_(_080116_, _083114_, _083115_);
  or g_138957_(_080113_, _083114_, _083116_);
  and g_138958_(_083115_, _083116_, _083117_);
  not g_138959_(_083117_, _083118_);
  and g_138960_(_080113_, _083114_, _083119_);
  and g_138961_(_080116_, _083119_, _083120_);
  or g_138962_(_083118_, _083120_, _083121_);
  or g_138963_(_080119_, _083121_, _083122_);
  xor g_138964_(_080119_, _083121_, _083124_);
  not g_138965_(_083124_, _083125_);
  or g_138966_(_080122_, _083125_, _083126_);
  xor g_138967_(_080122_, _083124_, _083127_);
  not g_138968_(_083127_, _083128_);
  and g_138969_(_080124_, _080127_, _083129_);
  xor g_138970_(_083128_, _083129_, _083130_);
  not g_138971_(_083130_, _083131_);
  or g_138972_(_080129_, _083130_, _083132_);
  xor g_138973_(_080129_, _083130_, _083133_);
  xor g_138974_(_080129_, _083131_, _083135_);
  and g_138975_(_080131_, _080134_, _083136_);
  xor g_138976_(_083133_, _083136_, _083137_);
  and g_138977_(_081026_, _083137_, _083138_);
  or g_138978_(_077358_, _080130_, _083139_);
  or g_138979_(_083137_, _083139_, _083140_);
  not g_138980_(_083140_, _083141_);
  or g_138981_(_083138_, _083141_, _083142_);
  or g_138982_(_080135_, _080137_, _083143_);
  and g_138983_(_080140_, _083143_, _083144_);
  xor g_138984_(_083142_, _083144_, _083146_);
  and g_138985_(_080142_, _083146_, _083147_);
  not g_138986_(_083147_, _083148_);
  xor g_138987_(_080144_, _083146_, _083149_);
  not g_138988_(_083149_, _083150_);
  or g_138989_(_080147_, _083149_, _083151_);
  not g_138990_(_083151_, _083152_);
  xor g_138991_(_080147_, _083149_, _083153_);
  xor g_138992_(_080147_, _083150_, _083154_);
  or g_138993_(_077368_, _080148_, _083155_);
  not g_138994_(_083155_, _083157_);
  and g_138995_(_083153_, _083157_, _083158_);
  or g_138996_(_083154_, _083155_, _083159_);
  xor g_138997_(_083153_, _083155_, _083160_);
  or g_138998_(_081024_, _083160_, _083161_);
  not g_138999_(_083161_, _083162_);
  xor g_139000_(_081025_, _083160_, _083163_);
  not g_139001_(_083163_, _083164_);
  or g_139002_(_080153_, _080156_, _083165_);
  and g_139003_(_080152_, _083165_, _083166_);
  xor g_139004_(_083163_, _083166_, _083168_);
  xor g_139005_(_083164_, _083166_, _083169_);
  or g_139006_(_081023_, _083169_, _083170_);
  xor g_139007_(_081023_, _083168_, _083171_);
  or g_139008_(_081021_, _083171_, _083172_);
  not g_139009_(_083172_, _083173_);
  xor g_139010_(_081021_, _083171_, _083174_);
  and g_139011_(_081020_, _083174_, _083175_);
  not g_139012_(_083175_, _083176_);
  xor g_139013_(_081020_, _083174_, _083177_);
  xor g_139014_(_081019_, _083174_, _083179_);
  or g_139015_(_078225_, _080158_, _083180_);
  and g_139016_(_080162_, _083180_, _083181_);
  xor g_139017_(_083177_, _083181_, _083182_);
  not g_139018_(_083182_, _083183_);
  or g_139019_(_081018_, _083182_, _083184_);
  xor g_139020_(_081018_, _083182_, _083185_);
  xor g_139021_(_081018_, _083183_, _083186_);
  or g_139022_(_081017_, _083186_, _083187_);
  not g_139023_(_083187_, _083188_);
  xor g_139024_(_081017_, _083185_, _083190_);
  or g_139025_(_080168_, _083190_, _083191_);
  xor g_139026_(_080169_, _083190_, _083192_);
  and g_139027_(_080172_, _083192_, _083193_);
  or g_139028_(_080172_, _083192_, _083194_);
  xor g_139029_(_080173_, _083192_, _083195_);
  not g_139030_(_083195_, _083196_);
  and g_139031_(_080177_, _080181_, _083197_);
  xor g_139032_(_083196_, _083197_, _083198_);
  or g_139033_(_080184_, _083198_, _083199_);
  xor g_139034_(_080184_, _083198_, _083201_);
  xor g_139035_(_080185_, _083198_, _083202_);
  and g_139036_(_080189_, _083201_, _083203_);
  or g_139037_(_080188_, _083202_, _083204_);
  xor g_139038_(_080189_, _083201_, _083205_);
  xor g_139039_(_080188_, _083201_, _083206_);
  and g_139040_(_080193_, _083205_, _083207_);
  or g_139041_(_080192_, _083206_, _083208_);
  xor g_139042_(_080192_, _083205_, _083209_);
  or g_139043_(_080196_, _083209_, _083210_);
  not g_139044_(_083210_, _083212_);
  xor g_139045_(_080196_, _083209_, _083213_);
  and g_139046_(_080201_, _083213_, _083214_);
  xor g_139047_(_080200_, _083213_, _083215_);
  or g_139048_(_080205_, _083215_, _083216_);
  xor g_139049_(_080205_, _083215_, _083217_);
  not g_139050_(_083217_, _083218_);
  or g_139051_(_080208_, _083218_, _083219_);
  not g_139052_(_083219_, _083220_);
  xor g_139053_(_080208_, _083217_, _083221_);
  or g_139054_(_080213_, _083221_, _083223_);
  not g_139055_(_083223_, _083224_);
  xor g_139056_(_080212_, _083221_, _083225_);
  not g_139057_(_083225_, _083226_);
  and g_139058_(_080216_, _083226_, _083227_);
  not g_139059_(_083227_, _083228_);
  xor g_139060_(_080216_, _083225_, _083229_);
  not g_139061_(_083229_, _083230_);
  or g_139062_(_081016_, _083229_, _083231_);
  xor g_139063_(_081016_, _083230_, _083232_);
  not g_139064_(_083232_, _083234_);
  or g_139065_(_081015_, _083232_, _083235_);
  xor g_139066_(_081015_, _083234_, _083236_);
  not g_139067_(_083236_, _083237_);
  or g_139068_(_080225_, _083236_, _083238_);
  not g_139069_(_083238_, _083239_);
  or g_139070_(_080222_, _083236_, _083240_);
  xor g_139071_(_080222_, _083237_, _083241_);
  and g_139072_(_080225_, _083241_, _083242_);
  or g_139073_(_083239_, _083242_, _083243_);
  and g_139074_(_080227_, _080229_, _083245_);
  xor g_139075_(_083243_, _083245_, _083246_);
  not g_139076_(_083246_, _083247_);
  or g_139077_(_080232_, _083247_, _083248_);
  xor g_139078_(_080232_, _083246_, _083249_);
  or g_139079_(_077461_, _080228_, _083250_);
  not g_139080_(_083250_, _083251_);
  or g_139081_(_083249_, _083250_, _083252_);
  xor g_139082_(_083249_, _083250_, _083253_);
  xor g_139083_(_083249_, _083251_, _083254_);
  or g_139084_(_081014_, _083254_, _083256_);
  xor g_139085_(_081014_, _083253_, _083257_);
  or g_139086_(_080240_, _083257_, _083258_);
  not g_139087_(_083258_, _083259_);
  and g_139088_(_080237_, _083257_, _083260_);
  and g_139089_(_080240_, _083260_, _083261_);
  or g_139090_(_080237_, _083257_, _083262_);
  not g_139091_(_083262_, _083263_);
  or g_139092_(_083261_, _083263_, _083264_);
  or g_139093_(_083259_, _083264_, _083265_);
  not g_139094_(_083265_, _083267_);
  xor g_139095_(_081013_, _083267_, _083268_);
  not g_139096_(_083268_, _083269_);
  or g_139097_(_081012_, _083268_, _083270_);
  xor g_139098_(_081012_, _083269_, _083271_);
  or g_139099_(_080255_, _083271_, _083272_);
  xor g_139100_(_080254_, _083271_, _083273_);
  not g_139101_(_083273_, _083274_);
  or g_139102_(_080261_, _083273_, _083275_);
  xor g_139103_(_080261_, _083273_, _083276_);
  xor g_139104_(_080261_, _083274_, _083278_);
  or g_139105_(_080260_, _083278_, _083279_);
  not g_139106_(_083279_, _083280_);
  xor g_139107_(_080260_, _083276_, _083281_);
  not g_139108_(_083281_, _083282_);
  and g_139109_(_080267_, _080269_, _083283_);
  xor g_139110_(_083281_, _083283_, _083284_);
  xor g_139111_(_083282_, _083283_, _083285_);
  or g_139112_(_080271_, _083285_, _083286_);
  xor g_139113_(_080271_, _083284_, _083287_);
  not g_139114_(_083287_, _083289_);
  or g_139115_(_080276_, _083287_, _083290_);
  xor g_139116_(_080276_, _083287_, _083291_);
  xor g_139117_(_080276_, _083289_, _083292_);
  or g_139118_(_080279_, _083292_, _083293_);
  xor g_139119_(_080279_, _083291_, _083294_);
  or g_139120_(_080285_, _083294_, _083295_);
  xor g_139121_(_080284_, _083294_, _083296_);
  not g_139122_(_083296_, _083297_);
  or g_139123_(_080289_, _083296_, _083298_);
  xor g_139124_(_080289_, _083297_, _083300_);
  or g_139125_(_080293_, _083300_, _083301_);
  xor g_139126_(_080292_, _083300_, _083302_);
  or g_139127_(_080296_, _083302_, _083303_);
  xor g_139128_(_080296_, _083302_, _083304_);
  xor g_139129_(_080304_, _083304_, _083305_);
  not g_139130_(_083305_, _083306_);
  or g_139131_(_080310_, _083305_, _083307_);
  xor g_139132_(_080310_, _083305_, _083308_);
  xor g_139133_(_080310_, _083306_, _083309_);
  or g_139134_(_080313_, _083309_, _083311_);
  xor g_139135_(_080313_, _083308_, _083312_);
  not g_139136_(_083312_, _083313_);
  and g_139137_(_080315_, _080317_, _083314_);
  xor g_139138_(_083313_, _083314_, _083315_);
  or g_139139_(_081010_, _083315_, _083316_);
  not g_139140_(_083316_, _083317_);
  xor g_139141_(_081010_, _083315_, _083318_);
  not g_139142_(_083318_, _083319_);
  or g_139143_(_081009_, _083319_, _083320_);
  xor g_139144_(_081009_, _083318_, _083322_);
  or g_139145_(_080323_, _083322_, _083323_);
  xor g_139146_(_080324_, _083322_, _083324_);
  and g_139147_(_081008_, _083324_, _083325_);
  or g_139148_(_081008_, _083324_, _083326_);
  not g_139149_(_083326_, _083327_);
  xor g_139150_(_081008_, _083324_, _083328_);
  or g_139151_(_083325_, _083327_, _083329_);
  or g_139152_(_081007_, _083329_, _083330_);
  xor g_139153_(_081007_, _083328_, _083331_);
  not g_139154_(_083331_, _083333_);
  or g_139155_(_081006_, _083331_, _083334_);
  xor g_139156_(_081006_, _083331_, _083335_);
  xor g_139157_(_081006_, _083333_, _083336_);
  and g_139158_(_080331_, _080334_, _083337_);
  xor g_139159_(_083335_, _083337_, _083338_);
  or g_139160_(_080339_, _080342_, _083339_);
  and g_139161_(_080338_, _083339_, _083340_);
  and g_139162_(_083338_, _083340_, _083341_);
  or g_139163_(_083338_, _083340_, _083342_);
  not g_139164_(_083342_, _083344_);
  xor g_139165_(_083338_, _083340_, _083345_);
  or g_139166_(_083341_, _083344_, _083346_);
  or g_139167_(_081005_, _083346_, _083347_);
  xor g_139168_(_081005_, _083345_, _083348_);
  not g_139169_(_083348_, _083349_);
  or g_139170_(_080345_, _083348_, _083350_);
  xor g_139171_(_080345_, _083348_, _083351_);
  xor g_139172_(_080345_, _083349_, _083352_);
  or g_139173_(_080351_, _083352_, _083353_);
  not g_139174_(_083353_, _083355_);
  and g_139175_(_080348_, _083349_, _083356_);
  or g_139176_(_080349_, _083348_, _083357_);
  and g_139177_(_080349_, _083352_, _083358_);
  or g_139178_(_080348_, _083351_, _083359_);
  and g_139179_(_083357_, _083359_, _083360_);
  or g_139180_(_083356_, _083358_, _083361_);
  or g_139181_(_080356_, _083361_, _083362_);
  xor g_139182_(_080356_, _083360_, _083363_);
  and g_139183_(_080351_, _083363_, _083364_);
  or g_139184_(_083355_, _083364_, _083366_);
  or g_139185_(_080365_, _083366_, _083367_);
  xor g_139186_(_080366_, _083366_, _083368_);
  not g_139187_(_083368_, _083369_);
  or g_139188_(_080364_, _083368_, _083370_);
  xor g_139189_(_080364_, _083368_, _083371_);
  xor g_139190_(_080364_, _083369_, _083372_);
  or g_139191_(_080371_, _083372_, _083373_);
  not g_139192_(_083373_, _083374_);
  xor g_139193_(_080371_, _083371_, _083375_);
  or g_139194_(_080373_, _083375_, _083377_);
  xor g_139195_(_080375_, _083375_, _083378_);
  and g_139196_(_080377_, _080381_, _083379_);
  xor g_139197_(_083378_, _083379_, _083380_);
  not g_139198_(_083380_, _083381_);
  or g_139199_(_080384_, _083381_, _083382_);
  xor g_139200_(_080384_, _083380_, _083383_);
  not g_139201_(_083383_, _083384_);
  or g_139202_(_080387_, _083383_, _083385_);
  xor g_139203_(_080387_, _083384_, _083386_);
  or g_139204_(_080390_, _083386_, _083388_);
  not g_139205_(_083388_, _083389_);
  xor g_139206_(_080391_, _083386_, _083390_);
  not g_139207_(_083390_, _083391_);
  and g_139208_(_080398_, _083391_, _083392_);
  not g_139209_(_083392_, _083393_);
  or g_139210_(_080394_, _083390_, _083394_);
  xor g_139211_(_080394_, _083390_, _083395_);
  not g_139212_(_083395_, _083396_);
  or g_139213_(_080402_, _083396_, _083397_);
  xor g_139214_(_080402_, _083395_, _083399_);
  and g_139215_(_080397_, _083399_, _083400_);
  or g_139216_(_083392_, _083400_, _083401_);
  not g_139217_(_083401_, _083402_);
  or g_139218_(_080404_, _083401_, _083403_);
  xor g_139219_(_080404_, _083402_, _083404_);
  or g_139220_(_080406_, _083404_, _083405_);
  xor g_139221_(_080408_, _083404_, _083406_);
  and g_139222_(_080410_, _080413_, _083407_);
  not g_139223_(_083407_, _083408_);
  xor g_139224_(_083406_, _083408_, _083410_);
  or g_139225_(_081004_, _083410_, _083411_);
  not g_139226_(_083411_, _083412_);
  xor g_139227_(_081004_, _083410_, _083413_);
  not g_139228_(_083413_, _083414_);
  and g_139229_(_081003_, _083413_, _083415_);
  or g_139230_(_081002_, _083414_, _083416_);
  xor g_139231_(_081002_, _083413_, _083417_);
  or g_139232_(_080419_, _083417_, _083418_);
  xor g_139233_(_080417_, _083417_, _083419_);
  not g_139234_(_083419_, _083421_);
  or g_139235_(_080421_, _083419_, _083422_);
  xor g_139236_(_080421_, _083419_, _083423_);
  xor g_139237_(_080421_, _083421_, _083424_);
  or g_139238_(_080424_, _083424_, _083425_);
  xor g_139239_(_080424_, _083423_, _083426_);
  or g_139240_(_081001_, _083426_, _083427_);
  xor g_139241_(_081001_, _083426_, _083428_);
  not g_139242_(_083428_, _083429_);
  or g_139243_(_077650_, _080426_, _083430_);
  or g_139244_(_083429_, _083430_, _083432_);
  not g_139245_(_083432_, _083433_);
  xor g_139246_(_083428_, _083430_, _083434_);
  not g_139247_(_083434_, _083435_);
  or g_139248_(_080999_, _083434_, _083436_);
  xor g_139249_(_080999_, _083434_, _083437_);
  xor g_139250_(_080999_, _083435_, _083438_);
  or g_139251_(_080998_, _083438_, _083439_);
  xor g_139252_(_080998_, _083437_, _083440_);
  not g_139253_(_083440_, _083441_);
  and g_139254_(_080431_, _080435_, _083443_);
  xor g_139255_(_083441_, _083443_, _083444_);
  xor g_139256_(_083440_, _083443_, _083445_);
  or g_139257_(_080438_, _083444_, _083446_);
  xor g_139258_(_080438_, _083445_, _083447_);
  not g_139259_(_083447_, _083448_);
  and g_139260_(_080442_, _080446_, _083449_);
  xor g_139261_(_083448_, _083449_, _083450_);
  or g_139262_(_080449_, _083450_, _083451_);
  xor g_139263_(_080450_, _083450_, _083452_);
  or g_139264_(_080453_, _083452_, _083454_);
  xor g_139265_(_080453_, _083452_, _083455_);
  not g_139266_(_083455_, _083456_);
  or g_139267_(_080457_, _083456_, _083457_);
  xor g_139268_(_080457_, _083455_, _083458_);
  not g_139269_(_083458_, _083459_);
  or g_139270_(_080461_, _083458_, _083460_);
  xor g_139271_(_080461_, _083459_, _083461_);
  or g_139272_(_080996_, _083461_, _083462_);
  xor g_139273_(_080997_, _083461_, _083463_);
  not g_139274_(_083463_, _083465_);
  or g_139275_(_080995_, _083463_, _083466_);
  xor g_139276_(_080995_, _083463_, _083467_);
  xor g_139277_(_080995_, _083465_, _083468_);
  and g_139278_(_080465_, _083467_, _083469_);
  or g_139279_(_080464_, _083468_, _083470_);
  xor g_139280_(_080464_, _083467_, _083471_);
  and g_139281_(_080469_, _080474_, _083472_);
  xor g_139282_(_083471_, _083472_, _083473_);
  not g_139283_(_083473_, _083474_);
  or g_139284_(_080477_, _083474_, _083476_);
  not g_139285_(_083476_, _083477_);
  xor g_139286_(_080477_, _083473_, _083478_);
  not g_139287_(_083478_, _083479_);
  or g_139288_(_080479_, _083478_, _083480_);
  xor g_139289_(_080479_, _083479_, _083481_);
  not g_139290_(_083481_, _083482_);
  and g_139291_(_080482_, _080485_, _083483_);
  xor g_139292_(_083481_, _083483_, _083484_);
  xor g_139293_(_083482_, _083483_, _083485_);
  or g_139294_(_080994_, _083485_, _083487_);
  xor g_139295_(_080994_, _083484_, _083488_);
  not g_139296_(_083488_, _083489_);
  or g_139297_(_080993_, _083488_, _083490_);
  xor g_139298_(_080993_, _083489_, _083491_);
  not g_139299_(_083491_, _083492_);
  and g_139300_(_080488_, _080491_, _083493_);
  xor g_139301_(_083491_, _083493_, _083494_);
  xor g_139302_(_083492_, _083493_, _083495_);
  or g_139303_(_080493_, _083495_, _083496_);
  xor g_139304_(_080493_, _083494_, _083498_);
  or g_139305_(_080498_, _083498_, _083499_);
  xor g_139306_(_080497_, _083498_, _083500_);
  or g_139307_(_080501_, _083500_, _083501_);
  xor g_139308_(_080501_, _083500_, _083502_);
  not g_139309_(_083502_, _083503_);
  or g_139310_(_080505_, _083503_, _083504_);
  xor g_139311_(_080505_, _083502_, _083505_);
  not g_139312_(_083505_, _083506_);
  or g_139313_(_080509_, _083505_, _083507_);
  xor g_139314_(_080509_, _083506_, _083509_);
  not g_139315_(_083509_, _083510_);
  and g_139316_(_080512_, _080515_, _083511_);
  xor g_139317_(_083509_, _083511_, _083512_);
  xor g_139318_(_083510_, _083511_, _083513_);
  or g_139319_(_077758_, _080521_, _083514_);
  and g_139320_(_080519_, _083514_, _083515_);
  not g_139321_(_083515_, _083516_);
  and g_139322_(_083512_, _083516_, _083517_);
  xor g_139323_(_083513_, _083515_, _083518_);
  xor g_139324_(_083512_, _083515_, _083520_);
  or g_139325_(_080992_, _083520_, _083521_);
  xor g_139326_(_080992_, _083518_, _083522_);
  or g_139327_(_080530_, _083522_, _083523_);
  xor g_139328_(_080529_, _083522_, _083524_);
  or g_139329_(_080526_, _083524_, _083525_);
  xor g_139330_(_080526_, _083524_, _083526_);
  xor g_139331_(_080527_, _083524_, _083527_);
  and g_139332_(_080533_, _080535_, _083528_);
  or g_139333_(_083527_, _083528_, _083529_);
  not g_139334_(_083529_, _083531_);
  xor g_139335_(_083527_, _083528_, _083532_);
  xor g_139336_(_083526_, _083528_, _083533_);
  or g_139337_(_080537_, _083533_, _083534_);
  not g_139338_(_083534_, _083535_);
  or g_139339_(_080541_, _083533_, _083536_);
  xor g_139340_(_080541_, _083532_, _083537_);
  and g_139341_(_080537_, _083537_, _083538_);
  or g_139342_(_083535_, _083538_, _083539_);
  or g_139343_(_080545_, _083539_, _083540_);
  xor g_139344_(_080544_, _083539_, _083542_);
  or g_139345_(_077795_, _080546_, _083543_);
  not g_139346_(_083543_, _083544_);
  or g_139347_(_083542_, _083543_, _083545_);
  xor g_139348_(_083542_, _083544_, _083546_);
  or g_139349_(_080990_, _083546_, _083547_);
  xor g_139350_(_080991_, _083546_, _083548_);
  not g_139351_(_083548_, _083549_);
  or g_139352_(_080988_, _083548_, _083550_);
  xor g_139353_(_080988_, _083549_, _083551_);
  or g_139354_(_077807_, _080552_, _083553_);
  and g_139355_(_080551_, _083553_, _083554_);
  or g_139356_(_083551_, _083554_, _083555_);
  xor g_139357_(_083551_, _083554_, _083556_);
  not g_139358_(_083556_, _083557_);
  or g_139359_(_080987_, _083557_, _083558_);
  not g_139360_(_083558_, _083559_);
  xor g_139361_(_080987_, _083556_, _083560_);
  or g_139362_(_080557_, _083560_, _083561_);
  not g_139363_(_083561_, _083562_);
  or g_139364_(_080566_, _083560_, _083564_);
  xor g_139365_(_080565_, _083560_, _083565_);
  and g_139366_(_080557_, _083565_, _083566_);
  or g_139367_(_083562_, _083566_, _083567_);
  or g_139368_(_080563_, _083567_, _083568_);
  xor g_139369_(_080563_, _083567_, _083569_);
  xor g_139370_(_080564_, _083567_, _083570_);
  or g_139371_(_077821_, _080568_, _083571_);
  or g_139372_(_083570_, _083571_, _083572_);
  xor g_139373_(_083569_, _083571_, _083573_);
  or g_139374_(_077822_, _080568_, _083575_);
  not g_139375_(_083575_, _083576_);
  or g_139376_(_083573_, _083575_, _083577_);
  xor g_139377_(_083573_, _083576_, _083578_);
  xor g_139378_(_080573_, _083578_, _083579_);
  not g_139379_(_083579_, _083580_);
  or g_139380_(_080579_, _083579_, _083581_);
  not g_139381_(_083581_, _083582_);
  and g_139382_(_080576_, _083579_, _083583_);
  and g_139383_(_080579_, _083583_, _083584_);
  and g_139384_(_080577_, _083580_, _083586_);
  not g_139385_(_083586_, _083587_);
  or g_139386_(_083584_, _083586_, _083588_);
  or g_139387_(_083582_, _083588_, _083589_);
  not g_139388_(_083589_, _083590_);
  or g_139389_(_080582_, _083589_, _083591_);
  xor g_139390_(_080582_, _083590_, _083592_);
  or g_139391_(_080589_, _083592_, _083593_);
  xor g_139392_(_080588_, _083592_, _083594_);
  or g_139393_(_080592_, _083594_, _083595_);
  xor g_139394_(_080593_, _083594_, _083597_);
  or g_139395_(_080601_, _083597_, _083598_);
  not g_139396_(_083598_, _083599_);
  xor g_139397_(_080602_, _083597_, _083600_);
  and g_139398_(_080606_, _083600_, _083601_);
  or g_139399_(_080606_, _083597_, _083602_);
  not g_139400_(_083602_, _083603_);
  or g_139401_(_083601_, _083603_, _083604_);
  not g_139402_(_083604_, _083605_);
  and g_139403_(_080609_, _080612_, _083606_);
  xor g_139404_(_083605_, _083606_, _083608_);
  or g_139405_(_080615_, _083608_, _083609_);
  xor g_139406_(_080615_, _083608_, _083610_);
  xor g_139407_(_080617_, _083608_, _083611_);
  and g_139408_(_080620_, _080622_, _083612_);
  xor g_139409_(_083610_, _083612_, _083613_);
  not g_139410_(_083613_, _083614_);
  or g_139411_(_080626_, _083613_, _083615_);
  xor g_139412_(_080626_, _083614_, _083616_);
  not g_139413_(_083616_, _083617_);
  and g_139414_(_080631_, _080633_, _083619_);
  xor g_139415_(_083617_, _083619_, _083620_);
  or g_139416_(_080635_, _083620_, _083621_);
  xor g_139417_(_080635_, _083620_, _083622_);
  not g_139418_(_083622_, _083623_);
  and g_139419_(_080637_, _080642_, _083624_);
  xor g_139420_(_083622_, _083624_, _083625_);
  not g_139421_(_083625_, _083626_);
  or g_139422_(_080645_, _083625_, _083627_);
  xor g_139423_(_080645_, _083625_, _083628_);
  xor g_139424_(_080645_, _083626_, _083630_);
  and g_139425_(_080647_, _080651_, _083631_);
  xor g_139426_(_083628_, _083631_, _083632_);
  or g_139427_(_080657_, _083632_, _083633_);
  not g_139428_(_083633_, _083634_);
  and g_139429_(_080655_, _083632_, _083635_);
  and g_139430_(_080657_, _083635_, _083636_);
  or g_139431_(_080655_, _083632_, _083637_);
  not g_139432_(_083637_, _083638_);
  or g_139433_(_083636_, _083638_, _083639_);
  or g_139434_(_083634_, _083639_, _083641_);
  not g_139435_(_083641_, _083642_);
  or g_139436_(_080659_, _083641_, _083643_);
  xor g_139437_(_080659_, _083641_, _083644_);
  xor g_139438_(_080659_, _083642_, _083645_);
  or g_139439_(_080667_, _083645_, _083646_);
  xor g_139440_(_080667_, _083644_, _083647_);
  or g_139441_(_080669_, _083647_, _083648_);
  xor g_139442_(_080670_, _083647_, _083649_);
  or g_139443_(_080985_, _083649_, _083650_);
  not g_139444_(_083650_, _083652_);
  xor g_139445_(_080986_, _083649_, _083653_);
  not g_139446_(_083653_, _083654_);
  or g_139447_(_080984_, _083653_, _083655_);
  xor g_139448_(_080984_, _083653_, _083656_);
  xor g_139449_(_080984_, _083654_, _083657_);
  or g_139450_(_080983_, _083657_, _083658_);
  not g_139451_(_083658_, _083659_);
  xor g_139452_(_080983_, _083656_, _083660_);
  and g_139453_(_080677_, _080680_, _083661_);
  or g_139454_(_083660_, _083661_, _083663_);
  xor g_139455_(_083660_, _083661_, _083664_);
  not g_139456_(_083664_, _083665_);
  or g_139457_(_080684_, _083665_, _083666_);
  not g_139458_(_083666_, _083667_);
  xor g_139459_(_080684_, _083664_, _083668_);
  not g_139460_(_083668_, _083669_);
  or g_139461_(_080686_, _083668_, _083670_);
  xor g_139462_(_080686_, _083669_, _083671_);
  or g_139463_(_080689_, _083671_, _083672_);
  not g_139464_(_083672_, _083674_);
  and g_139465_(_080689_, _083671_, _083675_);
  xor g_139466_(_080689_, _083671_, _083676_);
  or g_139467_(_083674_, _083675_, _083677_);
  or g_139468_(_080982_, _083677_, _083678_);
  not g_139469_(_083678_, _083679_);
  xor g_139470_(_080982_, _083676_, _083680_);
  not g_139471_(_083680_, _083681_);
  or g_139472_(_080981_, _083680_, _083682_);
  xor g_139473_(_080981_, _083680_, _083683_);
  xor g_139474_(_080981_, _083681_, _083685_);
  or g_139475_(_080695_, _083685_, _083686_);
  not g_139476_(_083686_, _083687_);
  xor g_139477_(_080695_, _083683_, _083688_);
  or g_139478_(_080697_, _083688_, _083689_);
  not g_139479_(_083689_, _083690_);
  and g_139480_(_080697_, _083688_, _083691_);
  xor g_139481_(_080697_, _083688_, _083692_);
  or g_139482_(_083690_, _083691_, _083693_);
  or g_139483_(_080701_, _083693_, _083694_);
  xor g_139484_(_080701_, _083692_, _083696_);
  or g_139485_(_080706_, _083696_, _083697_);
  xor g_139486_(_080707_, _083696_, _083698_);
  or g_139487_(_080709_, _083698_, _083699_);
  not g_139488_(_083699_, _083700_);
  xor g_139489_(_080710_, _083698_, _083701_);
  not g_139490_(_083701_, _083702_);
  or g_139491_(_080712_, _083701_, _083703_);
  xor g_139492_(_080712_, _083701_, _083704_);
  xor g_139493_(_080712_, _083702_, _083705_);
  and g_139494_(_080980_, _083704_, _083707_);
  or g_139495_(_080979_, _083705_, _083708_);
  or g_139496_(_080714_, _083705_, _083709_);
  xor g_139497_(_080714_, _083704_, _083710_);
  and g_139498_(_080979_, _083710_, _083711_);
  or g_139499_(_083707_, _083711_, _083712_);
  or g_139500_(_080977_, _083712_, _083713_);
  xor g_139501_(_080976_, _083712_, _083714_);
  or g_139502_(_080722_, _083714_, _083715_);
  xor g_139503_(_080722_, _083714_, _083716_);
  and g_139504_(_080725_, _083716_, _083718_);
  not g_139505_(_083718_, _083719_);
  xor g_139506_(_080724_, _083716_, _083720_);
  or g_139507_(_080730_, _083720_, _083721_);
  not g_139508_(_083721_, _083722_);
  xor g_139509_(_080729_, _083720_, _083723_);
  or g_139510_(_080734_, _083723_, _083724_);
  xor g_139511_(_080735_, _083723_, _083725_);
  not g_139512_(_083725_, _083726_);
  and g_139513_(_080739_, _080741_, _083727_);
  xor g_139514_(_083725_, _083727_, _083729_);
  xor g_139515_(_083726_, _083727_, _083730_);
  or g_139516_(_080745_, _083730_, _083731_);
  xor g_139517_(_080745_, _083729_, _083732_);
  and g_139518_(_080747_, _080750_, _083733_);
  not g_139519_(_083733_, _083734_);
  xor g_139520_(_083732_, _083733_, _083735_);
  xor g_139521_(_083732_, _083734_, _083736_);
  and g_139522_(_080752_, _083736_, _083737_);
  or g_139523_(_080753_, _083735_, _083738_);
  and g_139524_(_080756_, _083737_, _083740_);
  or g_139525_(_080757_, _083738_, _083741_);
  or g_139526_(_080756_, _083736_, _083742_);
  not g_139527_(_083742_, _083743_);
  or g_139528_(_080752_, _083736_, _083744_);
  not g_139529_(_083744_, _083745_);
  and g_139530_(_083742_, _083744_, _083746_);
  not g_139531_(_083746_, _083747_);
  and g_139532_(_083741_, _083746_, _083748_);
  or g_139533_(_083740_, _083747_, _083749_);
  or g_139534_(_080975_, _083749_, _083751_);
  xor g_139535_(_080975_, _083748_, _083752_);
  or g_139536_(_080974_, _083752_, _083753_);
  xor g_139537_(_080973_, _083752_, _083754_);
  or g_139538_(_080972_, _083754_, _083755_);
  xor g_139539_(_080971_, _083754_, _083756_);
  or g_139540_(_080970_, _083756_, _083757_);
  xor g_139541_(_080969_, _083756_, _083758_);
  or g_139542_(_080764_, _083758_, _083759_);
  xor g_139543_(_080765_, _083758_, _083760_);
  not g_139544_(_083760_, _083762_);
  and g_139545_(_080768_, _080772_, _083763_);
  xor g_139546_(_083760_, _083763_, _083764_);
  xor g_139547_(_083762_, _083763_, _083765_);
  or g_139548_(_080776_, _083765_, _083766_);
  not g_139549_(_083766_, _083767_);
  xor g_139550_(_080776_, _083764_, _083768_);
  or g_139551_(_080780_, _083768_, _083769_);
  xor g_139552_(_080779_, _083768_, _083770_);
  or g_139553_(_080783_, _083770_, _083771_);
  xor g_139554_(_080784_, _083770_, _083773_);
  and g_139555_(_080786_, _080788_, _083774_);
  or g_139556_(_083773_, _083774_, _083775_);
  xor g_139557_(_083773_, _083774_, _083776_);
  not g_139558_(_083776_, _083777_);
  and g_139559_(_080968_, _083776_, _083778_);
  or g_139560_(_080966_, _083777_, _083779_);
  xor g_139561_(_080966_, _083776_, _083780_);
  not g_139562_(_083780_, _083781_);
  or g_139563_(_080798_, _083780_, _083782_);
  xor g_139564_(_080798_, _083780_, _083784_);
  xor g_139565_(_080798_, _083781_, _083785_);
  and g_139566_(_080801_, _083784_, _083786_);
  or g_139567_(_080802_, _083785_, _083787_);
  xor g_139568_(_080802_, _083784_, _083788_);
  or g_139569_(_080805_, _083788_, _083789_);
  xor g_139570_(_080806_, _083788_, _083790_);
  or g_139571_(_078016_, _080804_, _083791_);
  and g_139572_(_083790_, _083791_, _083792_);
  or g_139573_(_083790_, _083791_, _083793_);
  not g_139574_(_083793_, _083795_);
  or g_139575_(_083792_, _083795_, _083796_);
  and g_139576_(_080810_, _080813_, _083797_);
  xor g_139577_(_083796_, _083797_, _083798_);
  not g_139578_(_083798_, _083799_);
  and g_139579_(_080817_, _083798_, _083800_);
  or g_139580_(_080816_, _083799_, _083801_);
  xor g_139581_(_080816_, _083798_, _083802_);
  and g_139582_(_080821_, _080827_, _083803_);
  not g_139583_(_083803_, _083804_);
  xor g_139584_(_083802_, _083804_, _083806_);
  or g_139585_(_080830_, _083806_, _083807_);
  xor g_139586_(_080830_, _083806_, _083808_);
  xor g_139587_(_080831_, _083806_, _083809_);
  and g_139588_(_080834_, _080839_, _083810_);
  not g_139589_(_083810_, _083811_);
  and g_139590_(_083808_, _083811_, _083812_);
  xor g_139591_(_083809_, _083810_, _083813_);
  and g_139592_(_080844_, _083813_, _083814_);
  xor g_139593_(_080843_, _083813_, _083815_);
  or g_139594_(_080965_, _083815_, _083817_);
  not g_139595_(_083817_, _083818_);
  and g_139596_(_080965_, _083815_, _083819_);
  xor g_139597_(_080965_, _083815_, _083820_);
  or g_139598_(_083818_, _083819_, _083821_);
  or g_139599_(_080964_, _083821_, _083822_);
  xor g_139600_(_080964_, _083820_, _083823_);
  or g_139601_(_080961_, _083823_, _083824_);
  not g_139602_(_083824_, _083825_);
  xor g_139603_(_080961_, _083823_, _083826_);
  xor g_139604_(_080962_, _083823_, _083828_);
  and g_139605_(_080850_, _083828_, _083829_);
  and g_139606_(_080959_, _083829_, _083830_);
  and g_139607_(_080851_, _083826_, _083831_);
  not g_139608_(_083831_, _083832_);
  and g_139609_(_080960_, _083826_, _083833_);
  or g_139610_(_083831_, _083833_, _083834_);
  or g_139611_(_083830_, _083834_, _083835_);
  not g_139612_(_083835_, _083836_);
  and g_139613_(_080957_, _083836_, _083837_);
  or g_139614_(_080958_, _083835_, _083839_);
  xor g_139615_(_080957_, _083835_, _083840_);
  or g_139616_(_080954_, _083840_, _083841_);
  not g_139617_(_083841_, _083842_);
  xor g_139618_(_080955_, _083840_, _083843_);
  not g_139619_(_083843_, _083844_);
  or g_139620_(_080953_, _083843_, _083845_);
  xor g_139621_(_080953_, _083844_, _083846_);
  and g_139622_(_080860_, _080863_, _083847_);
  not g_139623_(_083847_, _083848_);
  xor g_139624_(_083846_, _083848_, _083850_);
  not g_139625_(_083850_, _083851_);
  and g_139626_(_080872_, _083851_, _083852_);
  or g_139627_(_080871_, _083850_, _083853_);
  xor g_139628_(_080871_, _083850_, _083854_);
  and g_139629_(_080870_, _083854_, _083855_);
  not g_139630_(_083855_, _083856_);
  xor g_139631_(_080868_, _083854_, _083857_);
  and g_139632_(_080877_, _083857_, _083858_);
  and g_139633_(_080882_, _083858_, _083859_);
  or g_139634_(_080877_, _083857_, _083861_);
  not g_139635_(_083861_, _083862_);
  or g_139636_(_080882_, _083857_, _083863_);
  and g_139637_(_083861_, _083863_, _083864_);
  not g_139638_(_083864_, _083865_);
  or g_139639_(_083859_, _083865_, _083866_);
  not g_139640_(_083866_, _083867_);
  xor g_139641_(_080952_, _083867_, _083868_);
  or g_139642_(_080949_, _083868_, _083869_);
  xor g_139643_(_080950_, _083868_, _083870_);
  not g_139644_(_083870_, _083872_);
  or g_139645_(_080893_, _083870_, _083873_);
  not g_139646_(_083873_, _083874_);
  xor g_139647_(_080893_, _083872_, _083875_);
  or g_139648_(_080947_, _083875_, _083876_);
  xor g_139649_(_080948_, _083875_, _083877_);
  not g_139650_(_083877_, _083878_);
  or g_139651_(_078100_, _080895_, _083879_);
  and g_139652_(_080898_, _083879_, _083880_);
  xor g_139653_(_083878_, _083880_, _083881_);
  not g_139654_(_083881_, _083883_);
  or g_139655_(_080946_, _083881_, _083884_);
  xor g_139656_(_080946_, _083883_, _083885_);
  not g_139657_(_083885_, _083886_);
  or g_139658_(_080944_, _083885_, _083887_);
  xor g_139659_(_080944_, _083885_, _083888_);
  xor g_139660_(_080944_, _083886_, _083889_);
  or g_139661_(_078112_, _080899_, _083890_);
  not g_139662_(_083890_, _083891_);
  and g_139663_(_080904_, _083890_, _083892_);
  xor g_139664_(_083888_, _083892_, _083894_);
  xor g_139665_(_083889_, _083892_, _083895_);
  and g_139666_(_080909_, _083895_, _083896_);
  or g_139667_(_080908_, _083894_, _083897_);
  xor g_139668_(_080908_, _083894_, _083898_);
  xor g_139669_(_080909_, _083894_, _083899_);
  and g_139670_(_080912_, _083899_, _083900_);
  and g_139671_(_080918_, _083900_, _083901_);
  and g_139672_(_080917_, _083898_, _083902_);
  not g_139673_(_083902_, _083903_);
  and g_139674_(_080914_, _083898_, _083905_);
  or g_139675_(_080912_, _083899_, _083906_);
  or g_139676_(_083902_, _083905_, _083907_);
  or g_139677_(_083901_, _083907_, _083908_);
  or g_139678_(_080942_, _083908_, _083909_);
  xor g_139679_(_080942_, _083908_, _083910_);
  not g_139680_(_083910_, _083911_);
  or g_139681_(_080941_, _083911_, _083912_);
  xor g_139682_(_080941_, _083910_, _083913_);
  not g_139683_(_083913_, _083914_);
  and g_139684_(_080925_, _080928_, _083916_);
  xor g_139685_(_083914_, _083916_, _083917_);
  xor g_139686_(_083913_, _083916_, _083918_);
  or g_139687_(_080931_, _083917_, _083919_);
  xor g_139688_(_080931_, _083918_, _083920_);
  and g_139689_(_080933_, _083920_, _083921_);
  not g_139690_(_083921_, _083922_);
  or g_139691_(_078139_, _080929_, _083923_);
  or g_139692_(_083920_, _083923_, _083924_);
  and g_139693_(_083922_, _083924_, _083925_);
  not g_139694_(_083925_, _083927_);
  and g_139695_(_080938_, _083925_, _083928_);
  or g_139696_(_080937_, _083927_, _083929_);
  xor g_139697_(_080937_, _083925_, _083930_);
  or g_139698_(_080940_, _083930_, _083931_);
  xor g_139699_(_080940_, _083930_, out[963]);
  or g_139700_(_080928_, _083913_, _083932_);
  or g_139701_(_080925_, _083913_, _083933_);
  or g_139702_(_080904_, _083889_, _083934_);
  not g_139703_(_083934_, _083935_);
  and g_139704_(_083888_, _083891_, _083937_);
  or g_139705_(_083889_, _083890_, _083938_);
  or g_139706_(_080898_, _083877_, _083939_);
  or g_139707_(_083877_, _083879_, _083940_);
  or g_139708_(_080951_, _083866_, _083941_);
  not g_139709_(_083941_, _083942_);
  or g_139710_(_080860_, _083846_, _083943_);
  or g_139711_(_080827_, _083802_, _083944_);
  not g_139712_(_083944_, _083945_);
  or g_139713_(_080813_, _083796_, _083946_);
  not g_139714_(_083946_, _083948_);
  or g_139715_(_078018_, _080808_, _083949_);
  or g_139716_(_083796_, _083949_, _083950_);
  and g_139717_(_083789_, _083793_, _083951_);
  or g_139718_(_080772_, _083760_, _083952_);
  or g_139719_(_080768_, _083760_, _083953_);
  not g_139720_(_083953_, _083954_);
  or g_139721_(_080750_, _083732_, _083955_);
  or g_139722_(_080741_, _083725_, _083956_);
  and g_139723_(_083694_, _083697_, _083957_);
  or g_139724_(_080651_, _083630_, _083959_);
  or g_139725_(_080642_, _083623_, _083960_);
  not g_139726_(_083960_, _083961_);
  or g_139727_(_080633_, _083616_, _083962_);
  or g_139728_(_080622_, _083611_, _083963_);
  or g_139729_(_080620_, _083611_, _083964_);
  or g_139730_(_080612_, _083604_, _083965_);
  not g_139731_(_083965_, _083966_);
  and g_139732_(_083593_, _083595_, _083967_);
  or g_139733_(_080570_, _083578_, _083968_);
  or g_139734_(_077828_, _083968_, _083970_);
  not g_139735_(_083970_, _083971_);
  or g_139736_(_077826_, _083968_, _083972_);
  or g_139737_(_080515_, _083509_, _083973_);
  or g_139738_(_080512_, _083509_, _083974_);
  or g_139739_(_080491_, _083491_, _083975_);
  or g_139740_(_080485_, _083481_, _083976_);
  and g_139741_(_083487_, _083976_, _083977_);
  or g_139742_(_080474_, _083471_, _083978_);
  or g_139743_(_080469_, _083471_, _083979_);
  not g_139744_(_083979_, _083981_);
  and g_139745_(_083462_, _083466_, _083982_);
  not g_139746_(_083982_, _083983_);
  or g_139747_(_080442_, _083447_, _083984_);
  not g_139748_(_083984_, _083985_);
  or g_139749_(_080435_, _083440_, _083986_);
  and g_139750_(_083446_, _083986_, _083987_);
  and g_139751_(_083425_, _083427_, _083988_);
  not g_139752_(_083988_, _083989_);
  and g_139753_(_083388_, _083394_, _083990_);
  or g_139754_(_080381_, _083378_, _083992_);
  or g_139755_(_080377_, _083375_, _083993_);
  and g_139756_(_083347_, _083350_, _083994_);
  or g_139757_(_080334_, _083336_, _083995_);
  or g_139758_(_080317_, _083312_, _083996_);
  or g_139759_(_080315_, _083312_, _083997_);
  or g_139760_(_080301_, _083302_, _083998_);
  or g_139761_(_080303_, _083302_, _083999_);
  or g_139762_(_080269_, _083281_, _084000_);
  or g_139763_(_080267_, _083281_, _084001_);
  not g_139764_(_084001_, _084003_);
  or g_139765_(_080245_, _083265_, _084004_);
  or g_139766_(_080243_, _083265_, _084005_);
  and g_139767_(_083258_, _084005_, _084006_);
  and g_139768_(_083256_, _083262_, _084007_);
  or g_139769_(_080229_, _083243_, _084008_);
  or g_139770_(_080227_, _083241_, _084009_);
  or g_139771_(_080162_, _083179_, _084010_);
  or g_139772_(_083179_, _083180_, _084011_);
  or g_139773_(_080140_, _083142_, _084012_);
  or g_139774_(_080134_, _083135_, _084014_);
  or g_139775_(_080131_, _083135_, _084015_);
  or g_139776_(_080124_, _083127_, _084016_);
  or g_139777_(_080103_, _083099_, _084017_);
  and g_139778_(_080100_, _083098_, _084018_);
  and g_139779_(_080087_, _083093_, _084019_);
  or g_139780_(_080086_, _083094_, _084020_);
  or g_139781_(_077302_, _084020_, _084021_);
  and g_139782_(_077296_, _084019_, _084022_);
  or g_139783_(_077294_, _084020_, _084023_);
  or g_139784_(_080071_, _083080_, _084025_);
  or g_139785_(_077282_, _084025_, _084026_);
  not g_139786_(_084026_, _084027_);
  or g_139787_(_080068_, _083078_, _084028_);
  not g_139788_(_084028_, _084029_);
  or g_139789_(_081035_, _083078_, _084030_);
  or g_139790_(_083074_, _083076_, _084031_);
  not g_139791_(_084031_, _084032_);
  or g_139792_(_080059_, _083074_, _084033_);
  not g_139793_(_084033_, _084034_);
  and g_139794_(_083073_, _084033_, _084036_);
  or g_139795_(_080053_, _083067_, _084037_);
  not g_139796_(_084037_, _084038_);
  or g_139797_(_080051_, _083063_, _084039_);
  or g_139798_(_080048_, _083063_, _084040_);
  not g_139799_(_084040_, _084041_);
  or g_139800_(_080037_, _083045_, _084042_);
  not g_139801_(_084042_, _084043_);
  or g_139802_(_080025_, _083040_, _084044_);
  not g_139803_(_084044_, _084045_);
  or g_139804_(_080020_, _083040_, _084047_);
  not g_139805_(_084047_, _084048_);
  and g_139806_(_082986_, _082992_, _084049_);
  or g_139807_(_079955_, _082957_, _084050_);
  not g_139808_(_084050_, _084051_);
  or g_139809_(_079951_, _082957_, _084052_);
  and g_139810_(_079931_, _082935_, _084053_);
  or g_139811_(_079930_, _082937_, _084054_);
  or g_139812_(_077140_, _084054_, _084055_);
  not g_139813_(_084055_, _084056_);
  and g_139814_(_077133_, _084053_, _084058_);
  or g_139815_(_077132_, _084054_, _084059_);
  or g_139816_(_081050_, _082928_, _084060_);
  not g_139817_(_084060_, _084061_);
  or g_139818_(_079919_, _082920_, _084062_);
  not g_139819_(_084062_, _084063_);
  or g_139820_(_082912_, _082915_, _084064_);
  not g_139821_(_084064_, _084065_);
  or g_139822_(_079909_, _082912_, _084066_);
  or g_139823_(_079886_, _082893_, _084067_);
  not g_139824_(_084067_, _084069_);
  or g_139825_(_079884_, _082893_, _084070_);
  not g_139826_(_084070_, _084071_);
  or g_139827_(_082858_, _082860_, _084072_);
  or g_139828_(_082858_, _082861_, _084073_);
  and g_139829_(_082818_, _082823_, _084074_);
  or g_139830_(_082819_, _082822_, _084075_);
  or g_139831_(_082813_, _082816_, _084076_);
  and g_139832_(_079837_, _082814_, _084077_);
  or g_139833_(_079836_, _082813_, _084078_);
  or g_139834_(_081068_, _082811_, _084080_);
  not g_139835_(_084080_, _084081_);
  or g_139836_(_079822_, _082802_, _084082_);
  and g_139837_(_082785_, _082787_, _084083_);
  and g_139838_(_079805_, _082785_, _084084_);
  not g_139839_(_084084_, _084085_);
  or g_139840_(_079777_, _082757_, _084086_);
  or g_139841_(_079775_, _082752_, _084087_);
  or g_139842_(_079753_, _082731_, _084088_);
  or g_139843_(_079729_, _082697_, _084089_);
  not g_139844_(_084089_, _084091_);
  or g_139845_(_079727_, _082697_, _084092_);
  and g_139846_(_079685_, _082645_, _084093_);
  or g_139847_(_079684_, _082646_, _084094_);
  or g_139848_(_076860_, _084094_, _084095_);
  and g_139849_(_079662_, _082627_, _084096_);
  not g_139850_(_084096_, _084097_);
  or g_139851_(_079658_, _082629_, _084098_);
  and g_139852_(_082625_, _084098_, _084099_);
  or g_139853_(_079645_, _082603_, _084100_);
  and g_139854_(_082607_, _084100_, _084102_);
  not g_139855_(_084102_, _084103_);
  or g_139856_(_079635_, _082594_, _084104_);
  or g_139857_(_082594_, _082596_, _084105_);
  or g_139858_(_079630_, _082588_, _084106_);
  or g_139859_(_079628_, _082588_, _084107_);
  or g_139860_(_079621_, _082576_, _084108_);
  or g_139861_(_079619_, _082576_, _084109_);
  not g_139862_(_084109_, _084110_);
  or g_139863_(_079601_, _082549_, _084111_);
  not g_139864_(_084111_, _084113_);
  and g_139865_(_079584_, _082537_, _084114_);
  not g_139866_(_084114_, _084115_);
  or g_139867_(_079576_, _082538_, _084116_);
  not g_139868_(_084116_, _084117_);
  or g_139869_(_082487_, _082488_, _084118_);
  or g_139870_(_079532_, _082487_, _084119_);
  not g_139871_(_084119_, _084120_);
  or g_139872_(_079490_, _082437_, _084121_);
  not g_139873_(_084121_, _084122_);
  or g_139874_(_081122_, _082437_, _084124_);
  or g_139875_(_082433_, _082435_, _084125_);
  or g_139876_(_079485_, _082433_, _084126_);
  and g_139877_(_082432_, _084126_, _084127_);
  not g_139878_(_084127_, _084128_);
  or g_139879_(_081126_, _082411_, _084129_);
  not g_139880_(_084129_, _084130_);
  or g_139881_(_079454_, _082411_, _084131_);
  not g_139882_(_084131_, _084132_);
  or g_139883_(_079459_, _082406_, _084133_);
  not g_139884_(_084133_, _084135_);
  and g_139885_(_079432_, _082381_, _084136_);
  or g_139886_(_079433_, _082380_, _084137_);
  or g_139887_(_079429_, _082380_, _084138_);
  or g_139888_(_079413_, _082360_, _084139_);
  or g_139889_(_079379_, _082319_, _084140_);
  and g_139890_(_079375_, _082317_, _084141_);
  not g_139891_(_084141_, _084142_);
  or g_139892_(_079371_, _082316_, _084143_);
  or g_139893_(_079363_, _082307_, _084144_);
  or g_139894_(_079315_, _082268_, _084146_);
  or g_139895_(_082261_, _082262_, _084147_);
  not g_139896_(_084147_, _084148_);
  or g_139897_(_079309_, _082261_, _084149_);
  and g_139898_(_082240_, _082242_, _084150_);
  not g_139899_(_084150_, _084151_);
  or g_139900_(_079282_, _082239_, _084152_);
  or g_139901_(_079273_, _082233_, _084153_);
  not g_139902_(_084153_, _084154_);
  or g_139903_(_082195_, _082196_, _084155_);
  or g_139904_(_079264_, _082191_, _084157_);
  or g_139905_(_081163_, _082161_, _084158_);
  not g_139906_(_084158_, _084159_);
  or g_139907_(_079240_, _082159_, _084160_);
  and g_139908_(_082137_, _082140_, _084161_);
  or g_139909_(_079206_, _082123_, _084162_);
  and g_139910_(_079202_, _082121_, _084163_);
  or g_139911_(_079201_, _082123_, _084164_);
  or g_139912_(_079188_, _082109_, _084165_);
  not g_139913_(_084165_, _084166_);
  or g_139914_(_079182_, _082109_, _084168_);
  not g_139915_(_084168_, _084169_);
  or g_139916_(_079145_, _082075_, _084170_);
  not g_139917_(_084170_, _084171_);
  or g_139918_(_079140_, _082075_, _084172_);
  and g_139919_(_082074_, _084172_, _084173_);
  and g_139920_(_082052_, _082057_, _084174_);
  not g_139921_(_084174_, _084175_);
  and g_139922_(_081959_, _081961_, _084176_);
  or g_139923_(_079042_, _081929_, _084177_);
  or g_139924_(_079040_, _081929_, _084179_);
  or g_139925_(_079038_, _081926_, _084180_);
  or g_139926_(_079016_, _081903_, _084181_);
  or g_139927_(_079013_, _081903_, _084182_);
  or g_139928_(_078979_, _081866_, _084183_);
  not g_139929_(_084183_, _084184_);
  or g_139930_(_078961_, _081840_, _084185_);
  not g_139931_(_084185_, _084186_);
  or g_139932_(_078942_, _081821_, _084187_);
  or g_139933_(_078902_, _081779_, _084188_);
  not g_139934_(_084188_, _084190_);
  or g_139935_(_078899_, _081779_, _084191_);
  and g_139936_(_081776_, _081778_, _084192_);
  or g_139937_(_078877_, _081767_, _084193_);
  or g_139938_(_075973_, _084193_, _084194_);
  or g_139939_(_075970_, _084193_, _084195_);
  or g_139940_(_081760_, _081763_, _084196_);
  not g_139941_(_084196_, _084197_);
  or g_139942_(_078853_, _081740_, _084198_);
  not g_139943_(_084198_, _084199_);
  or g_139944_(_078826_, _081708_, _084201_);
  and g_139945_(_081667_, _081669_, _084202_);
  not g_139946_(_084202_, _084203_);
  or g_139947_(_081650_, _081651_, _084204_);
  or g_139948_(_078774_, _081646_, _084205_);
  not g_139949_(_084205_, _084206_);
  or g_139950_(_078760_, _081636_, _084207_);
  not g_139951_(_084207_, _084208_);
  or g_139952_(_078758_, _081636_, _084209_);
  not g_139953_(_084209_, _084210_);
  or g_139954_(_081565_, _081567_, _084212_);
  or g_139955_(_081565_, _081566_, _084213_);
  and g_139956_(_081537_, _081540_, _084214_);
  or g_139957_(_078683_, _081525_, _084215_);
  or g_139958_(_078677_, _081525_, _084216_);
  not g_139959_(_084216_, _084217_);
  or g_139960_(_078642_, _081460_, _084218_);
  or g_139961_(_078638_, _081460_, _084219_);
  not g_139962_(_084219_, _084220_);
  and g_139963_(_081456_, _081459_, _084221_);
  and g_139964_(_081449_, _081453_, _084223_);
  or g_139965_(_075642_, _078615_, _084224_);
  or g_139966_(_081437_, _084224_, _084225_);
  or g_139967_(_078615_, _078617_, _084226_);
  or g_139968_(_081437_, _084226_, _084227_);
  not g_139969_(_084227_, _084228_);
  and g_139970_(_081384_, _081386_, _084229_);
  or g_139971_(_078568_, _081381_, _084230_);
  not g_139972_(_084230_, _084231_);
  or g_139973_(_078564_, _081381_, _084232_);
  not g_139974_(_084232_, _084234_);
  or g_139975_(_075594_, _084232_, _084235_);
  and g_139976_(_075593_, _084234_, _084236_);
  not g_139977_(_084236_, _084237_);
  and g_139978_(_078563_, _081377_, _084238_);
  and g_139979_(_081377_, _081379_, _084239_);
  or g_139980_(_078552_, _081369_, _084240_);
  or g_139981_(_078545_, _081366_, _084241_);
  or g_139982_(_078543_, _081366_, _084242_);
  and g_139983_(_081365_, _084242_, _084243_);
  or g_139984_(_081350_, _081353_, _084245_);
  or g_139985_(_078529_, _081344_, _084246_);
  and g_139986_(_081346_, _084246_, _084247_);
  or g_139987_(_078525_, _081340_, _084248_);
  and g_139988_(_081336_, _084248_, _084249_);
  or g_139989_(_078496_, _081320_, _084250_);
  not g_139990_(_084250_, _084251_);
  and g_139991_(_081284_, _081288_, _084252_);
  and g_139992_(_081293_, _081300_, _084253_);
  and g_139993_(_081296_, _084252_, _084254_);
  and g_139994_(_084253_, _084254_, _084256_);
  and g_139995_(_081307_, _084256_, _084257_);
  and g_139996_(_081303_, _084257_, _084258_);
  or g_139997_(_078484_, _081309_, _084259_);
  and g_139998_(_084258_, _084259_, _084260_);
  or g_139999_(_078486_, _081309_, _084261_);
  and g_140000_(_084260_, _084261_, _084262_);
  and g_140001_(_081314_, _084262_, _084263_);
  or g_140002_(_078498_, _081316_, _084264_);
  and g_140003_(_081317_, _084264_, _084265_);
  and g_140004_(_084263_, _084265_, _084267_);
  or g_140005_(_084250_, _084267_, _084268_);
  xor g_140006_(_084251_, _084267_, _084269_);
  or g_140007_(_081325_, _084269_, _084270_);
  xor g_140008_(_081326_, _084269_, _084271_);
  or g_140009_(_081327_, _084271_, _084272_);
  not g_140010_(_084272_, _084273_);
  and g_140011_(_081327_, _084271_, _084274_);
  or g_140012_(_084273_, _084274_, _084275_);
  not g_140013_(_084275_, _084276_);
  and g_140014_(_081333_, _081338_, _084278_);
  xor g_140015_(_084275_, _084278_, _084279_);
  xor g_140016_(_084276_, _084278_, _084280_);
  or g_140017_(_084249_, _084280_, _084281_);
  xor g_140018_(_084249_, _084279_, _084282_);
  not g_140019_(_084282_, _084283_);
  or g_140020_(_084247_, _084282_, _084284_);
  xor g_140021_(_084247_, _084283_, _084285_);
  not g_140022_(_084285_, _084286_);
  or g_140023_(_078538_, _081350_, _084287_);
  and g_140024_(_081349_, _084287_, _084289_);
  or g_140025_(_084285_, _084289_, _084290_);
  xor g_140026_(_084286_, _084289_, _084291_);
  not g_140027_(_084291_, _084292_);
  and g_140028_(_084245_, _084291_, _084293_);
  or g_140029_(_084245_, _084291_, _084294_);
  xor g_140030_(_084245_, _084291_, _084295_);
  xor g_140031_(_084245_, _084292_, _084296_);
  xor g_140032_(_081358_, _084295_, _084297_);
  and g_140033_(_081361_, _084297_, _084298_);
  or g_140034_(_081361_, _084296_, _084300_);
  not g_140035_(_084300_, _084301_);
  or g_140036_(_084298_, _084301_, _084302_);
  not g_140037_(_084302_, _084303_);
  xor g_140038_(_084243_, _084302_, _084304_);
  xor g_140039_(_084243_, _084303_, _084305_);
  or g_140040_(_084241_, _084305_, _084306_);
  xor g_140041_(_084241_, _084304_, _084307_);
  not g_140042_(_084307_, _084308_);
  or g_140043_(_081370_, _084307_, _084309_);
  xor g_140044_(_081370_, _084307_, _084311_);
  xor g_140045_(_081370_, _084308_, _084312_);
  or g_140046_(_084240_, _084312_, _084313_);
  xor g_140047_(_084240_, _084311_, _084314_);
  or g_140048_(_078555_, _081372_, _084315_);
  not g_140049_(_084315_, _084316_);
  or g_140050_(_084314_, _084315_, _084317_);
  and g_140051_(_084314_, _084315_, _084318_);
  xor g_140052_(_084314_, _084316_, _084319_);
  xor g_140053_(_081376_, _084319_, _084320_);
  and g_140054_(_084239_, _084320_, _084322_);
  xor g_140055_(_084239_, _084320_, _084323_);
  and g_140056_(_084238_, _084323_, _084324_);
  or g_140057_(_084238_, _084323_, _084325_);
  xor g_140058_(_084238_, _084323_, _084326_);
  xor g_140059_(_084237_, _084326_, _084327_);
  or g_140060_(_084235_, _084327_, _084328_);
  and g_140061_(_084235_, _084327_, _084329_);
  xor g_140062_(_084235_, _084327_, _084330_);
  xor g_140063_(_084231_, _084330_, _084331_);
  xor g_140064_(_084230_, _084330_, _084333_);
  xor g_140065_(_084229_, _084331_, _084334_);
  not g_140066_(_084334_, _084335_);
  or g_140067_(_081388_, _084334_, _084336_);
  xor g_140068_(_081388_, _084335_, _084337_);
  not g_140069_(_084337_, _084338_);
  or g_140070_(_081393_, _084337_, _084339_);
  and g_140071_(_081393_, _084337_, _084340_);
  xor g_140072_(_081393_, _084338_, _084341_);
  and g_140073_(_081397_, _081403_, _084342_);
  xor g_140074_(_084341_, _084342_, _084344_);
  not g_140075_(_084344_, _084345_);
  or g_140076_(_081402_, _084345_, _084346_);
  xor g_140077_(_081402_, _084344_, _084347_);
  or g_140078_(_081409_, _084347_, _084348_);
  not g_140079_(_084348_, _084349_);
  xor g_140080_(_081409_, _084347_, _084350_);
  not g_140081_(_084350_, _084351_);
  and g_140082_(_081411_, _081419_, _084352_);
  xor g_140083_(_084350_, _084352_, _084353_);
  and g_140084_(_081421_, _081431_, _084355_);
  xor g_140085_(_084353_, _084355_, _084356_);
  and g_140086_(_081433_, _084356_, _084357_);
  not g_140087_(_084357_, _084358_);
  xor g_140088_(_081432_, _084356_, _084359_);
  not g_140089_(_084359_, _084360_);
  and g_140090_(_084228_, _084360_, _084361_);
  not g_140091_(_084361_, _084362_);
  and g_140092_(_084227_, _084359_, _084363_);
  or g_140093_(_084361_, _084363_, _084364_);
  or g_140094_(_084225_, _084364_, _084366_);
  xor g_140095_(_084225_, _084364_, _084367_);
  and g_140096_(_081441_, _081446_, _084368_);
  xor g_140097_(_084367_, _084368_, _084369_);
  or g_140098_(_084223_, _084369_, _084370_);
  xor g_140099_(_084223_, _084369_, _084371_);
  not g_140100_(_084371_, _084372_);
  xor g_140101_(_084221_, _084371_, _084373_);
  or g_140102_(_084219_, _084373_, _084374_);
  xor g_140103_(_084219_, _084373_, _084375_);
  xor g_140104_(_084220_, _084373_, _084377_);
  or g_140105_(_084218_, _084377_, _084378_);
  xor g_140106_(_084218_, _084375_, _084379_);
  not g_140107_(_084379_, _084380_);
  or g_140108_(_081467_, _084379_, _084381_);
  not g_140109_(_084381_, _084382_);
  xor g_140110_(_081467_, _084380_, _084383_);
  not g_140111_(_084383_, _084384_);
  or g_140112_(_081469_, _084383_, _084385_);
  xor g_140113_(_081469_, _084384_, _084386_);
  not g_140114_(_084386_, _084388_);
  and g_140115_(_081471_, _081475_, _084389_);
  xor g_140116_(_084388_, _084389_, _084390_);
  or g_140117_(_081485_, _084390_, _084391_);
  xor g_140118_(_081485_, _084390_, _084392_);
  not g_140119_(_084392_, _084393_);
  or g_140120_(_081478_, _084393_, _084394_);
  xor g_140121_(_081478_, _084392_, _084395_);
  not g_140122_(_084395_, _084396_);
  or g_140123_(_081491_, _084395_, _084397_);
  xor g_140124_(_081491_, _084395_, _084399_);
  xor g_140125_(_081491_, _084396_, _084400_);
  or g_140126_(_081493_, _084400_, _084401_);
  not g_140127_(_084401_, _084402_);
  xor g_140128_(_081493_, _084399_, _084403_);
  or g_140129_(_081496_, _084403_, _084404_);
  xor g_140130_(_081496_, _084403_, _084405_);
  not g_140131_(_084405_, _084406_);
  and g_140132_(_081500_, _084406_, _084407_);
  and g_140133_(_081504_, _084407_, _084408_);
  and g_140134_(_081499_, _084405_, _084410_);
  not g_140135_(_084410_, _084411_);
  and g_140136_(_081503_, _084405_, _084412_);
  or g_140137_(_081504_, _084406_, _084413_);
  or g_140138_(_084410_, _084412_, _084414_);
  or g_140139_(_084408_, _084414_, _084415_);
  and g_140140_(_081507_, _081510_, _084416_);
  or g_140141_(_084415_, _084416_, _084417_);
  xor g_140142_(_084415_, _084416_, _084418_);
  not g_140143_(_084418_, _084419_);
  or g_140144_(_081513_, _084419_, _084421_);
  and g_140145_(_081513_, _084419_, _084422_);
  xor g_140146_(_081513_, _084418_, _084423_);
  not g_140147_(_084423_, _084424_);
  and g_140148_(_081516_, _081520_, _084425_);
  xor g_140149_(_084424_, _084425_, _084426_);
  or g_140150_(_081524_, _084426_, _084427_);
  not g_140151_(_084427_, _084428_);
  xor g_140152_(_081524_, _084426_, _084429_);
  and g_140153_(_084217_, _084429_, _084430_);
  xor g_140154_(_084216_, _084429_, _084432_);
  not g_140155_(_084432_, _084433_);
  or g_140156_(_084215_, _084432_, _084434_);
  and g_140157_(_084215_, _084432_, _084435_);
  xor g_140158_(_084215_, _084433_, _084436_);
  and g_140159_(_081530_, _081533_, _084437_);
  xor g_140160_(_084436_, _084437_, _084438_);
  not g_140161_(_084438_, _084439_);
  or g_140162_(_084214_, _084439_, _084440_);
  xor g_140163_(_084214_, _084438_, _084441_);
  or g_140164_(_081546_, _084441_, _084443_);
  xor g_140165_(_081545_, _084441_, _084444_);
  or g_140166_(_081548_, _084444_, _084445_);
  xor g_140167_(_081549_, _084444_, _084446_);
  not g_140168_(_084446_, _084447_);
  and g_140169_(_081552_, _081560_, _084448_);
  xor g_140170_(_084447_, _084448_, _084449_);
  xor g_140171_(_084446_, _084448_, _084450_);
  or g_140172_(_081559_, _084449_, _084451_);
  xor g_140173_(_081559_, _084450_, _084452_);
  not g_140174_(_084452_, _084454_);
  or g_140175_(_084213_, _084452_, _084455_);
  xor g_140176_(_084213_, _084452_, _084456_);
  xor g_140177_(_084213_, _084454_, _084457_);
  or g_140178_(_084212_, _084457_, _084458_);
  xor g_140179_(_084212_, _084456_, _084459_);
  not g_140180_(_084459_, _084460_);
  or g_140181_(_081574_, _084459_, _084461_);
  not g_140182_(_084461_, _084462_);
  or g_140183_(_081570_, _084459_, _084463_);
  xor g_140184_(_081570_, _084460_, _084465_);
  not g_140185_(_084465_, _084466_);
  or g_140186_(_081576_, _084465_, _084467_);
  xor g_140187_(_081576_, _084466_, _084468_);
  and g_140188_(_081574_, _084468_, _084469_);
  or g_140189_(_084462_, _084469_, _084470_);
  not g_140190_(_084470_, _084471_);
  or g_140191_(_081579_, _084470_, _084472_);
  xor g_140192_(_081579_, _084470_, _084473_);
  xor g_140193_(_081579_, _084471_, _084474_);
  or g_140194_(_081582_, _084474_, _084476_);
  xor g_140195_(_081582_, _084473_, _084477_);
  or g_140196_(_081589_, _084477_, _084478_);
  not g_140197_(_084478_, _084479_);
  and g_140198_(_081589_, _084477_, _084480_);
  not g_140199_(_084480_, _084481_);
  and g_140200_(_084478_, _084481_, _084482_);
  or g_140201_(_084479_, _084480_, _084483_);
  or g_140202_(_081593_, _084483_, _084484_);
  not g_140203_(_084484_, _084485_);
  and g_140204_(_081586_, _084482_, _084487_);
  xor g_140205_(_081585_, _084482_, _084488_);
  and g_140206_(_081593_, _084488_, _084489_);
  or g_140207_(_084485_, _084489_, _084490_);
  or g_140208_(_081599_, _084490_, _084491_);
  not g_140209_(_084491_, _084492_);
  or g_140210_(_078733_, _081595_, _084493_);
  or g_140211_(_078730_, _081595_, _084494_);
  or g_140212_(_084490_, _084494_, _084495_);
  xor g_140213_(_084490_, _084494_, _084496_);
  not g_140214_(_084496_, _084498_);
  or g_140215_(_084493_, _084498_, _084499_);
  not g_140216_(_084499_, _084500_);
  xor g_140217_(_084493_, _084496_, _084501_);
  and g_140218_(_081599_, _084501_, _084502_);
  or g_140219_(_084492_, _084502_, _084503_);
  or g_140220_(_081606_, _084503_, _084504_);
  xor g_140221_(_081607_, _084503_, _084505_);
  or g_140222_(_081601_, _084505_, _084506_);
  xor g_140223_(_081602_, _084505_, _084507_);
  not g_140224_(_084507_, _084509_);
  or g_140225_(_081621_, _084507_, _084510_);
  not g_140226_(_084510_, _084511_);
  or g_140227_(_081611_, _084507_, _084512_);
  xor g_140228_(_081611_, _084507_, _084513_);
  xor g_140229_(_081611_, _084509_, _084514_);
  and g_140230_(_081621_, _084514_, _084515_);
  or g_140231_(_081620_, _084513_, _084516_);
  and g_140232_(_084510_, _084516_, _084517_);
  or g_140233_(_084511_, _084515_, _084518_);
  and g_140234_(_081629_, _084517_, _084520_);
  or g_140235_(_081628_, _084518_, _084521_);
  and g_140236_(_067877_, _084520_, _084522_);
  or g_140237_(_067876_, _084521_, _084523_);
  and g_140238_(_081630_, _084518_, _084524_);
  or g_140239_(_084522_, _084524_, _084525_);
  not g_140240_(_084525_, _084526_);
  and g_140241_(_081633_, _081635_, _084527_);
  xor g_140242_(_084526_, _084527_, _084528_);
  not g_140243_(_084528_, _084529_);
  and g_140244_(_084210_, _084529_, _084531_);
  not g_140245_(_084531_, _084532_);
  xor g_140246_(_084209_, _084528_, _084533_);
  and g_140247_(_084208_, _084533_, _084534_);
  xor g_140248_(_084207_, _084533_, _084535_);
  or g_140249_(_081643_, _084535_, _084536_);
  xor g_140250_(_081643_, _084535_, _084537_);
  not g_140251_(_084537_, _084538_);
  and g_140252_(_078770_, _081641_, _084539_);
  or g_140253_(_081645_, _084539_, _084540_);
  xor g_140254_(_084537_, _084540_, _084542_);
  or g_140255_(_084205_, _084542_, _084543_);
  xor g_140256_(_084206_, _084542_, _084544_);
  not g_140257_(_084544_, _084545_);
  or g_140258_(_084204_, _084544_, _084546_);
  xor g_140259_(_084204_, _084545_, _084547_);
  not g_140260_(_084547_, _084548_);
  and g_140261_(_081656_, _084548_, _084549_);
  or g_140262_(_081657_, _084547_, _084550_);
  xor g_140263_(_081656_, _084547_, _084551_);
  not g_140264_(_084551_, _084553_);
  or g_140265_(_081661_, _084551_, _084554_);
  xor g_140266_(_081661_, _084551_, _084555_);
  xor g_140267_(_081661_, _084553_, _084556_);
  xor g_140268_(_081664_, _084555_, _084557_);
  xor g_140269_(_084202_, _084557_, _084558_);
  xor g_140270_(_084203_, _084557_, _084559_);
  or g_140271_(_081672_, _084559_, _084560_);
  xor g_140272_(_081672_, _084558_, _084561_);
  not g_140273_(_084561_, _084562_);
  or g_140274_(_081678_, _084561_, _084564_);
  xor g_140275_(_081678_, _084561_, _084565_);
  xor g_140276_(_081678_, _084562_, _084566_);
  or g_140277_(_081676_, _084566_, _084567_);
  not g_140278_(_084567_, _084568_);
  or g_140279_(_081680_, _084561_, _084569_);
  not g_140280_(_084569_, _084570_);
  and g_140281_(_081680_, _084566_, _084571_);
  or g_140282_(_081681_, _084565_, _084572_);
  and g_140283_(_084569_, _084572_, _084573_);
  or g_140284_(_084570_, _084571_, _084575_);
  and g_140285_(_081676_, _084575_, _084576_);
  or g_140286_(_081677_, _084573_, _084577_);
  and g_140287_(_084567_, _084577_, _084578_);
  or g_140288_(_084568_, _084576_, _084579_);
  or g_140289_(_081686_, _084579_, _084580_);
  xor g_140290_(_081686_, _084578_, _084581_);
  or g_140291_(_081696_, _084581_, _084582_);
  not g_140292_(_084582_, _084583_);
  and g_140293_(_081694_, _084581_, _084584_);
  and g_140294_(_081696_, _084584_, _084586_);
  or g_140295_(_081694_, _084581_, _084587_);
  not g_140296_(_084587_, _084588_);
  or g_140297_(_084586_, _084588_, _084589_);
  or g_140298_(_084583_, _084589_, _084590_);
  and g_140299_(_081700_, _081705_, _084591_);
  not g_140300_(_084591_, _084592_);
  or g_140301_(_084590_, _084591_, _084593_);
  xor g_140302_(_084590_, _084592_, _084594_);
  and g_140303_(_081707_, _081709_, _084595_);
  not g_140304_(_084595_, _084597_);
  xor g_140305_(_084594_, _084597_, _084598_);
  not g_140306_(_084598_, _084599_);
  or g_140307_(_084201_, _084598_, _084600_);
  xor g_140308_(_084201_, _084598_, _084601_);
  xor g_140309_(_084201_, _084599_, _084602_);
  or g_140310_(_078830_, _081710_, _084603_);
  and g_140311_(_081716_, _084603_, _084604_);
  xor g_140312_(_084601_, _084604_, _084605_);
  or g_140313_(_081718_, _084605_, _084606_);
  xor g_140314_(_081719_, _084605_, _084608_);
  or g_140315_(_081722_, _084608_, _084609_);
  xor g_140316_(_081723_, _084608_, _084610_);
  and g_140317_(_081734_, _084610_, _084611_);
  or g_140318_(_081728_, _084608_, _084612_);
  or g_140319_(_081732_, _084610_, _084613_);
  and g_140320_(_084612_, _084613_, _084614_);
  not g_140321_(_084614_, _084615_);
  or g_140322_(_084611_, _084615_, _084616_);
  or g_140323_(_078850_, _081740_, _084617_);
  and g_140324_(_081739_, _084617_, _084619_);
  or g_140325_(_084616_, _084619_, _084620_);
  xor g_140326_(_084616_, _084619_, _084621_);
  not g_140327_(_084621_, _084622_);
  and g_140328_(_084199_, _084621_, _084623_);
  or g_140329_(_084198_, _084622_, _084624_);
  xor g_140330_(_084198_, _084621_, _084625_);
  not g_140331_(_084625_, _084626_);
  and g_140332_(_081744_, _081747_, _084627_);
  xor g_140333_(_084626_, _084627_, _084628_);
  xor g_140334_(_084625_, _084627_, _084630_);
  or g_140335_(_081751_, _084628_, _084631_);
  xor g_140336_(_081751_, _084630_, _084632_);
  not g_140337_(_084632_, _084633_);
  and g_140338_(_081753_, _081756_, _084634_);
  xor g_140339_(_084633_, _084634_, _084635_);
  or g_140340_(_081758_, _084635_, _084636_);
  xor g_140341_(_081758_, _084635_, _084637_);
  not g_140342_(_084637_, _084638_);
  and g_140343_(_084197_, _084637_, _084639_);
  or g_140344_(_084196_, _084638_, _084641_);
  xor g_140345_(_084196_, _084637_, _084642_);
  or g_140346_(_081760_, _081764_, _084643_);
  and g_140347_(_081768_, _084643_, _084644_);
  and g_140348_(_084642_, _084644_, _084645_);
  or g_140349_(_084642_, _084643_, _084646_);
  or g_140350_(_081768_, _084642_, _084647_);
  and g_140351_(_084646_, _084647_, _084648_);
  not g_140352_(_084648_, _084649_);
  or g_140353_(_084645_, _084649_, _084650_);
  and g_140354_(_084195_, _084650_, _084652_);
  or g_140355_(_084195_, _084650_, _084653_);
  not g_140356_(_084653_, _084654_);
  or g_140357_(_084652_, _084654_, _084655_);
  not g_140358_(_084655_, _084656_);
  or g_140359_(_084194_, _084655_, _084657_);
  xor g_140360_(_084194_, _084656_, _084658_);
  not g_140361_(_084658_, _084659_);
  or g_140362_(_078884_, _081771_, _084660_);
  and g_140363_(_081774_, _084660_, _084661_);
  xor g_140364_(_084659_, _084661_, _084663_);
  xor g_140365_(_084192_, _084663_, _084664_);
  not g_140366_(_084664_, _084665_);
  or g_140367_(_084191_, _084665_, _084666_);
  xor g_140368_(_084191_, _084664_, _084667_);
  or g_140369_(_084188_, _084667_, _084668_);
  xor g_140370_(_084190_, _084667_, _084669_);
  or g_140371_(_081786_, _084669_, _084670_);
  not g_140372_(_084670_, _084671_);
  xor g_140373_(_081785_, _084669_, _084672_);
  not g_140374_(_084672_, _084674_);
  and g_140375_(_081789_, _084674_, _084675_);
  or g_140376_(_081790_, _084672_, _084676_);
  xor g_140377_(_081790_, _084672_, _084677_);
  xor g_140378_(_081789_, _084672_, _084678_);
  or g_140379_(_081793_, _084678_, _084679_);
  xor g_140380_(_081793_, _084677_, _084680_);
  or g_140381_(_081797_, _084680_, _084681_);
  xor g_140382_(_081797_, _084680_, _084682_);
  xor g_140383_(_081796_, _084680_, _084683_);
  or g_140384_(_081798_, _084683_, _084685_);
  xor g_140385_(_081798_, _084682_, _084686_);
  not g_140386_(_084686_, _084687_);
  or g_140387_(_081802_, _084686_, _084688_);
  xor g_140388_(_081802_, _084687_, _084689_);
  or g_140389_(_078927_, _081805_, _084690_);
  and g_140390_(_081806_, _084690_, _084691_);
  xor g_140391_(_084689_, _084691_, _084692_);
  not g_140392_(_084692_, _084693_);
  or g_140393_(_081812_, _084693_, _084694_);
  not g_140394_(_084694_, _084696_);
  xor g_140395_(_081812_, _084692_, _084697_);
  and g_140396_(_081816_, _081818_, _084698_);
  not g_140397_(_084698_, _084699_);
  xor g_140398_(_084697_, _084699_, _084700_);
  not g_140399_(_084700_, _084701_);
  or g_140400_(_078940_, _081821_, _084702_);
  and g_140401_(_081820_, _084702_, _084703_);
  or g_140402_(_084700_, _084703_, _084704_);
  xor g_140403_(_084700_, _084703_, _084705_);
  xor g_140404_(_084701_, _084703_, _084707_);
  or g_140405_(_084187_, _084707_, _084708_);
  xor g_140406_(_084187_, _084705_, _084709_);
  or g_140407_(_081828_, _084709_, _084710_);
  not g_140408_(_084710_, _084711_);
  xor g_140409_(_081827_, _084709_, _084712_);
  not g_140410_(_084712_, _084713_);
  or g_140411_(_081833_, _084712_, _084714_);
  not g_140412_(_084714_, _084715_);
  and g_140413_(_081835_, _084713_, _084716_);
  xor g_140414_(_081835_, _084712_, _084718_);
  and g_140415_(_081833_, _084718_, _084719_);
  or g_140416_(_084715_, _084719_, _084720_);
  not g_140417_(_084720_, _084721_);
  and g_140418_(_081839_, _084721_, _084722_);
  xor g_140419_(_081839_, _084720_, _084723_);
  or g_140420_(_078958_, _081837_, _084724_);
  not g_140421_(_084724_, _084725_);
  or g_140422_(_084723_, _084724_, _084726_);
  xor g_140423_(_084723_, _084725_, _084727_);
  or g_140424_(_084185_, _084727_, _084729_);
  xor g_140425_(_084186_, _084727_, _084730_);
  or g_140426_(_081856_, _084730_, _084731_);
  not g_140427_(_084731_, _084732_);
  xor g_140428_(_081850_, _084730_, _084733_);
  xor g_140429_(_081851_, _084730_, _084734_);
  or g_140430_(_081860_, _084734_, _084735_);
  not g_140431_(_084735_, _084736_);
  xor g_140432_(_081860_, _084733_, _084737_);
  and g_140433_(_081856_, _084737_, _084738_);
  or g_140434_(_084732_, _084738_, _084740_);
  or g_140435_(_081863_, _084740_, _084741_);
  not g_140436_(_084741_, _084742_);
  xor g_140437_(_081864_, _084740_, _084743_);
  or g_140438_(_078976_, _081861_, _084744_);
  or g_140439_(_084743_, _084744_, _084745_);
  not g_140440_(_084745_, _084746_);
  xor g_140441_(_084743_, _084744_, _084747_);
  not g_140442_(_084747_, _084748_);
  and g_140443_(_084184_, _084747_, _084749_);
  or g_140444_(_084183_, _084748_, _084751_);
  xor g_140445_(_084183_, _084747_, _084752_);
  not g_140446_(_084752_, _084753_);
  or g_140447_(_081870_, _084752_, _084754_);
  xor g_140448_(_081870_, _084752_, _084755_);
  xor g_140449_(_081870_, _084753_, _084756_);
  and g_140450_(_081874_, _081875_, _084757_);
  xor g_140451_(_084755_, _084757_, _084758_);
  not g_140452_(_084758_, _084759_);
  and g_140453_(_081879_, _081883_, _084760_);
  xor g_140454_(_084759_, _084760_, _084762_);
  xor g_140455_(_084758_, _084760_, _084763_);
  or g_140456_(_081889_, _084762_, _084764_);
  not g_140457_(_084764_, _084765_);
  xor g_140458_(_081889_, _084763_, _084766_);
  or g_140459_(_079007_, _081894_, _084767_);
  and g_140460_(_081892_, _084767_, _084768_);
  xor g_140461_(_084766_, _084768_, _084769_);
  not g_140462_(_084769_, _084770_);
  or g_140463_(_081894_, _081896_, _084771_);
  and g_140464_(_081900_, _084771_, _084773_);
  xor g_140465_(_084769_, _084773_, _084774_);
  not g_140466_(_084774_, _084775_);
  or g_140467_(_084182_, _084774_, _084776_);
  xor g_140468_(_084182_, _084775_, _084777_);
  not g_140469_(_084777_, _084778_);
  or g_140470_(_084181_, _084777_, _084779_);
  xor g_140471_(_084181_, _084778_, _084780_);
  or g_140472_(_081907_, _084780_, _084781_);
  not g_140473_(_084781_, _084782_);
  or g_140474_(_081916_, _084780_, _084784_);
  xor g_140475_(_081915_, _084780_, _084785_);
  and g_140476_(_081907_, _084785_, _084786_);
  or g_140477_(_084782_, _084786_, _084787_);
  or g_140478_(_081920_, _084787_, _084788_);
  not g_140479_(_084788_, _084789_);
  or g_140480_(_081912_, _084787_, _084790_);
  xor g_140481_(_081914_, _084787_, _084791_);
  and g_140482_(_081920_, _084791_, _084792_);
  or g_140483_(_084789_, _084792_, _084793_);
  not g_140484_(_084793_, _084795_);
  or g_140485_(_079036_, _081926_, _084796_);
  and g_140486_(_081925_, _084796_, _084797_);
  xor g_140487_(_084793_, _084797_, _084798_);
  xor g_140488_(_084795_, _084797_, _084799_);
  or g_140489_(_084180_, _084799_, _084800_);
  xor g_140490_(_084180_, _084798_, _084801_);
  not g_140491_(_084801_, _084802_);
  or g_140492_(_084179_, _084801_, _084803_);
  xor g_140493_(_084179_, _084801_, _084804_);
  xor g_140494_(_084179_, _084802_, _084806_);
  or g_140495_(_084177_, _084806_, _084807_);
  xor g_140496_(_084177_, _084804_, _084808_);
  or g_140497_(_081936_, _084808_, _084809_);
  xor g_140498_(_081936_, _084808_, _084810_);
  xor g_140499_(_081937_, _084808_, _084811_);
  and g_140500_(_081940_, _081942_, _084812_);
  xor g_140501_(_084810_, _084812_, _084813_);
  or g_140502_(_081945_, _084813_, _084814_);
  not g_140503_(_084814_, _084815_);
  xor g_140504_(_081945_, _084813_, _084817_);
  not g_140505_(_084817_, _084818_);
  or g_140506_(_081950_, _084818_, _084819_);
  xor g_140507_(_081949_, _084817_, _084820_);
  not g_140508_(_084820_, _084821_);
  or g_140509_(_081952_, _084821_, _084822_);
  xor g_140510_(_081952_, _084820_, _084823_);
  not g_140511_(_084823_, _084824_);
  xor g_140512_(_081955_, _084824_, _084825_);
  xor g_140513_(_084176_, _084825_, _084826_);
  not g_140514_(_084826_, _084828_);
  or g_140515_(_081966_, _084828_, _084829_);
  xor g_140516_(_081966_, _084826_, _084830_);
  not g_140517_(_084830_, _084831_);
  or g_140518_(_081977_, _084830_, _084832_);
  xor g_140519_(_081977_, _084831_, _084833_);
  or g_140520_(_081976_, _084833_, _084834_);
  xor g_140521_(_081976_, _084833_, _084835_);
  not g_140522_(_084835_, _084836_);
  or g_140523_(_081983_, _084836_, _084837_);
  xor g_140524_(_081983_, _084835_, _084839_);
  not g_140525_(_084839_, _084840_);
  or g_140526_(_081985_, _084839_, _084841_);
  xor g_140527_(_081985_, _084840_, _084842_);
  or g_140528_(_081994_, _084842_, _084843_);
  not g_140529_(_084843_, _084844_);
  or g_140530_(_082002_, _084842_, _084845_);
  xor g_140531_(_082002_, _084842_, _084846_);
  or g_140532_(_081993_, _084846_, _084847_);
  not g_140533_(_084847_, _084848_);
  or g_140534_(_084844_, _084848_, _084850_);
  or g_140535_(_081999_, _084850_, _084851_);
  xor g_140536_(_082000_, _084850_, _084852_);
  not g_140537_(_084852_, _084853_);
  and g_140538_(_082006_, _082008_, _084854_);
  or g_140539_(_084852_, _084854_, _084855_);
  xor g_140540_(_084852_, _084854_, _084856_);
  xor g_140541_(_084853_, _084854_, _084857_);
  or g_140542_(_082014_, _084857_, _084858_);
  xor g_140543_(_082014_, _084856_, _084859_);
  not g_140544_(_084859_, _084861_);
  or g_140545_(_082015_, _084859_, _084862_);
  xor g_140546_(_082015_, _084859_, _084863_);
  xor g_140547_(_082015_, _084861_, _084864_);
  or g_140548_(_082019_, _084864_, _084865_);
  xor g_140549_(_082019_, _084863_, _084866_);
  not g_140550_(_084866_, _084867_);
  and g_140551_(_082028_, _084867_, _084868_);
  xor g_140552_(_082027_, _084866_, _084869_);
  xor g_140553_(_082028_, _084866_, _084870_);
  or g_140554_(_082036_, _084870_, _084872_);
  xor g_140555_(_082036_, _084869_, _084873_);
  not g_140556_(_084873_, _084874_);
  or g_140557_(_082038_, _084873_, _084875_);
  xor g_140558_(_082038_, _084873_, _084876_);
  xor g_140559_(_082038_, _084874_, _084877_);
  and g_140560_(_082041_, _082044_, _084878_);
  xor g_140561_(_084876_, _084878_, _084879_);
  not g_140562_(_084879_, _084880_);
  and g_140563_(_082047_, _082050_, _084881_);
  xor g_140564_(_084880_, _084881_, _084883_);
  or g_140565_(_084174_, _084883_, _084884_);
  xor g_140566_(_084174_, _084883_, _084885_);
  xor g_140567_(_084175_, _084883_, _084886_);
  or g_140568_(_082062_, _084886_, _084887_);
  not g_140569_(_084887_, _084888_);
  or g_140570_(_082059_, _084886_, _084889_);
  xor g_140571_(_082059_, _084885_, _084890_);
  or g_140572_(_082065_, _084890_, _084891_);
  xor g_140573_(_082066_, _084890_, _084892_);
  and g_140574_(_082062_, _084892_, _084894_);
  or g_140575_(_084888_, _084894_, _084895_);
  not g_140576_(_084895_, _084896_);
  and g_140577_(_082069_, _082071_, _084897_);
  xor g_140578_(_084895_, _084897_, _084898_);
  xor g_140579_(_084896_, _084897_, _084899_);
  xor g_140580_(_084173_, _084898_, _084900_);
  or g_140581_(_084170_, _084900_, _084901_);
  xor g_140582_(_084170_, _084900_, _084902_);
  xor g_140583_(_084171_, _084900_, _084903_);
  or g_140584_(_082081_, _084903_, _084905_);
  xor g_140585_(_082081_, _084902_, _084906_);
  xor g_140586_(_082085_, _084906_, _084907_);
  or g_140587_(_082090_, _084907_, _084908_);
  xor g_140588_(_082088_, _084907_, _084909_);
  or g_140589_(_082093_, _084909_, _084910_);
  xor g_140590_(_082094_, _084909_, _084911_);
  or g_140591_(_082097_, _084911_, _084912_);
  not g_140592_(_084912_, _084913_);
  or g_140593_(_082102_, _084911_, _084914_);
  not g_140594_(_084914_, _084916_);
  xor g_140595_(_082102_, _084911_, _084917_);
  xor g_140596_(_082103_, _084911_, _084918_);
  and g_140597_(_082097_, _084918_, _084919_);
  or g_140598_(_082098_, _084917_, _084920_);
  and g_140599_(_084912_, _084920_, _084921_);
  or g_140600_(_084913_, _084919_, _084922_);
  or g_140601_(_079176_, _082106_, _084923_);
  and g_140602_(_082105_, _084923_, _084924_);
  xor g_140603_(_084922_, _084924_, _084925_);
  xor g_140604_(_084921_, _084924_, _084927_);
  or g_140605_(_079179_, _082106_, _084928_);
  not g_140606_(_084928_, _084929_);
  and g_140607_(_084927_, _084928_, _084930_);
  and g_140608_(_084168_, _084930_, _084931_);
  and g_140609_(_084169_, _084925_, _084932_);
  or g_140610_(_084168_, _084927_, _084933_);
  and g_140611_(_084925_, _084929_, _084934_);
  not g_140612_(_084934_, _084935_);
  or g_140613_(_084932_, _084934_, _084936_);
  or g_140614_(_084931_, _084936_, _084938_);
  or g_140615_(_084165_, _084938_, _084939_);
  xor g_140616_(_084165_, _084938_, _084940_);
  xor g_140617_(_084166_, _084938_, _084941_);
  and g_140618_(_082113_, _082116_, _084942_);
  xor g_140619_(_084940_, _084942_, _084943_);
  not g_140620_(_084943_, _084944_);
  xor g_140621_(_082120_, _084944_, _084945_);
  or g_140622_(_084164_, _084945_, _084946_);
  not g_140623_(_084946_, _084947_);
  xor g_140624_(_084163_, _084945_, _084949_);
  not g_140625_(_084949_, _084950_);
  or g_140626_(_084162_, _084949_, _084951_);
  not g_140627_(_084951_, _084952_);
  xor g_140628_(_084162_, _084950_, _084953_);
  or g_140629_(_082125_, _084953_, _084954_);
  not g_140630_(_084954_, _084955_);
  xor g_140631_(_082126_, _084953_, _084956_);
  and g_140632_(_082130_, _082134_, _084957_);
  xor g_140633_(_084956_, _084957_, _084958_);
  not g_140634_(_084958_, _084960_);
  xor g_140635_(_084161_, _084958_, _084961_);
  or g_140636_(_082143_, _084961_, _084962_);
  xor g_140637_(_082145_, _084961_, _084963_);
  not g_140638_(_084963_, _084964_);
  and g_140639_(_082148_, _082151_, _084965_);
  xor g_140640_(_084964_, _084965_, _084966_);
  or g_140641_(_082153_, _084966_, _084967_);
  xor g_140642_(_082154_, _084966_, _084968_);
  not g_140643_(_084968_, _084969_);
  or g_140644_(_079236_, _082159_, _084971_);
  and g_140645_(_082157_, _084971_, _084972_);
  xor g_140646_(_084968_, _084972_, _084973_);
  xor g_140647_(_084969_, _084972_, _084974_);
  or g_140648_(_084160_, _084974_, _084975_);
  not g_140649_(_084975_, _084976_);
  xor g_140650_(_084160_, _084973_, _084977_);
  or g_140651_(_082162_, _084977_, _084978_);
  xor g_140652_(_082163_, _084977_, _084979_);
  or g_140653_(_084158_, _084979_, _084980_);
  xor g_140654_(_084158_, _084979_, _084982_);
  xor g_140655_(_084159_, _084979_, _084983_);
  and g_140656_(_082167_, _084983_, _084984_);
  and g_140657_(_082172_, _084984_, _084985_);
  and g_140658_(_082171_, _084982_, _084986_);
  or g_140659_(_082172_, _084983_, _084987_);
  and g_140660_(_082168_, _084982_, _084988_);
  or g_140661_(_084986_, _084988_, _084989_);
  or g_140662_(_084985_, _084989_, _084990_);
  xor g_140663_(_082179_, _084990_, _084991_);
  not g_140664_(_084991_, _084993_);
  or g_140665_(_082186_, _084991_, _084994_);
  xor g_140666_(_082186_, _084991_, _084995_);
  xor g_140667_(_082186_, _084993_, _084996_);
  and g_140668_(_082190_, _084995_, _084997_);
  or g_140669_(_082189_, _084996_, _084998_);
  or g_140670_(_082193_, _084996_, _084999_);
  not g_140671_(_084999_, _085000_);
  xor g_140672_(_082193_, _084995_, _085001_);
  and g_140673_(_082189_, _085001_, _085002_);
  or g_140674_(_084997_, _085002_, _085004_);
  or g_140675_(_084157_, _085004_, _085005_);
  not g_140676_(_085005_, _085006_);
  xor g_140677_(_084157_, _085004_, _085007_);
  not g_140678_(_085007_, _085008_);
  or g_140679_(_084155_, _085008_, _085009_);
  xor g_140680_(_084155_, _085007_, _085010_);
  or g_140681_(_082200_, _085010_, _085011_);
  xor g_140682_(_082201_, _085010_, _085012_);
  or g_140683_(_082204_, _085012_, _085013_);
  xor g_140684_(_082205_, _085012_, _085015_);
  and g_140685_(_082209_, _082212_, _085016_);
  xor g_140686_(_085015_, _085016_, _085017_);
  and g_140687_(_082217_, _085017_, _085018_);
  xor g_140688_(_082216_, _085017_, _085019_);
  or g_140689_(_082219_, _085019_, _085020_);
  xor g_140690_(_082220_, _085019_, _085021_);
  or g_140691_(_082227_, _085021_, _085022_);
  xor g_140692_(_082227_, _085021_, _085023_);
  xor g_140693_(_082226_, _085021_, _085024_);
  or g_140694_(_084153_, _085024_, _085026_);
  not g_140695_(_085026_, _085027_);
  and g_140696_(_082230_, _085024_, _085028_);
  or g_140697_(_082231_, _085023_, _085029_);
  and g_140698_(_084153_, _085028_, _085030_);
  or g_140699_(_084154_, _085029_, _085031_);
  or g_140700_(_082230_, _085024_, _085032_);
  not g_140701_(_085032_, _085033_);
  and g_140702_(_085031_, _085032_, _085034_);
  or g_140703_(_085030_, _085033_, _085035_);
  and g_140704_(_085026_, _085034_, _085037_);
  or g_140705_(_085027_, _085035_, _085038_);
  or g_140706_(_079277_, _082233_, _085039_);
  not g_140707_(_085039_, _085040_);
  and g_140708_(_085038_, _085039_, _085041_);
  or g_140709_(_085037_, _085040_, _085042_);
  and g_140710_(_082237_, _085041_, _085043_);
  or g_140711_(_082238_, _085042_, _085044_);
  or g_140712_(_082237_, _085038_, _085045_);
  not g_140713_(_085045_, _085046_);
  or g_140714_(_085038_, _085039_, _085048_);
  not g_140715_(_085048_, _085049_);
  and g_140716_(_085045_, _085048_, _085050_);
  not g_140717_(_085050_, _085051_);
  and g_140718_(_085044_, _085050_, _085052_);
  or g_140719_(_085043_, _085051_, _085053_);
  or g_140720_(_084152_, _085053_, _085054_);
  xor g_140721_(_084152_, _085052_, _085055_);
  or g_140722_(_084151_, _085055_, _085056_);
  xor g_140723_(_084150_, _085055_, _085057_);
  and g_140724_(_082247_, _085057_, _085059_);
  or g_140725_(_082247_, _085057_, _085060_);
  not g_140726_(_085060_, _085061_);
  xor g_140727_(_082247_, _085057_, _085062_);
  or g_140728_(_085059_, _085061_, _085063_);
  or g_140729_(_082251_, _085063_, _085064_);
  not g_140730_(_085064_, _085065_);
  xor g_140731_(_082251_, _085062_, _085066_);
  or g_140732_(_082253_, _085066_, _085067_);
  xor g_140733_(_082252_, _085066_, _085068_);
  and g_140734_(_082258_, _082260_, _085070_);
  xor g_140735_(_085068_, _085070_, _085071_);
  not g_140736_(_085071_, _085072_);
  or g_140737_(_084149_, _085072_, _085073_);
  not g_140738_(_085073_, _085074_);
  xor g_140739_(_084149_, _085071_, _085075_);
  or g_140740_(_084147_, _085075_, _085076_);
  xor g_140741_(_084148_, _085075_, _085077_);
  or g_140742_(_082267_, _085077_, _085078_);
  not g_140743_(_085078_, _085079_);
  xor g_140744_(_082266_, _085077_, _085081_);
  or g_140745_(_084146_, _085081_, _085082_);
  not g_140746_(_085082_, _085083_);
  xor g_140747_(_084146_, _085081_, _085084_);
  not g_140748_(_085084_, _085085_);
  or g_140749_(_082273_, _085085_, _085086_);
  not g_140750_(_085086_, _085087_);
  and g_140751_(_079320_, _082269_, _085088_);
  not g_140752_(_085088_, _085089_);
  or g_140753_(_085084_, _085088_, _085090_);
  or g_140754_(_085081_, _085089_, _085092_);
  not g_140755_(_085092_, _085093_);
  and g_140756_(_085090_, _085092_, _085094_);
  not g_140757_(_085094_, _085095_);
  or g_140758_(_082277_, _085095_, _085096_);
  xor g_140759_(_082275_, _085094_, _085097_);
  or g_140760_(_082272_, _085097_, _085098_);
  not g_140761_(_085098_, _085099_);
  and g_140762_(_085086_, _085098_, _085100_);
  or g_140763_(_085087_, _085099_, _085101_);
  or g_140764_(_082279_, _085101_, _085103_);
  not g_140765_(_085103_, _085104_);
  xor g_140766_(_082279_, _085100_, _085105_);
  not g_140767_(_085105_, _085106_);
  or g_140768_(_082282_, _085105_, _085107_);
  not g_140769_(_085107_, _085108_);
  xor g_140770_(_082282_, _085105_, _085109_);
  xor g_140771_(_082282_, _085106_, _085110_);
  or g_140772_(_082286_, _085110_, _085111_);
  xor g_140773_(_082286_, _085109_, _085112_);
  not g_140774_(_085112_, _085114_);
  or g_140775_(_082290_, _085112_, _085115_);
  xor g_140776_(_082290_, _085112_, _085116_);
  xor g_140777_(_082290_, _085114_, _085117_);
  or g_140778_(_082295_, _085117_, _085118_);
  xor g_140779_(_082295_, _085116_, _085119_);
  not g_140780_(_085119_, _085120_);
  and g_140781_(_082293_, _082297_, _085121_);
  not g_140782_(_085121_, _085122_);
  xor g_140783_(_085119_, _085122_, _085123_);
  or g_140784_(_079354_, _082304_, _085125_);
  and g_140785_(_082303_, _085125_, _085126_);
  not g_140786_(_085126_, _085127_);
  xor g_140787_(_085123_, _085127_, _085128_);
  or g_140788_(_079357_, _082304_, _085129_);
  or g_140789_(_079360_, _082307_, _085130_);
  and g_140790_(_085129_, _085130_, _085131_);
  xor g_140791_(_085128_, _085131_, _085132_);
  not g_140792_(_085132_, _085133_);
  or g_140793_(_084144_, _085133_, _085134_);
  not g_140794_(_085134_, _085136_);
  xor g_140795_(_084144_, _085132_, _085137_);
  not g_140796_(_085137_, _085138_);
  or g_140797_(_082311_, _085137_, _085139_);
  xor g_140798_(_082311_, _085137_, _085140_);
  xor g_140799_(_082311_, _085138_, _085141_);
  or g_140800_(_082313_, _085141_, _085142_);
  xor g_140801_(_082313_, _085140_, _085143_);
  or g_140802_(_082315_, _085143_, _085144_);
  not g_140803_(_085144_, _085145_);
  xor g_140804_(_082315_, _085143_, _085147_);
  not g_140805_(_085147_, _085148_);
  or g_140806_(_084143_, _085148_, _085149_);
  not g_140807_(_085149_, _085150_);
  xor g_140808_(_084143_, _085147_, _085151_);
  or g_140809_(_084142_, _085151_, _085152_);
  not g_140810_(_085152_, _085153_);
  xor g_140811_(_084141_, _085151_, _085154_);
  or g_140812_(_084140_, _085154_, _085155_);
  not g_140813_(_085155_, _085156_);
  and g_140814_(_084140_, _085154_, _085158_);
  xor g_140815_(_084140_, _085154_, _085159_);
  or g_140816_(_085156_, _085158_, _085160_);
  or g_140817_(_079382_, _082319_, _085161_);
  not g_140818_(_085161_, _085162_);
  and g_140819_(_082324_, _085161_, _085163_);
  xor g_140820_(_085159_, _085163_, _085164_);
  not g_140821_(_085164_, _085165_);
  and g_140822_(_082327_, _082329_, _085166_);
  xor g_140823_(_085165_, _085166_, _085167_);
  xor g_140824_(_085164_, _085166_, _085169_);
  or g_140825_(_082338_, _085169_, _085170_);
  and g_140826_(_082334_, _085169_, _085171_);
  or g_140827_(_082333_, _085167_, _085172_);
  or g_140828_(_082335_, _085167_, _085173_);
  not g_140829_(_085173_, _085174_);
  and g_140830_(_085172_, _085173_, _085175_);
  not g_140831_(_085175_, _085176_);
  and g_140832_(_085170_, _085175_, _085177_);
  and g_140833_(_082354_, _085177_, _085178_);
  xor g_140834_(_082352_, _085177_, _085180_);
  not g_140835_(_085180_, _085181_);
  and g_140836_(_082347_, _085181_, _085182_);
  not g_140837_(_085182_, _085183_);
  xor g_140838_(_082347_, _085180_, _085184_);
  not g_140839_(_085184_, _085185_);
  or g_140840_(_082360_, _082361_, _085186_);
  and g_140841_(_082359_, _085186_, _085187_);
  xor g_140842_(_085184_, _085187_, _085188_);
  xor g_140843_(_085185_, _085187_, _085189_);
  or g_140844_(_084139_, _085189_, _085191_);
  not g_140845_(_085191_, _085192_);
  xor g_140846_(_084139_, _085188_, _085193_);
  not g_140847_(_085193_, _085194_);
  and g_140848_(_082366_, _082368_, _085195_);
  xor g_140849_(_085193_, _085195_, _085196_);
  xor g_140850_(_085194_, _085195_, _085197_);
  xor g_140851_(_082376_, _085196_, _085198_);
  not g_140852_(_085198_, _085199_);
  or g_140853_(_084138_, _085198_, _085200_);
  xor g_140854_(_084138_, _085199_, _085202_);
  or g_140855_(_084137_, _085202_, _085203_);
  xor g_140856_(_084136_, _085202_, _085204_);
  and g_140857_(_082383_, _082387_, _085205_);
  not g_140858_(_085205_, _085206_);
  or g_140859_(_085204_, _085205_, _085207_);
  xor g_140860_(_085204_, _085206_, _085208_);
  or g_140861_(_082389_, _085208_, _085209_);
  xor g_140862_(_082390_, _085208_, _085210_);
  and g_140863_(_082392_, _082400_, _085211_);
  not g_140864_(_085211_, _085213_);
  xor g_140865_(_085210_, _085213_, _085214_);
  or g_140866_(_082394_, _085214_, _085215_);
  xor g_140867_(_082394_, _085214_, _085216_);
  xor g_140868_(_082395_, _085214_, _085217_);
  or g_140869_(_082404_, _085217_, _085218_);
  xor g_140870_(_082404_, _085216_, _085219_);
  and g_140871_(_082405_, _082409_, _085220_);
  not g_140872_(_085220_, _085221_);
  or g_140873_(_085219_, _085221_, _085222_);
  xor g_140874_(_085219_, _085220_, _085224_);
  or g_140875_(_084133_, _085224_, _085225_);
  xor g_140876_(_084135_, _085224_, _085226_);
  or g_140877_(_084131_, _085226_, _085227_);
  xor g_140878_(_084132_, _085226_, _085228_);
  or g_140879_(_084129_, _085228_, _085229_);
  xor g_140880_(_084130_, _085228_, _085230_);
  or g_140881_(_082414_, _085230_, _085231_);
  xor g_140882_(_082415_, _085230_, _085232_);
  or g_140883_(_082418_, _085232_, _085233_);
  xor g_140884_(_082420_, _085232_, _085235_);
  or g_140885_(_082424_, _085235_, _085236_);
  not g_140886_(_085236_, _085237_);
  and g_140887_(_082422_, _085235_, _085238_);
  and g_140888_(_082424_, _085238_, _085239_);
  or g_140889_(_082422_, _085232_, _085240_);
  not g_140890_(_085240_, _085241_);
  or g_140891_(_085239_, _085241_, _085242_);
  or g_140892_(_085237_, _085242_, _085243_);
  xor g_140893_(_082428_, _085243_, _085244_);
  xor g_140894_(_084128_, _085244_, _085246_);
  or g_140895_(_084125_, _085246_, _085247_);
  xor g_140896_(_084125_, _085246_, _085248_);
  not g_140897_(_085248_, _085249_);
  or g_140898_(_084124_, _085249_, _085250_);
  xor g_140899_(_084124_, _085248_, _085251_);
  or g_140900_(_084121_, _085251_, _085252_);
  not g_140901_(_085252_, _085253_);
  xor g_140902_(_084121_, _085251_, _085254_);
  xor g_140903_(_084122_, _085251_, _085255_);
  and g_140904_(_082440_, _085255_, _085257_);
  and g_140905_(_082444_, _085257_, _085258_);
  and g_140906_(_082445_, _085254_, _085259_);
  or g_140907_(_082444_, _085255_, _085260_);
  and g_140908_(_082442_, _085254_, _085261_);
  or g_140909_(_085259_, _085261_, _085262_);
  or g_140910_(_085258_, _085262_, _085263_);
  or g_140911_(_082448_, _085263_, _085264_);
  xor g_140912_(_082449_, _085263_, _085265_);
  or g_140913_(_082453_, _085265_, _085266_);
  xor g_140914_(_082453_, _085265_, _085268_);
  xor g_140915_(_082454_, _085265_, _085269_);
  or g_140916_(_082457_, _085269_, _085270_);
  xor g_140917_(_082457_, _085269_, _085271_);
  xor g_140918_(_082457_, _085268_, _085272_);
  or g_140919_(_082459_, _085272_, _085273_);
  xor g_140920_(_082459_, _085272_, _085274_);
  xor g_140921_(_082459_, _085271_, _085275_);
  and g_140922_(_082462_, _085275_, _085276_);
  and g_140923_(_082470_, _085276_, _085277_);
  and g_140924_(_082464_, _085271_, _085279_);
  not g_140925_(_085279_, _085280_);
  and g_140926_(_082469_, _085274_, _085281_);
  or g_140927_(_085279_, _085281_, _085282_);
  or g_140928_(_085277_, _085282_, _085283_);
  or g_140929_(_082467_, _085283_, _085284_);
  not g_140930_(_085284_, _085285_);
  xor g_140931_(_082468_, _085283_, _085286_);
  xor g_140932_(_082478_, _085286_, _085287_);
  xor g_140933_(_082481_, _085287_, _085288_);
  xor g_140934_(_082482_, _085287_, _085290_);
  and g_140935_(_082484_, _085290_, _085291_);
  or g_140936_(_082486_, _085288_, _085292_);
  and g_140937_(_084119_, _085291_, _085293_);
  or g_140938_(_084120_, _085292_, _085294_);
  or g_140939_(_082484_, _085287_, _085295_);
  not g_140940_(_085295_, _085296_);
  or g_140941_(_084119_, _085290_, _085297_);
  not g_140942_(_085297_, _085298_);
  and g_140943_(_085295_, _085297_, _085299_);
  not g_140944_(_085299_, _085301_);
  and g_140945_(_085294_, _085299_, _085302_);
  or g_140946_(_085293_, _085301_, _085303_);
  or g_140947_(_084118_, _085303_, _085304_);
  xor g_140948_(_084118_, _085302_, _085305_);
  or g_140949_(_082501_, _085305_, _085306_);
  not g_140950_(_085306_, _085307_);
  xor g_140951_(_082500_, _085305_, _085308_);
  or g_140952_(_082499_, _085308_, _085309_);
  xor g_140953_(_082499_, _085308_, _085310_);
  xor g_140954_(_082498_, _085308_, _085312_);
  and g_140955_(_082504_, _082506_, _085313_);
  or g_140956_(_085312_, _085313_, _085314_);
  xor g_140957_(_085312_, _085313_, _085315_);
  xor g_140958_(_085310_, _085313_, _085316_);
  and g_140959_(_082513_, _085315_, _085317_);
  not g_140960_(_085317_, _085318_);
  and g_140961_(_082510_, _085315_, _085319_);
  not g_140962_(_085319_, _085320_);
  and g_140963_(_085318_, _085320_, _085321_);
  or g_140964_(_085317_, _085319_, _085323_);
  and g_140965_(_082511_, _085316_, _085324_);
  and g_140966_(_082514_, _085324_, _085325_);
  or g_140967_(_085323_, _085325_, _085326_);
  or g_140968_(_082521_, _085326_, _085327_);
  not g_140969_(_085327_, _085328_);
  xor g_140970_(_082520_, _085326_, _085329_);
  or g_140971_(_082523_, _085329_, _085330_);
  not g_140972_(_085330_, _085331_);
  xor g_140973_(_082523_, _085329_, _085332_);
  xor g_140974_(_082522_, _085329_, _085334_);
  and g_140975_(_082532_, _085332_, _085335_);
  or g_140976_(_082533_, _085334_, _085336_);
  and g_140977_(_082527_, _085332_, _085337_);
  or g_140978_(_082528_, _085334_, _085338_);
  and g_140979_(_085336_, _085338_, _085339_);
  or g_140980_(_085335_, _085337_, _085340_);
  and g_140981_(_082528_, _085334_, _085341_);
  or g_140982_(_082527_, _085332_, _085342_);
  and g_140983_(_082533_, _085341_, _085343_);
  or g_140984_(_082532_, _085342_, _085345_);
  and g_140985_(_085339_, _085345_, _085346_);
  or g_140986_(_085340_, _085343_, _085347_);
  and g_140987_(_082535_, _085347_, _085348_);
  and g_140988_(_084116_, _085348_, _085349_);
  and g_140989_(_084117_, _085346_, _085350_);
  or g_140990_(_084116_, _085347_, _085351_);
  and g_140991_(_082536_, _085346_, _085352_);
  or g_140992_(_082535_, _085347_, _085353_);
  or g_140993_(_085350_, _085352_, _085354_);
  or g_140994_(_085349_, _085354_, _085356_);
  not g_140995_(_085356_, _085357_);
  and g_140996_(_084114_, _085357_, _085358_);
  or g_140997_(_084115_, _085356_, _085359_);
  xor g_140998_(_084114_, _085356_, _085360_);
  or g_140999_(_082542_, _085360_, _085361_);
  not g_141000_(_085361_, _085362_);
  xor g_141001_(_082543_, _085360_, _085363_);
  not g_141002_(_085363_, _085364_);
  or g_141003_(_079589_, _082548_, _085365_);
  or g_141004_(_085363_, _085365_, _085367_);
  not g_141005_(_085367_, _085368_);
  and g_141006_(_082546_, _085363_, _085369_);
  and g_141007_(_085365_, _085369_, _085370_);
  and g_141008_(_082547_, _085364_, _085371_);
  or g_141009_(_085370_, _085371_, _085372_);
  or g_141010_(_085368_, _085372_, _085373_);
  or g_141011_(_079599_, _082549_, _085374_);
  or g_141012_(_079591_, _082548_, _085375_);
  and g_141013_(_085374_, _085375_, _085376_);
  xor g_141014_(_085373_, _085376_, _085378_);
  not g_141015_(_085378_, _085379_);
  and g_141016_(_084113_, _085378_, _085380_);
  or g_141017_(_084111_, _085379_, _085381_);
  xor g_141018_(_084111_, _085378_, _085382_);
  or g_141019_(_082558_, _085382_, _085383_);
  xor g_141020_(_082558_, _085382_, _085384_);
  xor g_141021_(_082563_, _085384_, _085385_);
  not g_141022_(_085385_, _085386_);
  and g_141023_(_082566_, _085385_, _085387_);
  or g_141024_(_082567_, _085386_, _085389_);
  xor g_141025_(_082566_, _085385_, _085390_);
  xor g_141026_(_082567_, _085385_, _085391_);
  and g_141027_(_082570_, _085390_, _085392_);
  or g_141028_(_082569_, _085391_, _085393_);
  xor g_141029_(_082570_, _085390_, _085394_);
  xor g_141030_(_082569_, _085390_, _085395_);
  and g_141031_(_082575_, _085395_, _085396_);
  or g_141032_(_082574_, _085394_, _085397_);
  and g_141033_(_084109_, _085396_, _085398_);
  or g_141034_(_084110_, _085397_, _085400_);
  and g_141035_(_082574_, _085394_, _085401_);
  or g_141036_(_082575_, _085395_, _085402_);
  and g_141037_(_084110_, _085394_, _085403_);
  or g_141038_(_084109_, _085395_, _085404_);
  and g_141039_(_085402_, _085404_, _085405_);
  or g_141040_(_085401_, _085403_, _085406_);
  and g_141041_(_085400_, _085405_, _085407_);
  or g_141042_(_085398_, _085406_, _085408_);
  or g_141043_(_084108_, _085408_, _085409_);
  xor g_141044_(_084108_, _085407_, _085411_);
  or g_141045_(_082585_, _085411_, _085412_);
  xor g_141046_(_082586_, _085411_, _085413_);
  or g_141047_(_084107_, _085413_, _085414_);
  not g_141048_(_085414_, _085415_);
  xor g_141049_(_084107_, _085413_, _085416_);
  not g_141050_(_085416_, _085417_);
  or g_141051_(_084106_, _085417_, _085418_);
  xor g_141052_(_084106_, _085416_, _085419_);
  and g_141053_(_082592_, _085419_, _085420_);
  or g_141054_(_082592_, _085419_, _085422_);
  not g_141055_(_085422_, _085423_);
  xor g_141056_(_082592_, _085419_, _085424_);
  or g_141057_(_085420_, _085423_, _085425_);
  or g_141058_(_084105_, _085425_, _085426_);
  xor g_141059_(_084105_, _085424_, _085427_);
  or g_141060_(_084104_, _085427_, _085428_);
  xor g_141061_(_084104_, _085427_, _085429_);
  not g_141062_(_085429_, _085430_);
  or g_141063_(_079643_, _082603_, _085431_);
  and g_141064_(_082600_, _085431_, _085433_);
  xor g_141065_(_085429_, _085433_, _085434_);
  xor g_141066_(_084102_, _085434_, _085435_);
  xor g_141067_(_084103_, _085434_, _085436_);
  and g_141068_(_082611_, _085436_, _085437_);
  and g_141069_(_082613_, _085437_, _085438_);
  and g_141070_(_082614_, _085435_, _085439_);
  not g_141071_(_085439_, _085440_);
  and g_141072_(_082610_, _085435_, _085441_);
  or g_141073_(_085439_, _085441_, _085442_);
  or g_141074_(_085438_, _085442_, _085444_);
  or g_141075_(_082616_, _085444_, _085445_);
  xor g_141076_(_082618_, _085444_, _085446_);
  and g_141077_(_082621_, _082623_, _085447_);
  xor g_141078_(_085446_, _085447_, _085448_);
  not g_141079_(_085448_, _085449_);
  xor g_141080_(_084099_, _085448_, _085450_);
  not g_141081_(_085450_, _085451_);
  and g_141082_(_084096_, _085451_, _085452_);
  or g_141083_(_084097_, _085450_, _085453_);
  xor g_141084_(_084096_, _085450_, _085455_);
  not g_141085_(_085455_, _085456_);
  or g_141086_(_082632_, _085455_, _085457_);
  xor g_141087_(_082632_, _085455_, _085458_);
  xor g_141088_(_082632_, _085456_, _085459_);
  or g_141089_(_082637_, _085459_, _085460_);
  not g_141090_(_085460_, _085461_);
  and g_141091_(_082635_, _085459_, _085462_);
  or g_141092_(_082634_, _085458_, _085463_);
  and g_141093_(_082637_, _085462_, _085464_);
  or g_141094_(_082638_, _085463_, _085466_);
  and g_141095_(_082634_, _085456_, _085467_);
  not g_141096_(_085467_, _085468_);
  and g_141097_(_085466_, _085468_, _085469_);
  or g_141098_(_085464_, _085467_, _085470_);
  and g_141099_(_085460_, _085469_, _085471_);
  or g_141100_(_085461_, _085470_, _085472_);
  or g_141101_(_082644_, _085472_, _085473_);
  xor g_141102_(_082644_, _085472_, _085474_);
  xor g_141103_(_082644_, _085471_, _085475_);
  and g_141104_(_076856_, _084093_, _085477_);
  or g_141105_(_076854_, _084094_, _085478_);
  and g_141106_(_082642_, _085478_, _085479_);
  xor g_141107_(_085475_, _085479_, _085480_);
  xor g_141108_(_085474_, _085479_, _085481_);
  or g_141109_(_084095_, _085481_, _085482_);
  not g_141110_(_085482_, _085483_);
  xor g_141111_(_084095_, _085481_, _085484_);
  xor g_141112_(_084095_, _085480_, _085485_);
  or g_141113_(_082654_, _082658_, _085486_);
  or g_141114_(_085484_, _085486_, _085488_);
  or g_141115_(_082659_, _085485_, _085489_);
  not g_141116_(_085489_, _085490_);
  or g_141117_(_082655_, _085485_, _085491_);
  not g_141118_(_085491_, _085492_);
  and g_141119_(_085489_, _085491_, _085493_);
  and g_141120_(_085488_, _085493_, _085494_);
  not g_141121_(_085494_, _085495_);
  or g_141122_(_082665_, _085495_, _085496_);
  not g_141123_(_085496_, _085497_);
  or g_141124_(_082662_, _085495_, _085499_);
  not g_141125_(_085499_, _085500_);
  xor g_141126_(_082662_, _085494_, _085501_);
  or g_141127_(_082668_, _085501_, _085502_);
  not g_141128_(_085502_, _085503_);
  xor g_141129_(_082669_, _085501_, _085504_);
  and g_141130_(_082665_, _085504_, _085505_);
  or g_141131_(_085497_, _085505_, _085506_);
  or g_141132_(_082671_, _085506_, _085507_);
  xor g_141133_(_082671_, _085506_, _085508_);
  xor g_141134_(_082673_, _085506_, _085510_);
  and g_141135_(_082680_, _085510_, _085511_);
  or g_141136_(_082681_, _085508_, _085512_);
  and g_141137_(_082676_, _085508_, _085513_);
  or g_141138_(_082677_, _085510_, _085514_);
  or g_141139_(_082678_, _085506_, _085515_);
  not g_141140_(_085515_, _085516_);
  and g_141141_(_085514_, _085515_, _085517_);
  or g_141142_(_085513_, _085516_, _085518_);
  and g_141143_(_085512_, _085517_, _085519_);
  or g_141144_(_085511_, _085518_, _085521_);
  or g_141145_(_082693_, _085521_, _085522_);
  or g_141146_(_082690_, _085521_, _085523_);
  not g_141147_(_085523_, _085524_);
  and g_141148_(_085522_, _085523_, _085525_);
  not g_141149_(_085525_, _085526_);
  and g_141150_(_082690_, _085521_, _085527_);
  or g_141151_(_082689_, _085519_, _085528_);
  and g_141152_(_082693_, _085527_, _085529_);
  or g_141153_(_082695_, _085528_, _085530_);
  and g_141154_(_085525_, _085530_, _085532_);
  or g_141155_(_085526_, _085529_, _085533_);
  or g_141156_(_084092_, _085533_, _085534_);
  xor g_141157_(_084092_, _085532_, _085535_);
  or g_141158_(_084089_, _085535_, _085536_);
  xor g_141159_(_084091_, _085535_, _085537_);
  or g_141160_(_082707_, _085537_, _085538_);
  xor g_141161_(_082706_, _085537_, _085539_);
  or g_141162_(_082702_, _085539_, _085540_);
  xor g_141163_(_082701_, _085539_, _085541_);
  not g_141164_(_085541_, _085543_);
  and g_141165_(_082710_, _082712_, _085544_);
  xor g_141166_(_085541_, _085544_, _085545_);
  xor g_141167_(_085543_, _085544_, _085546_);
  or g_141168_(_082715_, _085546_, _085547_);
  xor g_141169_(_082715_, _085545_, _085548_);
  or g_141170_(_082719_, _085548_, _085549_);
  xor g_141171_(_082719_, _085548_, _085550_);
  not g_141172_(_085550_, _085551_);
  or g_141173_(_082721_, _085551_, _085552_);
  not g_141174_(_085552_, _085554_);
  xor g_141175_(_082721_, _085550_, _085555_);
  or g_141176_(_082724_, _085555_, _085556_);
  xor g_141177_(_082725_, _085555_, _085557_);
  or g_141178_(_079755_, _082731_, _085558_);
  and g_141179_(_082729_, _085558_, _085559_);
  not g_141180_(_085559_, _085560_);
  xor g_141181_(_085557_, _085560_, _085561_);
  or g_141182_(_084088_, _085561_, _085562_);
  not g_141183_(_085562_, _085563_);
  xor g_141184_(_084088_, _085561_, _085565_);
  not g_141185_(_085565_, _085566_);
  and g_141186_(_082735_, _085565_, _085567_);
  or g_141187_(_082734_, _085566_, _085568_);
  xor g_141188_(_082734_, _085565_, _085569_);
  not g_141189_(_085569_, _085570_);
  and g_141190_(_082739_, _085570_, _085571_);
  or g_141191_(_082740_, _085569_, _085572_);
  xor g_141192_(_082740_, _085569_, _085573_);
  not g_141193_(_085573_, _085574_);
  and g_141194_(_082742_, _082748_, _085576_);
  xor g_141195_(_085573_, _085576_, _085577_);
  or g_141196_(_082744_, _085577_, _085578_);
  xor g_141197_(_082745_, _085577_, _085579_);
  or g_141198_(_082754_, _085579_, _085580_);
  xor g_141199_(_082755_, _085579_, _085581_);
  or g_141200_(_084087_, _085581_, _085582_);
  not g_141201_(_085582_, _085583_);
  and g_141202_(_084087_, _085581_, _085584_);
  xor g_141203_(_084087_, _085581_, _085585_);
  or g_141204_(_085583_, _085584_, _085587_);
  or g_141205_(_084086_, _085587_, _085588_);
  xor g_141206_(_084086_, _085585_, _085589_);
  not g_141207_(_085589_, _085590_);
  or g_141208_(_082759_, _085589_, _085591_);
  not g_141209_(_085591_, _085592_);
  and g_141210_(_082765_, _085590_, _085593_);
  not g_141211_(_085593_, _085594_);
  xor g_141212_(_082766_, _085589_, _085595_);
  xor g_141213_(_082765_, _085589_, _085596_);
  and g_141214_(_082759_, _085596_, _085598_);
  or g_141215_(_082761_, _085595_, _085599_);
  and g_141216_(_085591_, _085599_, _085600_);
  or g_141217_(_085592_, _085598_, _085601_);
  and g_141218_(_082769_, _082772_, _085602_);
  xor g_141219_(_085600_, _085602_, _085603_);
  xor g_141220_(_082776_, _085603_, _085604_);
  xor g_141221_(_082777_, _085603_, _085605_);
  and g_141222_(_082779_, _085605_, _085606_);
  and g_141223_(_082784_, _085606_, _085607_);
  and g_141224_(_082783_, _085604_, _085609_);
  or g_141225_(_082784_, _085605_, _085610_);
  or g_141226_(_082779_, _085603_, _085611_);
  not g_141227_(_085611_, _085612_);
  or g_141228_(_085609_, _085612_, _085613_);
  or g_141229_(_085607_, _085613_, _085614_);
  or g_141230_(_084085_, _085614_, _085615_);
  not g_141231_(_085615_, _085616_);
  xor g_141232_(_084084_, _085614_, _085617_);
  not g_141233_(_085617_, _085618_);
  and g_141234_(_084083_, _085618_, _085620_);
  not g_141235_(_085620_, _085621_);
  xor g_141236_(_084083_, _085617_, _085622_);
  and g_141237_(_082790_, _082796_, _085623_);
  not g_141238_(_085623_, _085624_);
  or g_141239_(_085622_, _085623_, _085625_);
  not g_141240_(_085625_, _085626_);
  xor g_141241_(_085622_, _085624_, _085627_);
  or g_141242_(_082794_, _085627_, _085628_);
  xor g_141243_(_082795_, _085627_, _085629_);
  not g_141244_(_085629_, _085631_);
  or g_141245_(_079818_, _082798_, _085632_);
  or g_141246_(_085629_, _085632_, _085633_);
  xor g_141247_(_085629_, _085632_, _085634_);
  xor g_141248_(_085631_, _085632_, _085635_);
  or g_141249_(_084082_, _085635_, _085636_);
  xor g_141250_(_084082_, _085634_, _085637_);
  xor g_141251_(_082810_, _085637_, _085638_);
  or g_141252_(_084080_, _085638_, _085639_);
  xor g_141253_(_084080_, _085638_, _085640_);
  xor g_141254_(_084081_, _085638_, _085642_);
  or g_141255_(_079833_, _082811_, _085643_);
  not g_141256_(_085643_, _085644_);
  and g_141257_(_085642_, _085643_, _085645_);
  or g_141258_(_085640_, _085644_, _085646_);
  and g_141259_(_084078_, _085645_, _085647_);
  or g_141260_(_084077_, _085646_, _085648_);
  or g_141261_(_084078_, _085642_, _085649_);
  not g_141262_(_085649_, _085650_);
  or g_141263_(_085642_, _085643_, _085651_);
  and g_141264_(_085649_, _085651_, _085653_);
  not g_141265_(_085653_, _085654_);
  and g_141266_(_085648_, _085653_, _085655_);
  or g_141267_(_085647_, _085654_, _085656_);
  or g_141268_(_084076_, _085656_, _085657_);
  xor g_141269_(_084076_, _085655_, _085658_);
  or g_141270_(_084075_, _085658_, _085659_);
  not g_141271_(_085659_, _085660_);
  xor g_141272_(_084074_, _085658_, _085661_);
  and g_141273_(_082818_, _082821_, _085662_);
  or g_141274_(_082819_, _082820_, _085664_);
  and g_141275_(_082829_, _085664_, _085665_);
  or g_141276_(_085661_, _085665_, _085666_);
  not g_141277_(_085666_, _085667_);
  xor g_141278_(_085661_, _085665_, _085668_);
  not g_141279_(_085668_, _085669_);
  or g_141280_(_082827_, _085669_, _085670_);
  xor g_141281_(_082827_, _085668_, _085671_);
  and g_141282_(_081064_, _082830_, _085672_);
  or g_141283_(_081063_, _082831_, _085673_);
  or g_141284_(_085671_, _085673_, _085675_);
  xor g_141285_(_085671_, _085672_, _085676_);
  or g_141286_(_082836_, _085676_, _085677_);
  not g_141287_(_085677_, _085678_);
  and g_141288_(_082836_, _085676_, _085679_);
  xor g_141289_(_082836_, _085676_, _085680_);
  or g_141290_(_085678_, _085679_, _085681_);
  or g_141291_(_081061_, _082834_, _085682_);
  or g_141292_(_085681_, _085682_, _085683_);
  xor g_141293_(_085680_, _085682_, _085684_);
  or g_141294_(_082840_, _085684_, _085686_);
  not g_141295_(_085686_, _085687_);
  or g_141296_(_082845_, _085684_, _085688_);
  xor g_141297_(_082845_, _085684_, _085689_);
  xor g_141298_(_082844_, _085684_, _085690_);
  and g_141299_(_082840_, _085690_, _085691_);
  or g_141300_(_082841_, _085689_, _085692_);
  and g_141301_(_085686_, _085692_, _085693_);
  or g_141302_(_085687_, _085691_, _085694_);
  and g_141303_(_082849_, _085693_, _085695_);
  or g_141304_(_082847_, _085694_, _085697_);
  and g_141305_(_082852_, _085693_, _085698_);
  xor g_141306_(_082851_, _085693_, _085699_);
  and g_141307_(_082847_, _085699_, _085700_);
  or g_141308_(_085695_, _085700_, _085701_);
  or g_141309_(_082855_, _085701_, _085702_);
  xor g_141310_(_082856_, _085701_, _085703_);
  or g_141311_(_084073_, _085703_, _085704_);
  not g_141312_(_085704_, _085705_);
  xor g_141313_(_084073_, _085703_, _085706_);
  not g_141314_(_085706_, _085708_);
  or g_141315_(_084072_, _085708_, _085709_);
  not g_141316_(_085709_, _085710_);
  xor g_141317_(_084072_, _085706_, _085711_);
  and g_141318_(_082864_, _082867_, _085712_);
  or g_141319_(_085711_, _085712_, _085713_);
  not g_141320_(_085713_, _085714_);
  and g_141321_(_085711_, _085712_, _085715_);
  xor g_141322_(_085711_, _085712_, _085716_);
  or g_141323_(_085714_, _085715_, _085717_);
  or g_141324_(_082874_, _085717_, _085719_);
  not g_141325_(_085719_, _085720_);
  xor g_141326_(_082874_, _085716_, _085721_);
  or g_141327_(_082872_, _085721_, _085722_);
  not g_141328_(_085722_, _085723_);
  xor g_141329_(_082873_, _085721_, _085724_);
  or g_141330_(_082878_, _085724_, _085725_);
  not g_141331_(_085725_, _085726_);
  and g_141332_(_082880_, _085724_, _085727_);
  and g_141333_(_082878_, _085727_, _085728_);
  or g_141334_(_082880_, _085724_, _085730_);
  not g_141335_(_085730_, _085731_);
  or g_141336_(_085728_, _085731_, _085732_);
  or g_141337_(_085726_, _085732_, _085733_);
  or g_141338_(_082884_, _085733_, _085734_);
  xor g_141339_(_082884_, _085733_, _085735_);
  not g_141340_(_085735_, _085736_);
  or g_141341_(_082890_, _085736_, _085737_);
  xor g_141342_(_082889_, _085735_, _085738_);
  xor g_141343_(_082890_, _085735_, _085739_);
  and g_141344_(_084071_, _085738_, _085741_);
  or g_141345_(_084070_, _085739_, _085742_);
  xor g_141346_(_084070_, _085738_, _085743_);
  or g_141347_(_084067_, _085743_, _085744_);
  not g_141348_(_085744_, _085745_);
  xor g_141349_(_084069_, _085743_, _085746_);
  not g_141350_(_085746_, _085747_);
  and g_141351_(_082897_, _082900_, _085748_);
  xor g_141352_(_085746_, _085748_, _085749_);
  xor g_141353_(_085747_, _085748_, _085750_);
  and g_141354_(_082902_, _082906_, _085752_);
  xor g_141355_(_085749_, _085752_, _085753_);
  xor g_141356_(_082910_, _085753_, _085754_);
  xor g_141357_(_082911_, _085753_, _085755_);
  or g_141358_(_084066_, _085755_, _085756_);
  not g_141359_(_085756_, _085757_);
  xor g_141360_(_084066_, _085754_, _085758_);
  or g_141361_(_084064_, _085758_, _085759_);
  xor g_141362_(_084065_, _085758_, _085760_);
  or g_141363_(_079915_, _082920_, _085761_);
  and g_141364_(_082919_, _085761_, _085763_);
  or g_141365_(_085760_, _085763_, _085764_);
  xor g_141366_(_085760_, _085763_, _085765_);
  not g_141367_(_085765_, _085766_);
  and g_141368_(_084063_, _085765_, _085767_);
  or g_141369_(_084062_, _085766_, _085768_);
  xor g_141370_(_084063_, _085765_, _085769_);
  xor g_141371_(_084062_, _085765_, _085770_);
  and g_141372_(_082924_, _085770_, _085771_);
  and g_141373_(_082930_, _085771_, _085772_);
  and g_141374_(_082929_, _085769_, _085774_);
  or g_141375_(_082930_, _085770_, _085775_);
  and g_141376_(_082926_, _085765_, _085776_);
  not g_141377_(_085776_, _085777_);
  or g_141378_(_085774_, _085776_, _085778_);
  or g_141379_(_085772_, _085778_, _085779_);
  or g_141380_(_084060_, _085779_, _085780_);
  xor g_141381_(_084060_, _085779_, _085781_);
  xor g_141382_(_084061_, _085779_, _085782_);
  and g_141383_(_082933_, _085782_, _085783_);
  and g_141384_(_084059_, _085783_, _085785_);
  and g_141385_(_084058_, _085781_, _085786_);
  or g_141386_(_084059_, _085782_, _085787_);
  and g_141387_(_082934_, _085781_, _085788_);
  or g_141388_(_082933_, _085782_, _085789_);
  or g_141389_(_085786_, _085788_, _085790_);
  or g_141390_(_085785_, _085790_, _085791_);
  or g_141391_(_084055_, _085791_, _085792_);
  xor g_141392_(_084056_, _085791_, _085793_);
  or g_141393_(_082939_, _085793_, _085794_);
  xor g_141394_(_082940_, _085793_, _085796_);
  and g_141395_(_082944_, _082948_, _085797_);
  not g_141396_(_085797_, _085798_);
  xor g_141397_(_085796_, _085797_, _085799_);
  xor g_141398_(_085796_, _085798_, _085800_);
  or g_141399_(_079946_, _082945_, _085801_);
  or g_141400_(_085800_, _085801_, _085802_);
  not g_141401_(_085802_, _085803_);
  or g_141402_(_082955_, _085799_, _085804_);
  and g_141403_(_085802_, _085804_, _085805_);
  and g_141404_(_082951_, _085805_, _085807_);
  not g_141405_(_085807_, _085808_);
  xor g_141406_(_082951_, _085805_, _085809_);
  xor g_141407_(_082950_, _085805_, _085810_);
  or g_141408_(_084052_, _085810_, _085811_);
  xor g_141409_(_084052_, _085809_, _085812_);
  or g_141410_(_084050_, _085812_, _085813_);
  not g_141411_(_085813_, _085814_);
  xor g_141412_(_084051_, _085812_, _085815_);
  not g_141413_(_085815_, _085816_);
  and g_141414_(_082967_, _085816_, _085818_);
  not g_141415_(_085818_, _085819_);
  and g_141416_(_082962_, _085815_, _085820_);
  and g_141417_(_082966_, _085820_, _085821_);
  and g_141418_(_082963_, _085816_, _085822_);
  not g_141419_(_085822_, _085823_);
  or g_141420_(_085821_, _085822_, _085824_);
  or g_141421_(_085818_, _085824_, _085825_);
  and g_141422_(_082970_, _082973_, _085826_);
  and g_141423_(_085825_, _085826_, _085827_);
  or g_141424_(_085825_, _085826_, _085829_);
  not g_141425_(_085829_, _085830_);
  xor g_141426_(_085825_, _085826_, _085831_);
  or g_141427_(_085827_, _085830_, _085832_);
  or g_141428_(_082976_, _085832_, _085833_);
  xor g_141429_(_082976_, _085831_, _085834_);
  xor g_141430_(_082983_, _085834_, _085835_);
  xor g_141431_(_084049_, _085835_, _085836_);
  not g_141432_(_085836_, _085837_);
  or g_141433_(_082993_, _085837_, _085838_);
  xor g_141434_(_082994_, _085836_, _085840_);
  xor g_141435_(_082993_, _085836_, _085841_);
  or g_141436_(_082999_, _085841_, _085842_);
  xor g_141437_(_082999_, _085840_, _085843_);
  or g_141438_(_083007_, _085843_, _085844_);
  not g_141439_(_085844_, _085845_);
  and g_141440_(_083001_, _085843_, _085846_);
  and g_141441_(_083007_, _085846_, _085847_);
  or g_141442_(_083001_, _085843_, _085848_);
  not g_141443_(_085848_, _085849_);
  or g_141444_(_085847_, _085849_, _085851_);
  or g_141445_(_085845_, _085851_, _085852_);
  or g_141446_(_083010_, _085852_, _085853_);
  not g_141447_(_085853_, _085854_);
  xor g_141448_(_083010_, _085852_, _085855_);
  xor g_141449_(_083011_, _085852_, _085856_);
  or g_141450_(_083016_, _085855_, _085857_);
  or g_141451_(_083019_, _085857_, _085858_);
  or g_141452_(_083020_, _085856_, _085859_);
  or g_141453_(_083015_, _085852_, _085860_);
  not g_141454_(_085860_, _085862_);
  and g_141455_(_085859_, _085860_, _085863_);
  and g_141456_(_085858_, _085863_, _085864_);
  not g_141457_(_085864_, _085865_);
  or g_141458_(_080007_, _083023_, _085866_);
  not g_141459_(_085866_, _085867_);
  and g_141460_(_083022_, _085866_, _085868_);
  not g_141461_(_085868_, _085869_);
  xor g_141462_(_085864_, _085869_, _085870_);
  xor g_141463_(_085864_, _085868_, _085871_);
  or g_141464_(_080010_, _083023_, _085873_);
  not g_141465_(_085873_, _085874_);
  and g_141466_(_085871_, _085873_, _085875_);
  and g_141467_(_083028_, _085875_, _085876_);
  and g_141468_(_083029_, _085870_, _085877_);
  and g_141469_(_085870_, _085874_, _085878_);
  not g_141470_(_085878_, _085879_);
  or g_141471_(_085877_, _085878_, _085880_);
  or g_141472_(_085876_, _085880_, _085881_);
  or g_141473_(_083033_, _085881_, _085882_);
  xor g_141474_(_083034_, _085881_, _085884_);
  or g_141475_(_083038_, _085884_, _085885_);
  xor g_141476_(_083039_, _085884_, _085886_);
  or g_141477_(_084047_, _085886_, _085887_);
  xor g_141478_(_084048_, _085886_, _085888_);
  or g_141479_(_084044_, _085888_, _085889_);
  xor g_141480_(_084045_, _085888_, _085890_);
  not g_141481_(_085890_, _085891_);
  or g_141482_(_080032_, _083045_, _085892_);
  not g_141483_(_085892_, _085893_);
  and g_141484_(_083044_, _085892_, _085895_);
  xor g_141485_(_085890_, _085895_, _085896_);
  and g_141486_(_084043_, _085896_, _085897_);
  not g_141487_(_085897_, _085898_);
  xor g_141488_(_084043_, _085896_, _085899_);
  xor g_141489_(_084042_, _085896_, _085900_);
  and g_141490_(_083051_, _083054_, _085901_);
  xor g_141491_(_085899_, _085901_, _085902_);
  or g_141492_(_083056_, _085902_, _085903_);
  not g_141493_(_085903_, _085904_);
  xor g_141494_(_083056_, _085902_, _085906_);
  xor g_141495_(_083058_, _085902_, _085907_);
  and g_141496_(_083062_, _085907_, _085908_);
  or g_141497_(_083061_, _085906_, _085909_);
  and g_141498_(_084040_, _085908_, _085910_);
  or g_141499_(_084041_, _085909_, _085911_);
  or g_141500_(_084040_, _085907_, _085912_);
  or g_141501_(_083062_, _085902_, _085913_);
  not g_141502_(_085913_, _085914_);
  and g_141503_(_085912_, _085913_, _085915_);
  not g_141504_(_085915_, _085917_);
  and g_141505_(_085911_, _085915_, _085918_);
  or g_141506_(_085910_, _085917_, _085919_);
  or g_141507_(_084039_, _085919_, _085920_);
  xor g_141508_(_084039_, _085918_, _085921_);
  or g_141509_(_084037_, _085921_, _085922_);
  xor g_141510_(_084038_, _085921_, _085923_);
  or g_141511_(_081040_, _083067_, _085924_);
  and g_141512_(_083070_, _085924_, _085925_);
  not g_141513_(_085925_, _085926_);
  xor g_141514_(_085923_, _085926_, _085928_);
  not g_141515_(_085928_, _085929_);
  xor g_141516_(_084036_, _085928_, _085930_);
  and g_141517_(_084032_, _085930_, _085931_);
  xor g_141518_(_084031_, _085930_, _085932_);
  or g_141519_(_084030_, _085932_, _085933_);
  not g_141520_(_085933_, _085934_);
  xor g_141521_(_084030_, _085932_, _085935_);
  not g_141522_(_085935_, _085936_);
  and g_141523_(_084029_, _085935_, _085937_);
  or g_141524_(_084028_, _085936_, _085939_);
  xor g_141525_(_084028_, _085935_, _085940_);
  or g_141526_(_083081_, _085940_, _085941_);
  xor g_141527_(_083082_, _085940_, _085942_);
  or g_141528_(_077272_, _084025_, _085943_);
  not g_141529_(_085943_, _085944_);
  or g_141530_(_085942_, _085943_, _085945_);
  xor g_141531_(_085942_, _085944_, _085946_);
  or g_141532_(_084026_, _085946_, _085947_);
  xor g_141533_(_084027_, _085946_, _085948_);
  or g_141534_(_083086_, _085948_, _085950_);
  not g_141535_(_085950_, _085951_);
  xor g_141536_(_083087_, _085948_, _085952_);
  not g_141537_(_085952_, _085953_);
  and g_141538_(_083089_, _083092_, _085954_);
  xor g_141539_(_085952_, _085954_, _085955_);
  xor g_141540_(_085953_, _085954_, _085956_);
  or g_141541_(_084023_, _085956_, _085957_);
  not g_141542_(_085957_, _085958_);
  and g_141543_(_080085_, _083093_, _085959_);
  or g_141544_(_080084_, _083094_, _085961_);
  and g_141545_(_085956_, _085961_, _085962_);
  or g_141546_(_085955_, _085959_, _085963_);
  and g_141547_(_084023_, _085962_, _085964_);
  or g_141548_(_084022_, _085963_, _085965_);
  or g_141549_(_085956_, _085961_, _085966_);
  not g_141550_(_085966_, _085967_);
  and g_141551_(_085965_, _085966_, _085968_);
  or g_141552_(_085964_, _085967_, _085969_);
  and g_141553_(_085957_, _085968_, _085970_);
  or g_141554_(_085958_, _085969_, _085972_);
  or g_141555_(_084021_, _085972_, _085973_);
  xor g_141556_(_084021_, _085972_, _085974_);
  xor g_141557_(_084021_, _085970_, _085975_);
  xor g_141558_(_083097_, _085974_, _085976_);
  not g_141559_(_085976_, _085977_);
  and g_141560_(_084018_, _085977_, _085978_);
  not g_141561_(_085978_, _085979_);
  xor g_141562_(_084018_, _085976_, _085980_);
  or g_141563_(_084017_, _085980_, _085981_);
  not g_141564_(_085981_, _085983_);
  xor g_141565_(_084017_, _085980_, _085984_);
  not g_141566_(_085984_, _085985_);
  or g_141567_(_083102_, _085985_, _085986_);
  not g_141568_(_085986_, _085987_);
  xor g_141569_(_083102_, _085984_, _085988_);
  or g_141570_(_083106_, _085988_, _085989_);
  not g_141571_(_085989_, _085990_);
  xor g_141572_(_083105_, _085988_, _085991_);
  and g_141573_(_083109_, _085991_, _085992_);
  or g_141574_(_083109_, _085991_, _085994_);
  not g_141575_(_085994_, _085995_);
  xor g_141576_(_083109_, _085991_, _085996_);
  or g_141577_(_085992_, _085995_, _085997_);
  or g_141578_(_083113_, _085997_, _085998_);
  not g_141579_(_085998_, _085999_);
  xor g_141580_(_083113_, _085996_, _086000_);
  not g_141581_(_086000_, _086001_);
  and g_141582_(_083117_, _083122_, _086002_);
  xor g_141583_(_086001_, _086002_, _086003_);
  and g_141584_(_083126_, _086003_, _086005_);
  and g_141585_(_084016_, _086005_, _086006_);
  or g_141586_(_084016_, _086003_, _086007_);
  not g_141587_(_086007_, _086008_);
  or g_141588_(_083126_, _086003_, _086009_);
  not g_141589_(_086009_, _086010_);
  and g_141590_(_086007_, _086009_, _086011_);
  not g_141591_(_086011_, _086012_);
  or g_141592_(_086006_, _086012_, _086013_);
  not g_141593_(_086013_, _086014_);
  or g_141594_(_080127_, _083127_, _086016_);
  and g_141595_(_083132_, _086016_, _086017_);
  xor g_141596_(_086014_, _086017_, _086018_);
  xor g_141597_(_086013_, _086017_, _086019_);
  or g_141598_(_084015_, _086018_, _086020_);
  xor g_141599_(_084015_, _086019_, _086021_);
  not g_141600_(_086021_, _086022_);
  or g_141601_(_084014_, _086021_, _086023_);
  xor g_141602_(_084014_, _086021_, _086024_);
  xor g_141603_(_084014_, _086022_, _086025_);
  or g_141604_(_083142_, _083143_, _086027_);
  and g_141605_(_083140_, _086027_, _086028_);
  xor g_141606_(_086024_, _086028_, _086029_);
  or g_141607_(_084012_, _086029_, _086030_);
  xor g_141608_(_084012_, _086029_, _086031_);
  and g_141609_(_083148_, _083151_, _086032_);
  xor g_141610_(_086031_, _086032_, _086033_);
  not g_141611_(_086033_, _086034_);
  and g_141612_(_083158_, _086034_, _086035_);
  xor g_141613_(_083159_, _086033_, _086036_);
  not g_141614_(_086036_, _086038_);
  or g_141615_(_083161_, _086038_, _086039_);
  xor g_141616_(_083162_, _086036_, _086040_);
  xor g_141617_(_083161_, _086036_, _086041_);
  or g_141618_(_080152_, _083163_, _086042_);
  or g_141619_(_083163_, _083165_, _086043_);
  and g_141620_(_086042_, _086043_, _086044_);
  xor g_141621_(_086040_, _086044_, _086045_);
  or g_141622_(_083170_, _086045_, _086046_);
  xor g_141623_(_083170_, _086045_, _086047_);
  not g_141624_(_086047_, _086049_);
  and g_141625_(_083173_, _086047_, _086050_);
  or g_141626_(_083172_, _086049_, _086051_);
  xor g_141627_(_083172_, _086047_, _086052_);
  or g_141628_(_083176_, _086052_, _086053_);
  xor g_141629_(_083175_, _086052_, _086054_);
  or g_141630_(_084011_, _086054_, _086055_);
  xor g_141631_(_084011_, _086054_, _086056_);
  not g_141632_(_086056_, _086057_);
  or g_141633_(_084010_, _086057_, _086058_);
  not g_141634_(_086058_, _086060_);
  xor g_141635_(_084010_, _086056_, _086061_);
  not g_141636_(_086061_, _086062_);
  or g_141637_(_083184_, _086061_, _086063_);
  xor g_141638_(_083184_, _086061_, _086064_);
  xor g_141639_(_083184_, _086062_, _086065_);
  and g_141640_(_083187_, _083191_, _086066_);
  xor g_141641_(_086064_, _086066_, _086067_);
  not g_141642_(_086067_, _086068_);
  or g_141643_(_080177_, _083193_, _086069_);
  and g_141644_(_083194_, _086069_, _086071_);
  xor g_141645_(_086068_, _086071_, _086072_);
  not g_141646_(_086072_, _086073_);
  or g_141647_(_080181_, _083195_, _086074_);
  and g_141648_(_083199_, _086074_, _086075_);
  xor g_141649_(_086072_, _086075_, _086076_);
  xor g_141650_(_086073_, _086075_, _086077_);
  and g_141651_(_083207_, _086076_, _086078_);
  or g_141652_(_083208_, _086077_, _086079_);
  and g_141653_(_083203_, _086076_, _086080_);
  or g_141654_(_083204_, _086077_, _086082_);
  and g_141655_(_086079_, _086082_, _086083_);
  or g_141656_(_086078_, _086080_, _086084_);
  and g_141657_(_083204_, _086077_, _086085_);
  or g_141658_(_083203_, _086076_, _086086_);
  and g_141659_(_083208_, _086085_, _086087_);
  or g_141660_(_083207_, _086086_, _086088_);
  and g_141661_(_086083_, _086088_, _086089_);
  or g_141662_(_086084_, _086087_, _086090_);
  and g_141663_(_083214_, _086089_, _086091_);
  not g_141664_(_086091_, _086093_);
  and g_141665_(_083212_, _086089_, _086094_);
  or g_141666_(_083210_, _086090_, _086095_);
  xor g_141667_(_083210_, _086089_, _086096_);
  or g_141668_(_083216_, _086096_, _086097_);
  not g_141669_(_086097_, _086098_);
  xor g_141670_(_083216_, _086096_, _086099_);
  or g_141671_(_083214_, _086099_, _086100_);
  and g_141672_(_086093_, _086100_, _086101_);
  not g_141673_(_086101_, _086102_);
  and g_141674_(_083220_, _086101_, _086104_);
  not g_141675_(_086104_, _086105_);
  and g_141676_(_083224_, _086101_, _086106_);
  or g_141677_(_083223_, _086102_, _086107_);
  xor g_141678_(_083223_, _086101_, _086108_);
  and g_141679_(_083219_, _086108_, _086109_);
  or g_141680_(_086104_, _086109_, _086110_);
  or g_141681_(_083228_, _086110_, _086111_);
  xor g_141682_(_083227_, _086110_, _086112_);
  not g_141683_(_086112_, _086113_);
  or g_141684_(_083231_, _086112_, _086115_);
  xor g_141685_(_083231_, _086113_, _086116_);
  not g_141686_(_086116_, _086117_);
  or g_141687_(_083235_, _086116_, _086118_);
  xor g_141688_(_083235_, _086117_, _086119_);
  not g_141689_(_086119_, _086120_);
  and g_141690_(_083238_, _083240_, _086121_);
  xor g_141691_(_086119_, _086121_, _086122_);
  not g_141692_(_086122_, _086123_);
  or g_141693_(_084009_, _086123_, _086124_);
  xor g_141694_(_084009_, _086122_, _086126_);
  not g_141695_(_086126_, _086127_);
  or g_141696_(_084008_, _086126_, _086128_);
  xor g_141697_(_084008_, _086127_, _086129_);
  and g_141698_(_083248_, _086129_, _086130_);
  and g_141699_(_083252_, _086130_, _086131_);
  or g_141700_(_083248_, _086129_, _086132_);
  or g_141701_(_083252_, _086129_, _086133_);
  and g_141702_(_086132_, _086133_, _086134_);
  not g_141703_(_086134_, _086135_);
  or g_141704_(_086131_, _086135_, _086137_);
  not g_141705_(_086137_, _086138_);
  xor g_141706_(_084007_, _086138_, _086139_);
  not g_141707_(_086139_, _086140_);
  xor g_141708_(_084006_, _086140_, _086141_);
  or g_141709_(_084004_, _086141_, _086142_);
  xor g_141710_(_084004_, _086141_, _086143_);
  xor g_141711_(_083270_, _086143_, _086144_);
  not g_141712_(_086144_, _086145_);
  and g_141713_(_083272_, _083275_, _086146_);
  xor g_141714_(_086144_, _086146_, _086148_);
  xor g_141715_(_086145_, _086146_, _086149_);
  and g_141716_(_083279_, _086149_, _086150_);
  and g_141717_(_084001_, _086150_, _086151_);
  and g_141718_(_084003_, _086148_, _086152_);
  and g_141719_(_083280_, _086148_, _086153_);
  or g_141720_(_083279_, _086149_, _086154_);
  or g_141721_(_086152_, _086153_, _086155_);
  or g_141722_(_086151_, _086155_, _086156_);
  not g_141723_(_086156_, _086157_);
  or g_141724_(_084000_, _086156_, _086159_);
  not g_141725_(_086159_, _086160_);
  xor g_141726_(_084000_, _086157_, _086161_);
  not g_141727_(_086161_, _086162_);
  and g_141728_(_083286_, _083290_, _086163_);
  xor g_141729_(_086162_, _086163_, _086164_);
  not g_141730_(_086164_, _086165_);
  or g_141731_(_083293_, _086164_, _086166_);
  xor g_141732_(_083293_, _086165_, _086167_);
  not g_141733_(_086167_, _086168_);
  and g_141734_(_083295_, _083298_, _086170_);
  xor g_141735_(_086167_, _086170_, _086171_);
  xor g_141736_(_086168_, _086170_, _086172_);
  and g_141737_(_083301_, _083303_, _086173_);
  xor g_141738_(_086171_, _086173_, _086174_);
  or g_141739_(_083999_, _086174_, _086175_);
  not g_141740_(_086175_, _086176_);
  xor g_141741_(_083999_, _086174_, _086177_);
  not g_141742_(_086177_, _086178_);
  or g_141743_(_083998_, _086178_, _086179_);
  not g_141744_(_086179_, _086181_);
  xor g_141745_(_083998_, _086177_, _086182_);
  and g_141746_(_083307_, _083311_, _086183_);
  and g_141747_(_086182_, _086183_, _086184_);
  not g_141748_(_086184_, _086185_);
  or g_141749_(_083311_, _086182_, _086186_);
  or g_141750_(_083307_, _086182_, _086187_);
  and g_141751_(_086186_, _086187_, _086188_);
  and g_141752_(_086185_, _086188_, _086189_);
  not g_141753_(_086189_, _086190_);
  or g_141754_(_083997_, _086190_, _086192_);
  xor g_141755_(_083997_, _086189_, _086193_);
  not g_141756_(_086193_, _086194_);
  or g_141757_(_083996_, _086193_, _086195_);
  xor g_141758_(_083996_, _086194_, _086196_);
  or g_141759_(_083316_, _086196_, _086197_);
  xor g_141760_(_083317_, _086196_, _086198_);
  and g_141761_(_083320_, _083323_, _086199_);
  not g_141762_(_086199_, _086200_);
  xor g_141763_(_086198_, _086200_, _086201_);
  or g_141764_(_083326_, _086201_, _086203_);
  not g_141765_(_086203_, _086204_);
  xor g_141766_(_083326_, _086201_, _086205_);
  xor g_141767_(_083327_, _086201_, _086206_);
  or g_141768_(_083330_, _086206_, _086207_);
  not g_141769_(_086207_, _086208_);
  xor g_141770_(_083330_, _086205_, _086209_);
  or g_141771_(_080331_, _083336_, _086210_);
  and g_141772_(_083334_, _086210_, _086211_);
  xor g_141773_(_086209_, _086211_, _086212_);
  not g_141774_(_086212_, _086214_);
  or g_141775_(_083995_, _086214_, _086215_);
  xor g_141776_(_083995_, _086212_, _086216_);
  xor g_141777_(_083344_, _086216_, _086217_);
  or g_141778_(_083994_, _086217_, _086218_);
  not g_141779_(_086218_, _086219_);
  xor g_141780_(_083994_, _086217_, _086220_);
  and g_141781_(_083356_, _086220_, _086221_);
  not g_141782_(_086221_, _086222_);
  xor g_141783_(_083356_, _086220_, _086223_);
  not g_141784_(_086223_, _086225_);
  and g_141785_(_083355_, _086223_, _086226_);
  or g_141786_(_083353_, _086225_, _086227_);
  xor g_141787_(_083353_, _086223_, _086228_);
  or g_141788_(_083362_, _086228_, _086229_);
  not g_141789_(_086229_, _086230_);
  and g_141790_(_083362_, _086228_, _086231_);
  xor g_141791_(_083362_, _086228_, _086232_);
  or g_141792_(_086230_, _086231_, _086233_);
  or g_141793_(_083367_, _086233_, _086234_);
  not g_141794_(_086234_, _086236_);
  xor g_141795_(_083367_, _086232_, _086237_);
  not g_141796_(_086237_, _086238_);
  or g_141797_(_083373_, _086237_, _086239_);
  not g_141798_(_086239_, _086240_);
  or g_141799_(_083370_, _086237_, _086241_);
  xor g_141800_(_083370_, _086238_, _086242_);
  not g_141801_(_086242_, _086243_);
  or g_141802_(_083377_, _086242_, _086244_);
  xor g_141803_(_083377_, _086242_, _086245_);
  xor g_141804_(_083377_, _086243_, _086247_);
  and g_141805_(_083373_, _086247_, _086248_);
  or g_141806_(_083374_, _086245_, _086249_);
  and g_141807_(_086239_, _086249_, _086250_);
  or g_141808_(_086240_, _086248_, _086251_);
  or g_141809_(_083993_, _086251_, _086252_);
  xor g_141810_(_083993_, _086250_, _086253_);
  not g_141811_(_086253_, _086254_);
  or g_141812_(_083992_, _086253_, _086255_);
  xor g_141813_(_083992_, _086254_, _086256_);
  and g_141814_(_083382_, _083385_, _086258_);
  xor g_141815_(_086256_, _086258_, _086259_);
  not g_141816_(_086259_, _086260_);
  xor g_141817_(_083990_, _086259_, _086261_);
  or g_141818_(_083393_, _086261_, _086262_);
  xor g_141819_(_083393_, _086261_, _086263_);
  xor g_141820_(_083392_, _086261_, _086264_);
  or g_141821_(_083397_, _086264_, _086265_);
  not g_141822_(_086265_, _086266_);
  xor g_141823_(_083397_, _086263_, _086267_);
  not g_141824_(_086267_, _086269_);
  or g_141825_(_083403_, _086267_, _086270_);
  xor g_141826_(_083403_, _086269_, _086271_);
  not g_141827_(_086271_, _086272_);
  or g_141828_(_080410_, _083406_, _086273_);
  and g_141829_(_083405_, _086273_, _086274_);
  xor g_141830_(_086272_, _086274_, _086275_);
  not g_141831_(_086275_, _086276_);
  and g_141832_(_083412_, _086276_, _086277_);
  not g_141833_(_086277_, _086278_);
  or g_141834_(_080413_, _083406_, _086280_);
  or g_141835_(_086275_, _086280_, _086281_);
  xor g_141836_(_086275_, _086280_, _086282_);
  and g_141837_(_083415_, _086282_, _086283_);
  xor g_141838_(_083416_, _086282_, _086284_);
  and g_141839_(_083411_, _086284_, _086285_);
  or g_141840_(_086277_, _086285_, _086286_);
  not g_141841_(_086286_, _086287_);
  and g_141842_(_083418_, _083422_, _086288_);
  xor g_141843_(_086287_, _086288_, _086289_);
  xor g_141844_(_083989_, _086289_, _086291_);
  not g_141845_(_086291_, _086292_);
  or g_141846_(_083436_, _086291_, _086293_);
  not g_141847_(_086293_, _086294_);
  and g_141848_(_083432_, _086291_, _086295_);
  and g_141849_(_083436_, _086295_, _086296_);
  and g_141850_(_083433_, _086292_, _086297_);
  not g_141851_(_086297_, _086298_);
  or g_141852_(_086296_, _086297_, _086299_);
  or g_141853_(_086294_, _086299_, _086300_);
  not g_141854_(_086300_, _086302_);
  or g_141855_(_080431_, _083440_, _086303_);
  and g_141856_(_083439_, _086303_, _086304_);
  xor g_141857_(_086302_, _086304_, _086305_);
  xor g_141858_(_083987_, _086305_, _086306_);
  and g_141859_(_083985_, _086306_, _086307_);
  not g_141860_(_086307_, _086308_);
  xor g_141861_(_083984_, _086306_, _086309_);
  or g_141862_(_080446_, _083447_, _086310_);
  not g_141863_(_086310_, _086311_);
  or g_141864_(_086309_, _086310_, _086313_);
  xor g_141865_(_086309_, _086311_, _086314_);
  not g_141866_(_086314_, _086315_);
  and g_141867_(_083451_, _083454_, _086316_);
  xor g_141868_(_086315_, _086316_, _086317_);
  not g_141869_(_086317_, _086318_);
  and g_141870_(_083457_, _083460_, _086319_);
  xor g_141871_(_086318_, _086319_, _086320_);
  xor g_141872_(_083982_, _086320_, _086321_);
  xor g_141873_(_083983_, _086320_, _086322_);
  and g_141874_(_083470_, _086322_, _086324_);
  and g_141875_(_083979_, _086324_, _086325_);
  and g_141876_(_083981_, _086321_, _086326_);
  or g_141877_(_083979_, _086322_, _086327_);
  and g_141878_(_083469_, _086321_, _086328_);
  or g_141879_(_086326_, _086328_, _086329_);
  or g_141880_(_086325_, _086329_, _086330_);
  not g_141881_(_086330_, _086331_);
  or g_141882_(_083978_, _086330_, _086332_);
  xor g_141883_(_083978_, _086331_, _086333_);
  or g_141884_(_083476_, _086333_, _086335_);
  not g_141885_(_086335_, _086336_);
  xor g_141886_(_083477_, _086333_, _086337_);
  not g_141887_(_086337_, _086338_);
  or g_141888_(_080482_, _083481_, _086339_);
  and g_141889_(_083480_, _086339_, _086340_);
  xor g_141890_(_086337_, _086340_, _086341_);
  xor g_141891_(_086338_, _086340_, _086342_);
  xor g_141892_(_083977_, _086341_, _086343_);
  or g_141893_(_083490_, _086343_, _086344_);
  not g_141894_(_086344_, _086346_);
  xor g_141895_(_083490_, _086343_, _086347_);
  not g_141896_(_086347_, _086348_);
  or g_141897_(_080488_, _083491_, _086349_);
  or g_141898_(_086348_, _086349_, _086350_);
  xor g_141899_(_086347_, _086349_, _086351_);
  not g_141900_(_086351_, _086352_);
  or g_141901_(_083975_, _086351_, _086353_);
  xor g_141902_(_083975_, _086351_, _086354_);
  xor g_141903_(_083975_, _086352_, _086355_);
  or g_141904_(_083496_, _086355_, _086357_);
  xor g_141905_(_083496_, _086354_, _086358_);
  or g_141906_(_083501_, _086358_, _086359_);
  not g_141907_(_086359_, _086360_);
  or g_141908_(_083499_, _086355_, _086361_);
  not g_141909_(_086361_, _086362_);
  and g_141910_(_083499_, _086358_, _086363_);
  or g_141911_(_086362_, _086363_, _086364_);
  and g_141912_(_083501_, _086364_, _086365_);
  or g_141913_(_086360_, _086365_, _086366_);
  not g_141914_(_086366_, _086368_);
  and g_141915_(_083504_, _083507_, _086369_);
  xor g_141916_(_086366_, _086369_, _086370_);
  xor g_141917_(_086368_, _086369_, _086371_);
  or g_141918_(_083974_, _086371_, _086372_);
  xor g_141919_(_083974_, _086370_, _086373_);
  not g_141920_(_086373_, _086374_);
  or g_141921_(_083973_, _086373_, _086375_);
  xor g_141922_(_083973_, _086374_, _086376_);
  xor g_141923_(_083517_, _086376_, _086377_);
  or g_141924_(_083521_, _086377_, _086379_);
  not g_141925_(_086379_, _086380_);
  and g_141926_(_083521_, _086377_, _086381_);
  xor g_141927_(_083521_, _086377_, _086382_);
  or g_141928_(_086380_, _086381_, _086383_);
  or g_141929_(_083523_, _086383_, _086384_);
  not g_141930_(_086384_, _086385_);
  xor g_141931_(_083523_, _086382_, _086386_);
  or g_141932_(_083525_, _086386_, _086387_);
  xor g_141933_(_083525_, _086386_, _086388_);
  and g_141934_(_083529_, _086388_, _086390_);
  and g_141935_(_083531_, _086386_, _086391_);
  or g_141936_(_086390_, _086391_, _086392_);
  not g_141937_(_086392_, _086393_);
  or g_141938_(_083534_, _086393_, _086394_);
  xor g_141939_(_083534_, _086392_, _086395_);
  not g_141940_(_086395_, _086396_);
  or g_141941_(_083536_, _086395_, _086397_);
  xor g_141942_(_083536_, _086396_, _086398_);
  not g_141943_(_086398_, _086399_);
  and g_141944_(_083540_, _083545_, _086401_);
  xor g_141945_(_086398_, _086401_, _086402_);
  xor g_141946_(_086399_, _086401_, _086403_);
  or g_141947_(_083547_, _086403_, _086404_);
  xor g_141948_(_083547_, _086402_, _086405_);
  not g_141949_(_086405_, _086406_);
  or g_141950_(_083550_, _086405_, _086407_);
  xor g_141951_(_083550_, _086406_, _086408_);
  and g_141952_(_083555_, _086408_, _086409_);
  or g_141953_(_083551_, _086405_, _086410_);
  or g_141954_(_083553_, _086410_, _086412_);
  not g_141955_(_086412_, _086413_);
  or g_141956_(_080551_, _086410_, _086414_);
  not g_141957_(_086414_, _086415_);
  and g_141958_(_086412_, _086414_, _086416_);
  not g_141959_(_086416_, _086417_);
  or g_141960_(_086409_, _086417_, _086418_);
  or g_141961_(_083558_, _086418_, _086419_);
  not g_141962_(_086419_, _086420_);
  xor g_141963_(_083559_, _086418_, _086421_);
  or g_141964_(_083561_, _086421_, _086423_);
  xor g_141965_(_083562_, _086421_, _086424_);
  not g_141966_(_086424_, _086425_);
  and g_141967_(_083564_, _083568_, _086426_);
  xor g_141968_(_086425_, _086426_, _086427_);
  not g_141969_(_086427_, _086428_);
  and g_141970_(_083572_, _083577_, _086429_);
  xor g_141971_(_086428_, _086429_, _086430_);
  or g_141972_(_083972_, _086430_, _086431_);
  xor g_141973_(_083972_, _086430_, _086432_);
  and g_141974_(_083971_, _086432_, _086434_);
  not g_141975_(_086434_, _086435_);
  xor g_141976_(_083970_, _086432_, _086436_);
  or g_141977_(_083587_, _086436_, _086437_);
  xor g_141978_(_083586_, _086436_, _086438_);
  not g_141979_(_086438_, _086439_);
  and g_141980_(_083581_, _083591_, _086440_);
  xor g_141981_(_086439_, _086440_, _086441_);
  xor g_141982_(_083967_, _086441_, _086442_);
  not g_141983_(_086442_, _086443_);
  and g_141984_(_083599_, _086442_, _086445_);
  or g_141985_(_083598_, _086443_, _086446_);
  xor g_141986_(_083598_, _086442_, _086447_);
  not g_141987_(_086447_, _086448_);
  or g_141988_(_080609_, _083604_, _086449_);
  and g_141989_(_083602_, _086449_, _086450_);
  xor g_141990_(_086448_, _086450_, _086451_);
  or g_141991_(_083965_, _086451_, _086452_);
  xor g_141992_(_083966_, _086451_, _086453_);
  and g_141993_(_083609_, _086453_, _086454_);
  and g_141994_(_083964_, _086454_, _086456_);
  not g_141995_(_086456_, _086457_);
  or g_141996_(_083609_, _086453_, _086458_);
  or g_141997_(_083964_, _086453_, _086459_);
  not g_141998_(_086459_, _086460_);
  and g_141999_(_086458_, _086459_, _086461_);
  not g_142000_(_086461_, _086462_);
  and g_142001_(_086457_, _086461_, _086463_);
  or g_142002_(_086456_, _086462_, _086464_);
  or g_142003_(_083963_, _086464_, _086465_);
  xor g_142004_(_083963_, _086463_, _086467_);
  not g_142005_(_086467_, _086468_);
  or g_142006_(_080631_, _083616_, _086469_);
  and g_142007_(_083615_, _086469_, _086470_);
  xor g_142008_(_086467_, _086470_, _086471_);
  xor g_142009_(_086468_, _086470_, _086472_);
  or g_142010_(_083962_, _086472_, _086473_);
  xor g_142011_(_083962_, _086471_, _086474_);
  or g_142012_(_080637_, _083620_, _086475_);
  and g_142013_(_083621_, _086475_, _086476_);
  xor g_142014_(_086474_, _086476_, _086478_);
  and g_142015_(_083961_, _086478_, _086479_);
  not g_142016_(_086479_, _086480_);
  xor g_142017_(_083960_, _086478_, _086481_);
  not g_142018_(_086481_, _086482_);
  or g_142019_(_080647_, _083630_, _086483_);
  and g_142020_(_083627_, _086483_, _086484_);
  xor g_142021_(_086482_, _086484_, _086485_);
  or g_142022_(_083959_, _086485_, _086486_);
  xor g_142023_(_083959_, _086485_, _086487_);
  not g_142024_(_086487_, _086489_);
  or g_142025_(_083637_, _086489_, _086490_);
  xor g_142026_(_083637_, _086487_, _086491_);
  or g_142027_(_083643_, _086491_, _086492_);
  not g_142028_(_086492_, _086493_);
  or g_142029_(_083633_, _086491_, _086494_);
  not g_142030_(_086494_, _086495_);
  xor g_142031_(_083634_, _086491_, _086496_);
  and g_142032_(_083643_, _086496_, _086497_);
  or g_142033_(_086493_, _086497_, _086498_);
  not g_142034_(_086498_, _086500_);
  and g_142035_(_083646_, _083648_, _086501_);
  xor g_142036_(_086500_, _086501_, _086502_);
  or g_142037_(_083650_, _086502_, _086503_);
  not g_142038_(_086503_, _086504_);
  xor g_142039_(_083652_, _086502_, _086505_);
  or g_142040_(_083655_, _086505_, _086506_);
  not g_142041_(_086506_, _086507_);
  or g_142042_(_083658_, _086505_, _086508_);
  not g_142043_(_086508_, _086509_);
  xor g_142044_(_083659_, _086505_, _086511_);
  and g_142045_(_083655_, _086511_, _086512_);
  or g_142046_(_086507_, _086512_, _086513_);
  not g_142047_(_086513_, _086514_);
  or g_142048_(_083666_, _086513_, _086515_);
  xor g_142049_(_083663_, _086514_, _086516_);
  or g_142050_(_083670_, _086516_, _086517_);
  xor g_142051_(_083670_, _086516_, _086518_);
  or g_142052_(_083667_, _086518_, _086519_);
  and g_142053_(_086515_, _086519_, _086520_);
  not g_142054_(_086520_, _086522_);
  and g_142055_(_083674_, _086520_, _086523_);
  or g_142056_(_083672_, _086522_, _086524_);
  xor g_142057_(_083672_, _086520_, _086525_);
  and g_142058_(_083678_, _083682_, _086526_);
  xor g_142059_(_086525_, _086526_, _086527_);
  and g_142060_(_083686_, _083689_, _086528_);
  xor g_142061_(_086527_, _086528_, _086529_);
  xor g_142062_(_083957_, _086529_, _086530_);
  not g_142063_(_086530_, _086531_);
  and g_142064_(_083699_, _083703_, _086533_);
  xor g_142065_(_086530_, _086533_, _086534_);
  or g_142066_(_083708_, _086534_, _086535_);
  not g_142067_(_086535_, _086536_);
  and g_142068_(_083709_, _086534_, _086537_);
  and g_142069_(_083708_, _086537_, _086538_);
  or g_142070_(_083709_, _086534_, _086539_);
  not g_142071_(_086539_, _086540_);
  or g_142072_(_086538_, _086540_, _086541_);
  or g_142073_(_086536_, _086541_, _086542_);
  not g_142074_(_086542_, _086544_);
  or g_142075_(_083713_, _086542_, _086545_);
  not g_142076_(_086545_, _086546_);
  or g_142077_(_083715_, _086542_, _086547_);
  xor g_142078_(_083715_, _086544_, _086548_);
  and g_142079_(_083713_, _086548_, _086549_);
  or g_142080_(_086546_, _086549_, _086550_);
  or g_142081_(_083719_, _086550_, _086551_);
  xor g_142082_(_083718_, _086550_, _086552_);
  or g_142083_(_083721_, _086552_, _086553_);
  xor g_142084_(_083721_, _086552_, _086555_);
  xor g_142085_(_083722_, _086552_, _086556_);
  or g_142086_(_080739_, _083725_, _086557_);
  not g_142087_(_086557_, _086558_);
  and g_142088_(_083724_, _086557_, _086559_);
  xor g_142089_(_086556_, _086559_, _086560_);
  xor g_142090_(_086555_, _086559_, _086561_);
  or g_142091_(_083956_, _086561_, _086562_);
  xor g_142092_(_083956_, _086560_, _086563_);
  not g_142093_(_086563_, _086564_);
  or g_142094_(_080747_, _083732_, _086566_);
  and g_142095_(_083731_, _086566_, _086567_);
  xor g_142096_(_086563_, _086567_, _086568_);
  xor g_142097_(_086564_, _086567_, _086569_);
  or g_142098_(_083955_, _086569_, _086570_);
  xor g_142099_(_083955_, _086568_, _086571_);
  or g_142100_(_083744_, _086571_, _086572_);
  xor g_142101_(_083745_, _086571_, _086573_);
  or g_142102_(_083742_, _086573_, _086574_);
  xor g_142103_(_083743_, _086573_, _086575_);
  and g_142104_(_083751_, _083753_, _086577_);
  xor g_142105_(_086575_, _086577_, _086578_);
  not g_142106_(_086578_, _086579_);
  or g_142107_(_083755_, _086579_, _086580_);
  not g_142108_(_086580_, _086581_);
  xor g_142109_(_083755_, _086578_, _086582_);
  and g_142110_(_083757_, _083759_, _086583_);
  xor g_142111_(_086582_, _086583_, _086584_);
  not g_142112_(_086584_, _086585_);
  or g_142113_(_083953_, _086585_, _086586_);
  not g_142114_(_086586_, _086588_);
  xor g_142115_(_083954_, _086584_, _086589_);
  not g_142116_(_086589_, _086590_);
  or g_142117_(_083952_, _086590_, _086591_);
  not g_142118_(_086591_, _086592_);
  xor g_142119_(_083952_, _086589_, _086593_);
  or g_142120_(_083766_, _086593_, _086594_);
  xor g_142121_(_083766_, _086593_, _086595_);
  xor g_142122_(_083767_, _086593_, _086596_);
  and g_142123_(_083769_, _083771_, _086597_);
  xor g_142124_(_086596_, _086597_, _086599_);
  xor g_142125_(_086595_, _086597_, _086600_);
  and g_142126_(_083776_, _086599_, _086601_);
  or g_142127_(_083777_, _086600_, _086602_);
  and g_142128_(_080968_, _086601_, _086603_);
  or g_142129_(_080966_, _086602_, _086604_);
  xor g_142130_(_083775_, _086600_, _086605_);
  xor g_142131_(_083775_, _086599_, _086606_);
  and g_142132_(_083779_, _086606_, _086607_);
  or g_142133_(_083778_, _086605_, _086608_);
  and g_142134_(_086604_, _086608_, _086610_);
  or g_142135_(_086603_, _086607_, _086611_);
  and g_142136_(_083786_, _086610_, _086612_);
  or g_142137_(_083787_, _086611_, _086613_);
  or g_142138_(_083782_, _086606_, _086614_);
  not g_142139_(_086614_, _086615_);
  and g_142140_(_086613_, _086614_, _086616_);
  or g_142141_(_086612_, _086615_, _086617_);
  and g_142142_(_083782_, _086611_, _086618_);
  and g_142143_(_083787_, _086618_, _086619_);
  not g_142144_(_086619_, _086621_);
  and g_142145_(_086616_, _086621_, _086622_);
  or g_142146_(_086617_, _086619_, _086623_);
  xor g_142147_(_083951_, _086623_, _086624_);
  xor g_142148_(_083951_, _086622_, _086625_);
  or g_142149_(_083950_, _086625_, _086626_);
  xor g_142150_(_083950_, _086624_, _086627_);
  or g_142151_(_083946_, _086627_, _086628_);
  not g_142152_(_086628_, _086629_);
  xor g_142153_(_083946_, _086627_, _086630_);
  xor g_142154_(_083948_, _086627_, _086632_);
  and g_142155_(_080822_, _083798_, _086633_);
  or g_142156_(_080821_, _083799_, _086634_);
  and g_142157_(_086630_, _086633_, _086635_);
  and g_142158_(_083800_, _086630_, _086636_);
  not g_142159_(_086636_, _086637_);
  or g_142160_(_086635_, _086636_, _086638_);
  and g_142161_(_083801_, _086632_, _086639_);
  and g_142162_(_086634_, _086639_, _086640_);
  or g_142163_(_086638_, _086640_, _086641_);
  or g_142164_(_083944_, _086641_, _086643_);
  xor g_142165_(_083945_, _086641_, _086644_);
  or g_142166_(_083809_, _086644_, _086645_);
  or g_142167_(_083810_, _086645_, _086646_);
  or g_142168_(_083807_, _086644_, _086647_);
  xor g_142169_(_083807_, _086644_, _086648_);
  or g_142170_(_083812_, _086648_, _086649_);
  and g_142171_(_086646_, _086649_, _086650_);
  or g_142172_(_083814_, _083818_, _086651_);
  and g_142173_(_086650_, _086651_, _086652_);
  not g_142174_(_086652_, _086654_);
  xor g_142175_(_086650_, _086651_, _086655_);
  not g_142176_(_086655_, _086656_);
  or g_142177_(_083822_, _086656_, _086657_);
  xor g_142178_(_083822_, _086655_, _086658_);
  or g_142179_(_083824_, _086658_, _086659_);
  xor g_142180_(_083825_, _086658_, _086660_);
  or g_142181_(_083832_, _086660_, _086661_);
  xor g_142182_(_083831_, _086660_, _086662_);
  not g_142183_(_086662_, _086663_);
  and g_142184_(_083833_, _086663_, _086665_);
  not g_142185_(_086665_, _086666_);
  xor g_142186_(_083833_, _086662_, _086667_);
  or g_142187_(_083839_, _086667_, _086668_);
  not g_142188_(_086668_, _086669_);
  xor g_142189_(_083839_, _086667_, _086670_);
  xor g_142190_(_083837_, _086667_, _086671_);
  and g_142191_(_083841_, _083845_, _086672_);
  xor g_142192_(_086671_, _086672_, _086673_);
  xor g_142193_(_086670_, _086672_, _086674_);
  or g_142194_(_083943_, _086674_, _086676_);
  xor g_142195_(_083943_, _086674_, _086677_);
  xor g_142196_(_083943_, _086673_, _086678_);
  or g_142197_(_080863_, _083846_, _086679_);
  not g_142198_(_086679_, _086680_);
  or g_142199_(_086677_, _086680_, _086681_);
  not g_142200_(_086681_, _086682_);
  and g_142201_(_083853_, _086682_, _086683_);
  or g_142202_(_083852_, _086681_, _086684_);
  and g_142203_(_083852_, _086677_, _086685_);
  or g_142204_(_083853_, _086678_, _086687_);
  and g_142205_(_086677_, _086680_, _086688_);
  or g_142206_(_086678_, _086679_, _086689_);
  and g_142207_(_086687_, _086689_, _086690_);
  or g_142208_(_086685_, _086688_, _086691_);
  and g_142209_(_086684_, _086690_, _086692_);
  or g_142210_(_086683_, _086691_, _086693_);
  or g_142211_(_083861_, _086693_, _086694_);
  not g_142212_(_086694_, _086695_);
  and g_142213_(_083856_, _086693_, _086696_);
  or g_142214_(_083855_, _086692_, _086698_);
  and g_142215_(_083861_, _086696_, _086699_);
  or g_142216_(_083862_, _086698_, _086700_);
  and g_142217_(_083855_, _086692_, _086701_);
  not g_142218_(_086701_, _086702_);
  and g_142219_(_086700_, _086702_, _086703_);
  or g_142220_(_086699_, _086701_, _086704_);
  and g_142221_(_086694_, _086703_, _086705_);
  or g_142222_(_086695_, _086704_, _086706_);
  or g_142223_(_080886_, _083866_, _086707_);
  and g_142224_(_083863_, _086707_, _086709_);
  xor g_142225_(_086705_, _086709_, _086710_);
  xor g_142226_(_086706_, _086709_, _086711_);
  and g_142227_(_083942_, _086711_, _086712_);
  not g_142228_(_086712_, _086713_);
  xor g_142229_(_083941_, _086710_, _086714_);
  xor g_142230_(_083942_, _086710_, _086715_);
  or g_142231_(_083869_, _086715_, _086716_);
  xor g_142232_(_083869_, _086714_, _086717_);
  or g_142233_(_083876_, _086717_, _086718_);
  not g_142234_(_086718_, _086720_);
  and g_142235_(_083874_, _086714_, _086721_);
  not g_142236_(_086721_, _086722_);
  and g_142237_(_083873_, _086717_, _086723_);
  or g_142238_(_086721_, _086723_, _086724_);
  and g_142239_(_083876_, _086724_, _086725_);
  or g_142240_(_086720_, _086725_, _086726_);
  not g_142241_(_086726_, _086727_);
  xor g_142242_(_083940_, _086727_, _086728_);
  xor g_142243_(_083940_, _086726_, _086729_);
  or g_142244_(_083939_, _086728_, _086731_);
  xor g_142245_(_083939_, _086729_, _086732_);
  not g_142246_(_086732_, _086733_);
  or g_142247_(_083884_, _086732_, _086734_);
  xor g_142248_(_083884_, _086732_, _086735_);
  xor g_142249_(_083884_, _086733_, _086736_);
  or g_142250_(_083887_, _086736_, _086737_);
  xor g_142251_(_083887_, _086735_, _086738_);
  or g_142252_(_083938_, _086738_, _086739_);
  xor g_142253_(_083938_, _086738_, _086740_);
  xor g_142254_(_083937_, _086738_, _086742_);
  and g_142255_(_083935_, _086740_, _086743_);
  or g_142256_(_083934_, _086742_, _086744_);
  xor g_142257_(_083935_, _086740_, _086745_);
  xor g_142258_(_083934_, _086740_, _086746_);
  and g_142259_(_083897_, _086746_, _086747_);
  or g_142260_(_083896_, _086745_, _086748_);
  and g_142261_(_083906_, _086747_, _086749_);
  or g_142262_(_083905_, _086748_, _086750_);
  and g_142263_(_083905_, _086745_, _086751_);
  or g_142264_(_083906_, _086746_, _086753_);
  and g_142265_(_083896_, _086745_, _086754_);
  or g_142266_(_083897_, _086746_, _086755_);
  and g_142267_(_086753_, _086755_, _086756_);
  or g_142268_(_086751_, _086754_, _086757_);
  and g_142269_(_086750_, _086756_, _086758_);
  or g_142270_(_086749_, _086757_, _086759_);
  and g_142271_(_083902_, _086758_, _086760_);
  or g_142272_(_083903_, _086759_, _086761_);
  xor g_142273_(_083903_, _086758_, _086762_);
  or g_142274_(_083912_, _086762_, _086764_);
  not g_142275_(_086764_, _086765_);
  or g_142276_(_083909_, _086762_, _086766_);
  not g_142277_(_086766_, _086767_);
  and g_142278_(_083909_, _086762_, _086768_);
  and g_142279_(_083912_, _086768_, _086769_);
  or g_142280_(_086767_, _086769_, _086770_);
  or g_142281_(_086765_, _086770_, _086771_);
  not g_142282_(_086771_, _086772_);
  or g_142283_(_083933_, _086771_, _086773_);
  xor g_142284_(_083933_, _086771_, _086775_);
  xor g_142285_(_083933_, _086772_, _086776_);
  or g_142286_(_083932_, _086776_, _086777_);
  xor g_142287_(_083932_, _086775_, _086778_);
  not g_142288_(_086778_, _086779_);
  or g_142289_(_083919_, _086778_, _086780_);
  xor g_142290_(_083919_, _086779_, _086781_);
  not g_142291_(_086781_, _086782_);
  and g_142292_(_083928_, _086782_, _086783_);
  or g_142293_(_083929_, _086781_, _086784_);
  or g_142294_(_083924_, _086781_, _086786_);
  xor g_142295_(_083924_, _086782_, _086787_);
  or g_142296_(_083931_, _086787_, _086788_);
  xor g_142297_(_083931_, _086787_, _086789_);
  or g_142298_(_083928_, _086789_, _086790_);
  and g_142299_(_086784_, _086790_, out[964]);
  or g_142300_(_086706_, _086707_, _086791_);
  or g_142301_(_083845_, _086671_, _086792_);
  and g_142302_(_086657_, _086659_, _086793_);
  and g_142303_(_086643_, _086647_, _086794_);
  and g_142304_(_083795_, _086622_, _086796_);
  not g_142305_(_086796_, _086797_);
  or g_142306_(_083789_, _086623_, _086798_);
  or g_142307_(_080788_, _083773_, _086799_);
  or g_142308_(_086600_, _086799_, _086800_);
  or g_142309_(_080786_, _083773_, _086801_);
  not g_142310_(_086801_, _086802_);
  and g_142311_(_086599_, _086802_, _086803_);
  not g_142312_(_086803_, _086804_);
  or g_142313_(_083771_, _086596_, _086805_);
  not g_142314_(_086805_, _086807_);
  or g_142315_(_083759_, _086582_, _086808_);
  or g_142316_(_083757_, _086582_, _086809_);
  not g_142317_(_086809_, _086810_);
  or g_142318_(_083753_, _086575_, _086811_);
  not g_142319_(_086811_, _086812_);
  or g_142320_(_086563_, _086566_, _086813_);
  not g_142321_(_086813_, _086814_);
  or g_142322_(_083731_, _086563_, _086815_);
  and g_142323_(_086555_, _086558_, _086816_);
  or g_142324_(_086556_, _086557_, _086818_);
  or g_142325_(_083724_, _086552_, _086819_);
  or g_142326_(_083703_, _086531_, _086820_);
  and g_142327_(_083700_, _086530_, _086821_);
  or g_142328_(_083699_, _086531_, _086822_);
  or g_142329_(_083697_, _086529_, _086823_);
  or g_142330_(_083694_, _086529_, _086824_);
  and g_142331_(_083690_, _086527_, _086825_);
  and g_142332_(_083687_, _086527_, _086826_);
  not g_142333_(_086826_, _086827_);
  or g_142334_(_083682_, _086525_, _086829_);
  or g_142335_(_080680_, _083660_, _086830_);
  or g_142336_(_086513_, _086830_, _086831_);
  or g_142337_(_080677_, _083660_, _086832_);
  or g_142338_(_086513_, _086832_, _086833_);
  not g_142339_(_086833_, _086834_);
  or g_142340_(_083648_, _086498_, _086835_);
  not g_142341_(_086835_, _086836_);
  or g_142342_(_086481_, _086483_, _086837_);
  not g_142343_(_086837_, _086838_);
  or g_142344_(_083627_, _086481_, _086840_);
  or g_142345_(_086474_, _086475_, _086841_);
  not g_142346_(_086841_, _086842_);
  or g_142347_(_083621_, _086474_, _086843_);
  or g_142348_(_086467_, _086469_, _086844_);
  or g_142349_(_086447_, _086449_, _086845_);
  or g_142350_(_083602_, _086447_, _086846_);
  or g_142351_(_083595_, _086441_, _086847_);
  not g_142352_(_086847_, _086848_);
  or g_142353_(_083593_, _086441_, _086849_);
  or g_142354_(_083591_, _086438_, _086851_);
  or g_142355_(_083581_, _086438_, _086852_);
  or g_142356_(_083572_, _086427_, _086853_);
  or g_142357_(_083568_, _086424_, _086854_);
  or g_142358_(_083564_, _086424_, _086855_);
  or g_142359_(_083545_, _086398_, _086856_);
  not g_142360_(_086856_, _086857_);
  or g_142361_(_083527_, _086386_, _086858_);
  or g_142362_(_080535_, _086858_, _086859_);
  not g_142363_(_086859_, _086860_);
  or g_142364_(_080533_, _086858_, _086862_);
  or g_142365_(_083513_, _086376_, _086863_);
  or g_142366_(_080519_, _086863_, _086864_);
  not g_142367_(_086864_, _086865_);
  or g_142368_(_083507_, _086366_, _086866_);
  or g_142369_(_083487_, _086342_, _086867_);
  not g_142370_(_086867_, _086868_);
  or g_142371_(_083466_, _086320_, _086869_);
  or g_142372_(_083457_, _086317_, _086870_);
  not g_142373_(_086870_, _086871_);
  or g_142374_(_083454_, _086314_, _086873_);
  or g_142375_(_083446_, _086305_, _086874_);
  or g_142376_(_083986_, _086305_, _086875_);
  or g_142377_(_083427_, _086289_, _086876_);
  or g_142378_(_083425_, _086289_, _086877_);
  or g_142379_(_083422_, _086286_, _086878_);
  or g_142380_(_083418_, _086286_, _086879_);
  or g_142381_(_086271_, _086273_, _086880_);
  or g_142382_(_083405_, _086271_, _086881_);
  and g_142383_(_086270_, _086881_, _086882_);
  or g_142384_(_083394_, _086260_, _086884_);
  not g_142385_(_086884_, _086885_);
  and g_142386_(_083389_, _086259_, _086886_);
  or g_142387_(_083388_, _086260_, _086887_);
  or g_142388_(_083385_, _086256_, _086888_);
  or g_142389_(_083382_, _086256_, _086889_);
  or g_142390_(_080338_, _083338_, _086890_);
  or g_142391_(_086216_, _086890_, _086891_);
  or g_142392_(_083323_, _086198_, _086892_);
  and g_142393_(_086203_, _086892_, _086893_);
  or g_142394_(_083303_, _086172_, _086895_);
  or g_142395_(_083298_, _086167_, _086896_);
  or g_142396_(_083295_, _086164_, _086897_);
  or g_142397_(_083290_, _086161_, _086898_);
  or g_142398_(_083275_, _086144_, _086899_);
  and g_142399_(_086154_, _086899_, _086900_);
  not g_142400_(_086900_, _086901_);
  or g_142401_(_083268_, _086141_, _086902_);
  or g_142402_(_080248_, _086902_, _086903_);
  not g_142403_(_086903_, _086904_);
  or g_142404_(_084005_, _086139_, _086906_);
  or g_142405_(_083258_, _086139_, _086907_);
  or g_142406_(_083262_, _086137_, _086908_);
  or g_142407_(_083256_, _086137_, _086909_);
  not g_142408_(_086909_, _086910_);
  and g_142409_(_083239_, _086120_, _086911_);
  not g_142410_(_086911_, _086912_);
  or g_142411_(_083240_, _086119_, _086913_);
  or g_142412_(_083199_, _086072_, _086914_);
  not g_142413_(_086914_, _086915_);
  or g_142414_(_086072_, _086074_, _086917_);
  not g_142415_(_086917_, _086918_);
  or g_142416_(_083194_, _086067_, _086919_);
  not g_142417_(_086919_, _086920_);
  or g_142418_(_083191_, _086065_, _086921_);
  not g_142419_(_086921_, _086922_);
  and g_142420_(_083188_, _086064_, _086923_);
  or g_142421_(_083187_, _086065_, _086924_);
  and g_142422_(_086053_, _086055_, _086925_);
  or g_142423_(_086041_, _086043_, _086926_);
  and g_142424_(_083152_, _086031_, _086928_);
  and g_142425_(_083147_, _086031_, _086929_);
  or g_142426_(_086025_, _086027_, _086930_);
  or g_142427_(_083140_, _086025_, _086931_);
  or g_142428_(_083132_, _086013_, _086932_);
  not g_142429_(_086932_, _086933_);
  or g_142430_(_086013_, _086016_, _086934_);
  not g_142431_(_086934_, _086935_);
  or g_142432_(_083122_, _086000_, _086936_);
  not g_142433_(_086936_, _086937_);
  or g_142434_(_083115_, _086000_, _086939_);
  not g_142435_(_086939_, _086940_);
  or g_142436_(_083116_, _086000_, _086941_);
  not g_142437_(_086941_, _086942_);
  or g_142438_(_083096_, _085975_, _086943_);
  or g_142439_(_080096_, _086943_, _086944_);
  or g_142440_(_080093_, _086943_, _086945_);
  or g_142441_(_083092_, _085952_, _086946_);
  and g_142442_(_084034_, _085929_, _086947_);
  or g_142443_(_083073_, _085928_, _086948_);
  or g_142444_(_083070_, _085923_, _086950_);
  and g_142445_(_085891_, _085893_, _086951_);
  not g_142446_(_086951_, _086952_);
  or g_142447_(_083044_, _085890_, _086953_);
  and g_142448_(_085889_, _086953_, _086954_);
  and g_142449_(_085885_, _085887_, _086955_);
  and g_142450_(_085864_, _085867_, _086956_);
  or g_142451_(_083022_, _085865_, _086957_);
  or g_142452_(_082992_, _085835_, _086958_);
  or g_142453_(_082986_, _085834_, _086959_);
  or g_142454_(_082977_, _082978_, _086961_);
  or g_142455_(_085834_, _086961_, _086962_);
  not g_142456_(_086962_, _086963_);
  or g_142457_(_079973_, _082977_, _086964_);
  or g_142458_(_085834_, _086964_, _086965_);
  or g_142459_(_082948_, _085796_, _086966_);
  or g_142460_(_082944_, _085793_, _086967_);
  or g_142461_(_082907_, _085753_, _086968_);
  or g_142462_(_079905_, _086968_, _086969_);
  not g_142463_(_086969_, _086970_);
  or g_142464_(_079900_, _086968_, _086972_);
  or g_142465_(_082906_, _085750_, _086973_);
  and g_142466_(_082904_, _085749_, _086974_);
  or g_142467_(_082902_, _085750_, _086975_);
  or g_142468_(_082900_, _085746_, _086976_);
  and g_142469_(_085719_, _085722_, _086977_);
  and g_142470_(_085670_, _085675_, _086978_);
  not g_142471_(_086978_, _086979_);
  or g_142472_(_082805_, _082807_, _086980_);
  or g_142473_(_085637_, _086980_, _086981_);
  not g_142474_(_086981_, _086983_);
  or g_142475_(_079826_, _082805_, _086984_);
  or g_142476_(_085637_, _086984_, _086985_);
  and g_142477_(_085628_, _085633_, _086986_);
  not g_142478_(_086986_, _086987_);
  or g_142479_(_082773_, _085603_, _086988_);
  or g_142480_(_079794_, _086988_, _086989_);
  or g_142481_(_079789_, _086988_, _086990_);
  or g_142482_(_082772_, _085601_, _086991_);
  not g_142483_(_086991_, _086992_);
  or g_142484_(_082769_, _085601_, _086994_);
  not g_142485_(_086994_, _086995_);
  and g_142486_(_082750_, _085573_, _086996_);
  or g_142487_(_082742_, _085574_, _086997_);
  not g_142488_(_086997_, _086998_);
  or g_142489_(_085557_, _085558_, _086999_);
  not g_142490_(_086999_, _087000_);
  or g_142491_(_082712_, _085541_, _087001_);
  and g_142492_(_085474_, _085477_, _087002_);
  or g_142493_(_084098_, _085449_, _087003_);
  not g_142494_(_087003_, _087005_);
  and g_142495_(_082626_, _085448_, _087006_);
  or g_142496_(_082623_, _085446_, _087007_);
  not g_142497_(_087007_, _087008_);
  or g_142498_(_082607_, _085434_, _087009_);
  and g_142499_(_082601_, _085429_, _087010_);
  not g_142500_(_087010_, _087011_);
  or g_142501_(_082553_, _085383_, _087012_);
  or g_142502_(_082560_, _087012_, _087013_);
  not g_142503_(_087013_, _087014_);
  or g_142504_(_079610_, _087012_, _087016_);
  or g_142505_(_082554_, _085382_, _087017_);
  or g_142506_(_082556_, _085382_, _087018_);
  or g_142507_(_085373_, _085374_, _087019_);
  or g_142508_(_085373_, _085375_, _087020_);
  or g_142509_(_079524_, _082479_, _087021_);
  or g_142510_(_085287_, _087021_, _087022_);
  or g_142511_(_079522_, _085286_, _087023_);
  or g_142512_(_082479_, _087023_, _087024_);
  or g_142513_(_079519_, _082473_, _087025_);
  or g_142514_(_085286_, _087025_, _087027_);
  and g_142515_(_085270_, _085273_, _087028_);
  not g_142516_(_087028_, _087029_);
  or g_142517_(_084126_, _085244_, _087030_);
  or g_142518_(_082400_, _085210_, _087031_);
  or g_142519_(_082392_, _085210_, _087032_);
  and g_142520_(_085209_, _087032_, _087033_);
  or g_142521_(_082372_, _085197_, _087034_);
  or g_142522_(_082374_, _085197_, _087035_);
  not g_142523_(_087035_, _087036_);
  or g_142524_(_082368_, _085193_, _087038_);
  or g_142525_(_082366_, _085193_, _087039_);
  or g_142526_(_085184_, _085186_, _087040_);
  not g_142527_(_087040_, _087041_);
  or g_142528_(_082359_, _085184_, _087042_);
  or g_142529_(_082329_, _085164_, _087043_);
  or g_142530_(_082327_, _085164_, _087044_);
  not g_142531_(_087044_, _087045_);
  or g_142532_(_082324_, _085160_, _087046_);
  not g_142533_(_087046_, _087047_);
  and g_142534_(_085159_, _085162_, _087049_);
  or g_142535_(_085160_, _085161_, _087050_);
  or g_142536_(_085128_, _085130_, _087051_);
  not g_142537_(_087051_, _087052_);
  or g_142538_(_085128_, _085129_, _087053_);
  or g_142539_(_085123_, _085125_, _087054_);
  and g_142540_(_082299_, _085120_, _087055_);
  not g_142541_(_087055_, _087056_);
  or g_142542_(_082293_, _085119_, _087057_);
  and g_142543_(_085118_, _087057_, _087058_);
  and g_142544_(_085111_, _085115_, _087060_);
  not g_142545_(_087060_, _087061_);
  or g_142546_(_082260_, _085068_, _087062_);
  not g_142547_(_087062_, _087063_);
  or g_142548_(_082212_, _085015_, _087064_);
  or g_142549_(_082209_, _085015_, _087065_);
  not g_142550_(_087065_, _087066_);
  and g_142551_(_085013_, _087065_, _087067_);
  or g_142552_(_082175_, _084990_, _087068_);
  or g_142553_(_082176_, _084990_, _087069_);
  or g_142554_(_082157_, _084966_, _087071_);
  or g_142555_(_082151_, _084963_, _087072_);
  and g_142556_(_084967_, _087072_, _087073_);
  or g_142557_(_082140_, _084960_, _087074_);
  not g_142558_(_087074_, _087075_);
  and g_142559_(_082138_, _084958_, _087076_);
  not g_142560_(_087076_, _087077_);
  or g_142561_(_082134_, _084956_, _087078_);
  not g_142562_(_087078_, _087079_);
  or g_142563_(_082130_, _084953_, _087080_);
  or g_142564_(_079199_, _082117_, _087082_);
  or g_142565_(_084943_, _087082_, _087083_);
  or g_142566_(_084922_, _084923_, _087084_);
  not g_142567_(_087084_, _087085_);
  or g_142568_(_082105_, _084922_, _087086_);
  or g_142569_(_079154_, _082082_, _087087_);
  or g_142570_(_084906_, _087087_, _087088_);
  and g_142571_(_079151_, _084902_, _087089_);
  not g_142572_(_087089_, _087090_);
  or g_142573_(_082082_, _087090_, _087091_);
  or g_142574_(_084172_, _084899_, _087093_);
  not g_142575_(_087093_, _087094_);
  or g_142576_(_082074_, _084899_, _087095_);
  and g_142577_(_082072_, _084896_, _087096_);
  not g_142578_(_087096_, _087097_);
  or g_142579_(_082069_, _084895_, _087098_);
  and g_142580_(_084884_, _084889_, _087099_);
  or g_142581_(_082044_, _084877_, _087100_);
  or g_142582_(_082041_, _084877_, _087101_);
  and g_142583_(_084872_, _084875_, _087102_);
  or g_142584_(_081961_, _084825_, _087104_);
  not g_142585_(_087104_, _087105_);
  or g_142586_(_081959_, _084825_, _087106_);
  not g_142587_(_087106_, _087107_);
  or g_142588_(_079053_, _081953_, _087108_);
  or g_142589_(_084823_, _087108_, _087109_);
  or g_142590_(_079050_, _081953_, _087110_);
  or g_142591_(_084823_, _087110_, _087111_);
  not g_142592_(_087111_, _087112_);
  or g_142593_(_081940_, _084811_, _087113_);
  not g_142594_(_087113_, _087115_);
  and g_142595_(_084807_, _084809_, _087116_);
  or g_142596_(_084793_, _084796_, _087117_);
  or g_142597_(_081925_, _084793_, _087118_);
  and g_142598_(_081901_, _084769_, _087119_);
  not g_142599_(_087119_, _087120_);
  or g_142600_(_084770_, _084771_, _087121_);
  or g_142601_(_084766_, _084767_, _087122_);
  not g_142602_(_087122_, _087123_);
  or g_142603_(_081892_, _084766_, _087124_);
  not g_142604_(_087124_, _087126_);
  or g_142605_(_081883_, _084758_, _087127_);
  not g_142606_(_087127_, _087128_);
  or g_142607_(_081879_, _084758_, _087129_);
  or g_142608_(_081875_, _084756_, _087130_);
  or g_142609_(_081874_, _084752_, _087131_);
  or g_142610_(_081846_, _084727_, _087132_);
  not g_142611_(_087132_, _087133_);
  or g_142612_(_081849_, _084727_, _087134_);
  not g_142613_(_087134_, _087135_);
  or g_142614_(_081818_, _084697_, _087137_);
  or g_142615_(_081816_, _084697_, _087138_);
  not g_142616_(_087138_, _087139_);
  or g_142617_(_081809_, _084689_, _087140_);
  not g_142618_(_087140_, _087141_);
  or g_142619_(_081806_, _084686_, _087142_);
  or g_142620_(_081778_, _084663_, _087143_);
  not g_142621_(_087143_, _087144_);
  or g_142622_(_081776_, _084663_, _087145_);
  or g_142623_(_081774_, _084658_, _087146_);
  or g_142624_(_081756_, _084632_, _087148_);
  or g_142625_(_081753_, _084632_, _087149_);
  not g_142626_(_087149_, _087150_);
  or g_142627_(_084602_, _084603_, _087151_);
  not g_142628_(_087151_, _087152_);
  or g_142629_(_081709_, _084594_, _087153_);
  or g_142630_(_081707_, _084594_, _087154_);
  not g_142631_(_087154_, _087155_);
  or g_142632_(_081669_, _084557_, _087156_);
  or g_142633_(_081667_, _084557_, _087157_);
  or g_142634_(_081662_, _084556_, _087159_);
  or g_142635_(_078783_, _087159_, _087160_);
  or g_142636_(_078780_, _087159_, _087161_);
  and g_142637_(_081648_, _084537_, _087162_);
  or g_142638_(_081647_, _084538_, _087163_);
  or g_142639_(_081635_, _084525_, _087164_);
  or g_142640_(_081633_, _084525_, _087165_);
  or g_142641_(_081560_, _084446_, _087166_);
  or g_142642_(_081552_, _084446_, _087167_);
  not g_142643_(_087167_, _087168_);
  and g_142644_(_084443_, _084445_, _087170_);
  not g_142645_(_087170_, _087171_);
  or g_142646_(_081533_, _084436_, _087172_);
  not g_142647_(_087172_, _087173_);
  and g_142648_(_084394_, _084397_, _087174_);
  or g_142649_(_081475_, _084386_, _087175_);
  or g_142650_(_081471_, _084386_, _087176_);
  or g_142651_(_081459_, _084372_, _087177_);
  or g_142652_(_081453_, _084369_, _087178_);
  and g_142653_(_081457_, _084371_, _087179_);
  or g_142654_(_081456_, _084372_, _087181_);
  and g_142655_(_087178_, _087181_, _087182_);
  or g_142656_(_081449_, _084369_, _087183_);
  and g_142657_(_081447_, _084367_, _087184_);
  not g_142658_(_087184_, _087185_);
  and g_142659_(_081442_, _084367_, _087186_);
  or g_142660_(_081431_, _084353_, _087187_);
  not g_142661_(_087187_, _087188_);
  or g_142662_(_081421_, _084353_, _087189_);
  or g_142663_(_081419_, _084351_, _087190_);
  not g_142664_(_087190_, _087192_);
  and g_142665_(_081412_, _084350_, _087193_);
  or g_142666_(_081403_, _084341_, _087194_);
  or g_142667_(_081384_, _084333_, _087195_);
  and g_142668_(_081386_, _084230_, _087196_);
  or g_142669_(_084329_, _087196_, _087197_);
  and g_142670_(_084328_, _087197_, _087198_);
  and g_142671_(_084236_, _084325_, _087199_);
  or g_142672_(_084324_, _087199_, _087200_);
  and g_142673_(_084309_, _084313_, _087201_);
  or g_142674_(_084242_, _084302_, _087203_);
  or g_142675_(_081338_, _084275_, _087204_);
  or g_142676_(_078511_, _084274_, _087205_);
  or g_142677_(_078513_, _084269_, _087206_);
  and g_142678_(_087205_, _087206_, _087207_);
  or g_142679_(_081331_, _087207_, _087208_);
  and g_142680_(_084268_, _084270_, _087209_);
  and g_142681_(_084272_, _087209_, _087210_);
  and g_142682_(_087208_, _087210_, _087211_);
  and g_142683_(_087204_, _087211_, _087212_);
  and g_142684_(_084281_, _087212_, _087214_);
  and g_142685_(_084284_, _087214_, _087215_);
  and g_142686_(_084290_, _087215_, _087216_);
  or g_142687_(_081358_, _084293_, _087217_);
  and g_142688_(_084294_, _087217_, _087218_);
  and g_142689_(_087216_, _087218_, _087219_);
  or g_142690_(_081365_, _084298_, _087220_);
  and g_142691_(_084300_, _087220_, _087221_);
  and g_142692_(_087219_, _087221_, _087222_);
  and g_142693_(_087203_, _087222_, _087223_);
  xor g_142694_(_084306_, _087223_, _087225_);
  xor g_142695_(_087201_, _087225_, _087226_);
  or g_142696_(_081376_, _084318_, _087227_);
  and g_142697_(_084317_, _087227_, _087228_);
  xor g_142698_(_087226_, _087228_, _087229_);
  xor g_142699_(_084322_, _087229_, _087230_);
  xor g_142700_(_087200_, _087230_, _087231_);
  xor g_142701_(_087198_, _087231_, _087232_);
  xor g_142702_(_087195_, _087232_, _087233_);
  xor g_142703_(_084336_, _087233_, _087234_);
  and g_142704_(_081397_, _084339_, _087236_);
  or g_142705_(_084340_, _087236_, _087237_);
  not g_142706_(_087237_, _087238_);
  xor g_142707_(_087234_, _087237_, _087239_);
  xor g_142708_(_087234_, _087238_, _087240_);
  or g_142709_(_087194_, _087240_, _087241_);
  xor g_142710_(_087194_, _087239_, _087242_);
  or g_142711_(_084346_, _087242_, _087243_);
  xor g_142712_(_084346_, _087242_, _087244_);
  and g_142713_(_087193_, _087244_, _087245_);
  not g_142714_(_087245_, _087247_);
  or g_142715_(_084349_, _087244_, _087248_);
  or g_142716_(_084348_, _087242_, _087249_);
  and g_142717_(_087248_, _087249_, _087250_);
  or g_142718_(_087193_, _087250_, _087251_);
  and g_142719_(_087247_, _087251_, _087252_);
  xor g_142720_(_087190_, _087252_, _087253_);
  or g_142721_(_087189_, _087253_, _087254_);
  and g_142722_(_087189_, _087253_, _087255_);
  xor g_142723_(_087189_, _087253_, _087256_);
  xor g_142724_(_087188_, _087256_, _087258_);
  and g_142725_(_084357_, _087258_, _087259_);
  or g_142726_(_084357_, _087258_, _087260_);
  xor g_142727_(_084358_, _087258_, _087261_);
  or g_142728_(_084225_, _084363_, _087262_);
  and g_142729_(_084362_, _087262_, _087263_);
  xor g_142730_(_087261_, _087263_, _087264_);
  or g_142731_(_087186_, _087264_, _087265_);
  and g_142732_(_087186_, _087264_, _087266_);
  xor g_142733_(_087186_, _087264_, _087267_);
  xor g_142734_(_087185_, _087267_, _087269_);
  xor g_142735_(_087183_, _087269_, _087270_);
  not g_142736_(_087270_, _087271_);
  xor g_142737_(_087182_, _087271_, _087272_);
  xor g_142738_(_087182_, _087270_, _087273_);
  or g_142739_(_087177_, _087273_, _087274_);
  and g_142740_(_087177_, _087273_, _087275_);
  xor g_142741_(_087177_, _087272_, _087276_);
  not g_142742_(_087276_, _087277_);
  and g_142743_(_084374_, _084378_, _087278_);
  xor g_142744_(_087277_, _087278_, _087280_);
  or g_142745_(_084381_, _087280_, _087281_);
  xor g_142746_(_084382_, _087280_, _087282_);
  not g_142747_(_087282_, _087283_);
  or g_142748_(_084385_, _087282_, _087284_);
  xor g_142749_(_084385_, _087283_, _087285_);
  and g_142750_(_087176_, _087285_, _087286_);
  and g_142751_(_087175_, _087286_, _087287_);
  or g_142752_(_087176_, _087282_, _087288_);
  and g_142753_(_087175_, _087288_, _087289_);
  or g_142754_(_087286_, _087289_, _087291_);
  not g_142755_(_087291_, _087292_);
  or g_142756_(_087287_, _087292_, _087293_);
  not g_142757_(_087293_, _087294_);
  xor g_142758_(_084391_, _087294_, _087295_);
  not g_142759_(_087295_, _087296_);
  xor g_142760_(_087174_, _087296_, _087297_);
  or g_142761_(_084401_, _087297_, _087298_);
  xor g_142762_(_084401_, _087297_, _087299_);
  xor g_142763_(_084402_, _087297_, _087300_);
  and g_142764_(_084410_, _087299_, _087302_);
  or g_142765_(_084411_, _087300_, _087303_);
  or g_142766_(_084404_, _087300_, _087304_);
  xor g_142767_(_084404_, _087300_, _087305_);
  or g_142768_(_084410_, _087305_, _087306_);
  and g_142769_(_087303_, _087306_, _087307_);
  xor g_142770_(_084413_, _087307_, _087308_);
  not g_142771_(_087308_, _087309_);
  or g_142772_(_084417_, _087308_, _087310_);
  and g_142773_(_084417_, _087308_, _087311_);
  xor g_142774_(_084417_, _087309_, _087313_);
  or g_142775_(_081516_, _084422_, _087314_);
  and g_142776_(_084421_, _087314_, _087315_);
  xor g_142777_(_087313_, _087315_, _087316_);
  and g_142778_(_084428_, _087316_, _087317_);
  or g_142779_(_081520_, _084423_, _087318_);
  not g_142780_(_087318_, _087319_);
  and g_142781_(_087316_, _087319_, _087320_);
  xor g_142782_(_087316_, _087318_, _087321_);
  and g_142783_(_084427_, _087321_, _087322_);
  not g_142784_(_087322_, _087324_);
  or g_142785_(_087317_, _087322_, _087325_);
  xor g_142786_(_084430_, _087325_, _087326_);
  and g_142787_(_081530_, _084434_, _087327_);
  or g_142788_(_084435_, _087327_, _087328_);
  or g_142789_(_087326_, _087328_, _087329_);
  xor g_142790_(_087326_, _087328_, _087330_);
  and g_142791_(_087173_, _087330_, _087331_);
  xor g_142792_(_087172_, _087330_, _087332_);
  or g_142793_(_084440_, _087332_, _087333_);
  xor g_142794_(_084440_, _087332_, _087335_);
  not g_142795_(_087335_, _087336_);
  and g_142796_(_087171_, _087335_, _087337_);
  xor g_142797_(_087170_, _087335_, _087338_);
  or g_142798_(_087167_, _087338_, _087339_);
  xor g_142799_(_087168_, _087338_, _087340_);
  and g_142800_(_087166_, _087340_, _087341_);
  or g_142801_(_087166_, _087338_, _087342_);
  not g_142802_(_087342_, _087343_);
  or g_142803_(_087341_, _087343_, _087344_);
  and g_142804_(_084451_, _087344_, _087346_);
  not g_142805_(_087346_, _087347_);
  or g_142806_(_084451_, _087340_, _087348_);
  not g_142807_(_087348_, _087349_);
  and g_142808_(_084455_, _087348_, _087350_);
  not g_142809_(_087350_, _087351_);
  or g_142810_(_087346_, _087351_, _087352_);
  and g_142811_(_087347_, _087348_, _087353_);
  or g_142812_(_087346_, _087349_, _087354_);
  or g_142813_(_084455_, _087353_, _087355_);
  and g_142814_(_084458_, _087355_, _087357_);
  and g_142815_(_087352_, _087357_, _087358_);
  or g_142816_(_084458_, _087354_, _087359_);
  not g_142817_(_087359_, _087360_);
  or g_142818_(_087358_, _087360_, _087361_);
  not g_142819_(_087361_, _087362_);
  and g_142820_(_084461_, _084463_, _087363_);
  xor g_142821_(_087362_, _087363_, _087364_);
  not g_142822_(_087364_, _087365_);
  or g_142823_(_084467_, _087364_, _087366_);
  and g_142824_(_084467_, _087364_, _087368_);
  xor g_142825_(_084467_, _087364_, _087369_);
  xor g_142826_(_084467_, _087365_, _087370_);
  or g_142827_(_084476_, _087370_, _087371_);
  xor g_142828_(_084472_, _087369_, _087372_);
  and g_142829_(_084476_, _087372_, _087373_);
  not g_142830_(_087373_, _087374_);
  and g_142831_(_087371_, _087374_, _087375_);
  or g_142832_(_081585_, _084480_, _087376_);
  and g_142833_(_084478_, _087376_, _087377_);
  xor g_142834_(_087375_, _087377_, _087379_);
  or g_142835_(_084484_, _087379_, _087380_);
  xor g_142836_(_084485_, _087379_, _087381_);
  not g_142837_(_087381_, _087382_);
  or g_142838_(_084495_, _087381_, _087383_);
  xor g_142839_(_084495_, _087381_, _087384_);
  xor g_142840_(_084495_, _087382_, _087385_);
  and g_142841_(_084499_, _087385_, _087386_);
  or g_142842_(_084500_, _087384_, _087387_);
  or g_142843_(_084499_, _087381_, _087388_);
  not g_142844_(_087388_, _087390_);
  and g_142845_(_087387_, _087388_, _087391_);
  or g_142846_(_087386_, _087390_, _087392_);
  and g_142847_(_084491_, _084504_, _087393_);
  xor g_142848_(_087391_, _087393_, _087394_);
  or g_142849_(_084506_, _087394_, _087395_);
  xor g_142850_(_084506_, _087394_, _087396_);
  not g_142851_(_087396_, _087397_);
  or g_142852_(_084512_, _087397_, _087398_);
  not g_142853_(_087398_, _087399_);
  xor g_142854_(_084512_, _087396_, _087401_);
  or g_142855_(_084523_, _087401_, _087402_);
  not g_142856_(_087402_, _087403_);
  xor g_142857_(_084511_, _087401_, _087404_);
  xor g_142858_(_084510_, _087401_, _087405_);
  and g_142859_(_084523_, _087404_, _087406_);
  or g_142860_(_084522_, _087405_, _087407_);
  and g_142861_(_087402_, _087407_, _087408_);
  or g_142862_(_087403_, _087406_, _087409_);
  or g_142863_(_087165_, _087409_, _087410_);
  xor g_142864_(_087165_, _087408_, _087412_);
  not g_142865_(_087412_, _087413_);
  or g_142866_(_087164_, _087412_, _087414_);
  xor g_142867_(_087164_, _087413_, _087415_);
  not g_142868_(_087415_, _087416_);
  and g_142869_(_084531_, _087416_, _087417_);
  or g_142870_(_084532_, _087415_, _087418_);
  xor g_142871_(_084531_, _087415_, _087419_);
  not g_142872_(_087419_, _087420_);
  and g_142873_(_084534_, _087420_, _087421_);
  not g_142874_(_087421_, _087423_);
  xor g_142875_(_084534_, _087419_, _087424_);
  or g_142876_(_084536_, _087424_, _087425_);
  xor g_142877_(_084536_, _087424_, _087426_);
  not g_142878_(_087426_, _087427_);
  or g_142879_(_075844_, _078761_, _087428_);
  or g_142880_(_081644_, _087428_, _087429_);
  or g_142881_(_084535_, _087429_, _087430_);
  or g_142882_(_087427_, _087430_, _087431_);
  not g_142883_(_087431_, _087432_);
  xor g_142884_(_087426_, _087430_, _087434_);
  or g_142885_(_087163_, _087434_, _087435_);
  xor g_142886_(_087162_, _087434_, _087436_);
  not g_142887_(_087436_, _087437_);
  or g_142888_(_084543_, _087436_, _087438_);
  xor g_142889_(_084543_, _087436_, _087439_);
  xor g_142890_(_084543_, _087437_, _087440_);
  or g_142891_(_084546_, _087440_, _087441_);
  xor g_142892_(_084546_, _087439_, _087442_);
  or g_142893_(_084554_, _087442_, _087443_);
  not g_142894_(_087443_, _087445_);
  and g_142895_(_084550_, _087442_, _087446_);
  and g_142896_(_084549_, _087439_, _087447_);
  or g_142897_(_087446_, _087447_, _087448_);
  and g_142898_(_084554_, _087448_, _087449_);
  not g_142899_(_087449_, _087450_);
  and g_142900_(_087443_, _087450_, _087451_);
  or g_142901_(_087445_, _087449_, _087452_);
  or g_142902_(_087161_, _087452_, _087453_);
  xor g_142903_(_087161_, _087451_, _087454_);
  not g_142904_(_087454_, _087456_);
  or g_142905_(_087160_, _087454_, _087457_);
  xor g_142906_(_087160_, _087456_, _087458_);
  and g_142907_(_087157_, _087458_, _087459_);
  or g_142908_(_087157_, _087458_, _087460_);
  not g_142909_(_087460_, _087461_);
  or g_142910_(_087459_, _087461_, _087462_);
  not g_142911_(_087462_, _087463_);
  or g_142912_(_087156_, _087462_, _087464_);
  xor g_142913_(_087156_, _087463_, _087465_);
  not g_142914_(_087465_, _087467_);
  and g_142915_(_084560_, _084564_, _087468_);
  xor g_142916_(_087467_, _087468_, _087469_);
  or g_142917_(_084569_, _087469_, _087470_);
  xor g_142918_(_084570_, _087469_, _087471_);
  or g_142919_(_084567_, _087471_, _087472_);
  xor g_142920_(_084568_, _087471_, _087473_);
  not g_142921_(_087473_, _087474_);
  and g_142922_(_084580_, _084587_, _087475_);
  xor g_142923_(_087474_, _087475_, _087476_);
  or g_142924_(_084582_, _087476_, _087478_);
  xor g_142925_(_084583_, _087476_, _087479_);
  not g_142926_(_087479_, _087480_);
  xor g_142927_(_084593_, _087480_, _087481_);
  or g_142928_(_087154_, _087481_, _087482_);
  not g_142929_(_087482_, _087483_);
  xor g_142930_(_087155_, _087481_, _087484_);
  or g_142931_(_087153_, _087484_, _087485_);
  not g_142932_(_087485_, _087486_);
  xor g_142933_(_087153_, _087484_, _087487_);
  not g_142934_(_087487_, _087489_);
  or g_142935_(_084600_, _087489_, _087490_);
  not g_142936_(_087490_, _087491_);
  xor g_142937_(_084600_, _087487_, _087492_);
  or g_142938_(_087151_, _087492_, _087493_);
  xor g_142939_(_087152_, _087492_, _087494_);
  not g_142940_(_087494_, _087495_);
  or g_142941_(_081716_, _084602_, _087496_);
  not g_142942_(_087496_, _087497_);
  and g_142943_(_084606_, _087496_, _087498_);
  not g_142944_(_087498_, _087500_);
  xor g_142945_(_087494_, _087500_, _087501_);
  or g_142946_(_084609_, _087501_, _087502_);
  not g_142947_(_087502_, _087503_);
  and g_142948_(_084609_, _087501_, _087504_);
  xor g_142949_(_084609_, _087501_, _087505_);
  not g_142950_(_087505_, _087506_);
  and g_142951_(_084613_, _087506_, _087507_);
  or g_142952_(_084613_, _087504_, _087508_);
  or g_142953_(_087503_, _087508_, _087509_);
  not g_142954_(_087509_, _087511_);
  or g_142955_(_087507_, _087511_, _087512_);
  or g_142956_(_084612_, _087512_, _087513_);
  and g_142957_(_084612_, _087512_, _087514_);
  xor g_142958_(_084612_, _087512_, _087515_);
  xor g_142959_(_084620_, _087515_, _087516_);
  or g_142960_(_081744_, _084625_, _087517_);
  not g_142961_(_087517_, _087518_);
  or g_142962_(_084623_, _087518_, _087519_);
  xor g_142963_(_087516_, _087519_, _087520_);
  or g_142964_(_081747_, _084625_, _087522_);
  and g_142965_(_084631_, _087522_, _087523_);
  xor g_142966_(_087520_, _087523_, _087524_);
  and g_142967_(_087150_, _087524_, _087525_);
  xor g_142968_(_087149_, _087524_, _087526_);
  and g_142969_(_087148_, _087526_, _087527_);
  or g_142970_(_087148_, _087526_, _087528_);
  xor g_142971_(_087148_, _087526_, _087529_);
  and g_142972_(_084636_, _084641_, _087530_);
  xor g_142973_(_087529_, _087530_, _087531_);
  or g_142974_(_084646_, _087531_, _087533_);
  xor g_142975_(_084646_, _087531_, _087534_);
  not g_142976_(_087534_, _087535_);
  or g_142977_(_084647_, _087535_, _087536_);
  xor g_142978_(_084647_, _087534_, _087537_);
  or g_142979_(_084653_, _087537_, _087538_);
  not g_142980_(_087538_, _087539_);
  xor g_142981_(_084654_, _087537_, _087540_);
  or g_142982_(_084658_, _084660_, _087541_);
  and g_142983_(_084657_, _087541_, _087542_);
  not g_142984_(_087542_, _087544_);
  or g_142985_(_087540_, _087542_, _087545_);
  xor g_142986_(_087540_, _087544_, _087546_);
  and g_142987_(_087146_, _087546_, _087547_);
  or g_142988_(_087146_, _087546_, _087548_);
  not g_142989_(_087548_, _087549_);
  xor g_142990_(_087146_, _087546_, _087550_);
  or g_142991_(_087547_, _087549_, _087551_);
  or g_142992_(_087145_, _087551_, _087552_);
  xor g_142993_(_087145_, _087550_, _087553_);
  or g_142994_(_087143_, _087553_, _087555_);
  xor g_142995_(_087144_, _087553_, _087556_);
  and g_142996_(_084666_, _084668_, _087557_);
  not g_142997_(_087557_, _087558_);
  or g_142998_(_087556_, _087557_, _087559_);
  xor g_142999_(_087556_, _087557_, _087560_);
  xor g_143000_(_087556_, _087558_, _087561_);
  or g_143001_(_084676_, _087561_, _087562_);
  or g_143002_(_084671_, _087560_, _087563_);
  or g_143003_(_084675_, _087563_, _087564_);
  or g_143004_(_084670_, _087561_, _087566_);
  not g_143005_(_087566_, _087567_);
  and g_143006_(_087564_, _087566_, _087568_);
  and g_143007_(_087562_, _087568_, _087569_);
  not g_143008_(_087569_, _087570_);
  and g_143009_(_084679_, _084681_, _087571_);
  not g_143010_(_087571_, _087572_);
  and g_143011_(_087569_, _087572_, _087573_);
  or g_143012_(_087570_, _087571_, _087574_);
  xor g_143013_(_087569_, _087571_, _087575_);
  and g_143014_(_084685_, _084688_, _087577_);
  xor g_143015_(_087575_, _087577_, _087578_);
  not g_143016_(_087578_, _087579_);
  or g_143017_(_087142_, _087579_, _087580_);
  not g_143018_(_087580_, _087581_);
  xor g_143019_(_087142_, _087578_, _087582_);
  or g_143020_(_087140_, _087582_, _087583_);
  xor g_143021_(_087140_, _087582_, _087584_);
  xor g_143022_(_087141_, _087582_, _087585_);
  and g_143023_(_084694_, _087585_, _087586_);
  and g_143024_(_087138_, _087586_, _087588_);
  and g_143025_(_084696_, _087584_, _087589_);
  or g_143026_(_084694_, _087585_, _087590_);
  and g_143027_(_087139_, _087584_, _087591_);
  or g_143028_(_087138_, _087585_, _087592_);
  or g_143029_(_087589_, _087591_, _087593_);
  or g_143030_(_087588_, _087593_, _087594_);
  not g_143031_(_087594_, _087595_);
  or g_143032_(_087137_, _087594_, _087596_);
  xor g_143033_(_087137_, _087594_, _087597_);
  xor g_143034_(_087137_, _087595_, _087599_);
  xor g_143035_(_084704_, _087597_, _087600_);
  not g_143036_(_087600_, _087601_);
  or g_143037_(_084708_, _087600_, _087602_);
  not g_143038_(_087602_, _087603_);
  xor g_143039_(_084708_, _087600_, _087604_);
  and g_143040_(_084710_, _084714_, _087605_);
  xor g_143041_(_087604_, _087605_, _087606_);
  not g_143042_(_087606_, _087607_);
  and g_143043_(_084716_, _087607_, _087608_);
  not g_143044_(_087608_, _087610_);
  xor g_143045_(_084716_, _087606_, _087611_);
  not g_143046_(_087611_, _087612_);
  and g_143047_(_084722_, _087612_, _087613_);
  not g_143048_(_087613_, _087614_);
  or g_143049_(_084722_, _087612_, _087615_);
  not g_143050_(_087615_, _087616_);
  xor g_143051_(_084722_, _087611_, _087617_);
  and g_143052_(_084726_, _084729_, _087618_);
  or g_143053_(_087617_, _087618_, _087619_);
  xor g_143054_(_087617_, _087618_, _087621_);
  not g_143055_(_087621_, _087622_);
  and g_143056_(_087135_, _087621_, _087623_);
  not g_143057_(_087623_, _087624_);
  xor g_143058_(_087134_, _087621_, _087625_);
  or g_143059_(_087132_, _087625_, _087626_);
  xor g_143060_(_087133_, _087625_, _087627_);
  not g_143061_(_087627_, _087628_);
  and g_143062_(_084732_, _087628_, _087629_);
  or g_143063_(_084731_, _087627_, _087630_);
  xor g_143064_(_084731_, _087627_, _087632_);
  and g_143065_(_084736_, _087632_, _087633_);
  not g_143066_(_087633_, _087634_);
  xor g_143067_(_084735_, _087632_, _087635_);
  or g_143068_(_084741_, _087635_, _087636_);
  xor g_143069_(_084741_, _087635_, _087637_);
  xor g_143070_(_084742_, _087635_, _087638_);
  and g_143071_(_084745_, _087638_, _087639_);
  and g_143072_(_084751_, _087639_, _087640_);
  and g_143073_(_084749_, _087637_, _087641_);
  or g_143074_(_084751_, _087638_, _087643_);
  and g_143075_(_084746_, _087637_, _087644_);
  or g_143076_(_084745_, _087638_, _087645_);
  or g_143077_(_087641_, _087644_, _087646_);
  or g_143078_(_087640_, _087646_, _087647_);
  or g_143079_(_084754_, _087647_, _087648_);
  xor g_143080_(_084754_, _087647_, _087649_);
  not g_143081_(_087649_, _087650_);
  or g_143082_(_087131_, _087650_, _087651_);
  not g_143083_(_087651_, _087652_);
  xor g_143084_(_087131_, _087649_, _087654_);
  not g_143085_(_087654_, _087655_);
  or g_143086_(_087130_, _087654_, _087656_);
  xor g_143087_(_087130_, _087654_, _087657_);
  xor g_143088_(_087130_, _087655_, _087658_);
  or g_143089_(_087129_, _087658_, _087659_);
  xor g_143090_(_087129_, _087657_, _087660_);
  or g_143091_(_087127_, _087660_, _087661_);
  xor g_143092_(_087127_, _087660_, _087662_);
  xor g_143093_(_087128_, _087660_, _087663_);
  and g_143094_(_084764_, _087663_, _087665_);
  and g_143095_(_087124_, _087665_, _087666_);
  and g_143096_(_087126_, _087662_, _087667_);
  not g_143097_(_087667_, _087668_);
  and g_143098_(_084765_, _087662_, _087669_);
  or g_143099_(_084764_, _087663_, _087670_);
  or g_143100_(_087667_, _087669_, _087671_);
  or g_143101_(_087666_, _087671_, _087672_);
  or g_143102_(_087122_, _087672_, _087673_);
  xor g_143103_(_087122_, _087672_, _087674_);
  xor g_143104_(_087123_, _087672_, _087676_);
  or g_143105_(_087121_, _087676_, _087677_);
  and g_143106_(_087121_, _087676_, _087678_);
  xor g_143107_(_087121_, _087674_, _087679_);
  not g_143108_(_087679_, _087680_);
  and g_143109_(_087119_, _087680_, _087681_);
  xor g_143110_(_087119_, _087679_, _087682_);
  not g_143111_(_087682_, _087683_);
  and g_143112_(_084776_, _084779_, _087684_);
  xor g_143113_(_087683_, _087684_, _087685_);
  or g_143114_(_084781_, _087685_, _087687_);
  and g_143115_(_084781_, _087685_, _087688_);
  xor g_143116_(_084781_, _087685_, _087689_);
  xor g_143117_(_084782_, _087685_, _087690_);
  and g_143118_(_084784_, _084790_, _087691_);
  xor g_143119_(_087689_, _087691_, _087692_);
  or g_143120_(_084788_, _087692_, _087693_);
  xor g_143121_(_084788_, _087692_, _087694_);
  xor g_143122_(_084789_, _087692_, _087695_);
  or g_143123_(_087118_, _087695_, _087696_);
  xor g_143124_(_087118_, _087694_, _087698_);
  not g_143125_(_087698_, _087699_);
  or g_143126_(_087117_, _087698_, _087700_);
  xor g_143127_(_087117_, _087699_, _087701_);
  and g_143128_(_084800_, _084803_, _087702_);
  not g_143129_(_087702_, _087703_);
  or g_143130_(_087701_, _087702_, _087704_);
  xor g_143131_(_087701_, _087702_, _087705_);
  xor g_143132_(_087701_, _087703_, _087706_);
  or g_143133_(_087116_, _087706_, _087707_);
  xor g_143134_(_087116_, _087705_, _087709_);
  or g_143135_(_087113_, _087709_, _087710_);
  xor g_143136_(_087113_, _087709_, _087711_);
  xor g_143137_(_087115_, _087709_, _087712_);
  or g_143138_(_081942_, _084811_, _087713_);
  and g_143139_(_084814_, _087713_, _087714_);
  xor g_143140_(_087711_, _087714_, _087715_);
  or g_143141_(_084822_, _087715_, _087716_);
  not g_143142_(_087716_, _087717_);
  and g_143143_(_084819_, _087715_, _087718_);
  and g_143144_(_084822_, _087718_, _087720_);
  or g_143145_(_084819_, _087715_, _087721_);
  not g_143146_(_087721_, _087722_);
  or g_143147_(_087720_, _087722_, _087723_);
  or g_143148_(_087717_, _087723_, _087724_);
  or g_143149_(_087111_, _087724_, _087725_);
  not g_143150_(_087725_, _087726_);
  xor g_143151_(_087112_, _087724_, _087727_);
  not g_143152_(_087727_, _087728_);
  or g_143153_(_087109_, _087727_, _087729_);
  xor g_143154_(_087109_, _087727_, _087731_);
  xor g_143155_(_087109_, _087728_, _087732_);
  and g_143156_(_087107_, _087731_, _087733_);
  or g_143157_(_087106_, _087732_, _087734_);
  xor g_143158_(_087107_, _087731_, _087735_);
  not g_143159_(_087735_, _087736_);
  and g_143160_(_087105_, _087735_, _087737_);
  or g_143161_(_087104_, _087736_, _087738_);
  xor g_143162_(_087104_, _087735_, _087739_);
  and g_143163_(_084829_, _084832_, _087740_);
  xor g_143164_(_087739_, _087740_, _087742_);
  not g_143165_(_087742_, _087743_);
  or g_143166_(_084834_, _087743_, _087744_);
  not g_143167_(_087744_, _087745_);
  xor g_143168_(_084834_, _087742_, _087746_);
  not g_143169_(_087746_, _087747_);
  and g_143170_(_084837_, _084841_, _087748_);
  xor g_143171_(_087747_, _087748_, _087749_);
  or g_143172_(_084843_, _087749_, _087750_);
  and g_143173_(_084843_, _087749_, _087751_);
  xor g_143174_(_084843_, _087749_, _087753_);
  xor g_143175_(_084844_, _087749_, _087754_);
  and g_143176_(_084845_, _084851_, _087755_);
  xor g_143177_(_087753_, _087755_, _087756_);
  xor g_143178_(_084855_, _087756_, _087757_);
  not g_143179_(_087757_, _087758_);
  or g_143180_(_084858_, _087758_, _087759_);
  xor g_143181_(_084858_, _087758_, _087760_);
  and g_143182_(_084862_, _084865_, _087761_);
  not g_143183_(_087761_, _087762_);
  and g_143184_(_087760_, _087762_, _087764_);
  not g_143185_(_087764_, _087765_);
  xor g_143186_(_087760_, _087761_, _087766_);
  xor g_143187_(_084868_, _087766_, _087767_);
  or g_143188_(_087102_, _087767_, _087768_);
  xor g_143189_(_087102_, _087767_, _087769_);
  not g_143190_(_087769_, _087770_);
  or g_143191_(_087101_, _087770_, _087771_);
  xor g_143192_(_087101_, _087770_, _087772_);
  xor g_143193_(_087101_, _087769_, _087773_);
  or g_143194_(_087100_, _087773_, _087775_);
  xor g_143195_(_087100_, _087772_, _087776_);
  or g_143196_(_082047_, _084879_, _087777_);
  or g_143197_(_082050_, _084879_, _087778_);
  and g_143198_(_087777_, _087778_, _087779_);
  not g_143199_(_087779_, _087780_);
  xor g_143200_(_087776_, _087780_, _087781_);
  xor g_143201_(_087099_, _087781_, _087782_);
  not g_143202_(_087782_, _087783_);
  or g_143203_(_084887_, _087783_, _087784_);
  xor g_143204_(_084887_, _087782_, _087786_);
  not g_143205_(_087786_, _087787_);
  or g_143206_(_084891_, _087786_, _087788_);
  xor g_143207_(_084891_, _087786_, _087789_);
  xor g_143208_(_084891_, _087787_, _087790_);
  or g_143209_(_087098_, _087790_, _087791_);
  xor g_143210_(_087098_, _087789_, _087792_);
  or g_143211_(_087097_, _087792_, _087793_);
  not g_143212_(_087793_, _087794_);
  xor g_143213_(_087096_, _087792_, _087795_);
  or g_143214_(_087095_, _087795_, _087797_);
  xor g_143215_(_087095_, _087795_, _087798_);
  and g_143216_(_087094_, _087798_, _087799_);
  not g_143217_(_087799_, _087800_);
  xor g_143218_(_087094_, _087798_, _087801_);
  xor g_143219_(_087093_, _087798_, _087802_);
  and g_143220_(_084901_, _084905_, _087803_);
  xor g_143221_(_087801_, _087803_, _087804_);
  not g_143222_(_087804_, _087805_);
  or g_143223_(_087091_, _087804_, _087806_);
  xor g_143224_(_087091_, _087804_, _087808_);
  xor g_143225_(_087091_, _087805_, _087809_);
  or g_143226_(_087088_, _087809_, _087810_);
  xor g_143227_(_087088_, _087808_, _087811_);
  not g_143228_(_087811_, _087812_);
  or g_143229_(_084908_, _087811_, _087813_);
  xor g_143230_(_084908_, _087811_, _087814_);
  xor g_143231_(_084908_, _087812_, _087815_);
  and g_143232_(_084910_, _084912_, _087816_);
  xor g_143233_(_087814_, _087816_, _087817_);
  or g_143234_(_084914_, _087817_, _087819_);
  xor g_143235_(_084916_, _087817_, _087820_);
  not g_143236_(_087820_, _087821_);
  or g_143237_(_087086_, _087820_, _087822_);
  xor g_143238_(_087086_, _087820_, _087823_);
  xor g_143239_(_087086_, _087821_, _087824_);
  or g_143240_(_087084_, _087824_, _087825_);
  and g_143241_(_087084_, _087824_, _087826_);
  or g_143242_(_087085_, _087823_, _087827_);
  and g_143243_(_084934_, _087827_, _087828_);
  or g_143244_(_084935_, _087826_, _087830_);
  and g_143245_(_087825_, _087828_, _087831_);
  xor g_143246_(_087084_, _087823_, _087832_);
  and g_143247_(_084935_, _087832_, _087833_);
  or g_143248_(_087831_, _087833_, _087834_);
  and g_143249_(_084933_, _087834_, _087835_);
  or g_143250_(_084933_, _087834_, _087836_);
  xor g_143251_(_084933_, _087834_, _087837_);
  xor g_143252_(_084932_, _087834_, _087838_);
  or g_143253_(_082113_, _084941_, _087839_);
  and g_143254_(_084939_, _087839_, _087841_);
  xor g_143255_(_087838_, _087841_, _087842_);
  xor g_143256_(_087837_, _087841_, _087843_);
  or g_143257_(_079196_, _082117_, _087844_);
  or g_143258_(_084943_, _087844_, _087845_);
  not g_143259_(_087845_, _087846_);
  or g_143260_(_082116_, _084941_, _087847_);
  not g_143261_(_087847_, _087848_);
  and g_143262_(_087845_, _087847_, _087849_);
  xor g_143263_(_087842_, _087849_, _087850_);
  xor g_143264_(_087843_, _087849_, _087852_);
  or g_143265_(_087083_, _087850_, _087853_);
  xor g_143266_(_087083_, _087850_, _087854_);
  xor g_143267_(_087083_, _087852_, _087855_);
  and g_143268_(_084952_, _087854_, _087856_);
  not g_143269_(_087856_, _087857_);
  and g_143270_(_084947_, _087852_, _087858_);
  or g_143271_(_084946_, _087850_, _087859_);
  and g_143272_(_084946_, _087855_, _087860_);
  or g_143273_(_087858_, _087860_, _087861_);
  not g_143274_(_087861_, _087863_);
  and g_143275_(_084951_, _087861_, _087864_);
  or g_143276_(_087856_, _087864_, _087865_);
  and g_143277_(_084954_, _087865_, _087866_);
  and g_143278_(_084955_, _087863_, _087867_);
  not g_143279_(_087867_, _087868_);
  or g_143280_(_087866_, _087867_, _087869_);
  or g_143281_(_087080_, _087869_, _087870_);
  xor g_143282_(_087080_, _087869_, _087871_);
  and g_143283_(_087079_, _087871_, _087872_);
  xor g_143284_(_087078_, _087871_, _087874_);
  not g_143285_(_087874_, _087875_);
  and g_143286_(_087076_, _087875_, _087876_);
  or g_143287_(_087077_, _087874_, _087877_);
  xor g_143288_(_087076_, _087874_, _087878_);
  or g_143289_(_087074_, _087878_, _087879_);
  xor g_143290_(_087075_, _087878_, _087880_);
  or g_143291_(_082148_, _084961_, _087881_);
  and g_143292_(_084962_, _087881_, _087882_);
  not g_143293_(_087882_, _087883_);
  xor g_143294_(_087880_, _087883_, _087885_);
  not g_143295_(_087885_, _087886_);
  xor g_143296_(_087073_, _087886_, _087887_);
  or g_143297_(_087071_, _087887_, _087888_);
  and g_143298_(_087071_, _087887_, _087889_);
  not g_143299_(_087889_, _087890_);
  and g_143300_(_087888_, _087890_, _087891_);
  not g_143301_(_087891_, _087892_);
  or g_143302_(_084968_, _084971_, _087893_);
  not g_143303_(_087893_, _087894_);
  and g_143304_(_084975_, _087893_, _087896_);
  xor g_143305_(_087891_, _087896_, _087897_);
  or g_143306_(_084980_, _087897_, _087898_);
  not g_143307_(_087898_, _087899_);
  and g_143308_(_084978_, _087897_, _087900_);
  and g_143309_(_084980_, _087900_, _087901_);
  or g_143310_(_084978_, _087897_, _087902_);
  not g_143311_(_087902_, _087903_);
  or g_143312_(_087901_, _087903_, _087904_);
  or g_143313_(_087899_, _087904_, _087905_);
  not g_143314_(_087905_, _087907_);
  and g_143315_(_084988_, _087907_, _087908_);
  not g_143316_(_087908_, _087909_);
  xor g_143317_(_084988_, _087905_, _087910_);
  or g_143318_(_084987_, _087910_, _087911_);
  not g_143319_(_087911_, _087912_);
  xor g_143320_(_084987_, _087910_, _087913_);
  xor g_143321_(_084986_, _087910_, _087914_);
  or g_143322_(_087069_, _087914_, _087915_);
  xor g_143323_(_087069_, _087913_, _087916_);
  not g_143324_(_087916_, _087918_);
  or g_143325_(_087068_, _087916_, _087919_);
  xor g_143326_(_087068_, _087918_, _087920_);
  and g_143327_(_084994_, _084998_, _087921_);
  not g_143328_(_087921_, _087922_);
  xor g_143329_(_087920_, _087922_, _087923_);
  or g_143330_(_084999_, _087923_, _087924_);
  xor g_143331_(_085000_, _087923_, _087925_);
  not g_143332_(_087925_, _087926_);
  and g_143333_(_085006_, _087926_, _087927_);
  or g_143334_(_085005_, _087925_, _087929_);
  xor g_143335_(_085006_, _087925_, _087930_);
  and g_143336_(_085009_, _085011_, _087931_);
  not g_143337_(_087931_, _087932_);
  xor g_143338_(_087930_, _087932_, _087933_);
  not g_143339_(_087933_, _087934_);
  xor g_143340_(_087067_, _087933_, _087935_);
  xor g_143341_(_087067_, _087934_, _087936_);
  or g_143342_(_087064_, _087936_, _087937_);
  not g_143343_(_087937_, _087938_);
  xor g_143344_(_087064_, _087935_, _087940_);
  not g_143345_(_087940_, _087941_);
  and g_143346_(_085018_, _087941_, _087942_);
  xor g_143347_(_085018_, _087940_, _087943_);
  and g_143348_(_085020_, _085022_, _087944_);
  and g_143349_(_087943_, _087944_, _087945_);
  not g_143350_(_087945_, _087946_);
  or g_143351_(_085022_, _087943_, _087947_);
  not g_143352_(_087947_, _087948_);
  or g_143353_(_085020_, _087940_, _087949_);
  not g_143354_(_087949_, _087951_);
  and g_143355_(_087947_, _087949_, _087952_);
  not g_143356_(_087952_, _087953_);
  and g_143357_(_087946_, _087952_, _087954_);
  or g_143358_(_087945_, _087953_, _087955_);
  or g_143359_(_085032_, _087955_, _087956_);
  xor g_143360_(_085032_, _087954_, _087957_);
  or g_143361_(_085026_, _087957_, _087958_);
  xor g_143362_(_085027_, _087957_, _087959_);
  or g_143363_(_085048_, _087959_, _087960_);
  xor g_143364_(_085049_, _087959_, _087962_);
  or g_143365_(_085045_, _087962_, _087963_);
  not g_143366_(_087963_, _087964_);
  xor g_143367_(_085046_, _087962_, _087965_);
  and g_143368_(_085054_, _085056_, _087966_);
  not g_143369_(_087966_, _087967_);
  xor g_143370_(_087965_, _087967_, _087968_);
  or g_143371_(_085060_, _087968_, _087969_);
  xor g_143372_(_085061_, _087968_, _087970_);
  and g_143373_(_085064_, _087970_, _087971_);
  or g_143374_(_085064_, _087970_, _087973_);
  xor g_143375_(_085065_, _087970_, _087974_);
  or g_143376_(_082258_, _085068_, _087975_);
  and g_143377_(_085067_, _087975_, _087976_);
  not g_143378_(_087976_, _087977_);
  xor g_143379_(_087974_, _087977_, _087978_);
  or g_143380_(_087062_, _087978_, _087979_);
  xor g_143381_(_087063_, _087978_, _087980_);
  or g_143382_(_085073_, _087980_, _087981_);
  or g_143383_(_085076_, _087980_, _087982_);
  xor g_143384_(_085076_, _087980_, _087984_);
  or g_143385_(_085074_, _087984_, _087985_);
  and g_143386_(_087981_, _087985_, _087986_);
  and g_143387_(_085079_, _087986_, _087987_);
  not g_143388_(_087987_, _087988_);
  and g_143389_(_085083_, _087986_, _087989_);
  not g_143390_(_087989_, _087990_);
  xor g_143391_(_085083_, _087986_, _087991_);
  xor g_143392_(_085082_, _087986_, _087992_);
  and g_143393_(_085078_, _087992_, _087993_);
  or g_143394_(_085079_, _087991_, _087995_);
  and g_143395_(_087988_, _087995_, _087996_);
  or g_143396_(_087987_, _087993_, _087997_);
  and g_143397_(_085093_, _087996_, _087998_);
  not g_143398_(_087998_, _087999_);
  and g_143399_(_085086_, _085092_, _088000_);
  and g_143400_(_087997_, _088000_, _088001_);
  and g_143401_(_085087_, _087996_, _088002_);
  or g_143402_(_085086_, _087997_, _088003_);
  or g_143403_(_088001_, _088002_, _088004_);
  or g_143404_(_087998_, _088004_, _088006_);
  or g_143405_(_085096_, _088006_, _088007_);
  xor g_143406_(_085096_, _088006_, _088008_);
  and g_143407_(_085103_, _085107_, _088009_);
  xor g_143408_(_088008_, _088009_, _088010_);
  xor g_143409_(_087061_, _088010_, _088011_);
  xor g_143410_(_087058_, _088011_, _088012_);
  and g_143411_(_087055_, _088012_, _088013_);
  not g_143412_(_088013_, _088014_);
  or g_143413_(_082303_, _085123_, _088015_);
  not g_143414_(_088015_, _088017_);
  or g_143415_(_087055_, _088012_, _088018_);
  and g_143416_(_088017_, _088018_, _088019_);
  not g_143417_(_088019_, _088020_);
  and g_143418_(_088014_, _088019_, _088021_);
  xor g_143419_(_087056_, _088012_, _088022_);
  and g_143420_(_088015_, _088022_, _088023_);
  or g_143421_(_088021_, _088023_, _088024_);
  or g_143422_(_087054_, _088024_, _088025_);
  xor g_143423_(_087054_, _088024_, _088026_);
  not g_143424_(_088026_, _088028_);
  or g_143425_(_087053_, _088028_, _088029_);
  xor g_143426_(_087053_, _088026_, _088030_);
  or g_143427_(_087051_, _088030_, _088031_);
  xor g_143428_(_087052_, _088030_, _088032_);
  or g_143429_(_085134_, _088032_, _088033_);
  and g_143430_(_085134_, _088032_, _088034_);
  xor g_143431_(_085136_, _088032_, _088035_);
  and g_143432_(_085139_, _085142_, _088036_);
  not g_143433_(_088036_, _088037_);
  xor g_143434_(_088035_, _088037_, _088039_);
  or g_143435_(_085144_, _088039_, _088040_);
  xor g_143436_(_085144_, _088039_, _088041_);
  xor g_143437_(_085145_, _088039_, _088042_);
  and g_143438_(_085149_, _088042_, _088043_);
  and g_143439_(_085152_, _088043_, _088044_);
  and g_143440_(_085150_, _088041_, _088045_);
  or g_143441_(_085149_, _088042_, _088046_);
  and g_143442_(_085153_, _088041_, _088047_);
  or g_143443_(_085152_, _088042_, _088048_);
  or g_143444_(_088045_, _088047_, _088050_);
  or g_143445_(_088044_, _088050_, _088051_);
  or g_143446_(_085155_, _088051_, _088052_);
  xor g_143447_(_085156_, _088051_, _088053_);
  or g_143448_(_087050_, _088053_, _088054_);
  xor g_143449_(_087049_, _088053_, _088055_);
  or g_143450_(_087046_, _088055_, _088056_);
  and g_143451_(_087046_, _088055_, _088057_);
  xor g_143452_(_087047_, _088055_, _088058_);
  or g_143453_(_087044_, _088058_, _088059_);
  xor g_143454_(_087045_, _088058_, _088061_);
  or g_143455_(_087043_, _088061_, _088062_);
  xor g_143456_(_087043_, _088061_, _088063_);
  xor g_143457_(_085176_, _088063_, _088064_);
  not g_143458_(_088064_, _088065_);
  or g_143459_(_085178_, _088064_, _088066_);
  or g_143460_(_085182_, _088066_, _088067_);
  or g_143461_(_085183_, _088065_, _088068_);
  and g_143462_(_085178_, _088063_, _088069_);
  not g_143463_(_088069_, _088070_);
  and g_143464_(_088068_, _088070_, _088072_);
  and g_143465_(_088067_, _088072_, _088073_);
  not g_143466_(_088073_, _088074_);
  or g_143467_(_087042_, _088074_, _088075_);
  xor g_143468_(_087042_, _088073_, _088076_);
  or g_143469_(_087040_, _088076_, _088077_);
  xor g_143470_(_087041_, _088076_, _088078_);
  or g_143471_(_085191_, _088078_, _088079_);
  xor g_143472_(_085192_, _088078_, _088080_);
  and g_143473_(_087039_, _088080_, _088081_);
  or g_143474_(_087039_, _088080_, _088083_);
  not g_143475_(_088083_, _088084_);
  xor g_143476_(_087039_, _088080_, _088085_);
  or g_143477_(_088081_, _088084_, _088086_);
  or g_143478_(_087038_, _088086_, _088087_);
  xor g_143479_(_087038_, _088085_, _088088_);
  or g_143480_(_087035_, _088088_, _088089_);
  xor g_143481_(_087036_, _088088_, _088090_);
  not g_143482_(_088090_, _088091_);
  or g_143483_(_087034_, _088090_, _088092_);
  xor g_143484_(_087034_, _088090_, _088094_);
  xor g_143485_(_087034_, _088091_, _088095_);
  or g_143486_(_085200_, _088095_, _088096_);
  xor g_143487_(_085200_, _088094_, _088097_);
  or g_143488_(_085203_, _088097_, _088098_);
  and g_143489_(_085203_, _088097_, _088099_);
  xor g_143490_(_085203_, _088097_, _088100_);
  xor g_143491_(_085207_, _088100_, _088101_);
  xor g_143492_(_087033_, _088101_, _088102_);
  not g_143493_(_088102_, _088103_);
  or g_143494_(_087031_, _088103_, _088105_);
  not g_143495_(_088105_, _088106_);
  xor g_143496_(_087031_, _088102_, _088107_);
  not g_143497_(_088107_, _088108_);
  and g_143498_(_085215_, _085218_, _088109_);
  xor g_143499_(_088107_, _088109_, _088110_);
  xor g_143500_(_088108_, _088109_, _088111_);
  or g_143501_(_085222_, _088111_, _088112_);
  xor g_143502_(_085222_, _088110_, _088113_);
  not g_143503_(_088113_, _088114_);
  or g_143504_(_085225_, _088113_, _088116_);
  xor g_143505_(_085225_, _088114_, _088117_);
  or g_143506_(_085227_, _088117_, _088118_);
  not g_143507_(_088118_, _088119_);
  and g_143508_(_085227_, _088117_, _088120_);
  or g_143509_(_088119_, _088120_, _088121_);
  not g_143510_(_088121_, _088122_);
  and g_143511_(_085229_, _085231_, _088123_);
  xor g_143512_(_088122_, _088123_, _088124_);
  not g_143513_(_088124_, _088125_);
  and g_143514_(_085233_, _085240_, _088127_);
  xor g_143515_(_088125_, _088127_, _088128_);
  or g_143516_(_085236_, _088128_, _088129_);
  not g_143517_(_088129_, _088130_);
  xor g_143518_(_085236_, _088128_, _088131_);
  xor g_143519_(_085237_, _088128_, _088132_);
  and g_143520_(_082427_, _082432_, _088133_);
  or g_143521_(_085243_, _088133_, _088134_);
  or g_143522_(_088132_, _088134_, _088135_);
  xor g_143523_(_088131_, _088134_, _088136_);
  or g_143524_(_087030_, _088136_, _088138_);
  xor g_143525_(_087030_, _088136_, _088139_);
  not g_143526_(_088139_, _088140_);
  or g_143527_(_085247_, _088140_, _088141_);
  not g_143528_(_088141_, _088142_);
  xor g_143529_(_085247_, _088139_, _088143_);
  or g_143530_(_085250_, _088143_, _088144_);
  not g_143531_(_088144_, _088145_);
  xor g_143532_(_085250_, _088143_, _088146_);
  and g_143533_(_085253_, _088146_, _088147_);
  not g_143534_(_088147_, _088149_);
  xor g_143535_(_085252_, _088146_, _088150_);
  not g_143536_(_088150_, _088151_);
  and g_143537_(_085261_, _088151_, _088152_);
  not g_143538_(_088152_, _088153_);
  xor g_143539_(_085261_, _088150_, _088154_);
  or g_143540_(_085260_, _088154_, _088155_);
  xor g_143541_(_085259_, _088154_, _088156_);
  not g_143542_(_088156_, _088157_);
  and g_143543_(_085264_, _085266_, _088158_);
  xor g_143544_(_088157_, _088158_, _088160_);
  not g_143545_(_088160_, _088161_);
  and g_143546_(_087029_, _088161_, _088162_);
  not g_143547_(_088162_, _088163_);
  xor g_143548_(_087028_, _088160_, _088164_);
  and g_143549_(_085279_, _088164_, _088165_);
  xor g_143550_(_085280_, _088164_, _088166_);
  not g_143551_(_088166_, _088167_);
  and g_143552_(_085281_, _088167_, _088168_);
  xor g_143553_(_085281_, _088166_, _088169_);
  or g_143554_(_085284_, _088169_, _088171_);
  not g_143555_(_088171_, _088172_);
  or g_143556_(_079515_, _082473_, _088173_);
  or g_143557_(_085283_, _088173_, _088174_);
  not g_143558_(_088174_, _088175_);
  or g_143559_(_088169_, _088174_, _088176_);
  xor g_143560_(_088169_, _088174_, _088177_);
  xor g_143561_(_088169_, _088175_, _088178_);
  and g_143562_(_085284_, _088178_, _088179_);
  or g_143563_(_085285_, _088177_, _088180_);
  and g_143564_(_088171_, _088180_, _088182_);
  or g_143565_(_088172_, _088179_, _088183_);
  or g_143566_(_087027_, _088183_, _088184_);
  xor g_143567_(_087027_, _088182_, _088185_);
  not g_143568_(_088185_, _088186_);
  or g_143569_(_087024_, _088185_, _088187_);
  xor g_143570_(_087024_, _088186_, _088188_);
  not g_143571_(_088188_, _088189_);
  or g_143572_(_087022_, _088188_, _088190_);
  xor g_143573_(_087022_, _088189_, _088191_);
  or g_143574_(_085295_, _088191_, _088193_);
  xor g_143575_(_085296_, _088191_, _088194_);
  or g_143576_(_085297_, _088194_, _088195_);
  xor g_143577_(_085297_, _088194_, _088196_);
  xor g_143578_(_085298_, _088194_, _088197_);
  or g_143579_(_085304_, _088197_, _088198_);
  xor g_143580_(_085304_, _088196_, _088199_);
  or g_143581_(_085306_, _088199_, _088200_);
  xor g_143582_(_085307_, _088199_, _088201_);
  and g_143583_(_085309_, _085314_, _088202_);
  xor g_143584_(_088201_, _088202_, _088204_);
  xor g_143585_(_085321_, _088204_, _088205_);
  not g_143586_(_088205_, _088206_);
  and g_143587_(_085328_, _088206_, _088207_);
  xor g_143588_(_085327_, _088205_, _088208_);
  and g_143589_(_085331_, _088208_, _088209_);
  xor g_143590_(_085330_, _088208_, _088210_);
  or g_143591_(_085340_, _085352_, _088211_);
  xor g_143592_(_088210_, _088211_, _088212_);
  or g_143593_(_085351_, _088212_, _088213_);
  xor g_143594_(_085351_, _088212_, _088215_);
  and g_143595_(_085358_, _088215_, _088216_);
  not g_143596_(_088216_, _088217_);
  and g_143597_(_085362_, _088215_, _088218_);
  xor g_143598_(_085361_, _088215_, _088219_);
  and g_143599_(_085359_, _088219_, _088220_);
  or g_143600_(_088216_, _088220_, _088221_);
  not g_143601_(_088221_, _088222_);
  and g_143602_(_085371_, _088222_, _088223_);
  xor g_143603_(_085371_, _088221_, _088224_);
  not g_143604_(_088224_, _088226_);
  and g_143605_(_085368_, _088226_, _088227_);
  or g_143606_(_085367_, _088224_, _088228_);
  xor g_143607_(_085368_, _088224_, _088229_);
  and g_143608_(_087020_, _088229_, _088230_);
  or g_143609_(_087020_, _088229_, _088231_);
  not g_143610_(_088231_, _088232_);
  xor g_143611_(_087020_, _088229_, _088233_);
  or g_143612_(_088230_, _088232_, _088234_);
  or g_143613_(_087019_, _088234_, _088235_);
  xor g_143614_(_087019_, _088233_, _088237_);
  or g_143615_(_085381_, _088237_, _088238_);
  xor g_143616_(_085380_, _088237_, _088239_);
  and g_143617_(_087018_, _088239_, _088240_);
  or g_143618_(_087018_, _088239_, _088241_);
  not g_143619_(_088241_, _088242_);
  xor g_143620_(_087018_, _088239_, _088243_);
  or g_143621_(_088240_, _088242_, _088244_);
  or g_143622_(_087017_, _088244_, _088245_);
  xor g_143623_(_087017_, _088243_, _088246_);
  not g_143624_(_088246_, _088248_);
  or g_143625_(_087016_, _088246_, _088249_);
  xor g_143626_(_087016_, _088248_, _088250_);
  or g_143627_(_087013_, _088250_, _088251_);
  xor g_143628_(_087014_, _088250_, _088252_);
  not g_143629_(_088252_, _088253_);
  and g_143630_(_085389_, _085393_, _088254_);
  or g_143631_(_085387_, _085392_, _088255_);
  and g_143632_(_088253_, _088255_, _088256_);
  xor g_143633_(_088252_, _088254_, _088257_);
  and g_143634_(_085401_, _088257_, _088259_);
  xor g_143635_(_085402_, _088257_, _088260_);
  not g_143636_(_088260_, _088261_);
  and g_143637_(_085403_, _088261_, _088262_);
  xor g_143638_(_085404_, _088260_, _088263_);
  xor g_143639_(_085403_, _088260_, _088264_);
  and g_143640_(_085409_, _085412_, _088265_);
  xor g_143641_(_088263_, _088265_, _088266_);
  or g_143642_(_085418_, _088266_, _088267_);
  not g_143643_(_088267_, _088268_);
  or g_143644_(_085414_, _088266_, _088270_);
  xor g_143645_(_085415_, _088266_, _088271_);
  or g_143646_(_085422_, _088271_, _088272_);
  xor g_143647_(_085423_, _088271_, _088273_);
  and g_143648_(_085418_, _088273_, _088274_);
  or g_143649_(_088268_, _088274_, _088275_);
  and g_143650_(_085426_, _085428_, _088276_);
  not g_143651_(_088276_, _088277_);
  or g_143652_(_088275_, _088276_, _088278_);
  xor g_143653_(_088275_, _088276_, _088279_);
  xor g_143654_(_088275_, _088277_, _088281_);
  and g_143655_(_087010_, _088279_, _088282_);
  or g_143656_(_087011_, _088281_, _088283_);
  or g_143657_(_087010_, _088279_, _088284_);
  not g_143658_(_088284_, _088285_);
  xor g_143659_(_087010_, _088279_, _088286_);
  or g_143660_(_088282_, _088285_, _088287_);
  or g_143661_(_085430_, _085431_, _088288_);
  not g_143662_(_088288_, _088289_);
  or g_143663_(_084100_, _085434_, _088290_);
  and g_143664_(_088288_, _088290_, _088292_);
  xor g_143665_(_088286_, _088292_, _088293_);
  or g_143666_(_087009_, _088293_, _088294_);
  xor g_143667_(_087009_, _088293_, _088295_);
  and g_143668_(_085441_, _088295_, _088296_);
  not g_143669_(_088296_, _088297_);
  xor g_143670_(_085441_, _088295_, _088298_);
  and g_143671_(_085439_, _088298_, _088299_);
  xor g_143672_(_085440_, _088298_, _088300_);
  or g_143673_(_082621_, _085446_, _088301_);
  and g_143674_(_085445_, _088301_, _088303_);
  xor g_143675_(_088300_, _088303_, _088304_);
  and g_143676_(_087008_, _088304_, _088305_);
  not g_143677_(_088305_, _088306_);
  xor g_143678_(_087007_, _088304_, _088307_);
  not g_143679_(_088307_, _088308_);
  and g_143680_(_087006_, _088308_, _088309_);
  not g_143681_(_088309_, _088310_);
  xor g_143682_(_087006_, _088308_, _088311_);
  and g_143683_(_087005_, _088311_, _088312_);
  xor g_143684_(_087003_, _088311_, _088314_);
  not g_143685_(_088314_, _088315_);
  or g_143686_(_085457_, _088314_, _088316_);
  not g_143687_(_088316_, _088317_);
  and g_143688_(_085453_, _088314_, _088318_);
  and g_143689_(_085457_, _088318_, _088319_);
  and g_143690_(_085452_, _088315_, _088320_);
  not g_143691_(_088320_, _088321_);
  or g_143692_(_088319_, _088320_, _088322_);
  or g_143693_(_088317_, _088322_, _088323_);
  or g_143694_(_085468_, _088323_, _088325_);
  xor g_143695_(_085467_, _088323_, _088326_);
  or g_143696_(_085460_, _088326_, _088327_);
  xor g_143697_(_085461_, _088326_, _088328_);
  or g_143698_(_082642_, _085472_, _088329_);
  and g_143699_(_085473_, _088329_, _088330_);
  xor g_143700_(_088328_, _088330_, _088331_);
  and g_143701_(_087002_, _088331_, _088332_);
  xor g_143702_(_087002_, _088331_, _088333_);
  or g_143703_(_085483_, _085492_, _088334_);
  xor g_143704_(_088333_, _088334_, _088336_);
  and g_143705_(_085490_, _088336_, _088337_);
  not g_143706_(_088337_, _088338_);
  xor g_143707_(_085490_, _088336_, _088339_);
  not g_143708_(_088339_, _088340_);
  and g_143709_(_085496_, _085499_, _088341_);
  xor g_143710_(_088339_, _088341_, _088342_);
  xor g_143711_(_088340_, _088341_, _088343_);
  and g_143712_(_085503_, _088343_, _088344_);
  or g_143713_(_085502_, _088342_, _088345_);
  xor g_143714_(_085503_, _088342_, _088347_);
  not g_143715_(_088347_, _088348_);
  and g_143716_(_085507_, _088347_, _088349_);
  and g_143717_(_085515_, _088349_, _088350_);
  and g_143718_(_085516_, _088348_, _088351_);
  not g_143719_(_088351_, _088352_);
  or g_143720_(_085507_, _088347_, _088353_);
  not g_143721_(_088353_, _088354_);
  or g_143722_(_088351_, _088354_, _088355_);
  or g_143723_(_088350_, _088355_, _088356_);
  not g_143724_(_088356_, _088358_);
  and g_143725_(_085513_, _088358_, _088359_);
  not g_143726_(_088359_, _088360_);
  xor g_143727_(_085513_, _088356_, _088361_);
  not g_143728_(_088361_, _088362_);
  and g_143729_(_085525_, _088361_, _088363_);
  and g_143730_(_085524_, _088362_, _088364_);
  or g_143731_(_085522_, _088361_, _088365_);
  not g_143732_(_088365_, _088366_);
  or g_143733_(_088364_, _088366_, _088367_);
  or g_143734_(_088363_, _088367_, _088369_);
  not g_143735_(_088369_, _088370_);
  or g_143736_(_085534_, _088369_, _088371_);
  xor g_143737_(_085534_, _088369_, _088372_);
  xor g_143738_(_085534_, _088370_, _088373_);
  or g_143739_(_085536_, _088373_, _088374_);
  xor g_143740_(_085536_, _088372_, _088375_);
  not g_143741_(_088375_, _088376_);
  or g_143742_(_085538_, _088375_, _088377_);
  and g_143743_(_085538_, _088375_, _088378_);
  xor g_143744_(_085538_, _088376_, _088380_);
  not g_143745_(_088380_, _088381_);
  or g_143746_(_082710_, _085539_, _088382_);
  and g_143747_(_085540_, _088382_, _088383_);
  xor g_143748_(_088380_, _088383_, _088384_);
  xor g_143749_(_088381_, _088383_, _088385_);
  or g_143750_(_087001_, _088385_, _088386_);
  xor g_143751_(_087001_, _088384_, _088387_);
  or g_143752_(_085547_, _088387_, _088388_);
  not g_143753_(_088388_, _088389_);
  and g_143754_(_085547_, _088387_, _088391_);
  xor g_143755_(_085547_, _088387_, _088392_);
  or g_143756_(_088389_, _088391_, _088393_);
  and g_143757_(_085549_, _088393_, _088394_);
  and g_143758_(_085552_, _088394_, _088395_);
  or g_143759_(_085549_, _088387_, _088396_);
  not g_143760_(_088396_, _088397_);
  and g_143761_(_085554_, _088392_, _088398_);
  not g_143762_(_088398_, _088399_);
  or g_143763_(_088397_, _088398_, _088400_);
  or g_143764_(_088395_, _088400_, _088402_);
  or g_143765_(_082729_, _085557_, _088403_);
  and g_143766_(_085556_, _088403_, _088404_);
  or g_143767_(_088402_, _088404_, _088405_);
  xor g_143768_(_088402_, _088404_, _088406_);
  not g_143769_(_088406_, _088407_);
  and g_143770_(_087000_, _088406_, _088408_);
  or g_143771_(_086999_, _088407_, _088409_);
  xor g_143772_(_086999_, _088406_, _088410_);
  or g_143773_(_085562_, _088410_, _088411_);
  not g_143774_(_088411_, _088413_);
  xor g_143775_(_085562_, _088410_, _088414_);
  xor g_143776_(_085563_, _088410_, _088415_);
  or g_143777_(_085567_, _088414_, _088416_);
  or g_143778_(_085571_, _088416_, _088417_);
  or g_143779_(_085568_, _088415_, _088418_);
  or g_143780_(_085572_, _088415_, _088419_);
  not g_143781_(_088419_, _088420_);
  and g_143782_(_088418_, _088419_, _088421_);
  and g_143783_(_088417_, _088421_, _088422_);
  and g_143784_(_086998_, _088422_, _088424_);
  xor g_143785_(_086997_, _088422_, _088425_);
  not g_143786_(_088425_, _088426_);
  and g_143787_(_086996_, _088426_, _088427_);
  not g_143788_(_088427_, _088428_);
  xor g_143789_(_086996_, _088426_, _088429_);
  xor g_143790_(_086996_, _088425_, _088430_);
  or g_143791_(_085578_, _088430_, _088431_);
  xor g_143792_(_085578_, _088429_, _088432_);
  or g_143793_(_085580_, _088432_, _088433_);
  xor g_143794_(_085580_, _088432_, _088435_);
  and g_143795_(_085583_, _088435_, _088436_);
  xor g_143796_(_085582_, _088435_, _088437_);
  and g_143797_(_085588_, _085591_, _088438_);
  xor g_143798_(_088437_, _088438_, _088439_);
  and g_143799_(_085593_, _088439_, _088440_);
  not g_143800_(_088440_, _088441_);
  xor g_143801_(_085594_, _088439_, _088442_);
  not g_143802_(_088442_, _088443_);
  and g_143803_(_086995_, _088443_, _088444_);
  or g_143804_(_086995_, _088443_, _088446_);
  xor g_143805_(_086995_, _088442_, _088447_);
  or g_143806_(_086991_, _088447_, _088448_);
  xor g_143807_(_086992_, _088447_, _088449_);
  or g_143808_(_086990_, _088449_, _088450_);
  not g_143809_(_088450_, _088451_);
  and g_143810_(_086990_, _088449_, _088452_);
  xor g_143811_(_086990_, _088449_, _088453_);
  or g_143812_(_088451_, _088452_, _088454_);
  or g_143813_(_086989_, _088454_, _088455_);
  xor g_143814_(_086989_, _088453_, _088457_);
  or g_143815_(_085611_, _088457_, _088458_);
  xor g_143816_(_085612_, _088457_, _088459_);
  or g_143817_(_085610_, _088459_, _088460_);
  not g_143818_(_088460_, _088461_);
  xor g_143819_(_085610_, _088459_, _088462_);
  not g_143820_(_088462_, _088463_);
  and g_143821_(_085616_, _088462_, _088464_);
  or g_143822_(_085615_, _088463_, _088465_);
  xor g_143823_(_085615_, _088462_, _088466_);
  or g_143824_(_085621_, _088466_, _088468_);
  xor g_143825_(_085620_, _088466_, _088469_);
  xor g_143826_(_085626_, _088469_, _088470_);
  xor g_143827_(_086987_, _088470_, _088471_);
  and g_143828_(_085636_, _088471_, _088472_);
  or g_143829_(_085636_, _088471_, _088473_);
  not g_143830_(_088473_, _088474_);
  xor g_143831_(_085636_, _088471_, _088475_);
  or g_143832_(_088472_, _088474_, _088476_);
  or g_143833_(_086985_, _088476_, _088477_);
  xor g_143834_(_086985_, _088475_, _088479_);
  and g_143835_(_086981_, _088479_, _088480_);
  or g_143836_(_086981_, _088479_, _088481_);
  xor g_143837_(_086983_, _088479_, _088482_);
  and g_143838_(_085639_, _085651_, _088483_);
  xor g_143839_(_088482_, _088483_, _088484_);
  and g_143840_(_085650_, _088484_, _088485_);
  xor g_143841_(_085649_, _088484_, _088486_);
  or g_143842_(_085657_, _088486_, _088487_);
  not g_143843_(_088487_, _088488_);
  xor g_143844_(_085657_, _088486_, _088490_);
  not g_143845_(_088490_, _088491_);
  and g_143846_(_085660_, _088490_, _088492_);
  or g_143847_(_085659_, _088491_, _088493_);
  xor g_143848_(_085659_, _088490_, _088494_);
  xor g_143849_(_085667_, _088494_, _088495_);
  xor g_143850_(_086979_, _088495_, _088496_);
  or g_143851_(_085677_, _088496_, _088497_);
  xor g_143852_(_085678_, _088496_, _088498_);
  not g_143853_(_088498_, _088499_);
  and g_143854_(_085683_, _085686_, _088501_);
  xor g_143855_(_088498_, _088501_, _088502_);
  xor g_143856_(_088499_, _088501_, _088503_);
  and g_143857_(_085695_, _088502_, _088504_);
  or g_143858_(_085697_, _088503_, _088505_);
  or g_143859_(_085688_, _088503_, _088506_);
  xor g_143860_(_085688_, _088502_, _088507_);
  and g_143861_(_085697_, _088507_, _088508_);
  or g_143862_(_088504_, _088508_, _088509_);
  not g_143863_(_088509_, _088510_);
  and g_143864_(_085698_, _088510_, _088512_);
  not g_143865_(_088512_, _088513_);
  xor g_143866_(_085698_, _088510_, _088514_);
  xor g_143867_(_085698_, _088509_, _088515_);
  or g_143868_(_085702_, _088515_, _088516_);
  not g_143869_(_088516_, _088517_);
  xor g_143870_(_085702_, _088515_, _088518_);
  xor g_143871_(_085702_, _088514_, _088519_);
  and g_143872_(_085704_, _088519_, _088520_);
  and g_143873_(_085709_, _088520_, _088521_);
  and g_143874_(_085710_, _088518_, _088523_);
  or g_143875_(_085709_, _088519_, _088524_);
  and g_143876_(_085705_, _088514_, _088525_);
  not g_143877_(_088525_, _088526_);
  or g_143878_(_088523_, _088525_, _088527_);
  or g_143879_(_088521_, _088527_, _088528_);
  xor g_143880_(_085714_, _088528_, _088529_);
  xor g_143881_(_085713_, _088528_, _088530_);
  xor g_143882_(_086977_, _088529_, _088531_);
  not g_143883_(_088531_, _088532_);
  or g_143884_(_085730_, _088532_, _088534_);
  xor g_143885_(_085730_, _088531_, _088535_);
  or g_143886_(_085725_, _088535_, _088536_);
  xor g_143887_(_085726_, _088535_, _088537_);
  and g_143888_(_085734_, _088537_, _088538_);
  and g_143889_(_085737_, _088538_, _088539_);
  or g_143890_(_085734_, _088537_, _088540_);
  not g_143891_(_088540_, _088541_);
  or g_143892_(_085737_, _088537_, _088542_);
  and g_143893_(_088540_, _088542_, _088543_);
  not g_143894_(_088543_, _088545_);
  or g_143895_(_088539_, _088545_, _088546_);
  or g_143896_(_085742_, _088546_, _088547_);
  xor g_143897_(_085741_, _088546_, _088548_);
  or g_143898_(_085744_, _088548_, _088549_);
  xor g_143899_(_085745_, _088548_, _088550_);
  or g_143900_(_082897_, _085746_, _088551_);
  not g_143901_(_088551_, _088552_);
  or g_143902_(_088550_, _088551_, _088553_);
  xor g_143903_(_088550_, _088551_, _088554_);
  xor g_143904_(_088550_, _088552_, _088556_);
  or g_143905_(_086976_, _088556_, _088557_);
  not g_143906_(_088557_, _088558_);
  xor g_143907_(_086976_, _088554_, _088559_);
  or g_143908_(_086975_, _088559_, _088560_);
  not g_143909_(_088560_, _088561_);
  xor g_143910_(_086974_, _088559_, _088562_);
  and g_143911_(_086973_, _088562_, _088563_);
  or g_143912_(_086973_, _088562_, _088564_);
  not g_143913_(_088564_, _088565_);
  xor g_143914_(_086973_, _088562_, _088567_);
  or g_143915_(_088563_, _088565_, _088568_);
  or g_143916_(_086972_, _088568_, _088569_);
  xor g_143917_(_086972_, _088567_, _088570_);
  or g_143918_(_086969_, _088570_, _088571_);
  and g_143919_(_086969_, _088570_, _088572_);
  xor g_143920_(_086970_, _088570_, _088573_);
  or g_143921_(_085756_, _088573_, _088574_);
  xor g_143922_(_085757_, _088573_, _088575_);
  or g_143923_(_085759_, _088575_, _088576_);
  not g_143924_(_088576_, _088578_);
  xor g_143925_(_085759_, _088575_, _088579_);
  not g_143926_(_088579_, _088580_);
  xor g_143927_(_085764_, _088579_, _088581_);
  or g_143928_(_085768_, _088581_, _088582_);
  not g_143929_(_088582_, _088583_);
  xor g_143930_(_085767_, _088581_, _088584_);
  or g_143931_(_085777_, _088584_, _088585_);
  not g_143932_(_088585_, _088586_);
  xor g_143933_(_085776_, _088584_, _088587_);
  or g_143934_(_085775_, _088587_, _088589_);
  and g_143935_(_085775_, _088587_, _088590_);
  xor g_143936_(_085774_, _088587_, _088591_);
  and g_143937_(_085780_, _085789_, _088592_);
  xor g_143938_(_088591_, _088592_, _088593_);
  not g_143939_(_088593_, _088594_);
  or g_143940_(_085787_, _088594_, _088595_);
  xor g_143941_(_085787_, _088593_, _088596_);
  and g_143942_(_085792_, _085794_, _088597_);
  not g_143943_(_088597_, _088598_);
  xor g_143944_(_088596_, _088598_, _088600_);
  or g_143945_(_086967_, _088600_, _088601_);
  not g_143946_(_088601_, _088602_);
  and g_143947_(_086967_, _088600_, _088603_);
  xor g_143948_(_086967_, _088600_, _088604_);
  or g_143949_(_088602_, _088603_, _088605_);
  or g_143950_(_086966_, _088605_, _088606_);
  xor g_143951_(_086966_, _088604_, _088607_);
  not g_143952_(_088607_, _088608_);
  and g_143953_(_085803_, _088608_, _088609_);
  not g_143954_(_088609_, _088611_);
  or g_143955_(_085808_, _088607_, _088612_);
  not g_143956_(_088612_, _088613_);
  xor g_143957_(_085807_, _088607_, _088614_);
  and g_143958_(_085802_, _088614_, _088615_);
  or g_143959_(_088609_, _088615_, _088616_);
  or g_143960_(_085811_, _088616_, _088617_);
  not g_143961_(_088617_, _088618_);
  xor g_143962_(_085811_, _088616_, _088619_);
  and g_143963_(_085814_, _088619_, _088620_);
  xor g_143964_(_085813_, _088619_, _088622_);
  not g_143965_(_088622_, _088623_);
  and g_143966_(_085822_, _088623_, _088624_);
  or g_143967_(_085823_, _088622_, _088625_);
  xor g_143968_(_085822_, _088622_, _088626_);
  not g_143969_(_088626_, _088627_);
  or g_143970_(_085819_, _088626_, _088628_);
  not g_143971_(_088628_, _088629_);
  xor g_143972_(_085818_, _088626_, _088630_);
  or g_143973_(_085830_, _088630_, _088631_);
  or g_143974_(_085829_, _088627_, _088633_);
  and g_143975_(_088631_, _088633_, _088634_);
  not g_143976_(_088634_, _088635_);
  or g_143977_(_085833_, _088634_, _088636_);
  xor g_143978_(_085833_, _088634_, _088637_);
  xor g_143979_(_085833_, _088635_, _088638_);
  or g_143980_(_086965_, _088638_, _088639_);
  xor g_143981_(_086965_, _088637_, _088640_);
  or g_143982_(_086962_, _088640_, _088641_);
  xor g_143983_(_086963_, _088640_, _088642_);
  or g_143984_(_086959_, _088642_, _088644_);
  xor g_143985_(_086959_, _088642_, _088645_);
  not g_143986_(_088645_, _088646_);
  or g_143987_(_086958_, _088646_, _088647_);
  not g_143988_(_088647_, _088648_);
  xor g_143989_(_086958_, _088645_, _088649_);
  not g_143990_(_088649_, _088650_);
  or g_143991_(_085838_, _088649_, _088651_);
  and g_143992_(_085838_, _088649_, _088652_);
  xor g_143993_(_085838_, _088649_, _088653_);
  xor g_143994_(_085838_, _088650_, _088655_);
  and g_143995_(_085842_, _085848_, _088656_);
  xor g_143996_(_088653_, _088656_, _088657_);
  or g_143997_(_085844_, _088657_, _088658_);
  not g_143998_(_088658_, _088659_);
  xor g_143999_(_085844_, _088657_, _088660_);
  and g_144000_(_085854_, _088660_, _088661_);
  and g_144001_(_085862_, _088660_, _088662_);
  not g_144002_(_088662_, _088663_);
  xor g_144003_(_085860_, _088660_, _088664_);
  and g_144004_(_085853_, _088664_, _088666_);
  or g_144005_(_088661_, _088666_, _088667_);
  not g_144006_(_088667_, _088668_);
  or g_144007_(_085859_, _088667_, _088669_);
  xor g_144008_(_085859_, _088667_, _088670_);
  xor g_144009_(_085859_, _088668_, _088671_);
  or g_144010_(_086957_, _088671_, _088672_);
  xor g_144011_(_086957_, _088670_, _088673_);
  not g_144012_(_088673_, _088674_);
  and g_144013_(_086956_, _088674_, _088675_);
  not g_144014_(_088675_, _088677_);
  xor g_144015_(_086956_, _088673_, _088678_);
  not g_144016_(_088678_, _088679_);
  and g_144017_(_085878_, _088679_, _088680_);
  and g_144018_(_085879_, _088678_, _088681_);
  not g_144019_(_088681_, _088682_);
  xor g_144020_(_085878_, _088678_, _088683_);
  not g_144021_(_088683_, _088684_);
  and g_144022_(_085877_, _088684_, _088685_);
  xor g_144023_(_085877_, _088683_, _088686_);
  not g_144024_(_088686_, _088688_);
  xor g_144025_(_085882_, _088686_, _088689_);
  xor g_144026_(_085882_, _088688_, _088690_);
  xor g_144027_(_086955_, _088689_, _088691_);
  xor g_144028_(_086954_, _088691_, _088692_);
  or g_144029_(_086951_, _088692_, _088693_);
  not g_144030_(_088693_, _088694_);
  and g_144031_(_086951_, _088692_, _088695_);
  xor g_144032_(_086951_, _088692_, _088696_);
  xor g_144033_(_086952_, _088692_, _088697_);
  or g_144034_(_083051_, _085900_, _088699_);
  and g_144035_(_085898_, _088699_, _088700_);
  xor g_144036_(_088696_, _088700_, _088701_);
  xor g_144037_(_088697_, _088700_, _088702_);
  or g_144038_(_083054_, _085900_, _088703_);
  not g_144039_(_088703_, _088704_);
  and g_144040_(_088701_, _088703_, _088705_);
  and g_144041_(_085903_, _088705_, _088706_);
  and g_144042_(_085904_, _088702_, _088707_);
  and g_144043_(_088702_, _088704_, _088708_);
  or g_144044_(_088707_, _088708_, _088710_);
  or g_144045_(_088706_, _088710_, _088711_);
  or g_144046_(_085913_, _088711_, _088712_);
  not g_144047_(_088712_, _088713_);
  xor g_144048_(_085914_, _088711_, _088714_);
  or g_144049_(_085912_, _088714_, _088715_);
  not g_144050_(_088715_, _088716_);
  and g_144051_(_085912_, _088714_, _088717_);
  xor g_144052_(_085912_, _088714_, _088718_);
  or g_144053_(_088716_, _088717_, _088719_);
  or g_144054_(_085920_, _088719_, _088721_);
  xor g_144055_(_085920_, _088718_, _088722_);
  not g_144056_(_088722_, _088723_);
  or g_144057_(_085923_, _085924_, _088724_);
  and g_144058_(_085922_, _088724_, _088725_);
  xor g_144059_(_088722_, _088725_, _088726_);
  xor g_144060_(_088723_, _088725_, _088727_);
  or g_144061_(_086950_, _088727_, _088728_);
  xor g_144062_(_086950_, _088726_, _088729_);
  or g_144063_(_086948_, _088729_, _088730_);
  xor g_144064_(_086948_, _088729_, _088732_);
  and g_144065_(_086947_, _088732_, _088733_);
  xor g_144066_(_086947_, _088732_, _088734_);
  and g_144067_(_085931_, _088734_, _088735_);
  xor g_144068_(_085931_, _088734_, _088736_);
  not g_144069_(_088736_, _088737_);
  and g_144070_(_085933_, _085939_, _088738_);
  and g_144071_(_088737_, _088738_, _088739_);
  and g_144072_(_085934_, _088736_, _088740_);
  not g_144073_(_088740_, _088741_);
  and g_144074_(_085937_, _088736_, _088743_);
  or g_144075_(_088740_, _088743_, _088744_);
  or g_144076_(_088739_, _088744_, _088745_);
  and g_144077_(_085941_, _085945_, _088746_);
  not g_144078_(_088746_, _088747_);
  or g_144079_(_088745_, _088746_, _088748_);
  not g_144080_(_088748_, _088749_);
  xor g_144081_(_088745_, _088747_, _088750_);
  or g_144082_(_085947_, _088750_, _088751_);
  xor g_144083_(_085947_, _088750_, _088752_);
  or g_144084_(_083089_, _085952_, _088754_);
  not g_144085_(_088754_, _088755_);
  and g_144086_(_085950_, _088754_, _088756_);
  not g_144087_(_088756_, _088757_);
  xor g_144088_(_088752_, _088757_, _088758_);
  xor g_144089_(_088752_, _088756_, _088759_);
  or g_144090_(_086946_, _088759_, _088760_);
  xor g_144091_(_086946_, _088758_, _088761_);
  or g_144092_(_085966_, _088761_, _088762_);
  not g_144093_(_088762_, _088763_);
  xor g_144094_(_085966_, _088761_, _088765_);
  and g_144095_(_085958_, _088765_, _088766_);
  not g_144096_(_088766_, _088767_);
  xor g_144097_(_085958_, _088765_, _088768_);
  xor g_144098_(_085957_, _088765_, _088769_);
  or g_144099_(_085973_, _088769_, _088770_);
  xor g_144100_(_085973_, _088768_, _088771_);
  not g_144101_(_088771_, _088772_);
  or g_144102_(_086945_, _088771_, _088773_);
  xor g_144103_(_086945_, _088771_, _088774_);
  xor g_144104_(_086945_, _088772_, _088776_);
  or g_144105_(_086944_, _088776_, _088777_);
  not g_144106_(_088777_, _088778_);
  xor g_144107_(_086944_, _088774_, _088779_);
  or g_144108_(_085979_, _088779_, _088780_);
  not g_144109_(_088780_, _088781_);
  xor g_144110_(_085978_, _088779_, _088782_);
  or g_144111_(_085981_, _088782_, _088783_);
  xor g_144112_(_085983_, _088782_, _088784_);
  not g_144113_(_088784_, _088785_);
  and g_144114_(_085990_, _088785_, _088787_);
  and g_144115_(_085986_, _088784_, _088788_);
  and g_144116_(_085989_, _088788_, _088789_);
  and g_144117_(_085987_, _088785_, _088790_);
  not g_144118_(_088790_, _088791_);
  or g_144119_(_088789_, _088790_, _088792_);
  or g_144120_(_088787_, _088792_, _088793_);
  not g_144121_(_088793_, _088794_);
  and g_144122_(_085999_, _088794_, _088795_);
  or g_144123_(_085998_, _088793_, _088796_);
  and g_144124_(_085994_, _088793_, _088798_);
  and g_144125_(_085998_, _088798_, _088799_);
  and g_144126_(_085995_, _088794_, _088800_);
  or g_144127_(_088799_, _088800_, _088801_);
  or g_144128_(_088795_, _088801_, _088802_);
  or g_144129_(_086941_, _088802_, _088803_);
  xor g_144130_(_086942_, _088802_, _088804_);
  or g_144131_(_086939_, _088804_, _088805_);
  xor g_144132_(_086940_, _088804_, _088806_);
  or g_144133_(_086936_, _088806_, _088807_);
  xor g_144134_(_086937_, _088806_, _088809_);
  or g_144135_(_086009_, _088809_, _088810_);
  xor g_144136_(_086010_, _088809_, _088811_);
  or g_144137_(_086007_, _088811_, _088812_);
  xor g_144138_(_086008_, _088811_, _088813_);
  or g_144139_(_086934_, _088813_, _088814_);
  not g_144140_(_088814_, _088815_);
  xor g_144141_(_086935_, _088813_, _088816_);
  or g_144142_(_086932_, _088816_, _088817_);
  not g_144143_(_088817_, _088818_);
  and g_144144_(_086932_, _088816_, _088820_);
  xor g_144145_(_086933_, _088816_, _088821_);
  and g_144146_(_086020_, _086023_, _088822_);
  not g_144147_(_088822_, _088823_);
  xor g_144148_(_088821_, _088823_, _088824_);
  not g_144149_(_088824_, _088825_);
  or g_144150_(_086931_, _088824_, _088826_);
  xor g_144151_(_086931_, _088824_, _088827_);
  xor g_144152_(_086931_, _088825_, _088828_);
  or g_144153_(_086930_, _088828_, _088829_);
  xor g_144154_(_086930_, _088827_, _088831_);
  or g_144155_(_086030_, _088831_, _088832_);
  xor g_144156_(_086030_, _088831_, _088833_);
  and g_144157_(_086929_, _088833_, _088834_);
  xor g_144158_(_086929_, _088833_, _088835_);
  and g_144159_(_086928_, _088835_, _088836_);
  or g_144160_(_086928_, _088835_, _088837_);
  xor g_144161_(_086928_, _088835_, _088838_);
  not g_144162_(_088838_, _088839_);
  and g_144163_(_086035_, _088838_, _088840_);
  xor g_144164_(_086035_, _088838_, _088842_);
  xor g_144165_(_086035_, _088839_, _088843_);
  or g_144166_(_086041_, _086042_, _088844_);
  and g_144167_(_086039_, _088844_, _088845_);
  xor g_144168_(_088842_, _088845_, _088846_);
  or g_144169_(_086926_, _088846_, _088847_);
  xor g_144170_(_086926_, _088846_, _088848_);
  not g_144171_(_088848_, _088849_);
  and g_144172_(_086046_, _086051_, _088850_);
  xor g_144173_(_088848_, _088850_, _088851_);
  xor g_144174_(_086925_, _088851_, _088853_);
  not g_144175_(_088853_, _088854_);
  and g_144176_(_086060_, _088853_, _088855_);
  not g_144177_(_088855_, _088856_);
  or g_144178_(_086063_, _088854_, _088857_);
  not g_144179_(_088857_, _088858_);
  xor g_144180_(_086063_, _088853_, _088859_);
  and g_144181_(_086058_, _088859_, _088860_);
  or g_144182_(_088855_, _088860_, _088861_);
  or g_144183_(_086924_, _088861_, _088862_);
  xor g_144184_(_086923_, _088861_, _088864_);
  or g_144185_(_086921_, _088864_, _088865_);
  xor g_144186_(_086922_, _088864_, _088866_);
  or g_144187_(_086919_, _088866_, _088867_);
  xor g_144188_(_086920_, _088866_, _088868_);
  or g_144189_(_078222_, _080171_, _088869_);
  or g_144190_(_083195_, _088869_, _088870_);
  or g_144191_(_086067_, _088870_, _088871_);
  or g_144192_(_088868_, _088871_, _088872_);
  xor g_144193_(_088868_, _088871_, _088873_);
  not g_144194_(_088873_, _088875_);
  and g_144195_(_086918_, _088873_, _088876_);
  or g_144196_(_086917_, _088875_, _088877_);
  xor g_144197_(_086917_, _088873_, _088878_);
  or g_144198_(_086914_, _088878_, _088879_);
  xor g_144199_(_086914_, _088878_, _088880_);
  xor g_144200_(_086915_, _088878_, _088881_);
  xor g_144201_(_086083_, _088880_, _088882_);
  xor g_144202_(_086084_, _088880_, _088883_);
  or g_144203_(_086093_, _088882_, _088884_);
  not g_144204_(_088884_, _088886_);
  and g_144205_(_086095_, _088882_, _088887_);
  or g_144206_(_086094_, _088883_, _088888_);
  and g_144207_(_086093_, _088887_, _088889_);
  or g_144208_(_086091_, _088888_, _088890_);
  and g_144209_(_086094_, _088883_, _088891_);
  not g_144210_(_088891_, _088892_);
  and g_144211_(_088890_, _088892_, _088893_);
  or g_144212_(_088889_, _088891_, _088894_);
  and g_144213_(_088884_, _088893_, _088895_);
  or g_144214_(_088886_, _088894_, _088897_);
  and g_144215_(_086098_, _088895_, _088898_);
  or g_144216_(_086097_, _088897_, _088899_);
  xor g_144217_(_086097_, _088895_, _088900_);
  or g_144218_(_086105_, _088900_, _088901_);
  not g_144219_(_088901_, _088902_);
  xor g_144220_(_086104_, _088900_, _088903_);
  or g_144221_(_086107_, _088903_, _088904_);
  xor g_144222_(_086106_, _088903_, _088905_);
  or g_144223_(_086111_, _088905_, _088906_);
  not g_144224_(_088906_, _088908_);
  and g_144225_(_086111_, _088905_, _088909_);
  or g_144226_(_088908_, _088909_, _088910_);
  not g_144227_(_088910_, _088911_);
  and g_144228_(_086115_, _086118_, _088912_);
  xor g_144229_(_088911_, _088912_, _088913_);
  or g_144230_(_086913_, _088913_, _088914_);
  not g_144231_(_088914_, _088915_);
  xor g_144232_(_086913_, _088913_, _088916_);
  and g_144233_(_086911_, _088916_, _088917_);
  not g_144234_(_088917_, _088919_);
  xor g_144235_(_086911_, _088916_, _088920_);
  xor g_144236_(_086912_, _088916_, _088921_);
  or g_144237_(_086124_, _088921_, _088922_);
  xor g_144238_(_086124_, _088920_, _088923_);
  not g_144239_(_088923_, _088924_);
  or g_144240_(_086128_, _088923_, _088925_);
  xor g_144241_(_086128_, _088924_, _088926_);
  or g_144242_(_086132_, _088926_, _088927_);
  not g_144243_(_088927_, _088928_);
  and g_144244_(_086132_, _088926_, _088930_);
  or g_144245_(_088928_, _088930_, _088931_);
  or g_144246_(_086133_, _088931_, _088932_);
  not g_144247_(_088932_, _088933_);
  xor g_144248_(_086133_, _088931_, _088934_);
  and g_144249_(_086910_, _088934_, _088935_);
  not g_144250_(_088935_, _088936_);
  xor g_144251_(_086909_, _088934_, _088937_);
  or g_144252_(_086908_, _088937_, _088938_);
  not g_144253_(_088938_, _088939_);
  xor g_144254_(_086908_, _088937_, _088941_);
  not g_144255_(_088941_, _088942_);
  or g_144256_(_086907_, _088942_, _088943_);
  not g_144257_(_088943_, _088944_);
  xor g_144258_(_086907_, _088941_, _088945_);
  not g_144259_(_088945_, _088946_);
  or g_144260_(_086906_, _088945_, _088947_);
  xor g_144261_(_086906_, _088946_, _088948_);
  or g_144262_(_086142_, _088948_, _088949_);
  not g_144263_(_088949_, _088950_);
  xor g_144264_(_086142_, _088948_, _088952_);
  and g_144265_(_086904_, _088952_, _088953_);
  not g_144266_(_088953_, _088954_);
  xor g_144267_(_086904_, _088952_, _088955_);
  or g_144268_(_083272_, _086144_, _088956_);
  not g_144269_(_088956_, _088957_);
  or g_144270_(_080250_, _086902_, _088958_);
  not g_144271_(_088958_, _088959_);
  and g_144272_(_088956_, _088958_, _088960_);
  xor g_144273_(_088955_, _088960_, _088961_);
  not g_144274_(_088961_, _088963_);
  and g_144275_(_086901_, _088963_, _088964_);
  not g_144276_(_088964_, _088965_);
  xor g_144277_(_086900_, _088961_, _088966_);
  and g_144278_(_086152_, _088966_, _088967_);
  not g_144279_(_088967_, _088968_);
  xor g_144280_(_086152_, _088966_, _088969_);
  not g_144281_(_088969_, _088970_);
  or g_144282_(_083286_, _086161_, _088971_);
  not g_144283_(_088971_, _088972_);
  and g_144284_(_086159_, _088971_, _088974_);
  xor g_144285_(_088970_, _088974_, _088975_);
  xor g_144286_(_088969_, _088974_, _088976_);
  or g_144287_(_086898_, _088976_, _088977_);
  not g_144288_(_088977_, _088978_);
  xor g_144289_(_086898_, _088975_, _088979_);
  or g_144290_(_086166_, _088979_, _088980_);
  not g_144291_(_088980_, _088981_);
  xor g_144292_(_086166_, _088979_, _088982_);
  not g_144293_(_088982_, _088983_);
  or g_144294_(_086897_, _088983_, _088985_);
  not g_144295_(_088985_, _088986_);
  xor g_144296_(_086897_, _088982_, _088987_);
  or g_144297_(_086896_, _088987_, _088988_);
  not g_144298_(_088988_, _088989_);
  and g_144299_(_086896_, _088987_, _088990_);
  xor g_144300_(_086896_, _088987_, _088991_);
  or g_144301_(_088989_, _088990_, _088992_);
  or g_144302_(_086895_, _088992_, _088993_);
  or g_144303_(_083301_, _086172_, _088994_);
  or g_144304_(_088992_, _088994_, _088996_);
  not g_144305_(_088996_, _088997_);
  xor g_144306_(_088991_, _088994_, _088998_);
  and g_144307_(_086895_, _088998_, _088999_);
  not g_144308_(_088999_, _089000_);
  and g_144309_(_088993_, _089000_, _089001_);
  and g_144310_(_086176_, _089001_, _089002_);
  xor g_144311_(_086175_, _089001_, _089003_);
  not g_144312_(_089003_, _089004_);
  and g_144313_(_086179_, _086187_, _089005_);
  xor g_144314_(_089004_, _089005_, _089007_);
  or g_144315_(_086186_, _089007_, _089008_);
  not g_144316_(_089008_, _089009_);
  and g_144317_(_086186_, _089007_, _089010_);
  xor g_144318_(_086186_, _089007_, _089011_);
  or g_144319_(_089009_, _089010_, _089012_);
  or g_144320_(_086192_, _089012_, _089013_);
  xor g_144321_(_086192_, _089011_, _089014_);
  not g_144322_(_089014_, _089015_);
  or g_144323_(_086195_, _089014_, _089016_);
  xor g_144324_(_086195_, _089015_, _089018_);
  or g_144325_(_083320_, _086198_, _089019_);
  and g_144326_(_086197_, _089019_, _089020_);
  xor g_144327_(_089018_, _089020_, _089021_);
  not g_144328_(_089021_, _089022_);
  xor g_144329_(_086893_, _089021_, _089023_);
  and g_144330_(_086207_, _089023_, _089024_);
  or g_144331_(_086207_, _089023_, _089025_);
  xor g_144332_(_086207_, _089023_, _089026_);
  xor g_144333_(_086208_, _089023_, _089027_);
  or g_144334_(_083334_, _086209_, _089029_);
  or g_144335_(_086209_, _086210_, _089030_);
  and g_144336_(_089029_, _089030_, _089031_);
  xor g_144337_(_089026_, _089031_, _089032_);
  xor g_144338_(_089027_, _089031_, _089033_);
  or g_144339_(_086215_, _089032_, _089034_);
  not g_144340_(_089034_, _089035_);
  xor g_144341_(_086215_, _089033_, _089036_);
  or g_144342_(_086891_, _089036_, _089037_);
  or g_144343_(_083338_, _083339_, _089038_);
  or g_144344_(_086216_, _089038_, _089040_);
  not g_144345_(_089040_, _089041_);
  and g_144346_(_086891_, _089036_, _089042_);
  not g_144347_(_089042_, _089043_);
  or g_144348_(_089040_, _089042_, _089044_);
  not g_144349_(_089044_, _089045_);
  and g_144350_(_089037_, _089045_, _089046_);
  not g_144351_(_089046_, _089047_);
  and g_144352_(_089037_, _089043_, _089048_);
  or g_144353_(_089041_, _089048_, _089049_);
  and g_144354_(_089047_, _089049_, _089051_);
  xor g_144355_(_086219_, _089051_, _089052_);
  xor g_144356_(_086218_, _089051_, _089053_);
  and g_144357_(_086222_, _089053_, _089054_);
  or g_144358_(_086221_, _089052_, _089055_);
  and g_144359_(_086227_, _089054_, _089056_);
  or g_144360_(_086226_, _089055_, _089057_);
  and g_144361_(_086221_, _089051_, _089058_);
  not g_144362_(_089058_, _089059_);
  and g_144363_(_086226_, _089052_, _089060_);
  or g_144364_(_086227_, _089053_, _089062_);
  and g_144365_(_089059_, _089062_, _089063_);
  or g_144366_(_089058_, _089060_, _089064_);
  and g_144367_(_089057_, _089063_, _089065_);
  or g_144368_(_089056_, _089064_, _089066_);
  and g_144369_(_086229_, _086234_, _089067_);
  xor g_144370_(_089065_, _089067_, _089068_);
  and g_144371_(_086241_, _089068_, _089069_);
  or g_144372_(_086241_, _089068_, _089070_);
  not g_144373_(_089070_, _089071_);
  xor g_144374_(_086241_, _089068_, _089073_);
  or g_144375_(_089069_, _089071_, _089074_);
  and g_144376_(_086239_, _086244_, _089075_);
  xor g_144377_(_089073_, _089075_, _089076_);
  or g_144378_(_086252_, _089076_, _089077_);
  xor g_144379_(_086252_, _089076_, _089078_);
  not g_144380_(_089078_, _089079_);
  or g_144381_(_086255_, _089079_, _089080_);
  xor g_144382_(_086255_, _089078_, _089081_);
  not g_144383_(_089081_, _089082_);
  or g_144384_(_086889_, _089081_, _089084_);
  xor g_144385_(_086889_, _089082_, _089085_);
  not g_144386_(_089085_, _089086_);
  or g_144387_(_086888_, _089085_, _089087_);
  not g_144388_(_089087_, _089088_);
  xor g_144389_(_086888_, _089086_, _089089_);
  or g_144390_(_086887_, _089089_, _089090_);
  xor g_144391_(_086886_, _089089_, _089091_);
  or g_144392_(_086884_, _089091_, _089092_);
  xor g_144393_(_086885_, _089091_, _089093_);
  not g_144394_(_089093_, _089095_);
  and g_144395_(_086262_, _086265_, _089096_);
  xor g_144396_(_089093_, _089096_, _089097_);
  xor g_144397_(_089095_, _089096_, _089098_);
  xor g_144398_(_086882_, _089097_, _089099_);
  or g_144399_(_086880_, _089099_, _089100_);
  not g_144400_(_089100_, _089101_);
  xor g_144401_(_086880_, _089099_, _089102_);
  not g_144402_(_089102_, _089103_);
  or g_144403_(_086281_, _089103_, _089104_);
  xor g_144404_(_086281_, _089102_, _089106_);
  not g_144405_(_089106_, _089107_);
  and g_144406_(_086277_, _089107_, _089108_);
  xor g_144407_(_086278_, _089106_, _089109_);
  not g_144408_(_089109_, _089110_);
  and g_144409_(_086283_, _089109_, _089111_);
  xor g_144410_(_086283_, _089109_, _089112_);
  xor g_144411_(_086283_, _089110_, _089113_);
  or g_144412_(_086879_, _089113_, _089114_);
  not g_144413_(_089114_, _089115_);
  xor g_144414_(_086879_, _089112_, _089117_);
  not g_144415_(_089117_, _089118_);
  or g_144416_(_086878_, _089117_, _089119_);
  xor g_144417_(_086878_, _089118_, _089120_);
  not g_144418_(_089120_, _089121_);
  or g_144419_(_086877_, _089120_, _089122_);
  xor g_144420_(_086877_, _089121_, _089123_);
  not g_144421_(_089123_, _089124_);
  or g_144422_(_086876_, _089123_, _089125_);
  not g_144423_(_089125_, _089126_);
  xor g_144424_(_086876_, _089124_, _089128_);
  or g_144425_(_086298_, _089128_, _089129_);
  not g_144426_(_089129_, _089130_);
  xor g_144427_(_086297_, _089128_, _089131_);
  not g_144428_(_089131_, _089132_);
  or g_144429_(_086300_, _086303_, _089133_);
  or g_144430_(_083439_, _086300_, _089134_);
  and g_144431_(_086293_, _089134_, _089135_);
  and g_144432_(_089133_, _089135_, _089136_);
  xor g_144433_(_089131_, _089136_, _089137_);
  xor g_144434_(_089132_, _089136_, _089139_);
  or g_144435_(_086875_, _089139_, _089140_);
  xor g_144436_(_086875_, _089137_, _089141_);
  not g_144437_(_089141_, _089142_);
  or g_144438_(_086874_, _089141_, _089143_);
  xor g_144439_(_086874_, _089142_, _089144_);
  or g_144440_(_086308_, _089144_, _089145_);
  xor g_144441_(_086308_, _089144_, _089146_);
  xor g_144442_(_086307_, _089144_, _089147_);
  or g_144443_(_083451_, _086314_, _089148_);
  and g_144444_(_086313_, _089148_, _089150_);
  xor g_144445_(_089146_, _089150_, _089151_);
  or g_144446_(_086873_, _089151_, _089152_);
  xor g_144447_(_086873_, _089151_, _089153_);
  not g_144448_(_089153_, _089154_);
  and g_144449_(_086871_, _089153_, _089155_);
  or g_144450_(_086870_, _089154_, _089156_);
  xor g_144451_(_086870_, _089153_, _089157_);
  not g_144452_(_089157_, _089158_);
  or g_144453_(_083460_, _086317_, _089159_);
  or g_144454_(_083462_, _086320_, _089161_);
  and g_144455_(_089159_, _089161_, _089162_);
  xor g_144456_(_089158_, _089162_, _089163_);
  or g_144457_(_086869_, _089163_, _089164_);
  xor g_144458_(_086869_, _089163_, _089165_);
  or g_144459_(_086328_, _089165_, _089166_);
  or g_144460_(_077692_, _080466_, _089167_);
  or g_144461_(_083468_, _089167_, _089168_);
  or g_144462_(_086322_, _089168_, _089169_);
  or g_144463_(_089163_, _089169_, _089170_);
  and g_144464_(_089166_, _089170_, _089172_);
  not g_144465_(_089172_, _089173_);
  or g_144466_(_086327_, _089173_, _089174_);
  not g_144467_(_089174_, _089175_);
  xor g_144468_(_086327_, _089172_, _089176_);
  or g_144469_(_086332_, _089176_, _089177_);
  xor g_144470_(_086332_, _089176_, _089178_);
  not g_144471_(_089178_, _089179_);
  or g_144472_(_083480_, _086333_, _089180_);
  not g_144473_(_089180_, _089181_);
  and g_144474_(_086335_, _089180_, _089183_);
  xor g_144475_(_089178_, _089183_, _089184_);
  or g_144476_(_083976_, _086342_, _089185_);
  or g_144477_(_086337_, _086339_, _089186_);
  and g_144478_(_089185_, _089186_, _089187_);
  xor g_144479_(_089184_, _089187_, _089188_);
  and g_144480_(_086868_, _089188_, _089189_);
  not g_144481_(_089189_, _089190_);
  xor g_144482_(_086867_, _089188_, _089191_);
  not g_144483_(_089191_, _089192_);
  and g_144484_(_086346_, _089192_, _089194_);
  not g_144485_(_089194_, _089195_);
  and g_144486_(_086344_, _089191_, _089196_);
  or g_144487_(_089194_, _089196_, _089197_);
  not g_144488_(_089197_, _089198_);
  or g_144489_(_086350_, _089197_, _089199_);
  xor g_144490_(_086350_, _089198_, _089200_);
  not g_144491_(_089200_, _089201_);
  and g_144492_(_086353_, _086357_, _089202_);
  xor g_144493_(_089201_, _089202_, _089203_);
  or g_144494_(_086361_, _089203_, _089205_);
  not g_144495_(_089205_, _089206_);
  xor g_144496_(_086361_, _089203_, _089207_);
  not g_144497_(_089207_, _089208_);
  or g_144498_(_083504_, _086366_, _089209_);
  and g_144499_(_086359_, _089209_, _089210_);
  xor g_144500_(_089207_, _089210_, _089211_);
  or g_144501_(_086866_, _089211_, _089212_);
  xor g_144502_(_086866_, _089211_, _089213_);
  not g_144503_(_089213_, _089214_);
  or g_144504_(_086372_, _089214_, _089216_);
  xor g_144505_(_086372_, _089213_, _089217_);
  not g_144506_(_089217_, _089218_);
  or g_144507_(_086375_, _089217_, _089219_);
  xor g_144508_(_086375_, _089218_, _089220_);
  not g_144509_(_089220_, _089221_);
  and g_144510_(_086865_, _089221_, _089222_);
  xor g_144511_(_086864_, _089220_, _089223_);
  not g_144512_(_089223_, _089224_);
  or g_144513_(_083514_, _086863_, _089225_);
  not g_144514_(_089225_, _089227_);
  and g_144515_(_086379_, _089225_, _089228_);
  xor g_144516_(_089224_, _089228_, _089229_);
  xor g_144517_(_089223_, _089228_, _089230_);
  and g_144518_(_086384_, _086387_, _089231_);
  xor g_144519_(_089229_, _089231_, _089232_);
  or g_144520_(_086862_, _089232_, _089233_);
  xor g_144521_(_086862_, _089232_, _089234_);
  and g_144522_(_086860_, _089234_, _089235_);
  not g_144523_(_089235_, _089236_);
  xor g_144524_(_086859_, _089234_, _089238_);
  and g_144525_(_086394_, _089238_, _089239_);
  or g_144526_(_086394_, _089238_, _089240_);
  not g_144527_(_089240_, _089241_);
  or g_144528_(_089239_, _089241_, _089242_);
  or g_144529_(_083540_, _086398_, _089243_);
  and g_144530_(_086397_, _089243_, _089244_);
  xor g_144531_(_089242_, _089244_, _089245_);
  not g_144532_(_089245_, _089246_);
  and g_144533_(_086857_, _089245_, _089247_);
  or g_144534_(_086856_, _089246_, _089249_);
  xor g_144535_(_086856_, _089245_, _089250_);
  and g_144536_(_086404_, _086407_, _089251_);
  xor g_144537_(_089250_, _089251_, _089252_);
  and g_144538_(_086415_, _089252_, _089253_);
  xor g_144539_(_086415_, _089252_, _089254_);
  and g_144540_(_086413_, _089254_, _089255_);
  xor g_144541_(_086413_, _089254_, _089256_);
  xor g_144542_(_086412_, _089254_, _089257_);
  and g_144543_(_086419_, _086423_, _089258_);
  xor g_144544_(_089257_, _089258_, _089260_);
  xor g_144545_(_089256_, _089258_, _089261_);
  or g_144546_(_086855_, _089261_, _089262_);
  xor g_144547_(_086855_, _089260_, _089263_);
  not g_144548_(_089263_, _089264_);
  or g_144549_(_086854_, _089263_, _089265_);
  xor g_144550_(_086854_, _089264_, _089266_);
  not g_144551_(_089266_, _089267_);
  or g_144552_(_086853_, _089266_, _089268_);
  xor g_144553_(_086853_, _089267_, _089269_);
  or g_144554_(_083577_, _086427_, _089271_);
  and g_144555_(_086431_, _089271_, _089272_);
  or g_144556_(_089269_, _089272_, _089273_);
  xor g_144557_(_089269_, _089272_, _089274_);
  and g_144558_(_086434_, _089274_, _089275_);
  not g_144559_(_089275_, _089276_);
  xor g_144560_(_086434_, _089274_, _089277_);
  xor g_144561_(_086435_, _089274_, _089278_);
  or g_144562_(_086437_, _089278_, _089279_);
  xor g_144563_(_086437_, _089277_, _089280_);
  not g_144564_(_089280_, _089282_);
  or g_144565_(_086852_, _089280_, _089283_);
  xor g_144566_(_086852_, _089280_, _089284_);
  xor g_144567_(_086852_, _089282_, _089285_);
  or g_144568_(_086851_, _089285_, _089286_);
  not g_144569_(_089286_, _089287_);
  xor g_144570_(_086851_, _089284_, _089288_);
  not g_144571_(_089288_, _089289_);
  or g_144572_(_086849_, _089288_, _089290_);
  not g_144573_(_089290_, _089291_);
  xor g_144574_(_086849_, _089289_, _089293_);
  or g_144575_(_086847_, _089293_, _089294_);
  not g_144576_(_089294_, _089295_);
  xor g_144577_(_086848_, _089293_, _089296_);
  or g_144578_(_086446_, _089296_, _089297_);
  xor g_144579_(_086445_, _089296_, _089298_);
  not g_144580_(_089298_, _089299_);
  or g_144581_(_086846_, _089298_, _089300_);
  xor g_144582_(_086846_, _089298_, _089301_);
  xor g_144583_(_086846_, _089299_, _089302_);
  or g_144584_(_086845_, _089302_, _089304_);
  not g_144585_(_089304_, _089305_);
  xor g_144586_(_086845_, _089301_, _089306_);
  and g_144587_(_086452_, _086458_, _089307_);
  and g_144588_(_089306_, _089307_, _089308_);
  or g_144589_(_086458_, _089306_, _089309_);
  or g_144590_(_086452_, _089306_, _089310_);
  and g_144591_(_089309_, _089310_, _089311_);
  not g_144592_(_089311_, _089312_);
  or g_144593_(_089308_, _089312_, _089313_);
  or g_144594_(_086459_, _089313_, _089315_);
  not g_144595_(_089315_, _089316_);
  xor g_144596_(_086460_, _089313_, _089317_);
  not g_144597_(_089317_, _089318_);
  or g_144598_(_083615_, _086467_, _089319_);
  and g_144599_(_086465_, _089319_, _089320_);
  xor g_144600_(_089317_, _089320_, _089321_);
  xor g_144601_(_089318_, _089320_, _089322_);
  or g_144602_(_086844_, _089322_, _089323_);
  not g_144603_(_089323_, _089324_);
  xor g_144604_(_086844_, _089321_, _089326_);
  not g_144605_(_089326_, _089327_);
  or g_144606_(_086473_, _089326_, _089328_);
  xor g_144607_(_086473_, _089327_, _089329_);
  not g_144608_(_089329_, _089330_);
  or g_144609_(_086843_, _089329_, _089331_);
  xor g_144610_(_086843_, _089330_, _089332_);
  or g_144611_(_086841_, _089332_, _089333_);
  xor g_144612_(_086841_, _089332_, _089334_);
  xor g_144613_(_086842_, _089332_, _089335_);
  and g_144614_(_086479_, _089334_, _089337_);
  or g_144615_(_086480_, _089335_, _089338_);
  xor g_144616_(_086480_, _089334_, _089339_);
  or g_144617_(_086840_, _089339_, _089340_);
  not g_144618_(_089340_, _089341_);
  and g_144619_(_086840_, _089339_, _089342_);
  xor g_144620_(_086840_, _089339_, _089343_);
  or g_144621_(_089341_, _089342_, _089344_);
  and g_144622_(_086838_, _089343_, _089345_);
  or g_144623_(_086837_, _089344_, _089346_);
  xor g_144624_(_086838_, _089343_, _089348_);
  xor g_144625_(_086837_, _089343_, _089349_);
  or g_144626_(_086486_, _089349_, _089350_);
  not g_144627_(_089350_, _089351_);
  xor g_144628_(_086486_, _089348_, _089352_);
  or g_144629_(_086490_, _089352_, _089353_);
  not g_144630_(_089353_, _089354_);
  xor g_144631_(_086490_, _089352_, _089355_);
  not g_144632_(_089355_, _089356_);
  and g_144633_(_086495_, _089355_, _089357_);
  or g_144634_(_086494_, _089356_, _089359_);
  xor g_144635_(_086495_, _089355_, _089360_);
  xor g_144636_(_086494_, _089355_, _089361_);
  or g_144637_(_083646_, _086498_, _089362_);
  not g_144638_(_089362_, _089363_);
  and g_144639_(_086492_, _089362_, _089364_);
  xor g_144640_(_089360_, _089364_, _089365_);
  or g_144641_(_086835_, _089365_, _089366_);
  not g_144642_(_089366_, _089367_);
  xor g_144643_(_086835_, _089365_, _089368_);
  xor g_144644_(_086836_, _089365_, _089370_);
  and g_144645_(_086503_, _086506_, _089371_);
  xor g_144646_(_089370_, _089371_, _089372_);
  and g_144647_(_086509_, _089372_, _089373_);
  xor g_144648_(_086509_, _089372_, _089374_);
  xor g_144649_(_086508_, _089372_, _089375_);
  and g_144650_(_086834_, _089374_, _089376_);
  xor g_144651_(_086833_, _089375_, _089377_);
  not g_144652_(_089377_, _089378_);
  or g_144653_(_086831_, _089378_, _089379_);
  xor g_144654_(_086831_, _089377_, _089381_);
  not g_144655_(_089381_, _089382_);
  or g_144656_(_086515_, _089381_, _089383_);
  not g_144657_(_089383_, _089384_);
  xor g_144658_(_086515_, _089382_, _089385_);
  not g_144659_(_089385_, _089386_);
  or g_144660_(_086517_, _089385_, _089387_);
  and g_144661_(_086517_, _089385_, _089388_);
  xor g_144662_(_086517_, _089386_, _089389_);
  and g_144663_(_083679_, _086520_, _089390_);
  or g_144664_(_083678_, _086522_, _089392_);
  or g_144665_(_086523_, _089390_, _089393_);
  xor g_144666_(_089389_, _089393_, _089394_);
  or g_144667_(_086829_, _089394_, _089395_);
  xor g_144668_(_086829_, _089394_, _089396_);
  and g_144669_(_086826_, _089396_, _089397_);
  xor g_144670_(_086827_, _089396_, _089398_);
  not g_144671_(_089398_, _089399_);
  and g_144672_(_086825_, _089399_, _089400_);
  not g_144673_(_089400_, _089401_);
  xor g_144674_(_086825_, _089398_, _089403_);
  or g_144675_(_086824_, _089403_, _089404_);
  not g_144676_(_089404_, _089405_);
  and g_144677_(_086824_, _089403_, _089406_);
  or g_144678_(_089405_, _089406_, _089407_);
  not g_144679_(_089407_, _089408_);
  or g_144680_(_086823_, _089407_, _089409_);
  xor g_144681_(_086823_, _089408_, _089410_);
  or g_144682_(_086822_, _089410_, _089411_);
  xor g_144683_(_086821_, _089410_, _089412_);
  or g_144684_(_086820_, _089412_, _089414_);
  not g_144685_(_089414_, _089415_);
  xor g_144686_(_086820_, _089412_, _089416_);
  not g_144687_(_089416_, _089417_);
  or g_144688_(_086539_, _089417_, _089418_);
  not g_144689_(_089418_, _089419_);
  xor g_144690_(_086539_, _089416_, _089420_);
  or g_144691_(_086535_, _089420_, _089421_);
  xor g_144692_(_086536_, _089420_, _089422_);
  not g_144693_(_089422_, _089423_);
  and g_144694_(_086545_, _086547_, _089425_);
  xor g_144695_(_089423_, _089425_, _089426_);
  and g_144696_(_086551_, _089426_, _089427_);
  and g_144697_(_086553_, _089427_, _089428_);
  not g_144698_(_089428_, _089429_);
  or g_144699_(_086553_, _089426_, _089430_);
  or g_144700_(_086551_, _089426_, _089431_);
  not g_144701_(_089431_, _089432_);
  and g_144702_(_089430_, _089431_, _089433_);
  not g_144703_(_089433_, _089434_);
  and g_144704_(_089429_, _089433_, _089436_);
  or g_144705_(_089428_, _089434_, _089437_);
  or g_144706_(_086819_, _089437_, _089438_);
  xor g_144707_(_086819_, _089436_, _089439_);
  or g_144708_(_086818_, _089439_, _089440_);
  xor g_144709_(_086816_, _089439_, _089441_);
  not g_144710_(_089441_, _089442_);
  or g_144711_(_086562_, _089441_, _089443_);
  xor g_144712_(_086562_, _089441_, _089444_);
  xor g_144713_(_086562_, _089442_, _089445_);
  or g_144714_(_086815_, _089445_, _089447_);
  xor g_144715_(_086815_, _089444_, _089448_);
  or g_144716_(_086813_, _089448_, _089449_);
  xor g_144717_(_086814_, _089448_, _089450_);
  and g_144718_(_086570_, _086572_, _089451_);
  xor g_144719_(_089450_, _089451_, _089452_);
  not g_144720_(_089452_, _089453_);
  or g_144721_(_086574_, _089453_, _089454_);
  not g_144722_(_089454_, _089455_);
  xor g_144723_(_086574_, _089452_, _089456_);
  not g_144724_(_089456_, _089458_);
  or g_144725_(_083751_, _086575_, _089459_);
  not g_144726_(_089459_, _089460_);
  and g_144727_(_089458_, _089460_, _089461_);
  xor g_144728_(_089456_, _089459_, _089462_);
  xor g_144729_(_089456_, _089460_, _089463_);
  and g_144730_(_086812_, _089462_, _089464_);
  or g_144731_(_086811_, _089463_, _089465_);
  xor g_144732_(_086812_, _089462_, _089466_);
  xor g_144733_(_086811_, _089462_, _089467_);
  and g_144734_(_086580_, _089467_, _089469_);
  or g_144735_(_086581_, _089466_, _089470_);
  and g_144736_(_086809_, _089469_, _089471_);
  or g_144737_(_086810_, _089470_, _089472_);
  or g_144738_(_086809_, _089467_, _089473_);
  not g_144739_(_089473_, _089474_);
  or g_144740_(_086580_, _089467_, _089475_);
  and g_144741_(_089473_, _089475_, _089476_);
  not g_144742_(_089476_, _089477_);
  and g_144743_(_089472_, _089476_, _089478_);
  or g_144744_(_089471_, _089477_, _089480_);
  or g_144745_(_086808_, _089480_, _089481_);
  xor g_144746_(_086808_, _089478_, _089482_);
  or g_144747_(_086586_, _089482_, _089483_);
  xor g_144748_(_086588_, _089482_, _089484_);
  and g_144749_(_086591_, _089484_, _089485_);
  or g_144750_(_086591_, _089484_, _089486_);
  xor g_144751_(_086592_, _089484_, _089487_);
  or g_144752_(_083769_, _086596_, _089488_);
  and g_144753_(_086594_, _089488_, _089489_);
  xor g_144754_(_089487_, _089489_, _089491_);
  and g_144755_(_086807_, _089491_, _089492_);
  xor g_144756_(_086805_, _089491_, _089493_);
  not g_144757_(_089493_, _089494_);
  and g_144758_(_086803_, _089494_, _089495_);
  or g_144759_(_086804_, _089493_, _089496_);
  xor g_144760_(_086803_, _089493_, _089497_);
  not g_144761_(_089497_, _089498_);
  or g_144762_(_086800_, _089497_, _089499_);
  xor g_144763_(_086800_, _089498_, _089500_);
  not g_144764_(_089500_, _089502_);
  xor g_144765_(_086603_, _089500_, _089503_);
  xor g_144766_(_086617_, _089503_, _089504_);
  or g_144767_(_086798_, _089504_, _089505_);
  xor g_144768_(_086798_, _089504_, _089506_);
  not g_144769_(_089506_, _089507_);
  or g_144770_(_086797_, _089507_, _089508_);
  xor g_144771_(_086796_, _089506_, _089509_);
  xor g_144772_(_086797_, _089506_, _089510_);
  or g_144773_(_086626_, _089510_, _089511_);
  xor g_144774_(_086626_, _089509_, _089513_);
  or g_144775_(_086628_, _089513_, _089514_);
  xor g_144776_(_086629_, _089513_, _089515_);
  not g_144777_(_089515_, _089516_);
  xor g_144778_(_086638_, _089515_, _089517_);
  xor g_144779_(_086794_, _089517_, _089518_);
  not g_144780_(_089518_, _089519_);
  xor g_144781_(_086646_, _089518_, _089520_);
  and g_144782_(_086654_, _089520_, _089521_);
  and g_144783_(_086652_, _089518_, _089522_);
  or g_144784_(_089521_, _089522_, _089524_);
  not g_144785_(_089524_, _089525_);
  xor g_144786_(_086793_, _089525_, _089526_);
  not g_144787_(_089526_, _089527_);
  or g_144788_(_086661_, _089526_, _089528_);
  xor g_144789_(_086661_, _089526_, _089529_);
  and g_144790_(_086669_, _089529_, _089530_);
  and g_144791_(_083842_, _086670_, _089531_);
  not g_144792_(_089531_, _089532_);
  or g_144793_(_086665_, _089529_, _089533_);
  and g_144794_(_086665_, _089527_, _089535_);
  or g_144795_(_086666_, _089526_, _089536_);
  and g_144796_(_089533_, _089536_, _089537_);
  and g_144797_(_089531_, _089537_, _089538_);
  xor g_144798_(_089532_, _089537_, _089539_);
  and g_144799_(_086668_, _089539_, _089540_);
  or g_144800_(_089530_, _089540_, _089541_);
  or g_144801_(_086792_, _089541_, _089542_);
  not g_144802_(_089542_, _089543_);
  xor g_144803_(_086792_, _089541_, _089544_);
  xor g_144804_(_086676_, _089544_, _089546_);
  not g_144805_(_089546_, _089547_);
  and g_144806_(_086688_, _089547_, _089548_);
  not g_144807_(_089548_, _089549_);
  xor g_144808_(_086689_, _089546_, _089550_);
  and g_144809_(_086685_, _089550_, _089551_);
  xor g_144810_(_086687_, _089550_, _089552_);
  not g_144811_(_089552_, _089553_);
  and g_144812_(_086701_, _089553_, _089554_);
  xor g_144813_(_086702_, _089552_, _089555_);
  not g_144814_(_089555_, _089557_);
  or g_144815_(_083863_, _086706_, _089558_);
  and g_144816_(_086694_, _089558_, _089559_);
  xor g_144817_(_089555_, _089559_, _089560_);
  or g_144818_(_086791_, _089560_, _089561_);
  xor g_144819_(_086791_, _089560_, _089562_);
  not g_144820_(_089562_, _089563_);
  and g_144821_(_086713_, _086716_, _089564_);
  xor g_144822_(_089562_, _089564_, _089565_);
  or g_144823_(_086722_, _089565_, _089566_);
  xor g_144824_(_086721_, _089565_, _089568_);
  or g_144825_(_086718_, _089568_, _089569_);
  xor g_144826_(_086720_, _089568_, _089570_);
  or g_144827_(_083940_, _086724_, _089571_);
  not g_144828_(_089571_, _089572_);
  or g_144829_(_089570_, _089571_, _089573_);
  not g_144830_(_089573_, _089574_);
  xor g_144831_(_089570_, _089572_, _089575_);
  and g_144832_(_086731_, _086734_, _089576_);
  not g_144833_(_089576_, _089577_);
  xor g_144834_(_089575_, _089577_, _089579_);
  not g_144835_(_089579_, _089580_);
  or g_144836_(_086737_, _089579_, _089581_);
  xor g_144837_(_086737_, _089580_, _089582_);
  and g_144838_(_086739_, _089582_, _089583_);
  or g_144839_(_086739_, _089582_, _089584_);
  xor g_144840_(_086739_, _089582_, _089585_);
  or g_144841_(_086743_, _086754_, _089586_);
  xor g_144842_(_089585_, _089586_, _089587_);
  not g_144843_(_089587_, _089588_);
  and g_144844_(_086751_, _089587_, _089590_);
  xor g_144845_(_086751_, _089587_, _089591_);
  xor g_144846_(_086753_, _089587_, _089592_);
  and g_144847_(_086761_, _089592_, _089593_);
  or g_144848_(_086760_, _089591_, _089594_);
  and g_144849_(_086760_, _089587_, _089595_);
  or g_144850_(_086761_, _089588_, _089596_);
  and g_144851_(_089594_, _089596_, _089597_);
  or g_144852_(_089593_, _089595_, _089598_);
  and g_144853_(_086767_, _089597_, _089599_);
  or g_144854_(_086766_, _089598_, _089601_);
  xor g_144855_(_086767_, _089597_, _089602_);
  not g_144856_(_089602_, _089603_);
  and g_144857_(_086765_, _089602_, _089604_);
  or g_144858_(_086764_, _089603_, _089605_);
  xor g_144859_(_086764_, _089602_, _089606_);
  not g_144860_(_089606_, _089607_);
  and g_144861_(_086773_, _086777_, _089608_);
  xor g_144862_(_089607_, _089608_, _089609_);
  not g_144863_(_089609_, _089610_);
  and g_144864_(_086780_, _086786_, _089612_);
  xor g_144865_(_089610_, _089612_, _089613_);
  or g_144866_(_086784_, _089613_, _089614_);
  xor g_144867_(_086783_, _089613_, _089615_);
  or g_144868_(_086788_, _089615_, _089616_);
  xor g_144869_(_086788_, _089615_, out[965]);
  or g_144870_(_086786_, _089609_, _089617_);
  or g_144871_(_086780_, _089609_, _089618_);
  or g_144872_(_086777_, _089606_, _089619_);
  or g_144873_(_086773_, _089606_, _089620_);
  or g_144874_(_086734_, _089575_, _089622_);
  and g_144875_(_089581_, _089622_, _089623_);
  or g_144876_(_086731_, _089575_, _089624_);
  not g_144877_(_089624_, _089625_);
  or g_144878_(_086716_, _089563_, _089626_);
  not g_144879_(_089626_, _089627_);
  and g_144880_(_086712_, _089562_, _089628_);
  or g_144881_(_086713_, _089563_, _089629_);
  or g_144882_(_089557_, _089558_, _089630_);
  and g_144883_(_089561_, _089630_, _089631_);
  not g_144884_(_089631_, _089633_);
  and g_144885_(_086695_, _089555_, _089634_);
  or g_144886_(_086676_, _089541_, _089635_);
  not g_144887_(_089635_, _089636_);
  or g_144888_(_086659_, _089524_, _089637_);
  or g_144889_(_086657_, _089520_, _089638_);
  and g_144890_(_086650_, _089518_, _089639_);
  not g_144891_(_089639_, _089640_);
  and g_144892_(_083818_, _089639_, _089641_);
  or g_144893_(_083817_, _089640_, _089642_);
  and g_144894_(_083814_, _089639_, _089644_);
  or g_144895_(_086645_, _089519_, _089645_);
  or g_144896_(_080839_, _089645_, _089646_);
  not g_144897_(_089646_, _089647_);
  or g_144898_(_080834_, _089645_, _089648_);
  or g_144899_(_086647_, _089517_, _089649_);
  or g_144900_(_086643_, _089517_, _089650_);
  not g_144901_(_089650_, _089651_);
  and g_144902_(_086636_, _089516_, _089652_);
  or g_144903_(_086637_, _089515_, _089653_);
  and g_144904_(_089511_, _089514_, _089655_);
  and g_144905_(_086612_, _089502_, _089656_);
  or g_144906_(_086613_, _089500_, _089657_);
  or g_144907_(_086614_, _089500_, _089658_);
  not g_144908_(_089658_, _089659_);
  and g_144909_(_080795_, _086601_, _089660_);
  and g_144910_(_089502_, _089660_, _089661_);
  and g_144911_(_080791_, _086601_, _089662_);
  not g_144912_(_089662_, _089663_);
  and g_144913_(_089502_, _089662_, _089664_);
  or g_144914_(_089500_, _089663_, _089666_);
  or g_144915_(_089487_, _089488_, _089667_);
  not g_144916_(_089667_, _089668_);
  or g_144917_(_086572_, _089450_, _089669_);
  or g_144918_(_086570_, _089450_, _089670_);
  or g_144919_(_086547_, _089422_, _089671_);
  or g_144920_(_089389_, _089392_, _089672_);
  and g_144921_(_086507_, _089368_, _089673_);
  or g_144922_(_086506_, _089370_, _089674_);
  and g_144923_(_086504_, _089368_, _089675_);
  not g_144924_(_089675_, _089677_);
  and g_144925_(_089360_, _089363_, _089678_);
  or g_144926_(_089317_, _089319_, _089679_);
  not g_144927_(_089679_, _089680_);
  or g_144928_(_086465_, _089317_, _089681_);
  not g_144929_(_089681_, _089682_);
  or g_144930_(_089269_, _089271_, _089683_);
  not g_144931_(_089683_, _089684_);
  or g_144932_(_086423_, _089257_, _089685_);
  and g_144933_(_089262_, _089685_, _089686_);
  not g_144934_(_089686_, _089688_);
  and g_144935_(_086420_, _089256_, _089689_);
  or g_144936_(_086407_, _089250_, _089690_);
  or g_144937_(_086404_, _089246_, _089691_);
  not g_144938_(_089691_, _089692_);
  or g_144939_(_089242_, _089243_, _089693_);
  not g_144940_(_089693_, _089694_);
  or g_144941_(_086387_, _089230_, _089695_);
  and g_144942_(_086385_, _089229_, _089696_);
  and g_144943_(_086380_, _089223_, _089697_);
  and g_144944_(_089223_, _089227_, _089699_);
  not g_144945_(_089699_, _089700_);
  or g_144946_(_086359_, _089208_, _089701_);
  or g_144947_(_086357_, _089200_, _089702_);
  or g_144948_(_086353_, _089200_, _089703_);
  or g_144949_(_089184_, _089185_, _089704_);
  or g_144950_(_089184_, _089186_, _089705_);
  not g_144951_(_089705_, _089706_);
  and g_144952_(_089178_, _089181_, _089707_);
  or g_144953_(_089179_, _089180_, _089708_);
  or g_144954_(_089157_, _089161_, _089710_);
  or g_144955_(_089157_, _089159_, _089711_);
  or g_144956_(_089147_, _089148_, _089712_);
  or g_144957_(_086313_, _089144_, _089713_);
  not g_144958_(_089713_, _089714_);
  or g_144959_(_089131_, _089133_, _089715_);
  not g_144960_(_089715_, _089716_);
  or g_144961_(_089131_, _089134_, _089717_);
  or g_144962_(_086881_, _089098_, _089718_);
  or g_144963_(_086270_, _089098_, _089719_);
  and g_144964_(_086266_, _089095_, _089721_);
  or g_144965_(_086244_, _089074_, _089722_);
  and g_144966_(_089077_, _089722_, _089723_);
  not g_144967_(_089723_, _089724_);
  and g_144968_(_086240_, _089073_, _089725_);
  or g_144969_(_086239_, _089074_, _089726_);
  and g_144970_(_086236_, _089065_, _089727_);
  not g_144971_(_089727_, _089728_);
  and g_144972_(_086230_, _089065_, _089729_);
  or g_144973_(_086229_, _089066_, _089730_);
  or g_144974_(_083350_, _086217_, _089732_);
  not g_144975_(_089732_, _089733_);
  and g_144976_(_089051_, _089733_, _089734_);
  or g_144977_(_083347_, _086217_, _089735_);
  not g_144978_(_089735_, _089736_);
  and g_144979_(_089048_, _089736_, _089737_);
  not g_144980_(_089737_, _089738_);
  and g_144981_(_086204_, _089021_, _089739_);
  not g_144982_(_089739_, _089740_);
  or g_144983_(_086892_, _089022_, _089741_);
  or g_144984_(_089018_, _089019_, _089743_);
  or g_144985_(_086187_, _089003_, _089744_);
  not g_144986_(_089744_, _089745_);
  and g_144987_(_086181_, _089001_, _089746_);
  and g_144988_(_088969_, _088972_, _089747_);
  or g_144989_(_088970_, _088971_, _089748_);
  and g_144990_(_086160_, _088969_, _089749_);
  not g_144991_(_089749_, _089750_);
  and g_144992_(_088955_, _088957_, _089751_);
  and g_144993_(_088955_, _088959_, _089752_);
  not g_144994_(_089752_, _089754_);
  or g_144995_(_086118_, _088910_, _089755_);
  or g_144996_(_086115_, _088910_, _089756_);
  not g_144997_(_089756_, _089757_);
  and g_144998_(_086078_, _088880_, _089758_);
  and g_144999_(_088867_, _088872_, _089759_);
  and g_145000_(_088862_, _088865_, _089760_);
  not g_145001_(_089760_, _089761_);
  or g_145002_(_086055_, _088851_, _089762_);
  and g_145003_(_086050_, _088848_, _089763_);
  or g_145004_(_088843_, _088844_, _089765_);
  or g_145005_(_086039_, _088839_, _089766_);
  and g_145006_(_088807_, _088810_, _089767_);
  or g_145007_(_088787_, _088800_, _089768_);
  not g_145008_(_089768_, _089769_);
  and g_145009_(_088752_, _088755_, _089770_);
  not g_145010_(_089770_, _089771_);
  and g_145011_(_085951_, _088752_, _089772_);
  not g_145012_(_089772_, _089773_);
  or g_145013_(_088733_, _088735_, _089774_);
  or g_145014_(_088722_, _088724_, _089776_);
  not g_145015_(_089776_, _089777_);
  or g_145016_(_085922_, _088722_, _089778_);
  and g_145017_(_088721_, _089778_, _089779_);
  or g_145018_(_088697_, _088699_, _089780_);
  not g_145019_(_089780_, _089781_);
  or g_145020_(_086953_, _088691_, _089782_);
  or g_145021_(_085889_, _088691_, _089783_);
  or g_145022_(_085887_, _088690_, _089784_);
  and g_145023_(_085882_, _085885_, _089785_);
  or g_145024_(_088686_, _089785_, _089787_);
  or g_145025_(_085848_, _088655_, _089788_);
  or g_145026_(_082973_, _085825_, _089789_);
  or g_145027_(_088630_, _089789_, _089790_);
  not g_145028_(_089790_, _089791_);
  or g_145029_(_082970_, _085825_, _089792_);
  or g_145030_(_088626_, _089792_, _089793_);
  and g_145031_(_088606_, _088611_, _089794_);
  or g_145032_(_085794_, _088596_, _089795_);
  or g_145033_(_085792_, _088596_, _089796_);
  not g_145034_(_089796_, _089798_);
  or g_145035_(_085789_, _088591_, _089799_);
  not g_145036_(_089799_, _089800_);
  or g_145037_(_085780_, _088590_, _089801_);
  and g_145038_(_088589_, _089801_, _089802_);
  not g_145039_(_089802_, _089803_);
  or g_145040_(_085760_, _085761_, _089804_);
  not g_145041_(_089804_, _089805_);
  and g_145042_(_088579_, _089805_, _089806_);
  or g_145043_(_088580_, _089804_, _089807_);
  or g_145044_(_082919_, _085760_, _089809_);
  not g_145045_(_089809_, _089810_);
  and g_145046_(_088579_, _089810_, _089811_);
  and g_145047_(_088549_, _088553_, _089812_);
  and g_145048_(_088534_, _088536_, _089813_);
  not g_145049_(_089813_, _089814_);
  and g_145050_(_085723_, _088530_, _089815_);
  or g_145051_(_085722_, _088529_, _089816_);
  and g_145052_(_085720_, _088530_, _089817_);
  or g_145053_(_085711_, _088528_, _089818_);
  or g_145054_(_082867_, _089818_, _089820_);
  or g_145055_(_082864_, _089818_, _089821_);
  or g_145056_(_085683_, _088498_, _089822_);
  or g_145057_(_085675_, _088495_, _089823_);
  not g_145058_(_089823_, _089824_);
  or g_145059_(_085670_, _088495_, _089825_);
  or g_145060_(_085661_, _088494_, _089826_);
  not g_145061_(_089826_, _089827_);
  or g_145062_(_082829_, _089826_, _089828_);
  and g_145063_(_089825_, _089828_, _089829_);
  not g_145064_(_089829_, _089831_);
  and g_145065_(_085662_, _089827_, _089832_);
  or g_145066_(_085651_, _088482_, _089833_);
  or g_145067_(_085633_, _088470_, _089834_);
  not g_145068_(_089834_, _089835_);
  or g_145069_(_082796_, _085622_, _089836_);
  or g_145070_(_088469_, _089836_, _089837_);
  not g_145071_(_089837_, _089838_);
  or g_145072_(_082790_, _085622_, _089839_);
  or g_145073_(_088469_, _089839_, _089840_);
  not g_145074_(_089840_, _089842_);
  or g_145075_(_085591_, _088437_, _089843_);
  or g_145076_(_085588_, _088437_, _089844_);
  not g_145077_(_089844_, _089845_);
  and g_145078_(_088431_, _088433_, _089846_);
  and g_145079_(_088409_, _088411_, _089847_);
  or g_145080_(_088408_, _088413_, _089848_);
  or g_145081_(_088380_, _088382_, _089849_);
  and g_145082_(_088371_, _088374_, _089850_);
  not g_145083_(_089850_, _089851_);
  and g_145084_(_085483_, _088333_, _089853_);
  or g_145085_(_088328_, _088329_, _089854_);
  not g_145086_(_089854_, _089855_);
  or g_145087_(_088300_, _088301_, _089856_);
  not g_145088_(_089856_, _089857_);
  or g_145089_(_088287_, _088290_, _089858_);
  not g_145090_(_089858_, _089859_);
  or g_145091_(_085409_, _088264_, _089860_);
  not g_145092_(_089860_, _089861_);
  or g_145093_(_085336_, _088210_, _089862_);
  or g_145094_(_085338_, _088210_, _089864_);
  not g_145095_(_089864_, _089865_);
  and g_145096_(_085317_, _088204_, _089866_);
  not g_145097_(_089866_, _089867_);
  and g_145098_(_085319_, _088204_, _089868_);
  not g_145099_(_089868_, _089869_);
  or g_145100_(_085312_, _088201_, _089870_);
  or g_145101_(_082506_, _089870_, _089871_);
  not g_145102_(_089871_, _089872_);
  or g_145103_(_082504_, _089870_, _089873_);
  or g_145104_(_085309_, _088201_, _089875_);
  not g_145105_(_089875_, _089876_);
  and g_145106_(_088195_, _088198_, _089877_);
  not g_145107_(_089877_, _089878_);
  and g_145108_(_088171_, _088176_, _089879_);
  not g_145109_(_089879_, _089880_);
  or g_145110_(_085266_, _088156_, _089881_);
  not g_145111_(_089881_, _089882_);
  or g_145112_(_085264_, _088156_, _089883_);
  or g_145113_(_085240_, _088124_, _089884_);
  or g_145114_(_085231_, _088121_, _089886_);
  or g_145115_(_085233_, _088124_, _089887_);
  and g_145116_(_089886_, _089887_, _089888_);
  or g_145117_(_085229_, _088121_, _089889_);
  or g_145118_(_085215_, _088107_, _089890_);
  or g_145119_(_087032_, _088101_, _089891_);
  not g_145120_(_089891_, _089892_);
  or g_145121_(_085209_, _088101_, _089893_);
  not g_145122_(_089893_, _089894_);
  or g_145123_(_082387_, _085204_, _089895_);
  not g_145124_(_089895_, _089897_);
  and g_145125_(_088100_, _089897_, _089898_);
  and g_145126_(_088092_, _088096_, _089899_);
  not g_145127_(_089899_, _089900_);
  and g_145128_(_088077_, _088079_, _089901_);
  not g_145129_(_089901_, _089902_);
  and g_145130_(_085171_, _088063_, _089903_);
  and g_145131_(_085174_, _088063_, _089904_);
  or g_145132_(_085142_, _088035_, _089905_);
  and g_145133_(_088040_, _089905_, _089906_);
  or g_145134_(_087057_, _088011_, _089908_);
  or g_145135_(_085111_, _088010_, _089909_);
  not g_145136_(_089909_, _089910_);
  and g_145137_(_085104_, _088008_, _089911_);
  not g_145138_(_089911_, _089912_);
  or g_145139_(_087974_, _087975_, _089913_);
  not g_145140_(_089913_, _089914_);
  or g_145141_(_085056_, _087965_, _089915_);
  not g_145142_(_089915_, _089916_);
  or g_145143_(_085054_, _087965_, _089917_);
  and g_145144_(_087066_, _087934_, _089919_);
  or g_145145_(_085013_, _087933_, _089920_);
  or g_145146_(_085011_, _087930_, _089921_);
  or g_145147_(_085009_, _087930_, _089922_);
  not g_145148_(_089922_, _089923_);
  or g_145149_(_084998_, _087920_, _089924_);
  not g_145150_(_089924_, _089925_);
  or g_145151_(_084994_, _087920_, _089926_);
  not g_145152_(_089926_, _089927_);
  and g_145153_(_084976_, _087891_, _089928_);
  or g_145154_(_084975_, _087892_, _089930_);
  or g_145155_(_084967_, _087885_, _089931_);
  not g_145156_(_089931_, _089932_);
  or g_145157_(_087072_, _087885_, _089933_);
  not g_145158_(_089933_, _089934_);
  or g_145159_(_087880_, _087881_, _089935_);
  or g_145160_(_084962_, _087880_, _089936_);
  not g_145161_(_089936_, _089937_);
  and g_145162_(_087853_, _087859_, _089938_);
  and g_145163_(_087842_, _087846_, _089939_);
  not g_145164_(_089939_, _089941_);
  and g_145165_(_087842_, _087848_, _089942_);
  or g_145166_(_087838_, _087839_, _089943_);
  not g_145167_(_089943_, _089944_);
  or g_145168_(_084912_, _087815_, _089945_);
  or g_145169_(_084910_, _087811_, _089946_);
  and g_145170_(_087813_, _089946_, _089947_);
  or g_145171_(_084905_, _087802_, _089948_);
  or g_145172_(_084901_, _087802_, _089949_);
  not g_145173_(_089949_, _089950_);
  or g_145174_(_084889_, _087781_, _089952_);
  and g_145175_(_087784_, _089952_, _089953_);
  not g_145176_(_089953_, _089954_);
  or g_145177_(_084883_, _087781_, _089955_);
  or g_145178_(_082057_, _089955_, _089956_);
  or g_145179_(_082052_, _089955_, _089957_);
  or g_145180_(_087776_, _087778_, _089958_);
  or g_145181_(_087776_, _087777_, _089959_);
  and g_145182_(_087771_, _087775_, _089960_);
  not g_145183_(_089960_, _089961_);
  or g_145184_(_082025_, _084866_, _089963_);
  or g_145185_(_087766_, _089963_, _089964_);
  or g_145186_(_082026_, _084864_, _089965_);
  or g_145187_(_087766_, _089965_, _089966_);
  not g_145188_(_089966_, _089967_);
  or g_145189_(_084852_, _087756_, _089968_);
  or g_145190_(_082008_, _089968_, _089969_);
  not g_145191_(_089969_, _089970_);
  or g_145192_(_082006_, _089968_, _089971_);
  not g_145193_(_089971_, _089972_);
  or g_145194_(_084851_, _087754_, _089974_);
  not g_145195_(_089974_, _089975_);
  or g_145196_(_084841_, _087746_, _089976_);
  or g_145197_(_084832_, _087739_, _089977_);
  not g_145198_(_089977_, _089978_);
  or g_145199_(_084829_, _087739_, _089979_);
  and g_145200_(_084815_, _087711_, _089980_);
  or g_145201_(_084814_, _087712_, _089981_);
  or g_145202_(_087712_, _087713_, _089982_);
  not g_145203_(_089982_, _089983_);
  and g_145204_(_087696_, _087700_, _089985_);
  not g_145205_(_089985_, _089986_);
  or g_145206_(_084790_, _087690_, _089987_);
  or g_145207_(_084784_, _087688_, _089988_);
  and g_145208_(_087687_, _089988_, _089989_);
  not g_145209_(_089989_, _089990_);
  or g_145210_(_084779_, _087682_, _089991_);
  or g_145211_(_084776_, _087682_, _089992_);
  not g_145212_(_089992_, _089993_);
  and g_145213_(_087643_, _087648_, _089994_);
  or g_145214_(_081849_, _084730_, _089996_);
  or g_145215_(_087622_, _089996_, _089997_);
  and g_145216_(_087626_, _089997_, _089998_);
  and g_145217_(_084715_, _087604_, _089999_);
  and g_145218_(_084711_, _087601_, _090000_);
  or g_145219_(_084700_, _087599_, _090001_);
  or g_145220_(_084702_, _090001_, _090002_);
  or g_145221_(_081820_, _090001_, _090003_);
  not g_145222_(_090003_, _090004_);
  or g_145223_(_084688_, _087575_, _090005_);
  not g_145224_(_090005_, _090007_);
  or g_145225_(_084685_, _087575_, _090008_);
  not g_145226_(_090008_, _090009_);
  and g_145227_(_084639_, _087529_, _090010_);
  not g_145228_(_090010_, _090011_);
  or g_145229_(_084631_, _087520_, _090012_);
  not g_145230_(_090012_, _090013_);
  or g_145231_(_087520_, _087522_, _090014_);
  or g_145232_(_087516_, _087517_, _090015_);
  or g_145233_(_084624_, _087516_, _090016_);
  or g_145234_(_081739_, _084616_, _090018_);
  or g_145235_(_087514_, _090018_, _090019_);
  and g_145236_(_087513_, _090019_, _090020_);
  or g_145237_(_084606_, _087494_, _090021_);
  not g_145238_(_090021_, _090022_);
  and g_145239_(_087495_, _087497_, _090023_);
  or g_145240_(_081705_, _084590_, _090024_);
  or g_145241_(_087479_, _090024_, _090025_);
  or g_145242_(_084587_, _087473_, _090026_);
  not g_145243_(_090026_, _090027_);
  or g_145244_(_084560_, _087465_, _090029_);
  and g_145245_(_087438_, _087441_, _090030_);
  and g_145246_(_087414_, _087418_, _090031_);
  or g_145247_(_081619_, _084514_, _090032_);
  or g_145248_(_087397_, _090032_, _090033_);
  or g_145249_(_067914_, _090033_, _090034_);
  or g_145250_(_078742_, _081598_, _090035_);
  or g_145251_(_087392_, _090035_, _090036_);
  or g_145252_(_084503_, _090036_, _090037_);
  or g_145253_(_068025_, _090037_, _090038_);
  and g_145254_(_087395_, _090038_, _090040_);
  or g_145255_(_084491_, _087385_, _090041_);
  and g_145256_(_087380_, _087383_, _090042_);
  and g_145257_(_084487_, _087375_, _090043_);
  and g_145258_(_084478_, _087371_, _090044_);
  or g_145259_(_087373_, _090044_, _090045_);
  or g_145260_(_084472_, _087368_, _090046_);
  and g_145261_(_087366_, _090046_, _090047_);
  and g_145262_(_084462_, _087362_, _090048_);
  and g_145263_(_084463_, _087359_, _090049_);
  or g_145264_(_087358_, _090049_, _090051_);
  or g_145265_(_087346_, _087350_, _090052_);
  and g_145266_(_084430_, _087324_, _090053_);
  or g_145267_(_087317_, _090053_, _090054_);
  and g_145268_(_087310_, _087315_, _090055_);
  or g_145269_(_087311_, _090055_, _090056_);
  or g_145270_(_084397_, _087295_, _090057_);
  and g_145271_(_087281_, _087284_, _090058_);
  or g_145272_(_084378_, _087276_, _090059_);
  or g_145273_(_084374_, _087275_, _090060_);
  and g_145274_(_087274_, _090060_, _090062_);
  and g_145275_(_087179_, _087270_, _090063_);
  or g_145276_(_084370_, _087269_, _090064_);
  or g_145277_(_087184_, _087266_, _090065_);
  and g_145278_(_087265_, _090065_, _090066_);
  or g_145279_(_084366_, _087261_, _090067_);
  or g_145280_(_084361_, _087259_, _090068_);
  and g_145281_(_087260_, _090068_, _090069_);
  and g_145282_(_087241_, _087243_, _090070_);
  and g_145283_(_087249_, _090070_, _090071_);
  or g_145284_(_087192_, _087245_, _090073_);
  and g_145285_(_087251_, _090073_, _090074_);
  xor g_145286_(_090071_, _090074_, _090075_);
  or g_145287_(_087187_, _087255_, _090076_);
  and g_145288_(_087254_, _090076_, _090077_);
  xor g_145289_(_090075_, _090077_, _090078_);
  xor g_145290_(_090069_, _090078_, _090079_);
  xor g_145291_(_090067_, _090079_, _090080_);
  xor g_145292_(_090066_, _090080_, _090081_);
  xor g_145293_(_090064_, _090081_, _090082_);
  xor g_145294_(_090063_, _090082_, _090084_);
  xor g_145295_(_090062_, _090084_, _090085_);
  xor g_145296_(_090059_, _090085_, _090086_);
  xor g_145297_(_090058_, _090086_, _090087_);
  xor g_145298_(_090057_, _090087_, _090088_);
  and g_145299_(_084391_, _084394_, _090089_);
  or g_145300_(_087293_, _090089_, _090090_);
  and g_145301_(_087291_, _090090_, _090091_);
  xor g_145302_(_090088_, _090091_, _090092_);
  and g_145303_(_087298_, _087304_, _090093_);
  or g_145304_(_084412_, _087302_, _090095_);
  and g_145305_(_087306_, _090095_, _090096_);
  xor g_145306_(_090093_, _090096_, _090097_);
  xor g_145307_(_090092_, _090097_, _090098_);
  xor g_145308_(_090056_, _090098_, _090099_);
  xor g_145309_(_087320_, _090099_, _090100_);
  xor g_145310_(_090054_, _090100_, _090101_);
  xor g_145311_(_087329_, _090101_, _090102_);
  or g_145312_(_087333_, _090102_, _090103_);
  not g_145313_(_090103_, _090104_);
  or g_145314_(_087331_, _090102_, _090106_);
  and g_145315_(_087333_, _090106_, _090107_);
  not g_145316_(_090107_, _090108_);
  and g_145317_(_090103_, _090108_, _090109_);
  or g_145318_(_090104_, _090107_, _090110_);
  or g_145319_(_087337_, _090110_, _090111_);
  and g_145320_(_084443_, _090109_, _090112_);
  or g_145321_(_084445_, _087336_, _090113_);
  or g_145322_(_090112_, _090113_, _090114_);
  and g_145323_(_090111_, _090114_, _090115_);
  and g_145324_(_087168_, _087343_, _090117_);
  and g_145325_(_087339_, _087342_, _090118_);
  or g_145326_(_090117_, _090118_, _090119_);
  xor g_145327_(_090115_, _090119_, _090120_);
  xor g_145328_(_090052_, _090120_, _090121_);
  xor g_145329_(_090051_, _090121_, _090122_);
  xor g_145330_(_090048_, _090122_, _090123_);
  xor g_145331_(_090047_, _090123_, _090124_);
  xor g_145332_(_090045_, _090124_, _090125_);
  xor g_145333_(_090043_, _090125_, _090126_);
  xor g_145334_(_090042_, _090126_, _090128_);
  not g_145335_(_090128_, _090129_);
  or g_145336_(_087388_, _090129_, _090130_);
  and g_145337_(_087388_, _090129_, _090131_);
  xor g_145338_(_087388_, _090128_, _090132_);
  not g_145339_(_090132_, _090133_);
  xor g_145340_(_090041_, _090132_, _090134_);
  xor g_145341_(_090041_, _090133_, _090135_);
  xor g_145342_(_090040_, _090134_, _090136_);
  or g_145343_(_087398_, _090136_, _090137_);
  xor g_145344_(_087399_, _090136_, _090139_);
  and g_145345_(_090034_, _090139_, _090140_);
  or g_145346_(_090033_, _090139_, _090141_);
  or g_145347_(_067914_, _090141_, _090142_);
  not g_145348_(_090142_, _090143_);
  or g_145349_(_090140_, _090143_, _090144_);
  or g_145350_(_087410_, _090144_, _090145_);
  xor g_145351_(_087403_, _090144_, _090146_);
  and g_145352_(_087410_, _090146_, _090147_);
  not g_145353_(_090147_, _090148_);
  and g_145354_(_090145_, _090148_, _090150_);
  xor g_145355_(_090031_, _090150_, _090151_);
  or g_145356_(_087423_, _090151_, _090152_);
  xor g_145357_(_087421_, _090151_, _090153_);
  not g_145358_(_090153_, _090154_);
  or g_145359_(_087425_, _090153_, _090155_);
  xor g_145360_(_087425_, _090153_, _090156_);
  xor g_145361_(_087425_, _090154_, _090157_);
  and g_145362_(_087431_, _090157_, _090158_);
  or g_145363_(_087432_, _090156_, _090159_);
  or g_145364_(_087431_, _090153_, _090161_);
  and g_145365_(_090159_, _090161_, _090162_);
  xor g_145366_(_087435_, _090162_, _090163_);
  or g_145367_(_090030_, _090163_, _090164_);
  xor g_145368_(_090030_, _090163_, _090165_);
  and g_145369_(_087447_, _090165_, _090166_);
  xor g_145370_(_087447_, _090165_, _090167_);
  not g_145371_(_090167_, _090168_);
  or g_145372_(_087453_, _090168_, _090169_);
  and g_145373_(_087445_, _090167_, _090170_);
  xor g_145374_(_087443_, _090167_, _090172_);
  and g_145375_(_087453_, _090172_, _090173_);
  not g_145376_(_090173_, _090174_);
  and g_145377_(_090169_, _090174_, _090175_);
  xor g_145378_(_087457_, _090175_, _090176_);
  and g_145379_(_087460_, _090176_, _090177_);
  or g_145380_(_087460_, _090176_, _090178_);
  xor g_145381_(_087460_, _090176_, _090179_);
  xor g_145382_(_087461_, _090176_, _090180_);
  or g_145383_(_090029_, _090180_, _090181_);
  not g_145384_(_090181_, _090183_);
  xor g_145385_(_087464_, _090179_, _090184_);
  and g_145386_(_090029_, _090184_, _090185_);
  or g_145387_(_090183_, _090185_, _090186_);
  not g_145388_(_090186_, _090187_);
  or g_145389_(_087470_, _090186_, _090188_);
  or g_145390_(_084564_, _087465_, _090189_);
  not g_145391_(_090189_, _090190_);
  or g_145392_(_090187_, _090189_, _090191_);
  or g_145393_(_090186_, _090190_, _090192_);
  and g_145394_(_087470_, _090192_, _090194_);
  and g_145395_(_090191_, _090194_, _090195_);
  not g_145396_(_090195_, _090196_);
  and g_145397_(_090188_, _090196_, _090197_);
  or g_145398_(_084580_, _087473_, _090198_);
  not g_145399_(_090198_, _090199_);
  and g_145400_(_087472_, _090198_, _090200_);
  xor g_145401_(_090197_, _090200_, _090201_);
  or g_145402_(_090026_, _090201_, _090202_);
  and g_145403_(_090026_, _090201_, _090203_);
  xor g_145404_(_090027_, _090201_, _090205_);
  not g_145405_(_090205_, _090206_);
  or g_145406_(_081700_, _084590_, _090207_);
  or g_145407_(_087479_, _090207_, _090208_);
  and g_145408_(_087478_, _090208_, _090209_);
  xor g_145409_(_090206_, _090209_, _090210_);
  not g_145410_(_090210_, _090211_);
  or g_145411_(_090025_, _090210_, _090212_);
  xor g_145412_(_090025_, _090210_, _090213_);
  xor g_145413_(_090025_, _090211_, _090214_);
  and g_145414_(_087482_, _090214_, _090216_);
  or g_145415_(_087483_, _090213_, _090217_);
  or g_145416_(_087482_, _090210_, _090218_);
  not g_145417_(_090218_, _090219_);
  or g_145418_(_090216_, _090219_, _090220_);
  not g_145419_(_090220_, _090221_);
  or g_145420_(_087490_, _090220_, _090222_);
  and g_145421_(_087486_, _090220_, _090223_);
  or g_145422_(_087485_, _090221_, _090224_);
  and g_145423_(_087485_, _090218_, _090225_);
  not g_145424_(_090225_, _090227_);
  and g_145425_(_090217_, _090225_, _090228_);
  or g_145426_(_090216_, _090227_, _090229_);
  and g_145427_(_087490_, _090229_, _090230_);
  or g_145428_(_087491_, _090228_, _090231_);
  and g_145429_(_090224_, _090230_, _090232_);
  or g_145430_(_090223_, _090231_, _090233_);
  and g_145431_(_090222_, _090233_, _090234_);
  xor g_145432_(_087493_, _090234_, _090235_);
  not g_145433_(_090235_, _090236_);
  and g_145434_(_090023_, _090236_, _090238_);
  xor g_145435_(_090023_, _090235_, _090239_);
  and g_145436_(_090021_, _090239_, _090240_);
  or g_145437_(_090021_, _090239_, _090241_);
  xor g_145438_(_090022_, _090239_, _090242_);
  and g_145439_(_087502_, _087508_, _090243_);
  not g_145440_(_090243_, _090244_);
  xor g_145441_(_090242_, _090243_, _090245_);
  xor g_145442_(_090242_, _090244_, _090246_);
  or g_145443_(_090020_, _090246_, _090247_);
  xor g_145444_(_090020_, _090245_, _090249_);
  or g_145445_(_084616_, _087512_, _090250_);
  or g_145446_(_084617_, _090250_, _090251_);
  not g_145447_(_090251_, _090252_);
  or g_145448_(_090249_, _090251_, _090253_);
  xor g_145449_(_090249_, _090252_, _090254_);
  not g_145450_(_090254_, _090255_);
  or g_145451_(_090016_, _090254_, _090256_);
  xor g_145452_(_090016_, _090254_, _090257_);
  xor g_145453_(_090016_, _090255_, _090258_);
  or g_145454_(_090015_, _090258_, _090260_);
  xor g_145455_(_090015_, _090257_, _090261_);
  or g_145456_(_090014_, _090261_, _090262_);
  xor g_145457_(_090014_, _090261_, _090263_);
  and g_145458_(_090013_, _090263_, _090264_);
  xor g_145459_(_090012_, _090263_, _090265_);
  not g_145460_(_090265_, _090266_);
  and g_145461_(_087525_, _090266_, _090267_);
  xor g_145462_(_087525_, _090265_, _090268_);
  and g_145463_(_084636_, _087528_, _090269_);
  or g_145464_(_087527_, _090269_, _090271_);
  or g_145465_(_090268_, _090271_, _090272_);
  xor g_145466_(_090268_, _090271_, _090273_);
  and g_145467_(_090010_, _090273_, _090274_);
  xor g_145468_(_090011_, _090273_, _090275_);
  and g_145469_(_087533_, _087536_, _090276_);
  or g_145470_(_090275_, _090276_, _090277_);
  and g_145471_(_090275_, _090276_, _090278_);
  xor g_145472_(_090275_, _090276_, _090279_);
  xor g_145473_(_087539_, _090279_, _090280_);
  xor g_145474_(_087545_, _090280_, _090282_);
  or g_145475_(_087548_, _090282_, _090283_);
  xor g_145476_(_087549_, _090282_, _090284_);
  not g_145477_(_090284_, _090285_);
  and g_145478_(_087552_, _087555_, _090286_);
  or g_145479_(_090284_, _090286_, _090287_);
  xor g_145480_(_090284_, _090286_, _090288_);
  xor g_145481_(_090285_, _090286_, _090289_);
  or g_145482_(_087559_, _090289_, _090290_);
  xor g_145483_(_087559_, _090288_, _090291_);
  or g_145484_(_087566_, _090291_, _090293_);
  xor g_145485_(_087567_, _090291_, _090294_);
  or g_145486_(_087562_, _090294_, _090295_);
  xor g_145487_(_087562_, _090294_, _090296_);
  and g_145488_(_087573_, _090296_, _090297_);
  xor g_145489_(_087574_, _090296_, _090298_);
  or g_145490_(_090008_, _090298_, _090299_);
  xor g_145491_(_090009_, _090298_, _090300_);
  or g_145492_(_090005_, _090300_, _090301_);
  xor g_145493_(_090007_, _090300_, _090302_);
  and g_145494_(_087580_, _090302_, _090304_);
  or g_145495_(_087580_, _090302_, _090305_);
  xor g_145496_(_087581_, _090302_, _090306_);
  and g_145497_(_087583_, _087590_, _090307_);
  xor g_145498_(_090306_, _090307_, _090308_);
  not g_145499_(_090308_, _090309_);
  or g_145500_(_087592_, _090309_, _090310_);
  not g_145501_(_090310_, _090311_);
  xor g_145502_(_087592_, _090308_, _090312_);
  or g_145503_(_087596_, _090312_, _090313_);
  xor g_145504_(_087596_, _090312_, _090315_);
  not g_145505_(_090315_, _090316_);
  and g_145506_(_090004_, _090315_, _090317_);
  or g_145507_(_090003_, _090316_, _090318_);
  xor g_145508_(_090003_, _090315_, _090319_);
  and g_145509_(_090002_, _090319_, _090320_);
  or g_145510_(_090002_, _090319_, _090321_);
  xor g_145511_(_090002_, _090319_, _090322_);
  xor g_145512_(_087603_, _090322_, _090323_);
  or g_145513_(_090000_, _090323_, _090324_);
  and g_145514_(_090000_, _090323_, _090326_);
  xor g_145515_(_090000_, _090323_, _090327_);
  xor g_145516_(_089999_, _090327_, _090328_);
  or g_145517_(_087608_, _090328_, _090329_);
  and g_145518_(_087608_, _090328_, _090330_);
  xor g_145519_(_087608_, _090328_, _090331_);
  xor g_145520_(_087610_, _090328_, _090332_);
  and g_145521_(_087614_, _087618_, _090333_);
  or g_145522_(_087616_, _090333_, _090334_);
  xor g_145523_(_090331_, _090334_, _090335_);
  or g_145524_(_089998_, _090335_, _090337_);
  not g_145525_(_090337_, _090338_);
  and g_145526_(_087624_, _090335_, _090339_);
  and g_145527_(_087626_, _090339_, _090340_);
  or g_145528_(_090338_, _090340_, _090341_);
  and g_145529_(_087630_, _090341_, _090342_);
  or g_145530_(_087630_, _090341_, _090343_);
  xor g_145531_(_087630_, _090341_, _090344_);
  xor g_145532_(_087629_, _090341_, _090345_);
  or g_145533_(_087633_, _090345_, _090346_);
  or g_145534_(_087634_, _090344_, _090348_);
  and g_145535_(_087636_, _090348_, _090349_);
  and g_145536_(_090346_, _090349_, _090350_);
  or g_145537_(_087636_, _090345_, _090351_);
  not g_145538_(_090351_, _090352_);
  or g_145539_(_090350_, _090352_, _090353_);
  xor g_145540_(_087645_, _090353_, _090354_);
  xor g_145541_(_087644_, _090353_, _090355_);
  or g_145542_(_089994_, _090355_, _090356_);
  xor g_145543_(_089994_, _090354_, _090357_);
  and g_145544_(_087651_, _090357_, _090359_);
  or g_145545_(_087651_, _090357_, _090360_);
  xor g_145546_(_087652_, _090357_, _090361_);
  not g_145547_(_090361_, _090362_);
  and g_145548_(_087656_, _087659_, _090363_);
  xor g_145549_(_090361_, _090363_, _090364_);
  xor g_145550_(_090362_, _090363_, _090365_);
  or g_145551_(_087661_, _090365_, _090366_);
  xor g_145552_(_087661_, _090364_, _090367_);
  and g_145553_(_087670_, _090367_, _090368_);
  and g_145554_(_087669_, _090364_, _090370_);
  or g_145555_(_087670_, _090365_, _090371_);
  or g_145556_(_090368_, _090370_, _090372_);
  xor g_145557_(_087667_, _090372_, _090373_);
  or g_145558_(_087673_, _090373_, _090374_);
  and g_145559_(_087673_, _090373_, _090375_);
  xor g_145560_(_087673_, _090373_, _090376_);
  or g_145561_(_087120_, _087678_, _090377_);
  and g_145562_(_087677_, _090377_, _090378_);
  xor g_145563_(_090376_, _090378_, _090379_);
  and g_145564_(_089992_, _090379_, _090381_);
  or g_145565_(_089992_, _090379_, _090382_);
  xor g_145566_(_089993_, _090379_, _090383_);
  xor g_145567_(_089991_, _090383_, _090384_);
  and g_145568_(_089990_, _090384_, _090385_);
  xor g_145569_(_089989_, _090384_, _090386_);
  and g_145570_(_089987_, _090386_, _090387_);
  or g_145571_(_089987_, _090386_, _090388_);
  xor g_145572_(_089987_, _090386_, _090389_);
  xor g_145573_(_087693_, _090389_, _090390_);
  or g_145574_(_089985_, _090390_, _090392_);
  xor g_145575_(_089985_, _090390_, _090393_);
  xor g_145576_(_089986_, _090390_, _090394_);
  or g_145577_(_087704_, _090394_, _090395_);
  xor g_145578_(_087704_, _090393_, _090396_);
  not g_145579_(_090396_, _090397_);
  or g_145580_(_087707_, _090396_, _090398_);
  xor g_145581_(_087707_, _090396_, _090399_);
  xor g_145582_(_087707_, _090397_, _090400_);
  and g_145583_(_087710_, _090400_, _090401_);
  or g_145584_(_087710_, _090400_, _090403_);
  xor g_145585_(_087710_, _090399_, _090404_);
  xor g_145586_(_089982_, _090404_, _090405_);
  xor g_145587_(_089983_, _090404_, _090406_);
  or g_145588_(_089980_, _090405_, _090407_);
  or g_145589_(_089981_, _090404_, _090408_);
  not g_145590_(_090408_, _090409_);
  and g_145591_(_090407_, _090408_, _090410_);
  or g_145592_(_087722_, _090410_, _090411_);
  or g_145593_(_087721_, _090406_, _090412_);
  or g_145594_(_090409_, _090412_, _090414_);
  and g_145595_(_090411_, _090414_, _090415_);
  and g_145596_(_087717_, _090415_, _090416_);
  xor g_145597_(_087716_, _090415_, _090417_);
  or g_145598_(_087725_, _090417_, _090418_);
  xor g_145599_(_087726_, _090417_, _090419_);
  not g_145600_(_090419_, _090420_);
  or g_145601_(_087729_, _090419_, _090421_);
  xor g_145602_(_087729_, _090419_, _090422_);
  xor g_145603_(_087729_, _090420_, _090423_);
  and g_145604_(_087734_, _090423_, _090425_);
  or g_145605_(_087733_, _090422_, _090426_);
  and g_145606_(_087733_, _090420_, _090427_);
  or g_145607_(_087734_, _090419_, _090428_);
  and g_145608_(_090426_, _090428_, _090429_);
  or g_145609_(_090425_, _090427_, _090430_);
  or g_145610_(_089979_, _090430_, _090431_);
  not g_145611_(_090431_, _090432_);
  or g_145612_(_087737_, _090427_, _090433_);
  or g_145613_(_090425_, _090433_, _090434_);
  or g_145614_(_087738_, _090429_, _090436_);
  and g_145615_(_089979_, _090436_, _090437_);
  and g_145616_(_090434_, _090437_, _090438_);
  or g_145617_(_090432_, _090438_, _090439_);
  xor g_145618_(_089978_, _090439_, _090440_);
  xor g_145619_(_089977_, _090439_, _090441_);
  and g_145620_(_087744_, _090440_, _090442_);
  or g_145621_(_087745_, _090441_, _090443_);
  or g_145622_(_084837_, _087743_, _090444_);
  not g_145623_(_090444_, _090445_);
  and g_145624_(_090442_, _090444_, _090447_);
  or g_145625_(_090443_, _090445_, _090448_);
  or g_145626_(_087744_, _090439_, _090449_);
  and g_145627_(_090444_, _090449_, _090450_);
  not g_145628_(_090450_, _090451_);
  and g_145629_(_090443_, _090451_, _090452_);
  or g_145630_(_090442_, _090450_, _090453_);
  and g_145631_(_090448_, _090453_, _090454_);
  or g_145632_(_090447_, _090452_, _090455_);
  or g_145633_(_089976_, _090455_, _090456_);
  xor g_145634_(_089976_, _090455_, _090458_);
  xor g_145635_(_089976_, _090454_, _090459_);
  or g_145636_(_084845_, _087751_, _090460_);
  and g_145637_(_087750_, _090460_, _090461_);
  not g_145638_(_090461_, _090462_);
  and g_145639_(_090458_, _090462_, _090463_);
  not g_145640_(_090463_, _090464_);
  xor g_145641_(_090459_, _090461_, _090465_);
  and g_145642_(_089975_, _090465_, _090466_);
  xor g_145643_(_089975_, _090465_, _090467_);
  and g_145644_(_089972_, _090467_, _090469_);
  xor g_145645_(_089971_, _090467_, _090470_);
  or g_145646_(_089969_, _090470_, _090471_);
  and g_145647_(_089969_, _090470_, _090472_);
  xor g_145648_(_089970_, _090470_, _090473_);
  not g_145649_(_090473_, _090474_);
  and g_145650_(_087764_, _090474_, _090475_);
  or g_145651_(_087765_, _090473_, _090476_);
  xor g_145652_(_087759_, _090473_, _090477_);
  or g_145653_(_087764_, _090477_, _090478_);
  and g_145654_(_090476_, _090478_, _090480_);
  xor g_145655_(_089966_, _090480_, _090481_);
  not g_145656_(_090481_, _090482_);
  or g_145657_(_089964_, _090481_, _090483_);
  xor g_145658_(_089964_, _090481_, _090484_);
  xor g_145659_(_089964_, _090482_, _090485_);
  or g_145660_(_087768_, _090485_, _090486_);
  xor g_145661_(_087768_, _090484_, _090487_);
  or g_145662_(_089960_, _090487_, _090488_);
  xor g_145663_(_089961_, _090487_, _090489_);
  or g_145664_(_089959_, _090489_, _090491_);
  and g_145665_(_089959_, _090489_, _090492_);
  xor g_145666_(_089959_, _090489_, _090493_);
  xor g_145667_(_089958_, _090493_, _090494_);
  or g_145668_(_089957_, _090494_, _090495_);
  and g_145669_(_089957_, _090494_, _090496_);
  xor g_145670_(_089957_, _090494_, _090497_);
  xor g_145671_(_089956_, _090497_, _090498_);
  or g_145672_(_089953_, _090498_, _090499_);
  xor g_145673_(_089954_, _090498_, _090500_);
  and g_145674_(_087788_, _090500_, _090502_);
  or g_145675_(_087788_, _090500_, _090503_);
  xor g_145676_(_087788_, _090500_, _090504_);
  not g_145677_(_090504_, _090505_);
  and g_145678_(_087794_, _090504_, _090506_);
  or g_145679_(_087793_, _090505_, _090507_);
  xor g_145680_(_087791_, _090504_, _090508_);
  and g_145681_(_087793_, _090508_, _090509_);
  or g_145682_(_090506_, _090509_, _090510_);
  not g_145683_(_090510_, _090511_);
  and g_145684_(_087799_, _090511_, _090513_);
  or g_145685_(_087800_, _090510_, _090514_);
  xor g_145686_(_087797_, _090510_, _090515_);
  or g_145687_(_087799_, _090515_, _090516_);
  and g_145688_(_090514_, _090516_, _090517_);
  xor g_145689_(_089949_, _090517_, _090518_);
  xor g_145690_(_089948_, _090518_, _090519_);
  xor g_145691_(_087806_, _090519_, _090520_);
  not g_145692_(_090520_, _090521_);
  xor g_145693_(_087810_, _090520_, _090522_);
  xor g_145694_(_087810_, _090521_, _090524_);
  xor g_145695_(_089947_, _090522_, _090525_);
  or g_145696_(_089945_, _090525_, _090526_);
  and g_145697_(_089945_, _090525_, _090527_);
  xor g_145698_(_089945_, _090525_, _090528_);
  xor g_145699_(_087819_, _090528_, _090529_);
  or g_145700_(_087822_, _090529_, _090530_);
  and g_145701_(_087822_, _090529_, _090531_);
  xor g_145702_(_087822_, _090529_, _090532_);
  and g_145703_(_087825_, _087830_, _090533_);
  xor g_145704_(_090532_, _090533_, _090535_);
  or g_145705_(_084939_, _087835_, _090536_);
  and g_145706_(_087836_, _090536_, _090537_);
  or g_145707_(_090535_, _090537_, _090538_);
  and g_145708_(_090535_, _090537_, _090539_);
  xor g_145709_(_090535_, _090537_, _090540_);
  xor g_145710_(_089944_, _090540_, _090541_);
  and g_145711_(_089942_, _090541_, _090542_);
  or g_145712_(_089942_, _090541_, _090543_);
  xor g_145713_(_089942_, _090541_, _090544_);
  xor g_145714_(_089941_, _090544_, _090546_);
  or g_145715_(_089938_, _090546_, _090547_);
  xor g_145716_(_089938_, _090546_, _090548_);
  or g_145717_(_087856_, _090548_, _090549_);
  and g_145718_(_087856_, _090548_, _090550_);
  xor g_145719_(_087857_, _090548_, _090551_);
  and g_145720_(_087868_, _087870_, _090552_);
  xor g_145721_(_090551_, _090552_, _090553_);
  or g_145722_(_087872_, _090553_, _090554_);
  not g_145723_(_090554_, _090555_);
  and g_145724_(_087872_, _090553_, _090557_);
  not g_145725_(_090557_, _090558_);
  and g_145726_(_090554_, _090558_, _090559_);
  or g_145727_(_090555_, _090557_, _090560_);
  or g_145728_(_087877_, _090559_, _090561_);
  or g_145729_(_087876_, _090557_, _090562_);
  or g_145730_(_090555_, _090562_, _090563_);
  and g_145731_(_087879_, _090563_, _090564_);
  and g_145732_(_090561_, _090564_, _090565_);
  or g_145733_(_087879_, _090560_, _090566_);
  not g_145734_(_090566_, _090568_);
  or g_145735_(_090565_, _090568_, _090569_);
  xor g_145736_(_089937_, _090569_, _090570_);
  and g_145737_(_089935_, _090570_, _090571_);
  or g_145738_(_089935_, _090569_, _090572_);
  not g_145739_(_090572_, _090573_);
  or g_145740_(_090571_, _090573_, _090574_);
  xor g_145741_(_089934_, _090574_, _090575_);
  and g_145742_(_089931_, _090575_, _090576_);
  or g_145743_(_089931_, _090575_, _090577_);
  xor g_145744_(_089931_, _090575_, _090579_);
  xor g_145745_(_089932_, _090575_, _090580_);
  and g_145746_(_087888_, _087893_, _090581_);
  or g_145747_(_087889_, _090581_, _090582_);
  xor g_145748_(_090580_, _090582_, _090583_);
  and g_145749_(_089928_, _090583_, _090584_);
  xor g_145750_(_089930_, _090583_, _090585_);
  and g_145751_(_087902_, _090585_, _090586_);
  or g_145752_(_087902_, _090585_, _090587_);
  xor g_145753_(_087903_, _090585_, _090588_);
  not g_145754_(_090588_, _090590_);
  and g_145755_(_087908_, _090590_, _090591_);
  or g_145756_(_087909_, _090588_, _090592_);
  xor g_145757_(_087898_, _090588_, _090593_);
  or g_145758_(_087908_, _090593_, _090594_);
  not g_145759_(_090594_, _090595_);
  and g_145760_(_090592_, _090594_, _090596_);
  or g_145761_(_090591_, _090595_, _090597_);
  and g_145762_(_087911_, _087915_, _090598_);
  xor g_145763_(_090596_, _090598_, _090599_);
  or g_145764_(_087919_, _090599_, _090601_);
  xor g_145765_(_087919_, _090599_, _090602_);
  and g_145766_(_089927_, _090602_, _090603_);
  xor g_145767_(_089926_, _090602_, _090604_);
  or g_145768_(_089924_, _090604_, _090605_);
  and g_145769_(_089924_, _090604_, _090606_);
  xor g_145770_(_089925_, _090604_, _090607_);
  not g_145771_(_090607_, _090608_);
  xor g_145772_(_087924_, _090608_, _090609_);
  xor g_145773_(_087924_, _090607_, _090610_);
  or g_145774_(_089922_, _090609_, _090612_);
  and g_145775_(_087929_, _090609_, _090613_);
  or g_145776_(_087927_, _090610_, _090614_);
  and g_145777_(_087927_, _090608_, _090615_);
  or g_145778_(_087929_, _090607_, _090616_);
  and g_145779_(_090614_, _090616_, _090617_);
  or g_145780_(_090613_, _090615_, _090618_);
  and g_145781_(_089922_, _090618_, _090619_);
  or g_145782_(_089923_, _090617_, _090620_);
  and g_145783_(_090612_, _090620_, _090621_);
  xor g_145784_(_089921_, _090621_, _090623_);
  or g_145785_(_089920_, _090623_, _090624_);
  xor g_145786_(_089920_, _090623_, _090625_);
  and g_145787_(_089919_, _090625_, _090626_);
  or g_145788_(_089919_, _090625_, _090627_);
  xor g_145789_(_089919_, _090625_, _090628_);
  xor g_145790_(_087938_, _090628_, _090629_);
  or g_145791_(_087942_, _090629_, _090630_);
  and g_145792_(_087942_, _090628_, _090631_);
  not g_145793_(_090631_, _090632_);
  and g_145794_(_090630_, _090632_, _090634_);
  not g_145795_(_090634_, _090635_);
  xor g_145796_(_087949_, _090634_, _090636_);
  and g_145797_(_087947_, _090636_, _090637_);
  and g_145798_(_087948_, _090634_, _090638_);
  or g_145799_(_087947_, _090635_, _090639_);
  or g_145800_(_090637_, _090638_, _090640_);
  not g_145801_(_090640_, _090641_);
  and g_145802_(_087956_, _087958_, _090642_);
  xor g_145803_(_090640_, _090642_, _090643_);
  xor g_145804_(_090641_, _090642_, _090645_);
  and g_145805_(_087964_, _090643_, _090646_);
  or g_145806_(_087963_, _090645_, _090647_);
  or g_145807_(_087960_, _090645_, _090648_);
  xor g_145808_(_087960_, _090643_, _090649_);
  and g_145809_(_087963_, _090649_, _090650_);
  or g_145810_(_090646_, _090650_, _090651_);
  not g_145811_(_090651_, _090652_);
  xor g_145812_(_089917_, _090651_, _090653_);
  xor g_145813_(_089917_, _090652_, _090654_);
  and g_145814_(_089915_, _090654_, _090656_);
  or g_145815_(_089916_, _090653_, _090657_);
  or g_145816_(_089915_, _090651_, _090658_);
  not g_145817_(_090658_, _090659_);
  and g_145818_(_090657_, _090658_, _090660_);
  or g_145819_(_090656_, _090659_, _090661_);
  xor g_145820_(_087969_, _090660_, _090662_);
  xor g_145821_(_087969_, _090661_, _090663_);
  or g_145822_(_085067_, _087971_, _090664_);
  and g_145823_(_087973_, _090664_, _090665_);
  not g_145824_(_090665_, _090667_);
  and g_145825_(_090663_, _090667_, _090668_);
  xor g_145826_(_090662_, _090667_, _090669_);
  and g_145827_(_089913_, _090669_, _090670_);
  or g_145828_(_089913_, _090669_, _090671_);
  xor g_145829_(_089914_, _090669_, _090672_);
  and g_145830_(_087979_, _087981_, _090673_);
  not g_145831_(_090673_, _090674_);
  xor g_145832_(_090672_, _090674_, _090675_);
  or g_145833_(_087982_, _090675_, _090676_);
  xor g_145834_(_087982_, _090675_, _090678_);
  and g_145835_(_087987_, _090678_, _090679_);
  xor g_145836_(_087987_, _090678_, _090680_);
  and g_145837_(_087989_, _090680_, _090681_);
  xor g_145838_(_087990_, _090680_, _090682_);
  or g_145839_(_087999_, _090682_, _090683_);
  xor g_145840_(_087998_, _090682_, _090684_);
  and g_145841_(_088003_, _088007_, _090685_);
  or g_145842_(_090684_, _090685_, _090686_);
  xor g_145843_(_090684_, _090685_, _090687_);
  and g_145844_(_089911_, _090687_, _090689_);
  or g_145845_(_089911_, _090687_, _090690_);
  xor g_145846_(_089911_, _090687_, _090691_);
  xor g_145847_(_089912_, _090687_, _090692_);
  or g_145848_(_089909_, _090692_, _090693_);
  not g_145849_(_090693_, _090694_);
  and g_145850_(_085108_, _088008_, _090695_);
  not g_145851_(_090695_, _090696_);
  and g_145852_(_090692_, _090695_, _090697_);
  not g_145853_(_090697_, _090698_);
  and g_145854_(_090691_, _090696_, _090700_);
  or g_145855_(_090692_, _090695_, _090701_);
  and g_145856_(_089909_, _090701_, _090702_);
  or g_145857_(_089910_, _090700_, _090703_);
  and g_145858_(_090698_, _090702_, _090704_);
  or g_145859_(_090697_, _090703_, _090705_);
  or g_145860_(_090694_, _090704_, _090706_);
  or g_145861_(_085115_, _088010_, _090707_);
  or g_145862_(_085118_, _088011_, _090708_);
  and g_145863_(_090707_, _090708_, _090709_);
  not g_145864_(_090709_, _090711_);
  and g_145865_(_090706_, _090709_, _090712_);
  and g_145866_(_090705_, _090711_, _090713_);
  and g_145867_(_090693_, _090713_, _090714_);
  or g_145868_(_090712_, _090714_, _090715_);
  and g_145869_(_089908_, _090715_, _090716_);
  or g_145870_(_089908_, _090715_, _090717_);
  xor g_145871_(_089908_, _090715_, _090718_);
  and g_145872_(_088014_, _088020_, _090719_);
  xor g_145873_(_090718_, _090719_, _090720_);
  or g_145874_(_088025_, _090720_, _090722_);
  and g_145875_(_088025_, _090720_, _090723_);
  xor g_145876_(_088025_, _090720_, _090724_);
  xor g_145877_(_088029_, _090724_, _090725_);
  or g_145878_(_088031_, _090725_, _090726_);
  xor g_145879_(_088031_, _090725_, _090727_);
  or g_145880_(_085139_, _088034_, _090728_);
  and g_145881_(_088033_, _090728_, _090729_);
  not g_145882_(_090729_, _090730_);
  and g_145883_(_090727_, _090730_, _090731_);
  xor g_145884_(_090727_, _090729_, _090733_);
  and g_145885_(_089906_, _090733_, _090734_);
  or g_145886_(_089906_, _090733_, _090735_);
  xor g_145887_(_089906_, _090733_, _090736_);
  xor g_145888_(_088046_, _090736_, _090737_);
  and g_145889_(_088048_, _090737_, _090738_);
  or g_145890_(_088048_, _090737_, _090739_);
  xor g_145891_(_088048_, _090737_, _090740_);
  not g_145892_(_090740_, _090741_);
  and g_145893_(_088052_, _090740_, _090742_);
  not g_145894_(_090742_, _090744_);
  or g_145895_(_088052_, _090740_, _090745_);
  and g_145896_(_088054_, _090745_, _090746_);
  and g_145897_(_090744_, _090746_, _090747_);
  or g_145898_(_088054_, _090741_, _090748_);
  not g_145899_(_090748_, _090749_);
  or g_145900_(_090747_, _090749_, _090750_);
  or g_145901_(_087044_, _088057_, _090751_);
  and g_145902_(_088056_, _090751_, _090752_);
  not g_145903_(_090752_, _090753_);
  xor g_145904_(_090750_, _090753_, _090755_);
  or g_145905_(_088062_, _090755_, _090756_);
  xor g_145906_(_088062_, _090755_, _090757_);
  and g_145907_(_089904_, _090757_, _090758_);
  xor g_145908_(_089904_, _090757_, _090759_);
  and g_145909_(_089903_, _090759_, _090760_);
  or g_145910_(_089903_, _090759_, _090761_);
  xor g_145911_(_089903_, _090759_, _090762_);
  xor g_145912_(_088070_, _090762_, _090763_);
  and g_145913_(_088068_, _090763_, _090764_);
  or g_145914_(_088068_, _090763_, _090766_);
  xor g_145915_(_088068_, _090763_, _090767_);
  xor g_145916_(_088075_, _090767_, _090768_);
  or g_145917_(_089901_, _090768_, _090769_);
  xor g_145918_(_089902_, _090768_, _090770_);
  or g_145919_(_088083_, _090770_, _090771_);
  and g_145920_(_088083_, _090770_, _090772_);
  xor g_145921_(_088084_, _090770_, _090773_);
  not g_145922_(_090773_, _090774_);
  and g_145923_(_088087_, _088089_, _090775_);
  xor g_145924_(_090774_, _090775_, _090777_);
  or g_145925_(_089899_, _090777_, _090778_);
  xor g_145926_(_089899_, _090777_, _090779_);
  xor g_145927_(_089900_, _090777_, _090780_);
  or g_145928_(_082383_, _085204_, _090781_);
  or g_145929_(_088099_, _090781_, _090782_);
  and g_145930_(_088098_, _090782_, _090783_);
  or g_145931_(_090780_, _090783_, _090784_);
  xor g_145932_(_090779_, _090783_, _090785_);
  not g_145933_(_090785_, _090786_);
  and g_145934_(_089898_, _090786_, _090788_);
  xor g_145935_(_089898_, _090785_, _090789_);
  or g_145936_(_089893_, _090789_, _090790_);
  xor g_145937_(_089894_, _090789_, _090791_);
  or g_145938_(_089891_, _090791_, _090792_);
  xor g_145939_(_089892_, _090791_, _090793_);
  or g_145940_(_089890_, _090793_, _090794_);
  not g_145941_(_090794_, _090795_);
  or g_145942_(_088105_, _090793_, _090796_);
  xor g_145943_(_088106_, _090793_, _090797_);
  and g_145944_(_089890_, _090797_, _090799_);
  or g_145945_(_090795_, _090799_, _090800_);
  not g_145946_(_090800_, _090801_);
  or g_145947_(_088112_, _090800_, _090802_);
  not g_145948_(_090802_, _090803_);
  or g_145949_(_085218_, _088107_, _090804_);
  not g_145950_(_090804_, _090805_);
  or g_145951_(_090801_, _090804_, _090806_);
  or g_145952_(_090800_, _090805_, _090807_);
  and g_145953_(_088112_, _090807_, _090808_);
  and g_145954_(_090806_, _090808_, _090810_);
  or g_145955_(_090803_, _090810_, _090811_);
  not g_145956_(_090811_, _090812_);
  or g_145957_(_088118_, _090811_, _090813_);
  xor g_145958_(_088116_, _090811_, _090814_);
  xor g_145959_(_088116_, _090812_, _090815_);
  and g_145960_(_088118_, _090815_, _090816_);
  or g_145961_(_088119_, _090814_, _090817_);
  and g_145962_(_090813_, _090817_, _090818_);
  xor g_145963_(_089889_, _090818_, _090819_);
  or g_145964_(_089888_, _090819_, _090821_);
  xor g_145965_(_089888_, _090819_, _090822_);
  not g_145966_(_090822_, _090823_);
  or g_145967_(_089884_, _090823_, _090824_);
  xor g_145968_(_089884_, _090822_, _090825_);
  or g_145969_(_088135_, _090825_, _090826_);
  not g_145970_(_090826_, _090827_);
  or g_145971_(_088129_, _090825_, _090828_);
  xor g_145972_(_088130_, _090825_, _090829_);
  and g_145973_(_088135_, _090829_, _090830_);
  or g_145974_(_090827_, _090830_, _090832_);
  not g_145975_(_090832_, _090833_);
  xor g_145976_(_088138_, _090833_, _090834_);
  xor g_145977_(_088138_, _090832_, _090835_);
  and g_145978_(_088141_, _090834_, _090836_);
  or g_145979_(_088142_, _090835_, _090837_);
  or g_145980_(_088141_, _090832_, _090838_);
  and g_145981_(_090837_, _090838_, _090839_);
  xor g_145982_(_088144_, _090839_, _090840_);
  xor g_145983_(_088145_, _090839_, _090841_);
  and g_145984_(_088149_, _090840_, _090843_);
  or g_145985_(_088147_, _090841_, _090844_);
  and g_145986_(_088147_, _090839_, _090845_);
  not g_145987_(_090845_, _090846_);
  or g_145988_(_088152_, _090845_, _090847_);
  not g_145989_(_090847_, _090848_);
  and g_145990_(_090844_, _090848_, _090849_);
  not g_145991_(_090849_, _090850_);
  and g_145992_(_090844_, _090846_, _090851_);
  or g_145993_(_090843_, _090845_, _090852_);
  or g_145994_(_088153_, _090851_, _090854_);
  and g_145995_(_088155_, _090854_, _090855_);
  and g_145996_(_090850_, _090855_, _090856_);
  or g_145997_(_088155_, _090852_, _090857_);
  not g_145998_(_090857_, _090858_);
  or g_145999_(_090856_, _090858_, _090859_);
  xor g_146000_(_089883_, _090859_, _090860_);
  and g_146001_(_089882_, _090860_, _090861_);
  xor g_146002_(_089882_, _090860_, _090862_);
  and g_146003_(_088162_, _090862_, _090863_);
  or g_146004_(_088162_, _090862_, _090865_);
  xor g_146005_(_088163_, _090862_, _090866_);
  not g_146006_(_090866_, _090867_);
  or g_146007_(_088165_, _088168_, _090868_);
  xor g_146008_(_090867_, _090868_, _090869_);
  and g_146009_(_089880_, _090869_, _090870_);
  xor g_146010_(_089879_, _090869_, _090871_);
  and g_146011_(_088184_, _088187_, _090872_);
  not g_146012_(_090872_, _090873_);
  or g_146013_(_090871_, _090872_, _090874_);
  xor g_146014_(_090871_, _090873_, _090876_);
  and g_146015_(_088190_, _088193_, _090877_);
  or g_146016_(_090876_, _090877_, _090878_);
  xor g_146017_(_090876_, _090877_, _090879_);
  and g_146018_(_089878_, _090879_, _090880_);
  xor g_146019_(_089878_, _090879_, _090881_);
  xor g_146020_(_089877_, _090879_, _090882_);
  or g_146021_(_089875_, _090882_, _090883_);
  or g_146022_(_088200_, _090882_, _090884_);
  xor g_146023_(_088200_, _090882_, _090885_);
  xor g_146024_(_088200_, _090881_, _090887_);
  and g_146025_(_089875_, _090887_, _090888_);
  or g_146026_(_089876_, _090885_, _090889_);
  and g_146027_(_090883_, _090889_, _090890_);
  xor g_146028_(_089873_, _090890_, _090891_);
  or g_146029_(_089871_, _090891_, _090892_);
  xor g_146030_(_089872_, _090891_, _090893_);
  or g_146031_(_089869_, _090893_, _090894_);
  and g_146032_(_089869_, _090893_, _090895_);
  xor g_146033_(_089869_, _090893_, _090896_);
  xor g_146034_(_089866_, _090896_, _090898_);
  and g_146035_(_088207_, _090898_, _090899_);
  xor g_146036_(_088207_, _090898_, _090900_);
  or g_146037_(_088209_, _090900_, _090901_);
  and g_146038_(_088209_, _090898_, _090902_);
  not g_146039_(_090902_, _090903_);
  and g_146040_(_090901_, _090903_, _090904_);
  xor g_146041_(_089864_, _090904_, _090905_);
  or g_146042_(_089862_, _090905_, _090906_);
  xor g_146043_(_089862_, _090905_, _090907_);
  not g_146044_(_090907_, _090909_);
  or g_146045_(_085353_, _088210_, _090910_);
  and g_146046_(_088213_, _090910_, _090911_);
  or g_146047_(_090909_, _090911_, _090912_);
  xor g_146048_(_090907_, _090911_, _090913_);
  or g_146049_(_088217_, _090913_, _090914_);
  xor g_146050_(_088217_, _090913_, _090915_);
  xor g_146051_(_088216_, _090913_, _090916_);
  and g_146052_(_088218_, _090915_, _090917_);
  or g_146053_(_088218_, _090915_, _090918_);
  xor g_146054_(_088218_, _090916_, _090920_);
  or g_146055_(_088223_, _088227_, _090921_);
  xor g_146056_(_090920_, _090921_, _090922_);
  or g_146057_(_088231_, _090922_, _090923_);
  xor g_146058_(_088232_, _090922_, _090924_);
  or g_146059_(_088235_, _090924_, _090925_);
  and g_146060_(_088235_, _090924_, _090926_);
  xor g_146061_(_088235_, _090924_, _090927_);
  and g_146062_(_088238_, _088241_, _090928_);
  xor g_146063_(_090927_, _090928_, _090929_);
  or g_146064_(_088245_, _090929_, _090931_);
  and g_146065_(_088245_, _090929_, _090932_);
  xor g_146066_(_088245_, _090929_, _090933_);
  not g_146067_(_090933_, _090934_);
  and g_146068_(_088249_, _088251_, _090935_);
  xor g_146069_(_090934_, _090935_, _090936_);
  and g_146070_(_088256_, _090936_, _090937_);
  or g_146071_(_088256_, _090936_, _090938_);
  xor g_146072_(_088256_, _090936_, _090939_);
  xor g_146073_(_088259_, _090939_, _090940_);
  or g_146074_(_088262_, _090940_, _090942_);
  and g_146075_(_088262_, _090939_, _090943_);
  not g_146076_(_090943_, _090944_);
  and g_146077_(_090942_, _090944_, _090945_);
  xor g_146078_(_089861_, _090945_, _090946_);
  or g_146079_(_085412_, _088264_, _090947_);
  and g_146080_(_088270_, _090947_, _090948_);
  not g_146081_(_090948_, _090949_);
  and g_146082_(_090946_, _090949_, _090950_);
  xor g_146083_(_090946_, _090948_, _090951_);
  and g_146084_(_088267_, _090951_, _090953_);
  or g_146085_(_088267_, _090951_, _090954_);
  xor g_146086_(_088267_, _090951_, _090955_);
  xor g_146087_(_088272_, _090955_, _090956_);
  or g_146088_(_088278_, _090956_, _090957_);
  not g_146089_(_090957_, _090958_);
  and g_146090_(_088278_, _090956_, _090959_);
  xor g_146091_(_088278_, _090956_, _090960_);
  and g_146092_(_088283_, _088288_, _090961_);
  or g_146093_(_088282_, _088289_, _090962_);
  and g_146094_(_088284_, _090962_, _090964_);
  or g_146095_(_088285_, _090961_, _090965_);
  or g_146096_(_090960_, _090964_, _090966_);
  or g_146097_(_090959_, _090965_, _090967_);
  or g_146098_(_090958_, _090967_, _090968_);
  and g_146099_(_090966_, _090968_, _090969_);
  and g_146100_(_089859_, _090969_, _090970_);
  xor g_146101_(_089858_, _090969_, _090971_);
  or g_146102_(_088294_, _090971_, _090972_);
  xor g_146103_(_088294_, _090971_, _090973_);
  or g_146104_(_088296_, _090973_, _090975_);
  or g_146105_(_088297_, _090971_, _090976_);
  and g_146106_(_090975_, _090976_, _090977_);
  or g_146107_(_085445_, _088300_, _090978_);
  not g_146108_(_090978_, _090979_);
  or g_146109_(_088299_, _090979_, _090980_);
  not g_146110_(_090980_, _090981_);
  and g_146111_(_090977_, _090980_, _090982_);
  xor g_146112_(_090977_, _090981_, _090983_);
  or g_146113_(_089856_, _090983_, _090984_);
  xor g_146114_(_089856_, _090983_, _090986_);
  xor g_146115_(_089857_, _090983_, _090987_);
  and g_146116_(_088305_, _090986_, _090988_);
  and g_146117_(_088306_, _090987_, _090989_);
  or g_146118_(_088305_, _090986_, _090990_);
  xor g_146119_(_088305_, _090986_, _090991_);
  or g_146120_(_088309_, _090991_, _090992_);
  and g_146121_(_088309_, _090990_, _090993_);
  or g_146122_(_088310_, _090989_, _090994_);
  or g_146123_(_090988_, _090994_, _090995_);
  and g_146124_(_090992_, _090995_, _090997_);
  or g_146125_(_088312_, _090997_, _090998_);
  and g_146126_(_088312_, _090991_, _090999_);
  not g_146127_(_090999_, _091000_);
  and g_146128_(_090998_, _091000_, _091001_);
  xor g_146129_(_088321_, _091001_, _091002_);
  or g_146130_(_088316_, _091002_, _091003_);
  xor g_146131_(_088317_, _091002_, _091004_);
  or g_146132_(_088325_, _091004_, _091005_);
  and g_146133_(_088325_, _091004_, _091006_);
  xor g_146134_(_088325_, _091004_, _091008_);
  not g_146135_(_091008_, _091009_);
  or g_146136_(_085473_, _088328_, _091010_);
  not g_146137_(_091010_, _091011_);
  and g_146138_(_088327_, _091010_, _091012_);
  xor g_146139_(_091009_, _091012_, _091013_);
  and g_146140_(_089855_, _091013_, _091014_);
  xor g_146141_(_089855_, _091013_, _091015_);
  xor g_146142_(_089854_, _091013_, _091016_);
  or g_146143_(_088332_, _091015_, _091017_);
  and g_146144_(_088332_, _091015_, _091019_);
  xor g_146145_(_088332_, _091015_, _091020_);
  xor g_146146_(_088332_, _091016_, _091021_);
  or g_146147_(_089853_, _091021_, _091022_);
  not g_146148_(_091022_, _091023_);
  and g_146149_(_089853_, _091021_, _091024_);
  and g_146150_(_085492_, _088333_, _091025_);
  or g_146151_(_091024_, _091025_, _091026_);
  or g_146152_(_091023_, _091026_, _091027_);
  and g_146153_(_091020_, _091025_, _091028_);
  not g_146154_(_091028_, _091030_);
  and g_146155_(_091027_, _091030_, _091031_);
  and g_146156_(_088338_, _091031_, _091032_);
  not g_146157_(_091032_, _091033_);
  or g_146158_(_088338_, _091031_, _091034_);
  and g_146159_(_085500_, _088339_, _091035_);
  not g_146160_(_091035_, _091036_);
  and g_146161_(_091034_, _091036_, _091037_);
  and g_146162_(_091033_, _091037_, _091038_);
  or g_146163_(_085496_, _088340_, _091039_);
  and g_146164_(_091031_, _091035_, _091041_);
  not g_146165_(_091041_, _091042_);
  and g_146166_(_091039_, _091042_, _091043_);
  or g_146167_(_091038_, _091043_, _091044_);
  not g_146168_(_091044_, _091045_);
  and g_146169_(_091038_, _091039_, _091046_);
  or g_146170_(_091045_, _091046_, _091047_);
  or g_146171_(_088352_, _091047_, _091048_);
  not g_146172_(_091048_, _091049_);
  or g_146173_(_088345_, _091047_, _091050_);
  xor g_146174_(_088344_, _091047_, _091052_);
  or g_146175_(_088353_, _091052_, _091053_);
  xor g_146176_(_088353_, _091052_, _091054_);
  xor g_146177_(_088354_, _091052_, _091055_);
  and g_146178_(_088352_, _091055_, _091056_);
  or g_146179_(_088351_, _091054_, _091057_);
  and g_146180_(_091048_, _091057_, _091058_);
  or g_146181_(_091049_, _091056_, _091059_);
  and g_146182_(_088359_, _091059_, _091060_);
  and g_146183_(_088360_, _091048_, _091061_);
  and g_146184_(_091057_, _091061_, _091063_);
  or g_146185_(_088364_, _091063_, _091064_);
  or g_146186_(_091060_, _091064_, _091065_);
  and g_146187_(_088364_, _091058_, _091066_);
  not g_146188_(_091066_, _091067_);
  and g_146189_(_091065_, _091067_, _091068_);
  xor g_146190_(_088365_, _091068_, _091069_);
  or g_146191_(_089850_, _091069_, _091070_);
  xor g_146192_(_089851_, _091069_, _091071_);
  or g_146193_(_085540_, _088378_, _091072_);
  and g_146194_(_088377_, _091072_, _091074_);
  or g_146195_(_091071_, _091074_, _091075_);
  xor g_146196_(_091071_, _091074_, _091076_);
  not g_146197_(_091076_, _091077_);
  or g_146198_(_089849_, _091077_, _091078_);
  xor g_146199_(_089849_, _091076_, _091079_);
  and g_146200_(_088386_, _091079_, _091080_);
  not g_146201_(_091080_, _091081_);
  or g_146202_(_088386_, _091079_, _091082_);
  and g_146203_(_088388_, _091082_, _091083_);
  and g_146204_(_091081_, _091083_, _091085_);
  and g_146205_(_088389_, _091079_, _091086_);
  or g_146206_(_091085_, _091086_, _091087_);
  xor g_146207_(_088397_, _091087_, _091088_);
  and g_146208_(_088398_, _091088_, _091089_);
  xor g_146209_(_088398_, _091088_, _091090_);
  xor g_146210_(_088399_, _091088_, _091091_);
  or g_146211_(_088405_, _091091_, _091092_);
  xor g_146212_(_088405_, _091090_, _091093_);
  or g_146213_(_089847_, _091093_, _091094_);
  xor g_146214_(_089848_, _091093_, _091096_);
  or g_146215_(_088418_, _091096_, _091097_);
  and g_146216_(_088418_, _091096_, _091098_);
  xor g_146217_(_088418_, _091096_, _091099_);
  xor g_146218_(_088420_, _091099_, _091100_);
  and g_146219_(_088424_, _091100_, _091101_);
  or g_146220_(_088424_, _091100_, _091102_);
  xor g_146221_(_088424_, _091100_, _091103_);
  xor g_146222_(_088428_, _091103_, _091104_);
  or g_146223_(_089846_, _091104_, _091105_);
  xor g_146224_(_089846_, _091104_, _091107_);
  and g_146225_(_088436_, _091107_, _091108_);
  or g_146226_(_088436_, _091107_, _091109_);
  xor g_146227_(_088436_, _091107_, _091110_);
  xor g_146228_(_089844_, _091110_, _091111_);
  or g_146229_(_089843_, _091111_, _091112_);
  xor g_146230_(_089843_, _091111_, _091113_);
  or g_146231_(_088440_, _091113_, _091114_);
  and g_146232_(_088440_, _091113_, _091115_);
  xor g_146233_(_088441_, _091113_, _091116_);
  and g_146234_(_086992_, _088446_, _091118_);
  or g_146235_(_088444_, _091118_, _091119_);
  xor g_146236_(_091116_, _091119_, _091120_);
  or g_146237_(_088450_, _091120_, _091121_);
  and g_146238_(_088450_, _091120_, _091122_);
  xor g_146239_(_088451_, _091120_, _091123_);
  and g_146240_(_088455_, _088458_, _091124_);
  not g_146241_(_091124_, _091125_);
  xor g_146242_(_091123_, _091125_, _091126_);
  not g_146243_(_091126_, _091127_);
  and g_146244_(_088464_, _091127_, _091129_);
  or g_146245_(_088460_, _091126_, _091130_);
  xor g_146246_(_088461_, _091126_, _091131_);
  and g_146247_(_088465_, _091131_, _091132_);
  or g_146248_(_091129_, _091132_, _091133_);
  and g_146249_(_088468_, _091133_, _091134_);
  or g_146250_(_088468_, _091131_, _091135_);
  not g_146251_(_091135_, _091136_);
  or g_146252_(_091134_, _091136_, _091137_);
  xor g_146253_(_089842_, _091137_, _091138_);
  or g_146254_(_089837_, _091138_, _091140_);
  xor g_146255_(_089837_, _091138_, _091141_);
  xor g_146256_(_089838_, _091138_, _091142_);
  and g_146257_(_089835_, _091141_, _091143_);
  or g_146258_(_089834_, _091142_, _091144_);
  or g_146259_(_085628_, _088470_, _091145_);
  not g_146260_(_091145_, _091146_);
  or g_146261_(_091138_, _091145_, _091147_);
  not g_146262_(_091147_, _091148_);
  and g_146263_(_091142_, _091145_, _091149_);
  or g_146264_(_091141_, _091146_, _091151_);
  and g_146265_(_091147_, _091151_, _091152_);
  or g_146266_(_091148_, _091149_, _091153_);
  and g_146267_(_088474_, _091152_, _091154_);
  or g_146268_(_088473_, _091153_, _091155_);
  and g_146269_(_091144_, _091155_, _091156_);
  or g_146270_(_091143_, _091154_, _091157_);
  and g_146271_(_089834_, _091153_, _091158_);
  and g_146272_(_088473_, _091158_, _091159_);
  or g_146273_(_091157_, _091159_, _091160_);
  not g_146274_(_091160_, _091162_);
  or g_146275_(_088477_, _091160_, _091163_);
  xor g_146276_(_088477_, _091160_, _091164_);
  xor g_146277_(_088477_, _091162_, _091165_);
  and g_146278_(_085639_, _088481_, _091166_);
  or g_146279_(_088480_, _091166_, _091167_);
  or g_146280_(_091165_, _091167_, _091168_);
  xor g_146281_(_091164_, _091167_, _091169_);
  or g_146282_(_089833_, _091169_, _091170_);
  xor g_146283_(_089833_, _091169_, _091171_);
  and g_146284_(_088485_, _091171_, _091173_);
  or g_146285_(_088485_, _091171_, _091174_);
  xor g_146286_(_088485_, _091171_, _091175_);
  xor g_146287_(_088488_, _091175_, _091176_);
  xor g_146288_(_088487_, _091175_, _091177_);
  and g_146289_(_088493_, _091177_, _091178_);
  and g_146290_(_088492_, _091175_, _091179_);
  or g_146291_(_091178_, _091179_, _091180_);
  xor g_146292_(_089832_, _091180_, _091181_);
  or g_146293_(_089829_, _091181_, _091182_);
  xor g_146294_(_089831_, _091181_, _091184_);
  and g_146295_(_089823_, _091184_, _091185_);
  or g_146296_(_089823_, _091184_, _091186_);
  xor g_146297_(_089823_, _091184_, _091187_);
  xor g_146298_(_089824_, _091184_, _091188_);
  or g_146299_(_089822_, _091188_, _091189_);
  not g_146300_(_091189_, _091190_);
  xor g_146301_(_088497_, _091187_, _091191_);
  and g_146302_(_089822_, _091191_, _091192_);
  or g_146303_(_091190_, _091192_, _091193_);
  or g_146304_(_088506_, _091193_, _091195_);
  not g_146305_(_091195_, _091196_);
  or g_146306_(_085686_, _088498_, _091197_);
  not g_146307_(_091197_, _091198_);
  xor g_146308_(_091193_, _091198_, _091199_);
  and g_146309_(_088506_, _091199_, _091200_);
  or g_146310_(_091196_, _091200_, _091201_);
  not g_146311_(_091201_, _091202_);
  xor g_146312_(_088505_, _091201_, _091203_);
  or g_146313_(_088512_, _091203_, _091204_);
  and g_146314_(_088512_, _091202_, _091206_);
  or g_146315_(_088513_, _091201_, _091207_);
  and g_146316_(_091204_, _091207_, _091208_);
  and g_146317_(_088516_, _088526_, _091209_);
  xor g_146318_(_091208_, _091209_, _091210_);
  or g_146319_(_088524_, _091210_, _091211_);
  xor g_146320_(_088524_, _091210_, _091212_);
  xor g_146321_(_088523_, _091210_, _091213_);
  or g_146322_(_089821_, _091213_, _091214_);
  xor g_146323_(_089821_, _091212_, _091215_);
  or g_146324_(_089820_, _091215_, _091217_);
  xor g_146325_(_089820_, _091215_, _091218_);
  and g_146326_(_089817_, _091218_, _091219_);
  or g_146327_(_089817_, _091218_, _091220_);
  xor g_146328_(_089817_, _091218_, _091221_);
  xor g_146329_(_089816_, _091221_, _091222_);
  or g_146330_(_089813_, _091222_, _091223_);
  xor g_146331_(_089814_, _091222_, _091224_);
  or g_146332_(_088540_, _091224_, _091225_);
  and g_146333_(_088540_, _091224_, _091226_);
  xor g_146334_(_088541_, _091224_, _091228_);
  not g_146335_(_091228_, _091229_);
  and g_146336_(_088542_, _088547_, _091230_);
  xor g_146337_(_091228_, _091230_, _091231_);
  xor g_146338_(_091229_, _091230_, _091232_);
  or g_146339_(_089812_, _091232_, _091233_);
  xor g_146340_(_089812_, _091231_, _091234_);
  and g_146341_(_088557_, _091234_, _091235_);
  or g_146342_(_088557_, _091234_, _091236_);
  xor g_146343_(_088558_, _091234_, _091237_);
  xor g_146344_(_088561_, _091237_, _091239_);
  xor g_146345_(_088560_, _091237_, _091240_);
  and g_146346_(_088565_, _091240_, _091241_);
  xor g_146347_(_088565_, _091239_, _091242_);
  and g_146348_(_088569_, _091242_, _091243_);
  or g_146349_(_088569_, _091239_, _091244_);
  not g_146350_(_091244_, _091245_);
  or g_146351_(_091243_, _091245_, _091246_);
  or g_146352_(_085756_, _088572_, _091247_);
  and g_146353_(_088571_, _091247_, _091248_);
  xor g_146354_(_091246_, _091248_, _091250_);
  and g_146355_(_088578_, _091250_, _091251_);
  xor g_146356_(_088578_, _091250_, _091252_);
  or g_146357_(_089811_, _091252_, _091253_);
  and g_146358_(_089811_, _091250_, _091254_);
  not g_146359_(_091254_, _091255_);
  and g_146360_(_091253_, _091255_, _091256_);
  not g_146361_(_091256_, _091257_);
  xor g_146362_(_089807_, _091256_, _091258_);
  and g_146363_(_088582_, _091258_, _091259_);
  and g_146364_(_088583_, _091256_, _091261_);
  or g_146365_(_088582_, _091257_, _091262_);
  or g_146366_(_091259_, _091261_, _091263_);
  xor g_146367_(_088586_, _091263_, _091264_);
  or g_146368_(_089802_, _091264_, _091265_);
  xor g_146369_(_089803_, _091264_, _091266_);
  or g_146370_(_089799_, _091266_, _091267_);
  and g_146371_(_089799_, _091266_, _091268_);
  xor g_146372_(_089799_, _091266_, _091269_);
  xor g_146373_(_089800_, _091266_, _091270_);
  and g_146374_(_089798_, _091269_, _091272_);
  or g_146375_(_089796_, _091270_, _091273_);
  xor g_146376_(_088595_, _091269_, _091274_);
  and g_146377_(_089796_, _091274_, _091275_);
  or g_146378_(_091272_, _091275_, _091276_);
  xor g_146379_(_089795_, _091276_, _091277_);
  xor g_146380_(_088602_, _091277_, _091278_);
  not g_146381_(_091278_, _091279_);
  xor g_146382_(_089794_, _091278_, _091280_);
  and g_146383_(_088612_, _091280_, _091281_);
  not g_146384_(_091281_, _091283_);
  and g_146385_(_088613_, _091278_, _091284_);
  or g_146386_(_088612_, _091279_, _091285_);
  and g_146387_(_091283_, _091285_, _091286_);
  or g_146388_(_091281_, _091284_, _091287_);
  and g_146389_(_088620_, _091286_, _091288_);
  not g_146390_(_091288_, _091289_);
  and g_146391_(_088617_, _091286_, _091290_);
  and g_146392_(_088618_, _091287_, _091291_);
  or g_146393_(_088620_, _091291_, _091292_);
  or g_146394_(_091290_, _091292_, _091294_);
  and g_146395_(_091289_, _091294_, _091295_);
  xor g_146396_(_088625_, _091295_, _091296_);
  or g_146397_(_088628_, _091296_, _091297_);
  xor g_146398_(_088628_, _091296_, _091298_);
  xor g_146399_(_088629_, _091296_, _091299_);
  or g_146400_(_089793_, _091299_, _091300_);
  xor g_146401_(_089793_, _091298_, _091301_);
  or g_146402_(_089790_, _091301_, _091302_);
  xor g_146403_(_089791_, _091301_, _091303_);
  not g_146404_(_091303_, _091305_);
  or g_146405_(_088636_, _091303_, _091306_);
  xor g_146406_(_088636_, _091303_, _091307_);
  xor g_146407_(_088636_, _091305_, _091308_);
  or g_146408_(_088639_, _091308_, _091309_);
  xor g_146409_(_088639_, _091307_, _091310_);
  and g_146410_(_088641_, _088644_, _091311_);
  not g_146411_(_091311_, _091312_);
  or g_146412_(_091310_, _091311_, _091313_);
  xor g_146413_(_091310_, _091311_, _091314_);
  xor g_146414_(_091310_, _091312_, _091316_);
  or g_146415_(_088647_, _091316_, _091317_);
  and g_146416_(_088647_, _091316_, _091318_);
  or g_146417_(_088648_, _091314_, _091319_);
  xor g_146418_(_088647_, _091314_, _091320_);
  and g_146419_(_085842_, _088651_, _091321_);
  or g_146420_(_088652_, _091321_, _091322_);
  not g_146421_(_091322_, _091323_);
  and g_146422_(_091320_, _091322_, _091324_);
  and g_146423_(_091319_, _091323_, _091325_);
  or g_146424_(_091318_, _091322_, _091327_);
  and g_146425_(_091317_, _091325_, _091328_);
  or g_146426_(_091324_, _091328_, _091329_);
  or g_146427_(_089788_, _091329_, _091330_);
  and g_146428_(_089788_, _091329_, _091331_);
  xor g_146429_(_089788_, _091329_, _091332_);
  or g_146430_(_088659_, _088661_, _091333_);
  xor g_146431_(_091332_, _091333_, _091334_);
  and g_146432_(_088662_, _091334_, _091335_);
  xor g_146433_(_088663_, _091334_, _091336_);
  and g_146434_(_088669_, _091336_, _091338_);
  or g_146435_(_088669_, _091336_, _091339_);
  xor g_146436_(_088669_, _091336_, _091340_);
  and g_146437_(_088672_, _091340_, _091341_);
  not g_146438_(_091341_, _091342_);
  or g_146439_(_088672_, _091340_, _091343_);
  not g_146440_(_091343_, _091344_);
  and g_146441_(_088677_, _091343_, _091345_);
  or g_146442_(_088675_, _091344_, _091346_);
  and g_146443_(_091342_, _091345_, _091347_);
  or g_146444_(_091341_, _091346_, _091349_);
  and g_146445_(_088675_, _091340_, _091350_);
  not g_146446_(_091350_, _091351_);
  and g_146447_(_091349_, _091351_, _091352_);
  or g_146448_(_091347_, _091350_, _091353_);
  and g_146449_(_085877_, _088682_, _091354_);
  or g_146450_(_088680_, _091354_, _091355_);
  xor g_146451_(_091353_, _091355_, _091356_);
  or g_146452_(_089787_, _091356_, _091357_);
  and g_146453_(_089787_, _091356_, _091358_);
  xor g_146454_(_089787_, _091356_, _091360_);
  xor g_146455_(_089784_, _091360_, _091361_);
  and g_146456_(_089783_, _091361_, _091362_);
  or g_146457_(_089783_, _091361_, _091363_);
  xor g_146458_(_089783_, _091361_, _091364_);
  xor g_146459_(_089782_, _091364_, _091365_);
  or g_146460_(_085897_, _088695_, _091366_);
  not g_146461_(_091366_, _091367_);
  or g_146462_(_088694_, _091367_, _091368_);
  or g_146463_(_091365_, _091368_, _091369_);
  xor g_146464_(_091365_, _091368_, _091371_);
  or g_146465_(_089781_, _091371_, _091372_);
  and g_146466_(_089781_, _091371_, _091373_);
  xor g_146467_(_089780_, _091371_, _091374_);
  or g_146468_(_088707_, _088713_, _091375_);
  not g_146469_(_091375_, _091376_);
  or g_146470_(_088708_, _091375_, _091377_);
  not g_146471_(_091377_, _091378_);
  xor g_146472_(_091374_, _091378_, _091379_);
  xor g_146473_(_088716_, _091379_, _091380_);
  xor g_146474_(_088715_, _091379_, _091382_);
  xor g_146475_(_089779_, _091380_, _091383_);
  and g_146476_(_089776_, _091383_, _091384_);
  or g_146477_(_089776_, _091383_, _091385_);
  xor g_146478_(_089777_, _091383_, _091386_);
  and g_146479_(_088728_, _088730_, _091387_);
  xor g_146480_(_091386_, _091387_, _091388_);
  and g_146481_(_089774_, _091388_, _091389_);
  xor g_146482_(_089774_, _091388_, _091390_);
  and g_146483_(_088740_, _091390_, _091391_);
  or g_146484_(_088740_, _091390_, _091393_);
  xor g_146485_(_088741_, _091390_, _091394_);
  xor g_146486_(_088743_, _091394_, _091395_);
  or g_146487_(_088748_, _091395_, _091396_);
  xor g_146488_(_088749_, _091395_, _091397_);
  not g_146489_(_091397_, _091398_);
  or g_146490_(_088751_, _091397_, _091399_);
  xor g_146491_(_088751_, _091397_, _091400_);
  or g_146492_(_089772_, _091400_, _091401_);
  and g_146493_(_089772_, _091398_, _091402_);
  or g_146494_(_089773_, _091397_, _091404_);
  and g_146495_(_091401_, _091404_, _091405_);
  xor g_146496_(_089771_, _091405_, _091406_);
  or g_146497_(_088760_, _091406_, _091407_);
  xor g_146498_(_088760_, _091406_, _091408_);
  and g_146499_(_088763_, _091408_, _091409_);
  xor g_146500_(_088762_, _091408_, _091410_);
  not g_146501_(_091410_, _091411_);
  and g_146502_(_088766_, _091411_, _091412_);
  xor g_146503_(_088767_, _091410_, _091413_);
  and g_146504_(_088770_, _088773_, _091415_);
  not g_146505_(_091415_, _091416_);
  and g_146506_(_091413_, _091416_, _091417_);
  xor g_146507_(_091413_, _091416_, _091418_);
  not g_146508_(_091418_, _091419_);
  and g_146509_(_088781_, _091418_, _091420_);
  or g_146510_(_088780_, _091419_, _091421_);
  and g_146511_(_088778_, _091418_, _091422_);
  xor g_146512_(_088777_, _091418_, _091423_);
  and g_146513_(_088780_, _091423_, _091424_);
  not g_146514_(_091424_, _091426_);
  and g_146515_(_091421_, _091426_, _091427_);
  or g_146516_(_091420_, _091424_, _091428_);
  and g_146517_(_088783_, _088791_, _091429_);
  xor g_146518_(_091428_, _091429_, _091430_);
  and g_146519_(_089768_, _091430_, _091431_);
  xor g_146520_(_089769_, _091430_, _091432_);
  and g_146521_(_088796_, _091432_, _091433_);
  or g_146522_(_088796_, _091432_, _091434_);
  xor g_146523_(_088795_, _091432_, _091435_);
  and g_146524_(_088803_, _088805_, _091437_);
  xor g_146525_(_091435_, _091437_, _091438_);
  not g_146526_(_091438_, _091439_);
  or g_146527_(_089767_, _091439_, _091440_);
  xor g_146528_(_089767_, _091438_, _091441_);
  and g_146529_(_088812_, _091441_, _091442_);
  or g_146530_(_088812_, _091441_, _091443_);
  xor g_146531_(_088812_, _091441_, _091444_);
  xor g_146532_(_088815_, _091444_, _091445_);
  or g_146533_(_086020_, _088820_, _091446_);
  not g_146534_(_091446_, _091448_);
  or g_146535_(_088818_, _091448_, _091449_);
  and g_146536_(_091445_, _091449_, _091450_);
  xor g_146537_(_091445_, _091449_, _091451_);
  or g_146538_(_086023_, _088821_, _091452_);
  and g_146539_(_088826_, _091452_, _091453_);
  not g_146540_(_091453_, _091454_);
  and g_146541_(_091451_, _091454_, _091455_);
  xor g_146542_(_091451_, _091453_, _091456_);
  and g_146543_(_088829_, _088832_, _091457_);
  or g_146544_(_091456_, _091457_, _091459_);
  xor g_146545_(_091456_, _091457_, _091460_);
  and g_146546_(_088834_, _091460_, _091461_);
  or g_146547_(_088834_, _091460_, _091462_);
  xor g_146548_(_088834_, _091460_, _091463_);
  and g_146549_(_086035_, _088837_, _091464_);
  or g_146550_(_088836_, _091464_, _091465_);
  not g_146551_(_091465_, _091466_);
  xor g_146552_(_091463_, _091466_, _091467_);
  or g_146553_(_089766_, _091467_, _091468_);
  xor g_146554_(_089766_, _091467_, _091470_);
  not g_146555_(_091470_, _091471_);
  or g_146556_(_089765_, _091471_, _091472_);
  xor g_146557_(_089765_, _091470_, _091473_);
  or g_146558_(_086046_, _088849_, _091474_);
  and g_146559_(_088847_, _091474_, _091475_);
  xor g_146560_(_091473_, _091475_, _091476_);
  and g_146561_(_089763_, _091476_, _091477_);
  xor g_146562_(_089763_, _091476_, _091478_);
  or g_146563_(_086053_, _088851_, _091479_);
  not g_146564_(_091479_, _091481_);
  and g_146565_(_091478_, _091481_, _091482_);
  xor g_146566_(_091478_, _091479_, _091483_);
  and g_146567_(_089762_, _091483_, _091484_);
  or g_146568_(_089762_, _091483_, _091485_);
  xor g_146569_(_089762_, _091483_, _091486_);
  xor g_146570_(_088856_, _091486_, _091487_);
  xor g_146571_(_088858_, _091487_, _091488_);
  xor g_146572_(_089760_, _091488_, _091489_);
  xor g_146573_(_089761_, _091488_, _091490_);
  or g_146574_(_089759_, _091490_, _091492_);
  xor g_146575_(_089759_, _091489_, _091493_);
  and g_146576_(_088877_, _091493_, _091494_);
  xor g_146577_(_088867_, _091490_, _091495_);
  xor g_146578_(_088867_, _091489_, _091496_);
  and g_146579_(_088876_, _091495_, _091497_);
  or g_146580_(_088877_, _091496_, _091498_);
  or g_146581_(_091494_, _091497_, _091499_);
  or g_146582_(_086082_, _088881_, _091500_);
  and g_146583_(_088879_, _091500_, _091501_);
  xor g_146584_(_091499_, _091501_, _091503_);
  or g_146585_(_089758_, _091503_, _091504_);
  and g_146586_(_089758_, _091503_, _091505_);
  xor g_146587_(_089758_, _091503_, _091506_);
  xor g_146588_(_088892_, _091506_, _091507_);
  not g_146589_(_091507_, _091508_);
  or g_146590_(_088899_, _091508_, _091509_);
  or g_146591_(_088884_, _091507_, _091510_);
  xor g_146592_(_088886_, _091507_, _091511_);
  or g_146593_(_088898_, _091511_, _091512_);
  and g_146594_(_091509_, _091512_, _091514_);
  not g_146595_(_091514_, _091515_);
  or g_146596_(_088904_, _091514_, _091516_);
  not g_146597_(_091516_, _091517_);
  or g_146598_(_088901_, _091515_, _091518_);
  or g_146599_(_088902_, _091514_, _091519_);
  and g_146600_(_088904_, _091519_, _091520_);
  and g_146601_(_091518_, _091520_, _091521_);
  or g_146602_(_091517_, _091521_, _091522_);
  not g_146603_(_091522_, _091523_);
  or g_146604_(_089756_, _091522_, _091525_);
  and g_146605_(_088906_, _091523_, _091526_);
  or g_146606_(_088908_, _091522_, _091527_);
  and g_146607_(_088908_, _091522_, _091528_);
  or g_146608_(_088906_, _091523_, _091529_);
  and g_146609_(_089756_, _091529_, _091530_);
  or g_146610_(_089757_, _091528_, _091531_);
  and g_146611_(_091527_, _091530_, _091532_);
  or g_146612_(_091526_, _091531_, _091533_);
  and g_146613_(_091525_, _091533_, _091534_);
  xor g_146614_(_089755_, _091534_, _091536_);
  or g_146615_(_088914_, _091536_, _091537_);
  xor g_146616_(_088915_, _091536_, _091538_);
  or g_146617_(_088919_, _091538_, _091539_);
  xor g_146618_(_088917_, _091538_, _091540_);
  and g_146619_(_088922_, _091540_, _091541_);
  or g_146620_(_088922_, _091538_, _091542_);
  not g_146621_(_091542_, _091543_);
  or g_146622_(_091541_, _091543_, _091544_);
  not g_146623_(_091544_, _091545_);
  xor g_146624_(_088925_, _091544_, _091547_);
  or g_146625_(_088928_, _091547_, _091548_);
  and g_146626_(_088928_, _091545_, _091549_);
  or g_146627_(_088927_, _091544_, _091550_);
  and g_146628_(_091548_, _091550_, _091551_);
  xor g_146629_(_088933_, _091551_, _091552_);
  xor g_146630_(_088932_, _091551_, _091553_);
  and g_146631_(_088936_, _091553_, _091554_);
  or g_146632_(_088935_, _091552_, _091555_);
  and g_146633_(_088935_, _091551_, _091556_);
  or g_146634_(_091554_, _091556_, _091558_);
  or g_146635_(_088943_, _091558_, _091559_);
  not g_146636_(_091559_, _091560_);
  xor g_146637_(_088938_, _091558_, _091561_);
  xor g_146638_(_088939_, _091558_, _091562_);
  and g_146639_(_088943_, _091562_, _091563_);
  or g_146640_(_088944_, _091561_, _091564_);
  and g_146641_(_091559_, _091564_, _091565_);
  or g_146642_(_091560_, _091563_, _091566_);
  or g_146643_(_088949_, _091566_, _091567_);
  not g_146644_(_091567_, _091569_);
  xor g_146645_(_088947_, _091565_, _091570_);
  xor g_146646_(_088947_, _091566_, _091571_);
  and g_146647_(_088949_, _091570_, _091572_);
  or g_146648_(_088950_, _091571_, _091573_);
  and g_146649_(_088953_, _091573_, _091574_);
  or g_146650_(_088954_, _091572_, _091575_);
  and g_146651_(_091567_, _091575_, _091576_);
  or g_146652_(_091569_, _091574_, _091577_);
  or g_146653_(_088953_, _091573_, _091578_);
  and g_146654_(_091576_, _091578_, _091580_);
  and g_146655_(_089752_, _091580_, _091581_);
  or g_146656_(_089752_, _091580_, _091582_);
  xor g_146657_(_089754_, _091580_, _091583_);
  xor g_146658_(_089751_, _091583_, _091584_);
  or g_146659_(_088965_, _091584_, _091585_);
  xor g_146660_(_088965_, _091584_, _091586_);
  and g_146661_(_088967_, _091586_, _091587_);
  xor g_146662_(_088967_, _091586_, _091588_);
  xor g_146663_(_088968_, _091586_, _091589_);
  and g_146664_(_089750_, _091589_, _091591_);
  or g_146665_(_089749_, _091588_, _091592_);
  and g_146666_(_089748_, _091591_, _091593_);
  and g_146667_(_089749_, _091586_, _091594_);
  or g_146668_(_089747_, _091594_, _091595_);
  and g_146669_(_091592_, _091595_, _091596_);
  or g_146670_(_091593_, _091596_, _091597_);
  or g_146671_(_088977_, _091597_, _091598_);
  xor g_146672_(_088978_, _091597_, _091599_);
  not g_146673_(_091599_, _091600_);
  or g_146674_(_088980_, _091599_, _091602_);
  xor g_146675_(_088981_, _091599_, _091603_);
  or g_146676_(_088986_, _091603_, _091604_);
  or g_146677_(_088985_, _091600_, _091605_);
  and g_146678_(_091604_, _091605_, _091606_);
  xor g_146679_(_088988_, _091606_, _091607_);
  xor g_146680_(_088989_, _091606_, _091608_);
  and g_146681_(_088996_, _091608_, _091609_);
  or g_146682_(_088997_, _091607_, _091610_);
  or g_146683_(_088996_, _091606_, _091611_);
  and g_146684_(_091610_, _091611_, _091613_);
  or g_146685_(_086175_, _088999_, _091614_);
  and g_146686_(_088993_, _091614_, _091615_);
  xor g_146687_(_091613_, _091615_, _091616_);
  not g_146688_(_091616_, _091617_);
  and g_146689_(_089746_, _091617_, _091618_);
  xor g_146690_(_089746_, _091616_, _091619_);
  and g_146691_(_089744_, _091619_, _091620_);
  or g_146692_(_089744_, _091619_, _091621_);
  xor g_146693_(_089745_, _091619_, _091622_);
  xor g_146694_(_089009_, _091622_, _091624_);
  and g_146695_(_089013_, _091624_, _091625_);
  or g_146696_(_089013_, _091622_, _091626_);
  not g_146697_(_091626_, _091627_);
  or g_146698_(_091625_, _091627_, _091628_);
  or g_146699_(_086197_, _089014_, _091629_);
  and g_146700_(_089016_, _091629_, _091630_);
  not g_146701_(_091630_, _091631_);
  xor g_146702_(_091628_, _091631_, _091632_);
  or g_146703_(_089743_, _091632_, _091633_);
  and g_146704_(_089743_, _091632_, _091635_);
  xor g_146705_(_089743_, _091632_, _091636_);
  xor g_146706_(_089741_, _091636_, _091637_);
  or g_146707_(_089740_, _091637_, _091638_);
  xor g_146708_(_089739_, _091637_, _091639_);
  and g_146709_(_089025_, _089029_, _091640_);
  or g_146710_(_089024_, _091640_, _091641_);
  or g_146711_(_091639_, _091641_, _091642_);
  xor g_146712_(_091639_, _091641_, _091643_);
  not g_146713_(_091643_, _091644_);
  and g_146714_(_089035_, _091643_, _091646_);
  or g_146715_(_089034_, _091644_, _091647_);
  or g_146716_(_089027_, _089030_, _091648_);
  or g_146717_(_091644_, _091648_, _091649_);
  xor g_146718_(_091643_, _091648_, _091650_);
  and g_146719_(_089034_, _091650_, _091651_);
  or g_146720_(_091646_, _091651_, _091652_);
  and g_146721_(_089037_, _089044_, _091653_);
  xor g_146722_(_091652_, _091653_, _091654_);
  or g_146723_(_089737_, _091654_, _091655_);
  and g_146724_(_089737_, _091654_, _091657_);
  xor g_146725_(_089738_, _091654_, _091658_);
  xor g_146726_(_089734_, _091658_, _091659_);
  or g_146727_(_089059_, _091659_, _091660_);
  and g_146728_(_089059_, _091659_, _091661_);
  xor g_146729_(_089059_, _091659_, _091662_);
  xor g_146730_(_089062_, _091662_, _091663_);
  or g_146731_(_089730_, _091663_, _091664_);
  and g_146732_(_089730_, _091663_, _091665_);
  not g_146733_(_091665_, _091666_);
  xor g_146734_(_089729_, _091663_, _091668_);
  and g_146735_(_089727_, _091668_, _091669_);
  not g_146736_(_091669_, _091670_);
  and g_146737_(_089728_, _091664_, _091671_);
  not g_146738_(_091671_, _091672_);
  and g_146739_(_091666_, _091671_, _091673_);
  or g_146740_(_091665_, _091672_, _091674_);
  and g_146741_(_091670_, _091674_, _091675_);
  or g_146742_(_091669_, _091673_, _091676_);
  and g_146743_(_089070_, _091675_, _091677_);
  or g_146744_(_089071_, _091676_, _091679_);
  or g_146745_(_089070_, _091668_, _091680_);
  and g_146746_(_091679_, _091680_, _091681_);
  xor g_146747_(_089725_, _091681_, _091682_);
  and g_146748_(_089724_, _091682_, _091683_);
  xor g_146749_(_089723_, _091682_, _091684_);
  and g_146750_(_089080_, _091684_, _091685_);
  or g_146751_(_089080_, _091684_, _091686_);
  xor g_146752_(_089080_, _091684_, _091687_);
  xor g_146753_(_089084_, _091687_, _091688_);
  or g_146754_(_089087_, _091688_, _091690_);
  xor g_146755_(_089088_, _091688_, _091691_);
  or g_146756_(_089090_, _091691_, _091692_);
  and g_146757_(_089090_, _091691_, _091693_);
  xor g_146758_(_089090_, _091691_, _091694_);
  and g_146759_(_089092_, _091694_, _091695_);
  not g_146760_(_091695_, _091696_);
  or g_146761_(_089092_, _091694_, _091697_);
  or g_146762_(_086262_, _089093_, _091698_);
  not g_146763_(_091698_, _091699_);
  and g_146764_(_091697_, _091698_, _091701_);
  not g_146765_(_091701_, _091702_);
  and g_146766_(_091696_, _091701_, _091703_);
  or g_146767_(_091695_, _091702_, _091704_);
  and g_146768_(_091694_, _091699_, _091705_);
  or g_146769_(_091703_, _091705_, _091706_);
  xor g_146770_(_089721_, _091706_, _091707_);
  and g_146771_(_089719_, _091707_, _091708_);
  or g_146772_(_089719_, _091707_, _091709_);
  xor g_146773_(_089719_, _091707_, _091710_);
  xor g_146774_(_089718_, _091710_, _091712_);
  and g_146775_(_089100_, _091712_, _091713_);
  or g_146776_(_089100_, _091712_, _091714_);
  xor g_146777_(_089101_, _091712_, _091715_);
  xor g_146778_(_089104_, _091715_, _091716_);
  or g_146779_(_089108_, _089111_, _091717_);
  and g_146780_(_091716_, _091717_, _091718_);
  xor g_146781_(_091716_, _091717_, _091719_);
  and g_146782_(_089115_, _091719_, _091720_);
  xor g_146783_(_089114_, _091719_, _091721_);
  and g_146784_(_089119_, _089122_, _091723_);
  not g_146785_(_091723_, _091724_);
  xor g_146786_(_091721_, _091724_, _091725_);
  or g_146787_(_089125_, _091725_, _091726_);
  and g_146788_(_089125_, _091725_, _091727_);
  xor g_146789_(_089125_, _091725_, _091728_);
  xor g_146790_(_089126_, _091725_, _091729_);
  and g_146791_(_089129_, _091728_, _091730_);
  not g_146792_(_091730_, _091731_);
  and g_146793_(_089130_, _091729_, _091732_);
  or g_146794_(_089129_, _091728_, _091734_);
  or g_146795_(_086293_, _089131_, _091735_);
  not g_146796_(_091735_, _091736_);
  and g_146797_(_091734_, _091735_, _091737_);
  or g_146798_(_091732_, _091736_, _091738_);
  and g_146799_(_091731_, _091737_, _091739_);
  or g_146800_(_091730_, _091738_, _091740_);
  and g_146801_(_089717_, _091739_, _091741_);
  or g_146802_(_091729_, _091735_, _091742_);
  and g_146803_(_089717_, _091742_, _091743_);
  not g_146804_(_091743_, _091745_);
  and g_146805_(_091740_, _091745_, _091746_);
  or g_146806_(_091739_, _091743_, _091747_);
  or g_146807_(_091741_, _091746_, _091748_);
  or g_146808_(_089715_, _091748_, _091749_);
  xor g_146809_(_089716_, _091748_, _091750_);
  and g_146810_(_089140_, _091750_, _091751_);
  or g_146811_(_089140_, _091750_, _091752_);
  xor g_146812_(_089140_, _091750_, _091753_);
  not g_146813_(_091753_, _091754_);
  or g_146814_(_089145_, _091754_, _091756_);
  not g_146815_(_091756_, _091757_);
  and g_146816_(_089143_, _091753_, _091758_);
  not g_146817_(_091758_, _091759_);
  or g_146818_(_089143_, _091753_, _091760_);
  and g_146819_(_089145_, _091760_, _091761_);
  and g_146820_(_091759_, _091761_, _091762_);
  or g_146821_(_091757_, _091762_, _091763_);
  xor g_146822_(_089714_, _091763_, _091764_);
  or g_146823_(_089712_, _091764_, _091765_);
  and g_146824_(_089712_, _091764_, _091767_);
  xor g_146825_(_089712_, _091764_, _091768_);
  and g_146826_(_089152_, _089156_, _091769_);
  xor g_146827_(_091768_, _091769_, _091770_);
  or g_146828_(_089711_, _091770_, _091771_);
  and g_146829_(_089711_, _091770_, _091772_);
  xor g_146830_(_089711_, _091770_, _091773_);
  xor g_146831_(_089710_, _091773_, _091774_);
  and g_146832_(_089164_, _091774_, _091775_);
  or g_146833_(_089164_, _091774_, _091776_);
  xor g_146834_(_089164_, _091774_, _091778_);
  not g_146835_(_091778_, _091779_);
  xor g_146836_(_089170_, _091778_, _091780_);
  and g_146837_(_089174_, _091780_, _091781_);
  not g_146838_(_091781_, _091782_);
  and g_146839_(_089175_, _091778_, _091783_);
  or g_146840_(_089174_, _091779_, _091784_);
  and g_146841_(_091782_, _091784_, _091785_);
  or g_146842_(_091781_, _091783_, _091786_);
  and g_146843_(_086336_, _089178_, _091787_);
  or g_146844_(_086335_, _089179_, _091789_);
  and g_146845_(_089177_, _091789_, _091790_);
  xor g_146846_(_091786_, _091790_, _091791_);
  and g_146847_(_089707_, _091791_, _091792_);
  xor g_146848_(_089708_, _091791_, _091793_);
  or g_146849_(_089705_, _091793_, _091794_);
  and g_146850_(_089705_, _091793_, _091795_);
  xor g_146851_(_089706_, _091793_, _091796_);
  xor g_146852_(_089704_, _091796_, _091797_);
  and g_146853_(_089189_, _091797_, _091798_);
  or g_146854_(_089189_, _091797_, _091800_);
  xor g_146855_(_089190_, _091797_, _091801_);
  or g_146856_(_086350_, _089196_, _091802_);
  and g_146857_(_089195_, _091802_, _091803_);
  not g_146858_(_091803_, _091804_);
  xor g_146859_(_091801_, _091804_, _091805_);
  and g_146860_(_089703_, _091805_, _091806_);
  or g_146861_(_089703_, _091805_, _091807_);
  xor g_146862_(_089703_, _091805_, _091808_);
  xor g_146863_(_089702_, _091808_, _091809_);
  or g_146864_(_089701_, _091809_, _091811_);
  or g_146865_(_089205_, _091809_, _091812_);
  xor g_146866_(_089206_, _091809_, _091813_);
  and g_146867_(_089701_, _091813_, _091814_);
  or g_146868_(_089208_, _089209_, _091815_);
  or g_146869_(_091814_, _091815_, _091816_);
  and g_146870_(_091811_, _091816_, _091817_);
  not g_146871_(_091817_, _091818_);
  and g_146872_(_091814_, _091815_, _091819_);
  not g_146873_(_091819_, _091820_);
  and g_146874_(_091817_, _091820_, _091822_);
  or g_146875_(_091818_, _091819_, _091823_);
  or g_146876_(_089212_, _091823_, _091824_);
  xor g_146877_(_089212_, _091822_, _091825_);
  and g_146878_(_089216_, _089219_, _091826_);
  or g_146879_(_091825_, _091826_, _091827_);
  xor g_146880_(_091825_, _091826_, _091828_);
  and g_146881_(_089222_, _091828_, _091829_);
  xor g_146882_(_089222_, _091828_, _091830_);
  and g_146883_(_089699_, _091830_, _091831_);
  or g_146884_(_089699_, _091830_, _091833_);
  xor g_146885_(_089700_, _091830_, _091834_);
  xor g_146886_(_089697_, _091834_, _091835_);
  not g_146887_(_091835_, _091836_);
  and g_146888_(_089696_, _091836_, _091837_);
  xor g_146889_(_089696_, _091835_, _091838_);
  or g_146890_(_089695_, _091838_, _091839_);
  and g_146891_(_089695_, _091838_, _091840_);
  xor g_146892_(_089695_, _091838_, _091841_);
  xor g_146893_(_089233_, _091841_, _091842_);
  not g_146894_(_091842_, _091844_);
  or g_146895_(_089240_, _091842_, _091845_);
  not g_146896_(_091845_, _091846_);
  and g_146897_(_089235_, _091844_, _091847_);
  xor g_146898_(_089236_, _091842_, _091848_);
  xor g_146899_(_089235_, _091842_, _091849_);
  and g_146900_(_089240_, _091849_, _091850_);
  or g_146901_(_089241_, _091848_, _091851_);
  and g_146902_(_091845_, _091851_, _091852_);
  or g_146903_(_086397_, _089242_, _091853_);
  not g_146904_(_091853_, _091855_);
  or g_146905_(_091852_, _091855_, _091856_);
  or g_146906_(_091850_, _091853_, _091857_);
  or g_146907_(_091846_, _091857_, _091858_);
  and g_146908_(_091856_, _091858_, _091859_);
  and g_146909_(_089694_, _091859_, _091860_);
  xor g_146910_(_089694_, _091859_, _091861_);
  and g_146911_(_089247_, _091861_, _091862_);
  xor g_146912_(_089249_, _091861_, _091863_);
  or g_146913_(_089691_, _091863_, _091864_);
  xor g_146914_(_089692_, _091863_, _091866_);
  or g_146915_(_089690_, _091866_, _091867_);
  xor g_146916_(_089690_, _091866_, _091868_);
  and g_146917_(_089253_, _091868_, _091869_);
  xor g_146918_(_089253_, _091868_, _091870_);
  or g_146919_(_089255_, _091870_, _091871_);
  and g_146920_(_089255_, _091868_, _091872_);
  not g_146921_(_091872_, _091873_);
  and g_146922_(_091871_, _091873_, _091874_);
  xor g_146923_(_089689_, _091874_, _091875_);
  and g_146924_(_089688_, _091875_, _091877_);
  xor g_146925_(_089686_, _091875_, _091878_);
  or g_146926_(_089265_, _091878_, _091879_);
  and g_146927_(_089265_, _091878_, _091880_);
  xor g_146928_(_089265_, _091878_, _091881_);
  xor g_146929_(_089268_, _091881_, _091882_);
  xor g_146930_(_089683_, _091882_, _091883_);
  xor g_146931_(_089684_, _091882_, _091884_);
  and g_146932_(_089275_, _091883_, _091885_);
  or g_146933_(_089276_, _091884_, _091886_);
  or g_146934_(_089273_, _091882_, _091888_);
  xor g_146935_(_089273_, _091882_, _091889_);
  or g_146936_(_089275_, _091889_, _091890_);
  and g_146937_(_091886_, _091890_, _091891_);
  and g_146938_(_089279_, _089283_, _091892_);
  not g_146939_(_091892_, _091893_);
  and g_146940_(_091891_, _091893_, _091894_);
  xor g_146941_(_091891_, _091892_, _091895_);
  or g_146942_(_089286_, _091895_, _091896_);
  xor g_146943_(_089287_, _091895_, _091897_);
  or g_146944_(_089290_, _091897_, _091899_);
  and g_146945_(_089290_, _091897_, _091900_);
  xor g_146946_(_089291_, _091897_, _091901_);
  xor g_146947_(_089295_, _091901_, _091902_);
  and g_146948_(_089297_, _091902_, _091903_);
  or g_146949_(_089297_, _091901_, _091904_);
  not g_146950_(_091904_, _091905_);
  or g_146951_(_091903_, _091905_, _091906_);
  not g_146952_(_091906_, _091907_);
  or g_146953_(_089304_, _091906_, _091908_);
  xor g_146954_(_089300_, _091906_, _091910_);
  xor g_146955_(_089300_, _091907_, _091911_);
  and g_146956_(_089304_, _091911_, _091912_);
  or g_146957_(_089305_, _091910_, _091913_);
  and g_146958_(_091908_, _091913_, _091914_);
  xor g_146959_(_089310_, _091914_, _091915_);
  or g_146960_(_089309_, _091915_, _091916_);
  and g_146961_(_089309_, _091915_, _091917_);
  xor g_146962_(_089309_, _091915_, _091918_);
  xor g_146963_(_089316_, _091918_, _091919_);
  and g_146964_(_089682_, _091919_, _091921_);
  xor g_146965_(_089681_, _091919_, _091922_);
  or g_146966_(_089679_, _091922_, _091923_);
  xor g_146967_(_089680_, _091922_, _091924_);
  or g_146968_(_089323_, _091924_, _091925_);
  xor g_146969_(_089324_, _091924_, _091926_);
  and g_146970_(_089328_, _089331_, _091927_);
  or g_146971_(_091926_, _091927_, _091928_);
  xor g_146972_(_091926_, _091927_, _091929_);
  not g_146973_(_091929_, _091930_);
  and g_146974_(_089337_, _091929_, _091932_);
  or g_146975_(_089338_, _091930_, _091933_);
  or g_146976_(_089333_, _091930_, _091934_);
  xor g_146977_(_089333_, _091929_, _091935_);
  and g_146978_(_089338_, _091935_, _091936_);
  or g_146979_(_091932_, _091936_, _091937_);
  not g_146980_(_091937_, _091938_);
  xor g_146981_(_089340_, _091937_, _091939_);
  xor g_146982_(_089341_, _091937_, _091940_);
  and g_146983_(_089346_, _091940_, _091941_);
  or g_146984_(_089345_, _091939_, _091943_);
  and g_146985_(_089345_, _091938_, _091944_);
  or g_146986_(_089346_, _091937_, _091945_);
  and g_146987_(_091943_, _091945_, _091946_);
  or g_146988_(_091941_, _091944_, _091947_);
  and g_146989_(_089354_, _091946_, _091948_);
  or g_146990_(_089353_, _091947_, _091949_);
  or g_146991_(_089351_, _091943_, _091950_);
  or g_146992_(_089350_, _091940_, _091951_);
  and g_146993_(_091945_, _091951_, _091952_);
  and g_146994_(_091950_, _091952_, _091954_);
  or g_146995_(_089354_, _091954_, _091955_);
  and g_146996_(_091949_, _091955_, _091956_);
  or g_146997_(_086492_, _089361_, _091957_);
  not g_146998_(_091957_, _091958_);
  and g_146999_(_089359_, _091957_, _091959_);
  not g_147000_(_091959_, _091960_);
  xor g_147001_(_091956_, _091960_, _091961_);
  or g_147002_(_089678_, _091961_, _091962_);
  and g_147003_(_089678_, _091961_, _091963_);
  xor g_147004_(_089678_, _091961_, _091965_);
  xor g_147005_(_089367_, _091965_, _091966_);
  xor g_147006_(_089366_, _091965_, _091967_);
  and g_147007_(_089677_, _091967_, _091968_);
  or g_147008_(_089675_, _091966_, _091969_);
  and g_147009_(_089674_, _091968_, _091970_);
  and g_147010_(_089675_, _091965_, _091971_);
  or g_147011_(_089673_, _091971_, _091972_);
  and g_147012_(_091969_, _091972_, _091973_);
  or g_147013_(_091970_, _091973_, _091974_);
  not g_147014_(_091974_, _091976_);
  and g_147015_(_089373_, _091976_, _091977_);
  xor g_147016_(_089373_, _091974_, _091978_);
  not g_147017_(_091978_, _091979_);
  or g_147018_(_089379_, _091978_, _091980_);
  not g_147019_(_091980_, _091981_);
  and g_147020_(_089376_, _091979_, _091982_);
  xor g_147021_(_089376_, _091978_, _091983_);
  and g_147022_(_089379_, _091983_, _091984_);
  or g_147023_(_091981_, _091984_, _091985_);
  xor g_147024_(_089384_, _091985_, _091987_);
  not g_147025_(_091987_, _091988_);
  or g_147026_(_086524_, _089388_, _091989_);
  and g_147027_(_089387_, _091989_, _091990_);
  or g_147028_(_091987_, _091990_, _091991_);
  xor g_147029_(_091987_, _091990_, _091992_);
  xor g_147030_(_091988_, _091990_, _091993_);
  or g_147031_(_089672_, _091993_, _091994_);
  xor g_147032_(_089672_, _091992_, _091995_);
  or g_147033_(_089395_, _091995_, _091996_);
  xor g_147034_(_089395_, _091995_, _091998_);
  and g_147035_(_089397_, _091998_, _091999_);
  or g_147036_(_089397_, _091998_, _092000_);
  xor g_147037_(_089397_, _091998_, _092001_);
  xor g_147038_(_089401_, _092001_, _092002_);
  or g_147039_(_089404_, _092002_, _092003_);
  and g_147040_(_089404_, _092002_, _092004_);
  xor g_147041_(_089404_, _092002_, _092005_);
  xor g_147042_(_089405_, _092002_, _092006_);
  or g_147043_(_089411_, _092006_, _092007_);
  not g_147044_(_092007_, _092009_);
  xor g_147045_(_089409_, _092005_, _092010_);
  and g_147046_(_089411_, _092010_, _092011_);
  or g_147047_(_092009_, _092011_, _092012_);
  not g_147048_(_092012_, _092013_);
  or g_147049_(_089418_, _092012_, _092014_);
  and g_147050_(_089414_, _092013_, _092015_);
  or g_147051_(_089415_, _092012_, _092016_);
  and g_147052_(_089415_, _092012_, _092017_);
  or g_147053_(_089414_, _092013_, _092018_);
  and g_147054_(_089418_, _092018_, _092020_);
  or g_147055_(_089419_, _092017_, _092021_);
  and g_147056_(_092016_, _092020_, _092022_);
  or g_147057_(_092015_, _092021_, _092023_);
  and g_147058_(_092014_, _092023_, _092024_);
  not g_147059_(_092024_, _092025_);
  or g_147060_(_086545_, _089422_, _092026_);
  not g_147061_(_092026_, _092027_);
  and g_147062_(_092024_, _092027_, _092028_);
  or g_147063_(_092025_, _092026_, _092029_);
  xor g_147064_(_089421_, _092024_, _092031_);
  and g_147065_(_092026_, _092031_, _092032_);
  or g_147066_(_092028_, _092032_, _092033_);
  xor g_147067_(_089671_, _092033_, _092034_);
  and g_147068_(_089432_, _092034_, _092035_);
  xor g_147069_(_089431_, _092034_, _092036_);
  and g_147070_(_089430_, _092036_, _092037_);
  or g_147071_(_089430_, _092036_, _092038_);
  xor g_147072_(_089430_, _092036_, _092039_);
  and g_147073_(_089438_, _089440_, _092040_);
  xor g_147074_(_092039_, _092040_, _092042_);
  or g_147075_(_089443_, _092042_, _092043_);
  and g_147076_(_089443_, _092042_, _092044_);
  xor g_147077_(_089443_, _092042_, _092045_);
  xor g_147078_(_089447_, _092045_, _092046_);
  or g_147079_(_089449_, _092046_, _092047_);
  and g_147080_(_089449_, _092046_, _092048_);
  xor g_147081_(_089449_, _092046_, _092049_);
  xor g_147082_(_089670_, _092049_, _092050_);
  or g_147083_(_089669_, _092050_, _092051_);
  and g_147084_(_089669_, _092050_, _092053_);
  xor g_147085_(_089669_, _092050_, _092054_);
  xor g_147086_(_089455_, _092054_, _092055_);
  and g_147087_(_089461_, _092055_, _092056_);
  xor g_147088_(_089461_, _092055_, _092057_);
  not g_147089_(_092057_, _092058_);
  and g_147090_(_089464_, _092057_, _092059_);
  xor g_147091_(_089465_, _092057_, _092060_);
  not g_147092_(_092060_, _092061_);
  or g_147093_(_089475_, _092060_, _092062_);
  xor g_147094_(_089475_, _092060_, _092064_);
  xor g_147095_(_089475_, _092061_, _092065_);
  and g_147096_(_089473_, _092065_, _092066_);
  or g_147097_(_089474_, _092064_, _092067_);
  or g_147098_(_089473_, _092058_, _092068_);
  not g_147099_(_092068_, _092069_);
  and g_147100_(_092067_, _092068_, _092070_);
  or g_147101_(_092066_, _092069_, _092071_);
  and g_147102_(_089481_, _089483_, _092072_);
  xor g_147103_(_092070_, _092072_, _092073_);
  and g_147104_(_086594_, _089486_, _092075_);
  or g_147105_(_089485_, _092075_, _092076_);
  or g_147106_(_092073_, _092076_, _092077_);
  xor g_147107_(_092073_, _092076_, _092078_);
  and g_147108_(_089668_, _092078_, _092079_);
  xor g_147109_(_089668_, _092078_, _092080_);
  xor g_147110_(_089667_, _092078_, _092081_);
  or g_147111_(_089492_, _092080_, _092082_);
  and g_147112_(_089492_, _092080_, _092083_);
  xor g_147113_(_089492_, _092081_, _092084_);
  and g_147114_(_089496_, _089499_, _092086_);
  xor g_147115_(_092084_, _092086_, _092087_);
  or g_147116_(_089664_, _092087_, _092088_);
  and g_147117_(_089664_, _092087_, _092089_);
  xor g_147118_(_089666_, _092087_, _092090_);
  xor g_147119_(_089661_, _092090_, _092091_);
  or g_147120_(_089658_, _092091_, _092092_);
  xor g_147121_(_089659_, _092091_, _092093_);
  or g_147122_(_089657_, _092093_, _092094_);
  xor g_147123_(_089656_, _092093_, _092095_);
  or g_147124_(_089505_, _092095_, _092097_);
  and g_147125_(_089505_, _092095_, _092098_);
  xor g_147126_(_089505_, _092095_, _092099_);
  xor g_147127_(_089508_, _092099_, _092100_);
  or g_147128_(_089655_, _092100_, _092101_);
  xor g_147129_(_089655_, _092100_, _092102_);
  and g_147130_(_089652_, _092102_, _092103_);
  or g_147131_(_089652_, _092102_, _092104_);
  xor g_147132_(_089653_, _092102_, _092105_);
  or g_147133_(_089650_, _092105_, _092106_);
  and g_147134_(_086635_, _089516_, _092108_);
  not g_147135_(_092108_, _092109_);
  xor g_147136_(_092105_, _092109_, _092110_);
  xor g_147137_(_092105_, _092108_, _092111_);
  and g_147138_(_089650_, _092111_, _092112_);
  or g_147139_(_089651_, _092110_, _092113_);
  and g_147140_(_092106_, _092113_, _092114_);
  xor g_147141_(_089649_, _092114_, _092115_);
  and g_147142_(_089648_, _092115_, _092116_);
  or g_147143_(_089648_, _092115_, _092117_);
  xor g_147144_(_089648_, _092115_, _092119_);
  xor g_147145_(_089647_, _092119_, _092120_);
  or g_147146_(_089644_, _092120_, _092121_);
  and g_147147_(_089644_, _092120_, _092122_);
  xor g_147148_(_089644_, _092120_, _092123_);
  xor g_147149_(_089642_, _092123_, _092124_);
  or g_147150_(_089638_, _092124_, _092125_);
  and g_147151_(_089638_, _092124_, _092126_);
  xor g_147152_(_089638_, _092124_, _092127_);
  xor g_147153_(_089637_, _092127_, _092128_);
  or g_147154_(_089528_, _092128_, _092130_);
  xor g_147155_(_089528_, _092128_, _092131_);
  and g_147156_(_089535_, _092131_, _092132_);
  xor g_147157_(_089535_, _092131_, _092133_);
  and g_147158_(_089530_, _092133_, _092134_);
  xor g_147159_(_089530_, _092133_, _092135_);
  and g_147160_(_089538_, _092135_, _092136_);
  xor g_147161_(_089538_, _092135_, _092137_);
  and g_147162_(_089543_, _092137_, _092138_);
  xor g_147163_(_089542_, _092137_, _092139_);
  or g_147164_(_089635_, _092139_, _092141_);
  xor g_147165_(_089636_, _092139_, _092142_);
  not g_147166_(_092142_, _092143_);
  and g_147167_(_089548_, _092143_, _092144_);
  xor g_147168_(_089549_, _092142_, _092145_);
  and g_147169_(_089554_, _092145_, _092146_);
  not g_147170_(_092146_, _092147_);
  and g_147171_(_089551_, _092145_, _092148_);
  xor g_147172_(_089551_, _092145_, _092149_);
  or g_147173_(_089554_, _092149_, _092150_);
  and g_147174_(_092147_, _092150_, _092152_);
  xor g_147175_(_089634_, _092152_, _092153_);
  and g_147176_(_089633_, _092153_, _092154_);
  xor g_147177_(_089633_, _092153_, _092155_);
  and g_147178_(_089628_, _092155_, _092156_);
  xor g_147179_(_089629_, _092155_, _092157_);
  or g_147180_(_089626_, _092157_, _092158_);
  xor g_147181_(_089627_, _092157_, _092159_);
  and g_147182_(_089566_, _089569_, _092160_);
  not g_147183_(_092160_, _092161_);
  or g_147184_(_092159_, _092160_, _092163_);
  xor g_147185_(_092159_, _092161_, _092164_);
  and g_147186_(_089573_, _092164_, _092165_);
  or g_147187_(_089573_, _092164_, _092166_);
  xor g_147188_(_089574_, _092164_, _092167_);
  xor g_147189_(_089625_, _092167_, _092168_);
  xor g_147190_(_089624_, _092167_, _092169_);
  or g_147191_(_089623_, _092168_, _092170_);
  xor g_147192_(_089623_, _092169_, _092171_);
  and g_147193_(_086744_, _089584_, _092172_);
  or g_147194_(_089583_, _092172_, _092174_);
  or g_147195_(_092171_, _092174_, _092175_);
  xor g_147196_(_092171_, _092174_, _092176_);
  and g_147197_(_086754_, _089585_, _092177_);
  or g_147198_(_089590_, _092177_, _092178_);
  not g_147199_(_092178_, _092179_);
  and g_147200_(_092176_, _092178_, _092180_);
  xor g_147201_(_092176_, _092178_, _092181_);
  xor g_147202_(_092176_, _092179_, _092182_);
  and g_147203_(_089596_, _089601_, _092183_);
  or g_147204_(_089595_, _089599_, _092185_);
  and g_147205_(_092182_, _092183_, _092186_);
  or g_147206_(_092181_, _092185_, _092187_);
  and g_147207_(_092181_, _092185_, _092188_);
  xor g_147208_(_092182_, _092183_, _092189_);
  not g_147209_(_092189_, _092190_);
  or g_147210_(_089620_, _092190_, _092191_);
  not g_147211_(_092191_, _092192_);
  or g_147212_(_089604_, _092188_, _092193_);
  or g_147213_(_092186_, _092193_, _092194_);
  or g_147214_(_089605_, _092189_, _092196_);
  and g_147215_(_089620_, _092196_, _092197_);
  and g_147216_(_092194_, _092197_, _092198_);
  not g_147217_(_092198_, _092199_);
  and g_147218_(_092191_, _092199_, _092200_);
  or g_147219_(_092192_, _092198_, _092201_);
  xor g_147220_(_089619_, _092201_, _092202_);
  xor g_147221_(_089619_, _092200_, _092203_);
  or g_147222_(_089618_, _092203_, _092204_);
  xor g_147223_(_089618_, _092202_, _092205_);
  and g_147224_(_089617_, _092205_, _092207_);
  or g_147225_(_089617_, _092205_, _092208_);
  xor g_147226_(_089617_, _092205_, _092209_);
  xor g_147227_(_089614_, _092209_, _092210_);
  or g_147228_(_089616_, _092210_, _092211_);
  xor g_147229_(_089616_, _092210_, out[966]);
  and g_147230_(_089614_, _092208_, _092212_);
  or g_147231_(_092207_, _092212_, _092213_);
  and g_147232_(_092187_, _092193_, _092214_);
  or g_147233_(_089624_, _092165_, _092215_);
  and g_147234_(_092166_, _092215_, _092217_);
  and g_147235_(_092158_, _092163_, _092218_);
  or g_147236_(_092154_, _092156_, _092219_);
  and g_147237_(_089634_, _092150_, _092220_);
  or g_147238_(_092146_, _092220_, _092221_);
  or g_147239_(_092144_, _092148_, _092222_);
  or g_147240_(_092136_, _092138_, _092223_);
  or g_147241_(_092132_, _092134_, _092224_);
  and g_147242_(_089637_, _092125_, _092225_);
  or g_147243_(_092126_, _092225_, _092226_);
  and g_147244_(_089641_, _092121_, _092228_);
  or g_147245_(_092122_, _092228_, _092229_);
  or g_147246_(_089646_, _092116_, _092230_);
  and g_147247_(_092117_, _092230_, _092231_);
  and g_147248_(_092092_, _092094_, _092232_);
  and g_147249_(_089661_, _092088_, _092233_);
  or g_147250_(_092089_, _092233_, _092234_);
  or g_147251_(_089499_, _092084_, _092235_);
  or g_147252_(_092056_, _092059_, _092236_);
  or g_147253_(_089454_, _092053_, _092237_);
  and g_147254_(_092051_, _092237_, _092239_);
  or g_147255_(_089670_, _092048_, _092240_);
  and g_147256_(_092047_, _092240_, _092241_);
  or g_147257_(_092037_, _092040_, _092242_);
  and g_147258_(_092038_, _092242_, _092243_);
  or g_147259_(_089671_, _092032_, _092244_);
  and g_147260_(_092029_, _092244_, _092245_);
  or g_147261_(_089421_, _092022_, _092246_);
  and g_147262_(_092014_, _092246_, _092247_);
  and g_147263_(_089414_, _092007_, _092248_);
  or g_147264_(_092011_, _092248_, _092250_);
  and g_147265_(_089409_, _092003_, _092251_);
  or g_147266_(_092004_, _092251_, _092252_);
  and g_147267_(_089400_, _092000_, _092253_);
  or g_147268_(_091999_, _092253_, _092254_);
  and g_147269_(_091994_, _091996_, _092255_);
  or g_147270_(_091977_, _091982_, _092256_);
  and g_147271_(_091956_, _091958_, _092257_);
  and g_147272_(_089357_, _091955_, _092258_);
  or g_147273_(_091948_, _092258_, _092259_);
  and g_147274_(_091925_, _091928_, _092261_);
  or g_147275_(_089315_, _091917_, _092262_);
  and g_147276_(_091916_, _092262_, _092263_);
  and g_147277_(_089310_, _091908_, _092264_);
  or g_147278_(_091912_, _092264_, _092265_);
  and g_147279_(_089300_, _091904_, _092266_);
  or g_147280_(_091903_, _092266_, _092267_);
  or g_147281_(_089294_, _091900_, _092268_);
  and g_147282_(_091899_, _092268_, _092269_);
  or g_147283_(_091885_, _091894_, _092270_);
  or g_147284_(_089689_, _091872_, _092272_);
  and g_147285_(_091871_, _092272_, _092273_);
  or g_147286_(_091860_, _091862_, _092274_);
  or g_147287_(_089233_, _091840_, _092275_);
  and g_147288_(_091839_, _092275_, _092276_);
  and g_147289_(_089697_, _091833_, _092277_);
  or g_147290_(_091831_, _092277_, _092278_);
  and g_147291_(_091824_, _091827_, _092279_);
  and g_147292_(_089702_, _091807_, _092280_);
  or g_147293_(_091806_, _092280_, _092281_);
  or g_147294_(_089199_, _091801_, _092283_);
  and g_147295_(_089194_, _091800_, _092284_);
  or g_147296_(_091798_, _092284_, _092285_);
  and g_147297_(_089704_, _091794_, _092286_);
  or g_147298_(_091795_, _092286_, _092287_);
  and g_147299_(_091785_, _091787_, _092288_);
  or g_147300_(_091792_, _092288_, _092289_);
  or g_147301_(_089177_, _091781_, _092290_);
  and g_147302_(_091784_, _092290_, _092291_);
  and g_147303_(_089710_, _091771_, _092292_);
  or g_147304_(_091772_, _092292_, _092294_);
  or g_147305_(_089170_, _091775_, _092295_);
  and g_147306_(_091776_, _092295_, _092296_);
  and g_147307_(_089155_, _091768_, _092297_);
  or g_147308_(_089713_, _091762_, _092298_);
  and g_147309_(_091756_, _092298_, _092299_);
  and g_147310_(_089129_, _091726_, _092300_);
  or g_147311_(_091727_, _092300_, _092301_);
  or g_147312_(_091721_, _091723_, _092302_);
  or g_147313_(_089104_, _091713_, _092303_);
  and g_147314_(_091714_, _092303_, _092305_);
  and g_147315_(_089721_, _091704_, _092306_);
  or g_147316_(_091705_, _092306_, _092307_);
  or g_147317_(_089084_, _091685_, _092308_);
  and g_147318_(_091686_, _092308_, _092309_);
  and g_147319_(_089726_, _091680_, _092310_);
  or g_147320_(_091677_, _092310_, _092311_);
  and g_147321_(_091666_, _091672_, _092312_);
  or g_147322_(_089062_, _091661_, _092313_);
  and g_147323_(_091660_, _092313_, _092314_);
  and g_147324_(_089734_, _091655_, _092316_);
  or g_147325_(_091657_, _092316_, _092317_);
  or g_147326_(_089047_, _091652_, _092318_);
  and g_147327_(_091638_, _091642_, _092319_);
  or g_147328_(_089741_, _091635_, _092320_);
  and g_147329_(_091633_, _092320_, _092321_);
  or g_147330_(_089008_, _091620_, _092322_);
  and g_147331_(_091621_, _092322_, _092323_);
  and g_147332_(_089002_, _091613_, _092324_);
  or g_147333_(_091618_, _092324_, _092325_);
  and g_147334_(_088993_, _091611_, _092327_);
  or g_147335_(_091609_, _092327_, _092328_);
  and g_147336_(_088985_, _088988_, _092329_);
  or g_147337_(_091603_, _092329_, _092330_);
  and g_147338_(_091598_, _091602_, _092331_);
  and g_147339_(_089751_, _091582_, _092332_);
  or g_147340_(_091581_, _092332_, _092333_);
  and g_147341_(_088939_, _091555_, _092334_);
  or g_147342_(_091556_, _092334_, _092335_);
  and g_147343_(_088933_, _091547_, _092336_);
  or g_147344_(_091549_, _092336_, _092338_);
  and g_147345_(_088925_, _091542_, _092339_);
  or g_147346_(_091541_, _092339_, _092340_);
  and g_147347_(_091537_, _091539_, _092341_);
  or g_147348_(_089755_, _091532_, _092342_);
  and g_147349_(_091525_, _092342_, _092343_);
  and g_147350_(_088906_, _091516_, _092344_);
  or g_147351_(_091521_, _092344_, _092345_);
  and g_147352_(_088891_, _091504_, _092346_);
  or g_147353_(_091505_, _092346_, _092347_);
  or g_147354_(_091499_, _091500_, _092349_);
  or g_147355_(_088879_, _091494_, _092350_);
  and g_147356_(_091498_, _092350_, _092351_);
  or g_147357_(_088865_, _091488_, _092352_);
  and g_147358_(_088857_, _088862_, _092353_);
  or g_147359_(_091487_, _092353_, _092354_);
  or g_147360_(_088856_, _091484_, _092355_);
  and g_147361_(_091485_, _092355_, _092356_);
  or g_147362_(_091477_, _091482_, _092357_);
  or g_147363_(_091473_, _091475_, _092358_);
  and g_147364_(_091468_, _091472_, _092360_);
  and g_147365_(_088840_, _091463_, _092361_);
  or g_147366_(_091450_, _091455_, _092362_);
  or g_147367_(_091433_, _091437_, _092363_);
  and g_147368_(_091434_, _092363_, _092364_);
  or g_147369_(_091409_, _091412_, _092365_);
  and g_147370_(_089770_, _091401_, _092366_);
  or g_147371_(_091402_, _092366_, _092367_);
  or g_147372_(_088743_, _091391_, _092368_);
  and g_147373_(_091393_, _092368_, _092369_);
  or g_147374_(_091384_, _091387_, _092371_);
  and g_147375_(_091385_, _092371_, _092372_);
  or g_147376_(_089778_, _091382_, _092373_);
  or g_147377_(_091374_, _091376_, _092374_);
  and g_147378_(_088708_, _091372_, _092375_);
  or g_147379_(_091373_, _092375_, _092376_);
  or g_147380_(_089782_, _091362_, _092377_);
  and g_147381_(_091363_, _092377_, _092378_);
  and g_147382_(_089784_, _091357_, _092379_);
  or g_147383_(_091358_, _092379_, _092380_);
  and g_147384_(_088685_, _091352_, _092382_);
  or g_147385_(_088680_, _091350_, _092383_);
  and g_147386_(_091349_, _092383_, _092384_);
  and g_147387_(_088672_, _091339_, _092385_);
  or g_147388_(_091338_, _092385_, _092386_);
  and g_147389_(_088661_, _091332_, _092387_);
  and g_147390_(_091306_, _091309_, _092388_);
  and g_147391_(_088624_, _091294_, _092389_);
  or g_147392_(_091288_, _092389_, _092390_);
  and g_147393_(_088617_, _091285_, _092391_);
  or g_147394_(_091281_, _092391_, _092393_);
  and g_147395_(_088609_, _091278_, _092394_);
  and g_147396_(_088601_, _088606_, _092395_);
  not g_147397_(_092395_, _092396_);
  and g_147398_(_091277_, _092396_, _092397_);
  and g_147399_(_089795_, _091273_, _092398_);
  or g_147400_(_091275_, _092398_, _092399_);
  or g_147401_(_088595_, _091268_, _092400_);
  and g_147402_(_091267_, _092400_, _092401_);
  or g_147403_(_088585_, _091259_, _092402_);
  and g_147404_(_091262_, _092402_, _092404_);
  and g_147405_(_089806_, _091253_, _092405_);
  or g_147406_(_091254_, _092405_, _092406_);
  or g_147407_(_088574_, _091246_, _092407_);
  or g_147408_(_088571_, _091243_, _092408_);
  and g_147409_(_091244_, _092408_, _092409_);
  or g_147410_(_088560_, _091235_, _092410_);
  and g_147411_(_091236_, _092410_, _092411_);
  or g_147412_(_088542_, _091226_, _092412_);
  and g_147413_(_091225_, _092412_, _092413_);
  and g_147414_(_089815_, _091220_, _092415_);
  or g_147415_(_091219_, _092415_, _092416_);
  and g_147416_(_088525_, _091208_, _092417_);
  and g_147417_(_088517_, _091204_, _092418_);
  or g_147418_(_091206_, _092418_, _092419_);
  or g_147419_(_088497_, _091185_, _092420_);
  and g_147420_(_091186_, _092420_, _092421_);
  and g_147421_(_089832_, _091176_, _092422_);
  or g_147422_(_091179_, _092422_, _092423_);
  and g_147423_(_091140_, _091147_, _092424_);
  or g_147424_(_089840_, _091134_, _092426_);
  and g_147425_(_091135_, _092426_, _092427_);
  or g_147426_(_088448_, _091116_, _092428_);
  and g_147427_(_088444_, _091114_, _092429_);
  or g_147428_(_091115_, _092429_, _092430_);
  and g_147429_(_089845_, _091109_, _092431_);
  or g_147430_(_091108_, _092431_, _092432_);
  and g_147431_(_088427_, _091102_, _092433_);
  or g_147432_(_091101_, _092433_, _092434_);
  or g_147433_(_088419_, _091098_, _092435_);
  and g_147434_(_091097_, _092435_, _092437_);
  and g_147435_(_088388_, _088396_, _092438_);
  or g_147436_(_091079_, _092438_, _092439_);
  and g_147437_(_091075_, _091078_, _092440_);
  or g_147438_(_088366_, _091066_, _092441_);
  and g_147439_(_091065_, _092441_, _092442_);
  or g_147440_(_091056_, _091061_, _092443_);
  and g_147441_(_091050_, _091053_, _092444_);
  and g_147442_(_089853_, _091017_, _092445_);
  or g_147443_(_091019_, _092445_, _092446_);
  and g_147444_(_091008_, _091011_, _092448_);
  or g_147445_(_091014_, _092448_, _092449_);
  and g_147446_(_088327_, _091005_, _092450_);
  or g_147447_(_091006_, _092450_, _092451_);
  and g_147448_(_088320_, _090998_, _092452_);
  or g_147449_(_090999_, _092452_, _092453_);
  or g_147450_(_090988_, _090993_, _092454_);
  and g_147451_(_090957_, _090967_, _092455_);
  or g_147452_(_088272_, _090953_, _092456_);
  and g_147453_(_090954_, _092456_, _092457_);
  and g_147454_(_089861_, _090942_, _092459_);
  or g_147455_(_090943_, _092459_, _092460_);
  and g_147456_(_088259_, _090938_, _092461_);
  or g_147457_(_090937_, _092461_, _092462_);
  or g_147458_(_088251_, _090934_, _092463_);
  and g_147459_(_088242_, _090927_, _092464_);
  or g_147460_(_088228_, _090920_, _092465_);
  or g_147461_(_088223_, _090917_, _092466_);
  and g_147462_(_090918_, _092466_, _092467_);
  and g_147463_(_090912_, _090914_, _092468_);
  and g_147464_(_089865_, _090901_, _092470_);
  or g_147465_(_090902_, _092470_, _092471_);
  and g_147466_(_088168_, _090867_, _092472_);
  or g_147467_(_090870_, _092472_, _092473_);
  or g_147468_(_088165_, _090863_, _092474_);
  and g_147469_(_090865_, _092474_, _092475_);
  and g_147470_(_089883_, _090857_, _092476_);
  or g_147471_(_090856_, _092476_, _092477_);
  and g_147472_(_090844_, _090847_, _092478_);
  and g_147473_(_088144_, _090838_, _092479_);
  or g_147474_(_090836_, _092479_, _092481_);
  or g_147475_(_088138_, _090830_, _092482_);
  and g_147476_(_090826_, _092482_, _092483_);
  and g_147477_(_090824_, _090828_, _092484_);
  and g_147478_(_089889_, _090813_, _092485_);
  or g_147479_(_090816_, _092485_, _092486_);
  or g_147480_(_088116_, _090810_, _092487_);
  and g_147481_(_090802_, _092487_, _092488_);
  and g_147482_(_090794_, _090804_, _092489_);
  or g_147483_(_090799_, _092489_, _092490_);
  and g_147484_(_090790_, _090792_, _092492_);
  and g_147485_(_090778_, _090784_, _092493_);
  or g_147486_(_088089_, _090773_, _092494_);
  or g_147487_(_088075_, _090764_, _092495_);
  and g_147488_(_090766_, _092495_, _092496_);
  and g_147489_(_088069_, _090761_, _092497_);
  or g_147490_(_090760_, _092497_, _092498_);
  or g_147491_(_088052_, _090738_, _092499_);
  and g_147492_(_090739_, _092499_, _092500_);
  and g_147493_(_088046_, _090735_, _092501_);
  or g_147494_(_090734_, _092501_, _092503_);
  or g_147495_(_088029_, _090723_, _092504_);
  and g_147496_(_090722_, _092504_, _092505_);
  and g_147497_(_088021_, _090718_, _092506_);
  or g_147498_(_090694_, _090713_, _092507_);
  and g_147499_(_090690_, _090695_, _092508_);
  or g_147500_(_090689_, _092508_, _092509_);
  or g_147501_(_090679_, _090681_, _092510_);
  or g_147502_(_087981_, _090672_, _092511_);
  and g_147503_(_087979_, _090671_, _092512_);
  or g_147504_(_090670_, _092512_, _092514_);
  or g_147505_(_087969_, _090656_, _092515_);
  and g_147506_(_090658_, _092515_, _092516_);
  and g_147507_(_089917_, _090647_, _092517_);
  or g_147508_(_090650_, _092517_, _092518_);
  or g_147509_(_087958_, _090640_, _092519_);
  or g_147510_(_087956_, _090636_, _092520_);
  and g_147511_(_090639_, _092520_, _092521_);
  and g_147512_(_087951_, _090630_, _092522_);
  or g_147513_(_090631_, _092522_, _092523_);
  or g_147514_(_087938_, _090626_, _092525_);
  and g_147515_(_090627_, _092525_, _092526_);
  or g_147516_(_089921_, _090619_, _092527_);
  and g_147517_(_090612_, _092527_, _092528_);
  and g_147518_(_087924_, _090605_, _092529_);
  or g_147519_(_090606_, _092529_, _092530_);
  or g_147520_(_087915_, _090597_, _092531_);
  and g_147521_(_090601_, _092531_, _092532_);
  and g_147522_(_087912_, _090594_, _092533_);
  or g_147523_(_090591_, _092533_, _092534_);
  or g_147524_(_087898_, _090586_, _092536_);
  and g_147525_(_090587_, _092536_, _092537_);
  and g_147526_(_087888_, _090577_, _092538_);
  or g_147527_(_090576_, _092538_, _092539_);
  or g_147528_(_089933_, _090571_, _092540_);
  and g_147529_(_090572_, _092540_, _092541_);
  or g_147530_(_087870_, _090551_, _092542_);
  and g_147531_(_087867_, _090549_, _092543_);
  or g_147532_(_090550_, _092543_, _092544_);
  and g_147533_(_089939_, _090543_, _092545_);
  or g_147534_(_090542_, _092545_, _092547_);
  and g_147535_(_089943_, _090538_, _092548_);
  or g_147536_(_090539_, _092548_, _092549_);
  and g_147537_(_087831_, _090532_, _092550_);
  or g_147538_(_087825_, _090531_, _092551_);
  and g_147539_(_090530_, _092551_, _092552_);
  or g_147540_(_087819_, _090527_, _092553_);
  and g_147541_(_090526_, _092553_, _092554_);
  or g_147542_(_089946_, _090524_, _092555_);
  and g_147543_(_087810_, _087813_, _092556_);
  or g_147544_(_090520_, _092556_, _092558_);
  or g_147545_(_089950_, _090513_, _092559_);
  and g_147546_(_090516_, _092559_, _092560_);
  or g_147547_(_087797_, _090509_, _092561_);
  and g_147548_(_090507_, _092561_, _092562_);
  or g_147549_(_089958_, _090492_, _092563_);
  and g_147550_(_090491_, _092563_, _092564_);
  and g_147551_(_090486_, _090488_, _092565_);
  or g_147552_(_089967_, _090475_, _092566_);
  and g_147553_(_090478_, _092566_, _092567_);
  and g_147554_(_087759_, _090471_, _092569_);
  or g_147555_(_090472_, _092569_, _092570_);
  or g_147556_(_090466_, _090469_, _092571_);
  and g_147557_(_090456_, _090464_, _092572_);
  and g_147558_(_089977_, _090431_, _092573_);
  or g_147559_(_090438_, _092573_, _092574_);
  and g_147560_(_090426_, _090433_, _092575_);
  and g_147561_(_090418_, _090421_, _092576_);
  and g_147562_(_090408_, _090412_, _092577_);
  or g_147563_(_089982_, _090401_, _092578_);
  and g_147564_(_090403_, _092578_, _092580_);
  or g_147565_(_087693_, _090387_, _092581_);
  and g_147566_(_090388_, _092581_, _092582_);
  or g_147567_(_089991_, _090381_, _092583_);
  and g_147568_(_090382_, _092583_, _092584_);
  and g_147569_(_087681_, _090376_, _092585_);
  or g_147570_(_087677_, _090375_, _092586_);
  and g_147571_(_090374_, _092586_, _092587_);
  and g_147572_(_087668_, _090371_, _092588_);
  or g_147573_(_090368_, _092588_, _092589_);
  and g_147574_(_087656_, _090360_, _092591_);
  or g_147575_(_090359_, _092591_, _092592_);
  or g_147576_(_087645_, _090350_, _092593_);
  and g_147577_(_090351_, _092593_, _092594_);
  or g_147578_(_087634_, _090342_, _092595_);
  and g_147579_(_090343_, _092595_, _092596_);
  or g_147580_(_087619_, _090332_, _092597_);
  or g_147581_(_087613_, _090330_, _092598_);
  and g_147582_(_090329_, _092598_, _092599_);
  and g_147583_(_090299_, _090301_, _092600_);
  and g_147584_(_090293_, _090295_, _092602_);
  and g_147585_(_090287_, _090290_, _092603_);
  or g_147586_(_087540_, _087541_, _092604_);
  not g_147587_(_092604_, _092605_);
  and g_147588_(_090280_, _092605_, _092606_);
  or g_147589_(_084657_, _087540_, _092607_);
  and g_147590_(_087538_, _090277_, _092608_);
  and g_147591_(_092607_, _092608_, _092609_);
  or g_147592_(_090278_, _092609_, _092610_);
  or g_147593_(_090264_, _090267_, _092611_);
  and g_147594_(_090260_, _090262_, _092613_);
  and g_147595_(_090253_, _090256_, _092614_);
  or g_147596_(_087502_, _090240_, _092615_);
  and g_147597_(_090241_, _092615_, _092616_);
  and g_147598_(_087493_, _090222_, _092617_);
  or g_147599_(_090232_, _092617_, _092618_);
  or g_147600_(_090216_, _090225_, _092619_);
  or g_147601_(_090205_, _090208_, _092620_);
  and g_147602_(_090197_, _090199_, _092621_);
  or g_147603_(_087472_, _090195_, _092622_);
  and g_147604_(_090188_, _092622_, _092624_);
  or g_147605_(_090185_, _090189_, _092625_);
  and g_147606_(_090181_, _092625_, _092626_);
  or g_147607_(_087464_, _090177_, _092627_);
  and g_147608_(_090178_, _092627_, _092628_);
  or g_147609_(_087457_, _090173_, _092629_);
  and g_147610_(_090169_, _092629_, _092630_);
  or g_147611_(_090166_, _090170_, _092631_);
  and g_147612_(_087417_, _090150_, _092632_);
  and g_147613_(_087410_, _087414_, _092633_);
  or g_147614_(_090146_, _092633_, _092635_);
  and g_147615_(_072873_, _075794_, _092636_);
  not g_147616_(_092636_, _092637_);
  or g_147617_(_078734_, _092637_, _092638_);
  or g_147618_(_084490_, _092638_, _092639_);
  or g_147619_(_081598_, _092639_, _092640_);
  or g_147620_(_087385_, _092640_, _092641_);
  and g_147621_(_090130_, _092641_, _092642_);
  or g_147622_(_068062_, _090131_, _092643_);
  or g_147623_(_092642_, _092643_, _092644_);
  and g_147624_(_090037_, _092644_, _092646_);
  not g_147625_(_092646_, _092647_);
  or g_147626_(_090037_, _092644_, _092648_);
  and g_147627_(_068026_, _092648_, _092649_);
  and g_147628_(_092647_, _092649_, _092650_);
  or g_147629_(_067951_, _090135_, _092651_);
  or g_147630_(_087395_, _092651_, _092652_);
  or g_147631_(_092650_, _092652_, _092653_);
  and g_147632_(_090137_, _092653_, _092654_);
  and g_147633_(_090141_, _092654_, _092655_);
  or g_147634_(_067914_, _092655_, _092657_);
  or g_147635_(_084521_, _087401_, _092658_);
  or g_147636_(_090144_, _092658_, _092659_);
  and g_147637_(_092657_, _092659_, _092660_);
  or g_147638_(_092657_, _092659_, _092661_);
  not g_147639_(_092661_, _092662_);
  or g_147640_(_067876_, _092662_, _092663_);
  or g_147641_(_092660_, _092663_, _092664_);
  xor g_147642_(_092635_, _092664_, _092665_);
  xor g_147643_(_092632_, _092665_, _092666_);
  xor g_147644_(_090152_, _092666_, _092668_);
  and g_147645_(_090155_, _092668_, _092669_);
  or g_147646_(_087435_, _090158_, _092670_);
  and g_147647_(_090161_, _092670_, _092671_);
  xor g_147648_(_092669_, _092671_, _092672_);
  xor g_147649_(_090164_, _092672_, _092673_);
  xor g_147650_(_092631_, _092673_, _092674_);
  xor g_147651_(_092630_, _092674_, _092675_);
  xor g_147652_(_092628_, _092675_, _092676_);
  xor g_147653_(_092626_, _092676_, _092677_);
  xor g_147654_(_092624_, _092677_, _092679_);
  xor g_147655_(_092621_, _092679_, _092680_);
  or g_147656_(_087478_, _090203_, _092681_);
  and g_147657_(_090202_, _092681_, _092682_);
  xor g_147658_(_092680_, _092682_, _092683_);
  xor g_147659_(_092620_, _092683_, _092684_);
  xor g_147660_(_090212_, _092684_, _092685_);
  xor g_147661_(_092619_, _092685_, _092686_);
  xor g_147662_(_092618_, _092686_, _092687_);
  xor g_147663_(_090238_, _092687_, _092688_);
  xor g_147664_(_092616_, _092688_, _092690_);
  or g_147665_(_087509_, _090242_, _092691_);
  and g_147666_(_090247_, _092691_, _092692_);
  xor g_147667_(_092690_, _092692_, _092693_);
  xor g_147668_(_092614_, _092693_, _092694_);
  xor g_147669_(_092613_, _092694_, _092695_);
  xor g_147670_(_092611_, _092695_, _092696_);
  xor g_147671_(_090272_, _092696_, _092697_);
  xor g_147672_(_090274_, _092697_, _092698_);
  xor g_147673_(_092610_, _092698_, _092699_);
  xor g_147674_(_092606_, _092699_, _092701_);
  xor g_147675_(_090283_, _092701_, _092702_);
  xor g_147676_(_092603_, _092702_, _092703_);
  xor g_147677_(_092602_, _092703_, _092704_);
  xor g_147678_(_090297_, _092704_, _092705_);
  xor g_147679_(_092600_, _092705_, _092706_);
  or g_147680_(_090304_, _090307_, _092707_);
  and g_147681_(_090305_, _092707_, _092708_);
  xor g_147682_(_092706_, _092708_, _092709_);
  and g_147683_(_090313_, _090318_, _092710_);
  or g_147684_(_090311_, _092710_, _092712_);
  or g_147685_(_090310_, _090317_, _092713_);
  and g_147686_(_092712_, _092713_, _092714_);
  xor g_147687_(_092709_, _092714_, _092715_);
  and g_147688_(_089999_, _090324_, _092716_);
  or g_147689_(_090326_, _092716_, _092717_);
  and g_147690_(_087602_, _090321_, _092718_);
  or g_147691_(_090320_, _092718_, _092719_);
  xor g_147692_(_092717_, _092719_, _092720_);
  xor g_147693_(_092715_, _092720_, _092721_);
  xor g_147694_(_092599_, _092721_, _092723_);
  xor g_147695_(_092597_, _092723_, _092724_);
  xor g_147696_(_090338_, _092724_, _092725_);
  xor g_147697_(_092596_, _092725_, _092726_);
  xor g_147698_(_092594_, _092726_, _092727_);
  xor g_147699_(_090356_, _092727_, _092728_);
  xor g_147700_(_092592_, _092728_, _092729_);
  or g_147701_(_087659_, _090361_, _092730_);
  and g_147702_(_090366_, _092730_, _092731_);
  xor g_147703_(_092729_, _092731_, _092732_);
  xor g_147704_(_092589_, _092732_, _092734_);
  xor g_147705_(_092587_, _092734_, _092735_);
  xor g_147706_(_092585_, _092735_, _092736_);
  xor g_147707_(_092584_, _092736_, _092737_);
  xor g_147708_(_090385_, _092737_, _092738_);
  xor g_147709_(_092582_, _092738_, _092739_);
  xor g_147710_(_090392_, _092739_, _092740_);
  and g_147711_(_090395_, _090398_, _092741_);
  xor g_147712_(_092740_, _092741_, _092742_);
  xor g_147713_(_092580_, _092742_, _092743_);
  xor g_147714_(_092577_, _092743_, _092745_);
  xor g_147715_(_090416_, _092745_, _092746_);
  xor g_147716_(_092576_, _092746_, _092747_);
  xor g_147717_(_092575_, _092747_, _092748_);
  xor g_147718_(_092574_, _092748_, _092749_);
  xor g_147719_(_090452_, _092749_, _092750_);
  xor g_147720_(_092572_, _092750_, _092751_);
  xor g_147721_(_092571_, _092751_, _092752_);
  xor g_147722_(_092570_, _092752_, _092753_);
  xor g_147723_(_092567_, _092753_, _092754_);
  xor g_147724_(_090483_, _092754_, _092756_);
  xor g_147725_(_092565_, _092756_, _092757_);
  xor g_147726_(_092564_, _092757_, _092758_);
  or g_147727_(_089956_, _090496_, _092759_);
  and g_147728_(_090495_, _092759_, _092760_);
  xor g_147729_(_092758_, _092760_, _092761_);
  xor g_147730_(_090499_, _092761_, _092762_);
  and g_147731_(_087791_, _090503_, _092763_);
  or g_147732_(_090502_, _092763_, _092764_);
  xor g_147733_(_092762_, _092764_, _092765_);
  xor g_147734_(_092562_, _092765_, _092767_);
  xor g_147735_(_092560_, _092767_, _092768_);
  and g_147736_(_087806_, _089948_, _092769_);
  or g_147737_(_090518_, _092769_, _092770_);
  xor g_147738_(_092768_, _092770_, _092771_);
  xor g_147739_(_092558_, _092771_, _092772_);
  xor g_147740_(_092555_, _092772_, _092773_);
  xor g_147741_(_092554_, _092773_, _092774_);
  xor g_147742_(_092552_, _092774_, _092775_);
  xor g_147743_(_092550_, _092775_, _092776_);
  xor g_147744_(_092549_, _092776_, _092778_);
  xor g_147745_(_092547_, _092778_, _092779_);
  xor g_147746_(_090547_, _092779_, _092780_);
  xor g_147747_(_092544_, _092780_, _092781_);
  xor g_147748_(_092542_, _092781_, _092782_);
  and g_147749_(_089936_, _090566_, _092783_);
  or g_147750_(_090565_, _092783_, _092784_);
  and g_147751_(_090554_, _090562_, _092785_);
  xor g_147752_(_092784_, _092785_, _092786_);
  xor g_147753_(_092782_, _092786_, _092787_);
  xor g_147754_(_092541_, _092787_, _092789_);
  xor g_147755_(_092539_, _092789_, _092790_);
  and g_147756_(_087891_, _087894_, _092791_);
  and g_147757_(_090579_, _092791_, _092792_);
  or g_147758_(_090584_, _092792_, _092793_);
  xor g_147759_(_092790_, _092793_, _092794_);
  xor g_147760_(_092537_, _092794_, _092795_);
  xor g_147761_(_092534_, _092795_, _092796_);
  xor g_147762_(_092532_, _092796_, _092797_);
  xor g_147763_(_090603_, _092797_, _092798_);
  xor g_147764_(_092530_, _092798_, _092800_);
  xor g_147765_(_090615_, _092800_, _092801_);
  xor g_147766_(_092528_, _092801_, _092802_);
  xor g_147767_(_090624_, _092802_, _092803_);
  xor g_147768_(_092526_, _092803_, _092804_);
  xor g_147769_(_092523_, _092804_, _092805_);
  xor g_147770_(_092521_, _092805_, _092806_);
  xor g_147771_(_092519_, _092806_, _092807_);
  xor g_147772_(_090648_, _092807_, _092808_);
  xor g_147773_(_092518_, _092808_, _092809_);
  xor g_147774_(_092516_, _092809_, _092811_);
  xor g_147775_(_090668_, _092811_, _092812_);
  xor g_147776_(_092514_, _092812_, _092813_);
  xor g_147777_(_092511_, _092813_, _092814_);
  xor g_147778_(_090676_, _092814_, _092815_);
  xor g_147779_(_092510_, _092815_, _092816_);
  xor g_147780_(_090683_, _092816_, _092817_);
  xor g_147781_(_090686_, _092817_, _092818_);
  xor g_147782_(_092509_, _092818_, _092819_);
  xor g_147783_(_092507_, _092819_, _092820_);
  or g_147784_(_088014_, _090716_, _092822_);
  and g_147785_(_090717_, _092822_, _092823_);
  xor g_147786_(_092820_, _092823_, _092824_);
  xor g_147787_(_092506_, _092824_, _092825_);
  xor g_147788_(_092505_, _092825_, _092826_);
  xor g_147789_(_090726_, _092826_, _092827_);
  xor g_147790_(_090731_, _092827_, _092828_);
  xor g_147791_(_092503_, _092828_, _092829_);
  xor g_147792_(_092500_, _092829_, _092830_);
  or g_147793_(_088056_, _090747_, _092831_);
  and g_147794_(_090748_, _092831_, _092833_);
  xor g_147795_(_092830_, _092833_, _092834_);
  or g_147796_(_088059_, _090750_, _092835_);
  and g_147797_(_090756_, _092835_, _092836_);
  xor g_147798_(_090758_, _092836_, _092837_);
  xor g_147799_(_092834_, _092837_, _092838_);
  xor g_147800_(_092498_, _092838_, _092839_);
  xor g_147801_(_092496_, _092839_, _092840_);
  xor g_147802_(_090769_, _092840_, _092841_);
  or g_147803_(_088087_, _090772_, _092842_);
  and g_147804_(_090771_, _092842_, _092844_);
  xor g_147805_(_092841_, _092844_, _092845_);
  xor g_147806_(_092494_, _092845_, _092846_);
  xor g_147807_(_092493_, _092846_, _092847_);
  xor g_147808_(_090788_, _092847_, _092848_);
  xor g_147809_(_092492_, _092848_, _092849_);
  xor g_147810_(_090796_, _092849_, _092850_);
  xor g_147811_(_092490_, _092850_, _092851_);
  xor g_147812_(_092488_, _092851_, _092852_);
  xor g_147813_(_092486_, _092852_, _092853_);
  xor g_147814_(_090821_, _092853_, _092855_);
  xor g_147815_(_092484_, _092855_, _092856_);
  xor g_147816_(_092483_, _092856_, _092857_);
  xor g_147817_(_092481_, _092857_, _092858_);
  xor g_147818_(_092478_, _092858_, _092859_);
  xor g_147819_(_090861_, _092859_, _092860_);
  xor g_147820_(_092477_, _092860_, _092861_);
  xor g_147821_(_092475_, _092861_, _092862_);
  xor g_147822_(_092473_, _092862_, _092863_);
  and g_147823_(_090874_, _090878_, _092864_);
  xor g_147824_(_092863_, _092864_, _092866_);
  xor g_147825_(_090880_, _092866_, _092867_);
  xor g_147826_(_090884_, _092867_, _092868_);
  or g_147827_(_089873_, _090888_, _092869_);
  and g_147828_(_090883_, _092869_, _092870_);
  xor g_147829_(_092868_, _092870_, _092871_);
  xor g_147830_(_090892_, _092871_, _092872_);
  and g_147831_(_089867_, _090894_, _092873_);
  or g_147832_(_090895_, _092873_, _092874_);
  xor g_147833_(_092872_, _092874_, _092875_);
  xor g_147834_(_090899_, _092875_, _092877_);
  xor g_147835_(_092471_, _092877_, _092878_);
  xor g_147836_(_090906_, _092878_, _092879_);
  xor g_147837_(_092468_, _092879_, _092880_);
  xor g_147838_(_092467_, _092880_, _092881_);
  xor g_147839_(_092465_, _092881_, _092882_);
  xor g_147840_(_090923_, _092882_, _092883_);
  or g_147841_(_088238_, _090926_, _092884_);
  and g_147842_(_090925_, _092884_, _092885_);
  xor g_147843_(_092883_, _092885_, _092886_);
  xor g_147844_(_092464_, _092886_, _092888_);
  or g_147845_(_088249_, _090932_, _092889_);
  and g_147846_(_090931_, _092889_, _092890_);
  xor g_147847_(_092888_, _092890_, _092891_);
  xor g_147848_(_092463_, _092891_, _092892_);
  xor g_147849_(_092462_, _092892_, _092893_);
  xor g_147850_(_092460_, _092893_, _092894_);
  xor g_147851_(_090950_, _092894_, _092895_);
  xor g_147852_(_092457_, _092895_, _092896_);
  xor g_147853_(_092455_, _092896_, _092897_);
  and g_147854_(_090972_, _090976_, _092899_);
  xor g_147855_(_090970_, _092899_, _092900_);
  xor g_147856_(_092897_, _092900_, _092901_);
  xor g_147857_(_090982_, _092901_, _092902_);
  xor g_147858_(_090984_, _092902_, _092903_);
  xor g_147859_(_092454_, _092903_, _092904_);
  xor g_147860_(_092453_, _092904_, _092905_);
  xor g_147861_(_091003_, _092905_, _092906_);
  xor g_147862_(_092451_, _092906_, _092907_);
  xor g_147863_(_092449_, _092907_, _092908_);
  xor g_147864_(_092446_, _092908_, _092910_);
  or g_147865_(_088337_, _091028_, _092911_);
  and g_147866_(_091027_, _092911_, _092912_);
  xor g_147867_(_092910_, _092912_, _092913_);
  xor g_147868_(_091044_, _092913_, _092914_);
  xor g_147869_(_092444_, _092914_, _092915_);
  xor g_147870_(_092443_, _092915_, _092916_);
  xor g_147871_(_092442_, _092916_, _092917_);
  xor g_147872_(_091070_, _092917_, _092918_);
  xor g_147873_(_092440_, _092918_, _092919_);
  xor g_147874_(_091082_, _092919_, _092921_);
  xor g_147875_(_092439_, _092921_, _092922_);
  xor g_147876_(_091089_, _092922_, _092923_);
  and g_147877_(_091092_, _091094_, _092924_);
  xor g_147878_(_092923_, _092924_, _092925_);
  xor g_147879_(_092437_, _092925_, _092926_);
  xor g_147880_(_092434_, _092926_, _092927_);
  xor g_147881_(_091105_, _092927_, _092928_);
  xor g_147882_(_092432_, _092928_, _092929_);
  xor g_147883_(_091112_, _092929_, _092930_);
  xor g_147884_(_092430_, _092930_, _092932_);
  xor g_147885_(_092428_, _092932_, _092933_);
  or g_147886_(_088455_, _091122_, _092934_);
  and g_147887_(_091121_, _092934_, _092935_);
  xor g_147888_(_092933_, _092935_, _092936_);
  or g_147889_(_088458_, _091123_, _092937_);
  and g_147890_(_091130_, _092937_, _092938_);
  xor g_147891_(_091129_, _092938_, _092939_);
  xor g_147892_(_092936_, _092939_, _092940_);
  xor g_147893_(_092427_, _092940_, _092941_);
  xor g_147894_(_092424_, _092941_, _092943_);
  and g_147895_(_091156_, _091163_, _092944_);
  xor g_147896_(_092943_, _092944_, _092945_);
  and g_147897_(_091168_, _091170_, _092946_);
  xor g_147898_(_092945_, _092946_, _092947_);
  or g_147899_(_088488_, _091173_, _092948_);
  and g_147900_(_091174_, _092948_, _092949_);
  xor g_147901_(_092947_, _092949_, _092950_);
  xor g_147902_(_092423_, _092950_, _092951_);
  xor g_147903_(_091182_, _092951_, _092952_);
  xor g_147904_(_092421_, _092952_, _092954_);
  and g_147905_(_088505_, _091195_, _092955_);
  or g_147906_(_091200_, _092955_, _092956_);
  and g_147907_(_091189_, _091197_, _092957_);
  or g_147908_(_091192_, _092957_, _092958_);
  xor g_147909_(_092956_, _092958_, _092959_);
  xor g_147910_(_092954_, _092959_, _092960_);
  xor g_147911_(_092419_, _092960_, _092961_);
  xor g_147912_(_092417_, _092961_, _092962_);
  xor g_147913_(_091211_, _092962_, _092963_);
  xor g_147914_(_091214_, _092963_, _092965_);
  xor g_147915_(_091217_, _092965_, _092966_);
  xor g_147916_(_092416_, _092966_, _092967_);
  xor g_147917_(_091223_, _092967_, _092968_);
  xor g_147918_(_092413_, _092968_, _092969_);
  or g_147919_(_088547_, _091228_, _092970_);
  and g_147920_(_091233_, _092970_, _092971_);
  xor g_147921_(_092969_, _092971_, _092972_);
  xor g_147922_(_092411_, _092972_, _092973_);
  xor g_147923_(_091241_, _092973_, _092974_);
  xor g_147924_(_092409_, _092974_, _092976_);
  xor g_147925_(_092407_, _092976_, _092977_);
  xor g_147926_(_091251_, _092977_, _092978_);
  xor g_147927_(_092406_, _092978_, _092979_);
  xor g_147928_(_092404_, _092979_, _092980_);
  xor g_147929_(_091265_, _092980_, _092981_);
  xor g_147930_(_092401_, _092981_, _092982_);
  xor g_147931_(_092399_, _092982_, _092983_);
  xor g_147932_(_092397_, _092983_, _092984_);
  xor g_147933_(_092394_, _092984_, _092985_);
  xor g_147934_(_092393_, _092985_, _092987_);
  xor g_147935_(_092390_, _092987_, _092988_);
  and g_147936_(_091297_, _091300_, _092989_);
  xor g_147937_(_092988_, _092989_, _092990_);
  xor g_147938_(_091302_, _092990_, _092991_);
  xor g_147939_(_092388_, _092991_, _092992_);
  xor g_147940_(_091313_, _092992_, _092993_);
  and g_147941_(_091317_, _091327_, _092994_);
  xor g_147942_(_092993_, _092994_, _092995_);
  or g_147943_(_088658_, _091331_, _092996_);
  and g_147944_(_091330_, _092996_, _092998_);
  xor g_147945_(_092995_, _092998_, _092999_);
  xor g_147946_(_092387_, _092999_, _093000_);
  xor g_147947_(_091335_, _093000_, _093001_);
  xor g_147948_(_092386_, _093001_, _093002_);
  xor g_147949_(_092384_, _093002_, _093003_);
  xor g_147950_(_092382_, _093003_, _093004_);
  xor g_147951_(_092380_, _093004_, _093005_);
  xor g_147952_(_092378_, _093005_, _093006_);
  xor g_147953_(_091369_, _093006_, _093007_);
  xor g_147954_(_092376_, _093007_, _093009_);
  xor g_147955_(_092374_, _093009_, _093010_);
  and g_147956_(_088715_, _088721_, _093011_);
  not g_147957_(_093011_, _093012_);
  and g_147958_(_091379_, _093012_, _093013_);
  xor g_147959_(_093010_, _093013_, _093014_);
  xor g_147960_(_092373_, _093014_, _093015_);
  xor g_147961_(_092372_, _093015_, _093016_);
  xor g_147962_(_091389_, _093016_, _093017_);
  xor g_147963_(_092369_, _093017_, _093018_);
  xor g_147964_(_091396_, _093018_, _093020_);
  xor g_147965_(_091399_, _093020_, _093021_);
  xor g_147966_(_092367_, _093021_, _093022_);
  xor g_147967_(_091407_, _093022_, _093023_);
  xor g_147968_(_092365_, _093023_, _093024_);
  xor g_147969_(_091417_, _093024_, _093025_);
  xor g_147970_(_091422_, _093025_, _093026_);
  and g_147971_(_088783_, _091421_, _093027_);
  or g_147972_(_091424_, _093027_, _093028_);
  and g_147973_(_088790_, _091427_, _093029_);
  or g_147974_(_091431_, _093029_, _093031_);
  xor g_147975_(_093028_, _093031_, _093032_);
  xor g_147976_(_093026_, _093032_, _093033_);
  xor g_147977_(_092364_, _093033_, _093034_);
  xor g_147978_(_091440_, _093034_, _093035_);
  or g_147979_(_088814_, _091442_, _093036_);
  and g_147980_(_091443_, _093036_, _093037_);
  xor g_147981_(_093035_, _093037_, _093038_);
  xor g_147982_(_092362_, _093038_, _093039_);
  xor g_147983_(_091459_, _093039_, _093040_);
  or g_147984_(_088836_, _091461_, _093042_);
  and g_147985_(_091462_, _093042_, _093043_);
  xor g_147986_(_093040_, _093043_, _093044_);
  xor g_147987_(_092361_, _093044_, _093045_);
  xor g_147988_(_092360_, _093045_, _093046_);
  xor g_147989_(_092358_, _093046_, _093047_);
  xor g_147990_(_092357_, _093047_, _093048_);
  xor g_147991_(_092356_, _093048_, _093049_);
  xor g_147992_(_092354_, _093049_, _093050_);
  xor g_147993_(_092352_, _093050_, _093051_);
  xor g_147994_(_091492_, _093051_, _093053_);
  xor g_147995_(_092351_, _093053_, _093054_);
  xor g_147996_(_092349_, _093054_, _093055_);
  xor g_147997_(_092347_, _093055_, _093056_);
  or g_147998_(_088898_, _088902_, _093057_);
  not g_147999_(_093057_, _093058_);
  or g_148000_(_091511_, _093058_, _093059_);
  and g_148001_(_091510_, _093059_, _093060_);
  xor g_148002_(_093056_, _093060_, _093061_);
  xor g_148003_(_092345_, _093061_, _093062_);
  xor g_148004_(_092343_, _093062_, _093064_);
  xor g_148005_(_092341_, _093064_, _093065_);
  xor g_148006_(_092340_, _093065_, _093066_);
  xor g_148007_(_092338_, _093066_, _093067_);
  xor g_148008_(_092335_, _093067_, _093068_);
  and g_148009_(_088947_, _091559_, _093069_);
  or g_148010_(_091563_, _093069_, _093070_);
  xor g_148011_(_091577_, _093070_, _093071_);
  xor g_148012_(_093068_, _093071_, _093072_);
  xor g_148013_(_092333_, _093072_, _093073_);
  xor g_148014_(_091585_, _093073_, _093075_);
  xor g_148015_(_091587_, _093075_, _093076_);
  xor g_148016_(_091596_, _093076_, _093077_);
  xor g_148017_(_092331_, _093077_, _093078_);
  xor g_148018_(_092330_, _093078_, _093079_);
  xor g_148019_(_092328_, _093079_, _093080_);
  xor g_148020_(_092325_, _093080_, _093081_);
  xor g_148021_(_092323_, _093081_, _093082_);
  or g_148022_(_091628_, _091629_, _093083_);
  or g_148023_(_089016_, _091624_, _093084_);
  and g_148024_(_091626_, _093084_, _093086_);
  xor g_148025_(_093083_, _093086_, _093087_);
  xor g_148026_(_093082_, _093087_, _093088_);
  xor g_148027_(_092321_, _093088_, _093089_);
  xor g_148028_(_092319_, _093089_, _093090_);
  xor g_148029_(_091649_, _093090_, _093091_);
  or g_148030_(_089037_, _091651_, _093092_);
  and g_148031_(_091647_, _093092_, _093093_);
  xor g_148032_(_093091_, _093093_, _093094_);
  xor g_148033_(_092318_, _093094_, _093095_);
  xor g_148034_(_092317_, _093095_, _093097_);
  xor g_148035_(_092314_, _093097_, _093098_);
  xor g_148036_(_092312_, _093098_, _093099_);
  xor g_148037_(_092311_, _093099_, _093100_);
  xor g_148038_(_091683_, _093100_, _093101_);
  xor g_148039_(_092309_, _093101_, _093102_);
  xor g_148040_(_091690_, _093102_, _093103_);
  or g_148041_(_089092_, _091693_, _093104_);
  and g_148042_(_091692_, _093104_, _093105_);
  xor g_148043_(_093103_, _093105_, _093106_);
  xor g_148044_(_092307_, _093106_, _093108_);
  and g_148045_(_089718_, _091709_, _093109_);
  or g_148046_(_091708_, _093109_, _093110_);
  xor g_148047_(_093108_, _093110_, _093111_);
  xor g_148048_(_092305_, _093111_, _093112_);
  xor g_148049_(_091718_, _093112_, _093113_);
  xor g_148050_(_091720_, _093113_, _093114_);
  xor g_148051_(_092302_, _093114_, _093115_);
  xor g_148052_(_092301_, _093115_, _093116_);
  xor g_148053_(_091747_, _093116_, _093117_);
  xor g_148054_(_091749_, _093117_, _093119_);
  or g_148055_(_089143_, _091751_, _093120_);
  and g_148056_(_091752_, _093120_, _093121_);
  xor g_148057_(_093119_, _093121_, _093122_);
  xor g_148058_(_092299_, _093122_, _093123_);
  or g_148059_(_089152_, _091767_, _093124_);
  and g_148060_(_091765_, _093124_, _093125_);
  xor g_148061_(_093123_, _093125_, _093126_);
  xor g_148062_(_092297_, _093126_, _093127_);
  xor g_148063_(_092296_, _093127_, _093128_);
  xor g_148064_(_092294_, _093128_, _093130_);
  xor g_148065_(_092291_, _093130_, _093131_);
  xor g_148066_(_092289_, _093131_, _093132_);
  xor g_148067_(_092287_, _093132_, _093133_);
  xor g_148068_(_092285_, _093133_, _093134_);
  xor g_148069_(_092283_, _093134_, _093135_);
  xor g_148070_(_092281_, _093135_, _093136_);
  xor g_148071_(_091812_, _093136_, _093137_);
  xor g_148072_(_091817_, _093137_, _093138_);
  xor g_148073_(_092279_, _093138_, _093139_);
  xor g_148074_(_091829_, _093139_, _093141_);
  xor g_148075_(_092278_, _093141_, _093142_);
  xor g_148076_(_091837_, _093142_, _093143_);
  xor g_148077_(_092276_, _093143_, _093144_);
  xor g_148078_(_091847_, _093144_, _093145_);
  and g_148079_(_091845_, _091857_, _093146_);
  xor g_148080_(_093145_, _093146_, _093147_);
  xor g_148081_(_092274_, _093147_, _093148_);
  and g_148082_(_091864_, _091867_, _093149_);
  xor g_148083_(_093148_, _093149_, _093150_);
  xor g_148084_(_091869_, _093150_, _093152_);
  xor g_148085_(_092273_, _093152_, _093153_);
  xor g_148086_(_091877_, _093153_, _093154_);
  or g_148087_(_089268_, _091880_, _093155_);
  and g_148088_(_091879_, _093155_, _093156_);
  xor g_148089_(_093154_, _093156_, _093157_);
  xor g_148090_(_091888_, _093157_, _093158_);
  xor g_148091_(_092270_, _093158_, _093159_);
  xor g_148092_(_091896_, _093159_, _093160_);
  xor g_148093_(_092269_, _093160_, _093161_);
  xor g_148094_(_092267_, _093161_, _093163_);
  xor g_148095_(_092265_, _093163_, _093164_);
  xor g_148096_(_092263_, _093164_, _093165_);
  xor g_148097_(_091921_, _093165_, _093166_);
  xor g_148098_(_091923_, _093166_, _093167_);
  xor g_148099_(_092261_, _093167_, _093168_);
  xor g_148100_(_091934_, _093168_, _093169_);
  or g_148101_(_089340_, _091936_, _093170_);
  and g_148102_(_091933_, _093170_, _093171_);
  xor g_148103_(_093169_, _093171_, _093172_);
  xor g_148104_(_091952_, _093172_, _093174_);
  xor g_148105_(_092259_, _093174_, _093175_);
  xor g_148106_(_092257_, _093175_, _093176_);
  or g_148107_(_089367_, _091963_, _093177_);
  and g_148108_(_091962_, _093177_, _093178_);
  xor g_148109_(_093176_, _093178_, _093179_);
  xor g_148110_(_091973_, _093179_, _093180_);
  xor g_148111_(_092256_, _093180_, _093181_);
  or g_148112_(_089383_, _091984_, _093182_);
  and g_148113_(_091980_, _093182_, _093183_);
  xor g_148114_(_093181_, _093183_, _093185_);
  xor g_148115_(_091991_, _093185_, _093186_);
  xor g_148116_(_092255_, _093186_, _093187_);
  xor g_148117_(_092254_, _093187_, _093188_);
  xor g_148118_(_092252_, _093188_, _093189_);
  xor g_148119_(_092250_, _093189_, _093190_);
  xor g_148120_(_092247_, _093190_, _093191_);
  xor g_148121_(_092245_, _093191_, _093192_);
  xor g_148122_(_092035_, _093192_, _093193_);
  xor g_148123_(_092243_, _093193_, _093194_);
  or g_148124_(_089447_, _092044_, _093196_);
  and g_148125_(_092043_, _093196_, _093197_);
  xor g_148126_(_093194_, _093197_, _093198_);
  xor g_148127_(_092241_, _093198_, _093199_);
  xor g_148128_(_092239_, _093199_, _093200_);
  xor g_148129_(_092236_, _093200_, _093201_);
  or g_148130_(_089481_, _092066_, _093202_);
  and g_148131_(_092068_, _093202_, _093203_);
  xor g_148132_(_093201_, _093203_, _093204_);
  or g_148133_(_089483_, _092071_, _093205_);
  xor g_148134_(_092062_, _093205_, _093207_);
  xor g_148135_(_093204_, _093207_, _093208_);
  xor g_148136_(_092077_, _093208_, _093209_);
  xor g_148137_(_092079_, _093209_, _093210_);
  or g_148138_(_089495_, _092083_, _093211_);
  and g_148139_(_092082_, _093211_, _093212_);
  xor g_148140_(_093210_, _093212_, _093213_);
  xor g_148141_(_092235_, _093213_, _093214_);
  xor g_148142_(_092234_, _093214_, _093215_);
  xor g_148143_(_092232_, _093215_, _093216_);
  or g_148144_(_089508_, _092098_, _093218_);
  and g_148145_(_092097_, _093218_, _093219_);
  xor g_148146_(_093216_, _093219_, _093220_);
  xor g_148147_(_092101_, _093220_, _093221_);
  and g_148148_(_089649_, _092106_, _093222_);
  or g_148149_(_092112_, _093222_, _093223_);
  and g_148150_(_092104_, _092108_, _093224_);
  or g_148151_(_092103_, _093224_, _093225_);
  xor g_148152_(_093223_, _093225_, _093226_);
  xor g_148153_(_093221_, _093226_, _093227_);
  xor g_148154_(_092231_, _093227_, _093229_);
  xor g_148155_(_092229_, _093229_, _093230_);
  xor g_148156_(_092226_, _093230_, _093231_);
  xor g_148157_(_092130_, _093231_, _093232_);
  xor g_148158_(_092224_, _093232_, _093233_);
  xor g_148159_(_092223_, _093233_, _093234_);
  xor g_148160_(_092141_, _093234_, _093235_);
  xor g_148161_(_092222_, _093235_, _093236_);
  xor g_148162_(_092221_, _093236_, _093237_);
  xor g_148163_(_092219_, _093237_, _093238_);
  xor g_148164_(_092218_, _093238_, _093240_);
  xor g_148165_(_092217_, _093240_, _093241_);
  and g_148166_(_092170_, _092175_, _093242_);
  xor g_148167_(_092180_, _093242_, _093243_);
  xor g_148168_(_093241_, _093243_, _093244_);
  xor g_148169_(_092214_, _093244_, _093245_);
  or g_148170_(_089619_, _092198_, _093246_);
  and g_148171_(_092191_, _093246_, _093247_);
  xor g_148172_(_093245_, _093247_, _093248_);
  xor g_148173_(_092204_, _093248_, _093249_);
  xor g_148174_(_092213_, _093249_, _093251_);
  xor g_148175_(_092211_, _093251_, out[967]);
  buf b_0_(set2[375], out[375]);
  buf b_1_(set2[91], out[91]);
  buf b_2_(set2[377], out[377]);
  buf b_3_(set1[191], out[671]);
  buf b_4_(set1[234], out[714]);
  buf b_5_(set1[235], out[715]);
  buf b_6_(set2[417], out[417]);
  buf b_7_(set1[268], out[748]);
  buf b_8_(set2[337], out[337]);
  buf b_9_(set2[349], out[349]);
  buf b_10_(set2[138], out[138]);
  buf b_11_(set2[212], out[212]);
  buf b_12_(set1[208], out[688]);
  buf b_13_(set1[447], out[927]);
  buf b_14_(set1[427], out[907]);
  buf b_15_(set1[85], out[565]);
  buf b_16_(set2[233], out[233]);
  buf b_17_(set1[413], out[893]);
  buf b_18_(set1[120], out[600]);
  buf b_19_(set1[437], out[917]);
  buf b_20_(set1[178], out[658]);
  buf b_21_(set2[92], out[92]);
  buf b_22_(set1[374], out[854]);
  buf b_23_(set2[323], out[323]);
  buf b_24_(set2[177], out[177]);
  buf b_25_(set1[101], out[581]);
  buf b_26_(set1[302], out[782]);
  buf b_27_(set2[400], out[400]);
  buf b_28_(set2[34], out[34]);
  buf b_29_(set1[100], out[580]);
  buf b_30_(set1[329], out[809]);
  buf b_31_(set2[199], out[199]);
  buf b_32_(set2[289], out[289]);
  buf b_33_(set2[242], out[242]);
  buf b_34_(set2[344], out[344]);
  buf b_35_(set1[190], out[670]);
  buf b_36_(set2[146], out[146]);
  buf b_37_(set1[358], out[838]);
  buf b_38_(set1[198], out[678]);
  buf b_39_(set1[147], out[627]);
  buf b_40_(set2[90], out[90]);
  buf b_41_(set1[119], out[599]);
  buf b_42_(set2[359], out[359]);
  buf b_43_(set2[347], out[347]);
  buf b_44_(set1[2], out[482]);
  buf b_45_(set1[376], out[856]);
  buf b_46_(set2[27], out[27]);
  buf b_47_(set2[23], out[23]);
  buf b_48_(set2[187], out[187]);
  buf b_49_(set2[468], out[468]);
  buf b_50_(set1[383], out[863]);
  buf b_51_(set1[40], out[520]);
  buf b_52_(set2[271], out[271]);
  buf b_53_(set2[179], out[179]);
  buf b_54_(set1[291], out[771]);
  buf b_55_(set2[18], out[18]);
  buf b_56_(set2[25], out[25]);
  buf b_57_(set2[208], out[208]);
  buf b_58_(set1[197], out[677]);
  buf b_59_(set2[304], out[304]);
  buf b_60_(set2[124], out[124]);
  buf b_61_(set1[157], out[637]);
  buf b_62_(set1[353], out[833]);
  buf b_63_(set1[28], out[508]);
  buf b_64_(set2[290], out[290]);
  buf b_65_(set2[389], out[389]);
  buf b_66_(set2[231], out[231]);
  buf b_67_(set1[328], out[808]);
  buf b_68_(set1[303], out[783]);
  buf b_69_(set1[49], out[529]);
  buf b_70_(set2[416], out[416]);
  buf b_71_(set1[74], out[554]);
  buf b_72_(set1[248], out[728]);
  buf b_73_(set2[38], out[38]);
  buf b_74_(set1[343], out[823]);
  buf b_75_(set2[430], out[430]);
  buf b_76_(set2[19], out[19]);
  buf b_77_(set2[350], out[350]);
  buf b_78_(set1[176], out[656]);
  buf b_79_(set1[209], out[689]);
  buf b_80_(set1[431], out[911]);
  buf b_81_(set1[267], out[747]);
  buf b_82_(set1[395], out[875]);
  buf b_83_(set2[75], out[75]);
  buf b_84_(set1[443], out[923]);
  buf b_85_(set2[232], out[232]);
  buf b_86_(set2[469], out[469]);
  buf b_87_(set1[394], out[874]);
  buf b_88_(set1[98], out[578]);
  buf b_89_(set2[110], out[110]);
  buf b_90_(set2[306], out[306]);
  buf b_91_(set2[40], out[40]);
  buf b_92_(set1[106], out[586]);
  buf b_93_(set2[246], out[246]);
  buf b_94_(set2[123], out[123]);
  buf b_95_(set1[454], out[934]);
  buf b_96_(set2[315], out[315]);
  buf b_97_(set2[425], out[425]);
  buf b_98_(set2[153], out[153]);
  buf b_99_(set2[3], out[3]);
  buf b_100_(set2[4], out[4]);
  buf b_101_(set1[420], out[900]);
  buf b_102_(set1[149], out[629]);
  buf b_103_(set2[111], out[111]);
  buf b_104_(set2[443], out[443]);
  buf b_105_(set2[135], out[135]);
  buf b_106_(set2[161], out[161]);
  buf b_107_(set2[453], out[453]);
  buf b_108_(set1[250], out[730]);
  buf b_109_(set2[478], out[478]);
  buf b_110_(set2[81], out[81]);
  buf b_111_(set1[449], out[929]);
  buf b_112_(set1[154], out[634]);
  buf b_113_(set1[232], out[712]);
  buf b_114_(set1[206], out[686]);
  buf b_115_(set1[476], out[956]);
  buf b_116_(set1[50], out[530]);
  buf b_117_(set2[48], out[48]);
  buf b_118_(set1[103], out[583]);
  buf b_119_(set2[279], out[279]);
  buf b_120_(set1[270], out[750]);
  buf b_121_(set2[403], out[403]);
  buf b_122_(set2[100], out[100]);
  buf b_123_(set2[145], out[145]);
  buf b_124_(set2[392], out[392]);
  buf b_125_(set2[472], out[472]);
  buf b_126_(set1[19], out[499]);
  buf b_127_(set2[78], out[78]);
  buf b_128_(set2[96], out[96]);
  buf b_129_(set1[419], out[899]);
  buf b_130_(set2[288], out[288]);
  buf b_131_(set1[249], out[729]);
  buf b_132_(set1[299], out[779]);
  buf b_133_(set2[310], out[310]);
  buf b_134_(set1[111], out[591]);
  buf b_135_(set2[158], out[158]);
  buf b_136_(set2[459], out[459]);
  buf b_137_(set2[131], out[131]);
  buf b_138_(set2[357], out[357]);
  buf b_139_(set1[41], out[521]);
  buf b_140_(set1[14], out[494]);
  buf b_141_(set2[421], out[421]);
  buf b_142_(set2[1], out[1]);
  buf b_143_(set2[385], out[385]);
  buf b_144_(set2[354], out[354]);
  buf b_145_(set1[217], out[697]);
  buf b_146_(set2[137], out[137]);
  buf b_147_(set2[296], out[296]);
  buf b_148_(set2[159], out[159]);
  buf b_149_(set1[458], out[938]);
  buf b_150_(set2[374], out[374]);
  buf b_151_(set2[118], out[118]);
  buf b_152_(set1[368], out[848]);
  buf b_153_(set1[324], out[804]);
  buf b_154_(set1[409], out[889]);
  buf b_155_(set2[422], out[422]);
  buf b_156_(set1[269], out[749]);
  buf b_157_(set1[18], out[498]);
  buf b_158_(set1[22], out[502]);
  buf b_159_(set2[450], out[450]);
  buf b_160_(set1[201], out[681]);
  buf b_161_(set2[446], out[446]);
  buf b_162_(set1[364], out[844]);
  buf b_163_(set1[123], out[603]);
  buf b_164_(set1[401], out[881]);
  buf b_165_(set1[417], out[897]);
  buf b_166_(set1[59], out[539]);
  buf b_167_(set1[367], out[847]);
  buf b_168_(set1[153], out[633]);
  buf b_169_(set2[141], out[141]);
  buf b_170_(set2[442], out[442]);
  buf b_171_(set2[228], out[228]);
  buf b_172_(set2[217], out[217]);
  buf b_173_(set1[45], out[525]);
  buf b_174_(set1[426], out[906]);
  buf b_175_(set1[246], out[726]);
  buf b_176_(set2[335], out[335]);
  buf b_177_(set2[284], out[284]);
  buf b_178_(set2[183], out[183]);
  buf b_179_(set1[117], out[597]);
  buf b_180_(set1[405], out[885]);
  buf b_181_(set1[371], out[851]);
  buf b_182_(set1[425], out[905]);
  buf b_183_(set2[86], out[86]);
  buf b_184_(set1[195], out[675]);
  buf b_185_(set1[169], out[649]);
  buf b_186_(set2[174], out[174]);
  buf b_187_(set2[454], out[454]);
  buf b_188_(set1[381], out[861]);
  buf b_189_(set2[407], out[407]);
  buf b_190_(set1[57], out[537]);
  buf b_191_(set1[273], out[753]);
  buf b_192_(set2[342], out[342]);
  buf b_193_(set1[172], out[652]);
  buf b_194_(set1[300], out[780]);
  buf b_195_(set2[175], out[175]);
  buf b_196_(set1[465], out[945]);
  buf b_197_(set2[45], out[45]);
  buf b_198_(set2[299], out[299]);
  buf b_199_(set1[286], out[766]);
  buf b_200_(set1[4], out[484]);
  buf b_201_(set1[142], out[622]);
  buf b_202_(set1[171], out[651]);
  buf b_203_(set2[170], out[170]);
  buf b_204_(set1[52], out[532]);
  buf b_205_(set2[195], out[195]);
  buf b_206_(set2[268], out[268]);
  buf b_207_(set1[433], out[913]);
  buf b_208_(set1[115], out[595]);
  buf b_209_(set2[24], out[24]);
  buf b_210_(set2[340], out[340]);
  buf b_211_(set1[204], out[684]);
  buf b_212_(set1[212], out[692]);
  buf b_213_(set1[393], out[873]);
  buf b_214_(set2[426], out[426]);
  buf b_215_(set1[292], out[772]);
  buf b_216_(set1[361], out[841]);
  buf b_217_(set1[313], out[793]);
  buf b_218_(set2[447], out[447]);
  buf b_219_(set1[216], out[696]);
  buf b_220_(set1[360], out[840]);
  buf b_221_(set1[48], out[528]);
  buf b_222_(set2[411], out[411]);
  buf b_223_(set1[460], out[940]);
  buf b_224_(set1[386], out[866]);
  buf b_225_(set2[281], out[281]);
  buf b_226_(set1[346], out[826]);
  buf b_227_(set1[13], out[493]);
  buf b_228_(set2[102], out[102]);
  buf b_229_(set2[151], out[151]);
  buf b_230_(set1[390], out[870]);
  buf b_231_(set2[432], out[432]);
  buf b_232_(set1[320], out[800]);
  buf b_233_(set1[63], out[543]);
  buf b_234_(set1[180], out[660]);
  buf b_235_(set1[266], out[746]);
  buf b_236_(set1[205], out[685]);
  buf b_237_(set2[241], out[241]);
  buf b_238_(set2[236], out[236]);
  buf b_239_(set2[66], out[66]);
  buf b_240_(set1[423], out[903]);
  buf b_241_(set2[178], out[178]);
  buf b_242_(set1[43], out[523]);
  buf b_243_(set1[434], out[914]);
  buf b_244_(set2[223], out[223]);
  buf b_245_(set1[424], out[904]);
  buf b_246_(set1[233], out[713]);
  buf b_247_(set2[316], out[316]);
  buf b_248_(set2[353], out[353]);
  buf b_249_(set1[173], out[653]);
  buf b_250_(set1[479], out[959]);
  buf b_251_(set2[324], out[324]);
  buf b_252_(set2[235], out[235]);
  buf b_253_(set2[140], out[140]);
  buf b_254_(set2[429], out[429]);
  buf b_255_(set2[104], out[104]);
  buf b_256_(set2[33], out[33]);
  buf b_257_(set1[75], out[555]);
  buf b_258_(set2[456], out[456]);
  buf b_259_(set1[415], out[895]);
  buf b_260_(set2[465], out[465]);
  buf b_261_(set1[323], out[803]);
  buf b_262_(set1[220], out[700]);
  buf b_263_(set2[172], out[172]);
  buf b_264_(set1[325], out[805]);
  buf b_265_(set1[472], out[952]);
  buf b_266_(set2[479], out[479]);
  buf b_267_(set2[258], out[258]);
  buf b_268_(set2[54], out[54]);
  buf b_269_(set2[263], out[263]);
  buf b_270_(set1[442], out[922]);
  buf b_271_(set1[474], out[954]);
  buf b_272_(set1[397], out[877]);
  buf b_273_(set1[134], out[614]);
  buf b_274_(set1[392], out[872]);
  buf b_275_(set2[98], out[98]);
  buf b_276_(set1[65], out[545]);
  buf b_277_(set1[399], out[879]);
  buf b_278_(set1[344], out[824]);
  buf b_279_(set1[231], out[711]);
  buf b_280_(set1[228], out[708]);
  buf b_281_(set2[402], out[402]);
  buf b_282_(set2[95], out[95]);
  buf b_283_(set1[416], out[896]);
  buf b_284_(set1[287], out[767]);
  buf b_285_(set1[196], out[676]);
  buf b_286_(set2[364], out[364]);
  buf b_287_(set2[192], out[192]);
  buf b_288_(set2[383], out[383]);
  buf b_289_(set1[152], out[632]);
  buf b_290_(set1[466], out[946]);
  buf b_291_(set2[132], out[132]);
  buf b_292_(set2[214], out[214]);
  buf b_293_(set2[371], out[371]);
  buf b_294_(set1[92], out[572]);
  buf b_295_(set1[69], out[549]);
  buf b_296_(set1[36], out[516]);
  buf b_297_(set1[242], out[722]);
  buf b_298_(set2[382], out[382]);
  buf b_299_(set1[352], out[832]);
  buf b_300_(set1[288], out[768]);
  buf b_301_(set1[305], out[785]);
  buf b_302_(set2[395], out[395]);
  buf b_303_(set2[318], out[318]);
  buf b_304_(set2[218], out[218]);
  buf b_305_(set1[400], out[880]);
  buf b_306_(set2[355], out[355]);
  buf b_307_(set1[192], out[672]);
  buf b_308_(set2[108], out[108]);
  buf b_309_(set2[107], out[107]);
  buf b_310_(set1[83], out[563]);
  buf b_311_(set1[271], out[751]);
  buf b_312_(set2[7], out[7]);
  buf b_313_(set1[239], out[719]);
  buf b_314_(set1[306], out[786]);
  buf b_315_(set1[359], out[839]);
  buf b_316_(set2[51], out[51]);
  buf b_317_(set2[303], out[303]);
  buf b_318_(set1[55], out[535]);
  buf b_319_(set1[281], out[761]);
  buf b_320_(set2[106], out[106]);
  buf b_321_(set2[5], out[5]);
  buf b_322_(set1[71], out[551]);
  buf b_323_(set1[398], out[878]);
  buf b_324_(set2[467], out[467]);
  buf b_325_(set2[444], out[444]);
  buf b_326_(set1[441], out[921]);
  buf b_327_(set2[317], out[317]);
  buf b_328_(set1[349], out[829]);
  buf b_329_(set1[319], out[799]);
  buf b_330_(set2[29], out[29]);
  buf b_331_(set2[282], out[282]);
  buf b_332_(set2[457], out[457]);
  buf b_333_(set2[293], out[293]);
  buf b_334_(set2[272], out[272]);
  buf b_335_(set1[184], out[664]);
  buf b_336_(set2[88], out[88]);
  buf b_337_(set1[452], out[932]);
  buf b_338_(set1[156], out[636]);
  buf b_339_(set1[136], out[616]);
  buf b_340_(set1[372], out[852]);
  buf b_341_(set1[194], out[674]);
  buf b_342_(set1[336], out[816]);
  buf b_343_(set2[473], out[473]);
  buf b_344_(set2[169], out[169]);
  buf b_345_(set2[149], out[149]);
  buf b_346_(set2[190], out[190]);
  buf b_347_(set1[430], out[910]);
  buf b_348_(set2[64], out[64]);
  buf b_349_(set1[124], out[604]);
  buf b_350_(set2[266], out[266]);
  buf b_351_(set2[87], out[87]);
  buf b_352_(set2[380], out[380]);
  buf b_353_(set2[80], out[80]);
  buf b_354_(set2[68], out[68]);
  buf b_355_(set2[31], out[31]);
  buf b_356_(set1[15], out[495]);
  buf b_357_(set1[185], out[665]);
  buf b_358_(set2[112], out[112]);
  buf b_359_(set2[298], out[298]);
  buf b_360_(set1[450], out[930]);
  buf b_361_(set1[357], out[837]);
  buf b_362_(set1[129], out[609]);
  buf b_363_(set2[186], out[186]);
  buf b_364_(set2[334], out[334]);
  buf b_365_(set1[280], out[760]);
  buf b_366_(set2[409], out[409]);
  buf b_367_(set1[164], out[644]);
  buf b_368_(set1[38], out[518]);
  buf b_369_(set1[451], out[931]);
  buf b_370_(set2[339], out[339]);
  buf b_371_(set2[274], out[274]);
  buf b_372_(set2[391], out[391]);
  buf b_373_(set1[365], out[845]);
  buf b_374_(set2[82], out[82]);
  buf b_375_(set1[279], out[759]);
  buf b_376_(set1[304], out[784]);
  buf b_377_(set2[204], out[204]);
  buf b_378_(set1[167], out[647]);
  buf b_379_(set1[414], out[894]);
  buf b_380_(set2[160], out[160]);
  buf b_381_(set2[294], out[294]);
  buf b_382_(set1[406], out[886]);
  buf b_383_(set1[145], out[625]);
  buf b_384_(set2[14], out[14]);
  buf b_385_(set2[185], out[185]);
  buf b_386_(set2[401], out[401]);
  buf b_387_(set1[265], out[745]);
  buf b_388_(set1[432], out[912]);
  buf b_389_(set2[15], out[15]);
  buf b_390_(set2[370], out[370]);
  buf b_391_(set2[273], out[273]);
  buf b_392_(set1[121], out[601]);
  buf b_393_(set2[259], out[259]);
  buf b_394_(set2[203], out[203]);
  buf b_395_(set1[81], out[561]);
  buf b_396_(set1[261], out[741]);
  buf b_397_(set1[66], out[546]);
  buf b_398_(set1[264], out[744]);
  buf b_399_(set1[202], out[682]);
  buf b_400_(set1[410], out[890]);
  buf b_401_(set2[207], out[207]);
  buf b_402_(set1[293], out[773]);
  buf b_403_(set1[199], out[679]);
  buf b_404_(set1[245], out[725]);
  buf b_405_(set2[394], out[394]);
  buf b_406_(set2[269], out[269]);
  buf b_407_(set1[282], out[762]);
  buf b_408_(set2[210], out[210]);
  buf b_409_(set2[439], out[439]);
  buf b_410_(set1[345], out[825]);
  buf b_411_(set2[388], out[388]);
  buf b_412_(set1[237], out[717]);
  buf b_413_(set2[99], out[99]);
  buf b_414_(set2[79], out[79]);
  buf b_415_(set2[84], out[84]);
  buf b_416_(set1[94], out[574]);
  buf b_417_(set1[470], out[950]);
  buf b_418_(set1[34], out[514]);
  buf b_419_(set1[139], out[619]);
  buf b_420_(set2[136], out[136]);
  buf b_421_(set2[189], out[189]);
  buf b_422_(set2[36], out[36]);
  buf b_423_(set1[96], out[576]);
  buf b_424_(set2[143], out[143]);
  buf b_425_(set2[360], out[360]);
  buf b_426_(set2[345], out[345]);
  buf b_427_(set1[166], out[646]);
  buf b_428_(set2[441], out[441]);
  buf b_429_(set1[203], out[683]);
  buf b_430_(set1[348], out[828]);
  buf b_431_(set2[423], out[423]);
  buf b_432_(set1[110], out[590]);
  buf b_433_(set1[351], out[831]);
  buf b_434_(set2[56], out[56]);
  buf b_435_(set2[180], out[180]);
  buf b_436_(set2[408], out[408]);
  buf b_437_(set1[226], out[706]);
  buf b_438_(set1[444], out[924]);
  buf b_439_(set1[445], out[925]);
  buf b_440_(set2[0], out[0]);
  buf b_441_(set1[283], out[763]);
  buf b_442_(set2[103], out[103]);
  buf b_443_(set2[50], out[50]);
  buf b_444_(set1[477], out[957]);
  buf b_445_(set2[399], out[399]);
  buf b_446_(set2[35], out[35]);
  buf b_447_(set2[448], out[448]);
  buf b_448_(set1[422], out[902]);
  buf b_449_(set1[138], out[618]);
  buf b_450_(set2[182], out[182]);
  buf b_451_(set2[6], out[6]);
  buf b_452_(set2[363], out[363]);
  buf b_453_(set1[403], out[883]);
  buf b_454_(set1[84], out[564]);
  buf b_455_(set2[26], out[26]);
  buf b_456_(set2[329], out[329]);
  buf b_457_(set2[94], out[94]);
  buf b_458_(set2[440], out[440]);
  buf b_459_(set2[134], out[134]);
  buf b_460_(set2[396], out[396]);
  buf b_461_(set1[122], out[602]);
  buf b_462_(set2[278], out[278]);
  buf b_463_(set2[209], out[209]);
  buf b_464_(set1[140], out[620]);
  buf b_465_(set1[9], out[489]);
  buf b_466_(set1[144], out[624]);
  buf b_467_(set2[59], out[59]);
  buf b_468_(set2[384], out[384]);
  buf b_469_(set2[428], out[428]);
  buf b_470_(set2[121], out[121]);
  buf b_471_(set2[461], out[461]);
  buf b_472_(set1[3], out[483]);
  buf b_473_(set1[298], out[778]);
  buf b_474_(set2[206], out[206]);
  buf b_475_(set2[455], out[455]);
  buf b_476_(set1[131], out[611]);
  buf b_477_(set2[37], out[37]);
  buf b_478_(set2[168], out[168]);
  buf b_479_(set2[130], out[130]);
  buf b_480_(set1[26], out[506]);
  buf b_481_(set2[264], out[264]);
  buf b_482_(set1[182], out[662]);
  buf b_483_(set2[291], out[291]);
  buf b_484_(set1[259], out[739]);
  buf b_485_(set2[431], out[431]);
  buf b_486_(set1[210], out[690]);
  buf b_487_(set1[255], out[735]);
  buf b_488_(set1[218], out[698]);
  buf b_489_(set2[332], out[332]);
  buf b_490_(set1[241], out[721]);
  buf b_491_(set1[148], out[628]);
  buf b_492_(set2[470], out[470]);
  buf b_493_(set1[20], out[500]);
  buf b_494_(set2[22], out[22]);
  buf b_495_(set1[70], out[550]);
  buf b_496_(set2[11], out[11]);
  buf b_497_(set1[339], out[819]);
  buf b_498_(set2[115], out[115]);
  buf b_499_(set1[5], out[485]);
  buf b_500_(set1[301], out[781]);
  buf b_501_(set1[163], out[643]);
  buf b_502_(set2[125], out[125]);
  buf b_503_(set1[127], out[607]);
  buf b_504_(set1[295], out[775]);
  buf b_505_(set2[234], out[234]);
  buf b_506_(set2[476], out[476]);
  buf b_507_(set1[133], out[613]);
  buf b_508_(set1[396], out[876]);
  buf b_509_(set1[42], out[522]);
  buf b_510_(set2[393], out[393]);
  buf b_511_(set1[104], out[584]);
  buf b_512_(set1[459], out[939]);
  buf b_513_(set1[21], out[501]);
  buf b_514_(set2[267], out[267]);
  buf b_515_(set1[289], out[769]);
  buf b_516_(set2[471], out[471]);
  buf b_517_(set2[122], out[122]);
  buf b_518_(set1[312], out[792]);
  buf b_519_(set1[407], out[887]);
  buf b_520_(set2[362], out[362]);
  buf b_521_(set2[74], out[74]);
  buf b_522_(set2[283], out[283]);
  buf b_523_(set2[101], out[101]);
  buf b_524_(set2[265], out[265]);
  buf b_525_(set1[99], out[579]);
  buf b_526_(set1[380], out[860]);
  buf b_527_(set1[308], out[788]);
  buf b_528_(set2[254], out[254]);
  buf b_529_(set2[67], out[67]);
  buf b_530_(set1[97], out[577]);
  buf b_531_(set1[30], out[510]);
  buf b_532_(set2[341], out[341]);
  buf b_533_(set2[415], out[415]);
  buf b_534_(set2[405], out[405]);
  buf b_535_(set2[114], out[114]);
  buf b_536_(set2[378], out[378]);
  buf b_537_(set1[143], out[623]);
  buf b_538_(set1[25], out[505]);
  buf b_539_(set2[126], out[126]);
  buf b_540_(set1[377], out[857]);
  buf b_541_(set1[236], out[716]);
  buf b_542_(set1[107], out[587]);
  buf b_543_(set2[435], out[435]);
  buf b_544_(set2[85], out[85]);
  buf b_545_(set2[93], out[93]);
  buf b_546_(set2[325], out[325]);
  buf b_547_(set2[286], out[286]);
  buf b_548_(set1[332], out[812]);
  buf b_549_(set1[183], out[663]);
  buf b_550_(set2[445], out[445]);
  buf b_551_(set2[83], out[83]);
  buf b_552_(set1[389], out[869]);
  buf b_553_(set1[438], out[918]);
  buf b_554_(set1[39], out[519]);
  buf b_555_(set2[16], out[16]);
  buf b_556_(set1[331], out[811]);
  buf b_557_(set2[433], out[433]);
  buf b_558_(set2[253], out[253]);
  buf b_559_(set1[189], out[669]);
  buf b_560_(set2[181], out[181]);
  buf b_561_(set2[167], out[167]);
  buf b_562_(set1[193], out[673]);
  buf b_563_(set2[70], out[70]);
  buf b_564_(set1[146], out[626]);
  buf b_565_(set2[346], out[346]);
  buf b_566_(set2[420], out[420]);
  buf b_567_(set2[261], out[261]);
  buf b_568_(set1[112], out[592]);
  buf b_569_(set2[224], out[224]);
  buf b_570_(set2[462], out[462]);
  buf b_571_(set2[188], out[188]);
  buf b_572_(set1[109], out[589]);
  buf b_573_(set1[162], out[642]);
  buf b_574_(set2[184], out[184]);
  buf b_575_(set1[6], out[486]);
  buf b_576_(set1[227], out[707]);
  buf b_577_(set2[387], out[387]);
  buf b_578_(set2[376], out[376]);
  buf b_579_(set2[250], out[250]);
  buf b_580_(set1[446], out[926]);
  buf b_581_(set1[330], out[810]);
  buf b_582_(set1[257], out[737]);
  buf b_583_(set2[348], out[348]);
  buf b_584_(set2[76], out[76]);
  buf b_585_(set2[331], out[331]);
  buf b_586_(set2[73], out[73]);
  buf b_587_(set1[307], out[787]);
  buf b_588_(set2[128], out[128]);
  buf b_589_(set2[343], out[343]);
  buf b_590_(set2[166], out[166]);
  buf b_591_(set2[449], out[449]);
  buf b_592_(set1[89], out[569]);
  buf b_593_(set2[368], out[368]);
  buf b_594_(set2[451], out[451]);
  buf b_595_(set1[175], out[655]);
  buf b_596_(set1[230], out[710]);
  buf b_597_(set2[320], out[320]);
  buf b_598_(set2[436], out[436]);
  buf b_599_(set1[384], out[864]);
  buf b_600_(set2[285], out[285]);
  buf b_601_(set2[418], out[418]);
  buf b_602_(set1[32], out[512]);
  buf b_603_(set2[152], out[152]);
  buf b_604_(set1[347], out[827]);
  buf b_605_(set1[46], out[526]);
  buf b_606_(set1[54], out[534]);
  buf b_607_(set2[17], out[17]);
  buf b_608_(set1[87], out[567]);
  buf b_609_(set1[88], out[568]);
  buf b_610_(set2[406], out[406]);
  buf b_611_(set1[174], out[654]);
  buf b_612_(set1[215], out[695]);
  buf b_613_(set1[296], out[776]);
  buf b_614_(set2[147], out[147]);
  buf b_615_(set2[358], out[358]);
  buf b_616_(set1[80], out[560]);
  buf b_617_(set1[256], out[736]);
  buf b_618_(set1[263], out[743]);
  buf b_619_(set1[219], out[699]);
  buf b_620_(set1[391], out[871]);
  buf b_621_(set1[375], out[855]);
  buf b_622_(set2[193], out[193]);
  buf b_623_(set1[225], out[705]);
  buf b_624_(set1[62], out[542]);
  buf b_625_(set1[79], out[559]);
  buf b_626_(set1[243], out[723]);
  buf b_627_(set2[47], out[47]);
  buf b_628_(set1[82], out[562]);
  buf b_629_(set2[215], out[215]);
  buf b_630_(set1[207], out[687]);
  buf b_631_(set2[44], out[44]);
  buf b_632_(set1[161], out[641]);
  buf b_633_(set1[354], out[834]);
  buf b_634_(set1[284], out[764]);
  buf b_635_(set2[42], out[42]);
  buf b_636_(set1[251], out[731]);
  buf b_637_(set1[23], out[503]);
  buf b_638_(set1[342], out[822]);
  buf b_639_(set1[478], out[958]);
  buf b_640_(set2[427], out[427]);
  buf b_641_(set1[10], out[490]);
  buf b_642_(set2[338], out[338]);
  buf b_643_(set1[238], out[718]);
  buf b_644_(set2[352], out[352]);
  buf b_645_(set2[55], out[55]);
  buf b_646_(set1[402], out[882]);
  buf b_647_(set2[326], out[326]);
  buf b_648_(set1[258], out[738]);
  buf b_649_(set1[418], out[898]);
  buf b_650_(set1[404], out[884]);
  buf b_651_(set2[277], out[277]);
  buf b_652_(set1[1], out[481]);
  buf b_653_(set1[160], out[640]);
  buf b_654_(set2[142], out[142]);
  buf b_655_(set2[243], out[243]);
  buf b_656_(set2[301], out[301]);
  buf b_657_(set1[311], out[791]);
  buf b_658_(set2[49], out[49]);
  buf b_659_(set2[397], out[397]);
  buf b_660_(set2[237], out[237]);
  buf b_661_(set2[308], out[308]);
  buf b_662_(set2[438], out[438]);
  buf b_663_(set2[295], out[295]);
  buf b_664_(set1[150], out[630]);
  buf b_665_(set1[411], out[891]);
  buf b_666_(set2[9], out[9]);
  buf b_667_(set2[220], out[220]);
  buf b_668_(set2[20], out[20]);
  buf b_669_(set1[128], out[608]);
  buf b_670_(set1[130], out[610]);
  buf b_671_(set1[382], out[862]);
  buf b_672_(set1[179], out[659]);
  buf b_673_(set1[16], out[496]);
  buf b_674_(set2[154], out[154]);
  buf b_675_(set1[132], out[612]);
  buf b_676_(set1[317], out[797]);
  buf b_677_(set1[262], out[742]);
  buf b_678_(set1[456], out[936]);
  buf b_679_(set2[328], out[328]);
  buf b_680_(set1[333], out[813]);
  buf b_681_(set2[270], out[270]);
  buf b_682_(set2[367], out[367]);
  buf b_683_(set2[201], out[201]);
  buf b_684_(set1[93], out[573]);
  buf b_685_(set2[63], out[63]);
  buf b_686_(set2[127], out[127]);
  buf b_687_(set2[58], out[58]);
  buf b_688_(set1[44], out[524]);
  buf b_689_(set2[248], out[248]);
  buf b_690_(set1[213], out[693]);
  buf b_691_(set2[52], out[52]);
  buf b_692_(set1[334], out[814]);
  buf b_693_(set1[316], out[796]);
  buf b_694_(set1[118], out[598]);
  buf b_695_(set2[150], out[150]);
  buf b_696_(set2[386], out[386]);
  buf b_697_(set2[300], out[300]);
  buf b_698_(set2[164], out[164]);
  buf b_699_(set2[8], out[8]);
  buf b_700_(set2[252], out[252]);
  buf b_701_(set1[53], out[533]);
  buf b_702_(set2[120], out[120]);
  buf b_703_(set2[255], out[255]);
  buf b_704_(set1[105], out[585]);
  buf b_705_(set2[369], out[369]);
  buf b_706_(set2[230], out[230]);
  buf b_707_(set1[272], out[752]);
  buf b_708_(set1[385], out[865]);
  buf b_709_(set1[448], out[928]);
  buf b_710_(set1[47], out[527]);
  buf b_711_(set1[290], out[770]);
  buf b_712_(set2[148], out[148]);
  buf b_713_(set1[155], out[635]);
  buf b_714_(set1[429], out[909]);
  buf b_715_(set1[467], out[947]);
  buf b_716_(set1[126], out[606]);
  buf b_717_(set1[463], out[943]);
  buf b_718_(set2[133], out[133]);
  buf b_719_(set1[462], out[942]);
  buf b_720_(set1[297], out[777]);
  buf b_721_(set2[116], out[116]);
  buf b_722_(set2[157], out[157]);
  buf b_723_(set1[412], out[892]);
  buf b_724_(set1[8], out[488]);
  buf b_725_(set1[188], out[668]);
  buf b_726_(set1[91], out[571]);
  buf b_727_(set1[165], out[645]);
  buf b_728_(set2[113], out[113]);
  buf b_729_(set1[461], out[941]);
  buf b_730_(set1[177], out[657]);
  buf b_731_(set2[314], out[314]);
  buf b_732_(set2[162], out[162]);
  buf b_733_(set1[51], out[531]);
  buf b_734_(set1[61], out[541]);
  buf b_735_(set2[398], out[398]);
  buf b_736_(set1[321], out[801]);
  buf b_737_(set2[65], out[65]);
  buf b_738_(set2[119], out[119]);
  buf b_739_(set2[463], out[463]);
  buf b_740_(set2[105], out[105]);
  buf b_741_(set2[327], out[327]);
  buf b_742_(set2[155], out[155]);
  buf b_743_(set2[46], out[46]);
  buf b_744_(set2[171], out[171]);
  buf b_745_(set1[86], out[566]);
  buf b_746_(set1[24], out[504]);
  buf b_747_(set2[176], out[176]);
  buf b_748_(set2[366], out[366]);
  buf b_749_(set1[222], out[702]);
  buf b_750_(set2[173], out[173]);
  buf b_751_(set1[211], out[691]);
  buf b_752_(set1[200], out[680]);
  buf b_753_(set1[285], out[765]);
  buf b_754_(set1[37], out[517]);
  buf b_755_(set1[72], out[552]);
  buf b_756_(set1[310], out[790]);
  buf b_757_(set2[424], out[424]);
  buf b_758_(set1[322], out[802]);
  buf b_759_(set1[338], out[818]);
  buf b_760_(set2[311], out[311]);
  buf b_761_(set1[294], out[774]);
  buf b_762_(set1[335], out[815]);
  buf b_763_(set2[72], out[72]);
  buf b_764_(set2[43], out[43]);
  buf b_765_(set1[455], out[935]);
  buf b_766_(set1[277], out[757]);
  buf b_767_(set1[314], out[794]);
  buf b_768_(set1[221], out[701]);
  buf b_769_(set2[219], out[219]);
  buf b_770_(set2[117], out[117]);
  buf b_771_(set2[458], out[458]);
  buf b_772_(set2[191], out[191]);
  buf b_773_(set2[245], out[245]);
  buf b_774_(set2[412], out[412]);
  buf b_775_(set2[226], out[226]);
  buf b_776_(set2[373], out[373]);
  buf b_777_(set1[363], out[843]);
  buf b_778_(set1[224], out[704]);
  buf b_779_(set2[194], out[194]);
  buf b_780_(set2[297], out[297]);
  buf b_781_(set2[213], out[213]);
  buf b_782_(set2[251], out[251]);
  buf b_783_(set2[97], out[97]);
  buf b_784_(set1[90], out[570]);
  buf b_785_(set1[326], out[806]);
  buf b_786_(set1[350], out[830]);
  buf b_787_(set2[32], out[32]);
  buf b_788_(set2[62], out[62]);
  buf b_789_(set1[379], out[859]);
  buf b_790_(set2[305], out[305]);
  buf b_791_(set1[435], out[915]);
  buf b_792_(set2[60], out[60]);
  buf b_793_(set2[2], out[2]);
  buf b_794_(set2[216], out[216]);
  buf b_795_(set2[221], out[221]);
  buf b_796_(set2[312], out[312]);
  buf b_797_(set1[137], out[617]);
  buf b_798_(set2[437], out[437]);
  buf b_799_(set2[333], out[333]);
  buf b_800_(set1[33], out[513]);
  buf b_801_(set1[370], out[850]);
  buf b_802_(set2[244], out[244]);
  buf b_803_(set2[200], out[200]);
  buf b_804_(set1[77], out[557]);
  buf b_805_(set2[211], out[211]);
  buf b_806_(set2[77], out[77]);
  buf b_807_(set2[292], out[292]);
  buf b_808_(set2[229], out[229]);
  buf b_809_(set2[330], out[330]);
  buf b_810_(set2[61], out[61]);
  buf b_811_(set2[109], out[109]);
  buf b_812_(set2[413], out[413]);
  buf b_813_(set2[240], out[240]);
  buf b_814_(set2[262], out[262]);
  buf b_815_(set1[67], out[547]);
  buf b_816_(set1[76], out[556]);
  buf b_817_(set2[89], out[89]);
  buf b_818_(set2[202], out[202]);
  buf b_819_(set2[247], out[247]);
  buf b_820_(set2[163], out[163]);
  buf b_821_(set2[156], out[156]);
  buf b_822_(set2[410], out[410]);
  buf b_823_(set2[275], out[275]);
  buf b_824_(set2[404], out[404]);
  buf b_825_(set1[78], out[558]);
  buf b_826_(set1[116], out[596]);
  buf b_827_(set1[186], out[666]);
  buf b_828_(set2[287], out[287]);
  buf b_829_(set1[337], out[817]);
  buf b_830_(set2[257], out[257]);
  buf b_831_(set1[181], out[661]);
  buf b_832_(set1[35], out[515]);
  buf b_833_(set1[387], out[867]);
  buf b_834_(set1[260], out[740]);
  buf b_835_(set1[158], out[638]);
  buf b_836_(set2[322], out[322]);
  buf b_837_(set2[13], out[13]);
  buf b_838_(set1[135], out[615]);
  buf b_839_(set2[302], out[302]);
  buf b_840_(set1[464], out[944]);
  buf b_841_(set2[129], out[129]);
  buf b_842_(set1[471], out[951]);
  buf b_843_(set2[198], out[198]);
  buf b_844_(set1[114], out[594]);
  buf b_845_(set2[260], out[260]);
  buf b_846_(set1[108], out[588]);
  buf b_847_(set2[309], out[309]);
  buf b_848_(set1[275], out[755]);
  buf b_849_(set1[362], out[842]);
  buf b_850_(set1[73], out[553]);
  buf b_851_(set2[239], out[239]);
  buf b_852_(set2[460], out[460]);
  buf b_853_(set1[421], out[901]);
  buf b_854_(set1[252], out[732]);
  buf b_855_(set2[313], out[313]);
  buf b_856_(set1[31], out[511]);
  buf b_857_(set1[436], out[916]);
  buf b_858_(set2[12], out[12]);
  buf b_859_(set1[113], out[593]);
  buf b_860_(set2[372], out[372]);
  buf b_861_(set2[419], out[419]);
  buf b_862_(set1[388], out[868]);
  buf b_863_(set1[278], out[758]);
  buf b_864_(set1[356], out[836]);
  buf b_865_(set1[68], out[548]);
  buf b_866_(set2[222], out[222]);
  buf b_867_(set1[318], out[798]);
  buf b_868_(set2[71], out[71]);
  buf b_869_(set1[309], out[789]);
  buf b_870_(set2[319], out[319]);
  buf b_871_(set1[439], out[919]);
  buf b_872_(set2[351], out[351]);
  buf b_873_(set2[238], out[238]);
  buf b_874_(set2[30], out[30]);
  buf b_875_(set1[56], out[536]);
  buf b_876_(set2[356], out[356]);
  buf b_877_(set1[141], out[621]);
  buf b_878_(set2[139], out[139]);
  buf b_879_(set2[256], out[256]);
  buf b_880_(set1[223], out[703]);
  buf b_881_(set1[341], out[821]);
  buf b_882_(set1[7], out[487]);
  buf b_883_(set1[253], out[733]);
  buf b_884_(set2[41], out[41]);
  buf b_885_(set2[452], out[452]);
  buf b_886_(set1[369], out[849]);
  buf b_887_(set2[69], out[69]);
  buf b_888_(set2[390], out[390]);
  buf b_889_(set1[187], out[667]);
  buf b_890_(set2[307], out[307]);
  buf b_891_(set1[428], out[908]);
  buf b_892_(set1[229], out[709]);
  buf b_893_(set1[276], out[756]);
  buf b_894_(set1[214], out[694]);
  buf b_895_(set1[17], out[497]);
  buf b_896_(set2[474], out[474]);
  buf b_897_(set1[102], out[582]);
  buf b_898_(set1[378], out[858]);
  buf b_899_(set1[457], out[937]);
  buf b_900_(set2[225], out[225]);
  buf b_901_(set2[361], out[361]);
  buf b_902_(set2[165], out[165]);
  buf b_903_(set1[373], out[853]);
  buf b_904_(set1[340], out[820]);
  buf b_905_(set1[440], out[920]);
  buf b_906_(set2[336], out[336]);
  buf b_907_(set1[58], out[538]);
  buf b_908_(set2[196], out[196]);
  buf b_909_(set1[475], out[955]);
  buf b_910_(set2[10], out[10]);
  buf b_911_(set2[227], out[227]);
  buf b_912_(set2[39], out[39]);
  buf b_913_(set2[249], out[249]);
  buf b_914_(set2[414], out[414]);
  buf b_915_(set1[11], out[491]);
  buf b_916_(set1[125], out[605]);
  buf b_917_(set2[379], out[379]);
  buf b_918_(set1[29], out[509]);
  buf b_919_(set1[244], out[724]);
  buf b_920_(set1[12], out[492]);
  buf b_921_(set2[57], out[57]);
  buf b_922_(set2[53], out[53]);
  buf b_923_(set1[170], out[650]);
  buf b_924_(set2[477], out[477]);
  buf b_925_(set1[159], out[639]);
  buf b_926_(set2[197], out[197]);
  buf b_927_(set2[321], out[321]);
  buf b_928_(set1[408], out[888]);
  buf b_929_(set2[28], out[28]);
  buf b_930_(set1[355], out[835]);
  buf b_931_(set1[468], out[948]);
  buf b_932_(set1[315], out[795]);
  buf b_933_(set1[0], out[480]);
  buf b_934_(set1[254], out[734]);
  buf b_935_(set1[151], out[631]);
  buf b_936_(set1[473], out[953]);
  buf b_937_(set2[464], out[464]);
  buf b_938_(set1[168], out[648]);
  buf b_939_(set2[205], out[205]);
  buf b_940_(set1[469], out[949]);
  buf b_941_(set1[274], out[754]);
  buf b_942_(set2[381], out[381]);
  buf b_943_(set2[466], out[466]);
  buf b_944_(set1[453], out[933]);
  buf b_945_(set1[64], out[544]);
  buf b_946_(set1[27], out[507]);
  buf b_947_(set2[144], out[144]);
  buf b_948_(set1[240], out[720]);
  buf b_949_(set2[365], out[365]);
  buf b_950_(set1[366], out[846]);
  buf b_951_(set2[276], out[276]);
  buf b_952_(set2[280], out[280]);
  buf b_953_(set1[247], out[727]);
  buf b_954_(set1[95], out[575]);
  buf b_955_(set2[21], out[21]);
  buf b_956_(set1[327], out[807]);
  buf b_957_(set1[60], out[540]);
  buf b_958_(set2[475], out[475]);
  buf b_959_(set2[434], out[434]);

endmodule
