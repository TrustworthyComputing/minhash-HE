module min_hash(
  input wire [3199:0] set1,
  input wire [3199:0] set2,
  output wire [6415:0] out
);
  wire [15:0] set1_unflattened[200];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  assign set1_unflattened[30] = set1[495:480];
  assign set1_unflattened[31] = set1[511:496];
  assign set1_unflattened[32] = set1[527:512];
  assign set1_unflattened[33] = set1[543:528];
  assign set1_unflattened[34] = set1[559:544];
  assign set1_unflattened[35] = set1[575:560];
  assign set1_unflattened[36] = set1[591:576];
  assign set1_unflattened[37] = set1[607:592];
  assign set1_unflattened[38] = set1[623:608];
  assign set1_unflattened[39] = set1[639:624];
  assign set1_unflattened[40] = set1[655:640];
  assign set1_unflattened[41] = set1[671:656];
  assign set1_unflattened[42] = set1[687:672];
  assign set1_unflattened[43] = set1[703:688];
  assign set1_unflattened[44] = set1[719:704];
  assign set1_unflattened[45] = set1[735:720];
  assign set1_unflattened[46] = set1[751:736];
  assign set1_unflattened[47] = set1[767:752];
  assign set1_unflattened[48] = set1[783:768];
  assign set1_unflattened[49] = set1[799:784];
  assign set1_unflattened[50] = set1[815:800];
  assign set1_unflattened[51] = set1[831:816];
  assign set1_unflattened[52] = set1[847:832];
  assign set1_unflattened[53] = set1[863:848];
  assign set1_unflattened[54] = set1[879:864];
  assign set1_unflattened[55] = set1[895:880];
  assign set1_unflattened[56] = set1[911:896];
  assign set1_unflattened[57] = set1[927:912];
  assign set1_unflattened[58] = set1[943:928];
  assign set1_unflattened[59] = set1[959:944];
  assign set1_unflattened[60] = set1[975:960];
  assign set1_unflattened[61] = set1[991:976];
  assign set1_unflattened[62] = set1[1007:992];
  assign set1_unflattened[63] = set1[1023:1008];
  assign set1_unflattened[64] = set1[1039:1024];
  assign set1_unflattened[65] = set1[1055:1040];
  assign set1_unflattened[66] = set1[1071:1056];
  assign set1_unflattened[67] = set1[1087:1072];
  assign set1_unflattened[68] = set1[1103:1088];
  assign set1_unflattened[69] = set1[1119:1104];
  assign set1_unflattened[70] = set1[1135:1120];
  assign set1_unflattened[71] = set1[1151:1136];
  assign set1_unflattened[72] = set1[1167:1152];
  assign set1_unflattened[73] = set1[1183:1168];
  assign set1_unflattened[74] = set1[1199:1184];
  assign set1_unflattened[75] = set1[1215:1200];
  assign set1_unflattened[76] = set1[1231:1216];
  assign set1_unflattened[77] = set1[1247:1232];
  assign set1_unflattened[78] = set1[1263:1248];
  assign set1_unflattened[79] = set1[1279:1264];
  assign set1_unflattened[80] = set1[1295:1280];
  assign set1_unflattened[81] = set1[1311:1296];
  assign set1_unflattened[82] = set1[1327:1312];
  assign set1_unflattened[83] = set1[1343:1328];
  assign set1_unflattened[84] = set1[1359:1344];
  assign set1_unflattened[85] = set1[1375:1360];
  assign set1_unflattened[86] = set1[1391:1376];
  assign set1_unflattened[87] = set1[1407:1392];
  assign set1_unflattened[88] = set1[1423:1408];
  assign set1_unflattened[89] = set1[1439:1424];
  assign set1_unflattened[90] = set1[1455:1440];
  assign set1_unflattened[91] = set1[1471:1456];
  assign set1_unflattened[92] = set1[1487:1472];
  assign set1_unflattened[93] = set1[1503:1488];
  assign set1_unflattened[94] = set1[1519:1504];
  assign set1_unflattened[95] = set1[1535:1520];
  assign set1_unflattened[96] = set1[1551:1536];
  assign set1_unflattened[97] = set1[1567:1552];
  assign set1_unflattened[98] = set1[1583:1568];
  assign set1_unflattened[99] = set1[1599:1584];
  assign set1_unflattened[100] = set1[1615:1600];
  assign set1_unflattened[101] = set1[1631:1616];
  assign set1_unflattened[102] = set1[1647:1632];
  assign set1_unflattened[103] = set1[1663:1648];
  assign set1_unflattened[104] = set1[1679:1664];
  assign set1_unflattened[105] = set1[1695:1680];
  assign set1_unflattened[106] = set1[1711:1696];
  assign set1_unflattened[107] = set1[1727:1712];
  assign set1_unflattened[108] = set1[1743:1728];
  assign set1_unflattened[109] = set1[1759:1744];
  assign set1_unflattened[110] = set1[1775:1760];
  assign set1_unflattened[111] = set1[1791:1776];
  assign set1_unflattened[112] = set1[1807:1792];
  assign set1_unflattened[113] = set1[1823:1808];
  assign set1_unflattened[114] = set1[1839:1824];
  assign set1_unflattened[115] = set1[1855:1840];
  assign set1_unflattened[116] = set1[1871:1856];
  assign set1_unflattened[117] = set1[1887:1872];
  assign set1_unflattened[118] = set1[1903:1888];
  assign set1_unflattened[119] = set1[1919:1904];
  assign set1_unflattened[120] = set1[1935:1920];
  assign set1_unflattened[121] = set1[1951:1936];
  assign set1_unflattened[122] = set1[1967:1952];
  assign set1_unflattened[123] = set1[1983:1968];
  assign set1_unflattened[124] = set1[1999:1984];
  assign set1_unflattened[125] = set1[2015:2000];
  assign set1_unflattened[126] = set1[2031:2016];
  assign set1_unflattened[127] = set1[2047:2032];
  assign set1_unflattened[128] = set1[2063:2048];
  assign set1_unflattened[129] = set1[2079:2064];
  assign set1_unflattened[130] = set1[2095:2080];
  assign set1_unflattened[131] = set1[2111:2096];
  assign set1_unflattened[132] = set1[2127:2112];
  assign set1_unflattened[133] = set1[2143:2128];
  assign set1_unflattened[134] = set1[2159:2144];
  assign set1_unflattened[135] = set1[2175:2160];
  assign set1_unflattened[136] = set1[2191:2176];
  assign set1_unflattened[137] = set1[2207:2192];
  assign set1_unflattened[138] = set1[2223:2208];
  assign set1_unflattened[139] = set1[2239:2224];
  assign set1_unflattened[140] = set1[2255:2240];
  assign set1_unflattened[141] = set1[2271:2256];
  assign set1_unflattened[142] = set1[2287:2272];
  assign set1_unflattened[143] = set1[2303:2288];
  assign set1_unflattened[144] = set1[2319:2304];
  assign set1_unflattened[145] = set1[2335:2320];
  assign set1_unflattened[146] = set1[2351:2336];
  assign set1_unflattened[147] = set1[2367:2352];
  assign set1_unflattened[148] = set1[2383:2368];
  assign set1_unflattened[149] = set1[2399:2384];
  assign set1_unflattened[150] = set1[2415:2400];
  assign set1_unflattened[151] = set1[2431:2416];
  assign set1_unflattened[152] = set1[2447:2432];
  assign set1_unflattened[153] = set1[2463:2448];
  assign set1_unflattened[154] = set1[2479:2464];
  assign set1_unflattened[155] = set1[2495:2480];
  assign set1_unflattened[156] = set1[2511:2496];
  assign set1_unflattened[157] = set1[2527:2512];
  assign set1_unflattened[158] = set1[2543:2528];
  assign set1_unflattened[159] = set1[2559:2544];
  assign set1_unflattened[160] = set1[2575:2560];
  assign set1_unflattened[161] = set1[2591:2576];
  assign set1_unflattened[162] = set1[2607:2592];
  assign set1_unflattened[163] = set1[2623:2608];
  assign set1_unflattened[164] = set1[2639:2624];
  assign set1_unflattened[165] = set1[2655:2640];
  assign set1_unflattened[166] = set1[2671:2656];
  assign set1_unflattened[167] = set1[2687:2672];
  assign set1_unflattened[168] = set1[2703:2688];
  assign set1_unflattened[169] = set1[2719:2704];
  assign set1_unflattened[170] = set1[2735:2720];
  assign set1_unflattened[171] = set1[2751:2736];
  assign set1_unflattened[172] = set1[2767:2752];
  assign set1_unflattened[173] = set1[2783:2768];
  assign set1_unflattened[174] = set1[2799:2784];
  assign set1_unflattened[175] = set1[2815:2800];
  assign set1_unflattened[176] = set1[2831:2816];
  assign set1_unflattened[177] = set1[2847:2832];
  assign set1_unflattened[178] = set1[2863:2848];
  assign set1_unflattened[179] = set1[2879:2864];
  assign set1_unflattened[180] = set1[2895:2880];
  assign set1_unflattened[181] = set1[2911:2896];
  assign set1_unflattened[182] = set1[2927:2912];
  assign set1_unflattened[183] = set1[2943:2928];
  assign set1_unflattened[184] = set1[2959:2944];
  assign set1_unflattened[185] = set1[2975:2960];
  assign set1_unflattened[186] = set1[2991:2976];
  assign set1_unflattened[187] = set1[3007:2992];
  assign set1_unflattened[188] = set1[3023:3008];
  assign set1_unflattened[189] = set1[3039:3024];
  assign set1_unflattened[190] = set1[3055:3040];
  assign set1_unflattened[191] = set1[3071:3056];
  assign set1_unflattened[192] = set1[3087:3072];
  assign set1_unflattened[193] = set1[3103:3088];
  assign set1_unflattened[194] = set1[3119:3104];
  assign set1_unflattened[195] = set1[3135:3120];
  assign set1_unflattened[196] = set1[3151:3136];
  assign set1_unflattened[197] = set1[3167:3152];
  assign set1_unflattened[198] = set1[3183:3168];
  assign set1_unflattened[199] = set1[3199:3184];
  wire [15:0] set2_unflattened[200];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  assign set2_unflattened[30] = set2[495:480];
  assign set2_unflattened[31] = set2[511:496];
  assign set2_unflattened[32] = set2[527:512];
  assign set2_unflattened[33] = set2[543:528];
  assign set2_unflattened[34] = set2[559:544];
  assign set2_unflattened[35] = set2[575:560];
  assign set2_unflattened[36] = set2[591:576];
  assign set2_unflattened[37] = set2[607:592];
  assign set2_unflattened[38] = set2[623:608];
  assign set2_unflattened[39] = set2[639:624];
  assign set2_unflattened[40] = set2[655:640];
  assign set2_unflattened[41] = set2[671:656];
  assign set2_unflattened[42] = set2[687:672];
  assign set2_unflattened[43] = set2[703:688];
  assign set2_unflattened[44] = set2[719:704];
  assign set2_unflattened[45] = set2[735:720];
  assign set2_unflattened[46] = set2[751:736];
  assign set2_unflattened[47] = set2[767:752];
  assign set2_unflattened[48] = set2[783:768];
  assign set2_unflattened[49] = set2[799:784];
  assign set2_unflattened[50] = set2[815:800];
  assign set2_unflattened[51] = set2[831:816];
  assign set2_unflattened[52] = set2[847:832];
  assign set2_unflattened[53] = set2[863:848];
  assign set2_unflattened[54] = set2[879:864];
  assign set2_unflattened[55] = set2[895:880];
  assign set2_unflattened[56] = set2[911:896];
  assign set2_unflattened[57] = set2[927:912];
  assign set2_unflattened[58] = set2[943:928];
  assign set2_unflattened[59] = set2[959:944];
  assign set2_unflattened[60] = set2[975:960];
  assign set2_unflattened[61] = set2[991:976];
  assign set2_unflattened[62] = set2[1007:992];
  assign set2_unflattened[63] = set2[1023:1008];
  assign set2_unflattened[64] = set2[1039:1024];
  assign set2_unflattened[65] = set2[1055:1040];
  assign set2_unflattened[66] = set2[1071:1056];
  assign set2_unflattened[67] = set2[1087:1072];
  assign set2_unflattened[68] = set2[1103:1088];
  assign set2_unflattened[69] = set2[1119:1104];
  assign set2_unflattened[70] = set2[1135:1120];
  assign set2_unflattened[71] = set2[1151:1136];
  assign set2_unflattened[72] = set2[1167:1152];
  assign set2_unflattened[73] = set2[1183:1168];
  assign set2_unflattened[74] = set2[1199:1184];
  assign set2_unflattened[75] = set2[1215:1200];
  assign set2_unflattened[76] = set2[1231:1216];
  assign set2_unflattened[77] = set2[1247:1232];
  assign set2_unflattened[78] = set2[1263:1248];
  assign set2_unflattened[79] = set2[1279:1264];
  assign set2_unflattened[80] = set2[1295:1280];
  assign set2_unflattened[81] = set2[1311:1296];
  assign set2_unflattened[82] = set2[1327:1312];
  assign set2_unflattened[83] = set2[1343:1328];
  assign set2_unflattened[84] = set2[1359:1344];
  assign set2_unflattened[85] = set2[1375:1360];
  assign set2_unflattened[86] = set2[1391:1376];
  assign set2_unflattened[87] = set2[1407:1392];
  assign set2_unflattened[88] = set2[1423:1408];
  assign set2_unflattened[89] = set2[1439:1424];
  assign set2_unflattened[90] = set2[1455:1440];
  assign set2_unflattened[91] = set2[1471:1456];
  assign set2_unflattened[92] = set2[1487:1472];
  assign set2_unflattened[93] = set2[1503:1488];
  assign set2_unflattened[94] = set2[1519:1504];
  assign set2_unflattened[95] = set2[1535:1520];
  assign set2_unflattened[96] = set2[1551:1536];
  assign set2_unflattened[97] = set2[1567:1552];
  assign set2_unflattened[98] = set2[1583:1568];
  assign set2_unflattened[99] = set2[1599:1584];
  assign set2_unflattened[100] = set2[1615:1600];
  assign set2_unflattened[101] = set2[1631:1616];
  assign set2_unflattened[102] = set2[1647:1632];
  assign set2_unflattened[103] = set2[1663:1648];
  assign set2_unflattened[104] = set2[1679:1664];
  assign set2_unflattened[105] = set2[1695:1680];
  assign set2_unflattened[106] = set2[1711:1696];
  assign set2_unflattened[107] = set2[1727:1712];
  assign set2_unflattened[108] = set2[1743:1728];
  assign set2_unflattened[109] = set2[1759:1744];
  assign set2_unflattened[110] = set2[1775:1760];
  assign set2_unflattened[111] = set2[1791:1776];
  assign set2_unflattened[112] = set2[1807:1792];
  assign set2_unflattened[113] = set2[1823:1808];
  assign set2_unflattened[114] = set2[1839:1824];
  assign set2_unflattened[115] = set2[1855:1840];
  assign set2_unflattened[116] = set2[1871:1856];
  assign set2_unflattened[117] = set2[1887:1872];
  assign set2_unflattened[118] = set2[1903:1888];
  assign set2_unflattened[119] = set2[1919:1904];
  assign set2_unflattened[120] = set2[1935:1920];
  assign set2_unflattened[121] = set2[1951:1936];
  assign set2_unflattened[122] = set2[1967:1952];
  assign set2_unflattened[123] = set2[1983:1968];
  assign set2_unflattened[124] = set2[1999:1984];
  assign set2_unflattened[125] = set2[2015:2000];
  assign set2_unflattened[126] = set2[2031:2016];
  assign set2_unflattened[127] = set2[2047:2032];
  assign set2_unflattened[128] = set2[2063:2048];
  assign set2_unflattened[129] = set2[2079:2064];
  assign set2_unflattened[130] = set2[2095:2080];
  assign set2_unflattened[131] = set2[2111:2096];
  assign set2_unflattened[132] = set2[2127:2112];
  assign set2_unflattened[133] = set2[2143:2128];
  assign set2_unflattened[134] = set2[2159:2144];
  assign set2_unflattened[135] = set2[2175:2160];
  assign set2_unflattened[136] = set2[2191:2176];
  assign set2_unflattened[137] = set2[2207:2192];
  assign set2_unflattened[138] = set2[2223:2208];
  assign set2_unflattened[139] = set2[2239:2224];
  assign set2_unflattened[140] = set2[2255:2240];
  assign set2_unflattened[141] = set2[2271:2256];
  assign set2_unflattened[142] = set2[2287:2272];
  assign set2_unflattened[143] = set2[2303:2288];
  assign set2_unflattened[144] = set2[2319:2304];
  assign set2_unflattened[145] = set2[2335:2320];
  assign set2_unflattened[146] = set2[2351:2336];
  assign set2_unflattened[147] = set2[2367:2352];
  assign set2_unflattened[148] = set2[2383:2368];
  assign set2_unflattened[149] = set2[2399:2384];
  assign set2_unflattened[150] = set2[2415:2400];
  assign set2_unflattened[151] = set2[2431:2416];
  assign set2_unflattened[152] = set2[2447:2432];
  assign set2_unflattened[153] = set2[2463:2448];
  assign set2_unflattened[154] = set2[2479:2464];
  assign set2_unflattened[155] = set2[2495:2480];
  assign set2_unflattened[156] = set2[2511:2496];
  assign set2_unflattened[157] = set2[2527:2512];
  assign set2_unflattened[158] = set2[2543:2528];
  assign set2_unflattened[159] = set2[2559:2544];
  assign set2_unflattened[160] = set2[2575:2560];
  assign set2_unflattened[161] = set2[2591:2576];
  assign set2_unflattened[162] = set2[2607:2592];
  assign set2_unflattened[163] = set2[2623:2608];
  assign set2_unflattened[164] = set2[2639:2624];
  assign set2_unflattened[165] = set2[2655:2640];
  assign set2_unflattened[166] = set2[2671:2656];
  assign set2_unflattened[167] = set2[2687:2672];
  assign set2_unflattened[168] = set2[2703:2688];
  assign set2_unflattened[169] = set2[2719:2704];
  assign set2_unflattened[170] = set2[2735:2720];
  assign set2_unflattened[171] = set2[2751:2736];
  assign set2_unflattened[172] = set2[2767:2752];
  assign set2_unflattened[173] = set2[2783:2768];
  assign set2_unflattened[174] = set2[2799:2784];
  assign set2_unflattened[175] = set2[2815:2800];
  assign set2_unflattened[176] = set2[2831:2816];
  assign set2_unflattened[177] = set2[2847:2832];
  assign set2_unflattened[178] = set2[2863:2848];
  assign set2_unflattened[179] = set2[2879:2864];
  assign set2_unflattened[180] = set2[2895:2880];
  assign set2_unflattened[181] = set2[2911:2896];
  assign set2_unflattened[182] = set2[2927:2912];
  assign set2_unflattened[183] = set2[2943:2928];
  assign set2_unflattened[184] = set2[2959:2944];
  assign set2_unflattened[185] = set2[2975:2960];
  assign set2_unflattened[186] = set2[2991:2976];
  assign set2_unflattened[187] = set2[3007:2992];
  assign set2_unflattened[188] = set2[3023:3008];
  assign set2_unflattened[189] = set2[3039:3024];
  assign set2_unflattened[190] = set2[3055:3040];
  assign set2_unflattened[191] = set2[3071:3056];
  assign set2_unflattened[192] = set2[3087:3072];
  assign set2_unflattened[193] = set2[3103:3088];
  assign set2_unflattened[194] = set2[3119:3104];
  assign set2_unflattened[195] = set2[3135:3120];
  assign set2_unflattened[196] = set2[3151:3136];
  assign set2_unflattened[197] = set2[3167:3152];
  assign set2_unflattened[198] = set2[3183:3168];
  assign set2_unflattened[199] = set2[3199:3184];
  wire [15:0] array_index_292858;
  wire [15:0] array_index_292859;
  wire [11:0] add_292866;
  wire [11:0] add_292869;
  wire [15:0] array_index_292874;
  wire [15:0] array_index_292877;
  wire [10:0] add_292881;
  wire [10:0] add_292884;
  wire [11:0] add_292900;
  wire [11:0] sel_292902;
  wire [11:0] add_292905;
  wire [11:0] sel_292907;
  wire [15:0] array_index_292922;
  wire [15:0] array_index_292925;
  wire [8:0] add_292929;
  wire [8:0] add_292932;
  wire [10:0] add_292935;
  wire [11:0] sel_292938;
  wire [10:0] add_292940;
  wire [11:0] sel_292943;
  wire [11:0] add_292960;
  wire [11:0] sel_292962;
  wire [11:0] add_292965;
  wire [11:0] sel_292967;
  wire [15:0] array_index_292988;
  wire [15:0] array_index_292991;
  wire [10:0] add_292995;
  wire [10:0] add_292997;
  wire [8:0] add_292999;
  wire [11:0] sel_293002;
  wire [8:0] add_293004;
  wire [11:0] sel_293007;
  wire [10:0] add_293009;
  wire [11:0] sel_293012;
  wire [10:0] add_293014;
  wire [11:0] sel_293017;
  wire [11:0] add_293038;
  wire [11:0] sel_293040;
  wire [11:0] add_293043;
  wire [11:0] sel_293045;
  wire [15:0] array_index_293072;
  wire [15:0] array_index_293075;
  wire [10:0] add_293079;
  wire [10:0] add_293081;
  wire [10:0] add_293083;
  wire [11:0] sel_293085;
  wire [10:0] add_293087;
  wire [11:0] sel_293089;
  wire [8:0] add_293091;
  wire [11:0] sel_293094;
  wire [8:0] add_293096;
  wire [11:0] sel_293099;
  wire [10:0] add_293101;
  wire [11:0] sel_293104;
  wire [10:0] add_293106;
  wire [11:0] sel_293109;
  wire [11:0] add_293134;
  wire [11:0] sel_293136;
  wire [11:0] add_293139;
  wire [11:0] sel_293141;
  wire [15:0] array_index_293172;
  wire [15:0] array_index_293175;
  wire [10:0] add_293179;
  wire [11:0] sel_293181;
  wire [10:0] add_293183;
  wire [11:0] sel_293185;
  wire [10:0] add_293187;
  wire [11:0] sel_293189;
  wire [10:0] add_293191;
  wire [11:0] sel_293193;
  wire [8:0] add_293195;
  wire [11:0] sel_293198;
  wire [8:0] add_293200;
  wire [11:0] sel_293203;
  wire [10:0] add_293205;
  wire [11:0] sel_293208;
  wire [10:0] add_293210;
  wire [11:0] sel_293213;
  wire [11:0] add_293238;
  wire [11:0] sel_293240;
  wire [11:0] add_293243;
  wire [11:0] sel_293245;
  wire [15:0] array_index_293274;
  wire [15:0] array_index_293277;
  wire [10:0] add_293281;
  wire [11:0] sel_293283;
  wire [10:0] add_293285;
  wire [11:0] sel_293287;
  wire [10:0] add_293289;
  wire [11:0] sel_293291;
  wire [10:0] add_293293;
  wire [11:0] sel_293295;
  wire [8:0] add_293297;
  wire [11:0] sel_293300;
  wire [8:0] add_293302;
  wire [11:0] sel_293305;
  wire [10:0] add_293307;
  wire [11:0] sel_293310;
  wire [10:0] add_293312;
  wire [11:0] sel_293315;
  wire [11:0] add_293340;
  wire [11:0] sel_293342;
  wire [11:0] add_293345;
  wire [11:0] sel_293347;
  wire [15:0] array_index_293376;
  wire [15:0] array_index_293379;
  wire [10:0] add_293383;
  wire [11:0] sel_293385;
  wire [10:0] add_293387;
  wire [11:0] sel_293389;
  wire [10:0] add_293391;
  wire [11:0] sel_293393;
  wire [10:0] add_293395;
  wire [11:0] sel_293397;
  wire [8:0] add_293399;
  wire [11:0] sel_293402;
  wire [8:0] add_293404;
  wire [11:0] sel_293407;
  wire [10:0] add_293409;
  wire [11:0] sel_293412;
  wire [10:0] add_293414;
  wire [11:0] sel_293417;
  wire [11:0] add_293442;
  wire [11:0] sel_293444;
  wire [11:0] add_293447;
  wire [11:0] sel_293449;
  wire [15:0] array_index_293478;
  wire [15:0] array_index_293481;
  wire [10:0] add_293485;
  wire [11:0] sel_293487;
  wire [10:0] add_293489;
  wire [11:0] sel_293491;
  wire [10:0] add_293493;
  wire [11:0] sel_293495;
  wire [10:0] add_293497;
  wire [11:0] sel_293499;
  wire [8:0] add_293501;
  wire [11:0] sel_293504;
  wire [8:0] add_293506;
  wire [11:0] sel_293509;
  wire [10:0] add_293511;
  wire [11:0] sel_293514;
  wire [10:0] add_293516;
  wire [11:0] sel_293519;
  wire [11:0] add_293544;
  wire [11:0] sel_293546;
  wire [11:0] add_293549;
  wire [11:0] sel_293551;
  wire [15:0] array_index_293580;
  wire [15:0] array_index_293583;
  wire [10:0] add_293587;
  wire [11:0] sel_293589;
  wire [10:0] add_293591;
  wire [11:0] sel_293593;
  wire [10:0] add_293595;
  wire [11:0] sel_293597;
  wire [10:0] add_293599;
  wire [11:0] sel_293601;
  wire [8:0] add_293603;
  wire [11:0] sel_293606;
  wire [8:0] add_293608;
  wire [11:0] sel_293611;
  wire [10:0] add_293613;
  wire [11:0] sel_293616;
  wire [10:0] add_293618;
  wire [11:0] sel_293621;
  wire [11:0] add_293646;
  wire [11:0] sel_293648;
  wire [11:0] add_293651;
  wire [11:0] sel_293653;
  wire [15:0] array_index_293682;
  wire [15:0] array_index_293685;
  wire [10:0] add_293689;
  wire [11:0] sel_293691;
  wire [10:0] add_293693;
  wire [11:0] sel_293695;
  wire [10:0] add_293697;
  wire [11:0] sel_293699;
  wire [10:0] add_293701;
  wire [11:0] sel_293703;
  wire [8:0] add_293705;
  wire [11:0] sel_293708;
  wire [8:0] add_293710;
  wire [11:0] sel_293713;
  wire [10:0] add_293715;
  wire [11:0] sel_293718;
  wire [10:0] add_293720;
  wire [11:0] sel_293723;
  wire [11:0] add_293748;
  wire [11:0] sel_293750;
  wire [11:0] add_293753;
  wire [11:0] sel_293755;
  wire [15:0] array_index_293784;
  wire [15:0] array_index_293787;
  wire [10:0] add_293791;
  wire [11:0] sel_293793;
  wire [10:0] add_293795;
  wire [11:0] sel_293797;
  wire [10:0] add_293799;
  wire [11:0] sel_293801;
  wire [10:0] add_293803;
  wire [11:0] sel_293805;
  wire [8:0] add_293807;
  wire [11:0] sel_293810;
  wire [8:0] add_293812;
  wire [11:0] sel_293815;
  wire [10:0] add_293817;
  wire [11:0] sel_293820;
  wire [10:0] add_293822;
  wire [11:0] sel_293825;
  wire [11:0] add_293850;
  wire [11:0] sel_293852;
  wire [11:0] add_293855;
  wire [11:0] sel_293857;
  wire [15:0] array_index_293886;
  wire [15:0] array_index_293889;
  wire [10:0] add_293893;
  wire [11:0] sel_293895;
  wire [10:0] add_293897;
  wire [11:0] sel_293899;
  wire [10:0] add_293901;
  wire [11:0] sel_293903;
  wire [10:0] add_293905;
  wire [11:0] sel_293907;
  wire [8:0] add_293909;
  wire [11:0] sel_293912;
  wire [8:0] add_293914;
  wire [11:0] sel_293917;
  wire [10:0] add_293919;
  wire [11:0] sel_293922;
  wire [10:0] add_293924;
  wire [11:0] sel_293927;
  wire [11:0] add_293952;
  wire [11:0] sel_293954;
  wire [11:0] add_293957;
  wire [11:0] sel_293959;
  wire [15:0] array_index_293988;
  wire [15:0] array_index_293991;
  wire [10:0] add_293995;
  wire [11:0] sel_293997;
  wire [10:0] add_293999;
  wire [11:0] sel_294001;
  wire [10:0] add_294003;
  wire [11:0] sel_294005;
  wire [10:0] add_294007;
  wire [11:0] sel_294009;
  wire [8:0] add_294011;
  wire [11:0] sel_294014;
  wire [8:0] add_294016;
  wire [11:0] sel_294019;
  wire [10:0] add_294021;
  wire [11:0] sel_294024;
  wire [10:0] add_294026;
  wire [11:0] sel_294029;
  wire [11:0] add_294054;
  wire [11:0] sel_294056;
  wire [11:0] add_294059;
  wire [11:0] sel_294061;
  wire [15:0] array_index_294090;
  wire [15:0] array_index_294093;
  wire [10:0] add_294097;
  wire [11:0] sel_294099;
  wire [10:0] add_294101;
  wire [11:0] sel_294103;
  wire [10:0] add_294105;
  wire [11:0] sel_294107;
  wire [10:0] add_294109;
  wire [11:0] sel_294111;
  wire [8:0] add_294113;
  wire [11:0] sel_294116;
  wire [8:0] add_294118;
  wire [11:0] sel_294121;
  wire [10:0] add_294123;
  wire [11:0] sel_294126;
  wire [10:0] add_294128;
  wire [11:0] sel_294131;
  wire [11:0] add_294156;
  wire [11:0] sel_294158;
  wire [11:0] add_294161;
  wire [11:0] sel_294163;
  wire [15:0] array_index_294192;
  wire [15:0] array_index_294195;
  wire [10:0] add_294199;
  wire [11:0] sel_294201;
  wire [10:0] add_294203;
  wire [11:0] sel_294205;
  wire [10:0] add_294207;
  wire [11:0] sel_294209;
  wire [10:0] add_294211;
  wire [11:0] sel_294213;
  wire [8:0] add_294215;
  wire [11:0] sel_294218;
  wire [8:0] add_294220;
  wire [11:0] sel_294223;
  wire [10:0] add_294225;
  wire [11:0] sel_294228;
  wire [10:0] add_294230;
  wire [11:0] sel_294233;
  wire [11:0] add_294258;
  wire [11:0] sel_294260;
  wire [11:0] add_294263;
  wire [11:0] sel_294265;
  wire [15:0] array_index_294294;
  wire [15:0] array_index_294297;
  wire [10:0] add_294301;
  wire [11:0] sel_294303;
  wire [10:0] add_294305;
  wire [11:0] sel_294307;
  wire [10:0] add_294309;
  wire [11:0] sel_294311;
  wire [10:0] add_294313;
  wire [11:0] sel_294315;
  wire [8:0] add_294317;
  wire [11:0] sel_294320;
  wire [8:0] add_294322;
  wire [11:0] sel_294325;
  wire [10:0] add_294327;
  wire [11:0] sel_294330;
  wire [10:0] add_294332;
  wire [11:0] sel_294335;
  wire [11:0] add_294360;
  wire [11:0] sel_294362;
  wire [11:0] add_294365;
  wire [11:0] sel_294367;
  wire [15:0] array_index_294396;
  wire [15:0] array_index_294399;
  wire [10:0] add_294403;
  wire [11:0] sel_294405;
  wire [10:0] add_294407;
  wire [11:0] sel_294409;
  wire [10:0] add_294411;
  wire [11:0] sel_294413;
  wire [10:0] add_294415;
  wire [11:0] sel_294417;
  wire [8:0] add_294419;
  wire [11:0] sel_294422;
  wire [8:0] add_294424;
  wire [11:0] sel_294427;
  wire [10:0] add_294429;
  wire [11:0] sel_294432;
  wire [10:0] add_294434;
  wire [11:0] sel_294437;
  wire [11:0] add_294462;
  wire [11:0] sel_294464;
  wire [11:0] add_294467;
  wire [11:0] sel_294469;
  wire [15:0] array_index_294498;
  wire [15:0] array_index_294501;
  wire [10:0] add_294505;
  wire [11:0] sel_294507;
  wire [10:0] add_294509;
  wire [11:0] sel_294511;
  wire [10:0] add_294513;
  wire [11:0] sel_294515;
  wire [10:0] add_294517;
  wire [11:0] sel_294519;
  wire [8:0] add_294521;
  wire [11:0] sel_294524;
  wire [8:0] add_294526;
  wire [11:0] sel_294529;
  wire [10:0] add_294531;
  wire [11:0] sel_294534;
  wire [10:0] add_294536;
  wire [11:0] sel_294539;
  wire [11:0] add_294564;
  wire [11:0] sel_294566;
  wire [11:0] add_294569;
  wire [11:0] sel_294571;
  wire [15:0] array_index_294600;
  wire [15:0] array_index_294603;
  wire [10:0] add_294607;
  wire [11:0] sel_294609;
  wire [10:0] add_294611;
  wire [11:0] sel_294613;
  wire [10:0] add_294615;
  wire [11:0] sel_294617;
  wire [10:0] add_294619;
  wire [11:0] sel_294621;
  wire [8:0] add_294623;
  wire [11:0] sel_294626;
  wire [8:0] add_294628;
  wire [11:0] sel_294631;
  wire [10:0] add_294633;
  wire [11:0] sel_294636;
  wire [10:0] add_294638;
  wire [11:0] sel_294641;
  wire [11:0] add_294666;
  wire [11:0] sel_294668;
  wire [11:0] add_294671;
  wire [11:0] sel_294673;
  wire [15:0] array_index_294702;
  wire [15:0] array_index_294705;
  wire [10:0] add_294709;
  wire [11:0] sel_294711;
  wire [10:0] add_294713;
  wire [11:0] sel_294715;
  wire [10:0] add_294717;
  wire [11:0] sel_294719;
  wire [10:0] add_294721;
  wire [11:0] sel_294723;
  wire [8:0] add_294725;
  wire [11:0] sel_294728;
  wire [8:0] add_294730;
  wire [11:0] sel_294733;
  wire [10:0] add_294735;
  wire [11:0] sel_294738;
  wire [10:0] add_294740;
  wire [11:0] sel_294743;
  wire [11:0] add_294768;
  wire [11:0] sel_294770;
  wire [11:0] add_294773;
  wire [11:0] sel_294775;
  wire [15:0] array_index_294804;
  wire [15:0] array_index_294807;
  wire [10:0] add_294811;
  wire [11:0] sel_294813;
  wire [10:0] add_294815;
  wire [11:0] sel_294817;
  wire [10:0] add_294819;
  wire [11:0] sel_294821;
  wire [10:0] add_294823;
  wire [11:0] sel_294825;
  wire [8:0] add_294827;
  wire [11:0] sel_294830;
  wire [8:0] add_294832;
  wire [11:0] sel_294835;
  wire [10:0] add_294837;
  wire [11:0] sel_294840;
  wire [10:0] add_294842;
  wire [11:0] sel_294845;
  wire [11:0] add_294870;
  wire [11:0] sel_294872;
  wire [11:0] add_294875;
  wire [11:0] sel_294877;
  wire [15:0] array_index_294906;
  wire [15:0] array_index_294909;
  wire [10:0] add_294913;
  wire [11:0] sel_294915;
  wire [10:0] add_294917;
  wire [11:0] sel_294919;
  wire [10:0] add_294921;
  wire [11:0] sel_294923;
  wire [10:0] add_294925;
  wire [11:0] sel_294927;
  wire [8:0] add_294929;
  wire [11:0] sel_294932;
  wire [8:0] add_294934;
  wire [11:0] sel_294937;
  wire [10:0] add_294939;
  wire [11:0] sel_294942;
  wire [10:0] add_294944;
  wire [11:0] sel_294947;
  wire [11:0] add_294972;
  wire [11:0] sel_294974;
  wire [11:0] add_294977;
  wire [11:0] sel_294979;
  wire [15:0] array_index_295008;
  wire [15:0] array_index_295011;
  wire [10:0] add_295015;
  wire [11:0] sel_295017;
  wire [10:0] add_295019;
  wire [11:0] sel_295021;
  wire [10:0] add_295023;
  wire [11:0] sel_295025;
  wire [10:0] add_295027;
  wire [11:0] sel_295029;
  wire [8:0] add_295031;
  wire [11:0] sel_295034;
  wire [8:0] add_295036;
  wire [11:0] sel_295039;
  wire [10:0] add_295041;
  wire [11:0] sel_295044;
  wire [10:0] add_295046;
  wire [11:0] sel_295049;
  wire [11:0] add_295074;
  wire [11:0] sel_295076;
  wire [11:0] add_295079;
  wire [11:0] sel_295081;
  wire [15:0] array_index_295110;
  wire [15:0] array_index_295113;
  wire [10:0] add_295117;
  wire [11:0] sel_295119;
  wire [10:0] add_295121;
  wire [11:0] sel_295123;
  wire [10:0] add_295125;
  wire [11:0] sel_295127;
  wire [10:0] add_295129;
  wire [11:0] sel_295131;
  wire [8:0] add_295133;
  wire [11:0] sel_295136;
  wire [8:0] add_295138;
  wire [11:0] sel_295141;
  wire [10:0] add_295143;
  wire [11:0] sel_295146;
  wire [10:0] add_295148;
  wire [11:0] sel_295151;
  wire [11:0] add_295176;
  wire [11:0] sel_295178;
  wire [11:0] add_295181;
  wire [11:0] sel_295183;
  wire [15:0] array_index_295212;
  wire [15:0] array_index_295215;
  wire [10:0] add_295219;
  wire [11:0] sel_295221;
  wire [10:0] add_295223;
  wire [11:0] sel_295225;
  wire [10:0] add_295227;
  wire [11:0] sel_295229;
  wire [10:0] add_295231;
  wire [11:0] sel_295233;
  wire [8:0] add_295235;
  wire [11:0] sel_295238;
  wire [8:0] add_295240;
  wire [11:0] sel_295243;
  wire [10:0] add_295245;
  wire [11:0] sel_295248;
  wire [10:0] add_295250;
  wire [11:0] sel_295253;
  wire [11:0] add_295278;
  wire [11:0] sel_295280;
  wire [11:0] add_295283;
  wire [11:0] sel_295285;
  wire [15:0] array_index_295314;
  wire [15:0] array_index_295317;
  wire [10:0] add_295321;
  wire [11:0] sel_295323;
  wire [10:0] add_295325;
  wire [11:0] sel_295327;
  wire [10:0] add_295329;
  wire [11:0] sel_295331;
  wire [10:0] add_295333;
  wire [11:0] sel_295335;
  wire [8:0] add_295337;
  wire [11:0] sel_295340;
  wire [8:0] add_295342;
  wire [11:0] sel_295345;
  wire [10:0] add_295347;
  wire [11:0] sel_295350;
  wire [10:0] add_295352;
  wire [11:0] sel_295355;
  wire [11:0] add_295380;
  wire [11:0] sel_295382;
  wire [11:0] add_295385;
  wire [11:0] sel_295387;
  wire [15:0] array_index_295416;
  wire [15:0] array_index_295419;
  wire [10:0] add_295423;
  wire [11:0] sel_295425;
  wire [10:0] add_295427;
  wire [11:0] sel_295429;
  wire [10:0] add_295431;
  wire [11:0] sel_295433;
  wire [10:0] add_295435;
  wire [11:0] sel_295437;
  wire [8:0] add_295439;
  wire [11:0] sel_295442;
  wire [8:0] add_295444;
  wire [11:0] sel_295447;
  wire [10:0] add_295449;
  wire [11:0] sel_295452;
  wire [10:0] add_295454;
  wire [11:0] sel_295457;
  wire [11:0] add_295482;
  wire [11:0] sel_295484;
  wire [11:0] add_295487;
  wire [11:0] sel_295489;
  wire [15:0] array_index_295518;
  wire [15:0] array_index_295521;
  wire [10:0] add_295525;
  wire [11:0] sel_295527;
  wire [10:0] add_295529;
  wire [11:0] sel_295531;
  wire [10:0] add_295533;
  wire [11:0] sel_295535;
  wire [10:0] add_295537;
  wire [11:0] sel_295539;
  wire [8:0] add_295541;
  wire [11:0] sel_295544;
  wire [8:0] add_295546;
  wire [11:0] sel_295549;
  wire [10:0] add_295551;
  wire [11:0] sel_295554;
  wire [10:0] add_295556;
  wire [11:0] sel_295559;
  wire [11:0] add_295584;
  wire [11:0] sel_295586;
  wire [11:0] add_295589;
  wire [11:0] sel_295591;
  wire [15:0] array_index_295620;
  wire [15:0] array_index_295623;
  wire [10:0] add_295627;
  wire [11:0] sel_295629;
  wire [10:0] add_295631;
  wire [11:0] sel_295633;
  wire [10:0] add_295635;
  wire [11:0] sel_295637;
  wire [10:0] add_295639;
  wire [11:0] sel_295641;
  wire [8:0] add_295643;
  wire [11:0] sel_295646;
  wire [8:0] add_295648;
  wire [11:0] sel_295651;
  wire [10:0] add_295653;
  wire [11:0] sel_295656;
  wire [10:0] add_295658;
  wire [11:0] sel_295661;
  wire [11:0] add_295686;
  wire [11:0] sel_295688;
  wire [11:0] add_295691;
  wire [11:0] sel_295693;
  wire [15:0] array_index_295722;
  wire [15:0] array_index_295725;
  wire [10:0] add_295729;
  wire [11:0] sel_295731;
  wire [10:0] add_295733;
  wire [11:0] sel_295735;
  wire [10:0] add_295737;
  wire [11:0] sel_295739;
  wire [10:0] add_295741;
  wire [11:0] sel_295743;
  wire [8:0] add_295745;
  wire [11:0] sel_295748;
  wire [8:0] add_295750;
  wire [11:0] sel_295753;
  wire [10:0] add_295755;
  wire [11:0] sel_295758;
  wire [10:0] add_295760;
  wire [11:0] sel_295763;
  wire [11:0] add_295788;
  wire [11:0] sel_295790;
  wire [11:0] add_295793;
  wire [11:0] sel_295795;
  wire [15:0] array_index_295824;
  wire [15:0] array_index_295827;
  wire [10:0] add_295831;
  wire [11:0] sel_295833;
  wire [10:0] add_295835;
  wire [11:0] sel_295837;
  wire [10:0] add_295839;
  wire [11:0] sel_295841;
  wire [10:0] add_295843;
  wire [11:0] sel_295845;
  wire [8:0] add_295847;
  wire [11:0] sel_295850;
  wire [8:0] add_295852;
  wire [11:0] sel_295855;
  wire [10:0] add_295857;
  wire [11:0] sel_295860;
  wire [10:0] add_295862;
  wire [11:0] sel_295865;
  wire [11:0] add_295890;
  wire [11:0] sel_295892;
  wire [11:0] add_295895;
  wire [11:0] sel_295897;
  wire [15:0] array_index_295926;
  wire [15:0] array_index_295929;
  wire [10:0] add_295933;
  wire [11:0] sel_295935;
  wire [10:0] add_295937;
  wire [11:0] sel_295939;
  wire [10:0] add_295941;
  wire [11:0] sel_295943;
  wire [10:0] add_295945;
  wire [11:0] sel_295947;
  wire [8:0] add_295949;
  wire [11:0] sel_295952;
  wire [8:0] add_295954;
  wire [11:0] sel_295957;
  wire [10:0] add_295959;
  wire [11:0] sel_295962;
  wire [10:0] add_295964;
  wire [11:0] sel_295967;
  wire [11:0] add_295992;
  wire [11:0] sel_295994;
  wire [11:0] add_295997;
  wire [11:0] sel_295999;
  wire [15:0] array_index_296028;
  wire [15:0] array_index_296031;
  wire [10:0] add_296035;
  wire [11:0] sel_296037;
  wire [10:0] add_296039;
  wire [11:0] sel_296041;
  wire [10:0] add_296043;
  wire [11:0] sel_296045;
  wire [10:0] add_296047;
  wire [11:0] sel_296049;
  wire [8:0] add_296051;
  wire [11:0] sel_296054;
  wire [8:0] add_296056;
  wire [11:0] sel_296059;
  wire [10:0] add_296061;
  wire [11:0] sel_296064;
  wire [10:0] add_296066;
  wire [11:0] sel_296069;
  wire [11:0] add_296094;
  wire [11:0] sel_296096;
  wire [11:0] add_296099;
  wire [11:0] sel_296101;
  wire [15:0] array_index_296130;
  wire [15:0] array_index_296133;
  wire [10:0] add_296137;
  wire [11:0] sel_296139;
  wire [10:0] add_296141;
  wire [11:0] sel_296143;
  wire [10:0] add_296145;
  wire [11:0] sel_296147;
  wire [10:0] add_296149;
  wire [11:0] sel_296151;
  wire [8:0] add_296153;
  wire [11:0] sel_296156;
  wire [8:0] add_296158;
  wire [11:0] sel_296161;
  wire [10:0] add_296163;
  wire [11:0] sel_296166;
  wire [10:0] add_296168;
  wire [11:0] sel_296171;
  wire [11:0] add_296196;
  wire [11:0] sel_296198;
  wire [11:0] add_296201;
  wire [11:0] sel_296203;
  wire [15:0] array_index_296232;
  wire [15:0] array_index_296235;
  wire [10:0] add_296239;
  wire [11:0] sel_296241;
  wire [10:0] add_296243;
  wire [11:0] sel_296245;
  wire [10:0] add_296247;
  wire [11:0] sel_296249;
  wire [10:0] add_296251;
  wire [11:0] sel_296253;
  wire [8:0] add_296255;
  wire [11:0] sel_296258;
  wire [8:0] add_296260;
  wire [11:0] sel_296263;
  wire [10:0] add_296265;
  wire [11:0] sel_296268;
  wire [10:0] add_296270;
  wire [11:0] sel_296273;
  wire [11:0] add_296298;
  wire [11:0] sel_296300;
  wire [11:0] add_296303;
  wire [11:0] sel_296305;
  wire [15:0] array_index_296334;
  wire [15:0] array_index_296337;
  wire [10:0] add_296341;
  wire [11:0] sel_296343;
  wire [10:0] add_296345;
  wire [11:0] sel_296347;
  wire [10:0] add_296349;
  wire [11:0] sel_296351;
  wire [10:0] add_296353;
  wire [11:0] sel_296355;
  wire [8:0] add_296357;
  wire [11:0] sel_296360;
  wire [8:0] add_296362;
  wire [11:0] sel_296365;
  wire [10:0] add_296367;
  wire [11:0] sel_296370;
  wire [10:0] add_296372;
  wire [11:0] sel_296375;
  wire [11:0] add_296400;
  wire [11:0] sel_296402;
  wire [11:0] add_296405;
  wire [11:0] sel_296407;
  wire [15:0] array_index_296436;
  wire [15:0] array_index_296439;
  wire [10:0] add_296443;
  wire [11:0] sel_296445;
  wire [10:0] add_296447;
  wire [11:0] sel_296449;
  wire [10:0] add_296451;
  wire [11:0] sel_296453;
  wire [10:0] add_296455;
  wire [11:0] sel_296457;
  wire [8:0] add_296459;
  wire [11:0] sel_296462;
  wire [8:0] add_296464;
  wire [11:0] sel_296467;
  wire [10:0] add_296469;
  wire [11:0] sel_296472;
  wire [10:0] add_296474;
  wire [11:0] sel_296477;
  wire [11:0] add_296502;
  wire [11:0] sel_296504;
  wire [11:0] add_296507;
  wire [11:0] sel_296509;
  wire [15:0] array_index_296538;
  wire [15:0] array_index_296541;
  wire [10:0] add_296545;
  wire [11:0] sel_296547;
  wire [10:0] add_296549;
  wire [11:0] sel_296551;
  wire [10:0] add_296553;
  wire [11:0] sel_296555;
  wire [10:0] add_296557;
  wire [11:0] sel_296559;
  wire [8:0] add_296561;
  wire [11:0] sel_296564;
  wire [8:0] add_296566;
  wire [11:0] sel_296569;
  wire [10:0] add_296571;
  wire [11:0] sel_296574;
  wire [10:0] add_296576;
  wire [11:0] sel_296579;
  wire [11:0] add_296604;
  wire [11:0] sel_296606;
  wire [11:0] add_296609;
  wire [11:0] sel_296611;
  wire [15:0] array_index_296640;
  wire [15:0] array_index_296643;
  wire [10:0] add_296647;
  wire [11:0] sel_296649;
  wire [10:0] add_296651;
  wire [11:0] sel_296653;
  wire [10:0] add_296655;
  wire [11:0] sel_296657;
  wire [10:0] add_296659;
  wire [11:0] sel_296661;
  wire [8:0] add_296663;
  wire [11:0] sel_296666;
  wire [8:0] add_296668;
  wire [11:0] sel_296671;
  wire [10:0] add_296673;
  wire [11:0] sel_296676;
  wire [10:0] add_296678;
  wire [11:0] sel_296681;
  wire [11:0] add_296706;
  wire [11:0] sel_296708;
  wire [11:0] add_296711;
  wire [11:0] sel_296713;
  wire [15:0] array_index_296742;
  wire [15:0] array_index_296745;
  wire [10:0] add_296749;
  wire [11:0] sel_296751;
  wire [10:0] add_296753;
  wire [11:0] sel_296755;
  wire [10:0] add_296757;
  wire [11:0] sel_296759;
  wire [10:0] add_296761;
  wire [11:0] sel_296763;
  wire [8:0] add_296765;
  wire [11:0] sel_296768;
  wire [8:0] add_296770;
  wire [11:0] sel_296773;
  wire [10:0] add_296775;
  wire [11:0] sel_296778;
  wire [10:0] add_296780;
  wire [11:0] sel_296783;
  wire [11:0] add_296808;
  wire [11:0] sel_296810;
  wire [11:0] add_296813;
  wire [11:0] sel_296815;
  wire [15:0] array_index_296844;
  wire [15:0] array_index_296847;
  wire [10:0] add_296851;
  wire [11:0] sel_296853;
  wire [10:0] add_296855;
  wire [11:0] sel_296857;
  wire [10:0] add_296859;
  wire [11:0] sel_296861;
  wire [10:0] add_296863;
  wire [11:0] sel_296865;
  wire [8:0] add_296867;
  wire [11:0] sel_296870;
  wire [8:0] add_296872;
  wire [11:0] sel_296875;
  wire [10:0] add_296877;
  wire [11:0] sel_296880;
  wire [10:0] add_296882;
  wire [11:0] sel_296885;
  wire [11:0] add_296910;
  wire [11:0] sel_296912;
  wire [11:0] add_296915;
  wire [11:0] sel_296917;
  wire [15:0] array_index_296946;
  wire [15:0] array_index_296949;
  wire [10:0] add_296953;
  wire [11:0] sel_296955;
  wire [10:0] add_296957;
  wire [11:0] sel_296959;
  wire [10:0] add_296961;
  wire [11:0] sel_296963;
  wire [10:0] add_296965;
  wire [11:0] sel_296967;
  wire [8:0] add_296969;
  wire [11:0] sel_296972;
  wire [8:0] add_296974;
  wire [11:0] sel_296977;
  wire [10:0] add_296979;
  wire [11:0] sel_296982;
  wire [10:0] add_296984;
  wire [11:0] sel_296987;
  wire [11:0] add_297012;
  wire [11:0] sel_297014;
  wire [11:0] add_297017;
  wire [11:0] sel_297019;
  wire [15:0] array_index_297048;
  wire [15:0] array_index_297051;
  wire [10:0] add_297055;
  wire [11:0] sel_297057;
  wire [10:0] add_297059;
  wire [11:0] sel_297061;
  wire [10:0] add_297063;
  wire [11:0] sel_297065;
  wire [10:0] add_297067;
  wire [11:0] sel_297069;
  wire [8:0] add_297071;
  wire [11:0] sel_297074;
  wire [8:0] add_297076;
  wire [11:0] sel_297079;
  wire [10:0] add_297081;
  wire [11:0] sel_297084;
  wire [10:0] add_297086;
  wire [11:0] sel_297089;
  wire [11:0] add_297114;
  wire [11:0] sel_297116;
  wire [11:0] add_297119;
  wire [11:0] sel_297121;
  wire [15:0] array_index_297150;
  wire [15:0] array_index_297153;
  wire [10:0] add_297157;
  wire [11:0] sel_297159;
  wire [10:0] add_297161;
  wire [11:0] sel_297163;
  wire [10:0] add_297165;
  wire [11:0] sel_297167;
  wire [10:0] add_297169;
  wire [11:0] sel_297171;
  wire [8:0] add_297173;
  wire [11:0] sel_297176;
  wire [8:0] add_297178;
  wire [11:0] sel_297181;
  wire [10:0] add_297183;
  wire [11:0] sel_297186;
  wire [10:0] add_297188;
  wire [11:0] sel_297191;
  wire [11:0] add_297216;
  wire [11:0] sel_297218;
  wire [11:0] add_297221;
  wire [11:0] sel_297223;
  wire [15:0] array_index_297252;
  wire [15:0] array_index_297255;
  wire [10:0] add_297259;
  wire [11:0] sel_297261;
  wire [10:0] add_297263;
  wire [11:0] sel_297265;
  wire [10:0] add_297267;
  wire [11:0] sel_297269;
  wire [10:0] add_297271;
  wire [11:0] sel_297273;
  wire [8:0] add_297275;
  wire [11:0] sel_297278;
  wire [8:0] add_297280;
  wire [11:0] sel_297283;
  wire [10:0] add_297285;
  wire [11:0] sel_297288;
  wire [10:0] add_297290;
  wire [11:0] sel_297293;
  wire [11:0] add_297318;
  wire [11:0] sel_297320;
  wire [11:0] add_297323;
  wire [11:0] sel_297325;
  wire [15:0] array_index_297354;
  wire [15:0] array_index_297357;
  wire [10:0] add_297361;
  wire [11:0] sel_297363;
  wire [10:0] add_297365;
  wire [11:0] sel_297367;
  wire [10:0] add_297369;
  wire [11:0] sel_297371;
  wire [10:0] add_297373;
  wire [11:0] sel_297375;
  wire [8:0] add_297377;
  wire [11:0] sel_297380;
  wire [8:0] add_297382;
  wire [11:0] sel_297385;
  wire [10:0] add_297387;
  wire [11:0] sel_297390;
  wire [10:0] add_297392;
  wire [11:0] sel_297395;
  wire [11:0] add_297420;
  wire [11:0] sel_297422;
  wire [11:0] add_297425;
  wire [11:0] sel_297427;
  wire [15:0] array_index_297456;
  wire [15:0] array_index_297459;
  wire [10:0] add_297463;
  wire [11:0] sel_297465;
  wire [10:0] add_297467;
  wire [11:0] sel_297469;
  wire [10:0] add_297471;
  wire [11:0] sel_297473;
  wire [10:0] add_297475;
  wire [11:0] sel_297477;
  wire [8:0] add_297479;
  wire [11:0] sel_297482;
  wire [8:0] add_297484;
  wire [11:0] sel_297487;
  wire [10:0] add_297489;
  wire [11:0] sel_297492;
  wire [10:0] add_297494;
  wire [11:0] sel_297497;
  wire [11:0] add_297522;
  wire [11:0] sel_297524;
  wire [11:0] add_297527;
  wire [11:0] sel_297529;
  wire [15:0] array_index_297558;
  wire [15:0] array_index_297561;
  wire [10:0] add_297565;
  wire [11:0] sel_297567;
  wire [10:0] add_297569;
  wire [11:0] sel_297571;
  wire [10:0] add_297573;
  wire [11:0] sel_297575;
  wire [10:0] add_297577;
  wire [11:0] sel_297579;
  wire [8:0] add_297581;
  wire [11:0] sel_297584;
  wire [8:0] add_297586;
  wire [11:0] sel_297589;
  wire [10:0] add_297591;
  wire [11:0] sel_297594;
  wire [10:0] add_297596;
  wire [11:0] sel_297599;
  wire [11:0] add_297624;
  wire [11:0] sel_297626;
  wire [11:0] add_297629;
  wire [11:0] sel_297631;
  wire [15:0] array_index_297660;
  wire [15:0] array_index_297663;
  wire [10:0] add_297667;
  wire [11:0] sel_297669;
  wire [10:0] add_297671;
  wire [11:0] sel_297673;
  wire [10:0] add_297675;
  wire [11:0] sel_297677;
  wire [10:0] add_297679;
  wire [11:0] sel_297681;
  wire [8:0] add_297683;
  wire [11:0] sel_297686;
  wire [8:0] add_297688;
  wire [11:0] sel_297691;
  wire [10:0] add_297693;
  wire [11:0] sel_297696;
  wire [10:0] add_297698;
  wire [11:0] sel_297701;
  wire [11:0] add_297726;
  wire [11:0] sel_297728;
  wire [11:0] add_297731;
  wire [11:0] sel_297733;
  wire [15:0] array_index_297762;
  wire [15:0] array_index_297765;
  wire [10:0] add_297769;
  wire [11:0] sel_297771;
  wire [10:0] add_297773;
  wire [11:0] sel_297775;
  wire [10:0] add_297777;
  wire [11:0] sel_297779;
  wire [10:0] add_297781;
  wire [11:0] sel_297783;
  wire [8:0] add_297785;
  wire [11:0] sel_297788;
  wire [8:0] add_297790;
  wire [11:0] sel_297793;
  wire [10:0] add_297795;
  wire [11:0] sel_297798;
  wire [10:0] add_297800;
  wire [11:0] sel_297803;
  wire [11:0] add_297828;
  wire [11:0] sel_297830;
  wire [11:0] add_297833;
  wire [11:0] sel_297835;
  wire [15:0] array_index_297864;
  wire [15:0] array_index_297867;
  wire [10:0] add_297871;
  wire [11:0] sel_297873;
  wire [10:0] add_297875;
  wire [11:0] sel_297877;
  wire [10:0] add_297879;
  wire [11:0] sel_297881;
  wire [10:0] add_297883;
  wire [11:0] sel_297885;
  wire [8:0] add_297887;
  wire [11:0] sel_297890;
  wire [8:0] add_297892;
  wire [11:0] sel_297895;
  wire [10:0] add_297897;
  wire [11:0] sel_297900;
  wire [10:0] add_297902;
  wire [11:0] sel_297905;
  wire [11:0] add_297930;
  wire [11:0] sel_297932;
  wire [11:0] add_297935;
  wire [11:0] sel_297937;
  wire [15:0] array_index_297966;
  wire [15:0] array_index_297969;
  wire [10:0] add_297973;
  wire [11:0] sel_297975;
  wire [10:0] add_297977;
  wire [11:0] sel_297979;
  wire [10:0] add_297981;
  wire [11:0] sel_297983;
  wire [10:0] add_297985;
  wire [11:0] sel_297987;
  wire [8:0] add_297989;
  wire [11:0] sel_297992;
  wire [8:0] add_297994;
  wire [11:0] sel_297997;
  wire [10:0] add_297999;
  wire [11:0] sel_298002;
  wire [10:0] add_298004;
  wire [11:0] sel_298007;
  wire [11:0] add_298032;
  wire [11:0] sel_298034;
  wire [11:0] add_298037;
  wire [11:0] sel_298039;
  wire [15:0] array_index_298068;
  wire [15:0] array_index_298071;
  wire [10:0] add_298075;
  wire [11:0] sel_298077;
  wire [10:0] add_298079;
  wire [11:0] sel_298081;
  wire [10:0] add_298083;
  wire [11:0] sel_298085;
  wire [10:0] add_298087;
  wire [11:0] sel_298089;
  wire [8:0] add_298091;
  wire [11:0] sel_298094;
  wire [8:0] add_298096;
  wire [11:0] sel_298099;
  wire [10:0] add_298101;
  wire [11:0] sel_298104;
  wire [10:0] add_298106;
  wire [11:0] sel_298109;
  wire [11:0] add_298134;
  wire [11:0] sel_298136;
  wire [11:0] add_298139;
  wire [11:0] sel_298141;
  wire [15:0] array_index_298170;
  wire [15:0] array_index_298173;
  wire [10:0] add_298177;
  wire [11:0] sel_298179;
  wire [10:0] add_298181;
  wire [11:0] sel_298183;
  wire [10:0] add_298185;
  wire [11:0] sel_298187;
  wire [10:0] add_298189;
  wire [11:0] sel_298191;
  wire [8:0] add_298193;
  wire [11:0] sel_298196;
  wire [8:0] add_298198;
  wire [11:0] sel_298201;
  wire [10:0] add_298203;
  wire [11:0] sel_298206;
  wire [10:0] add_298208;
  wire [11:0] sel_298211;
  wire [11:0] add_298236;
  wire [11:0] sel_298238;
  wire [11:0] add_298241;
  wire [11:0] sel_298243;
  wire [15:0] array_index_298272;
  wire [15:0] array_index_298275;
  wire [10:0] add_298279;
  wire [11:0] sel_298281;
  wire [10:0] add_298283;
  wire [11:0] sel_298285;
  wire [10:0] add_298287;
  wire [11:0] sel_298289;
  wire [10:0] add_298291;
  wire [11:0] sel_298293;
  wire [8:0] add_298295;
  wire [11:0] sel_298298;
  wire [8:0] add_298300;
  wire [11:0] sel_298303;
  wire [10:0] add_298305;
  wire [11:0] sel_298308;
  wire [10:0] add_298310;
  wire [11:0] sel_298313;
  wire [11:0] add_298338;
  wire [11:0] sel_298340;
  wire [11:0] add_298343;
  wire [11:0] sel_298345;
  wire [15:0] array_index_298374;
  wire [15:0] array_index_298377;
  wire [10:0] add_298381;
  wire [11:0] sel_298383;
  wire [10:0] add_298385;
  wire [11:0] sel_298387;
  wire [10:0] add_298389;
  wire [11:0] sel_298391;
  wire [10:0] add_298393;
  wire [11:0] sel_298395;
  wire [8:0] add_298397;
  wire [11:0] sel_298400;
  wire [8:0] add_298402;
  wire [11:0] sel_298405;
  wire [10:0] add_298407;
  wire [11:0] sel_298410;
  wire [10:0] add_298412;
  wire [11:0] sel_298415;
  wire [11:0] add_298440;
  wire [11:0] sel_298442;
  wire [11:0] add_298445;
  wire [11:0] sel_298447;
  wire [15:0] array_index_298476;
  wire [15:0] array_index_298479;
  wire [10:0] add_298483;
  wire [11:0] sel_298485;
  wire [10:0] add_298487;
  wire [11:0] sel_298489;
  wire [10:0] add_298491;
  wire [11:0] sel_298493;
  wire [10:0] add_298495;
  wire [11:0] sel_298497;
  wire [8:0] add_298499;
  wire [11:0] sel_298502;
  wire [8:0] add_298504;
  wire [11:0] sel_298507;
  wire [10:0] add_298509;
  wire [11:0] sel_298512;
  wire [10:0] add_298514;
  wire [11:0] sel_298517;
  wire [11:0] add_298542;
  wire [11:0] sel_298544;
  wire [11:0] add_298547;
  wire [11:0] sel_298549;
  wire [15:0] array_index_298578;
  wire [15:0] array_index_298581;
  wire [10:0] add_298585;
  wire [11:0] sel_298587;
  wire [10:0] add_298589;
  wire [11:0] sel_298591;
  wire [10:0] add_298593;
  wire [11:0] sel_298595;
  wire [10:0] add_298597;
  wire [11:0] sel_298599;
  wire [8:0] add_298601;
  wire [11:0] sel_298604;
  wire [8:0] add_298606;
  wire [11:0] sel_298609;
  wire [10:0] add_298611;
  wire [11:0] sel_298614;
  wire [10:0] add_298616;
  wire [11:0] sel_298619;
  wire [11:0] add_298644;
  wire [11:0] sel_298646;
  wire [11:0] add_298649;
  wire [11:0] sel_298651;
  wire [15:0] array_index_298680;
  wire [15:0] array_index_298683;
  wire [10:0] add_298687;
  wire [11:0] sel_298689;
  wire [10:0] add_298691;
  wire [11:0] sel_298693;
  wire [10:0] add_298695;
  wire [11:0] sel_298697;
  wire [10:0] add_298699;
  wire [11:0] sel_298701;
  wire [8:0] add_298703;
  wire [11:0] sel_298706;
  wire [8:0] add_298708;
  wire [11:0] sel_298711;
  wire [10:0] add_298713;
  wire [11:0] sel_298716;
  wire [10:0] add_298718;
  wire [11:0] sel_298721;
  wire [11:0] add_298746;
  wire [11:0] sel_298748;
  wire [11:0] add_298751;
  wire [11:0] sel_298753;
  wire [15:0] array_index_298782;
  wire [15:0] array_index_298785;
  wire [10:0] add_298789;
  wire [11:0] sel_298791;
  wire [10:0] add_298793;
  wire [11:0] sel_298795;
  wire [10:0] add_298797;
  wire [11:0] sel_298799;
  wire [10:0] add_298801;
  wire [11:0] sel_298803;
  wire [8:0] add_298805;
  wire [11:0] sel_298808;
  wire [8:0] add_298810;
  wire [11:0] sel_298813;
  wire [10:0] add_298815;
  wire [11:0] sel_298818;
  wire [10:0] add_298820;
  wire [11:0] sel_298823;
  wire [11:0] add_298848;
  wire [11:0] sel_298850;
  wire [11:0] add_298853;
  wire [11:0] sel_298855;
  wire [15:0] array_index_298884;
  wire [15:0] array_index_298887;
  wire [10:0] add_298891;
  wire [11:0] sel_298893;
  wire [10:0] add_298895;
  wire [11:0] sel_298897;
  wire [10:0] add_298899;
  wire [11:0] sel_298901;
  wire [10:0] add_298903;
  wire [11:0] sel_298905;
  wire [8:0] add_298907;
  wire [11:0] sel_298910;
  wire [8:0] add_298912;
  wire [11:0] sel_298915;
  wire [10:0] add_298917;
  wire [11:0] sel_298920;
  wire [10:0] add_298922;
  wire [11:0] sel_298925;
  wire [11:0] add_298950;
  wire [11:0] sel_298952;
  wire [11:0] add_298955;
  wire [11:0] sel_298957;
  wire [15:0] array_index_298986;
  wire [15:0] array_index_298989;
  wire [10:0] add_298993;
  wire [11:0] sel_298995;
  wire [10:0] add_298997;
  wire [11:0] sel_298999;
  wire [10:0] add_299001;
  wire [11:0] sel_299003;
  wire [10:0] add_299005;
  wire [11:0] sel_299007;
  wire [8:0] add_299009;
  wire [11:0] sel_299012;
  wire [8:0] add_299014;
  wire [11:0] sel_299017;
  wire [10:0] add_299019;
  wire [11:0] sel_299022;
  wire [10:0] add_299024;
  wire [11:0] sel_299027;
  wire [11:0] add_299052;
  wire [11:0] sel_299054;
  wire [11:0] add_299057;
  wire [11:0] sel_299059;
  wire [15:0] array_index_299088;
  wire [15:0] array_index_299091;
  wire [10:0] add_299095;
  wire [11:0] sel_299097;
  wire [10:0] add_299099;
  wire [11:0] sel_299101;
  wire [10:0] add_299103;
  wire [11:0] sel_299105;
  wire [10:0] add_299107;
  wire [11:0] sel_299109;
  wire [8:0] add_299111;
  wire [11:0] sel_299114;
  wire [8:0] add_299116;
  wire [11:0] sel_299119;
  wire [10:0] add_299121;
  wire [11:0] sel_299124;
  wire [10:0] add_299126;
  wire [11:0] sel_299129;
  wire [11:0] add_299154;
  wire [11:0] sel_299156;
  wire [11:0] add_299159;
  wire [11:0] sel_299161;
  wire [15:0] array_index_299190;
  wire [15:0] array_index_299193;
  wire [10:0] add_299197;
  wire [11:0] sel_299199;
  wire [10:0] add_299201;
  wire [11:0] sel_299203;
  wire [10:0] add_299205;
  wire [11:0] sel_299207;
  wire [10:0] add_299209;
  wire [11:0] sel_299211;
  wire [8:0] add_299213;
  wire [11:0] sel_299216;
  wire [8:0] add_299218;
  wire [11:0] sel_299221;
  wire [10:0] add_299223;
  wire [11:0] sel_299226;
  wire [10:0] add_299228;
  wire [11:0] sel_299231;
  wire [11:0] add_299256;
  wire [11:0] sel_299258;
  wire [11:0] add_299261;
  wire [11:0] sel_299263;
  wire [15:0] array_index_299292;
  wire [15:0] array_index_299295;
  wire [10:0] add_299299;
  wire [11:0] sel_299301;
  wire [10:0] add_299303;
  wire [11:0] sel_299305;
  wire [10:0] add_299307;
  wire [11:0] sel_299309;
  wire [10:0] add_299311;
  wire [11:0] sel_299313;
  wire [8:0] add_299315;
  wire [11:0] sel_299318;
  wire [8:0] add_299320;
  wire [11:0] sel_299323;
  wire [10:0] add_299325;
  wire [11:0] sel_299328;
  wire [10:0] add_299330;
  wire [11:0] sel_299333;
  wire [11:0] add_299358;
  wire [11:0] sel_299360;
  wire [11:0] add_299363;
  wire [11:0] sel_299365;
  wire [15:0] array_index_299394;
  wire [15:0] array_index_299397;
  wire [10:0] add_299401;
  wire [11:0] sel_299403;
  wire [10:0] add_299405;
  wire [11:0] sel_299407;
  wire [10:0] add_299409;
  wire [11:0] sel_299411;
  wire [10:0] add_299413;
  wire [11:0] sel_299415;
  wire [8:0] add_299417;
  wire [11:0] sel_299420;
  wire [8:0] add_299422;
  wire [11:0] sel_299425;
  wire [10:0] add_299427;
  wire [11:0] sel_299430;
  wire [10:0] add_299432;
  wire [11:0] sel_299435;
  wire [11:0] add_299460;
  wire [11:0] sel_299462;
  wire [11:0] add_299465;
  wire [11:0] sel_299467;
  wire [15:0] array_index_299496;
  wire [15:0] array_index_299499;
  wire [10:0] add_299503;
  wire [11:0] sel_299505;
  wire [10:0] add_299507;
  wire [11:0] sel_299509;
  wire [10:0] add_299511;
  wire [11:0] sel_299513;
  wire [10:0] add_299515;
  wire [11:0] sel_299517;
  wire [8:0] add_299519;
  wire [11:0] sel_299522;
  wire [8:0] add_299524;
  wire [11:0] sel_299527;
  wire [10:0] add_299529;
  wire [11:0] sel_299532;
  wire [10:0] add_299534;
  wire [11:0] sel_299537;
  wire [11:0] add_299562;
  wire [11:0] sel_299564;
  wire [11:0] add_299567;
  wire [11:0] sel_299569;
  wire [15:0] array_index_299598;
  wire [15:0] array_index_299601;
  wire [10:0] add_299605;
  wire [11:0] sel_299607;
  wire [10:0] add_299609;
  wire [11:0] sel_299611;
  wire [10:0] add_299613;
  wire [11:0] sel_299615;
  wire [10:0] add_299617;
  wire [11:0] sel_299619;
  wire [8:0] add_299621;
  wire [11:0] sel_299624;
  wire [8:0] add_299626;
  wire [11:0] sel_299629;
  wire [10:0] add_299631;
  wire [11:0] sel_299634;
  wire [10:0] add_299636;
  wire [11:0] sel_299639;
  wire [11:0] add_299664;
  wire [11:0] sel_299666;
  wire [11:0] add_299669;
  wire [11:0] sel_299671;
  wire [15:0] array_index_299700;
  wire [15:0] array_index_299703;
  wire [10:0] add_299707;
  wire [11:0] sel_299709;
  wire [10:0] add_299711;
  wire [11:0] sel_299713;
  wire [10:0] add_299715;
  wire [11:0] sel_299717;
  wire [10:0] add_299719;
  wire [11:0] sel_299721;
  wire [8:0] add_299723;
  wire [11:0] sel_299726;
  wire [8:0] add_299728;
  wire [11:0] sel_299731;
  wire [10:0] add_299733;
  wire [11:0] sel_299736;
  wire [10:0] add_299738;
  wire [11:0] sel_299741;
  wire [11:0] add_299766;
  wire [11:0] sel_299768;
  wire [11:0] add_299771;
  wire [11:0] sel_299773;
  wire [15:0] array_index_299802;
  wire [15:0] array_index_299805;
  wire [10:0] add_299809;
  wire [11:0] sel_299811;
  wire [10:0] add_299813;
  wire [11:0] sel_299815;
  wire [10:0] add_299817;
  wire [11:0] sel_299819;
  wire [10:0] add_299821;
  wire [11:0] sel_299823;
  wire [8:0] add_299825;
  wire [11:0] sel_299828;
  wire [8:0] add_299830;
  wire [11:0] sel_299833;
  wire [10:0] add_299835;
  wire [11:0] sel_299838;
  wire [10:0] add_299840;
  wire [11:0] sel_299843;
  wire [11:0] add_299868;
  wire [11:0] sel_299870;
  wire [11:0] add_299873;
  wire [11:0] sel_299875;
  wire [15:0] array_index_299904;
  wire [15:0] array_index_299907;
  wire [10:0] add_299911;
  wire [11:0] sel_299913;
  wire [10:0] add_299915;
  wire [11:0] sel_299917;
  wire [10:0] add_299919;
  wire [11:0] sel_299921;
  wire [10:0] add_299923;
  wire [11:0] sel_299925;
  wire [8:0] add_299927;
  wire [11:0] sel_299930;
  wire [8:0] add_299932;
  wire [11:0] sel_299935;
  wire [10:0] add_299937;
  wire [11:0] sel_299940;
  wire [10:0] add_299942;
  wire [11:0] sel_299945;
  wire [11:0] add_299970;
  wire [11:0] sel_299972;
  wire [11:0] add_299975;
  wire [11:0] sel_299977;
  wire [15:0] array_index_300006;
  wire [15:0] array_index_300009;
  wire [10:0] add_300013;
  wire [11:0] sel_300015;
  wire [10:0] add_300017;
  wire [11:0] sel_300019;
  wire [10:0] add_300021;
  wire [11:0] sel_300023;
  wire [10:0] add_300025;
  wire [11:0] sel_300027;
  wire [8:0] add_300029;
  wire [11:0] sel_300032;
  wire [8:0] add_300034;
  wire [11:0] sel_300037;
  wire [10:0] add_300039;
  wire [11:0] sel_300042;
  wire [10:0] add_300044;
  wire [11:0] sel_300047;
  wire [11:0] add_300072;
  wire [11:0] sel_300074;
  wire [11:0] add_300077;
  wire [11:0] sel_300079;
  wire [15:0] array_index_300108;
  wire [15:0] array_index_300111;
  wire [10:0] add_300115;
  wire [11:0] sel_300117;
  wire [10:0] add_300119;
  wire [11:0] sel_300121;
  wire [10:0] add_300123;
  wire [11:0] sel_300125;
  wire [10:0] add_300127;
  wire [11:0] sel_300129;
  wire [8:0] add_300131;
  wire [11:0] sel_300134;
  wire [8:0] add_300136;
  wire [11:0] sel_300139;
  wire [10:0] add_300141;
  wire [11:0] sel_300144;
  wire [10:0] add_300146;
  wire [11:0] sel_300149;
  wire [11:0] add_300174;
  wire [11:0] sel_300176;
  wire [11:0] add_300179;
  wire [11:0] sel_300181;
  wire [15:0] array_index_300210;
  wire [15:0] array_index_300213;
  wire [10:0] add_300217;
  wire [11:0] sel_300219;
  wire [10:0] add_300221;
  wire [11:0] sel_300223;
  wire [10:0] add_300225;
  wire [11:0] sel_300227;
  wire [10:0] add_300229;
  wire [11:0] sel_300231;
  wire [8:0] add_300233;
  wire [11:0] sel_300236;
  wire [8:0] add_300238;
  wire [11:0] sel_300241;
  wire [10:0] add_300243;
  wire [11:0] sel_300246;
  wire [10:0] add_300248;
  wire [11:0] sel_300251;
  wire [11:0] add_300276;
  wire [11:0] sel_300278;
  wire [11:0] add_300281;
  wire [11:0] sel_300283;
  wire [15:0] array_index_300312;
  wire [15:0] array_index_300315;
  wire [10:0] add_300319;
  wire [11:0] sel_300321;
  wire [10:0] add_300323;
  wire [11:0] sel_300325;
  wire [10:0] add_300327;
  wire [11:0] sel_300329;
  wire [10:0] add_300331;
  wire [11:0] sel_300333;
  wire [8:0] add_300335;
  wire [11:0] sel_300338;
  wire [8:0] add_300340;
  wire [11:0] sel_300343;
  wire [10:0] add_300345;
  wire [11:0] sel_300348;
  wire [10:0] add_300350;
  wire [11:0] sel_300353;
  wire [11:0] add_300378;
  wire [11:0] sel_300380;
  wire [11:0] add_300383;
  wire [11:0] sel_300385;
  wire [15:0] array_index_300414;
  wire [15:0] array_index_300417;
  wire [10:0] add_300421;
  wire [11:0] sel_300423;
  wire [10:0] add_300425;
  wire [11:0] sel_300427;
  wire [10:0] add_300429;
  wire [11:0] sel_300431;
  wire [10:0] add_300433;
  wire [11:0] sel_300435;
  wire [8:0] add_300437;
  wire [11:0] sel_300440;
  wire [8:0] add_300442;
  wire [11:0] sel_300445;
  wire [10:0] add_300447;
  wire [11:0] sel_300450;
  wire [10:0] add_300452;
  wire [11:0] sel_300455;
  wire [11:0] add_300480;
  wire [11:0] sel_300482;
  wire [11:0] add_300485;
  wire [11:0] sel_300487;
  wire [15:0] array_index_300516;
  wire [15:0] array_index_300519;
  wire [10:0] add_300523;
  wire [11:0] sel_300525;
  wire [10:0] add_300527;
  wire [11:0] sel_300529;
  wire [10:0] add_300531;
  wire [11:0] sel_300533;
  wire [10:0] add_300535;
  wire [11:0] sel_300537;
  wire [8:0] add_300539;
  wire [11:0] sel_300542;
  wire [8:0] add_300544;
  wire [11:0] sel_300547;
  wire [10:0] add_300549;
  wire [11:0] sel_300552;
  wire [10:0] add_300554;
  wire [11:0] sel_300557;
  wire [11:0] add_300582;
  wire [11:0] sel_300584;
  wire [11:0] add_300587;
  wire [11:0] sel_300589;
  wire [15:0] array_index_300618;
  wire [15:0] array_index_300621;
  wire [10:0] add_300625;
  wire [11:0] sel_300627;
  wire [10:0] add_300629;
  wire [11:0] sel_300631;
  wire [10:0] add_300633;
  wire [11:0] sel_300635;
  wire [10:0] add_300637;
  wire [11:0] sel_300639;
  wire [8:0] add_300641;
  wire [11:0] sel_300644;
  wire [8:0] add_300646;
  wire [11:0] sel_300649;
  wire [10:0] add_300651;
  wire [11:0] sel_300654;
  wire [10:0] add_300656;
  wire [11:0] sel_300659;
  wire [11:0] add_300684;
  wire [11:0] sel_300686;
  wire [11:0] add_300689;
  wire [11:0] sel_300691;
  wire [15:0] array_index_300720;
  wire [15:0] array_index_300723;
  wire [10:0] add_300727;
  wire [11:0] sel_300729;
  wire [10:0] add_300731;
  wire [11:0] sel_300733;
  wire [10:0] add_300735;
  wire [11:0] sel_300737;
  wire [10:0] add_300739;
  wire [11:0] sel_300741;
  wire [8:0] add_300743;
  wire [11:0] sel_300746;
  wire [8:0] add_300748;
  wire [11:0] sel_300751;
  wire [10:0] add_300753;
  wire [11:0] sel_300756;
  wire [10:0] add_300758;
  wire [11:0] sel_300761;
  wire [11:0] add_300786;
  wire [11:0] sel_300788;
  wire [11:0] add_300791;
  wire [11:0] sel_300793;
  wire [15:0] array_index_300822;
  wire [15:0] array_index_300825;
  wire [10:0] add_300829;
  wire [11:0] sel_300831;
  wire [10:0] add_300833;
  wire [11:0] sel_300835;
  wire [10:0] add_300837;
  wire [11:0] sel_300839;
  wire [10:0] add_300841;
  wire [11:0] sel_300843;
  wire [8:0] add_300845;
  wire [11:0] sel_300848;
  wire [8:0] add_300850;
  wire [11:0] sel_300853;
  wire [10:0] add_300855;
  wire [11:0] sel_300858;
  wire [10:0] add_300860;
  wire [11:0] sel_300863;
  wire [11:0] add_300888;
  wire [11:0] sel_300890;
  wire [11:0] add_300893;
  wire [11:0] sel_300895;
  wire [15:0] array_index_300924;
  wire [15:0] array_index_300927;
  wire [10:0] add_300931;
  wire [11:0] sel_300933;
  wire [10:0] add_300935;
  wire [11:0] sel_300937;
  wire [10:0] add_300939;
  wire [11:0] sel_300941;
  wire [10:0] add_300943;
  wire [11:0] sel_300945;
  wire [8:0] add_300947;
  wire [11:0] sel_300950;
  wire [8:0] add_300952;
  wire [11:0] sel_300955;
  wire [10:0] add_300957;
  wire [11:0] sel_300960;
  wire [10:0] add_300962;
  wire [11:0] sel_300965;
  wire [11:0] add_300990;
  wire [11:0] sel_300992;
  wire [11:0] add_300995;
  wire [11:0] sel_300997;
  wire [15:0] array_index_301026;
  wire [15:0] array_index_301029;
  wire [10:0] add_301033;
  wire [11:0] sel_301035;
  wire [10:0] add_301037;
  wire [11:0] sel_301039;
  wire [10:0] add_301041;
  wire [11:0] sel_301043;
  wire [10:0] add_301045;
  wire [11:0] sel_301047;
  wire [8:0] add_301049;
  wire [11:0] sel_301052;
  wire [8:0] add_301054;
  wire [11:0] sel_301057;
  wire [10:0] add_301059;
  wire [11:0] sel_301062;
  wire [10:0] add_301064;
  wire [11:0] sel_301067;
  wire [11:0] add_301092;
  wire [11:0] sel_301094;
  wire [11:0] add_301097;
  wire [11:0] sel_301099;
  wire [15:0] array_index_301128;
  wire [15:0] array_index_301131;
  wire [10:0] add_301135;
  wire [11:0] sel_301137;
  wire [10:0] add_301139;
  wire [11:0] sel_301141;
  wire [10:0] add_301143;
  wire [11:0] sel_301145;
  wire [10:0] add_301147;
  wire [11:0] sel_301149;
  wire [8:0] add_301151;
  wire [11:0] sel_301154;
  wire [8:0] add_301156;
  wire [11:0] sel_301159;
  wire [10:0] add_301161;
  wire [11:0] sel_301164;
  wire [10:0] add_301166;
  wire [11:0] sel_301169;
  wire [11:0] add_301194;
  wire [11:0] sel_301196;
  wire [11:0] add_301199;
  wire [11:0] sel_301201;
  wire [15:0] array_index_301230;
  wire [15:0] array_index_301233;
  wire [10:0] add_301237;
  wire [11:0] sel_301239;
  wire [10:0] add_301241;
  wire [11:0] sel_301243;
  wire [10:0] add_301245;
  wire [11:0] sel_301247;
  wire [10:0] add_301249;
  wire [11:0] sel_301251;
  wire [8:0] add_301253;
  wire [11:0] sel_301256;
  wire [8:0] add_301258;
  wire [11:0] sel_301261;
  wire [10:0] add_301263;
  wire [11:0] sel_301266;
  wire [10:0] add_301268;
  wire [11:0] sel_301271;
  wire [11:0] add_301296;
  wire [11:0] sel_301298;
  wire [11:0] add_301301;
  wire [11:0] sel_301303;
  wire [15:0] array_index_301332;
  wire [15:0] array_index_301335;
  wire [10:0] add_301339;
  wire [11:0] sel_301341;
  wire [10:0] add_301343;
  wire [11:0] sel_301345;
  wire [10:0] add_301347;
  wire [11:0] sel_301349;
  wire [10:0] add_301351;
  wire [11:0] sel_301353;
  wire [8:0] add_301355;
  wire [11:0] sel_301358;
  wire [8:0] add_301360;
  wire [11:0] sel_301363;
  wire [10:0] add_301365;
  wire [11:0] sel_301368;
  wire [10:0] add_301370;
  wire [11:0] sel_301373;
  wire [11:0] add_301398;
  wire [11:0] sel_301400;
  wire [11:0] add_301403;
  wire [11:0] sel_301405;
  wire [15:0] array_index_301434;
  wire [15:0] array_index_301437;
  wire [10:0] add_301441;
  wire [11:0] sel_301443;
  wire [10:0] add_301445;
  wire [11:0] sel_301447;
  wire [10:0] add_301449;
  wire [11:0] sel_301451;
  wire [10:0] add_301453;
  wire [11:0] sel_301455;
  wire [8:0] add_301457;
  wire [11:0] sel_301460;
  wire [8:0] add_301462;
  wire [11:0] sel_301465;
  wire [10:0] add_301467;
  wire [11:0] sel_301470;
  wire [10:0] add_301472;
  wire [11:0] sel_301475;
  wire [11:0] add_301500;
  wire [11:0] sel_301502;
  wire [11:0] add_301505;
  wire [11:0] sel_301507;
  wire [15:0] array_index_301536;
  wire [15:0] array_index_301539;
  wire [10:0] add_301543;
  wire [11:0] sel_301545;
  wire [10:0] add_301547;
  wire [11:0] sel_301549;
  wire [10:0] add_301551;
  wire [11:0] sel_301553;
  wire [10:0] add_301555;
  wire [11:0] sel_301557;
  wire [8:0] add_301559;
  wire [11:0] sel_301562;
  wire [8:0] add_301564;
  wire [11:0] sel_301567;
  wire [10:0] add_301569;
  wire [11:0] sel_301572;
  wire [10:0] add_301574;
  wire [11:0] sel_301577;
  wire [11:0] add_301602;
  wire [11:0] sel_301604;
  wire [11:0] add_301607;
  wire [11:0] sel_301609;
  wire [15:0] array_index_301638;
  wire [15:0] array_index_301641;
  wire [10:0] add_301645;
  wire [11:0] sel_301647;
  wire [10:0] add_301649;
  wire [11:0] sel_301651;
  wire [10:0] add_301653;
  wire [11:0] sel_301655;
  wire [10:0] add_301657;
  wire [11:0] sel_301659;
  wire [8:0] add_301661;
  wire [11:0] sel_301664;
  wire [8:0] add_301666;
  wire [11:0] sel_301669;
  wire [10:0] add_301671;
  wire [11:0] sel_301674;
  wire [10:0] add_301676;
  wire [11:0] sel_301679;
  wire [11:0] add_301704;
  wire [11:0] sel_301706;
  wire [11:0] add_301709;
  wire [11:0] sel_301711;
  wire [15:0] array_index_301740;
  wire [15:0] array_index_301743;
  wire [10:0] add_301747;
  wire [11:0] sel_301749;
  wire [10:0] add_301751;
  wire [11:0] sel_301753;
  wire [10:0] add_301755;
  wire [11:0] sel_301757;
  wire [10:0] add_301759;
  wire [11:0] sel_301761;
  wire [8:0] add_301763;
  wire [11:0] sel_301766;
  wire [8:0] add_301768;
  wire [11:0] sel_301771;
  wire [10:0] add_301773;
  wire [11:0] sel_301776;
  wire [10:0] add_301778;
  wire [11:0] sel_301781;
  wire [11:0] add_301806;
  wire [11:0] sel_301808;
  wire [11:0] add_301811;
  wire [11:0] sel_301813;
  wire [15:0] array_index_301842;
  wire [15:0] array_index_301845;
  wire [10:0] add_301849;
  wire [11:0] sel_301851;
  wire [10:0] add_301853;
  wire [11:0] sel_301855;
  wire [10:0] add_301857;
  wire [11:0] sel_301859;
  wire [10:0] add_301861;
  wire [11:0] sel_301863;
  wire [8:0] add_301865;
  wire [11:0] sel_301868;
  wire [8:0] add_301870;
  wire [11:0] sel_301873;
  wire [10:0] add_301875;
  wire [11:0] sel_301878;
  wire [10:0] add_301880;
  wire [11:0] sel_301883;
  wire [11:0] add_301908;
  wire [11:0] sel_301910;
  wire [11:0] add_301913;
  wire [11:0] sel_301915;
  wire [15:0] array_index_301944;
  wire [15:0] array_index_301947;
  wire [10:0] add_301951;
  wire [11:0] sel_301953;
  wire [10:0] add_301955;
  wire [11:0] sel_301957;
  wire [10:0] add_301959;
  wire [11:0] sel_301961;
  wire [10:0] add_301963;
  wire [11:0] sel_301965;
  wire [8:0] add_301967;
  wire [11:0] sel_301970;
  wire [8:0] add_301972;
  wire [11:0] sel_301975;
  wire [10:0] add_301977;
  wire [11:0] sel_301980;
  wire [10:0] add_301982;
  wire [11:0] sel_301985;
  wire [11:0] add_302010;
  wire [11:0] sel_302012;
  wire [11:0] add_302015;
  wire [11:0] sel_302017;
  wire [15:0] array_index_302046;
  wire [15:0] array_index_302049;
  wire [10:0] add_302053;
  wire [11:0] sel_302055;
  wire [10:0] add_302057;
  wire [11:0] sel_302059;
  wire [10:0] add_302061;
  wire [11:0] sel_302063;
  wire [10:0] add_302065;
  wire [11:0] sel_302067;
  wire [8:0] add_302069;
  wire [11:0] sel_302072;
  wire [8:0] add_302074;
  wire [11:0] sel_302077;
  wire [10:0] add_302079;
  wire [11:0] sel_302082;
  wire [10:0] add_302084;
  wire [11:0] sel_302087;
  wire [11:0] add_302112;
  wire [11:0] sel_302114;
  wire [11:0] add_302117;
  wire [11:0] sel_302119;
  wire [15:0] array_index_302148;
  wire [15:0] array_index_302151;
  wire [10:0] add_302155;
  wire [11:0] sel_302157;
  wire [10:0] add_302159;
  wire [11:0] sel_302161;
  wire [10:0] add_302163;
  wire [11:0] sel_302165;
  wire [10:0] add_302167;
  wire [11:0] sel_302169;
  wire [8:0] add_302171;
  wire [11:0] sel_302174;
  wire [8:0] add_302176;
  wire [11:0] sel_302179;
  wire [10:0] add_302181;
  wire [11:0] sel_302184;
  wire [10:0] add_302186;
  wire [11:0] sel_302189;
  wire [11:0] add_302214;
  wire [11:0] sel_302216;
  wire [11:0] add_302219;
  wire [11:0] sel_302221;
  wire [15:0] array_index_302250;
  wire [15:0] array_index_302253;
  wire [10:0] add_302257;
  wire [11:0] sel_302259;
  wire [10:0] add_302261;
  wire [11:0] sel_302263;
  wire [10:0] add_302265;
  wire [11:0] sel_302267;
  wire [10:0] add_302269;
  wire [11:0] sel_302271;
  wire [8:0] add_302273;
  wire [11:0] sel_302276;
  wire [8:0] add_302278;
  wire [11:0] sel_302281;
  wire [10:0] add_302283;
  wire [11:0] sel_302286;
  wire [10:0] add_302288;
  wire [11:0] sel_302291;
  wire [11:0] add_302316;
  wire [11:0] sel_302318;
  wire [11:0] add_302321;
  wire [11:0] sel_302323;
  wire [15:0] array_index_302352;
  wire [15:0] array_index_302355;
  wire [10:0] add_302359;
  wire [11:0] sel_302361;
  wire [10:0] add_302363;
  wire [11:0] sel_302365;
  wire [10:0] add_302367;
  wire [11:0] sel_302369;
  wire [10:0] add_302371;
  wire [11:0] sel_302373;
  wire [8:0] add_302375;
  wire [11:0] sel_302378;
  wire [8:0] add_302380;
  wire [11:0] sel_302383;
  wire [10:0] add_302385;
  wire [11:0] sel_302388;
  wire [10:0] add_302390;
  wire [11:0] sel_302393;
  wire [11:0] add_302418;
  wire [11:0] sel_302420;
  wire [11:0] add_302423;
  wire [11:0] sel_302425;
  wire [15:0] array_index_302454;
  wire [15:0] array_index_302457;
  wire [10:0] add_302461;
  wire [11:0] sel_302463;
  wire [10:0] add_302465;
  wire [11:0] sel_302467;
  wire [10:0] add_302469;
  wire [11:0] sel_302471;
  wire [10:0] add_302473;
  wire [11:0] sel_302475;
  wire [8:0] add_302477;
  wire [11:0] sel_302480;
  wire [8:0] add_302482;
  wire [11:0] sel_302485;
  wire [10:0] add_302487;
  wire [11:0] sel_302490;
  wire [10:0] add_302492;
  wire [11:0] sel_302495;
  wire [11:0] add_302520;
  wire [11:0] sel_302522;
  wire [11:0] add_302525;
  wire [11:0] sel_302527;
  wire [15:0] array_index_302556;
  wire [15:0] array_index_302559;
  wire [10:0] add_302563;
  wire [11:0] sel_302565;
  wire [10:0] add_302567;
  wire [11:0] sel_302569;
  wire [10:0] add_302571;
  wire [11:0] sel_302573;
  wire [10:0] add_302575;
  wire [11:0] sel_302577;
  wire [8:0] add_302579;
  wire [11:0] sel_302582;
  wire [8:0] add_302584;
  wire [11:0] sel_302587;
  wire [10:0] add_302589;
  wire [11:0] sel_302592;
  wire [10:0] add_302594;
  wire [11:0] sel_302597;
  wire [11:0] add_302622;
  wire [11:0] sel_302624;
  wire [11:0] add_302627;
  wire [11:0] sel_302629;
  wire [15:0] array_index_302658;
  wire [15:0] array_index_302661;
  wire [10:0] add_302665;
  wire [11:0] sel_302667;
  wire [10:0] add_302669;
  wire [11:0] sel_302671;
  wire [10:0] add_302673;
  wire [11:0] sel_302675;
  wire [10:0] add_302677;
  wire [11:0] sel_302679;
  wire [8:0] add_302681;
  wire [11:0] sel_302684;
  wire [8:0] add_302686;
  wire [11:0] sel_302689;
  wire [10:0] add_302691;
  wire [11:0] sel_302694;
  wire [10:0] add_302696;
  wire [11:0] sel_302699;
  wire [11:0] add_302724;
  wire [11:0] sel_302726;
  wire [11:0] add_302729;
  wire [11:0] sel_302731;
  wire [15:0] array_index_302760;
  wire [15:0] array_index_302763;
  wire [10:0] add_302767;
  wire [11:0] sel_302769;
  wire [10:0] add_302771;
  wire [11:0] sel_302773;
  wire [10:0] add_302775;
  wire [11:0] sel_302777;
  wire [10:0] add_302779;
  wire [11:0] sel_302781;
  wire [8:0] add_302783;
  wire [11:0] sel_302786;
  wire [8:0] add_302788;
  wire [11:0] sel_302791;
  wire [10:0] add_302793;
  wire [11:0] sel_302796;
  wire [10:0] add_302798;
  wire [11:0] sel_302801;
  wire [11:0] add_302825;
  wire [11:0] sel_302827;
  wire [11:0] add_302829;
  wire [11:0] sel_302831;
  wire [10:0] add_302865;
  wire [11:0] sel_302867;
  wire [10:0] add_302869;
  wire [11:0] sel_302871;
  wire [10:0] add_302873;
  wire [11:0] sel_302875;
  wire [10:0] add_302877;
  wire [11:0] sel_302879;
  wire [8:0] add_302881;
  wire [11:0] sel_302884;
  wire [8:0] add_302886;
  wire [11:0] sel_302889;
  wire [10:0] add_302891;
  wire [11:0] sel_302894;
  wire [10:0] add_302896;
  wire [11:0] sel_302899;
  wire [10:0] add_302947;
  wire [11:0] sel_302949;
  wire [10:0] add_302951;
  wire [11:0] sel_302953;
  wire [10:0] add_302955;
  wire [11:0] sel_302957;
  wire [10:0] add_302959;
  wire [11:0] sel_302961;
  wire [8:0] add_302963;
  wire [11:0] sel_302966;
  wire [8:0] add_302968;
  wire [11:0] sel_302971;
  wire [1:0] concat_302974;
  wire [1:0] add_302989;
  wire [10:0] add_303009;
  wire [11:0] sel_303011;
  wire [10:0] add_303013;
  wire [11:0] sel_303015;
  wire [10:0] add_303017;
  wire [11:0] sel_303019;
  wire [10:0] add_303021;
  wire [11:0] sel_303023;
  wire [2:0] concat_303026;
  wire [2:0] add_303037;
  wire [10:0] add_303051;
  wire [11:0] sel_303053;
  wire [10:0] add_303055;
  wire [11:0] sel_303057;
  wire [3:0] concat_303060;
  wire [3:0] add_303067;
  wire [4:0] concat_303076;
  wire [4:0] add_303079;
  assign array_index_292858 = set1_unflattened[8'h64];
  assign array_index_292859 = set2_unflattened[8'h64];
  assign add_292866 = array_index_292858[11:0] + 12'h247;
  assign add_292869 = array_index_292859[11:0] + 12'h247;
  assign array_index_292874 = set1_unflattened[8'h65];
  assign array_index_292877 = set2_unflattened[8'h65];
  assign add_292881 = array_index_292858[11:1] + 11'h247;
  assign add_292884 = array_index_292859[11:1] + 11'h247;
  assign add_292900 = array_index_292874[11:0] + 12'h247;
  assign sel_292902 = $signed({1'h0, add_292866}) < $signed(13'h0fff) ? add_292866 : 12'hfff;
  assign add_292905 = array_index_292877[11:0] + 12'h247;
  assign sel_292907 = $signed({1'h0, add_292869}) < $signed(13'h0fff) ? add_292869 : 12'hfff;
  assign array_index_292922 = set1_unflattened[8'h66];
  assign array_index_292925 = set2_unflattened[8'h66];
  assign add_292929 = array_index_292858[11:3] + 9'h0bd;
  assign add_292932 = array_index_292859[11:3] + 9'h0bd;
  assign add_292935 = array_index_292874[11:1] + 11'h247;
  assign sel_292938 = $signed({1'h0, add_292881, array_index_292858[0]}) < $signed(13'h0fff) ? {add_292881, array_index_292858[0]} : 12'hfff;
  assign add_292940 = array_index_292877[11:1] + 11'h247;
  assign sel_292943 = $signed({1'h0, add_292884, array_index_292859[0]}) < $signed(13'h0fff) ? {add_292884, array_index_292859[0]} : 12'hfff;
  assign add_292960 = array_index_292922[11:0] + 12'h247;
  assign sel_292962 = $signed({1'h0, add_292900}) < $signed({1'h0, sel_292902}) ? add_292900 : sel_292902;
  assign add_292965 = array_index_292925[11:0] + 12'h247;
  assign sel_292967 = $signed({1'h0, add_292905}) < $signed({1'h0, sel_292907}) ? add_292905 : sel_292907;
  assign array_index_292988 = set1_unflattened[8'h67];
  assign array_index_292991 = set2_unflattened[8'h67];
  assign add_292995 = array_index_292858[11:1] + 11'h347;
  assign add_292997 = array_index_292859[11:1] + 11'h347;
  assign add_292999 = array_index_292874[11:3] + 9'h0bd;
  assign sel_293002 = $signed({1'h0, add_292929, array_index_292858[2:0]}) < $signed(13'h0fff) ? {add_292929, array_index_292858[2:0]} : 12'hfff;
  assign add_293004 = array_index_292877[11:3] + 9'h0bd;
  assign sel_293007 = $signed({1'h0, add_292932, array_index_292859[2:0]}) < $signed(13'h0fff) ? {add_292932, array_index_292859[2:0]} : 12'hfff;
  assign add_293009 = array_index_292922[11:1] + 11'h247;
  assign sel_293012 = $signed({1'h0, add_292935, array_index_292874[0]}) < $signed({1'h0, sel_292938}) ? {add_292935, array_index_292874[0]} : sel_292938;
  assign add_293014 = array_index_292925[11:1] + 11'h247;
  assign sel_293017 = $signed({1'h0, add_292940, array_index_292877[0]}) < $signed({1'h0, sel_292943}) ? {add_292940, array_index_292877[0]} : sel_292943;
  assign add_293038 = array_index_292988[11:0] + 12'h247;
  assign sel_293040 = $signed({1'h0, add_292960}) < $signed({1'h0, sel_292962}) ? add_292960 : sel_292962;
  assign add_293043 = array_index_292991[11:0] + 12'h247;
  assign sel_293045 = $signed({1'h0, add_292965}) < $signed({1'h0, sel_292967}) ? add_292965 : sel_292967;
  assign array_index_293072 = set1_unflattened[8'h68];
  assign array_index_293075 = set2_unflattened[8'h68];
  assign add_293079 = array_index_292858[11:1] + 11'h79d;
  assign add_293081 = array_index_292859[11:1] + 11'h79d;
  assign add_293083 = array_index_292874[11:1] + 11'h347;
  assign sel_293085 = $signed({1'h0, add_292995, array_index_292858[0]}) < $signed(13'h0fff) ? {add_292995, array_index_292858[0]} : 12'hfff;
  assign add_293087 = array_index_292877[11:1] + 11'h347;
  assign sel_293089 = $signed({1'h0, add_292997, array_index_292859[0]}) < $signed(13'h0fff) ? {add_292997, array_index_292859[0]} : 12'hfff;
  assign add_293091 = array_index_292922[11:3] + 9'h0bd;
  assign sel_293094 = $signed({1'h0, add_292999, array_index_292874[2:0]}) < $signed({1'h0, sel_293002}) ? {add_292999, array_index_292874[2:0]} : sel_293002;
  assign add_293096 = array_index_292925[11:3] + 9'h0bd;
  assign sel_293099 = $signed({1'h0, add_293004, array_index_292877[2:0]}) < $signed({1'h0, sel_293007}) ? {add_293004, array_index_292877[2:0]} : sel_293007;
  assign add_293101 = array_index_292988[11:1] + 11'h247;
  assign sel_293104 = $signed({1'h0, add_293009, array_index_292922[0]}) < $signed({1'h0, sel_293012}) ? {add_293009, array_index_292922[0]} : sel_293012;
  assign add_293106 = array_index_292991[11:1] + 11'h247;
  assign sel_293109 = $signed({1'h0, add_293014, array_index_292925[0]}) < $signed({1'h0, sel_293017}) ? {add_293014, array_index_292925[0]} : sel_293017;
  assign add_293134 = array_index_293072[11:0] + 12'h247;
  assign sel_293136 = $signed({1'h0, add_293038}) < $signed({1'h0, sel_293040}) ? add_293038 : sel_293040;
  assign add_293139 = array_index_293075[11:0] + 12'h247;
  assign sel_293141 = $signed({1'h0, add_293043}) < $signed({1'h0, sel_293045}) ? add_293043 : sel_293045;
  assign array_index_293172 = set1_unflattened[8'h69];
  assign array_index_293175 = set2_unflattened[8'h69];
  assign add_293179 = array_index_292874[11:1] + 11'h79d;
  assign sel_293181 = $signed({1'h0, add_293079, array_index_292858[0]}) < $signed(13'h0fff) ? {add_293079, array_index_292858[0]} : 12'hfff;
  assign add_293183 = array_index_292877[11:1] + 11'h79d;
  assign sel_293185 = $signed({1'h0, add_293081, array_index_292859[0]}) < $signed(13'h0fff) ? {add_293081, array_index_292859[0]} : 12'hfff;
  assign add_293187 = array_index_292922[11:1] + 11'h347;
  assign sel_293189 = $signed({1'h0, add_293083, array_index_292874[0]}) < $signed({1'h0, sel_293085}) ? {add_293083, array_index_292874[0]} : sel_293085;
  assign add_293191 = array_index_292925[11:1] + 11'h347;
  assign sel_293193 = $signed({1'h0, add_293087, array_index_292877[0]}) < $signed({1'h0, sel_293089}) ? {add_293087, array_index_292877[0]} : sel_293089;
  assign add_293195 = array_index_292988[11:3] + 9'h0bd;
  assign sel_293198 = $signed({1'h0, add_293091, array_index_292922[2:0]}) < $signed({1'h0, sel_293094}) ? {add_293091, array_index_292922[2:0]} : sel_293094;
  assign add_293200 = array_index_292991[11:3] + 9'h0bd;
  assign sel_293203 = $signed({1'h0, add_293096, array_index_292925[2:0]}) < $signed({1'h0, sel_293099}) ? {add_293096, array_index_292925[2:0]} : sel_293099;
  assign add_293205 = array_index_293072[11:1] + 11'h247;
  assign sel_293208 = $signed({1'h0, add_293101, array_index_292988[0]}) < $signed({1'h0, sel_293104}) ? {add_293101, array_index_292988[0]} : sel_293104;
  assign add_293210 = array_index_293075[11:1] + 11'h247;
  assign sel_293213 = $signed({1'h0, add_293106, array_index_292991[0]}) < $signed({1'h0, sel_293109}) ? {add_293106, array_index_292991[0]} : sel_293109;
  assign add_293238 = array_index_293172[11:0] + 12'h247;
  assign sel_293240 = $signed({1'h0, add_293134}) < $signed({1'h0, sel_293136}) ? add_293134 : sel_293136;
  assign add_293243 = array_index_293175[11:0] + 12'h247;
  assign sel_293245 = $signed({1'h0, add_293139}) < $signed({1'h0, sel_293141}) ? add_293139 : sel_293141;
  assign array_index_293274 = set1_unflattened[8'h6a];
  assign array_index_293277 = set2_unflattened[8'h6a];
  assign add_293281 = array_index_292922[11:1] + 11'h79d;
  assign sel_293283 = $signed({1'h0, add_293179, array_index_292874[0]}) < $signed({1'h0, sel_293181}) ? {add_293179, array_index_292874[0]} : sel_293181;
  assign add_293285 = array_index_292925[11:1] + 11'h79d;
  assign sel_293287 = $signed({1'h0, add_293183, array_index_292877[0]}) < $signed({1'h0, sel_293185}) ? {add_293183, array_index_292877[0]} : sel_293185;
  assign add_293289 = array_index_292988[11:1] + 11'h347;
  assign sel_293291 = $signed({1'h0, add_293187, array_index_292922[0]}) < $signed({1'h0, sel_293189}) ? {add_293187, array_index_292922[0]} : sel_293189;
  assign add_293293 = array_index_292991[11:1] + 11'h347;
  assign sel_293295 = $signed({1'h0, add_293191, array_index_292925[0]}) < $signed({1'h0, sel_293193}) ? {add_293191, array_index_292925[0]} : sel_293193;
  assign add_293297 = array_index_293072[11:3] + 9'h0bd;
  assign sel_293300 = $signed({1'h0, add_293195, array_index_292988[2:0]}) < $signed({1'h0, sel_293198}) ? {add_293195, array_index_292988[2:0]} : sel_293198;
  assign add_293302 = array_index_293075[11:3] + 9'h0bd;
  assign sel_293305 = $signed({1'h0, add_293200, array_index_292991[2:0]}) < $signed({1'h0, sel_293203}) ? {add_293200, array_index_292991[2:0]} : sel_293203;
  assign add_293307 = array_index_293172[11:1] + 11'h247;
  assign sel_293310 = $signed({1'h0, add_293205, array_index_293072[0]}) < $signed({1'h0, sel_293208}) ? {add_293205, array_index_293072[0]} : sel_293208;
  assign add_293312 = array_index_293175[11:1] + 11'h247;
  assign sel_293315 = $signed({1'h0, add_293210, array_index_293075[0]}) < $signed({1'h0, sel_293213}) ? {add_293210, array_index_293075[0]} : sel_293213;
  assign add_293340 = array_index_293274[11:0] + 12'h247;
  assign sel_293342 = $signed({1'h0, add_293238}) < $signed({1'h0, sel_293240}) ? add_293238 : sel_293240;
  assign add_293345 = array_index_293277[11:0] + 12'h247;
  assign sel_293347 = $signed({1'h0, add_293243}) < $signed({1'h0, sel_293245}) ? add_293243 : sel_293245;
  assign array_index_293376 = set1_unflattened[8'h6b];
  assign array_index_293379 = set2_unflattened[8'h6b];
  assign add_293383 = array_index_292988[11:1] + 11'h79d;
  assign sel_293385 = $signed({1'h0, add_293281, array_index_292922[0]}) < $signed({1'h0, sel_293283}) ? {add_293281, array_index_292922[0]} : sel_293283;
  assign add_293387 = array_index_292991[11:1] + 11'h79d;
  assign sel_293389 = $signed({1'h0, add_293285, array_index_292925[0]}) < $signed({1'h0, sel_293287}) ? {add_293285, array_index_292925[0]} : sel_293287;
  assign add_293391 = array_index_293072[11:1] + 11'h347;
  assign sel_293393 = $signed({1'h0, add_293289, array_index_292988[0]}) < $signed({1'h0, sel_293291}) ? {add_293289, array_index_292988[0]} : sel_293291;
  assign add_293395 = array_index_293075[11:1] + 11'h347;
  assign sel_293397 = $signed({1'h0, add_293293, array_index_292991[0]}) < $signed({1'h0, sel_293295}) ? {add_293293, array_index_292991[0]} : sel_293295;
  assign add_293399 = array_index_293172[11:3] + 9'h0bd;
  assign sel_293402 = $signed({1'h0, add_293297, array_index_293072[2:0]}) < $signed({1'h0, sel_293300}) ? {add_293297, array_index_293072[2:0]} : sel_293300;
  assign add_293404 = array_index_293175[11:3] + 9'h0bd;
  assign sel_293407 = $signed({1'h0, add_293302, array_index_293075[2:0]}) < $signed({1'h0, sel_293305}) ? {add_293302, array_index_293075[2:0]} : sel_293305;
  assign add_293409 = array_index_293274[11:1] + 11'h247;
  assign sel_293412 = $signed({1'h0, add_293307, array_index_293172[0]}) < $signed({1'h0, sel_293310}) ? {add_293307, array_index_293172[0]} : sel_293310;
  assign add_293414 = array_index_293277[11:1] + 11'h247;
  assign sel_293417 = $signed({1'h0, add_293312, array_index_293175[0]}) < $signed({1'h0, sel_293315}) ? {add_293312, array_index_293175[0]} : sel_293315;
  assign add_293442 = array_index_293376[11:0] + 12'h247;
  assign sel_293444 = $signed({1'h0, add_293340}) < $signed({1'h0, sel_293342}) ? add_293340 : sel_293342;
  assign add_293447 = array_index_293379[11:0] + 12'h247;
  assign sel_293449 = $signed({1'h0, add_293345}) < $signed({1'h0, sel_293347}) ? add_293345 : sel_293347;
  assign array_index_293478 = set1_unflattened[8'h6c];
  assign array_index_293481 = set2_unflattened[8'h6c];
  assign add_293485 = array_index_293072[11:1] + 11'h79d;
  assign sel_293487 = $signed({1'h0, add_293383, array_index_292988[0]}) < $signed({1'h0, sel_293385}) ? {add_293383, array_index_292988[0]} : sel_293385;
  assign add_293489 = array_index_293075[11:1] + 11'h79d;
  assign sel_293491 = $signed({1'h0, add_293387, array_index_292991[0]}) < $signed({1'h0, sel_293389}) ? {add_293387, array_index_292991[0]} : sel_293389;
  assign add_293493 = array_index_293172[11:1] + 11'h347;
  assign sel_293495 = $signed({1'h0, add_293391, array_index_293072[0]}) < $signed({1'h0, sel_293393}) ? {add_293391, array_index_293072[0]} : sel_293393;
  assign add_293497 = array_index_293175[11:1] + 11'h347;
  assign sel_293499 = $signed({1'h0, add_293395, array_index_293075[0]}) < $signed({1'h0, sel_293397}) ? {add_293395, array_index_293075[0]} : sel_293397;
  assign add_293501 = array_index_293274[11:3] + 9'h0bd;
  assign sel_293504 = $signed({1'h0, add_293399, array_index_293172[2:0]}) < $signed({1'h0, sel_293402}) ? {add_293399, array_index_293172[2:0]} : sel_293402;
  assign add_293506 = array_index_293277[11:3] + 9'h0bd;
  assign sel_293509 = $signed({1'h0, add_293404, array_index_293175[2:0]}) < $signed({1'h0, sel_293407}) ? {add_293404, array_index_293175[2:0]} : sel_293407;
  assign add_293511 = array_index_293376[11:1] + 11'h247;
  assign sel_293514 = $signed({1'h0, add_293409, array_index_293274[0]}) < $signed({1'h0, sel_293412}) ? {add_293409, array_index_293274[0]} : sel_293412;
  assign add_293516 = array_index_293379[11:1] + 11'h247;
  assign sel_293519 = $signed({1'h0, add_293414, array_index_293277[0]}) < $signed({1'h0, sel_293417}) ? {add_293414, array_index_293277[0]} : sel_293417;
  assign add_293544 = array_index_293478[11:0] + 12'h247;
  assign sel_293546 = $signed({1'h0, add_293442}) < $signed({1'h0, sel_293444}) ? add_293442 : sel_293444;
  assign add_293549 = array_index_293481[11:0] + 12'h247;
  assign sel_293551 = $signed({1'h0, add_293447}) < $signed({1'h0, sel_293449}) ? add_293447 : sel_293449;
  assign array_index_293580 = set1_unflattened[8'h6d];
  assign array_index_293583 = set2_unflattened[8'h6d];
  assign add_293587 = array_index_293172[11:1] + 11'h79d;
  assign sel_293589 = $signed({1'h0, add_293485, array_index_293072[0]}) < $signed({1'h0, sel_293487}) ? {add_293485, array_index_293072[0]} : sel_293487;
  assign add_293591 = array_index_293175[11:1] + 11'h79d;
  assign sel_293593 = $signed({1'h0, add_293489, array_index_293075[0]}) < $signed({1'h0, sel_293491}) ? {add_293489, array_index_293075[0]} : sel_293491;
  assign add_293595 = array_index_293274[11:1] + 11'h347;
  assign sel_293597 = $signed({1'h0, add_293493, array_index_293172[0]}) < $signed({1'h0, sel_293495}) ? {add_293493, array_index_293172[0]} : sel_293495;
  assign add_293599 = array_index_293277[11:1] + 11'h347;
  assign sel_293601 = $signed({1'h0, add_293497, array_index_293175[0]}) < $signed({1'h0, sel_293499}) ? {add_293497, array_index_293175[0]} : sel_293499;
  assign add_293603 = array_index_293376[11:3] + 9'h0bd;
  assign sel_293606 = $signed({1'h0, add_293501, array_index_293274[2:0]}) < $signed({1'h0, sel_293504}) ? {add_293501, array_index_293274[2:0]} : sel_293504;
  assign add_293608 = array_index_293379[11:3] + 9'h0bd;
  assign sel_293611 = $signed({1'h0, add_293506, array_index_293277[2:0]}) < $signed({1'h0, sel_293509}) ? {add_293506, array_index_293277[2:0]} : sel_293509;
  assign add_293613 = array_index_293478[11:1] + 11'h247;
  assign sel_293616 = $signed({1'h0, add_293511, array_index_293376[0]}) < $signed({1'h0, sel_293514}) ? {add_293511, array_index_293376[0]} : sel_293514;
  assign add_293618 = array_index_293481[11:1] + 11'h247;
  assign sel_293621 = $signed({1'h0, add_293516, array_index_293379[0]}) < $signed({1'h0, sel_293519}) ? {add_293516, array_index_293379[0]} : sel_293519;
  assign add_293646 = array_index_293580[11:0] + 12'h247;
  assign sel_293648 = $signed({1'h0, add_293544}) < $signed({1'h0, sel_293546}) ? add_293544 : sel_293546;
  assign add_293651 = array_index_293583[11:0] + 12'h247;
  assign sel_293653 = $signed({1'h0, add_293549}) < $signed({1'h0, sel_293551}) ? add_293549 : sel_293551;
  assign array_index_293682 = set1_unflattened[8'h6e];
  assign array_index_293685 = set2_unflattened[8'h6e];
  assign add_293689 = array_index_293274[11:1] + 11'h79d;
  assign sel_293691 = $signed({1'h0, add_293587, array_index_293172[0]}) < $signed({1'h0, sel_293589}) ? {add_293587, array_index_293172[0]} : sel_293589;
  assign add_293693 = array_index_293277[11:1] + 11'h79d;
  assign sel_293695 = $signed({1'h0, add_293591, array_index_293175[0]}) < $signed({1'h0, sel_293593}) ? {add_293591, array_index_293175[0]} : sel_293593;
  assign add_293697 = array_index_293376[11:1] + 11'h347;
  assign sel_293699 = $signed({1'h0, add_293595, array_index_293274[0]}) < $signed({1'h0, sel_293597}) ? {add_293595, array_index_293274[0]} : sel_293597;
  assign add_293701 = array_index_293379[11:1] + 11'h347;
  assign sel_293703 = $signed({1'h0, add_293599, array_index_293277[0]}) < $signed({1'h0, sel_293601}) ? {add_293599, array_index_293277[0]} : sel_293601;
  assign add_293705 = array_index_293478[11:3] + 9'h0bd;
  assign sel_293708 = $signed({1'h0, add_293603, array_index_293376[2:0]}) < $signed({1'h0, sel_293606}) ? {add_293603, array_index_293376[2:0]} : sel_293606;
  assign add_293710 = array_index_293481[11:3] + 9'h0bd;
  assign sel_293713 = $signed({1'h0, add_293608, array_index_293379[2:0]}) < $signed({1'h0, sel_293611}) ? {add_293608, array_index_293379[2:0]} : sel_293611;
  assign add_293715 = array_index_293580[11:1] + 11'h247;
  assign sel_293718 = $signed({1'h0, add_293613, array_index_293478[0]}) < $signed({1'h0, sel_293616}) ? {add_293613, array_index_293478[0]} : sel_293616;
  assign add_293720 = array_index_293583[11:1] + 11'h247;
  assign sel_293723 = $signed({1'h0, add_293618, array_index_293481[0]}) < $signed({1'h0, sel_293621}) ? {add_293618, array_index_293481[0]} : sel_293621;
  assign add_293748 = array_index_293682[11:0] + 12'h247;
  assign sel_293750 = $signed({1'h0, add_293646}) < $signed({1'h0, sel_293648}) ? add_293646 : sel_293648;
  assign add_293753 = array_index_293685[11:0] + 12'h247;
  assign sel_293755 = $signed({1'h0, add_293651}) < $signed({1'h0, sel_293653}) ? add_293651 : sel_293653;
  assign array_index_293784 = set1_unflattened[8'h6f];
  assign array_index_293787 = set2_unflattened[8'h6f];
  assign add_293791 = array_index_293376[11:1] + 11'h79d;
  assign sel_293793 = $signed({1'h0, add_293689, array_index_293274[0]}) < $signed({1'h0, sel_293691}) ? {add_293689, array_index_293274[0]} : sel_293691;
  assign add_293795 = array_index_293379[11:1] + 11'h79d;
  assign sel_293797 = $signed({1'h0, add_293693, array_index_293277[0]}) < $signed({1'h0, sel_293695}) ? {add_293693, array_index_293277[0]} : sel_293695;
  assign add_293799 = array_index_293478[11:1] + 11'h347;
  assign sel_293801 = $signed({1'h0, add_293697, array_index_293376[0]}) < $signed({1'h0, sel_293699}) ? {add_293697, array_index_293376[0]} : sel_293699;
  assign add_293803 = array_index_293481[11:1] + 11'h347;
  assign sel_293805 = $signed({1'h0, add_293701, array_index_293379[0]}) < $signed({1'h0, sel_293703}) ? {add_293701, array_index_293379[0]} : sel_293703;
  assign add_293807 = array_index_293580[11:3] + 9'h0bd;
  assign sel_293810 = $signed({1'h0, add_293705, array_index_293478[2:0]}) < $signed({1'h0, sel_293708}) ? {add_293705, array_index_293478[2:0]} : sel_293708;
  assign add_293812 = array_index_293583[11:3] + 9'h0bd;
  assign sel_293815 = $signed({1'h0, add_293710, array_index_293481[2:0]}) < $signed({1'h0, sel_293713}) ? {add_293710, array_index_293481[2:0]} : sel_293713;
  assign add_293817 = array_index_293682[11:1] + 11'h247;
  assign sel_293820 = $signed({1'h0, add_293715, array_index_293580[0]}) < $signed({1'h0, sel_293718}) ? {add_293715, array_index_293580[0]} : sel_293718;
  assign add_293822 = array_index_293685[11:1] + 11'h247;
  assign sel_293825 = $signed({1'h0, add_293720, array_index_293583[0]}) < $signed({1'h0, sel_293723}) ? {add_293720, array_index_293583[0]} : sel_293723;
  assign add_293850 = array_index_293784[11:0] + 12'h247;
  assign sel_293852 = $signed({1'h0, add_293748}) < $signed({1'h0, sel_293750}) ? add_293748 : sel_293750;
  assign add_293855 = array_index_293787[11:0] + 12'h247;
  assign sel_293857 = $signed({1'h0, add_293753}) < $signed({1'h0, sel_293755}) ? add_293753 : sel_293755;
  assign array_index_293886 = set1_unflattened[8'h70];
  assign array_index_293889 = set2_unflattened[8'h70];
  assign add_293893 = array_index_293478[11:1] + 11'h79d;
  assign sel_293895 = $signed({1'h0, add_293791, array_index_293376[0]}) < $signed({1'h0, sel_293793}) ? {add_293791, array_index_293376[0]} : sel_293793;
  assign add_293897 = array_index_293481[11:1] + 11'h79d;
  assign sel_293899 = $signed({1'h0, add_293795, array_index_293379[0]}) < $signed({1'h0, sel_293797}) ? {add_293795, array_index_293379[0]} : sel_293797;
  assign add_293901 = array_index_293580[11:1] + 11'h347;
  assign sel_293903 = $signed({1'h0, add_293799, array_index_293478[0]}) < $signed({1'h0, sel_293801}) ? {add_293799, array_index_293478[0]} : sel_293801;
  assign add_293905 = array_index_293583[11:1] + 11'h347;
  assign sel_293907 = $signed({1'h0, add_293803, array_index_293481[0]}) < $signed({1'h0, sel_293805}) ? {add_293803, array_index_293481[0]} : sel_293805;
  assign add_293909 = array_index_293682[11:3] + 9'h0bd;
  assign sel_293912 = $signed({1'h0, add_293807, array_index_293580[2:0]}) < $signed({1'h0, sel_293810}) ? {add_293807, array_index_293580[2:0]} : sel_293810;
  assign add_293914 = array_index_293685[11:3] + 9'h0bd;
  assign sel_293917 = $signed({1'h0, add_293812, array_index_293583[2:0]}) < $signed({1'h0, sel_293815}) ? {add_293812, array_index_293583[2:0]} : sel_293815;
  assign add_293919 = array_index_293784[11:1] + 11'h247;
  assign sel_293922 = $signed({1'h0, add_293817, array_index_293682[0]}) < $signed({1'h0, sel_293820}) ? {add_293817, array_index_293682[0]} : sel_293820;
  assign add_293924 = array_index_293787[11:1] + 11'h247;
  assign sel_293927 = $signed({1'h0, add_293822, array_index_293685[0]}) < $signed({1'h0, sel_293825}) ? {add_293822, array_index_293685[0]} : sel_293825;
  assign add_293952 = array_index_293886[11:0] + 12'h247;
  assign sel_293954 = $signed({1'h0, add_293850}) < $signed({1'h0, sel_293852}) ? add_293850 : sel_293852;
  assign add_293957 = array_index_293889[11:0] + 12'h247;
  assign sel_293959 = $signed({1'h0, add_293855}) < $signed({1'h0, sel_293857}) ? add_293855 : sel_293857;
  assign array_index_293988 = set1_unflattened[8'h71];
  assign array_index_293991 = set2_unflattened[8'h71];
  assign add_293995 = array_index_293580[11:1] + 11'h79d;
  assign sel_293997 = $signed({1'h0, add_293893, array_index_293478[0]}) < $signed({1'h0, sel_293895}) ? {add_293893, array_index_293478[0]} : sel_293895;
  assign add_293999 = array_index_293583[11:1] + 11'h79d;
  assign sel_294001 = $signed({1'h0, add_293897, array_index_293481[0]}) < $signed({1'h0, sel_293899}) ? {add_293897, array_index_293481[0]} : sel_293899;
  assign add_294003 = array_index_293682[11:1] + 11'h347;
  assign sel_294005 = $signed({1'h0, add_293901, array_index_293580[0]}) < $signed({1'h0, sel_293903}) ? {add_293901, array_index_293580[0]} : sel_293903;
  assign add_294007 = array_index_293685[11:1] + 11'h347;
  assign sel_294009 = $signed({1'h0, add_293905, array_index_293583[0]}) < $signed({1'h0, sel_293907}) ? {add_293905, array_index_293583[0]} : sel_293907;
  assign add_294011 = array_index_293784[11:3] + 9'h0bd;
  assign sel_294014 = $signed({1'h0, add_293909, array_index_293682[2:0]}) < $signed({1'h0, sel_293912}) ? {add_293909, array_index_293682[2:0]} : sel_293912;
  assign add_294016 = array_index_293787[11:3] + 9'h0bd;
  assign sel_294019 = $signed({1'h0, add_293914, array_index_293685[2:0]}) < $signed({1'h0, sel_293917}) ? {add_293914, array_index_293685[2:0]} : sel_293917;
  assign add_294021 = array_index_293886[11:1] + 11'h247;
  assign sel_294024 = $signed({1'h0, add_293919, array_index_293784[0]}) < $signed({1'h0, sel_293922}) ? {add_293919, array_index_293784[0]} : sel_293922;
  assign add_294026 = array_index_293889[11:1] + 11'h247;
  assign sel_294029 = $signed({1'h0, add_293924, array_index_293787[0]}) < $signed({1'h0, sel_293927}) ? {add_293924, array_index_293787[0]} : sel_293927;
  assign add_294054 = array_index_293988[11:0] + 12'h247;
  assign sel_294056 = $signed({1'h0, add_293952}) < $signed({1'h0, sel_293954}) ? add_293952 : sel_293954;
  assign add_294059 = array_index_293991[11:0] + 12'h247;
  assign sel_294061 = $signed({1'h0, add_293957}) < $signed({1'h0, sel_293959}) ? add_293957 : sel_293959;
  assign array_index_294090 = set1_unflattened[8'h72];
  assign array_index_294093 = set2_unflattened[8'h72];
  assign add_294097 = array_index_293682[11:1] + 11'h79d;
  assign sel_294099 = $signed({1'h0, add_293995, array_index_293580[0]}) < $signed({1'h0, sel_293997}) ? {add_293995, array_index_293580[0]} : sel_293997;
  assign add_294101 = array_index_293685[11:1] + 11'h79d;
  assign sel_294103 = $signed({1'h0, add_293999, array_index_293583[0]}) < $signed({1'h0, sel_294001}) ? {add_293999, array_index_293583[0]} : sel_294001;
  assign add_294105 = array_index_293784[11:1] + 11'h347;
  assign sel_294107 = $signed({1'h0, add_294003, array_index_293682[0]}) < $signed({1'h0, sel_294005}) ? {add_294003, array_index_293682[0]} : sel_294005;
  assign add_294109 = array_index_293787[11:1] + 11'h347;
  assign sel_294111 = $signed({1'h0, add_294007, array_index_293685[0]}) < $signed({1'h0, sel_294009}) ? {add_294007, array_index_293685[0]} : sel_294009;
  assign add_294113 = array_index_293886[11:3] + 9'h0bd;
  assign sel_294116 = $signed({1'h0, add_294011, array_index_293784[2:0]}) < $signed({1'h0, sel_294014}) ? {add_294011, array_index_293784[2:0]} : sel_294014;
  assign add_294118 = array_index_293889[11:3] + 9'h0bd;
  assign sel_294121 = $signed({1'h0, add_294016, array_index_293787[2:0]}) < $signed({1'h0, sel_294019}) ? {add_294016, array_index_293787[2:0]} : sel_294019;
  assign add_294123 = array_index_293988[11:1] + 11'h247;
  assign sel_294126 = $signed({1'h0, add_294021, array_index_293886[0]}) < $signed({1'h0, sel_294024}) ? {add_294021, array_index_293886[0]} : sel_294024;
  assign add_294128 = array_index_293991[11:1] + 11'h247;
  assign sel_294131 = $signed({1'h0, add_294026, array_index_293889[0]}) < $signed({1'h0, sel_294029}) ? {add_294026, array_index_293889[0]} : sel_294029;
  assign add_294156 = array_index_294090[11:0] + 12'h247;
  assign sel_294158 = $signed({1'h0, add_294054}) < $signed({1'h0, sel_294056}) ? add_294054 : sel_294056;
  assign add_294161 = array_index_294093[11:0] + 12'h247;
  assign sel_294163 = $signed({1'h0, add_294059}) < $signed({1'h0, sel_294061}) ? add_294059 : sel_294061;
  assign array_index_294192 = set1_unflattened[8'h73];
  assign array_index_294195 = set2_unflattened[8'h73];
  assign add_294199 = array_index_293784[11:1] + 11'h79d;
  assign sel_294201 = $signed({1'h0, add_294097, array_index_293682[0]}) < $signed({1'h0, sel_294099}) ? {add_294097, array_index_293682[0]} : sel_294099;
  assign add_294203 = array_index_293787[11:1] + 11'h79d;
  assign sel_294205 = $signed({1'h0, add_294101, array_index_293685[0]}) < $signed({1'h0, sel_294103}) ? {add_294101, array_index_293685[0]} : sel_294103;
  assign add_294207 = array_index_293886[11:1] + 11'h347;
  assign sel_294209 = $signed({1'h0, add_294105, array_index_293784[0]}) < $signed({1'h0, sel_294107}) ? {add_294105, array_index_293784[0]} : sel_294107;
  assign add_294211 = array_index_293889[11:1] + 11'h347;
  assign sel_294213 = $signed({1'h0, add_294109, array_index_293787[0]}) < $signed({1'h0, sel_294111}) ? {add_294109, array_index_293787[0]} : sel_294111;
  assign add_294215 = array_index_293988[11:3] + 9'h0bd;
  assign sel_294218 = $signed({1'h0, add_294113, array_index_293886[2:0]}) < $signed({1'h0, sel_294116}) ? {add_294113, array_index_293886[2:0]} : sel_294116;
  assign add_294220 = array_index_293991[11:3] + 9'h0bd;
  assign sel_294223 = $signed({1'h0, add_294118, array_index_293889[2:0]}) < $signed({1'h0, sel_294121}) ? {add_294118, array_index_293889[2:0]} : sel_294121;
  assign add_294225 = array_index_294090[11:1] + 11'h247;
  assign sel_294228 = $signed({1'h0, add_294123, array_index_293988[0]}) < $signed({1'h0, sel_294126}) ? {add_294123, array_index_293988[0]} : sel_294126;
  assign add_294230 = array_index_294093[11:1] + 11'h247;
  assign sel_294233 = $signed({1'h0, add_294128, array_index_293991[0]}) < $signed({1'h0, sel_294131}) ? {add_294128, array_index_293991[0]} : sel_294131;
  assign add_294258 = array_index_294192[11:0] + 12'h247;
  assign sel_294260 = $signed({1'h0, add_294156}) < $signed({1'h0, sel_294158}) ? add_294156 : sel_294158;
  assign add_294263 = array_index_294195[11:0] + 12'h247;
  assign sel_294265 = $signed({1'h0, add_294161}) < $signed({1'h0, sel_294163}) ? add_294161 : sel_294163;
  assign array_index_294294 = set1_unflattened[8'h74];
  assign array_index_294297 = set2_unflattened[8'h74];
  assign add_294301 = array_index_293886[11:1] + 11'h79d;
  assign sel_294303 = $signed({1'h0, add_294199, array_index_293784[0]}) < $signed({1'h0, sel_294201}) ? {add_294199, array_index_293784[0]} : sel_294201;
  assign add_294305 = array_index_293889[11:1] + 11'h79d;
  assign sel_294307 = $signed({1'h0, add_294203, array_index_293787[0]}) < $signed({1'h0, sel_294205}) ? {add_294203, array_index_293787[0]} : sel_294205;
  assign add_294309 = array_index_293988[11:1] + 11'h347;
  assign sel_294311 = $signed({1'h0, add_294207, array_index_293886[0]}) < $signed({1'h0, sel_294209}) ? {add_294207, array_index_293886[0]} : sel_294209;
  assign add_294313 = array_index_293991[11:1] + 11'h347;
  assign sel_294315 = $signed({1'h0, add_294211, array_index_293889[0]}) < $signed({1'h0, sel_294213}) ? {add_294211, array_index_293889[0]} : sel_294213;
  assign add_294317 = array_index_294090[11:3] + 9'h0bd;
  assign sel_294320 = $signed({1'h0, add_294215, array_index_293988[2:0]}) < $signed({1'h0, sel_294218}) ? {add_294215, array_index_293988[2:0]} : sel_294218;
  assign add_294322 = array_index_294093[11:3] + 9'h0bd;
  assign sel_294325 = $signed({1'h0, add_294220, array_index_293991[2:0]}) < $signed({1'h0, sel_294223}) ? {add_294220, array_index_293991[2:0]} : sel_294223;
  assign add_294327 = array_index_294192[11:1] + 11'h247;
  assign sel_294330 = $signed({1'h0, add_294225, array_index_294090[0]}) < $signed({1'h0, sel_294228}) ? {add_294225, array_index_294090[0]} : sel_294228;
  assign add_294332 = array_index_294195[11:1] + 11'h247;
  assign sel_294335 = $signed({1'h0, add_294230, array_index_294093[0]}) < $signed({1'h0, sel_294233}) ? {add_294230, array_index_294093[0]} : sel_294233;
  assign add_294360 = array_index_294294[11:0] + 12'h247;
  assign sel_294362 = $signed({1'h0, add_294258}) < $signed({1'h0, sel_294260}) ? add_294258 : sel_294260;
  assign add_294365 = array_index_294297[11:0] + 12'h247;
  assign sel_294367 = $signed({1'h0, add_294263}) < $signed({1'h0, sel_294265}) ? add_294263 : sel_294265;
  assign array_index_294396 = set1_unflattened[8'h75];
  assign array_index_294399 = set2_unflattened[8'h75];
  assign add_294403 = array_index_293988[11:1] + 11'h79d;
  assign sel_294405 = $signed({1'h0, add_294301, array_index_293886[0]}) < $signed({1'h0, sel_294303}) ? {add_294301, array_index_293886[0]} : sel_294303;
  assign add_294407 = array_index_293991[11:1] + 11'h79d;
  assign sel_294409 = $signed({1'h0, add_294305, array_index_293889[0]}) < $signed({1'h0, sel_294307}) ? {add_294305, array_index_293889[0]} : sel_294307;
  assign add_294411 = array_index_294090[11:1] + 11'h347;
  assign sel_294413 = $signed({1'h0, add_294309, array_index_293988[0]}) < $signed({1'h0, sel_294311}) ? {add_294309, array_index_293988[0]} : sel_294311;
  assign add_294415 = array_index_294093[11:1] + 11'h347;
  assign sel_294417 = $signed({1'h0, add_294313, array_index_293991[0]}) < $signed({1'h0, sel_294315}) ? {add_294313, array_index_293991[0]} : sel_294315;
  assign add_294419 = array_index_294192[11:3] + 9'h0bd;
  assign sel_294422 = $signed({1'h0, add_294317, array_index_294090[2:0]}) < $signed({1'h0, sel_294320}) ? {add_294317, array_index_294090[2:0]} : sel_294320;
  assign add_294424 = array_index_294195[11:3] + 9'h0bd;
  assign sel_294427 = $signed({1'h0, add_294322, array_index_294093[2:0]}) < $signed({1'h0, sel_294325}) ? {add_294322, array_index_294093[2:0]} : sel_294325;
  assign add_294429 = array_index_294294[11:1] + 11'h247;
  assign sel_294432 = $signed({1'h0, add_294327, array_index_294192[0]}) < $signed({1'h0, sel_294330}) ? {add_294327, array_index_294192[0]} : sel_294330;
  assign add_294434 = array_index_294297[11:1] + 11'h247;
  assign sel_294437 = $signed({1'h0, add_294332, array_index_294195[0]}) < $signed({1'h0, sel_294335}) ? {add_294332, array_index_294195[0]} : sel_294335;
  assign add_294462 = array_index_294396[11:0] + 12'h247;
  assign sel_294464 = $signed({1'h0, add_294360}) < $signed({1'h0, sel_294362}) ? add_294360 : sel_294362;
  assign add_294467 = array_index_294399[11:0] + 12'h247;
  assign sel_294469 = $signed({1'h0, add_294365}) < $signed({1'h0, sel_294367}) ? add_294365 : sel_294367;
  assign array_index_294498 = set1_unflattened[8'h76];
  assign array_index_294501 = set2_unflattened[8'h76];
  assign add_294505 = array_index_294090[11:1] + 11'h79d;
  assign sel_294507 = $signed({1'h0, add_294403, array_index_293988[0]}) < $signed({1'h0, sel_294405}) ? {add_294403, array_index_293988[0]} : sel_294405;
  assign add_294509 = array_index_294093[11:1] + 11'h79d;
  assign sel_294511 = $signed({1'h0, add_294407, array_index_293991[0]}) < $signed({1'h0, sel_294409}) ? {add_294407, array_index_293991[0]} : sel_294409;
  assign add_294513 = array_index_294192[11:1] + 11'h347;
  assign sel_294515 = $signed({1'h0, add_294411, array_index_294090[0]}) < $signed({1'h0, sel_294413}) ? {add_294411, array_index_294090[0]} : sel_294413;
  assign add_294517 = array_index_294195[11:1] + 11'h347;
  assign sel_294519 = $signed({1'h0, add_294415, array_index_294093[0]}) < $signed({1'h0, sel_294417}) ? {add_294415, array_index_294093[0]} : sel_294417;
  assign add_294521 = array_index_294294[11:3] + 9'h0bd;
  assign sel_294524 = $signed({1'h0, add_294419, array_index_294192[2:0]}) < $signed({1'h0, sel_294422}) ? {add_294419, array_index_294192[2:0]} : sel_294422;
  assign add_294526 = array_index_294297[11:3] + 9'h0bd;
  assign sel_294529 = $signed({1'h0, add_294424, array_index_294195[2:0]}) < $signed({1'h0, sel_294427}) ? {add_294424, array_index_294195[2:0]} : sel_294427;
  assign add_294531 = array_index_294396[11:1] + 11'h247;
  assign sel_294534 = $signed({1'h0, add_294429, array_index_294294[0]}) < $signed({1'h0, sel_294432}) ? {add_294429, array_index_294294[0]} : sel_294432;
  assign add_294536 = array_index_294399[11:1] + 11'h247;
  assign sel_294539 = $signed({1'h0, add_294434, array_index_294297[0]}) < $signed({1'h0, sel_294437}) ? {add_294434, array_index_294297[0]} : sel_294437;
  assign add_294564 = array_index_294498[11:0] + 12'h247;
  assign sel_294566 = $signed({1'h0, add_294462}) < $signed({1'h0, sel_294464}) ? add_294462 : sel_294464;
  assign add_294569 = array_index_294501[11:0] + 12'h247;
  assign sel_294571 = $signed({1'h0, add_294467}) < $signed({1'h0, sel_294469}) ? add_294467 : sel_294469;
  assign array_index_294600 = set1_unflattened[8'h77];
  assign array_index_294603 = set2_unflattened[8'h77];
  assign add_294607 = array_index_294192[11:1] + 11'h79d;
  assign sel_294609 = $signed({1'h0, add_294505, array_index_294090[0]}) < $signed({1'h0, sel_294507}) ? {add_294505, array_index_294090[0]} : sel_294507;
  assign add_294611 = array_index_294195[11:1] + 11'h79d;
  assign sel_294613 = $signed({1'h0, add_294509, array_index_294093[0]}) < $signed({1'h0, sel_294511}) ? {add_294509, array_index_294093[0]} : sel_294511;
  assign add_294615 = array_index_294294[11:1] + 11'h347;
  assign sel_294617 = $signed({1'h0, add_294513, array_index_294192[0]}) < $signed({1'h0, sel_294515}) ? {add_294513, array_index_294192[0]} : sel_294515;
  assign add_294619 = array_index_294297[11:1] + 11'h347;
  assign sel_294621 = $signed({1'h0, add_294517, array_index_294195[0]}) < $signed({1'h0, sel_294519}) ? {add_294517, array_index_294195[0]} : sel_294519;
  assign add_294623 = array_index_294396[11:3] + 9'h0bd;
  assign sel_294626 = $signed({1'h0, add_294521, array_index_294294[2:0]}) < $signed({1'h0, sel_294524}) ? {add_294521, array_index_294294[2:0]} : sel_294524;
  assign add_294628 = array_index_294399[11:3] + 9'h0bd;
  assign sel_294631 = $signed({1'h0, add_294526, array_index_294297[2:0]}) < $signed({1'h0, sel_294529}) ? {add_294526, array_index_294297[2:0]} : sel_294529;
  assign add_294633 = array_index_294498[11:1] + 11'h247;
  assign sel_294636 = $signed({1'h0, add_294531, array_index_294396[0]}) < $signed({1'h0, sel_294534}) ? {add_294531, array_index_294396[0]} : sel_294534;
  assign add_294638 = array_index_294501[11:1] + 11'h247;
  assign sel_294641 = $signed({1'h0, add_294536, array_index_294399[0]}) < $signed({1'h0, sel_294539}) ? {add_294536, array_index_294399[0]} : sel_294539;
  assign add_294666 = array_index_294600[11:0] + 12'h247;
  assign sel_294668 = $signed({1'h0, add_294564}) < $signed({1'h0, sel_294566}) ? add_294564 : sel_294566;
  assign add_294671 = array_index_294603[11:0] + 12'h247;
  assign sel_294673 = $signed({1'h0, add_294569}) < $signed({1'h0, sel_294571}) ? add_294569 : sel_294571;
  assign array_index_294702 = set1_unflattened[8'h78];
  assign array_index_294705 = set2_unflattened[8'h78];
  assign add_294709 = array_index_294294[11:1] + 11'h79d;
  assign sel_294711 = $signed({1'h0, add_294607, array_index_294192[0]}) < $signed({1'h0, sel_294609}) ? {add_294607, array_index_294192[0]} : sel_294609;
  assign add_294713 = array_index_294297[11:1] + 11'h79d;
  assign sel_294715 = $signed({1'h0, add_294611, array_index_294195[0]}) < $signed({1'h0, sel_294613}) ? {add_294611, array_index_294195[0]} : sel_294613;
  assign add_294717 = array_index_294396[11:1] + 11'h347;
  assign sel_294719 = $signed({1'h0, add_294615, array_index_294294[0]}) < $signed({1'h0, sel_294617}) ? {add_294615, array_index_294294[0]} : sel_294617;
  assign add_294721 = array_index_294399[11:1] + 11'h347;
  assign sel_294723 = $signed({1'h0, add_294619, array_index_294297[0]}) < $signed({1'h0, sel_294621}) ? {add_294619, array_index_294297[0]} : sel_294621;
  assign add_294725 = array_index_294498[11:3] + 9'h0bd;
  assign sel_294728 = $signed({1'h0, add_294623, array_index_294396[2:0]}) < $signed({1'h0, sel_294626}) ? {add_294623, array_index_294396[2:0]} : sel_294626;
  assign add_294730 = array_index_294501[11:3] + 9'h0bd;
  assign sel_294733 = $signed({1'h0, add_294628, array_index_294399[2:0]}) < $signed({1'h0, sel_294631}) ? {add_294628, array_index_294399[2:0]} : sel_294631;
  assign add_294735 = array_index_294600[11:1] + 11'h247;
  assign sel_294738 = $signed({1'h0, add_294633, array_index_294498[0]}) < $signed({1'h0, sel_294636}) ? {add_294633, array_index_294498[0]} : sel_294636;
  assign add_294740 = array_index_294603[11:1] + 11'h247;
  assign sel_294743 = $signed({1'h0, add_294638, array_index_294501[0]}) < $signed({1'h0, sel_294641}) ? {add_294638, array_index_294501[0]} : sel_294641;
  assign add_294768 = array_index_294702[11:0] + 12'h247;
  assign sel_294770 = $signed({1'h0, add_294666}) < $signed({1'h0, sel_294668}) ? add_294666 : sel_294668;
  assign add_294773 = array_index_294705[11:0] + 12'h247;
  assign sel_294775 = $signed({1'h0, add_294671}) < $signed({1'h0, sel_294673}) ? add_294671 : sel_294673;
  assign array_index_294804 = set1_unflattened[8'h79];
  assign array_index_294807 = set2_unflattened[8'h79];
  assign add_294811 = array_index_294396[11:1] + 11'h79d;
  assign sel_294813 = $signed({1'h0, add_294709, array_index_294294[0]}) < $signed({1'h0, sel_294711}) ? {add_294709, array_index_294294[0]} : sel_294711;
  assign add_294815 = array_index_294399[11:1] + 11'h79d;
  assign sel_294817 = $signed({1'h0, add_294713, array_index_294297[0]}) < $signed({1'h0, sel_294715}) ? {add_294713, array_index_294297[0]} : sel_294715;
  assign add_294819 = array_index_294498[11:1] + 11'h347;
  assign sel_294821 = $signed({1'h0, add_294717, array_index_294396[0]}) < $signed({1'h0, sel_294719}) ? {add_294717, array_index_294396[0]} : sel_294719;
  assign add_294823 = array_index_294501[11:1] + 11'h347;
  assign sel_294825 = $signed({1'h0, add_294721, array_index_294399[0]}) < $signed({1'h0, sel_294723}) ? {add_294721, array_index_294399[0]} : sel_294723;
  assign add_294827 = array_index_294600[11:3] + 9'h0bd;
  assign sel_294830 = $signed({1'h0, add_294725, array_index_294498[2:0]}) < $signed({1'h0, sel_294728}) ? {add_294725, array_index_294498[2:0]} : sel_294728;
  assign add_294832 = array_index_294603[11:3] + 9'h0bd;
  assign sel_294835 = $signed({1'h0, add_294730, array_index_294501[2:0]}) < $signed({1'h0, sel_294733}) ? {add_294730, array_index_294501[2:0]} : sel_294733;
  assign add_294837 = array_index_294702[11:1] + 11'h247;
  assign sel_294840 = $signed({1'h0, add_294735, array_index_294600[0]}) < $signed({1'h0, sel_294738}) ? {add_294735, array_index_294600[0]} : sel_294738;
  assign add_294842 = array_index_294705[11:1] + 11'h247;
  assign sel_294845 = $signed({1'h0, add_294740, array_index_294603[0]}) < $signed({1'h0, sel_294743}) ? {add_294740, array_index_294603[0]} : sel_294743;
  assign add_294870 = array_index_294804[11:0] + 12'h247;
  assign sel_294872 = $signed({1'h0, add_294768}) < $signed({1'h0, sel_294770}) ? add_294768 : sel_294770;
  assign add_294875 = array_index_294807[11:0] + 12'h247;
  assign sel_294877 = $signed({1'h0, add_294773}) < $signed({1'h0, sel_294775}) ? add_294773 : sel_294775;
  assign array_index_294906 = set1_unflattened[8'h7a];
  assign array_index_294909 = set2_unflattened[8'h7a];
  assign add_294913 = array_index_294498[11:1] + 11'h79d;
  assign sel_294915 = $signed({1'h0, add_294811, array_index_294396[0]}) < $signed({1'h0, sel_294813}) ? {add_294811, array_index_294396[0]} : sel_294813;
  assign add_294917 = array_index_294501[11:1] + 11'h79d;
  assign sel_294919 = $signed({1'h0, add_294815, array_index_294399[0]}) < $signed({1'h0, sel_294817}) ? {add_294815, array_index_294399[0]} : sel_294817;
  assign add_294921 = array_index_294600[11:1] + 11'h347;
  assign sel_294923 = $signed({1'h0, add_294819, array_index_294498[0]}) < $signed({1'h0, sel_294821}) ? {add_294819, array_index_294498[0]} : sel_294821;
  assign add_294925 = array_index_294603[11:1] + 11'h347;
  assign sel_294927 = $signed({1'h0, add_294823, array_index_294501[0]}) < $signed({1'h0, sel_294825}) ? {add_294823, array_index_294501[0]} : sel_294825;
  assign add_294929 = array_index_294702[11:3] + 9'h0bd;
  assign sel_294932 = $signed({1'h0, add_294827, array_index_294600[2:0]}) < $signed({1'h0, sel_294830}) ? {add_294827, array_index_294600[2:0]} : sel_294830;
  assign add_294934 = array_index_294705[11:3] + 9'h0bd;
  assign sel_294937 = $signed({1'h0, add_294832, array_index_294603[2:0]}) < $signed({1'h0, sel_294835}) ? {add_294832, array_index_294603[2:0]} : sel_294835;
  assign add_294939 = array_index_294804[11:1] + 11'h247;
  assign sel_294942 = $signed({1'h0, add_294837, array_index_294702[0]}) < $signed({1'h0, sel_294840}) ? {add_294837, array_index_294702[0]} : sel_294840;
  assign add_294944 = array_index_294807[11:1] + 11'h247;
  assign sel_294947 = $signed({1'h0, add_294842, array_index_294705[0]}) < $signed({1'h0, sel_294845}) ? {add_294842, array_index_294705[0]} : sel_294845;
  assign add_294972 = array_index_294906[11:0] + 12'h247;
  assign sel_294974 = $signed({1'h0, add_294870}) < $signed({1'h0, sel_294872}) ? add_294870 : sel_294872;
  assign add_294977 = array_index_294909[11:0] + 12'h247;
  assign sel_294979 = $signed({1'h0, add_294875}) < $signed({1'h0, sel_294877}) ? add_294875 : sel_294877;
  assign array_index_295008 = set1_unflattened[8'h7b];
  assign array_index_295011 = set2_unflattened[8'h7b];
  assign add_295015 = array_index_294600[11:1] + 11'h79d;
  assign sel_295017 = $signed({1'h0, add_294913, array_index_294498[0]}) < $signed({1'h0, sel_294915}) ? {add_294913, array_index_294498[0]} : sel_294915;
  assign add_295019 = array_index_294603[11:1] + 11'h79d;
  assign sel_295021 = $signed({1'h0, add_294917, array_index_294501[0]}) < $signed({1'h0, sel_294919}) ? {add_294917, array_index_294501[0]} : sel_294919;
  assign add_295023 = array_index_294702[11:1] + 11'h347;
  assign sel_295025 = $signed({1'h0, add_294921, array_index_294600[0]}) < $signed({1'h0, sel_294923}) ? {add_294921, array_index_294600[0]} : sel_294923;
  assign add_295027 = array_index_294705[11:1] + 11'h347;
  assign sel_295029 = $signed({1'h0, add_294925, array_index_294603[0]}) < $signed({1'h0, sel_294927}) ? {add_294925, array_index_294603[0]} : sel_294927;
  assign add_295031 = array_index_294804[11:3] + 9'h0bd;
  assign sel_295034 = $signed({1'h0, add_294929, array_index_294702[2:0]}) < $signed({1'h0, sel_294932}) ? {add_294929, array_index_294702[2:0]} : sel_294932;
  assign add_295036 = array_index_294807[11:3] + 9'h0bd;
  assign sel_295039 = $signed({1'h0, add_294934, array_index_294705[2:0]}) < $signed({1'h0, sel_294937}) ? {add_294934, array_index_294705[2:0]} : sel_294937;
  assign add_295041 = array_index_294906[11:1] + 11'h247;
  assign sel_295044 = $signed({1'h0, add_294939, array_index_294804[0]}) < $signed({1'h0, sel_294942}) ? {add_294939, array_index_294804[0]} : sel_294942;
  assign add_295046 = array_index_294909[11:1] + 11'h247;
  assign sel_295049 = $signed({1'h0, add_294944, array_index_294807[0]}) < $signed({1'h0, sel_294947}) ? {add_294944, array_index_294807[0]} : sel_294947;
  assign add_295074 = array_index_295008[11:0] + 12'h247;
  assign sel_295076 = $signed({1'h0, add_294972}) < $signed({1'h0, sel_294974}) ? add_294972 : sel_294974;
  assign add_295079 = array_index_295011[11:0] + 12'h247;
  assign sel_295081 = $signed({1'h0, add_294977}) < $signed({1'h0, sel_294979}) ? add_294977 : sel_294979;
  assign array_index_295110 = set1_unflattened[8'h7c];
  assign array_index_295113 = set2_unflattened[8'h7c];
  assign add_295117 = array_index_294702[11:1] + 11'h79d;
  assign sel_295119 = $signed({1'h0, add_295015, array_index_294600[0]}) < $signed({1'h0, sel_295017}) ? {add_295015, array_index_294600[0]} : sel_295017;
  assign add_295121 = array_index_294705[11:1] + 11'h79d;
  assign sel_295123 = $signed({1'h0, add_295019, array_index_294603[0]}) < $signed({1'h0, sel_295021}) ? {add_295019, array_index_294603[0]} : sel_295021;
  assign add_295125 = array_index_294804[11:1] + 11'h347;
  assign sel_295127 = $signed({1'h0, add_295023, array_index_294702[0]}) < $signed({1'h0, sel_295025}) ? {add_295023, array_index_294702[0]} : sel_295025;
  assign add_295129 = array_index_294807[11:1] + 11'h347;
  assign sel_295131 = $signed({1'h0, add_295027, array_index_294705[0]}) < $signed({1'h0, sel_295029}) ? {add_295027, array_index_294705[0]} : sel_295029;
  assign add_295133 = array_index_294906[11:3] + 9'h0bd;
  assign sel_295136 = $signed({1'h0, add_295031, array_index_294804[2:0]}) < $signed({1'h0, sel_295034}) ? {add_295031, array_index_294804[2:0]} : sel_295034;
  assign add_295138 = array_index_294909[11:3] + 9'h0bd;
  assign sel_295141 = $signed({1'h0, add_295036, array_index_294807[2:0]}) < $signed({1'h0, sel_295039}) ? {add_295036, array_index_294807[2:0]} : sel_295039;
  assign add_295143 = array_index_295008[11:1] + 11'h247;
  assign sel_295146 = $signed({1'h0, add_295041, array_index_294906[0]}) < $signed({1'h0, sel_295044}) ? {add_295041, array_index_294906[0]} : sel_295044;
  assign add_295148 = array_index_295011[11:1] + 11'h247;
  assign sel_295151 = $signed({1'h0, add_295046, array_index_294909[0]}) < $signed({1'h0, sel_295049}) ? {add_295046, array_index_294909[0]} : sel_295049;
  assign add_295176 = array_index_295110[11:0] + 12'h247;
  assign sel_295178 = $signed({1'h0, add_295074}) < $signed({1'h0, sel_295076}) ? add_295074 : sel_295076;
  assign add_295181 = array_index_295113[11:0] + 12'h247;
  assign sel_295183 = $signed({1'h0, add_295079}) < $signed({1'h0, sel_295081}) ? add_295079 : sel_295081;
  assign array_index_295212 = set1_unflattened[8'h7d];
  assign array_index_295215 = set2_unflattened[8'h7d];
  assign add_295219 = array_index_294804[11:1] + 11'h79d;
  assign sel_295221 = $signed({1'h0, add_295117, array_index_294702[0]}) < $signed({1'h0, sel_295119}) ? {add_295117, array_index_294702[0]} : sel_295119;
  assign add_295223 = array_index_294807[11:1] + 11'h79d;
  assign sel_295225 = $signed({1'h0, add_295121, array_index_294705[0]}) < $signed({1'h0, sel_295123}) ? {add_295121, array_index_294705[0]} : sel_295123;
  assign add_295227 = array_index_294906[11:1] + 11'h347;
  assign sel_295229 = $signed({1'h0, add_295125, array_index_294804[0]}) < $signed({1'h0, sel_295127}) ? {add_295125, array_index_294804[0]} : sel_295127;
  assign add_295231 = array_index_294909[11:1] + 11'h347;
  assign sel_295233 = $signed({1'h0, add_295129, array_index_294807[0]}) < $signed({1'h0, sel_295131}) ? {add_295129, array_index_294807[0]} : sel_295131;
  assign add_295235 = array_index_295008[11:3] + 9'h0bd;
  assign sel_295238 = $signed({1'h0, add_295133, array_index_294906[2:0]}) < $signed({1'h0, sel_295136}) ? {add_295133, array_index_294906[2:0]} : sel_295136;
  assign add_295240 = array_index_295011[11:3] + 9'h0bd;
  assign sel_295243 = $signed({1'h0, add_295138, array_index_294909[2:0]}) < $signed({1'h0, sel_295141}) ? {add_295138, array_index_294909[2:0]} : sel_295141;
  assign add_295245 = array_index_295110[11:1] + 11'h247;
  assign sel_295248 = $signed({1'h0, add_295143, array_index_295008[0]}) < $signed({1'h0, sel_295146}) ? {add_295143, array_index_295008[0]} : sel_295146;
  assign add_295250 = array_index_295113[11:1] + 11'h247;
  assign sel_295253 = $signed({1'h0, add_295148, array_index_295011[0]}) < $signed({1'h0, sel_295151}) ? {add_295148, array_index_295011[0]} : sel_295151;
  assign add_295278 = array_index_295212[11:0] + 12'h247;
  assign sel_295280 = $signed({1'h0, add_295176}) < $signed({1'h0, sel_295178}) ? add_295176 : sel_295178;
  assign add_295283 = array_index_295215[11:0] + 12'h247;
  assign sel_295285 = $signed({1'h0, add_295181}) < $signed({1'h0, sel_295183}) ? add_295181 : sel_295183;
  assign array_index_295314 = set1_unflattened[8'h7e];
  assign array_index_295317 = set2_unflattened[8'h7e];
  assign add_295321 = array_index_294906[11:1] + 11'h79d;
  assign sel_295323 = $signed({1'h0, add_295219, array_index_294804[0]}) < $signed({1'h0, sel_295221}) ? {add_295219, array_index_294804[0]} : sel_295221;
  assign add_295325 = array_index_294909[11:1] + 11'h79d;
  assign sel_295327 = $signed({1'h0, add_295223, array_index_294807[0]}) < $signed({1'h0, sel_295225}) ? {add_295223, array_index_294807[0]} : sel_295225;
  assign add_295329 = array_index_295008[11:1] + 11'h347;
  assign sel_295331 = $signed({1'h0, add_295227, array_index_294906[0]}) < $signed({1'h0, sel_295229}) ? {add_295227, array_index_294906[0]} : sel_295229;
  assign add_295333 = array_index_295011[11:1] + 11'h347;
  assign sel_295335 = $signed({1'h0, add_295231, array_index_294909[0]}) < $signed({1'h0, sel_295233}) ? {add_295231, array_index_294909[0]} : sel_295233;
  assign add_295337 = array_index_295110[11:3] + 9'h0bd;
  assign sel_295340 = $signed({1'h0, add_295235, array_index_295008[2:0]}) < $signed({1'h0, sel_295238}) ? {add_295235, array_index_295008[2:0]} : sel_295238;
  assign add_295342 = array_index_295113[11:3] + 9'h0bd;
  assign sel_295345 = $signed({1'h0, add_295240, array_index_295011[2:0]}) < $signed({1'h0, sel_295243}) ? {add_295240, array_index_295011[2:0]} : sel_295243;
  assign add_295347 = array_index_295212[11:1] + 11'h247;
  assign sel_295350 = $signed({1'h0, add_295245, array_index_295110[0]}) < $signed({1'h0, sel_295248}) ? {add_295245, array_index_295110[0]} : sel_295248;
  assign add_295352 = array_index_295215[11:1] + 11'h247;
  assign sel_295355 = $signed({1'h0, add_295250, array_index_295113[0]}) < $signed({1'h0, sel_295253}) ? {add_295250, array_index_295113[0]} : sel_295253;
  assign add_295380 = array_index_295314[11:0] + 12'h247;
  assign sel_295382 = $signed({1'h0, add_295278}) < $signed({1'h0, sel_295280}) ? add_295278 : sel_295280;
  assign add_295385 = array_index_295317[11:0] + 12'h247;
  assign sel_295387 = $signed({1'h0, add_295283}) < $signed({1'h0, sel_295285}) ? add_295283 : sel_295285;
  assign array_index_295416 = set1_unflattened[8'h7f];
  assign array_index_295419 = set2_unflattened[8'h7f];
  assign add_295423 = array_index_295008[11:1] + 11'h79d;
  assign sel_295425 = $signed({1'h0, add_295321, array_index_294906[0]}) < $signed({1'h0, sel_295323}) ? {add_295321, array_index_294906[0]} : sel_295323;
  assign add_295427 = array_index_295011[11:1] + 11'h79d;
  assign sel_295429 = $signed({1'h0, add_295325, array_index_294909[0]}) < $signed({1'h0, sel_295327}) ? {add_295325, array_index_294909[0]} : sel_295327;
  assign add_295431 = array_index_295110[11:1] + 11'h347;
  assign sel_295433 = $signed({1'h0, add_295329, array_index_295008[0]}) < $signed({1'h0, sel_295331}) ? {add_295329, array_index_295008[0]} : sel_295331;
  assign add_295435 = array_index_295113[11:1] + 11'h347;
  assign sel_295437 = $signed({1'h0, add_295333, array_index_295011[0]}) < $signed({1'h0, sel_295335}) ? {add_295333, array_index_295011[0]} : sel_295335;
  assign add_295439 = array_index_295212[11:3] + 9'h0bd;
  assign sel_295442 = $signed({1'h0, add_295337, array_index_295110[2:0]}) < $signed({1'h0, sel_295340}) ? {add_295337, array_index_295110[2:0]} : sel_295340;
  assign add_295444 = array_index_295215[11:3] + 9'h0bd;
  assign sel_295447 = $signed({1'h0, add_295342, array_index_295113[2:0]}) < $signed({1'h0, sel_295345}) ? {add_295342, array_index_295113[2:0]} : sel_295345;
  assign add_295449 = array_index_295314[11:1] + 11'h247;
  assign sel_295452 = $signed({1'h0, add_295347, array_index_295212[0]}) < $signed({1'h0, sel_295350}) ? {add_295347, array_index_295212[0]} : sel_295350;
  assign add_295454 = array_index_295317[11:1] + 11'h247;
  assign sel_295457 = $signed({1'h0, add_295352, array_index_295215[0]}) < $signed({1'h0, sel_295355}) ? {add_295352, array_index_295215[0]} : sel_295355;
  assign add_295482 = array_index_295416[11:0] + 12'h247;
  assign sel_295484 = $signed({1'h0, add_295380}) < $signed({1'h0, sel_295382}) ? add_295380 : sel_295382;
  assign add_295487 = array_index_295419[11:0] + 12'h247;
  assign sel_295489 = $signed({1'h0, add_295385}) < $signed({1'h0, sel_295387}) ? add_295385 : sel_295387;
  assign array_index_295518 = set1_unflattened[8'h80];
  assign array_index_295521 = set2_unflattened[8'h80];
  assign add_295525 = array_index_295110[11:1] + 11'h79d;
  assign sel_295527 = $signed({1'h0, add_295423, array_index_295008[0]}) < $signed({1'h0, sel_295425}) ? {add_295423, array_index_295008[0]} : sel_295425;
  assign add_295529 = array_index_295113[11:1] + 11'h79d;
  assign sel_295531 = $signed({1'h0, add_295427, array_index_295011[0]}) < $signed({1'h0, sel_295429}) ? {add_295427, array_index_295011[0]} : sel_295429;
  assign add_295533 = array_index_295212[11:1] + 11'h347;
  assign sel_295535 = $signed({1'h0, add_295431, array_index_295110[0]}) < $signed({1'h0, sel_295433}) ? {add_295431, array_index_295110[0]} : sel_295433;
  assign add_295537 = array_index_295215[11:1] + 11'h347;
  assign sel_295539 = $signed({1'h0, add_295435, array_index_295113[0]}) < $signed({1'h0, sel_295437}) ? {add_295435, array_index_295113[0]} : sel_295437;
  assign add_295541 = array_index_295314[11:3] + 9'h0bd;
  assign sel_295544 = $signed({1'h0, add_295439, array_index_295212[2:0]}) < $signed({1'h0, sel_295442}) ? {add_295439, array_index_295212[2:0]} : sel_295442;
  assign add_295546 = array_index_295317[11:3] + 9'h0bd;
  assign sel_295549 = $signed({1'h0, add_295444, array_index_295215[2:0]}) < $signed({1'h0, sel_295447}) ? {add_295444, array_index_295215[2:0]} : sel_295447;
  assign add_295551 = array_index_295416[11:1] + 11'h247;
  assign sel_295554 = $signed({1'h0, add_295449, array_index_295314[0]}) < $signed({1'h0, sel_295452}) ? {add_295449, array_index_295314[0]} : sel_295452;
  assign add_295556 = array_index_295419[11:1] + 11'h247;
  assign sel_295559 = $signed({1'h0, add_295454, array_index_295317[0]}) < $signed({1'h0, sel_295457}) ? {add_295454, array_index_295317[0]} : sel_295457;
  assign add_295584 = array_index_295518[11:0] + 12'h247;
  assign sel_295586 = $signed({1'h0, add_295482}) < $signed({1'h0, sel_295484}) ? add_295482 : sel_295484;
  assign add_295589 = array_index_295521[11:0] + 12'h247;
  assign sel_295591 = $signed({1'h0, add_295487}) < $signed({1'h0, sel_295489}) ? add_295487 : sel_295489;
  assign array_index_295620 = set1_unflattened[8'h81];
  assign array_index_295623 = set2_unflattened[8'h81];
  assign add_295627 = array_index_295212[11:1] + 11'h79d;
  assign sel_295629 = $signed({1'h0, add_295525, array_index_295110[0]}) < $signed({1'h0, sel_295527}) ? {add_295525, array_index_295110[0]} : sel_295527;
  assign add_295631 = array_index_295215[11:1] + 11'h79d;
  assign sel_295633 = $signed({1'h0, add_295529, array_index_295113[0]}) < $signed({1'h0, sel_295531}) ? {add_295529, array_index_295113[0]} : sel_295531;
  assign add_295635 = array_index_295314[11:1] + 11'h347;
  assign sel_295637 = $signed({1'h0, add_295533, array_index_295212[0]}) < $signed({1'h0, sel_295535}) ? {add_295533, array_index_295212[0]} : sel_295535;
  assign add_295639 = array_index_295317[11:1] + 11'h347;
  assign sel_295641 = $signed({1'h0, add_295537, array_index_295215[0]}) < $signed({1'h0, sel_295539}) ? {add_295537, array_index_295215[0]} : sel_295539;
  assign add_295643 = array_index_295416[11:3] + 9'h0bd;
  assign sel_295646 = $signed({1'h0, add_295541, array_index_295314[2:0]}) < $signed({1'h0, sel_295544}) ? {add_295541, array_index_295314[2:0]} : sel_295544;
  assign add_295648 = array_index_295419[11:3] + 9'h0bd;
  assign sel_295651 = $signed({1'h0, add_295546, array_index_295317[2:0]}) < $signed({1'h0, sel_295549}) ? {add_295546, array_index_295317[2:0]} : sel_295549;
  assign add_295653 = array_index_295518[11:1] + 11'h247;
  assign sel_295656 = $signed({1'h0, add_295551, array_index_295416[0]}) < $signed({1'h0, sel_295554}) ? {add_295551, array_index_295416[0]} : sel_295554;
  assign add_295658 = array_index_295521[11:1] + 11'h247;
  assign sel_295661 = $signed({1'h0, add_295556, array_index_295419[0]}) < $signed({1'h0, sel_295559}) ? {add_295556, array_index_295419[0]} : sel_295559;
  assign add_295686 = array_index_295620[11:0] + 12'h247;
  assign sel_295688 = $signed({1'h0, add_295584}) < $signed({1'h0, sel_295586}) ? add_295584 : sel_295586;
  assign add_295691 = array_index_295623[11:0] + 12'h247;
  assign sel_295693 = $signed({1'h0, add_295589}) < $signed({1'h0, sel_295591}) ? add_295589 : sel_295591;
  assign array_index_295722 = set1_unflattened[8'h82];
  assign array_index_295725 = set2_unflattened[8'h82];
  assign add_295729 = array_index_295314[11:1] + 11'h79d;
  assign sel_295731 = $signed({1'h0, add_295627, array_index_295212[0]}) < $signed({1'h0, sel_295629}) ? {add_295627, array_index_295212[0]} : sel_295629;
  assign add_295733 = array_index_295317[11:1] + 11'h79d;
  assign sel_295735 = $signed({1'h0, add_295631, array_index_295215[0]}) < $signed({1'h0, sel_295633}) ? {add_295631, array_index_295215[0]} : sel_295633;
  assign add_295737 = array_index_295416[11:1] + 11'h347;
  assign sel_295739 = $signed({1'h0, add_295635, array_index_295314[0]}) < $signed({1'h0, sel_295637}) ? {add_295635, array_index_295314[0]} : sel_295637;
  assign add_295741 = array_index_295419[11:1] + 11'h347;
  assign sel_295743 = $signed({1'h0, add_295639, array_index_295317[0]}) < $signed({1'h0, sel_295641}) ? {add_295639, array_index_295317[0]} : sel_295641;
  assign add_295745 = array_index_295518[11:3] + 9'h0bd;
  assign sel_295748 = $signed({1'h0, add_295643, array_index_295416[2:0]}) < $signed({1'h0, sel_295646}) ? {add_295643, array_index_295416[2:0]} : sel_295646;
  assign add_295750 = array_index_295521[11:3] + 9'h0bd;
  assign sel_295753 = $signed({1'h0, add_295648, array_index_295419[2:0]}) < $signed({1'h0, sel_295651}) ? {add_295648, array_index_295419[2:0]} : sel_295651;
  assign add_295755 = array_index_295620[11:1] + 11'h247;
  assign sel_295758 = $signed({1'h0, add_295653, array_index_295518[0]}) < $signed({1'h0, sel_295656}) ? {add_295653, array_index_295518[0]} : sel_295656;
  assign add_295760 = array_index_295623[11:1] + 11'h247;
  assign sel_295763 = $signed({1'h0, add_295658, array_index_295521[0]}) < $signed({1'h0, sel_295661}) ? {add_295658, array_index_295521[0]} : sel_295661;
  assign add_295788 = array_index_295722[11:0] + 12'h247;
  assign sel_295790 = $signed({1'h0, add_295686}) < $signed({1'h0, sel_295688}) ? add_295686 : sel_295688;
  assign add_295793 = array_index_295725[11:0] + 12'h247;
  assign sel_295795 = $signed({1'h0, add_295691}) < $signed({1'h0, sel_295693}) ? add_295691 : sel_295693;
  assign array_index_295824 = set1_unflattened[8'h83];
  assign array_index_295827 = set2_unflattened[8'h83];
  assign add_295831 = array_index_295416[11:1] + 11'h79d;
  assign sel_295833 = $signed({1'h0, add_295729, array_index_295314[0]}) < $signed({1'h0, sel_295731}) ? {add_295729, array_index_295314[0]} : sel_295731;
  assign add_295835 = array_index_295419[11:1] + 11'h79d;
  assign sel_295837 = $signed({1'h0, add_295733, array_index_295317[0]}) < $signed({1'h0, sel_295735}) ? {add_295733, array_index_295317[0]} : sel_295735;
  assign add_295839 = array_index_295518[11:1] + 11'h347;
  assign sel_295841 = $signed({1'h0, add_295737, array_index_295416[0]}) < $signed({1'h0, sel_295739}) ? {add_295737, array_index_295416[0]} : sel_295739;
  assign add_295843 = array_index_295521[11:1] + 11'h347;
  assign sel_295845 = $signed({1'h0, add_295741, array_index_295419[0]}) < $signed({1'h0, sel_295743}) ? {add_295741, array_index_295419[0]} : sel_295743;
  assign add_295847 = array_index_295620[11:3] + 9'h0bd;
  assign sel_295850 = $signed({1'h0, add_295745, array_index_295518[2:0]}) < $signed({1'h0, sel_295748}) ? {add_295745, array_index_295518[2:0]} : sel_295748;
  assign add_295852 = array_index_295623[11:3] + 9'h0bd;
  assign sel_295855 = $signed({1'h0, add_295750, array_index_295521[2:0]}) < $signed({1'h0, sel_295753}) ? {add_295750, array_index_295521[2:0]} : sel_295753;
  assign add_295857 = array_index_295722[11:1] + 11'h247;
  assign sel_295860 = $signed({1'h0, add_295755, array_index_295620[0]}) < $signed({1'h0, sel_295758}) ? {add_295755, array_index_295620[0]} : sel_295758;
  assign add_295862 = array_index_295725[11:1] + 11'h247;
  assign sel_295865 = $signed({1'h0, add_295760, array_index_295623[0]}) < $signed({1'h0, sel_295763}) ? {add_295760, array_index_295623[0]} : sel_295763;
  assign add_295890 = array_index_295824[11:0] + 12'h247;
  assign sel_295892 = $signed({1'h0, add_295788}) < $signed({1'h0, sel_295790}) ? add_295788 : sel_295790;
  assign add_295895 = array_index_295827[11:0] + 12'h247;
  assign sel_295897 = $signed({1'h0, add_295793}) < $signed({1'h0, sel_295795}) ? add_295793 : sel_295795;
  assign array_index_295926 = set1_unflattened[8'h84];
  assign array_index_295929 = set2_unflattened[8'h84];
  assign add_295933 = array_index_295518[11:1] + 11'h79d;
  assign sel_295935 = $signed({1'h0, add_295831, array_index_295416[0]}) < $signed({1'h0, sel_295833}) ? {add_295831, array_index_295416[0]} : sel_295833;
  assign add_295937 = array_index_295521[11:1] + 11'h79d;
  assign sel_295939 = $signed({1'h0, add_295835, array_index_295419[0]}) < $signed({1'h0, sel_295837}) ? {add_295835, array_index_295419[0]} : sel_295837;
  assign add_295941 = array_index_295620[11:1] + 11'h347;
  assign sel_295943 = $signed({1'h0, add_295839, array_index_295518[0]}) < $signed({1'h0, sel_295841}) ? {add_295839, array_index_295518[0]} : sel_295841;
  assign add_295945 = array_index_295623[11:1] + 11'h347;
  assign sel_295947 = $signed({1'h0, add_295843, array_index_295521[0]}) < $signed({1'h0, sel_295845}) ? {add_295843, array_index_295521[0]} : sel_295845;
  assign add_295949 = array_index_295722[11:3] + 9'h0bd;
  assign sel_295952 = $signed({1'h0, add_295847, array_index_295620[2:0]}) < $signed({1'h0, sel_295850}) ? {add_295847, array_index_295620[2:0]} : sel_295850;
  assign add_295954 = array_index_295725[11:3] + 9'h0bd;
  assign sel_295957 = $signed({1'h0, add_295852, array_index_295623[2:0]}) < $signed({1'h0, sel_295855}) ? {add_295852, array_index_295623[2:0]} : sel_295855;
  assign add_295959 = array_index_295824[11:1] + 11'h247;
  assign sel_295962 = $signed({1'h0, add_295857, array_index_295722[0]}) < $signed({1'h0, sel_295860}) ? {add_295857, array_index_295722[0]} : sel_295860;
  assign add_295964 = array_index_295827[11:1] + 11'h247;
  assign sel_295967 = $signed({1'h0, add_295862, array_index_295725[0]}) < $signed({1'h0, sel_295865}) ? {add_295862, array_index_295725[0]} : sel_295865;
  assign add_295992 = array_index_295926[11:0] + 12'h247;
  assign sel_295994 = $signed({1'h0, add_295890}) < $signed({1'h0, sel_295892}) ? add_295890 : sel_295892;
  assign add_295997 = array_index_295929[11:0] + 12'h247;
  assign sel_295999 = $signed({1'h0, add_295895}) < $signed({1'h0, sel_295897}) ? add_295895 : sel_295897;
  assign array_index_296028 = set1_unflattened[8'h85];
  assign array_index_296031 = set2_unflattened[8'h85];
  assign add_296035 = array_index_295620[11:1] + 11'h79d;
  assign sel_296037 = $signed({1'h0, add_295933, array_index_295518[0]}) < $signed({1'h0, sel_295935}) ? {add_295933, array_index_295518[0]} : sel_295935;
  assign add_296039 = array_index_295623[11:1] + 11'h79d;
  assign sel_296041 = $signed({1'h0, add_295937, array_index_295521[0]}) < $signed({1'h0, sel_295939}) ? {add_295937, array_index_295521[0]} : sel_295939;
  assign add_296043 = array_index_295722[11:1] + 11'h347;
  assign sel_296045 = $signed({1'h0, add_295941, array_index_295620[0]}) < $signed({1'h0, sel_295943}) ? {add_295941, array_index_295620[0]} : sel_295943;
  assign add_296047 = array_index_295725[11:1] + 11'h347;
  assign sel_296049 = $signed({1'h0, add_295945, array_index_295623[0]}) < $signed({1'h0, sel_295947}) ? {add_295945, array_index_295623[0]} : sel_295947;
  assign add_296051 = array_index_295824[11:3] + 9'h0bd;
  assign sel_296054 = $signed({1'h0, add_295949, array_index_295722[2:0]}) < $signed({1'h0, sel_295952}) ? {add_295949, array_index_295722[2:0]} : sel_295952;
  assign add_296056 = array_index_295827[11:3] + 9'h0bd;
  assign sel_296059 = $signed({1'h0, add_295954, array_index_295725[2:0]}) < $signed({1'h0, sel_295957}) ? {add_295954, array_index_295725[2:0]} : sel_295957;
  assign add_296061 = array_index_295926[11:1] + 11'h247;
  assign sel_296064 = $signed({1'h0, add_295959, array_index_295824[0]}) < $signed({1'h0, sel_295962}) ? {add_295959, array_index_295824[0]} : sel_295962;
  assign add_296066 = array_index_295929[11:1] + 11'h247;
  assign sel_296069 = $signed({1'h0, add_295964, array_index_295827[0]}) < $signed({1'h0, sel_295967}) ? {add_295964, array_index_295827[0]} : sel_295967;
  assign add_296094 = array_index_296028[11:0] + 12'h247;
  assign sel_296096 = $signed({1'h0, add_295992}) < $signed({1'h0, sel_295994}) ? add_295992 : sel_295994;
  assign add_296099 = array_index_296031[11:0] + 12'h247;
  assign sel_296101 = $signed({1'h0, add_295997}) < $signed({1'h0, sel_295999}) ? add_295997 : sel_295999;
  assign array_index_296130 = set1_unflattened[8'h86];
  assign array_index_296133 = set2_unflattened[8'h86];
  assign add_296137 = array_index_295722[11:1] + 11'h79d;
  assign sel_296139 = $signed({1'h0, add_296035, array_index_295620[0]}) < $signed({1'h0, sel_296037}) ? {add_296035, array_index_295620[0]} : sel_296037;
  assign add_296141 = array_index_295725[11:1] + 11'h79d;
  assign sel_296143 = $signed({1'h0, add_296039, array_index_295623[0]}) < $signed({1'h0, sel_296041}) ? {add_296039, array_index_295623[0]} : sel_296041;
  assign add_296145 = array_index_295824[11:1] + 11'h347;
  assign sel_296147 = $signed({1'h0, add_296043, array_index_295722[0]}) < $signed({1'h0, sel_296045}) ? {add_296043, array_index_295722[0]} : sel_296045;
  assign add_296149 = array_index_295827[11:1] + 11'h347;
  assign sel_296151 = $signed({1'h0, add_296047, array_index_295725[0]}) < $signed({1'h0, sel_296049}) ? {add_296047, array_index_295725[0]} : sel_296049;
  assign add_296153 = array_index_295926[11:3] + 9'h0bd;
  assign sel_296156 = $signed({1'h0, add_296051, array_index_295824[2:0]}) < $signed({1'h0, sel_296054}) ? {add_296051, array_index_295824[2:0]} : sel_296054;
  assign add_296158 = array_index_295929[11:3] + 9'h0bd;
  assign sel_296161 = $signed({1'h0, add_296056, array_index_295827[2:0]}) < $signed({1'h0, sel_296059}) ? {add_296056, array_index_295827[2:0]} : sel_296059;
  assign add_296163 = array_index_296028[11:1] + 11'h247;
  assign sel_296166 = $signed({1'h0, add_296061, array_index_295926[0]}) < $signed({1'h0, sel_296064}) ? {add_296061, array_index_295926[0]} : sel_296064;
  assign add_296168 = array_index_296031[11:1] + 11'h247;
  assign sel_296171 = $signed({1'h0, add_296066, array_index_295929[0]}) < $signed({1'h0, sel_296069}) ? {add_296066, array_index_295929[0]} : sel_296069;
  assign add_296196 = array_index_296130[11:0] + 12'h247;
  assign sel_296198 = $signed({1'h0, add_296094}) < $signed({1'h0, sel_296096}) ? add_296094 : sel_296096;
  assign add_296201 = array_index_296133[11:0] + 12'h247;
  assign sel_296203 = $signed({1'h0, add_296099}) < $signed({1'h0, sel_296101}) ? add_296099 : sel_296101;
  assign array_index_296232 = set1_unflattened[8'h87];
  assign array_index_296235 = set2_unflattened[8'h87];
  assign add_296239 = array_index_295824[11:1] + 11'h79d;
  assign sel_296241 = $signed({1'h0, add_296137, array_index_295722[0]}) < $signed({1'h0, sel_296139}) ? {add_296137, array_index_295722[0]} : sel_296139;
  assign add_296243 = array_index_295827[11:1] + 11'h79d;
  assign sel_296245 = $signed({1'h0, add_296141, array_index_295725[0]}) < $signed({1'h0, sel_296143}) ? {add_296141, array_index_295725[0]} : sel_296143;
  assign add_296247 = array_index_295926[11:1] + 11'h347;
  assign sel_296249 = $signed({1'h0, add_296145, array_index_295824[0]}) < $signed({1'h0, sel_296147}) ? {add_296145, array_index_295824[0]} : sel_296147;
  assign add_296251 = array_index_295929[11:1] + 11'h347;
  assign sel_296253 = $signed({1'h0, add_296149, array_index_295827[0]}) < $signed({1'h0, sel_296151}) ? {add_296149, array_index_295827[0]} : sel_296151;
  assign add_296255 = array_index_296028[11:3] + 9'h0bd;
  assign sel_296258 = $signed({1'h0, add_296153, array_index_295926[2:0]}) < $signed({1'h0, sel_296156}) ? {add_296153, array_index_295926[2:0]} : sel_296156;
  assign add_296260 = array_index_296031[11:3] + 9'h0bd;
  assign sel_296263 = $signed({1'h0, add_296158, array_index_295929[2:0]}) < $signed({1'h0, sel_296161}) ? {add_296158, array_index_295929[2:0]} : sel_296161;
  assign add_296265 = array_index_296130[11:1] + 11'h247;
  assign sel_296268 = $signed({1'h0, add_296163, array_index_296028[0]}) < $signed({1'h0, sel_296166}) ? {add_296163, array_index_296028[0]} : sel_296166;
  assign add_296270 = array_index_296133[11:1] + 11'h247;
  assign sel_296273 = $signed({1'h0, add_296168, array_index_296031[0]}) < $signed({1'h0, sel_296171}) ? {add_296168, array_index_296031[0]} : sel_296171;
  assign add_296298 = array_index_296232[11:0] + 12'h247;
  assign sel_296300 = $signed({1'h0, add_296196}) < $signed({1'h0, sel_296198}) ? add_296196 : sel_296198;
  assign add_296303 = array_index_296235[11:0] + 12'h247;
  assign sel_296305 = $signed({1'h0, add_296201}) < $signed({1'h0, sel_296203}) ? add_296201 : sel_296203;
  assign array_index_296334 = set1_unflattened[8'h88];
  assign array_index_296337 = set2_unflattened[8'h88];
  assign add_296341 = array_index_295926[11:1] + 11'h79d;
  assign sel_296343 = $signed({1'h0, add_296239, array_index_295824[0]}) < $signed({1'h0, sel_296241}) ? {add_296239, array_index_295824[0]} : sel_296241;
  assign add_296345 = array_index_295929[11:1] + 11'h79d;
  assign sel_296347 = $signed({1'h0, add_296243, array_index_295827[0]}) < $signed({1'h0, sel_296245}) ? {add_296243, array_index_295827[0]} : sel_296245;
  assign add_296349 = array_index_296028[11:1] + 11'h347;
  assign sel_296351 = $signed({1'h0, add_296247, array_index_295926[0]}) < $signed({1'h0, sel_296249}) ? {add_296247, array_index_295926[0]} : sel_296249;
  assign add_296353 = array_index_296031[11:1] + 11'h347;
  assign sel_296355 = $signed({1'h0, add_296251, array_index_295929[0]}) < $signed({1'h0, sel_296253}) ? {add_296251, array_index_295929[0]} : sel_296253;
  assign add_296357 = array_index_296130[11:3] + 9'h0bd;
  assign sel_296360 = $signed({1'h0, add_296255, array_index_296028[2:0]}) < $signed({1'h0, sel_296258}) ? {add_296255, array_index_296028[2:0]} : sel_296258;
  assign add_296362 = array_index_296133[11:3] + 9'h0bd;
  assign sel_296365 = $signed({1'h0, add_296260, array_index_296031[2:0]}) < $signed({1'h0, sel_296263}) ? {add_296260, array_index_296031[2:0]} : sel_296263;
  assign add_296367 = array_index_296232[11:1] + 11'h247;
  assign sel_296370 = $signed({1'h0, add_296265, array_index_296130[0]}) < $signed({1'h0, sel_296268}) ? {add_296265, array_index_296130[0]} : sel_296268;
  assign add_296372 = array_index_296235[11:1] + 11'h247;
  assign sel_296375 = $signed({1'h0, add_296270, array_index_296133[0]}) < $signed({1'h0, sel_296273}) ? {add_296270, array_index_296133[0]} : sel_296273;
  assign add_296400 = array_index_296334[11:0] + 12'h247;
  assign sel_296402 = $signed({1'h0, add_296298}) < $signed({1'h0, sel_296300}) ? add_296298 : sel_296300;
  assign add_296405 = array_index_296337[11:0] + 12'h247;
  assign sel_296407 = $signed({1'h0, add_296303}) < $signed({1'h0, sel_296305}) ? add_296303 : sel_296305;
  assign array_index_296436 = set1_unflattened[8'h89];
  assign array_index_296439 = set2_unflattened[8'h89];
  assign add_296443 = array_index_296028[11:1] + 11'h79d;
  assign sel_296445 = $signed({1'h0, add_296341, array_index_295926[0]}) < $signed({1'h0, sel_296343}) ? {add_296341, array_index_295926[0]} : sel_296343;
  assign add_296447 = array_index_296031[11:1] + 11'h79d;
  assign sel_296449 = $signed({1'h0, add_296345, array_index_295929[0]}) < $signed({1'h0, sel_296347}) ? {add_296345, array_index_295929[0]} : sel_296347;
  assign add_296451 = array_index_296130[11:1] + 11'h347;
  assign sel_296453 = $signed({1'h0, add_296349, array_index_296028[0]}) < $signed({1'h0, sel_296351}) ? {add_296349, array_index_296028[0]} : sel_296351;
  assign add_296455 = array_index_296133[11:1] + 11'h347;
  assign sel_296457 = $signed({1'h0, add_296353, array_index_296031[0]}) < $signed({1'h0, sel_296355}) ? {add_296353, array_index_296031[0]} : sel_296355;
  assign add_296459 = array_index_296232[11:3] + 9'h0bd;
  assign sel_296462 = $signed({1'h0, add_296357, array_index_296130[2:0]}) < $signed({1'h0, sel_296360}) ? {add_296357, array_index_296130[2:0]} : sel_296360;
  assign add_296464 = array_index_296235[11:3] + 9'h0bd;
  assign sel_296467 = $signed({1'h0, add_296362, array_index_296133[2:0]}) < $signed({1'h0, sel_296365}) ? {add_296362, array_index_296133[2:0]} : sel_296365;
  assign add_296469 = array_index_296334[11:1] + 11'h247;
  assign sel_296472 = $signed({1'h0, add_296367, array_index_296232[0]}) < $signed({1'h0, sel_296370}) ? {add_296367, array_index_296232[0]} : sel_296370;
  assign add_296474 = array_index_296337[11:1] + 11'h247;
  assign sel_296477 = $signed({1'h0, add_296372, array_index_296235[0]}) < $signed({1'h0, sel_296375}) ? {add_296372, array_index_296235[0]} : sel_296375;
  assign add_296502 = array_index_296436[11:0] + 12'h247;
  assign sel_296504 = $signed({1'h0, add_296400}) < $signed({1'h0, sel_296402}) ? add_296400 : sel_296402;
  assign add_296507 = array_index_296439[11:0] + 12'h247;
  assign sel_296509 = $signed({1'h0, add_296405}) < $signed({1'h0, sel_296407}) ? add_296405 : sel_296407;
  assign array_index_296538 = set1_unflattened[8'h8a];
  assign array_index_296541 = set2_unflattened[8'h8a];
  assign add_296545 = array_index_296130[11:1] + 11'h79d;
  assign sel_296547 = $signed({1'h0, add_296443, array_index_296028[0]}) < $signed({1'h0, sel_296445}) ? {add_296443, array_index_296028[0]} : sel_296445;
  assign add_296549 = array_index_296133[11:1] + 11'h79d;
  assign sel_296551 = $signed({1'h0, add_296447, array_index_296031[0]}) < $signed({1'h0, sel_296449}) ? {add_296447, array_index_296031[0]} : sel_296449;
  assign add_296553 = array_index_296232[11:1] + 11'h347;
  assign sel_296555 = $signed({1'h0, add_296451, array_index_296130[0]}) < $signed({1'h0, sel_296453}) ? {add_296451, array_index_296130[0]} : sel_296453;
  assign add_296557 = array_index_296235[11:1] + 11'h347;
  assign sel_296559 = $signed({1'h0, add_296455, array_index_296133[0]}) < $signed({1'h0, sel_296457}) ? {add_296455, array_index_296133[0]} : sel_296457;
  assign add_296561 = array_index_296334[11:3] + 9'h0bd;
  assign sel_296564 = $signed({1'h0, add_296459, array_index_296232[2:0]}) < $signed({1'h0, sel_296462}) ? {add_296459, array_index_296232[2:0]} : sel_296462;
  assign add_296566 = array_index_296337[11:3] + 9'h0bd;
  assign sel_296569 = $signed({1'h0, add_296464, array_index_296235[2:0]}) < $signed({1'h0, sel_296467}) ? {add_296464, array_index_296235[2:0]} : sel_296467;
  assign add_296571 = array_index_296436[11:1] + 11'h247;
  assign sel_296574 = $signed({1'h0, add_296469, array_index_296334[0]}) < $signed({1'h0, sel_296472}) ? {add_296469, array_index_296334[0]} : sel_296472;
  assign add_296576 = array_index_296439[11:1] + 11'h247;
  assign sel_296579 = $signed({1'h0, add_296474, array_index_296337[0]}) < $signed({1'h0, sel_296477}) ? {add_296474, array_index_296337[0]} : sel_296477;
  assign add_296604 = array_index_296538[11:0] + 12'h247;
  assign sel_296606 = $signed({1'h0, add_296502}) < $signed({1'h0, sel_296504}) ? add_296502 : sel_296504;
  assign add_296609 = array_index_296541[11:0] + 12'h247;
  assign sel_296611 = $signed({1'h0, add_296507}) < $signed({1'h0, sel_296509}) ? add_296507 : sel_296509;
  assign array_index_296640 = set1_unflattened[8'h8b];
  assign array_index_296643 = set2_unflattened[8'h8b];
  assign add_296647 = array_index_296232[11:1] + 11'h79d;
  assign sel_296649 = $signed({1'h0, add_296545, array_index_296130[0]}) < $signed({1'h0, sel_296547}) ? {add_296545, array_index_296130[0]} : sel_296547;
  assign add_296651 = array_index_296235[11:1] + 11'h79d;
  assign sel_296653 = $signed({1'h0, add_296549, array_index_296133[0]}) < $signed({1'h0, sel_296551}) ? {add_296549, array_index_296133[0]} : sel_296551;
  assign add_296655 = array_index_296334[11:1] + 11'h347;
  assign sel_296657 = $signed({1'h0, add_296553, array_index_296232[0]}) < $signed({1'h0, sel_296555}) ? {add_296553, array_index_296232[0]} : sel_296555;
  assign add_296659 = array_index_296337[11:1] + 11'h347;
  assign sel_296661 = $signed({1'h0, add_296557, array_index_296235[0]}) < $signed({1'h0, sel_296559}) ? {add_296557, array_index_296235[0]} : sel_296559;
  assign add_296663 = array_index_296436[11:3] + 9'h0bd;
  assign sel_296666 = $signed({1'h0, add_296561, array_index_296334[2:0]}) < $signed({1'h0, sel_296564}) ? {add_296561, array_index_296334[2:0]} : sel_296564;
  assign add_296668 = array_index_296439[11:3] + 9'h0bd;
  assign sel_296671 = $signed({1'h0, add_296566, array_index_296337[2:0]}) < $signed({1'h0, sel_296569}) ? {add_296566, array_index_296337[2:0]} : sel_296569;
  assign add_296673 = array_index_296538[11:1] + 11'h247;
  assign sel_296676 = $signed({1'h0, add_296571, array_index_296436[0]}) < $signed({1'h0, sel_296574}) ? {add_296571, array_index_296436[0]} : sel_296574;
  assign add_296678 = array_index_296541[11:1] + 11'h247;
  assign sel_296681 = $signed({1'h0, add_296576, array_index_296439[0]}) < $signed({1'h0, sel_296579}) ? {add_296576, array_index_296439[0]} : sel_296579;
  assign add_296706 = array_index_296640[11:0] + 12'h247;
  assign sel_296708 = $signed({1'h0, add_296604}) < $signed({1'h0, sel_296606}) ? add_296604 : sel_296606;
  assign add_296711 = array_index_296643[11:0] + 12'h247;
  assign sel_296713 = $signed({1'h0, add_296609}) < $signed({1'h0, sel_296611}) ? add_296609 : sel_296611;
  assign array_index_296742 = set1_unflattened[8'h8c];
  assign array_index_296745 = set2_unflattened[8'h8c];
  assign add_296749 = array_index_296334[11:1] + 11'h79d;
  assign sel_296751 = $signed({1'h0, add_296647, array_index_296232[0]}) < $signed({1'h0, sel_296649}) ? {add_296647, array_index_296232[0]} : sel_296649;
  assign add_296753 = array_index_296337[11:1] + 11'h79d;
  assign sel_296755 = $signed({1'h0, add_296651, array_index_296235[0]}) < $signed({1'h0, sel_296653}) ? {add_296651, array_index_296235[0]} : sel_296653;
  assign add_296757 = array_index_296436[11:1] + 11'h347;
  assign sel_296759 = $signed({1'h0, add_296655, array_index_296334[0]}) < $signed({1'h0, sel_296657}) ? {add_296655, array_index_296334[0]} : sel_296657;
  assign add_296761 = array_index_296439[11:1] + 11'h347;
  assign sel_296763 = $signed({1'h0, add_296659, array_index_296337[0]}) < $signed({1'h0, sel_296661}) ? {add_296659, array_index_296337[0]} : sel_296661;
  assign add_296765 = array_index_296538[11:3] + 9'h0bd;
  assign sel_296768 = $signed({1'h0, add_296663, array_index_296436[2:0]}) < $signed({1'h0, sel_296666}) ? {add_296663, array_index_296436[2:0]} : sel_296666;
  assign add_296770 = array_index_296541[11:3] + 9'h0bd;
  assign sel_296773 = $signed({1'h0, add_296668, array_index_296439[2:0]}) < $signed({1'h0, sel_296671}) ? {add_296668, array_index_296439[2:0]} : sel_296671;
  assign add_296775 = array_index_296640[11:1] + 11'h247;
  assign sel_296778 = $signed({1'h0, add_296673, array_index_296538[0]}) < $signed({1'h0, sel_296676}) ? {add_296673, array_index_296538[0]} : sel_296676;
  assign add_296780 = array_index_296643[11:1] + 11'h247;
  assign sel_296783 = $signed({1'h0, add_296678, array_index_296541[0]}) < $signed({1'h0, sel_296681}) ? {add_296678, array_index_296541[0]} : sel_296681;
  assign add_296808 = array_index_296742[11:0] + 12'h247;
  assign sel_296810 = $signed({1'h0, add_296706}) < $signed({1'h0, sel_296708}) ? add_296706 : sel_296708;
  assign add_296813 = array_index_296745[11:0] + 12'h247;
  assign sel_296815 = $signed({1'h0, add_296711}) < $signed({1'h0, sel_296713}) ? add_296711 : sel_296713;
  assign array_index_296844 = set1_unflattened[8'h8d];
  assign array_index_296847 = set2_unflattened[8'h8d];
  assign add_296851 = array_index_296436[11:1] + 11'h79d;
  assign sel_296853 = $signed({1'h0, add_296749, array_index_296334[0]}) < $signed({1'h0, sel_296751}) ? {add_296749, array_index_296334[0]} : sel_296751;
  assign add_296855 = array_index_296439[11:1] + 11'h79d;
  assign sel_296857 = $signed({1'h0, add_296753, array_index_296337[0]}) < $signed({1'h0, sel_296755}) ? {add_296753, array_index_296337[0]} : sel_296755;
  assign add_296859 = array_index_296538[11:1] + 11'h347;
  assign sel_296861 = $signed({1'h0, add_296757, array_index_296436[0]}) < $signed({1'h0, sel_296759}) ? {add_296757, array_index_296436[0]} : sel_296759;
  assign add_296863 = array_index_296541[11:1] + 11'h347;
  assign sel_296865 = $signed({1'h0, add_296761, array_index_296439[0]}) < $signed({1'h0, sel_296763}) ? {add_296761, array_index_296439[0]} : sel_296763;
  assign add_296867 = array_index_296640[11:3] + 9'h0bd;
  assign sel_296870 = $signed({1'h0, add_296765, array_index_296538[2:0]}) < $signed({1'h0, sel_296768}) ? {add_296765, array_index_296538[2:0]} : sel_296768;
  assign add_296872 = array_index_296643[11:3] + 9'h0bd;
  assign sel_296875 = $signed({1'h0, add_296770, array_index_296541[2:0]}) < $signed({1'h0, sel_296773}) ? {add_296770, array_index_296541[2:0]} : sel_296773;
  assign add_296877 = array_index_296742[11:1] + 11'h247;
  assign sel_296880 = $signed({1'h0, add_296775, array_index_296640[0]}) < $signed({1'h0, sel_296778}) ? {add_296775, array_index_296640[0]} : sel_296778;
  assign add_296882 = array_index_296745[11:1] + 11'h247;
  assign sel_296885 = $signed({1'h0, add_296780, array_index_296643[0]}) < $signed({1'h0, sel_296783}) ? {add_296780, array_index_296643[0]} : sel_296783;
  assign add_296910 = array_index_296844[11:0] + 12'h247;
  assign sel_296912 = $signed({1'h0, add_296808}) < $signed({1'h0, sel_296810}) ? add_296808 : sel_296810;
  assign add_296915 = array_index_296847[11:0] + 12'h247;
  assign sel_296917 = $signed({1'h0, add_296813}) < $signed({1'h0, sel_296815}) ? add_296813 : sel_296815;
  assign array_index_296946 = set1_unflattened[8'h8e];
  assign array_index_296949 = set2_unflattened[8'h8e];
  assign add_296953 = array_index_296538[11:1] + 11'h79d;
  assign sel_296955 = $signed({1'h0, add_296851, array_index_296436[0]}) < $signed({1'h0, sel_296853}) ? {add_296851, array_index_296436[0]} : sel_296853;
  assign add_296957 = array_index_296541[11:1] + 11'h79d;
  assign sel_296959 = $signed({1'h0, add_296855, array_index_296439[0]}) < $signed({1'h0, sel_296857}) ? {add_296855, array_index_296439[0]} : sel_296857;
  assign add_296961 = array_index_296640[11:1] + 11'h347;
  assign sel_296963 = $signed({1'h0, add_296859, array_index_296538[0]}) < $signed({1'h0, sel_296861}) ? {add_296859, array_index_296538[0]} : sel_296861;
  assign add_296965 = array_index_296643[11:1] + 11'h347;
  assign sel_296967 = $signed({1'h0, add_296863, array_index_296541[0]}) < $signed({1'h0, sel_296865}) ? {add_296863, array_index_296541[0]} : sel_296865;
  assign add_296969 = array_index_296742[11:3] + 9'h0bd;
  assign sel_296972 = $signed({1'h0, add_296867, array_index_296640[2:0]}) < $signed({1'h0, sel_296870}) ? {add_296867, array_index_296640[2:0]} : sel_296870;
  assign add_296974 = array_index_296745[11:3] + 9'h0bd;
  assign sel_296977 = $signed({1'h0, add_296872, array_index_296643[2:0]}) < $signed({1'h0, sel_296875}) ? {add_296872, array_index_296643[2:0]} : sel_296875;
  assign add_296979 = array_index_296844[11:1] + 11'h247;
  assign sel_296982 = $signed({1'h0, add_296877, array_index_296742[0]}) < $signed({1'h0, sel_296880}) ? {add_296877, array_index_296742[0]} : sel_296880;
  assign add_296984 = array_index_296847[11:1] + 11'h247;
  assign sel_296987 = $signed({1'h0, add_296882, array_index_296745[0]}) < $signed({1'h0, sel_296885}) ? {add_296882, array_index_296745[0]} : sel_296885;
  assign add_297012 = array_index_296946[11:0] + 12'h247;
  assign sel_297014 = $signed({1'h0, add_296910}) < $signed({1'h0, sel_296912}) ? add_296910 : sel_296912;
  assign add_297017 = array_index_296949[11:0] + 12'h247;
  assign sel_297019 = $signed({1'h0, add_296915}) < $signed({1'h0, sel_296917}) ? add_296915 : sel_296917;
  assign array_index_297048 = set1_unflattened[8'h8f];
  assign array_index_297051 = set2_unflattened[8'h8f];
  assign add_297055 = array_index_296640[11:1] + 11'h79d;
  assign sel_297057 = $signed({1'h0, add_296953, array_index_296538[0]}) < $signed({1'h0, sel_296955}) ? {add_296953, array_index_296538[0]} : sel_296955;
  assign add_297059 = array_index_296643[11:1] + 11'h79d;
  assign sel_297061 = $signed({1'h0, add_296957, array_index_296541[0]}) < $signed({1'h0, sel_296959}) ? {add_296957, array_index_296541[0]} : sel_296959;
  assign add_297063 = array_index_296742[11:1] + 11'h347;
  assign sel_297065 = $signed({1'h0, add_296961, array_index_296640[0]}) < $signed({1'h0, sel_296963}) ? {add_296961, array_index_296640[0]} : sel_296963;
  assign add_297067 = array_index_296745[11:1] + 11'h347;
  assign sel_297069 = $signed({1'h0, add_296965, array_index_296643[0]}) < $signed({1'h0, sel_296967}) ? {add_296965, array_index_296643[0]} : sel_296967;
  assign add_297071 = array_index_296844[11:3] + 9'h0bd;
  assign sel_297074 = $signed({1'h0, add_296969, array_index_296742[2:0]}) < $signed({1'h0, sel_296972}) ? {add_296969, array_index_296742[2:0]} : sel_296972;
  assign add_297076 = array_index_296847[11:3] + 9'h0bd;
  assign sel_297079 = $signed({1'h0, add_296974, array_index_296745[2:0]}) < $signed({1'h0, sel_296977}) ? {add_296974, array_index_296745[2:0]} : sel_296977;
  assign add_297081 = array_index_296946[11:1] + 11'h247;
  assign sel_297084 = $signed({1'h0, add_296979, array_index_296844[0]}) < $signed({1'h0, sel_296982}) ? {add_296979, array_index_296844[0]} : sel_296982;
  assign add_297086 = array_index_296949[11:1] + 11'h247;
  assign sel_297089 = $signed({1'h0, add_296984, array_index_296847[0]}) < $signed({1'h0, sel_296987}) ? {add_296984, array_index_296847[0]} : sel_296987;
  assign add_297114 = array_index_297048[11:0] + 12'h247;
  assign sel_297116 = $signed({1'h0, add_297012}) < $signed({1'h0, sel_297014}) ? add_297012 : sel_297014;
  assign add_297119 = array_index_297051[11:0] + 12'h247;
  assign sel_297121 = $signed({1'h0, add_297017}) < $signed({1'h0, sel_297019}) ? add_297017 : sel_297019;
  assign array_index_297150 = set1_unflattened[8'h90];
  assign array_index_297153 = set2_unflattened[8'h90];
  assign add_297157 = array_index_296742[11:1] + 11'h79d;
  assign sel_297159 = $signed({1'h0, add_297055, array_index_296640[0]}) < $signed({1'h0, sel_297057}) ? {add_297055, array_index_296640[0]} : sel_297057;
  assign add_297161 = array_index_296745[11:1] + 11'h79d;
  assign sel_297163 = $signed({1'h0, add_297059, array_index_296643[0]}) < $signed({1'h0, sel_297061}) ? {add_297059, array_index_296643[0]} : sel_297061;
  assign add_297165 = array_index_296844[11:1] + 11'h347;
  assign sel_297167 = $signed({1'h0, add_297063, array_index_296742[0]}) < $signed({1'h0, sel_297065}) ? {add_297063, array_index_296742[0]} : sel_297065;
  assign add_297169 = array_index_296847[11:1] + 11'h347;
  assign sel_297171 = $signed({1'h0, add_297067, array_index_296745[0]}) < $signed({1'h0, sel_297069}) ? {add_297067, array_index_296745[0]} : sel_297069;
  assign add_297173 = array_index_296946[11:3] + 9'h0bd;
  assign sel_297176 = $signed({1'h0, add_297071, array_index_296844[2:0]}) < $signed({1'h0, sel_297074}) ? {add_297071, array_index_296844[2:0]} : sel_297074;
  assign add_297178 = array_index_296949[11:3] + 9'h0bd;
  assign sel_297181 = $signed({1'h0, add_297076, array_index_296847[2:0]}) < $signed({1'h0, sel_297079}) ? {add_297076, array_index_296847[2:0]} : sel_297079;
  assign add_297183 = array_index_297048[11:1] + 11'h247;
  assign sel_297186 = $signed({1'h0, add_297081, array_index_296946[0]}) < $signed({1'h0, sel_297084}) ? {add_297081, array_index_296946[0]} : sel_297084;
  assign add_297188 = array_index_297051[11:1] + 11'h247;
  assign sel_297191 = $signed({1'h0, add_297086, array_index_296949[0]}) < $signed({1'h0, sel_297089}) ? {add_297086, array_index_296949[0]} : sel_297089;
  assign add_297216 = array_index_297150[11:0] + 12'h247;
  assign sel_297218 = $signed({1'h0, add_297114}) < $signed({1'h0, sel_297116}) ? add_297114 : sel_297116;
  assign add_297221 = array_index_297153[11:0] + 12'h247;
  assign sel_297223 = $signed({1'h0, add_297119}) < $signed({1'h0, sel_297121}) ? add_297119 : sel_297121;
  assign array_index_297252 = set1_unflattened[8'h91];
  assign array_index_297255 = set2_unflattened[8'h91];
  assign add_297259 = array_index_296844[11:1] + 11'h79d;
  assign sel_297261 = $signed({1'h0, add_297157, array_index_296742[0]}) < $signed({1'h0, sel_297159}) ? {add_297157, array_index_296742[0]} : sel_297159;
  assign add_297263 = array_index_296847[11:1] + 11'h79d;
  assign sel_297265 = $signed({1'h0, add_297161, array_index_296745[0]}) < $signed({1'h0, sel_297163}) ? {add_297161, array_index_296745[0]} : sel_297163;
  assign add_297267 = array_index_296946[11:1] + 11'h347;
  assign sel_297269 = $signed({1'h0, add_297165, array_index_296844[0]}) < $signed({1'h0, sel_297167}) ? {add_297165, array_index_296844[0]} : sel_297167;
  assign add_297271 = array_index_296949[11:1] + 11'h347;
  assign sel_297273 = $signed({1'h0, add_297169, array_index_296847[0]}) < $signed({1'h0, sel_297171}) ? {add_297169, array_index_296847[0]} : sel_297171;
  assign add_297275 = array_index_297048[11:3] + 9'h0bd;
  assign sel_297278 = $signed({1'h0, add_297173, array_index_296946[2:0]}) < $signed({1'h0, sel_297176}) ? {add_297173, array_index_296946[2:0]} : sel_297176;
  assign add_297280 = array_index_297051[11:3] + 9'h0bd;
  assign sel_297283 = $signed({1'h0, add_297178, array_index_296949[2:0]}) < $signed({1'h0, sel_297181}) ? {add_297178, array_index_296949[2:0]} : sel_297181;
  assign add_297285 = array_index_297150[11:1] + 11'h247;
  assign sel_297288 = $signed({1'h0, add_297183, array_index_297048[0]}) < $signed({1'h0, sel_297186}) ? {add_297183, array_index_297048[0]} : sel_297186;
  assign add_297290 = array_index_297153[11:1] + 11'h247;
  assign sel_297293 = $signed({1'h0, add_297188, array_index_297051[0]}) < $signed({1'h0, sel_297191}) ? {add_297188, array_index_297051[0]} : sel_297191;
  assign add_297318 = array_index_297252[11:0] + 12'h247;
  assign sel_297320 = $signed({1'h0, add_297216}) < $signed({1'h0, sel_297218}) ? add_297216 : sel_297218;
  assign add_297323 = array_index_297255[11:0] + 12'h247;
  assign sel_297325 = $signed({1'h0, add_297221}) < $signed({1'h0, sel_297223}) ? add_297221 : sel_297223;
  assign array_index_297354 = set1_unflattened[8'h92];
  assign array_index_297357 = set2_unflattened[8'h92];
  assign add_297361 = array_index_296946[11:1] + 11'h79d;
  assign sel_297363 = $signed({1'h0, add_297259, array_index_296844[0]}) < $signed({1'h0, sel_297261}) ? {add_297259, array_index_296844[0]} : sel_297261;
  assign add_297365 = array_index_296949[11:1] + 11'h79d;
  assign sel_297367 = $signed({1'h0, add_297263, array_index_296847[0]}) < $signed({1'h0, sel_297265}) ? {add_297263, array_index_296847[0]} : sel_297265;
  assign add_297369 = array_index_297048[11:1] + 11'h347;
  assign sel_297371 = $signed({1'h0, add_297267, array_index_296946[0]}) < $signed({1'h0, sel_297269}) ? {add_297267, array_index_296946[0]} : sel_297269;
  assign add_297373 = array_index_297051[11:1] + 11'h347;
  assign sel_297375 = $signed({1'h0, add_297271, array_index_296949[0]}) < $signed({1'h0, sel_297273}) ? {add_297271, array_index_296949[0]} : sel_297273;
  assign add_297377 = array_index_297150[11:3] + 9'h0bd;
  assign sel_297380 = $signed({1'h0, add_297275, array_index_297048[2:0]}) < $signed({1'h0, sel_297278}) ? {add_297275, array_index_297048[2:0]} : sel_297278;
  assign add_297382 = array_index_297153[11:3] + 9'h0bd;
  assign sel_297385 = $signed({1'h0, add_297280, array_index_297051[2:0]}) < $signed({1'h0, sel_297283}) ? {add_297280, array_index_297051[2:0]} : sel_297283;
  assign add_297387 = array_index_297252[11:1] + 11'h247;
  assign sel_297390 = $signed({1'h0, add_297285, array_index_297150[0]}) < $signed({1'h0, sel_297288}) ? {add_297285, array_index_297150[0]} : sel_297288;
  assign add_297392 = array_index_297255[11:1] + 11'h247;
  assign sel_297395 = $signed({1'h0, add_297290, array_index_297153[0]}) < $signed({1'h0, sel_297293}) ? {add_297290, array_index_297153[0]} : sel_297293;
  assign add_297420 = array_index_297354[11:0] + 12'h247;
  assign sel_297422 = $signed({1'h0, add_297318}) < $signed({1'h0, sel_297320}) ? add_297318 : sel_297320;
  assign add_297425 = array_index_297357[11:0] + 12'h247;
  assign sel_297427 = $signed({1'h0, add_297323}) < $signed({1'h0, sel_297325}) ? add_297323 : sel_297325;
  assign array_index_297456 = set1_unflattened[8'h93];
  assign array_index_297459 = set2_unflattened[8'h93];
  assign add_297463 = array_index_297048[11:1] + 11'h79d;
  assign sel_297465 = $signed({1'h0, add_297361, array_index_296946[0]}) < $signed({1'h0, sel_297363}) ? {add_297361, array_index_296946[0]} : sel_297363;
  assign add_297467 = array_index_297051[11:1] + 11'h79d;
  assign sel_297469 = $signed({1'h0, add_297365, array_index_296949[0]}) < $signed({1'h0, sel_297367}) ? {add_297365, array_index_296949[0]} : sel_297367;
  assign add_297471 = array_index_297150[11:1] + 11'h347;
  assign sel_297473 = $signed({1'h0, add_297369, array_index_297048[0]}) < $signed({1'h0, sel_297371}) ? {add_297369, array_index_297048[0]} : sel_297371;
  assign add_297475 = array_index_297153[11:1] + 11'h347;
  assign sel_297477 = $signed({1'h0, add_297373, array_index_297051[0]}) < $signed({1'h0, sel_297375}) ? {add_297373, array_index_297051[0]} : sel_297375;
  assign add_297479 = array_index_297252[11:3] + 9'h0bd;
  assign sel_297482 = $signed({1'h0, add_297377, array_index_297150[2:0]}) < $signed({1'h0, sel_297380}) ? {add_297377, array_index_297150[2:0]} : sel_297380;
  assign add_297484 = array_index_297255[11:3] + 9'h0bd;
  assign sel_297487 = $signed({1'h0, add_297382, array_index_297153[2:0]}) < $signed({1'h0, sel_297385}) ? {add_297382, array_index_297153[2:0]} : sel_297385;
  assign add_297489 = array_index_297354[11:1] + 11'h247;
  assign sel_297492 = $signed({1'h0, add_297387, array_index_297252[0]}) < $signed({1'h0, sel_297390}) ? {add_297387, array_index_297252[0]} : sel_297390;
  assign add_297494 = array_index_297357[11:1] + 11'h247;
  assign sel_297497 = $signed({1'h0, add_297392, array_index_297255[0]}) < $signed({1'h0, sel_297395}) ? {add_297392, array_index_297255[0]} : sel_297395;
  assign add_297522 = array_index_297456[11:0] + 12'h247;
  assign sel_297524 = $signed({1'h0, add_297420}) < $signed({1'h0, sel_297422}) ? add_297420 : sel_297422;
  assign add_297527 = array_index_297459[11:0] + 12'h247;
  assign sel_297529 = $signed({1'h0, add_297425}) < $signed({1'h0, sel_297427}) ? add_297425 : sel_297427;
  assign array_index_297558 = set1_unflattened[8'h94];
  assign array_index_297561 = set2_unflattened[8'h94];
  assign add_297565 = array_index_297150[11:1] + 11'h79d;
  assign sel_297567 = $signed({1'h0, add_297463, array_index_297048[0]}) < $signed({1'h0, sel_297465}) ? {add_297463, array_index_297048[0]} : sel_297465;
  assign add_297569 = array_index_297153[11:1] + 11'h79d;
  assign sel_297571 = $signed({1'h0, add_297467, array_index_297051[0]}) < $signed({1'h0, sel_297469}) ? {add_297467, array_index_297051[0]} : sel_297469;
  assign add_297573 = array_index_297252[11:1] + 11'h347;
  assign sel_297575 = $signed({1'h0, add_297471, array_index_297150[0]}) < $signed({1'h0, sel_297473}) ? {add_297471, array_index_297150[0]} : sel_297473;
  assign add_297577 = array_index_297255[11:1] + 11'h347;
  assign sel_297579 = $signed({1'h0, add_297475, array_index_297153[0]}) < $signed({1'h0, sel_297477}) ? {add_297475, array_index_297153[0]} : sel_297477;
  assign add_297581 = array_index_297354[11:3] + 9'h0bd;
  assign sel_297584 = $signed({1'h0, add_297479, array_index_297252[2:0]}) < $signed({1'h0, sel_297482}) ? {add_297479, array_index_297252[2:0]} : sel_297482;
  assign add_297586 = array_index_297357[11:3] + 9'h0bd;
  assign sel_297589 = $signed({1'h0, add_297484, array_index_297255[2:0]}) < $signed({1'h0, sel_297487}) ? {add_297484, array_index_297255[2:0]} : sel_297487;
  assign add_297591 = array_index_297456[11:1] + 11'h247;
  assign sel_297594 = $signed({1'h0, add_297489, array_index_297354[0]}) < $signed({1'h0, sel_297492}) ? {add_297489, array_index_297354[0]} : sel_297492;
  assign add_297596 = array_index_297459[11:1] + 11'h247;
  assign sel_297599 = $signed({1'h0, add_297494, array_index_297357[0]}) < $signed({1'h0, sel_297497}) ? {add_297494, array_index_297357[0]} : sel_297497;
  assign add_297624 = array_index_297558[11:0] + 12'h247;
  assign sel_297626 = $signed({1'h0, add_297522}) < $signed({1'h0, sel_297524}) ? add_297522 : sel_297524;
  assign add_297629 = array_index_297561[11:0] + 12'h247;
  assign sel_297631 = $signed({1'h0, add_297527}) < $signed({1'h0, sel_297529}) ? add_297527 : sel_297529;
  assign array_index_297660 = set1_unflattened[8'h95];
  assign array_index_297663 = set2_unflattened[8'h95];
  assign add_297667 = array_index_297252[11:1] + 11'h79d;
  assign sel_297669 = $signed({1'h0, add_297565, array_index_297150[0]}) < $signed({1'h0, sel_297567}) ? {add_297565, array_index_297150[0]} : sel_297567;
  assign add_297671 = array_index_297255[11:1] + 11'h79d;
  assign sel_297673 = $signed({1'h0, add_297569, array_index_297153[0]}) < $signed({1'h0, sel_297571}) ? {add_297569, array_index_297153[0]} : sel_297571;
  assign add_297675 = array_index_297354[11:1] + 11'h347;
  assign sel_297677 = $signed({1'h0, add_297573, array_index_297252[0]}) < $signed({1'h0, sel_297575}) ? {add_297573, array_index_297252[0]} : sel_297575;
  assign add_297679 = array_index_297357[11:1] + 11'h347;
  assign sel_297681 = $signed({1'h0, add_297577, array_index_297255[0]}) < $signed({1'h0, sel_297579}) ? {add_297577, array_index_297255[0]} : sel_297579;
  assign add_297683 = array_index_297456[11:3] + 9'h0bd;
  assign sel_297686 = $signed({1'h0, add_297581, array_index_297354[2:0]}) < $signed({1'h0, sel_297584}) ? {add_297581, array_index_297354[2:0]} : sel_297584;
  assign add_297688 = array_index_297459[11:3] + 9'h0bd;
  assign sel_297691 = $signed({1'h0, add_297586, array_index_297357[2:0]}) < $signed({1'h0, sel_297589}) ? {add_297586, array_index_297357[2:0]} : sel_297589;
  assign add_297693 = array_index_297558[11:1] + 11'h247;
  assign sel_297696 = $signed({1'h0, add_297591, array_index_297456[0]}) < $signed({1'h0, sel_297594}) ? {add_297591, array_index_297456[0]} : sel_297594;
  assign add_297698 = array_index_297561[11:1] + 11'h247;
  assign sel_297701 = $signed({1'h0, add_297596, array_index_297459[0]}) < $signed({1'h0, sel_297599}) ? {add_297596, array_index_297459[0]} : sel_297599;
  assign add_297726 = array_index_297660[11:0] + 12'h247;
  assign sel_297728 = $signed({1'h0, add_297624}) < $signed({1'h0, sel_297626}) ? add_297624 : sel_297626;
  assign add_297731 = array_index_297663[11:0] + 12'h247;
  assign sel_297733 = $signed({1'h0, add_297629}) < $signed({1'h0, sel_297631}) ? add_297629 : sel_297631;
  assign array_index_297762 = set1_unflattened[8'h96];
  assign array_index_297765 = set2_unflattened[8'h96];
  assign add_297769 = array_index_297354[11:1] + 11'h79d;
  assign sel_297771 = $signed({1'h0, add_297667, array_index_297252[0]}) < $signed({1'h0, sel_297669}) ? {add_297667, array_index_297252[0]} : sel_297669;
  assign add_297773 = array_index_297357[11:1] + 11'h79d;
  assign sel_297775 = $signed({1'h0, add_297671, array_index_297255[0]}) < $signed({1'h0, sel_297673}) ? {add_297671, array_index_297255[0]} : sel_297673;
  assign add_297777 = array_index_297456[11:1] + 11'h347;
  assign sel_297779 = $signed({1'h0, add_297675, array_index_297354[0]}) < $signed({1'h0, sel_297677}) ? {add_297675, array_index_297354[0]} : sel_297677;
  assign add_297781 = array_index_297459[11:1] + 11'h347;
  assign sel_297783 = $signed({1'h0, add_297679, array_index_297357[0]}) < $signed({1'h0, sel_297681}) ? {add_297679, array_index_297357[0]} : sel_297681;
  assign add_297785 = array_index_297558[11:3] + 9'h0bd;
  assign sel_297788 = $signed({1'h0, add_297683, array_index_297456[2:0]}) < $signed({1'h0, sel_297686}) ? {add_297683, array_index_297456[2:0]} : sel_297686;
  assign add_297790 = array_index_297561[11:3] + 9'h0bd;
  assign sel_297793 = $signed({1'h0, add_297688, array_index_297459[2:0]}) < $signed({1'h0, sel_297691}) ? {add_297688, array_index_297459[2:0]} : sel_297691;
  assign add_297795 = array_index_297660[11:1] + 11'h247;
  assign sel_297798 = $signed({1'h0, add_297693, array_index_297558[0]}) < $signed({1'h0, sel_297696}) ? {add_297693, array_index_297558[0]} : sel_297696;
  assign add_297800 = array_index_297663[11:1] + 11'h247;
  assign sel_297803 = $signed({1'h0, add_297698, array_index_297561[0]}) < $signed({1'h0, sel_297701}) ? {add_297698, array_index_297561[0]} : sel_297701;
  assign add_297828 = array_index_297762[11:0] + 12'h247;
  assign sel_297830 = $signed({1'h0, add_297726}) < $signed({1'h0, sel_297728}) ? add_297726 : sel_297728;
  assign add_297833 = array_index_297765[11:0] + 12'h247;
  assign sel_297835 = $signed({1'h0, add_297731}) < $signed({1'h0, sel_297733}) ? add_297731 : sel_297733;
  assign array_index_297864 = set1_unflattened[8'h97];
  assign array_index_297867 = set2_unflattened[8'h97];
  assign add_297871 = array_index_297456[11:1] + 11'h79d;
  assign sel_297873 = $signed({1'h0, add_297769, array_index_297354[0]}) < $signed({1'h0, sel_297771}) ? {add_297769, array_index_297354[0]} : sel_297771;
  assign add_297875 = array_index_297459[11:1] + 11'h79d;
  assign sel_297877 = $signed({1'h0, add_297773, array_index_297357[0]}) < $signed({1'h0, sel_297775}) ? {add_297773, array_index_297357[0]} : sel_297775;
  assign add_297879 = array_index_297558[11:1] + 11'h347;
  assign sel_297881 = $signed({1'h0, add_297777, array_index_297456[0]}) < $signed({1'h0, sel_297779}) ? {add_297777, array_index_297456[0]} : sel_297779;
  assign add_297883 = array_index_297561[11:1] + 11'h347;
  assign sel_297885 = $signed({1'h0, add_297781, array_index_297459[0]}) < $signed({1'h0, sel_297783}) ? {add_297781, array_index_297459[0]} : sel_297783;
  assign add_297887 = array_index_297660[11:3] + 9'h0bd;
  assign sel_297890 = $signed({1'h0, add_297785, array_index_297558[2:0]}) < $signed({1'h0, sel_297788}) ? {add_297785, array_index_297558[2:0]} : sel_297788;
  assign add_297892 = array_index_297663[11:3] + 9'h0bd;
  assign sel_297895 = $signed({1'h0, add_297790, array_index_297561[2:0]}) < $signed({1'h0, sel_297793}) ? {add_297790, array_index_297561[2:0]} : sel_297793;
  assign add_297897 = array_index_297762[11:1] + 11'h247;
  assign sel_297900 = $signed({1'h0, add_297795, array_index_297660[0]}) < $signed({1'h0, sel_297798}) ? {add_297795, array_index_297660[0]} : sel_297798;
  assign add_297902 = array_index_297765[11:1] + 11'h247;
  assign sel_297905 = $signed({1'h0, add_297800, array_index_297663[0]}) < $signed({1'h0, sel_297803}) ? {add_297800, array_index_297663[0]} : sel_297803;
  assign add_297930 = array_index_297864[11:0] + 12'h247;
  assign sel_297932 = $signed({1'h0, add_297828}) < $signed({1'h0, sel_297830}) ? add_297828 : sel_297830;
  assign add_297935 = array_index_297867[11:0] + 12'h247;
  assign sel_297937 = $signed({1'h0, add_297833}) < $signed({1'h0, sel_297835}) ? add_297833 : sel_297835;
  assign array_index_297966 = set1_unflattened[8'h98];
  assign array_index_297969 = set2_unflattened[8'h98];
  assign add_297973 = array_index_297558[11:1] + 11'h79d;
  assign sel_297975 = $signed({1'h0, add_297871, array_index_297456[0]}) < $signed({1'h0, sel_297873}) ? {add_297871, array_index_297456[0]} : sel_297873;
  assign add_297977 = array_index_297561[11:1] + 11'h79d;
  assign sel_297979 = $signed({1'h0, add_297875, array_index_297459[0]}) < $signed({1'h0, sel_297877}) ? {add_297875, array_index_297459[0]} : sel_297877;
  assign add_297981 = array_index_297660[11:1] + 11'h347;
  assign sel_297983 = $signed({1'h0, add_297879, array_index_297558[0]}) < $signed({1'h0, sel_297881}) ? {add_297879, array_index_297558[0]} : sel_297881;
  assign add_297985 = array_index_297663[11:1] + 11'h347;
  assign sel_297987 = $signed({1'h0, add_297883, array_index_297561[0]}) < $signed({1'h0, sel_297885}) ? {add_297883, array_index_297561[0]} : sel_297885;
  assign add_297989 = array_index_297762[11:3] + 9'h0bd;
  assign sel_297992 = $signed({1'h0, add_297887, array_index_297660[2:0]}) < $signed({1'h0, sel_297890}) ? {add_297887, array_index_297660[2:0]} : sel_297890;
  assign add_297994 = array_index_297765[11:3] + 9'h0bd;
  assign sel_297997 = $signed({1'h0, add_297892, array_index_297663[2:0]}) < $signed({1'h0, sel_297895}) ? {add_297892, array_index_297663[2:0]} : sel_297895;
  assign add_297999 = array_index_297864[11:1] + 11'h247;
  assign sel_298002 = $signed({1'h0, add_297897, array_index_297762[0]}) < $signed({1'h0, sel_297900}) ? {add_297897, array_index_297762[0]} : sel_297900;
  assign add_298004 = array_index_297867[11:1] + 11'h247;
  assign sel_298007 = $signed({1'h0, add_297902, array_index_297765[0]}) < $signed({1'h0, sel_297905}) ? {add_297902, array_index_297765[0]} : sel_297905;
  assign add_298032 = array_index_297966[11:0] + 12'h247;
  assign sel_298034 = $signed({1'h0, add_297930}) < $signed({1'h0, sel_297932}) ? add_297930 : sel_297932;
  assign add_298037 = array_index_297969[11:0] + 12'h247;
  assign sel_298039 = $signed({1'h0, add_297935}) < $signed({1'h0, sel_297937}) ? add_297935 : sel_297937;
  assign array_index_298068 = set1_unflattened[8'h99];
  assign array_index_298071 = set2_unflattened[8'h99];
  assign add_298075 = array_index_297660[11:1] + 11'h79d;
  assign sel_298077 = $signed({1'h0, add_297973, array_index_297558[0]}) < $signed({1'h0, sel_297975}) ? {add_297973, array_index_297558[0]} : sel_297975;
  assign add_298079 = array_index_297663[11:1] + 11'h79d;
  assign sel_298081 = $signed({1'h0, add_297977, array_index_297561[0]}) < $signed({1'h0, sel_297979}) ? {add_297977, array_index_297561[0]} : sel_297979;
  assign add_298083 = array_index_297762[11:1] + 11'h347;
  assign sel_298085 = $signed({1'h0, add_297981, array_index_297660[0]}) < $signed({1'h0, sel_297983}) ? {add_297981, array_index_297660[0]} : sel_297983;
  assign add_298087 = array_index_297765[11:1] + 11'h347;
  assign sel_298089 = $signed({1'h0, add_297985, array_index_297663[0]}) < $signed({1'h0, sel_297987}) ? {add_297985, array_index_297663[0]} : sel_297987;
  assign add_298091 = array_index_297864[11:3] + 9'h0bd;
  assign sel_298094 = $signed({1'h0, add_297989, array_index_297762[2:0]}) < $signed({1'h0, sel_297992}) ? {add_297989, array_index_297762[2:0]} : sel_297992;
  assign add_298096 = array_index_297867[11:3] + 9'h0bd;
  assign sel_298099 = $signed({1'h0, add_297994, array_index_297765[2:0]}) < $signed({1'h0, sel_297997}) ? {add_297994, array_index_297765[2:0]} : sel_297997;
  assign add_298101 = array_index_297966[11:1] + 11'h247;
  assign sel_298104 = $signed({1'h0, add_297999, array_index_297864[0]}) < $signed({1'h0, sel_298002}) ? {add_297999, array_index_297864[0]} : sel_298002;
  assign add_298106 = array_index_297969[11:1] + 11'h247;
  assign sel_298109 = $signed({1'h0, add_298004, array_index_297867[0]}) < $signed({1'h0, sel_298007}) ? {add_298004, array_index_297867[0]} : sel_298007;
  assign add_298134 = array_index_298068[11:0] + 12'h247;
  assign sel_298136 = $signed({1'h0, add_298032}) < $signed({1'h0, sel_298034}) ? add_298032 : sel_298034;
  assign add_298139 = array_index_298071[11:0] + 12'h247;
  assign sel_298141 = $signed({1'h0, add_298037}) < $signed({1'h0, sel_298039}) ? add_298037 : sel_298039;
  assign array_index_298170 = set1_unflattened[8'h9a];
  assign array_index_298173 = set2_unflattened[8'h9a];
  assign add_298177 = array_index_297762[11:1] + 11'h79d;
  assign sel_298179 = $signed({1'h0, add_298075, array_index_297660[0]}) < $signed({1'h0, sel_298077}) ? {add_298075, array_index_297660[0]} : sel_298077;
  assign add_298181 = array_index_297765[11:1] + 11'h79d;
  assign sel_298183 = $signed({1'h0, add_298079, array_index_297663[0]}) < $signed({1'h0, sel_298081}) ? {add_298079, array_index_297663[0]} : sel_298081;
  assign add_298185 = array_index_297864[11:1] + 11'h347;
  assign sel_298187 = $signed({1'h0, add_298083, array_index_297762[0]}) < $signed({1'h0, sel_298085}) ? {add_298083, array_index_297762[0]} : sel_298085;
  assign add_298189 = array_index_297867[11:1] + 11'h347;
  assign sel_298191 = $signed({1'h0, add_298087, array_index_297765[0]}) < $signed({1'h0, sel_298089}) ? {add_298087, array_index_297765[0]} : sel_298089;
  assign add_298193 = array_index_297966[11:3] + 9'h0bd;
  assign sel_298196 = $signed({1'h0, add_298091, array_index_297864[2:0]}) < $signed({1'h0, sel_298094}) ? {add_298091, array_index_297864[2:0]} : sel_298094;
  assign add_298198 = array_index_297969[11:3] + 9'h0bd;
  assign sel_298201 = $signed({1'h0, add_298096, array_index_297867[2:0]}) < $signed({1'h0, sel_298099}) ? {add_298096, array_index_297867[2:0]} : sel_298099;
  assign add_298203 = array_index_298068[11:1] + 11'h247;
  assign sel_298206 = $signed({1'h0, add_298101, array_index_297966[0]}) < $signed({1'h0, sel_298104}) ? {add_298101, array_index_297966[0]} : sel_298104;
  assign add_298208 = array_index_298071[11:1] + 11'h247;
  assign sel_298211 = $signed({1'h0, add_298106, array_index_297969[0]}) < $signed({1'h0, sel_298109}) ? {add_298106, array_index_297969[0]} : sel_298109;
  assign add_298236 = array_index_298170[11:0] + 12'h247;
  assign sel_298238 = $signed({1'h0, add_298134}) < $signed({1'h0, sel_298136}) ? add_298134 : sel_298136;
  assign add_298241 = array_index_298173[11:0] + 12'h247;
  assign sel_298243 = $signed({1'h0, add_298139}) < $signed({1'h0, sel_298141}) ? add_298139 : sel_298141;
  assign array_index_298272 = set1_unflattened[8'h9b];
  assign array_index_298275 = set2_unflattened[8'h9b];
  assign add_298279 = array_index_297864[11:1] + 11'h79d;
  assign sel_298281 = $signed({1'h0, add_298177, array_index_297762[0]}) < $signed({1'h0, sel_298179}) ? {add_298177, array_index_297762[0]} : sel_298179;
  assign add_298283 = array_index_297867[11:1] + 11'h79d;
  assign sel_298285 = $signed({1'h0, add_298181, array_index_297765[0]}) < $signed({1'h0, sel_298183}) ? {add_298181, array_index_297765[0]} : sel_298183;
  assign add_298287 = array_index_297966[11:1] + 11'h347;
  assign sel_298289 = $signed({1'h0, add_298185, array_index_297864[0]}) < $signed({1'h0, sel_298187}) ? {add_298185, array_index_297864[0]} : sel_298187;
  assign add_298291 = array_index_297969[11:1] + 11'h347;
  assign sel_298293 = $signed({1'h0, add_298189, array_index_297867[0]}) < $signed({1'h0, sel_298191}) ? {add_298189, array_index_297867[0]} : sel_298191;
  assign add_298295 = array_index_298068[11:3] + 9'h0bd;
  assign sel_298298 = $signed({1'h0, add_298193, array_index_297966[2:0]}) < $signed({1'h0, sel_298196}) ? {add_298193, array_index_297966[2:0]} : sel_298196;
  assign add_298300 = array_index_298071[11:3] + 9'h0bd;
  assign sel_298303 = $signed({1'h0, add_298198, array_index_297969[2:0]}) < $signed({1'h0, sel_298201}) ? {add_298198, array_index_297969[2:0]} : sel_298201;
  assign add_298305 = array_index_298170[11:1] + 11'h247;
  assign sel_298308 = $signed({1'h0, add_298203, array_index_298068[0]}) < $signed({1'h0, sel_298206}) ? {add_298203, array_index_298068[0]} : sel_298206;
  assign add_298310 = array_index_298173[11:1] + 11'h247;
  assign sel_298313 = $signed({1'h0, add_298208, array_index_298071[0]}) < $signed({1'h0, sel_298211}) ? {add_298208, array_index_298071[0]} : sel_298211;
  assign add_298338 = array_index_298272[11:0] + 12'h247;
  assign sel_298340 = $signed({1'h0, add_298236}) < $signed({1'h0, sel_298238}) ? add_298236 : sel_298238;
  assign add_298343 = array_index_298275[11:0] + 12'h247;
  assign sel_298345 = $signed({1'h0, add_298241}) < $signed({1'h0, sel_298243}) ? add_298241 : sel_298243;
  assign array_index_298374 = set1_unflattened[8'h9c];
  assign array_index_298377 = set2_unflattened[8'h9c];
  assign add_298381 = array_index_297966[11:1] + 11'h79d;
  assign sel_298383 = $signed({1'h0, add_298279, array_index_297864[0]}) < $signed({1'h0, sel_298281}) ? {add_298279, array_index_297864[0]} : sel_298281;
  assign add_298385 = array_index_297969[11:1] + 11'h79d;
  assign sel_298387 = $signed({1'h0, add_298283, array_index_297867[0]}) < $signed({1'h0, sel_298285}) ? {add_298283, array_index_297867[0]} : sel_298285;
  assign add_298389 = array_index_298068[11:1] + 11'h347;
  assign sel_298391 = $signed({1'h0, add_298287, array_index_297966[0]}) < $signed({1'h0, sel_298289}) ? {add_298287, array_index_297966[0]} : sel_298289;
  assign add_298393 = array_index_298071[11:1] + 11'h347;
  assign sel_298395 = $signed({1'h0, add_298291, array_index_297969[0]}) < $signed({1'h0, sel_298293}) ? {add_298291, array_index_297969[0]} : sel_298293;
  assign add_298397 = array_index_298170[11:3] + 9'h0bd;
  assign sel_298400 = $signed({1'h0, add_298295, array_index_298068[2:0]}) < $signed({1'h0, sel_298298}) ? {add_298295, array_index_298068[2:0]} : sel_298298;
  assign add_298402 = array_index_298173[11:3] + 9'h0bd;
  assign sel_298405 = $signed({1'h0, add_298300, array_index_298071[2:0]}) < $signed({1'h0, sel_298303}) ? {add_298300, array_index_298071[2:0]} : sel_298303;
  assign add_298407 = array_index_298272[11:1] + 11'h247;
  assign sel_298410 = $signed({1'h0, add_298305, array_index_298170[0]}) < $signed({1'h0, sel_298308}) ? {add_298305, array_index_298170[0]} : sel_298308;
  assign add_298412 = array_index_298275[11:1] + 11'h247;
  assign sel_298415 = $signed({1'h0, add_298310, array_index_298173[0]}) < $signed({1'h0, sel_298313}) ? {add_298310, array_index_298173[0]} : sel_298313;
  assign add_298440 = array_index_298374[11:0] + 12'h247;
  assign sel_298442 = $signed({1'h0, add_298338}) < $signed({1'h0, sel_298340}) ? add_298338 : sel_298340;
  assign add_298445 = array_index_298377[11:0] + 12'h247;
  assign sel_298447 = $signed({1'h0, add_298343}) < $signed({1'h0, sel_298345}) ? add_298343 : sel_298345;
  assign array_index_298476 = set1_unflattened[8'h9d];
  assign array_index_298479 = set2_unflattened[8'h9d];
  assign add_298483 = array_index_298068[11:1] + 11'h79d;
  assign sel_298485 = $signed({1'h0, add_298381, array_index_297966[0]}) < $signed({1'h0, sel_298383}) ? {add_298381, array_index_297966[0]} : sel_298383;
  assign add_298487 = array_index_298071[11:1] + 11'h79d;
  assign sel_298489 = $signed({1'h0, add_298385, array_index_297969[0]}) < $signed({1'h0, sel_298387}) ? {add_298385, array_index_297969[0]} : sel_298387;
  assign add_298491 = array_index_298170[11:1] + 11'h347;
  assign sel_298493 = $signed({1'h0, add_298389, array_index_298068[0]}) < $signed({1'h0, sel_298391}) ? {add_298389, array_index_298068[0]} : sel_298391;
  assign add_298495 = array_index_298173[11:1] + 11'h347;
  assign sel_298497 = $signed({1'h0, add_298393, array_index_298071[0]}) < $signed({1'h0, sel_298395}) ? {add_298393, array_index_298071[0]} : sel_298395;
  assign add_298499 = array_index_298272[11:3] + 9'h0bd;
  assign sel_298502 = $signed({1'h0, add_298397, array_index_298170[2:0]}) < $signed({1'h0, sel_298400}) ? {add_298397, array_index_298170[2:0]} : sel_298400;
  assign add_298504 = array_index_298275[11:3] + 9'h0bd;
  assign sel_298507 = $signed({1'h0, add_298402, array_index_298173[2:0]}) < $signed({1'h0, sel_298405}) ? {add_298402, array_index_298173[2:0]} : sel_298405;
  assign add_298509 = array_index_298374[11:1] + 11'h247;
  assign sel_298512 = $signed({1'h0, add_298407, array_index_298272[0]}) < $signed({1'h0, sel_298410}) ? {add_298407, array_index_298272[0]} : sel_298410;
  assign add_298514 = array_index_298377[11:1] + 11'h247;
  assign sel_298517 = $signed({1'h0, add_298412, array_index_298275[0]}) < $signed({1'h0, sel_298415}) ? {add_298412, array_index_298275[0]} : sel_298415;
  assign add_298542 = array_index_298476[11:0] + 12'h247;
  assign sel_298544 = $signed({1'h0, add_298440}) < $signed({1'h0, sel_298442}) ? add_298440 : sel_298442;
  assign add_298547 = array_index_298479[11:0] + 12'h247;
  assign sel_298549 = $signed({1'h0, add_298445}) < $signed({1'h0, sel_298447}) ? add_298445 : sel_298447;
  assign array_index_298578 = set1_unflattened[8'h9e];
  assign array_index_298581 = set2_unflattened[8'h9e];
  assign add_298585 = array_index_298170[11:1] + 11'h79d;
  assign sel_298587 = $signed({1'h0, add_298483, array_index_298068[0]}) < $signed({1'h0, sel_298485}) ? {add_298483, array_index_298068[0]} : sel_298485;
  assign add_298589 = array_index_298173[11:1] + 11'h79d;
  assign sel_298591 = $signed({1'h0, add_298487, array_index_298071[0]}) < $signed({1'h0, sel_298489}) ? {add_298487, array_index_298071[0]} : sel_298489;
  assign add_298593 = array_index_298272[11:1] + 11'h347;
  assign sel_298595 = $signed({1'h0, add_298491, array_index_298170[0]}) < $signed({1'h0, sel_298493}) ? {add_298491, array_index_298170[0]} : sel_298493;
  assign add_298597 = array_index_298275[11:1] + 11'h347;
  assign sel_298599 = $signed({1'h0, add_298495, array_index_298173[0]}) < $signed({1'h0, sel_298497}) ? {add_298495, array_index_298173[0]} : sel_298497;
  assign add_298601 = array_index_298374[11:3] + 9'h0bd;
  assign sel_298604 = $signed({1'h0, add_298499, array_index_298272[2:0]}) < $signed({1'h0, sel_298502}) ? {add_298499, array_index_298272[2:0]} : sel_298502;
  assign add_298606 = array_index_298377[11:3] + 9'h0bd;
  assign sel_298609 = $signed({1'h0, add_298504, array_index_298275[2:0]}) < $signed({1'h0, sel_298507}) ? {add_298504, array_index_298275[2:0]} : sel_298507;
  assign add_298611 = array_index_298476[11:1] + 11'h247;
  assign sel_298614 = $signed({1'h0, add_298509, array_index_298374[0]}) < $signed({1'h0, sel_298512}) ? {add_298509, array_index_298374[0]} : sel_298512;
  assign add_298616 = array_index_298479[11:1] + 11'h247;
  assign sel_298619 = $signed({1'h0, add_298514, array_index_298377[0]}) < $signed({1'h0, sel_298517}) ? {add_298514, array_index_298377[0]} : sel_298517;
  assign add_298644 = array_index_298578[11:0] + 12'h247;
  assign sel_298646 = $signed({1'h0, add_298542}) < $signed({1'h0, sel_298544}) ? add_298542 : sel_298544;
  assign add_298649 = array_index_298581[11:0] + 12'h247;
  assign sel_298651 = $signed({1'h0, add_298547}) < $signed({1'h0, sel_298549}) ? add_298547 : sel_298549;
  assign array_index_298680 = set1_unflattened[8'h9f];
  assign array_index_298683 = set2_unflattened[8'h9f];
  assign add_298687 = array_index_298272[11:1] + 11'h79d;
  assign sel_298689 = $signed({1'h0, add_298585, array_index_298170[0]}) < $signed({1'h0, sel_298587}) ? {add_298585, array_index_298170[0]} : sel_298587;
  assign add_298691 = array_index_298275[11:1] + 11'h79d;
  assign sel_298693 = $signed({1'h0, add_298589, array_index_298173[0]}) < $signed({1'h0, sel_298591}) ? {add_298589, array_index_298173[0]} : sel_298591;
  assign add_298695 = array_index_298374[11:1] + 11'h347;
  assign sel_298697 = $signed({1'h0, add_298593, array_index_298272[0]}) < $signed({1'h0, sel_298595}) ? {add_298593, array_index_298272[0]} : sel_298595;
  assign add_298699 = array_index_298377[11:1] + 11'h347;
  assign sel_298701 = $signed({1'h0, add_298597, array_index_298275[0]}) < $signed({1'h0, sel_298599}) ? {add_298597, array_index_298275[0]} : sel_298599;
  assign add_298703 = array_index_298476[11:3] + 9'h0bd;
  assign sel_298706 = $signed({1'h0, add_298601, array_index_298374[2:0]}) < $signed({1'h0, sel_298604}) ? {add_298601, array_index_298374[2:0]} : sel_298604;
  assign add_298708 = array_index_298479[11:3] + 9'h0bd;
  assign sel_298711 = $signed({1'h0, add_298606, array_index_298377[2:0]}) < $signed({1'h0, sel_298609}) ? {add_298606, array_index_298377[2:0]} : sel_298609;
  assign add_298713 = array_index_298578[11:1] + 11'h247;
  assign sel_298716 = $signed({1'h0, add_298611, array_index_298476[0]}) < $signed({1'h0, sel_298614}) ? {add_298611, array_index_298476[0]} : sel_298614;
  assign add_298718 = array_index_298581[11:1] + 11'h247;
  assign sel_298721 = $signed({1'h0, add_298616, array_index_298479[0]}) < $signed({1'h0, sel_298619}) ? {add_298616, array_index_298479[0]} : sel_298619;
  assign add_298746 = array_index_298680[11:0] + 12'h247;
  assign sel_298748 = $signed({1'h0, add_298644}) < $signed({1'h0, sel_298646}) ? add_298644 : sel_298646;
  assign add_298751 = array_index_298683[11:0] + 12'h247;
  assign sel_298753 = $signed({1'h0, add_298649}) < $signed({1'h0, sel_298651}) ? add_298649 : sel_298651;
  assign array_index_298782 = set1_unflattened[8'ha0];
  assign array_index_298785 = set2_unflattened[8'ha0];
  assign add_298789 = array_index_298374[11:1] + 11'h79d;
  assign sel_298791 = $signed({1'h0, add_298687, array_index_298272[0]}) < $signed({1'h0, sel_298689}) ? {add_298687, array_index_298272[0]} : sel_298689;
  assign add_298793 = array_index_298377[11:1] + 11'h79d;
  assign sel_298795 = $signed({1'h0, add_298691, array_index_298275[0]}) < $signed({1'h0, sel_298693}) ? {add_298691, array_index_298275[0]} : sel_298693;
  assign add_298797 = array_index_298476[11:1] + 11'h347;
  assign sel_298799 = $signed({1'h0, add_298695, array_index_298374[0]}) < $signed({1'h0, sel_298697}) ? {add_298695, array_index_298374[0]} : sel_298697;
  assign add_298801 = array_index_298479[11:1] + 11'h347;
  assign sel_298803 = $signed({1'h0, add_298699, array_index_298377[0]}) < $signed({1'h0, sel_298701}) ? {add_298699, array_index_298377[0]} : sel_298701;
  assign add_298805 = array_index_298578[11:3] + 9'h0bd;
  assign sel_298808 = $signed({1'h0, add_298703, array_index_298476[2:0]}) < $signed({1'h0, sel_298706}) ? {add_298703, array_index_298476[2:0]} : sel_298706;
  assign add_298810 = array_index_298581[11:3] + 9'h0bd;
  assign sel_298813 = $signed({1'h0, add_298708, array_index_298479[2:0]}) < $signed({1'h0, sel_298711}) ? {add_298708, array_index_298479[2:0]} : sel_298711;
  assign add_298815 = array_index_298680[11:1] + 11'h247;
  assign sel_298818 = $signed({1'h0, add_298713, array_index_298578[0]}) < $signed({1'h0, sel_298716}) ? {add_298713, array_index_298578[0]} : sel_298716;
  assign add_298820 = array_index_298683[11:1] + 11'h247;
  assign sel_298823 = $signed({1'h0, add_298718, array_index_298581[0]}) < $signed({1'h0, sel_298721}) ? {add_298718, array_index_298581[0]} : sel_298721;
  assign add_298848 = array_index_298782[11:0] + 12'h247;
  assign sel_298850 = $signed({1'h0, add_298746}) < $signed({1'h0, sel_298748}) ? add_298746 : sel_298748;
  assign add_298853 = array_index_298785[11:0] + 12'h247;
  assign sel_298855 = $signed({1'h0, add_298751}) < $signed({1'h0, sel_298753}) ? add_298751 : sel_298753;
  assign array_index_298884 = set1_unflattened[8'ha1];
  assign array_index_298887 = set2_unflattened[8'ha1];
  assign add_298891 = array_index_298476[11:1] + 11'h79d;
  assign sel_298893 = $signed({1'h0, add_298789, array_index_298374[0]}) < $signed({1'h0, sel_298791}) ? {add_298789, array_index_298374[0]} : sel_298791;
  assign add_298895 = array_index_298479[11:1] + 11'h79d;
  assign sel_298897 = $signed({1'h0, add_298793, array_index_298377[0]}) < $signed({1'h0, sel_298795}) ? {add_298793, array_index_298377[0]} : sel_298795;
  assign add_298899 = array_index_298578[11:1] + 11'h347;
  assign sel_298901 = $signed({1'h0, add_298797, array_index_298476[0]}) < $signed({1'h0, sel_298799}) ? {add_298797, array_index_298476[0]} : sel_298799;
  assign add_298903 = array_index_298581[11:1] + 11'h347;
  assign sel_298905 = $signed({1'h0, add_298801, array_index_298479[0]}) < $signed({1'h0, sel_298803}) ? {add_298801, array_index_298479[0]} : sel_298803;
  assign add_298907 = array_index_298680[11:3] + 9'h0bd;
  assign sel_298910 = $signed({1'h0, add_298805, array_index_298578[2:0]}) < $signed({1'h0, sel_298808}) ? {add_298805, array_index_298578[2:0]} : sel_298808;
  assign add_298912 = array_index_298683[11:3] + 9'h0bd;
  assign sel_298915 = $signed({1'h0, add_298810, array_index_298581[2:0]}) < $signed({1'h0, sel_298813}) ? {add_298810, array_index_298581[2:0]} : sel_298813;
  assign add_298917 = array_index_298782[11:1] + 11'h247;
  assign sel_298920 = $signed({1'h0, add_298815, array_index_298680[0]}) < $signed({1'h0, sel_298818}) ? {add_298815, array_index_298680[0]} : sel_298818;
  assign add_298922 = array_index_298785[11:1] + 11'h247;
  assign sel_298925 = $signed({1'h0, add_298820, array_index_298683[0]}) < $signed({1'h0, sel_298823}) ? {add_298820, array_index_298683[0]} : sel_298823;
  assign add_298950 = array_index_298884[11:0] + 12'h247;
  assign sel_298952 = $signed({1'h0, add_298848}) < $signed({1'h0, sel_298850}) ? add_298848 : sel_298850;
  assign add_298955 = array_index_298887[11:0] + 12'h247;
  assign sel_298957 = $signed({1'h0, add_298853}) < $signed({1'h0, sel_298855}) ? add_298853 : sel_298855;
  assign array_index_298986 = set1_unflattened[8'ha2];
  assign array_index_298989 = set2_unflattened[8'ha2];
  assign add_298993 = array_index_298578[11:1] + 11'h79d;
  assign sel_298995 = $signed({1'h0, add_298891, array_index_298476[0]}) < $signed({1'h0, sel_298893}) ? {add_298891, array_index_298476[0]} : sel_298893;
  assign add_298997 = array_index_298581[11:1] + 11'h79d;
  assign sel_298999 = $signed({1'h0, add_298895, array_index_298479[0]}) < $signed({1'h0, sel_298897}) ? {add_298895, array_index_298479[0]} : sel_298897;
  assign add_299001 = array_index_298680[11:1] + 11'h347;
  assign sel_299003 = $signed({1'h0, add_298899, array_index_298578[0]}) < $signed({1'h0, sel_298901}) ? {add_298899, array_index_298578[0]} : sel_298901;
  assign add_299005 = array_index_298683[11:1] + 11'h347;
  assign sel_299007 = $signed({1'h0, add_298903, array_index_298581[0]}) < $signed({1'h0, sel_298905}) ? {add_298903, array_index_298581[0]} : sel_298905;
  assign add_299009 = array_index_298782[11:3] + 9'h0bd;
  assign sel_299012 = $signed({1'h0, add_298907, array_index_298680[2:0]}) < $signed({1'h0, sel_298910}) ? {add_298907, array_index_298680[2:0]} : sel_298910;
  assign add_299014 = array_index_298785[11:3] + 9'h0bd;
  assign sel_299017 = $signed({1'h0, add_298912, array_index_298683[2:0]}) < $signed({1'h0, sel_298915}) ? {add_298912, array_index_298683[2:0]} : sel_298915;
  assign add_299019 = array_index_298884[11:1] + 11'h247;
  assign sel_299022 = $signed({1'h0, add_298917, array_index_298782[0]}) < $signed({1'h0, sel_298920}) ? {add_298917, array_index_298782[0]} : sel_298920;
  assign add_299024 = array_index_298887[11:1] + 11'h247;
  assign sel_299027 = $signed({1'h0, add_298922, array_index_298785[0]}) < $signed({1'h0, sel_298925}) ? {add_298922, array_index_298785[0]} : sel_298925;
  assign add_299052 = array_index_298986[11:0] + 12'h247;
  assign sel_299054 = $signed({1'h0, add_298950}) < $signed({1'h0, sel_298952}) ? add_298950 : sel_298952;
  assign add_299057 = array_index_298989[11:0] + 12'h247;
  assign sel_299059 = $signed({1'h0, add_298955}) < $signed({1'h0, sel_298957}) ? add_298955 : sel_298957;
  assign array_index_299088 = set1_unflattened[8'ha3];
  assign array_index_299091 = set2_unflattened[8'ha3];
  assign add_299095 = array_index_298680[11:1] + 11'h79d;
  assign sel_299097 = $signed({1'h0, add_298993, array_index_298578[0]}) < $signed({1'h0, sel_298995}) ? {add_298993, array_index_298578[0]} : sel_298995;
  assign add_299099 = array_index_298683[11:1] + 11'h79d;
  assign sel_299101 = $signed({1'h0, add_298997, array_index_298581[0]}) < $signed({1'h0, sel_298999}) ? {add_298997, array_index_298581[0]} : sel_298999;
  assign add_299103 = array_index_298782[11:1] + 11'h347;
  assign sel_299105 = $signed({1'h0, add_299001, array_index_298680[0]}) < $signed({1'h0, sel_299003}) ? {add_299001, array_index_298680[0]} : sel_299003;
  assign add_299107 = array_index_298785[11:1] + 11'h347;
  assign sel_299109 = $signed({1'h0, add_299005, array_index_298683[0]}) < $signed({1'h0, sel_299007}) ? {add_299005, array_index_298683[0]} : sel_299007;
  assign add_299111 = array_index_298884[11:3] + 9'h0bd;
  assign sel_299114 = $signed({1'h0, add_299009, array_index_298782[2:0]}) < $signed({1'h0, sel_299012}) ? {add_299009, array_index_298782[2:0]} : sel_299012;
  assign add_299116 = array_index_298887[11:3] + 9'h0bd;
  assign sel_299119 = $signed({1'h0, add_299014, array_index_298785[2:0]}) < $signed({1'h0, sel_299017}) ? {add_299014, array_index_298785[2:0]} : sel_299017;
  assign add_299121 = array_index_298986[11:1] + 11'h247;
  assign sel_299124 = $signed({1'h0, add_299019, array_index_298884[0]}) < $signed({1'h0, sel_299022}) ? {add_299019, array_index_298884[0]} : sel_299022;
  assign add_299126 = array_index_298989[11:1] + 11'h247;
  assign sel_299129 = $signed({1'h0, add_299024, array_index_298887[0]}) < $signed({1'h0, sel_299027}) ? {add_299024, array_index_298887[0]} : sel_299027;
  assign add_299154 = array_index_299088[11:0] + 12'h247;
  assign sel_299156 = $signed({1'h0, add_299052}) < $signed({1'h0, sel_299054}) ? add_299052 : sel_299054;
  assign add_299159 = array_index_299091[11:0] + 12'h247;
  assign sel_299161 = $signed({1'h0, add_299057}) < $signed({1'h0, sel_299059}) ? add_299057 : sel_299059;
  assign array_index_299190 = set1_unflattened[8'ha4];
  assign array_index_299193 = set2_unflattened[8'ha4];
  assign add_299197 = array_index_298782[11:1] + 11'h79d;
  assign sel_299199 = $signed({1'h0, add_299095, array_index_298680[0]}) < $signed({1'h0, sel_299097}) ? {add_299095, array_index_298680[0]} : sel_299097;
  assign add_299201 = array_index_298785[11:1] + 11'h79d;
  assign sel_299203 = $signed({1'h0, add_299099, array_index_298683[0]}) < $signed({1'h0, sel_299101}) ? {add_299099, array_index_298683[0]} : sel_299101;
  assign add_299205 = array_index_298884[11:1] + 11'h347;
  assign sel_299207 = $signed({1'h0, add_299103, array_index_298782[0]}) < $signed({1'h0, sel_299105}) ? {add_299103, array_index_298782[0]} : sel_299105;
  assign add_299209 = array_index_298887[11:1] + 11'h347;
  assign sel_299211 = $signed({1'h0, add_299107, array_index_298785[0]}) < $signed({1'h0, sel_299109}) ? {add_299107, array_index_298785[0]} : sel_299109;
  assign add_299213 = array_index_298986[11:3] + 9'h0bd;
  assign sel_299216 = $signed({1'h0, add_299111, array_index_298884[2:0]}) < $signed({1'h0, sel_299114}) ? {add_299111, array_index_298884[2:0]} : sel_299114;
  assign add_299218 = array_index_298989[11:3] + 9'h0bd;
  assign sel_299221 = $signed({1'h0, add_299116, array_index_298887[2:0]}) < $signed({1'h0, sel_299119}) ? {add_299116, array_index_298887[2:0]} : sel_299119;
  assign add_299223 = array_index_299088[11:1] + 11'h247;
  assign sel_299226 = $signed({1'h0, add_299121, array_index_298986[0]}) < $signed({1'h0, sel_299124}) ? {add_299121, array_index_298986[0]} : sel_299124;
  assign add_299228 = array_index_299091[11:1] + 11'h247;
  assign sel_299231 = $signed({1'h0, add_299126, array_index_298989[0]}) < $signed({1'h0, sel_299129}) ? {add_299126, array_index_298989[0]} : sel_299129;
  assign add_299256 = array_index_299190[11:0] + 12'h247;
  assign sel_299258 = $signed({1'h0, add_299154}) < $signed({1'h0, sel_299156}) ? add_299154 : sel_299156;
  assign add_299261 = array_index_299193[11:0] + 12'h247;
  assign sel_299263 = $signed({1'h0, add_299159}) < $signed({1'h0, sel_299161}) ? add_299159 : sel_299161;
  assign array_index_299292 = set1_unflattened[8'ha5];
  assign array_index_299295 = set2_unflattened[8'ha5];
  assign add_299299 = array_index_298884[11:1] + 11'h79d;
  assign sel_299301 = $signed({1'h0, add_299197, array_index_298782[0]}) < $signed({1'h0, sel_299199}) ? {add_299197, array_index_298782[0]} : sel_299199;
  assign add_299303 = array_index_298887[11:1] + 11'h79d;
  assign sel_299305 = $signed({1'h0, add_299201, array_index_298785[0]}) < $signed({1'h0, sel_299203}) ? {add_299201, array_index_298785[0]} : sel_299203;
  assign add_299307 = array_index_298986[11:1] + 11'h347;
  assign sel_299309 = $signed({1'h0, add_299205, array_index_298884[0]}) < $signed({1'h0, sel_299207}) ? {add_299205, array_index_298884[0]} : sel_299207;
  assign add_299311 = array_index_298989[11:1] + 11'h347;
  assign sel_299313 = $signed({1'h0, add_299209, array_index_298887[0]}) < $signed({1'h0, sel_299211}) ? {add_299209, array_index_298887[0]} : sel_299211;
  assign add_299315 = array_index_299088[11:3] + 9'h0bd;
  assign sel_299318 = $signed({1'h0, add_299213, array_index_298986[2:0]}) < $signed({1'h0, sel_299216}) ? {add_299213, array_index_298986[2:0]} : sel_299216;
  assign add_299320 = array_index_299091[11:3] + 9'h0bd;
  assign sel_299323 = $signed({1'h0, add_299218, array_index_298989[2:0]}) < $signed({1'h0, sel_299221}) ? {add_299218, array_index_298989[2:0]} : sel_299221;
  assign add_299325 = array_index_299190[11:1] + 11'h247;
  assign sel_299328 = $signed({1'h0, add_299223, array_index_299088[0]}) < $signed({1'h0, sel_299226}) ? {add_299223, array_index_299088[0]} : sel_299226;
  assign add_299330 = array_index_299193[11:1] + 11'h247;
  assign sel_299333 = $signed({1'h0, add_299228, array_index_299091[0]}) < $signed({1'h0, sel_299231}) ? {add_299228, array_index_299091[0]} : sel_299231;
  assign add_299358 = array_index_299292[11:0] + 12'h247;
  assign sel_299360 = $signed({1'h0, add_299256}) < $signed({1'h0, sel_299258}) ? add_299256 : sel_299258;
  assign add_299363 = array_index_299295[11:0] + 12'h247;
  assign sel_299365 = $signed({1'h0, add_299261}) < $signed({1'h0, sel_299263}) ? add_299261 : sel_299263;
  assign array_index_299394 = set1_unflattened[8'ha6];
  assign array_index_299397 = set2_unflattened[8'ha6];
  assign add_299401 = array_index_298986[11:1] + 11'h79d;
  assign sel_299403 = $signed({1'h0, add_299299, array_index_298884[0]}) < $signed({1'h0, sel_299301}) ? {add_299299, array_index_298884[0]} : sel_299301;
  assign add_299405 = array_index_298989[11:1] + 11'h79d;
  assign sel_299407 = $signed({1'h0, add_299303, array_index_298887[0]}) < $signed({1'h0, sel_299305}) ? {add_299303, array_index_298887[0]} : sel_299305;
  assign add_299409 = array_index_299088[11:1] + 11'h347;
  assign sel_299411 = $signed({1'h0, add_299307, array_index_298986[0]}) < $signed({1'h0, sel_299309}) ? {add_299307, array_index_298986[0]} : sel_299309;
  assign add_299413 = array_index_299091[11:1] + 11'h347;
  assign sel_299415 = $signed({1'h0, add_299311, array_index_298989[0]}) < $signed({1'h0, sel_299313}) ? {add_299311, array_index_298989[0]} : sel_299313;
  assign add_299417 = array_index_299190[11:3] + 9'h0bd;
  assign sel_299420 = $signed({1'h0, add_299315, array_index_299088[2:0]}) < $signed({1'h0, sel_299318}) ? {add_299315, array_index_299088[2:0]} : sel_299318;
  assign add_299422 = array_index_299193[11:3] + 9'h0bd;
  assign sel_299425 = $signed({1'h0, add_299320, array_index_299091[2:0]}) < $signed({1'h0, sel_299323}) ? {add_299320, array_index_299091[2:0]} : sel_299323;
  assign add_299427 = array_index_299292[11:1] + 11'h247;
  assign sel_299430 = $signed({1'h0, add_299325, array_index_299190[0]}) < $signed({1'h0, sel_299328}) ? {add_299325, array_index_299190[0]} : sel_299328;
  assign add_299432 = array_index_299295[11:1] + 11'h247;
  assign sel_299435 = $signed({1'h0, add_299330, array_index_299193[0]}) < $signed({1'h0, sel_299333}) ? {add_299330, array_index_299193[0]} : sel_299333;
  assign add_299460 = array_index_299394[11:0] + 12'h247;
  assign sel_299462 = $signed({1'h0, add_299358}) < $signed({1'h0, sel_299360}) ? add_299358 : sel_299360;
  assign add_299465 = array_index_299397[11:0] + 12'h247;
  assign sel_299467 = $signed({1'h0, add_299363}) < $signed({1'h0, sel_299365}) ? add_299363 : sel_299365;
  assign array_index_299496 = set1_unflattened[8'ha7];
  assign array_index_299499 = set2_unflattened[8'ha7];
  assign add_299503 = array_index_299088[11:1] + 11'h79d;
  assign sel_299505 = $signed({1'h0, add_299401, array_index_298986[0]}) < $signed({1'h0, sel_299403}) ? {add_299401, array_index_298986[0]} : sel_299403;
  assign add_299507 = array_index_299091[11:1] + 11'h79d;
  assign sel_299509 = $signed({1'h0, add_299405, array_index_298989[0]}) < $signed({1'h0, sel_299407}) ? {add_299405, array_index_298989[0]} : sel_299407;
  assign add_299511 = array_index_299190[11:1] + 11'h347;
  assign sel_299513 = $signed({1'h0, add_299409, array_index_299088[0]}) < $signed({1'h0, sel_299411}) ? {add_299409, array_index_299088[0]} : sel_299411;
  assign add_299515 = array_index_299193[11:1] + 11'h347;
  assign sel_299517 = $signed({1'h0, add_299413, array_index_299091[0]}) < $signed({1'h0, sel_299415}) ? {add_299413, array_index_299091[0]} : sel_299415;
  assign add_299519 = array_index_299292[11:3] + 9'h0bd;
  assign sel_299522 = $signed({1'h0, add_299417, array_index_299190[2:0]}) < $signed({1'h0, sel_299420}) ? {add_299417, array_index_299190[2:0]} : sel_299420;
  assign add_299524 = array_index_299295[11:3] + 9'h0bd;
  assign sel_299527 = $signed({1'h0, add_299422, array_index_299193[2:0]}) < $signed({1'h0, sel_299425}) ? {add_299422, array_index_299193[2:0]} : sel_299425;
  assign add_299529 = array_index_299394[11:1] + 11'h247;
  assign sel_299532 = $signed({1'h0, add_299427, array_index_299292[0]}) < $signed({1'h0, sel_299430}) ? {add_299427, array_index_299292[0]} : sel_299430;
  assign add_299534 = array_index_299397[11:1] + 11'h247;
  assign sel_299537 = $signed({1'h0, add_299432, array_index_299295[0]}) < $signed({1'h0, sel_299435}) ? {add_299432, array_index_299295[0]} : sel_299435;
  assign add_299562 = array_index_299496[11:0] + 12'h247;
  assign sel_299564 = $signed({1'h0, add_299460}) < $signed({1'h0, sel_299462}) ? add_299460 : sel_299462;
  assign add_299567 = array_index_299499[11:0] + 12'h247;
  assign sel_299569 = $signed({1'h0, add_299465}) < $signed({1'h0, sel_299467}) ? add_299465 : sel_299467;
  assign array_index_299598 = set1_unflattened[8'ha8];
  assign array_index_299601 = set2_unflattened[8'ha8];
  assign add_299605 = array_index_299190[11:1] + 11'h79d;
  assign sel_299607 = $signed({1'h0, add_299503, array_index_299088[0]}) < $signed({1'h0, sel_299505}) ? {add_299503, array_index_299088[0]} : sel_299505;
  assign add_299609 = array_index_299193[11:1] + 11'h79d;
  assign sel_299611 = $signed({1'h0, add_299507, array_index_299091[0]}) < $signed({1'h0, sel_299509}) ? {add_299507, array_index_299091[0]} : sel_299509;
  assign add_299613 = array_index_299292[11:1] + 11'h347;
  assign sel_299615 = $signed({1'h0, add_299511, array_index_299190[0]}) < $signed({1'h0, sel_299513}) ? {add_299511, array_index_299190[0]} : sel_299513;
  assign add_299617 = array_index_299295[11:1] + 11'h347;
  assign sel_299619 = $signed({1'h0, add_299515, array_index_299193[0]}) < $signed({1'h0, sel_299517}) ? {add_299515, array_index_299193[0]} : sel_299517;
  assign add_299621 = array_index_299394[11:3] + 9'h0bd;
  assign sel_299624 = $signed({1'h0, add_299519, array_index_299292[2:0]}) < $signed({1'h0, sel_299522}) ? {add_299519, array_index_299292[2:0]} : sel_299522;
  assign add_299626 = array_index_299397[11:3] + 9'h0bd;
  assign sel_299629 = $signed({1'h0, add_299524, array_index_299295[2:0]}) < $signed({1'h0, sel_299527}) ? {add_299524, array_index_299295[2:0]} : sel_299527;
  assign add_299631 = array_index_299496[11:1] + 11'h247;
  assign sel_299634 = $signed({1'h0, add_299529, array_index_299394[0]}) < $signed({1'h0, sel_299532}) ? {add_299529, array_index_299394[0]} : sel_299532;
  assign add_299636 = array_index_299499[11:1] + 11'h247;
  assign sel_299639 = $signed({1'h0, add_299534, array_index_299397[0]}) < $signed({1'h0, sel_299537}) ? {add_299534, array_index_299397[0]} : sel_299537;
  assign add_299664 = array_index_299598[11:0] + 12'h247;
  assign sel_299666 = $signed({1'h0, add_299562}) < $signed({1'h0, sel_299564}) ? add_299562 : sel_299564;
  assign add_299669 = array_index_299601[11:0] + 12'h247;
  assign sel_299671 = $signed({1'h0, add_299567}) < $signed({1'h0, sel_299569}) ? add_299567 : sel_299569;
  assign array_index_299700 = set1_unflattened[8'ha9];
  assign array_index_299703 = set2_unflattened[8'ha9];
  assign add_299707 = array_index_299292[11:1] + 11'h79d;
  assign sel_299709 = $signed({1'h0, add_299605, array_index_299190[0]}) < $signed({1'h0, sel_299607}) ? {add_299605, array_index_299190[0]} : sel_299607;
  assign add_299711 = array_index_299295[11:1] + 11'h79d;
  assign sel_299713 = $signed({1'h0, add_299609, array_index_299193[0]}) < $signed({1'h0, sel_299611}) ? {add_299609, array_index_299193[0]} : sel_299611;
  assign add_299715 = array_index_299394[11:1] + 11'h347;
  assign sel_299717 = $signed({1'h0, add_299613, array_index_299292[0]}) < $signed({1'h0, sel_299615}) ? {add_299613, array_index_299292[0]} : sel_299615;
  assign add_299719 = array_index_299397[11:1] + 11'h347;
  assign sel_299721 = $signed({1'h0, add_299617, array_index_299295[0]}) < $signed({1'h0, sel_299619}) ? {add_299617, array_index_299295[0]} : sel_299619;
  assign add_299723 = array_index_299496[11:3] + 9'h0bd;
  assign sel_299726 = $signed({1'h0, add_299621, array_index_299394[2:0]}) < $signed({1'h0, sel_299624}) ? {add_299621, array_index_299394[2:0]} : sel_299624;
  assign add_299728 = array_index_299499[11:3] + 9'h0bd;
  assign sel_299731 = $signed({1'h0, add_299626, array_index_299397[2:0]}) < $signed({1'h0, sel_299629}) ? {add_299626, array_index_299397[2:0]} : sel_299629;
  assign add_299733 = array_index_299598[11:1] + 11'h247;
  assign sel_299736 = $signed({1'h0, add_299631, array_index_299496[0]}) < $signed({1'h0, sel_299634}) ? {add_299631, array_index_299496[0]} : sel_299634;
  assign add_299738 = array_index_299601[11:1] + 11'h247;
  assign sel_299741 = $signed({1'h0, add_299636, array_index_299499[0]}) < $signed({1'h0, sel_299639}) ? {add_299636, array_index_299499[0]} : sel_299639;
  assign add_299766 = array_index_299700[11:0] + 12'h247;
  assign sel_299768 = $signed({1'h0, add_299664}) < $signed({1'h0, sel_299666}) ? add_299664 : sel_299666;
  assign add_299771 = array_index_299703[11:0] + 12'h247;
  assign sel_299773 = $signed({1'h0, add_299669}) < $signed({1'h0, sel_299671}) ? add_299669 : sel_299671;
  assign array_index_299802 = set1_unflattened[8'haa];
  assign array_index_299805 = set2_unflattened[8'haa];
  assign add_299809 = array_index_299394[11:1] + 11'h79d;
  assign sel_299811 = $signed({1'h0, add_299707, array_index_299292[0]}) < $signed({1'h0, sel_299709}) ? {add_299707, array_index_299292[0]} : sel_299709;
  assign add_299813 = array_index_299397[11:1] + 11'h79d;
  assign sel_299815 = $signed({1'h0, add_299711, array_index_299295[0]}) < $signed({1'h0, sel_299713}) ? {add_299711, array_index_299295[0]} : sel_299713;
  assign add_299817 = array_index_299496[11:1] + 11'h347;
  assign sel_299819 = $signed({1'h0, add_299715, array_index_299394[0]}) < $signed({1'h0, sel_299717}) ? {add_299715, array_index_299394[0]} : sel_299717;
  assign add_299821 = array_index_299499[11:1] + 11'h347;
  assign sel_299823 = $signed({1'h0, add_299719, array_index_299397[0]}) < $signed({1'h0, sel_299721}) ? {add_299719, array_index_299397[0]} : sel_299721;
  assign add_299825 = array_index_299598[11:3] + 9'h0bd;
  assign sel_299828 = $signed({1'h0, add_299723, array_index_299496[2:0]}) < $signed({1'h0, sel_299726}) ? {add_299723, array_index_299496[2:0]} : sel_299726;
  assign add_299830 = array_index_299601[11:3] + 9'h0bd;
  assign sel_299833 = $signed({1'h0, add_299728, array_index_299499[2:0]}) < $signed({1'h0, sel_299731}) ? {add_299728, array_index_299499[2:0]} : sel_299731;
  assign add_299835 = array_index_299700[11:1] + 11'h247;
  assign sel_299838 = $signed({1'h0, add_299733, array_index_299598[0]}) < $signed({1'h0, sel_299736}) ? {add_299733, array_index_299598[0]} : sel_299736;
  assign add_299840 = array_index_299703[11:1] + 11'h247;
  assign sel_299843 = $signed({1'h0, add_299738, array_index_299601[0]}) < $signed({1'h0, sel_299741}) ? {add_299738, array_index_299601[0]} : sel_299741;
  assign add_299868 = array_index_299802[11:0] + 12'h247;
  assign sel_299870 = $signed({1'h0, add_299766}) < $signed({1'h0, sel_299768}) ? add_299766 : sel_299768;
  assign add_299873 = array_index_299805[11:0] + 12'h247;
  assign sel_299875 = $signed({1'h0, add_299771}) < $signed({1'h0, sel_299773}) ? add_299771 : sel_299773;
  assign array_index_299904 = set1_unflattened[8'hab];
  assign array_index_299907 = set2_unflattened[8'hab];
  assign add_299911 = array_index_299496[11:1] + 11'h79d;
  assign sel_299913 = $signed({1'h0, add_299809, array_index_299394[0]}) < $signed({1'h0, sel_299811}) ? {add_299809, array_index_299394[0]} : sel_299811;
  assign add_299915 = array_index_299499[11:1] + 11'h79d;
  assign sel_299917 = $signed({1'h0, add_299813, array_index_299397[0]}) < $signed({1'h0, sel_299815}) ? {add_299813, array_index_299397[0]} : sel_299815;
  assign add_299919 = array_index_299598[11:1] + 11'h347;
  assign sel_299921 = $signed({1'h0, add_299817, array_index_299496[0]}) < $signed({1'h0, sel_299819}) ? {add_299817, array_index_299496[0]} : sel_299819;
  assign add_299923 = array_index_299601[11:1] + 11'h347;
  assign sel_299925 = $signed({1'h0, add_299821, array_index_299499[0]}) < $signed({1'h0, sel_299823}) ? {add_299821, array_index_299499[0]} : sel_299823;
  assign add_299927 = array_index_299700[11:3] + 9'h0bd;
  assign sel_299930 = $signed({1'h0, add_299825, array_index_299598[2:0]}) < $signed({1'h0, sel_299828}) ? {add_299825, array_index_299598[2:0]} : sel_299828;
  assign add_299932 = array_index_299703[11:3] + 9'h0bd;
  assign sel_299935 = $signed({1'h0, add_299830, array_index_299601[2:0]}) < $signed({1'h0, sel_299833}) ? {add_299830, array_index_299601[2:0]} : sel_299833;
  assign add_299937 = array_index_299802[11:1] + 11'h247;
  assign sel_299940 = $signed({1'h0, add_299835, array_index_299700[0]}) < $signed({1'h0, sel_299838}) ? {add_299835, array_index_299700[0]} : sel_299838;
  assign add_299942 = array_index_299805[11:1] + 11'h247;
  assign sel_299945 = $signed({1'h0, add_299840, array_index_299703[0]}) < $signed({1'h0, sel_299843}) ? {add_299840, array_index_299703[0]} : sel_299843;
  assign add_299970 = array_index_299904[11:0] + 12'h247;
  assign sel_299972 = $signed({1'h0, add_299868}) < $signed({1'h0, sel_299870}) ? add_299868 : sel_299870;
  assign add_299975 = array_index_299907[11:0] + 12'h247;
  assign sel_299977 = $signed({1'h0, add_299873}) < $signed({1'h0, sel_299875}) ? add_299873 : sel_299875;
  assign array_index_300006 = set1_unflattened[8'hac];
  assign array_index_300009 = set2_unflattened[8'hac];
  assign add_300013 = array_index_299598[11:1] + 11'h79d;
  assign sel_300015 = $signed({1'h0, add_299911, array_index_299496[0]}) < $signed({1'h0, sel_299913}) ? {add_299911, array_index_299496[0]} : sel_299913;
  assign add_300017 = array_index_299601[11:1] + 11'h79d;
  assign sel_300019 = $signed({1'h0, add_299915, array_index_299499[0]}) < $signed({1'h0, sel_299917}) ? {add_299915, array_index_299499[0]} : sel_299917;
  assign add_300021 = array_index_299700[11:1] + 11'h347;
  assign sel_300023 = $signed({1'h0, add_299919, array_index_299598[0]}) < $signed({1'h0, sel_299921}) ? {add_299919, array_index_299598[0]} : sel_299921;
  assign add_300025 = array_index_299703[11:1] + 11'h347;
  assign sel_300027 = $signed({1'h0, add_299923, array_index_299601[0]}) < $signed({1'h0, sel_299925}) ? {add_299923, array_index_299601[0]} : sel_299925;
  assign add_300029 = array_index_299802[11:3] + 9'h0bd;
  assign sel_300032 = $signed({1'h0, add_299927, array_index_299700[2:0]}) < $signed({1'h0, sel_299930}) ? {add_299927, array_index_299700[2:0]} : sel_299930;
  assign add_300034 = array_index_299805[11:3] + 9'h0bd;
  assign sel_300037 = $signed({1'h0, add_299932, array_index_299703[2:0]}) < $signed({1'h0, sel_299935}) ? {add_299932, array_index_299703[2:0]} : sel_299935;
  assign add_300039 = array_index_299904[11:1] + 11'h247;
  assign sel_300042 = $signed({1'h0, add_299937, array_index_299802[0]}) < $signed({1'h0, sel_299940}) ? {add_299937, array_index_299802[0]} : sel_299940;
  assign add_300044 = array_index_299907[11:1] + 11'h247;
  assign sel_300047 = $signed({1'h0, add_299942, array_index_299805[0]}) < $signed({1'h0, sel_299945}) ? {add_299942, array_index_299805[0]} : sel_299945;
  assign add_300072 = array_index_300006[11:0] + 12'h247;
  assign sel_300074 = $signed({1'h0, add_299970}) < $signed({1'h0, sel_299972}) ? add_299970 : sel_299972;
  assign add_300077 = array_index_300009[11:0] + 12'h247;
  assign sel_300079 = $signed({1'h0, add_299975}) < $signed({1'h0, sel_299977}) ? add_299975 : sel_299977;
  assign array_index_300108 = set1_unflattened[8'had];
  assign array_index_300111 = set2_unflattened[8'had];
  assign add_300115 = array_index_299700[11:1] + 11'h79d;
  assign sel_300117 = $signed({1'h0, add_300013, array_index_299598[0]}) < $signed({1'h0, sel_300015}) ? {add_300013, array_index_299598[0]} : sel_300015;
  assign add_300119 = array_index_299703[11:1] + 11'h79d;
  assign sel_300121 = $signed({1'h0, add_300017, array_index_299601[0]}) < $signed({1'h0, sel_300019}) ? {add_300017, array_index_299601[0]} : sel_300019;
  assign add_300123 = array_index_299802[11:1] + 11'h347;
  assign sel_300125 = $signed({1'h0, add_300021, array_index_299700[0]}) < $signed({1'h0, sel_300023}) ? {add_300021, array_index_299700[0]} : sel_300023;
  assign add_300127 = array_index_299805[11:1] + 11'h347;
  assign sel_300129 = $signed({1'h0, add_300025, array_index_299703[0]}) < $signed({1'h0, sel_300027}) ? {add_300025, array_index_299703[0]} : sel_300027;
  assign add_300131 = array_index_299904[11:3] + 9'h0bd;
  assign sel_300134 = $signed({1'h0, add_300029, array_index_299802[2:0]}) < $signed({1'h0, sel_300032}) ? {add_300029, array_index_299802[2:0]} : sel_300032;
  assign add_300136 = array_index_299907[11:3] + 9'h0bd;
  assign sel_300139 = $signed({1'h0, add_300034, array_index_299805[2:0]}) < $signed({1'h0, sel_300037}) ? {add_300034, array_index_299805[2:0]} : sel_300037;
  assign add_300141 = array_index_300006[11:1] + 11'h247;
  assign sel_300144 = $signed({1'h0, add_300039, array_index_299904[0]}) < $signed({1'h0, sel_300042}) ? {add_300039, array_index_299904[0]} : sel_300042;
  assign add_300146 = array_index_300009[11:1] + 11'h247;
  assign sel_300149 = $signed({1'h0, add_300044, array_index_299907[0]}) < $signed({1'h0, sel_300047}) ? {add_300044, array_index_299907[0]} : sel_300047;
  assign add_300174 = array_index_300108[11:0] + 12'h247;
  assign sel_300176 = $signed({1'h0, add_300072}) < $signed({1'h0, sel_300074}) ? add_300072 : sel_300074;
  assign add_300179 = array_index_300111[11:0] + 12'h247;
  assign sel_300181 = $signed({1'h0, add_300077}) < $signed({1'h0, sel_300079}) ? add_300077 : sel_300079;
  assign array_index_300210 = set1_unflattened[8'hae];
  assign array_index_300213 = set2_unflattened[8'hae];
  assign add_300217 = array_index_299802[11:1] + 11'h79d;
  assign sel_300219 = $signed({1'h0, add_300115, array_index_299700[0]}) < $signed({1'h0, sel_300117}) ? {add_300115, array_index_299700[0]} : sel_300117;
  assign add_300221 = array_index_299805[11:1] + 11'h79d;
  assign sel_300223 = $signed({1'h0, add_300119, array_index_299703[0]}) < $signed({1'h0, sel_300121}) ? {add_300119, array_index_299703[0]} : sel_300121;
  assign add_300225 = array_index_299904[11:1] + 11'h347;
  assign sel_300227 = $signed({1'h0, add_300123, array_index_299802[0]}) < $signed({1'h0, sel_300125}) ? {add_300123, array_index_299802[0]} : sel_300125;
  assign add_300229 = array_index_299907[11:1] + 11'h347;
  assign sel_300231 = $signed({1'h0, add_300127, array_index_299805[0]}) < $signed({1'h0, sel_300129}) ? {add_300127, array_index_299805[0]} : sel_300129;
  assign add_300233 = array_index_300006[11:3] + 9'h0bd;
  assign sel_300236 = $signed({1'h0, add_300131, array_index_299904[2:0]}) < $signed({1'h0, sel_300134}) ? {add_300131, array_index_299904[2:0]} : sel_300134;
  assign add_300238 = array_index_300009[11:3] + 9'h0bd;
  assign sel_300241 = $signed({1'h0, add_300136, array_index_299907[2:0]}) < $signed({1'h0, sel_300139}) ? {add_300136, array_index_299907[2:0]} : sel_300139;
  assign add_300243 = array_index_300108[11:1] + 11'h247;
  assign sel_300246 = $signed({1'h0, add_300141, array_index_300006[0]}) < $signed({1'h0, sel_300144}) ? {add_300141, array_index_300006[0]} : sel_300144;
  assign add_300248 = array_index_300111[11:1] + 11'h247;
  assign sel_300251 = $signed({1'h0, add_300146, array_index_300009[0]}) < $signed({1'h0, sel_300149}) ? {add_300146, array_index_300009[0]} : sel_300149;
  assign add_300276 = array_index_300210[11:0] + 12'h247;
  assign sel_300278 = $signed({1'h0, add_300174}) < $signed({1'h0, sel_300176}) ? add_300174 : sel_300176;
  assign add_300281 = array_index_300213[11:0] + 12'h247;
  assign sel_300283 = $signed({1'h0, add_300179}) < $signed({1'h0, sel_300181}) ? add_300179 : sel_300181;
  assign array_index_300312 = set1_unflattened[8'haf];
  assign array_index_300315 = set2_unflattened[8'haf];
  assign add_300319 = array_index_299904[11:1] + 11'h79d;
  assign sel_300321 = $signed({1'h0, add_300217, array_index_299802[0]}) < $signed({1'h0, sel_300219}) ? {add_300217, array_index_299802[0]} : sel_300219;
  assign add_300323 = array_index_299907[11:1] + 11'h79d;
  assign sel_300325 = $signed({1'h0, add_300221, array_index_299805[0]}) < $signed({1'h0, sel_300223}) ? {add_300221, array_index_299805[0]} : sel_300223;
  assign add_300327 = array_index_300006[11:1] + 11'h347;
  assign sel_300329 = $signed({1'h0, add_300225, array_index_299904[0]}) < $signed({1'h0, sel_300227}) ? {add_300225, array_index_299904[0]} : sel_300227;
  assign add_300331 = array_index_300009[11:1] + 11'h347;
  assign sel_300333 = $signed({1'h0, add_300229, array_index_299907[0]}) < $signed({1'h0, sel_300231}) ? {add_300229, array_index_299907[0]} : sel_300231;
  assign add_300335 = array_index_300108[11:3] + 9'h0bd;
  assign sel_300338 = $signed({1'h0, add_300233, array_index_300006[2:0]}) < $signed({1'h0, sel_300236}) ? {add_300233, array_index_300006[2:0]} : sel_300236;
  assign add_300340 = array_index_300111[11:3] + 9'h0bd;
  assign sel_300343 = $signed({1'h0, add_300238, array_index_300009[2:0]}) < $signed({1'h0, sel_300241}) ? {add_300238, array_index_300009[2:0]} : sel_300241;
  assign add_300345 = array_index_300210[11:1] + 11'h247;
  assign sel_300348 = $signed({1'h0, add_300243, array_index_300108[0]}) < $signed({1'h0, sel_300246}) ? {add_300243, array_index_300108[0]} : sel_300246;
  assign add_300350 = array_index_300213[11:1] + 11'h247;
  assign sel_300353 = $signed({1'h0, add_300248, array_index_300111[0]}) < $signed({1'h0, sel_300251}) ? {add_300248, array_index_300111[0]} : sel_300251;
  assign add_300378 = array_index_300312[11:0] + 12'h247;
  assign sel_300380 = $signed({1'h0, add_300276}) < $signed({1'h0, sel_300278}) ? add_300276 : sel_300278;
  assign add_300383 = array_index_300315[11:0] + 12'h247;
  assign sel_300385 = $signed({1'h0, add_300281}) < $signed({1'h0, sel_300283}) ? add_300281 : sel_300283;
  assign array_index_300414 = set1_unflattened[8'hb0];
  assign array_index_300417 = set2_unflattened[8'hb0];
  assign add_300421 = array_index_300006[11:1] + 11'h79d;
  assign sel_300423 = $signed({1'h0, add_300319, array_index_299904[0]}) < $signed({1'h0, sel_300321}) ? {add_300319, array_index_299904[0]} : sel_300321;
  assign add_300425 = array_index_300009[11:1] + 11'h79d;
  assign sel_300427 = $signed({1'h0, add_300323, array_index_299907[0]}) < $signed({1'h0, sel_300325}) ? {add_300323, array_index_299907[0]} : sel_300325;
  assign add_300429 = array_index_300108[11:1] + 11'h347;
  assign sel_300431 = $signed({1'h0, add_300327, array_index_300006[0]}) < $signed({1'h0, sel_300329}) ? {add_300327, array_index_300006[0]} : sel_300329;
  assign add_300433 = array_index_300111[11:1] + 11'h347;
  assign sel_300435 = $signed({1'h0, add_300331, array_index_300009[0]}) < $signed({1'h0, sel_300333}) ? {add_300331, array_index_300009[0]} : sel_300333;
  assign add_300437 = array_index_300210[11:3] + 9'h0bd;
  assign sel_300440 = $signed({1'h0, add_300335, array_index_300108[2:0]}) < $signed({1'h0, sel_300338}) ? {add_300335, array_index_300108[2:0]} : sel_300338;
  assign add_300442 = array_index_300213[11:3] + 9'h0bd;
  assign sel_300445 = $signed({1'h0, add_300340, array_index_300111[2:0]}) < $signed({1'h0, sel_300343}) ? {add_300340, array_index_300111[2:0]} : sel_300343;
  assign add_300447 = array_index_300312[11:1] + 11'h247;
  assign sel_300450 = $signed({1'h0, add_300345, array_index_300210[0]}) < $signed({1'h0, sel_300348}) ? {add_300345, array_index_300210[0]} : sel_300348;
  assign add_300452 = array_index_300315[11:1] + 11'h247;
  assign sel_300455 = $signed({1'h0, add_300350, array_index_300213[0]}) < $signed({1'h0, sel_300353}) ? {add_300350, array_index_300213[0]} : sel_300353;
  assign add_300480 = array_index_300414[11:0] + 12'h247;
  assign sel_300482 = $signed({1'h0, add_300378}) < $signed({1'h0, sel_300380}) ? add_300378 : sel_300380;
  assign add_300485 = array_index_300417[11:0] + 12'h247;
  assign sel_300487 = $signed({1'h0, add_300383}) < $signed({1'h0, sel_300385}) ? add_300383 : sel_300385;
  assign array_index_300516 = set1_unflattened[8'hb1];
  assign array_index_300519 = set2_unflattened[8'hb1];
  assign add_300523 = array_index_300108[11:1] + 11'h79d;
  assign sel_300525 = $signed({1'h0, add_300421, array_index_300006[0]}) < $signed({1'h0, sel_300423}) ? {add_300421, array_index_300006[0]} : sel_300423;
  assign add_300527 = array_index_300111[11:1] + 11'h79d;
  assign sel_300529 = $signed({1'h0, add_300425, array_index_300009[0]}) < $signed({1'h0, sel_300427}) ? {add_300425, array_index_300009[0]} : sel_300427;
  assign add_300531 = array_index_300210[11:1] + 11'h347;
  assign sel_300533 = $signed({1'h0, add_300429, array_index_300108[0]}) < $signed({1'h0, sel_300431}) ? {add_300429, array_index_300108[0]} : sel_300431;
  assign add_300535 = array_index_300213[11:1] + 11'h347;
  assign sel_300537 = $signed({1'h0, add_300433, array_index_300111[0]}) < $signed({1'h0, sel_300435}) ? {add_300433, array_index_300111[0]} : sel_300435;
  assign add_300539 = array_index_300312[11:3] + 9'h0bd;
  assign sel_300542 = $signed({1'h0, add_300437, array_index_300210[2:0]}) < $signed({1'h0, sel_300440}) ? {add_300437, array_index_300210[2:0]} : sel_300440;
  assign add_300544 = array_index_300315[11:3] + 9'h0bd;
  assign sel_300547 = $signed({1'h0, add_300442, array_index_300213[2:0]}) < $signed({1'h0, sel_300445}) ? {add_300442, array_index_300213[2:0]} : sel_300445;
  assign add_300549 = array_index_300414[11:1] + 11'h247;
  assign sel_300552 = $signed({1'h0, add_300447, array_index_300312[0]}) < $signed({1'h0, sel_300450}) ? {add_300447, array_index_300312[0]} : sel_300450;
  assign add_300554 = array_index_300417[11:1] + 11'h247;
  assign sel_300557 = $signed({1'h0, add_300452, array_index_300315[0]}) < $signed({1'h0, sel_300455}) ? {add_300452, array_index_300315[0]} : sel_300455;
  assign add_300582 = array_index_300516[11:0] + 12'h247;
  assign sel_300584 = $signed({1'h0, add_300480}) < $signed({1'h0, sel_300482}) ? add_300480 : sel_300482;
  assign add_300587 = array_index_300519[11:0] + 12'h247;
  assign sel_300589 = $signed({1'h0, add_300485}) < $signed({1'h0, sel_300487}) ? add_300485 : sel_300487;
  assign array_index_300618 = set1_unflattened[8'hb2];
  assign array_index_300621 = set2_unflattened[8'hb2];
  assign add_300625 = array_index_300210[11:1] + 11'h79d;
  assign sel_300627 = $signed({1'h0, add_300523, array_index_300108[0]}) < $signed({1'h0, sel_300525}) ? {add_300523, array_index_300108[0]} : sel_300525;
  assign add_300629 = array_index_300213[11:1] + 11'h79d;
  assign sel_300631 = $signed({1'h0, add_300527, array_index_300111[0]}) < $signed({1'h0, sel_300529}) ? {add_300527, array_index_300111[0]} : sel_300529;
  assign add_300633 = array_index_300312[11:1] + 11'h347;
  assign sel_300635 = $signed({1'h0, add_300531, array_index_300210[0]}) < $signed({1'h0, sel_300533}) ? {add_300531, array_index_300210[0]} : sel_300533;
  assign add_300637 = array_index_300315[11:1] + 11'h347;
  assign sel_300639 = $signed({1'h0, add_300535, array_index_300213[0]}) < $signed({1'h0, sel_300537}) ? {add_300535, array_index_300213[0]} : sel_300537;
  assign add_300641 = array_index_300414[11:3] + 9'h0bd;
  assign sel_300644 = $signed({1'h0, add_300539, array_index_300312[2:0]}) < $signed({1'h0, sel_300542}) ? {add_300539, array_index_300312[2:0]} : sel_300542;
  assign add_300646 = array_index_300417[11:3] + 9'h0bd;
  assign sel_300649 = $signed({1'h0, add_300544, array_index_300315[2:0]}) < $signed({1'h0, sel_300547}) ? {add_300544, array_index_300315[2:0]} : sel_300547;
  assign add_300651 = array_index_300516[11:1] + 11'h247;
  assign sel_300654 = $signed({1'h0, add_300549, array_index_300414[0]}) < $signed({1'h0, sel_300552}) ? {add_300549, array_index_300414[0]} : sel_300552;
  assign add_300656 = array_index_300519[11:1] + 11'h247;
  assign sel_300659 = $signed({1'h0, add_300554, array_index_300417[0]}) < $signed({1'h0, sel_300557}) ? {add_300554, array_index_300417[0]} : sel_300557;
  assign add_300684 = array_index_300618[11:0] + 12'h247;
  assign sel_300686 = $signed({1'h0, add_300582}) < $signed({1'h0, sel_300584}) ? add_300582 : sel_300584;
  assign add_300689 = array_index_300621[11:0] + 12'h247;
  assign sel_300691 = $signed({1'h0, add_300587}) < $signed({1'h0, sel_300589}) ? add_300587 : sel_300589;
  assign array_index_300720 = set1_unflattened[8'hb3];
  assign array_index_300723 = set2_unflattened[8'hb3];
  assign add_300727 = array_index_300312[11:1] + 11'h79d;
  assign sel_300729 = $signed({1'h0, add_300625, array_index_300210[0]}) < $signed({1'h0, sel_300627}) ? {add_300625, array_index_300210[0]} : sel_300627;
  assign add_300731 = array_index_300315[11:1] + 11'h79d;
  assign sel_300733 = $signed({1'h0, add_300629, array_index_300213[0]}) < $signed({1'h0, sel_300631}) ? {add_300629, array_index_300213[0]} : sel_300631;
  assign add_300735 = array_index_300414[11:1] + 11'h347;
  assign sel_300737 = $signed({1'h0, add_300633, array_index_300312[0]}) < $signed({1'h0, sel_300635}) ? {add_300633, array_index_300312[0]} : sel_300635;
  assign add_300739 = array_index_300417[11:1] + 11'h347;
  assign sel_300741 = $signed({1'h0, add_300637, array_index_300315[0]}) < $signed({1'h0, sel_300639}) ? {add_300637, array_index_300315[0]} : sel_300639;
  assign add_300743 = array_index_300516[11:3] + 9'h0bd;
  assign sel_300746 = $signed({1'h0, add_300641, array_index_300414[2:0]}) < $signed({1'h0, sel_300644}) ? {add_300641, array_index_300414[2:0]} : sel_300644;
  assign add_300748 = array_index_300519[11:3] + 9'h0bd;
  assign sel_300751 = $signed({1'h0, add_300646, array_index_300417[2:0]}) < $signed({1'h0, sel_300649}) ? {add_300646, array_index_300417[2:0]} : sel_300649;
  assign add_300753 = array_index_300618[11:1] + 11'h247;
  assign sel_300756 = $signed({1'h0, add_300651, array_index_300516[0]}) < $signed({1'h0, sel_300654}) ? {add_300651, array_index_300516[0]} : sel_300654;
  assign add_300758 = array_index_300621[11:1] + 11'h247;
  assign sel_300761 = $signed({1'h0, add_300656, array_index_300519[0]}) < $signed({1'h0, sel_300659}) ? {add_300656, array_index_300519[0]} : sel_300659;
  assign add_300786 = array_index_300720[11:0] + 12'h247;
  assign sel_300788 = $signed({1'h0, add_300684}) < $signed({1'h0, sel_300686}) ? add_300684 : sel_300686;
  assign add_300791 = array_index_300723[11:0] + 12'h247;
  assign sel_300793 = $signed({1'h0, add_300689}) < $signed({1'h0, sel_300691}) ? add_300689 : sel_300691;
  assign array_index_300822 = set1_unflattened[8'hb4];
  assign array_index_300825 = set2_unflattened[8'hb4];
  assign add_300829 = array_index_300414[11:1] + 11'h79d;
  assign sel_300831 = $signed({1'h0, add_300727, array_index_300312[0]}) < $signed({1'h0, sel_300729}) ? {add_300727, array_index_300312[0]} : sel_300729;
  assign add_300833 = array_index_300417[11:1] + 11'h79d;
  assign sel_300835 = $signed({1'h0, add_300731, array_index_300315[0]}) < $signed({1'h0, sel_300733}) ? {add_300731, array_index_300315[0]} : sel_300733;
  assign add_300837 = array_index_300516[11:1] + 11'h347;
  assign sel_300839 = $signed({1'h0, add_300735, array_index_300414[0]}) < $signed({1'h0, sel_300737}) ? {add_300735, array_index_300414[0]} : sel_300737;
  assign add_300841 = array_index_300519[11:1] + 11'h347;
  assign sel_300843 = $signed({1'h0, add_300739, array_index_300417[0]}) < $signed({1'h0, sel_300741}) ? {add_300739, array_index_300417[0]} : sel_300741;
  assign add_300845 = array_index_300618[11:3] + 9'h0bd;
  assign sel_300848 = $signed({1'h0, add_300743, array_index_300516[2:0]}) < $signed({1'h0, sel_300746}) ? {add_300743, array_index_300516[2:0]} : sel_300746;
  assign add_300850 = array_index_300621[11:3] + 9'h0bd;
  assign sel_300853 = $signed({1'h0, add_300748, array_index_300519[2:0]}) < $signed({1'h0, sel_300751}) ? {add_300748, array_index_300519[2:0]} : sel_300751;
  assign add_300855 = array_index_300720[11:1] + 11'h247;
  assign sel_300858 = $signed({1'h0, add_300753, array_index_300618[0]}) < $signed({1'h0, sel_300756}) ? {add_300753, array_index_300618[0]} : sel_300756;
  assign add_300860 = array_index_300723[11:1] + 11'h247;
  assign sel_300863 = $signed({1'h0, add_300758, array_index_300621[0]}) < $signed({1'h0, sel_300761}) ? {add_300758, array_index_300621[0]} : sel_300761;
  assign add_300888 = array_index_300822[11:0] + 12'h247;
  assign sel_300890 = $signed({1'h0, add_300786}) < $signed({1'h0, sel_300788}) ? add_300786 : sel_300788;
  assign add_300893 = array_index_300825[11:0] + 12'h247;
  assign sel_300895 = $signed({1'h0, add_300791}) < $signed({1'h0, sel_300793}) ? add_300791 : sel_300793;
  assign array_index_300924 = set1_unflattened[8'hb5];
  assign array_index_300927 = set2_unflattened[8'hb5];
  assign add_300931 = array_index_300516[11:1] + 11'h79d;
  assign sel_300933 = $signed({1'h0, add_300829, array_index_300414[0]}) < $signed({1'h0, sel_300831}) ? {add_300829, array_index_300414[0]} : sel_300831;
  assign add_300935 = array_index_300519[11:1] + 11'h79d;
  assign sel_300937 = $signed({1'h0, add_300833, array_index_300417[0]}) < $signed({1'h0, sel_300835}) ? {add_300833, array_index_300417[0]} : sel_300835;
  assign add_300939 = array_index_300618[11:1] + 11'h347;
  assign sel_300941 = $signed({1'h0, add_300837, array_index_300516[0]}) < $signed({1'h0, sel_300839}) ? {add_300837, array_index_300516[0]} : sel_300839;
  assign add_300943 = array_index_300621[11:1] + 11'h347;
  assign sel_300945 = $signed({1'h0, add_300841, array_index_300519[0]}) < $signed({1'h0, sel_300843}) ? {add_300841, array_index_300519[0]} : sel_300843;
  assign add_300947 = array_index_300720[11:3] + 9'h0bd;
  assign sel_300950 = $signed({1'h0, add_300845, array_index_300618[2:0]}) < $signed({1'h0, sel_300848}) ? {add_300845, array_index_300618[2:0]} : sel_300848;
  assign add_300952 = array_index_300723[11:3] + 9'h0bd;
  assign sel_300955 = $signed({1'h0, add_300850, array_index_300621[2:0]}) < $signed({1'h0, sel_300853}) ? {add_300850, array_index_300621[2:0]} : sel_300853;
  assign add_300957 = array_index_300822[11:1] + 11'h247;
  assign sel_300960 = $signed({1'h0, add_300855, array_index_300720[0]}) < $signed({1'h0, sel_300858}) ? {add_300855, array_index_300720[0]} : sel_300858;
  assign add_300962 = array_index_300825[11:1] + 11'h247;
  assign sel_300965 = $signed({1'h0, add_300860, array_index_300723[0]}) < $signed({1'h0, sel_300863}) ? {add_300860, array_index_300723[0]} : sel_300863;
  assign add_300990 = array_index_300924[11:0] + 12'h247;
  assign sel_300992 = $signed({1'h0, add_300888}) < $signed({1'h0, sel_300890}) ? add_300888 : sel_300890;
  assign add_300995 = array_index_300927[11:0] + 12'h247;
  assign sel_300997 = $signed({1'h0, add_300893}) < $signed({1'h0, sel_300895}) ? add_300893 : sel_300895;
  assign array_index_301026 = set1_unflattened[8'hb6];
  assign array_index_301029 = set2_unflattened[8'hb6];
  assign add_301033 = array_index_300618[11:1] + 11'h79d;
  assign sel_301035 = $signed({1'h0, add_300931, array_index_300516[0]}) < $signed({1'h0, sel_300933}) ? {add_300931, array_index_300516[0]} : sel_300933;
  assign add_301037 = array_index_300621[11:1] + 11'h79d;
  assign sel_301039 = $signed({1'h0, add_300935, array_index_300519[0]}) < $signed({1'h0, sel_300937}) ? {add_300935, array_index_300519[0]} : sel_300937;
  assign add_301041 = array_index_300720[11:1] + 11'h347;
  assign sel_301043 = $signed({1'h0, add_300939, array_index_300618[0]}) < $signed({1'h0, sel_300941}) ? {add_300939, array_index_300618[0]} : sel_300941;
  assign add_301045 = array_index_300723[11:1] + 11'h347;
  assign sel_301047 = $signed({1'h0, add_300943, array_index_300621[0]}) < $signed({1'h0, sel_300945}) ? {add_300943, array_index_300621[0]} : sel_300945;
  assign add_301049 = array_index_300822[11:3] + 9'h0bd;
  assign sel_301052 = $signed({1'h0, add_300947, array_index_300720[2:0]}) < $signed({1'h0, sel_300950}) ? {add_300947, array_index_300720[2:0]} : sel_300950;
  assign add_301054 = array_index_300825[11:3] + 9'h0bd;
  assign sel_301057 = $signed({1'h0, add_300952, array_index_300723[2:0]}) < $signed({1'h0, sel_300955}) ? {add_300952, array_index_300723[2:0]} : sel_300955;
  assign add_301059 = array_index_300924[11:1] + 11'h247;
  assign sel_301062 = $signed({1'h0, add_300957, array_index_300822[0]}) < $signed({1'h0, sel_300960}) ? {add_300957, array_index_300822[0]} : sel_300960;
  assign add_301064 = array_index_300927[11:1] + 11'h247;
  assign sel_301067 = $signed({1'h0, add_300962, array_index_300825[0]}) < $signed({1'h0, sel_300965}) ? {add_300962, array_index_300825[0]} : sel_300965;
  assign add_301092 = array_index_301026[11:0] + 12'h247;
  assign sel_301094 = $signed({1'h0, add_300990}) < $signed({1'h0, sel_300992}) ? add_300990 : sel_300992;
  assign add_301097 = array_index_301029[11:0] + 12'h247;
  assign sel_301099 = $signed({1'h0, add_300995}) < $signed({1'h0, sel_300997}) ? add_300995 : sel_300997;
  assign array_index_301128 = set1_unflattened[8'hb7];
  assign array_index_301131 = set2_unflattened[8'hb7];
  assign add_301135 = array_index_300720[11:1] + 11'h79d;
  assign sel_301137 = $signed({1'h0, add_301033, array_index_300618[0]}) < $signed({1'h0, sel_301035}) ? {add_301033, array_index_300618[0]} : sel_301035;
  assign add_301139 = array_index_300723[11:1] + 11'h79d;
  assign sel_301141 = $signed({1'h0, add_301037, array_index_300621[0]}) < $signed({1'h0, sel_301039}) ? {add_301037, array_index_300621[0]} : sel_301039;
  assign add_301143 = array_index_300822[11:1] + 11'h347;
  assign sel_301145 = $signed({1'h0, add_301041, array_index_300720[0]}) < $signed({1'h0, sel_301043}) ? {add_301041, array_index_300720[0]} : sel_301043;
  assign add_301147 = array_index_300825[11:1] + 11'h347;
  assign sel_301149 = $signed({1'h0, add_301045, array_index_300723[0]}) < $signed({1'h0, sel_301047}) ? {add_301045, array_index_300723[0]} : sel_301047;
  assign add_301151 = array_index_300924[11:3] + 9'h0bd;
  assign sel_301154 = $signed({1'h0, add_301049, array_index_300822[2:0]}) < $signed({1'h0, sel_301052}) ? {add_301049, array_index_300822[2:0]} : sel_301052;
  assign add_301156 = array_index_300927[11:3] + 9'h0bd;
  assign sel_301159 = $signed({1'h0, add_301054, array_index_300825[2:0]}) < $signed({1'h0, sel_301057}) ? {add_301054, array_index_300825[2:0]} : sel_301057;
  assign add_301161 = array_index_301026[11:1] + 11'h247;
  assign sel_301164 = $signed({1'h0, add_301059, array_index_300924[0]}) < $signed({1'h0, sel_301062}) ? {add_301059, array_index_300924[0]} : sel_301062;
  assign add_301166 = array_index_301029[11:1] + 11'h247;
  assign sel_301169 = $signed({1'h0, add_301064, array_index_300927[0]}) < $signed({1'h0, sel_301067}) ? {add_301064, array_index_300927[0]} : sel_301067;
  assign add_301194 = array_index_301128[11:0] + 12'h247;
  assign sel_301196 = $signed({1'h0, add_301092}) < $signed({1'h0, sel_301094}) ? add_301092 : sel_301094;
  assign add_301199 = array_index_301131[11:0] + 12'h247;
  assign sel_301201 = $signed({1'h0, add_301097}) < $signed({1'h0, sel_301099}) ? add_301097 : sel_301099;
  assign array_index_301230 = set1_unflattened[8'hb8];
  assign array_index_301233 = set2_unflattened[8'hb8];
  assign add_301237 = array_index_300822[11:1] + 11'h79d;
  assign sel_301239 = $signed({1'h0, add_301135, array_index_300720[0]}) < $signed({1'h0, sel_301137}) ? {add_301135, array_index_300720[0]} : sel_301137;
  assign add_301241 = array_index_300825[11:1] + 11'h79d;
  assign sel_301243 = $signed({1'h0, add_301139, array_index_300723[0]}) < $signed({1'h0, sel_301141}) ? {add_301139, array_index_300723[0]} : sel_301141;
  assign add_301245 = array_index_300924[11:1] + 11'h347;
  assign sel_301247 = $signed({1'h0, add_301143, array_index_300822[0]}) < $signed({1'h0, sel_301145}) ? {add_301143, array_index_300822[0]} : sel_301145;
  assign add_301249 = array_index_300927[11:1] + 11'h347;
  assign sel_301251 = $signed({1'h0, add_301147, array_index_300825[0]}) < $signed({1'h0, sel_301149}) ? {add_301147, array_index_300825[0]} : sel_301149;
  assign add_301253 = array_index_301026[11:3] + 9'h0bd;
  assign sel_301256 = $signed({1'h0, add_301151, array_index_300924[2:0]}) < $signed({1'h0, sel_301154}) ? {add_301151, array_index_300924[2:0]} : sel_301154;
  assign add_301258 = array_index_301029[11:3] + 9'h0bd;
  assign sel_301261 = $signed({1'h0, add_301156, array_index_300927[2:0]}) < $signed({1'h0, sel_301159}) ? {add_301156, array_index_300927[2:0]} : sel_301159;
  assign add_301263 = array_index_301128[11:1] + 11'h247;
  assign sel_301266 = $signed({1'h0, add_301161, array_index_301026[0]}) < $signed({1'h0, sel_301164}) ? {add_301161, array_index_301026[0]} : sel_301164;
  assign add_301268 = array_index_301131[11:1] + 11'h247;
  assign sel_301271 = $signed({1'h0, add_301166, array_index_301029[0]}) < $signed({1'h0, sel_301169}) ? {add_301166, array_index_301029[0]} : sel_301169;
  assign add_301296 = array_index_301230[11:0] + 12'h247;
  assign sel_301298 = $signed({1'h0, add_301194}) < $signed({1'h0, sel_301196}) ? add_301194 : sel_301196;
  assign add_301301 = array_index_301233[11:0] + 12'h247;
  assign sel_301303 = $signed({1'h0, add_301199}) < $signed({1'h0, sel_301201}) ? add_301199 : sel_301201;
  assign array_index_301332 = set1_unflattened[8'hb9];
  assign array_index_301335 = set2_unflattened[8'hb9];
  assign add_301339 = array_index_300924[11:1] + 11'h79d;
  assign sel_301341 = $signed({1'h0, add_301237, array_index_300822[0]}) < $signed({1'h0, sel_301239}) ? {add_301237, array_index_300822[0]} : sel_301239;
  assign add_301343 = array_index_300927[11:1] + 11'h79d;
  assign sel_301345 = $signed({1'h0, add_301241, array_index_300825[0]}) < $signed({1'h0, sel_301243}) ? {add_301241, array_index_300825[0]} : sel_301243;
  assign add_301347 = array_index_301026[11:1] + 11'h347;
  assign sel_301349 = $signed({1'h0, add_301245, array_index_300924[0]}) < $signed({1'h0, sel_301247}) ? {add_301245, array_index_300924[0]} : sel_301247;
  assign add_301351 = array_index_301029[11:1] + 11'h347;
  assign sel_301353 = $signed({1'h0, add_301249, array_index_300927[0]}) < $signed({1'h0, sel_301251}) ? {add_301249, array_index_300927[0]} : sel_301251;
  assign add_301355 = array_index_301128[11:3] + 9'h0bd;
  assign sel_301358 = $signed({1'h0, add_301253, array_index_301026[2:0]}) < $signed({1'h0, sel_301256}) ? {add_301253, array_index_301026[2:0]} : sel_301256;
  assign add_301360 = array_index_301131[11:3] + 9'h0bd;
  assign sel_301363 = $signed({1'h0, add_301258, array_index_301029[2:0]}) < $signed({1'h0, sel_301261}) ? {add_301258, array_index_301029[2:0]} : sel_301261;
  assign add_301365 = array_index_301230[11:1] + 11'h247;
  assign sel_301368 = $signed({1'h0, add_301263, array_index_301128[0]}) < $signed({1'h0, sel_301266}) ? {add_301263, array_index_301128[0]} : sel_301266;
  assign add_301370 = array_index_301233[11:1] + 11'h247;
  assign sel_301373 = $signed({1'h0, add_301268, array_index_301131[0]}) < $signed({1'h0, sel_301271}) ? {add_301268, array_index_301131[0]} : sel_301271;
  assign add_301398 = array_index_301332[11:0] + 12'h247;
  assign sel_301400 = $signed({1'h0, add_301296}) < $signed({1'h0, sel_301298}) ? add_301296 : sel_301298;
  assign add_301403 = array_index_301335[11:0] + 12'h247;
  assign sel_301405 = $signed({1'h0, add_301301}) < $signed({1'h0, sel_301303}) ? add_301301 : sel_301303;
  assign array_index_301434 = set1_unflattened[8'hba];
  assign array_index_301437 = set2_unflattened[8'hba];
  assign add_301441 = array_index_301026[11:1] + 11'h79d;
  assign sel_301443 = $signed({1'h0, add_301339, array_index_300924[0]}) < $signed({1'h0, sel_301341}) ? {add_301339, array_index_300924[0]} : sel_301341;
  assign add_301445 = array_index_301029[11:1] + 11'h79d;
  assign sel_301447 = $signed({1'h0, add_301343, array_index_300927[0]}) < $signed({1'h0, sel_301345}) ? {add_301343, array_index_300927[0]} : sel_301345;
  assign add_301449 = array_index_301128[11:1] + 11'h347;
  assign sel_301451 = $signed({1'h0, add_301347, array_index_301026[0]}) < $signed({1'h0, sel_301349}) ? {add_301347, array_index_301026[0]} : sel_301349;
  assign add_301453 = array_index_301131[11:1] + 11'h347;
  assign sel_301455 = $signed({1'h0, add_301351, array_index_301029[0]}) < $signed({1'h0, sel_301353}) ? {add_301351, array_index_301029[0]} : sel_301353;
  assign add_301457 = array_index_301230[11:3] + 9'h0bd;
  assign sel_301460 = $signed({1'h0, add_301355, array_index_301128[2:0]}) < $signed({1'h0, sel_301358}) ? {add_301355, array_index_301128[2:0]} : sel_301358;
  assign add_301462 = array_index_301233[11:3] + 9'h0bd;
  assign sel_301465 = $signed({1'h0, add_301360, array_index_301131[2:0]}) < $signed({1'h0, sel_301363}) ? {add_301360, array_index_301131[2:0]} : sel_301363;
  assign add_301467 = array_index_301332[11:1] + 11'h247;
  assign sel_301470 = $signed({1'h0, add_301365, array_index_301230[0]}) < $signed({1'h0, sel_301368}) ? {add_301365, array_index_301230[0]} : sel_301368;
  assign add_301472 = array_index_301335[11:1] + 11'h247;
  assign sel_301475 = $signed({1'h0, add_301370, array_index_301233[0]}) < $signed({1'h0, sel_301373}) ? {add_301370, array_index_301233[0]} : sel_301373;
  assign add_301500 = array_index_301434[11:0] + 12'h247;
  assign sel_301502 = $signed({1'h0, add_301398}) < $signed({1'h0, sel_301400}) ? add_301398 : sel_301400;
  assign add_301505 = array_index_301437[11:0] + 12'h247;
  assign sel_301507 = $signed({1'h0, add_301403}) < $signed({1'h0, sel_301405}) ? add_301403 : sel_301405;
  assign array_index_301536 = set1_unflattened[8'hbb];
  assign array_index_301539 = set2_unflattened[8'hbb];
  assign add_301543 = array_index_301128[11:1] + 11'h79d;
  assign sel_301545 = $signed({1'h0, add_301441, array_index_301026[0]}) < $signed({1'h0, sel_301443}) ? {add_301441, array_index_301026[0]} : sel_301443;
  assign add_301547 = array_index_301131[11:1] + 11'h79d;
  assign sel_301549 = $signed({1'h0, add_301445, array_index_301029[0]}) < $signed({1'h0, sel_301447}) ? {add_301445, array_index_301029[0]} : sel_301447;
  assign add_301551 = array_index_301230[11:1] + 11'h347;
  assign sel_301553 = $signed({1'h0, add_301449, array_index_301128[0]}) < $signed({1'h0, sel_301451}) ? {add_301449, array_index_301128[0]} : sel_301451;
  assign add_301555 = array_index_301233[11:1] + 11'h347;
  assign sel_301557 = $signed({1'h0, add_301453, array_index_301131[0]}) < $signed({1'h0, sel_301455}) ? {add_301453, array_index_301131[0]} : sel_301455;
  assign add_301559 = array_index_301332[11:3] + 9'h0bd;
  assign sel_301562 = $signed({1'h0, add_301457, array_index_301230[2:0]}) < $signed({1'h0, sel_301460}) ? {add_301457, array_index_301230[2:0]} : sel_301460;
  assign add_301564 = array_index_301335[11:3] + 9'h0bd;
  assign sel_301567 = $signed({1'h0, add_301462, array_index_301233[2:0]}) < $signed({1'h0, sel_301465}) ? {add_301462, array_index_301233[2:0]} : sel_301465;
  assign add_301569 = array_index_301434[11:1] + 11'h247;
  assign sel_301572 = $signed({1'h0, add_301467, array_index_301332[0]}) < $signed({1'h0, sel_301470}) ? {add_301467, array_index_301332[0]} : sel_301470;
  assign add_301574 = array_index_301437[11:1] + 11'h247;
  assign sel_301577 = $signed({1'h0, add_301472, array_index_301335[0]}) < $signed({1'h0, sel_301475}) ? {add_301472, array_index_301335[0]} : sel_301475;
  assign add_301602 = array_index_301536[11:0] + 12'h247;
  assign sel_301604 = $signed({1'h0, add_301500}) < $signed({1'h0, sel_301502}) ? add_301500 : sel_301502;
  assign add_301607 = array_index_301539[11:0] + 12'h247;
  assign sel_301609 = $signed({1'h0, add_301505}) < $signed({1'h0, sel_301507}) ? add_301505 : sel_301507;
  assign array_index_301638 = set1_unflattened[8'hbc];
  assign array_index_301641 = set2_unflattened[8'hbc];
  assign add_301645 = array_index_301230[11:1] + 11'h79d;
  assign sel_301647 = $signed({1'h0, add_301543, array_index_301128[0]}) < $signed({1'h0, sel_301545}) ? {add_301543, array_index_301128[0]} : sel_301545;
  assign add_301649 = array_index_301233[11:1] + 11'h79d;
  assign sel_301651 = $signed({1'h0, add_301547, array_index_301131[0]}) < $signed({1'h0, sel_301549}) ? {add_301547, array_index_301131[0]} : sel_301549;
  assign add_301653 = array_index_301332[11:1] + 11'h347;
  assign sel_301655 = $signed({1'h0, add_301551, array_index_301230[0]}) < $signed({1'h0, sel_301553}) ? {add_301551, array_index_301230[0]} : sel_301553;
  assign add_301657 = array_index_301335[11:1] + 11'h347;
  assign sel_301659 = $signed({1'h0, add_301555, array_index_301233[0]}) < $signed({1'h0, sel_301557}) ? {add_301555, array_index_301233[0]} : sel_301557;
  assign add_301661 = array_index_301434[11:3] + 9'h0bd;
  assign sel_301664 = $signed({1'h0, add_301559, array_index_301332[2:0]}) < $signed({1'h0, sel_301562}) ? {add_301559, array_index_301332[2:0]} : sel_301562;
  assign add_301666 = array_index_301437[11:3] + 9'h0bd;
  assign sel_301669 = $signed({1'h0, add_301564, array_index_301335[2:0]}) < $signed({1'h0, sel_301567}) ? {add_301564, array_index_301335[2:0]} : sel_301567;
  assign add_301671 = array_index_301536[11:1] + 11'h247;
  assign sel_301674 = $signed({1'h0, add_301569, array_index_301434[0]}) < $signed({1'h0, sel_301572}) ? {add_301569, array_index_301434[0]} : sel_301572;
  assign add_301676 = array_index_301539[11:1] + 11'h247;
  assign sel_301679 = $signed({1'h0, add_301574, array_index_301437[0]}) < $signed({1'h0, sel_301577}) ? {add_301574, array_index_301437[0]} : sel_301577;
  assign add_301704 = array_index_301638[11:0] + 12'h247;
  assign sel_301706 = $signed({1'h0, add_301602}) < $signed({1'h0, sel_301604}) ? add_301602 : sel_301604;
  assign add_301709 = array_index_301641[11:0] + 12'h247;
  assign sel_301711 = $signed({1'h0, add_301607}) < $signed({1'h0, sel_301609}) ? add_301607 : sel_301609;
  assign array_index_301740 = set1_unflattened[8'hbd];
  assign array_index_301743 = set2_unflattened[8'hbd];
  assign add_301747 = array_index_301332[11:1] + 11'h79d;
  assign sel_301749 = $signed({1'h0, add_301645, array_index_301230[0]}) < $signed({1'h0, sel_301647}) ? {add_301645, array_index_301230[0]} : sel_301647;
  assign add_301751 = array_index_301335[11:1] + 11'h79d;
  assign sel_301753 = $signed({1'h0, add_301649, array_index_301233[0]}) < $signed({1'h0, sel_301651}) ? {add_301649, array_index_301233[0]} : sel_301651;
  assign add_301755 = array_index_301434[11:1] + 11'h347;
  assign sel_301757 = $signed({1'h0, add_301653, array_index_301332[0]}) < $signed({1'h0, sel_301655}) ? {add_301653, array_index_301332[0]} : sel_301655;
  assign add_301759 = array_index_301437[11:1] + 11'h347;
  assign sel_301761 = $signed({1'h0, add_301657, array_index_301335[0]}) < $signed({1'h0, sel_301659}) ? {add_301657, array_index_301335[0]} : sel_301659;
  assign add_301763 = array_index_301536[11:3] + 9'h0bd;
  assign sel_301766 = $signed({1'h0, add_301661, array_index_301434[2:0]}) < $signed({1'h0, sel_301664}) ? {add_301661, array_index_301434[2:0]} : sel_301664;
  assign add_301768 = array_index_301539[11:3] + 9'h0bd;
  assign sel_301771 = $signed({1'h0, add_301666, array_index_301437[2:0]}) < $signed({1'h0, sel_301669}) ? {add_301666, array_index_301437[2:0]} : sel_301669;
  assign add_301773 = array_index_301638[11:1] + 11'h247;
  assign sel_301776 = $signed({1'h0, add_301671, array_index_301536[0]}) < $signed({1'h0, sel_301674}) ? {add_301671, array_index_301536[0]} : sel_301674;
  assign add_301778 = array_index_301641[11:1] + 11'h247;
  assign sel_301781 = $signed({1'h0, add_301676, array_index_301539[0]}) < $signed({1'h0, sel_301679}) ? {add_301676, array_index_301539[0]} : sel_301679;
  assign add_301806 = array_index_301740[11:0] + 12'h247;
  assign sel_301808 = $signed({1'h0, add_301704}) < $signed({1'h0, sel_301706}) ? add_301704 : sel_301706;
  assign add_301811 = array_index_301743[11:0] + 12'h247;
  assign sel_301813 = $signed({1'h0, add_301709}) < $signed({1'h0, sel_301711}) ? add_301709 : sel_301711;
  assign array_index_301842 = set1_unflattened[8'hbe];
  assign array_index_301845 = set2_unflattened[8'hbe];
  assign add_301849 = array_index_301434[11:1] + 11'h79d;
  assign sel_301851 = $signed({1'h0, add_301747, array_index_301332[0]}) < $signed({1'h0, sel_301749}) ? {add_301747, array_index_301332[0]} : sel_301749;
  assign add_301853 = array_index_301437[11:1] + 11'h79d;
  assign sel_301855 = $signed({1'h0, add_301751, array_index_301335[0]}) < $signed({1'h0, sel_301753}) ? {add_301751, array_index_301335[0]} : sel_301753;
  assign add_301857 = array_index_301536[11:1] + 11'h347;
  assign sel_301859 = $signed({1'h0, add_301755, array_index_301434[0]}) < $signed({1'h0, sel_301757}) ? {add_301755, array_index_301434[0]} : sel_301757;
  assign add_301861 = array_index_301539[11:1] + 11'h347;
  assign sel_301863 = $signed({1'h0, add_301759, array_index_301437[0]}) < $signed({1'h0, sel_301761}) ? {add_301759, array_index_301437[0]} : sel_301761;
  assign add_301865 = array_index_301638[11:3] + 9'h0bd;
  assign sel_301868 = $signed({1'h0, add_301763, array_index_301536[2:0]}) < $signed({1'h0, sel_301766}) ? {add_301763, array_index_301536[2:0]} : sel_301766;
  assign add_301870 = array_index_301641[11:3] + 9'h0bd;
  assign sel_301873 = $signed({1'h0, add_301768, array_index_301539[2:0]}) < $signed({1'h0, sel_301771}) ? {add_301768, array_index_301539[2:0]} : sel_301771;
  assign add_301875 = array_index_301740[11:1] + 11'h247;
  assign sel_301878 = $signed({1'h0, add_301773, array_index_301638[0]}) < $signed({1'h0, sel_301776}) ? {add_301773, array_index_301638[0]} : sel_301776;
  assign add_301880 = array_index_301743[11:1] + 11'h247;
  assign sel_301883 = $signed({1'h0, add_301778, array_index_301641[0]}) < $signed({1'h0, sel_301781}) ? {add_301778, array_index_301641[0]} : sel_301781;
  assign add_301908 = array_index_301842[11:0] + 12'h247;
  assign sel_301910 = $signed({1'h0, add_301806}) < $signed({1'h0, sel_301808}) ? add_301806 : sel_301808;
  assign add_301913 = array_index_301845[11:0] + 12'h247;
  assign sel_301915 = $signed({1'h0, add_301811}) < $signed({1'h0, sel_301813}) ? add_301811 : sel_301813;
  assign array_index_301944 = set1_unflattened[8'hbf];
  assign array_index_301947 = set2_unflattened[8'hbf];
  assign add_301951 = array_index_301536[11:1] + 11'h79d;
  assign sel_301953 = $signed({1'h0, add_301849, array_index_301434[0]}) < $signed({1'h0, sel_301851}) ? {add_301849, array_index_301434[0]} : sel_301851;
  assign add_301955 = array_index_301539[11:1] + 11'h79d;
  assign sel_301957 = $signed({1'h0, add_301853, array_index_301437[0]}) < $signed({1'h0, sel_301855}) ? {add_301853, array_index_301437[0]} : sel_301855;
  assign add_301959 = array_index_301638[11:1] + 11'h347;
  assign sel_301961 = $signed({1'h0, add_301857, array_index_301536[0]}) < $signed({1'h0, sel_301859}) ? {add_301857, array_index_301536[0]} : sel_301859;
  assign add_301963 = array_index_301641[11:1] + 11'h347;
  assign sel_301965 = $signed({1'h0, add_301861, array_index_301539[0]}) < $signed({1'h0, sel_301863}) ? {add_301861, array_index_301539[0]} : sel_301863;
  assign add_301967 = array_index_301740[11:3] + 9'h0bd;
  assign sel_301970 = $signed({1'h0, add_301865, array_index_301638[2:0]}) < $signed({1'h0, sel_301868}) ? {add_301865, array_index_301638[2:0]} : sel_301868;
  assign add_301972 = array_index_301743[11:3] + 9'h0bd;
  assign sel_301975 = $signed({1'h0, add_301870, array_index_301641[2:0]}) < $signed({1'h0, sel_301873}) ? {add_301870, array_index_301641[2:0]} : sel_301873;
  assign add_301977 = array_index_301842[11:1] + 11'h247;
  assign sel_301980 = $signed({1'h0, add_301875, array_index_301740[0]}) < $signed({1'h0, sel_301878}) ? {add_301875, array_index_301740[0]} : sel_301878;
  assign add_301982 = array_index_301845[11:1] + 11'h247;
  assign sel_301985 = $signed({1'h0, add_301880, array_index_301743[0]}) < $signed({1'h0, sel_301883}) ? {add_301880, array_index_301743[0]} : sel_301883;
  assign add_302010 = array_index_301944[11:0] + 12'h247;
  assign sel_302012 = $signed({1'h0, add_301908}) < $signed({1'h0, sel_301910}) ? add_301908 : sel_301910;
  assign add_302015 = array_index_301947[11:0] + 12'h247;
  assign sel_302017 = $signed({1'h0, add_301913}) < $signed({1'h0, sel_301915}) ? add_301913 : sel_301915;
  assign array_index_302046 = set1_unflattened[8'hc0];
  assign array_index_302049 = set2_unflattened[8'hc0];
  assign add_302053 = array_index_301638[11:1] + 11'h79d;
  assign sel_302055 = $signed({1'h0, add_301951, array_index_301536[0]}) < $signed({1'h0, sel_301953}) ? {add_301951, array_index_301536[0]} : sel_301953;
  assign add_302057 = array_index_301641[11:1] + 11'h79d;
  assign sel_302059 = $signed({1'h0, add_301955, array_index_301539[0]}) < $signed({1'h0, sel_301957}) ? {add_301955, array_index_301539[0]} : sel_301957;
  assign add_302061 = array_index_301740[11:1] + 11'h347;
  assign sel_302063 = $signed({1'h0, add_301959, array_index_301638[0]}) < $signed({1'h0, sel_301961}) ? {add_301959, array_index_301638[0]} : sel_301961;
  assign add_302065 = array_index_301743[11:1] + 11'h347;
  assign sel_302067 = $signed({1'h0, add_301963, array_index_301641[0]}) < $signed({1'h0, sel_301965}) ? {add_301963, array_index_301641[0]} : sel_301965;
  assign add_302069 = array_index_301842[11:3] + 9'h0bd;
  assign sel_302072 = $signed({1'h0, add_301967, array_index_301740[2:0]}) < $signed({1'h0, sel_301970}) ? {add_301967, array_index_301740[2:0]} : sel_301970;
  assign add_302074 = array_index_301845[11:3] + 9'h0bd;
  assign sel_302077 = $signed({1'h0, add_301972, array_index_301743[2:0]}) < $signed({1'h0, sel_301975}) ? {add_301972, array_index_301743[2:0]} : sel_301975;
  assign add_302079 = array_index_301944[11:1] + 11'h247;
  assign sel_302082 = $signed({1'h0, add_301977, array_index_301842[0]}) < $signed({1'h0, sel_301980}) ? {add_301977, array_index_301842[0]} : sel_301980;
  assign add_302084 = array_index_301947[11:1] + 11'h247;
  assign sel_302087 = $signed({1'h0, add_301982, array_index_301845[0]}) < $signed({1'h0, sel_301985}) ? {add_301982, array_index_301845[0]} : sel_301985;
  assign add_302112 = array_index_302046[11:0] + 12'h247;
  assign sel_302114 = $signed({1'h0, add_302010}) < $signed({1'h0, sel_302012}) ? add_302010 : sel_302012;
  assign add_302117 = array_index_302049[11:0] + 12'h247;
  assign sel_302119 = $signed({1'h0, add_302015}) < $signed({1'h0, sel_302017}) ? add_302015 : sel_302017;
  assign array_index_302148 = set1_unflattened[8'hc1];
  assign array_index_302151 = set2_unflattened[8'hc1];
  assign add_302155 = array_index_301740[11:1] + 11'h79d;
  assign sel_302157 = $signed({1'h0, add_302053, array_index_301638[0]}) < $signed({1'h0, sel_302055}) ? {add_302053, array_index_301638[0]} : sel_302055;
  assign add_302159 = array_index_301743[11:1] + 11'h79d;
  assign sel_302161 = $signed({1'h0, add_302057, array_index_301641[0]}) < $signed({1'h0, sel_302059}) ? {add_302057, array_index_301641[0]} : sel_302059;
  assign add_302163 = array_index_301842[11:1] + 11'h347;
  assign sel_302165 = $signed({1'h0, add_302061, array_index_301740[0]}) < $signed({1'h0, sel_302063}) ? {add_302061, array_index_301740[0]} : sel_302063;
  assign add_302167 = array_index_301845[11:1] + 11'h347;
  assign sel_302169 = $signed({1'h0, add_302065, array_index_301743[0]}) < $signed({1'h0, sel_302067}) ? {add_302065, array_index_301743[0]} : sel_302067;
  assign add_302171 = array_index_301944[11:3] + 9'h0bd;
  assign sel_302174 = $signed({1'h0, add_302069, array_index_301842[2:0]}) < $signed({1'h0, sel_302072}) ? {add_302069, array_index_301842[2:0]} : sel_302072;
  assign add_302176 = array_index_301947[11:3] + 9'h0bd;
  assign sel_302179 = $signed({1'h0, add_302074, array_index_301845[2:0]}) < $signed({1'h0, sel_302077}) ? {add_302074, array_index_301845[2:0]} : sel_302077;
  assign add_302181 = array_index_302046[11:1] + 11'h247;
  assign sel_302184 = $signed({1'h0, add_302079, array_index_301944[0]}) < $signed({1'h0, sel_302082}) ? {add_302079, array_index_301944[0]} : sel_302082;
  assign add_302186 = array_index_302049[11:1] + 11'h247;
  assign sel_302189 = $signed({1'h0, add_302084, array_index_301947[0]}) < $signed({1'h0, sel_302087}) ? {add_302084, array_index_301947[0]} : sel_302087;
  assign add_302214 = array_index_302148[11:0] + 12'h247;
  assign sel_302216 = $signed({1'h0, add_302112}) < $signed({1'h0, sel_302114}) ? add_302112 : sel_302114;
  assign add_302219 = array_index_302151[11:0] + 12'h247;
  assign sel_302221 = $signed({1'h0, add_302117}) < $signed({1'h0, sel_302119}) ? add_302117 : sel_302119;
  assign array_index_302250 = set1_unflattened[8'hc2];
  assign array_index_302253 = set2_unflattened[8'hc2];
  assign add_302257 = array_index_301842[11:1] + 11'h79d;
  assign sel_302259 = $signed({1'h0, add_302155, array_index_301740[0]}) < $signed({1'h0, sel_302157}) ? {add_302155, array_index_301740[0]} : sel_302157;
  assign add_302261 = array_index_301845[11:1] + 11'h79d;
  assign sel_302263 = $signed({1'h0, add_302159, array_index_301743[0]}) < $signed({1'h0, sel_302161}) ? {add_302159, array_index_301743[0]} : sel_302161;
  assign add_302265 = array_index_301944[11:1] + 11'h347;
  assign sel_302267 = $signed({1'h0, add_302163, array_index_301842[0]}) < $signed({1'h0, sel_302165}) ? {add_302163, array_index_301842[0]} : sel_302165;
  assign add_302269 = array_index_301947[11:1] + 11'h347;
  assign sel_302271 = $signed({1'h0, add_302167, array_index_301845[0]}) < $signed({1'h0, sel_302169}) ? {add_302167, array_index_301845[0]} : sel_302169;
  assign add_302273 = array_index_302046[11:3] + 9'h0bd;
  assign sel_302276 = $signed({1'h0, add_302171, array_index_301944[2:0]}) < $signed({1'h0, sel_302174}) ? {add_302171, array_index_301944[2:0]} : sel_302174;
  assign add_302278 = array_index_302049[11:3] + 9'h0bd;
  assign sel_302281 = $signed({1'h0, add_302176, array_index_301947[2:0]}) < $signed({1'h0, sel_302179}) ? {add_302176, array_index_301947[2:0]} : sel_302179;
  assign add_302283 = array_index_302148[11:1] + 11'h247;
  assign sel_302286 = $signed({1'h0, add_302181, array_index_302046[0]}) < $signed({1'h0, sel_302184}) ? {add_302181, array_index_302046[0]} : sel_302184;
  assign add_302288 = array_index_302151[11:1] + 11'h247;
  assign sel_302291 = $signed({1'h0, add_302186, array_index_302049[0]}) < $signed({1'h0, sel_302189}) ? {add_302186, array_index_302049[0]} : sel_302189;
  assign add_302316 = array_index_302250[11:0] + 12'h247;
  assign sel_302318 = $signed({1'h0, add_302214}) < $signed({1'h0, sel_302216}) ? add_302214 : sel_302216;
  assign add_302321 = array_index_302253[11:0] + 12'h247;
  assign sel_302323 = $signed({1'h0, add_302219}) < $signed({1'h0, sel_302221}) ? add_302219 : sel_302221;
  assign array_index_302352 = set1_unflattened[8'hc3];
  assign array_index_302355 = set2_unflattened[8'hc3];
  assign add_302359 = array_index_301944[11:1] + 11'h79d;
  assign sel_302361 = $signed({1'h0, add_302257, array_index_301842[0]}) < $signed({1'h0, sel_302259}) ? {add_302257, array_index_301842[0]} : sel_302259;
  assign add_302363 = array_index_301947[11:1] + 11'h79d;
  assign sel_302365 = $signed({1'h0, add_302261, array_index_301845[0]}) < $signed({1'h0, sel_302263}) ? {add_302261, array_index_301845[0]} : sel_302263;
  assign add_302367 = array_index_302046[11:1] + 11'h347;
  assign sel_302369 = $signed({1'h0, add_302265, array_index_301944[0]}) < $signed({1'h0, sel_302267}) ? {add_302265, array_index_301944[0]} : sel_302267;
  assign add_302371 = array_index_302049[11:1] + 11'h347;
  assign sel_302373 = $signed({1'h0, add_302269, array_index_301947[0]}) < $signed({1'h0, sel_302271}) ? {add_302269, array_index_301947[0]} : sel_302271;
  assign add_302375 = array_index_302148[11:3] + 9'h0bd;
  assign sel_302378 = $signed({1'h0, add_302273, array_index_302046[2:0]}) < $signed({1'h0, sel_302276}) ? {add_302273, array_index_302046[2:0]} : sel_302276;
  assign add_302380 = array_index_302151[11:3] + 9'h0bd;
  assign sel_302383 = $signed({1'h0, add_302278, array_index_302049[2:0]}) < $signed({1'h0, sel_302281}) ? {add_302278, array_index_302049[2:0]} : sel_302281;
  assign add_302385 = array_index_302250[11:1] + 11'h247;
  assign sel_302388 = $signed({1'h0, add_302283, array_index_302148[0]}) < $signed({1'h0, sel_302286}) ? {add_302283, array_index_302148[0]} : sel_302286;
  assign add_302390 = array_index_302253[11:1] + 11'h247;
  assign sel_302393 = $signed({1'h0, add_302288, array_index_302151[0]}) < $signed({1'h0, sel_302291}) ? {add_302288, array_index_302151[0]} : sel_302291;
  assign add_302418 = array_index_302352[11:0] + 12'h247;
  assign sel_302420 = $signed({1'h0, add_302316}) < $signed({1'h0, sel_302318}) ? add_302316 : sel_302318;
  assign add_302423 = array_index_302355[11:0] + 12'h247;
  assign sel_302425 = $signed({1'h0, add_302321}) < $signed({1'h0, sel_302323}) ? add_302321 : sel_302323;
  assign array_index_302454 = set1_unflattened[8'hc4];
  assign array_index_302457 = set2_unflattened[8'hc4];
  assign add_302461 = array_index_302046[11:1] + 11'h79d;
  assign sel_302463 = $signed({1'h0, add_302359, array_index_301944[0]}) < $signed({1'h0, sel_302361}) ? {add_302359, array_index_301944[0]} : sel_302361;
  assign add_302465 = array_index_302049[11:1] + 11'h79d;
  assign sel_302467 = $signed({1'h0, add_302363, array_index_301947[0]}) < $signed({1'h0, sel_302365}) ? {add_302363, array_index_301947[0]} : sel_302365;
  assign add_302469 = array_index_302148[11:1] + 11'h347;
  assign sel_302471 = $signed({1'h0, add_302367, array_index_302046[0]}) < $signed({1'h0, sel_302369}) ? {add_302367, array_index_302046[0]} : sel_302369;
  assign add_302473 = array_index_302151[11:1] + 11'h347;
  assign sel_302475 = $signed({1'h0, add_302371, array_index_302049[0]}) < $signed({1'h0, sel_302373}) ? {add_302371, array_index_302049[0]} : sel_302373;
  assign add_302477 = array_index_302250[11:3] + 9'h0bd;
  assign sel_302480 = $signed({1'h0, add_302375, array_index_302148[2:0]}) < $signed({1'h0, sel_302378}) ? {add_302375, array_index_302148[2:0]} : sel_302378;
  assign add_302482 = array_index_302253[11:3] + 9'h0bd;
  assign sel_302485 = $signed({1'h0, add_302380, array_index_302151[2:0]}) < $signed({1'h0, sel_302383}) ? {add_302380, array_index_302151[2:0]} : sel_302383;
  assign add_302487 = array_index_302352[11:1] + 11'h247;
  assign sel_302490 = $signed({1'h0, add_302385, array_index_302250[0]}) < $signed({1'h0, sel_302388}) ? {add_302385, array_index_302250[0]} : sel_302388;
  assign add_302492 = array_index_302355[11:1] + 11'h247;
  assign sel_302495 = $signed({1'h0, add_302390, array_index_302253[0]}) < $signed({1'h0, sel_302393}) ? {add_302390, array_index_302253[0]} : sel_302393;
  assign add_302520 = array_index_302454[11:0] + 12'h247;
  assign sel_302522 = $signed({1'h0, add_302418}) < $signed({1'h0, sel_302420}) ? add_302418 : sel_302420;
  assign add_302525 = array_index_302457[11:0] + 12'h247;
  assign sel_302527 = $signed({1'h0, add_302423}) < $signed({1'h0, sel_302425}) ? add_302423 : sel_302425;
  assign array_index_302556 = set1_unflattened[8'hc5];
  assign array_index_302559 = set2_unflattened[8'hc5];
  assign add_302563 = array_index_302148[11:1] + 11'h79d;
  assign sel_302565 = $signed({1'h0, add_302461, array_index_302046[0]}) < $signed({1'h0, sel_302463}) ? {add_302461, array_index_302046[0]} : sel_302463;
  assign add_302567 = array_index_302151[11:1] + 11'h79d;
  assign sel_302569 = $signed({1'h0, add_302465, array_index_302049[0]}) < $signed({1'h0, sel_302467}) ? {add_302465, array_index_302049[0]} : sel_302467;
  assign add_302571 = array_index_302250[11:1] + 11'h347;
  assign sel_302573 = $signed({1'h0, add_302469, array_index_302148[0]}) < $signed({1'h0, sel_302471}) ? {add_302469, array_index_302148[0]} : sel_302471;
  assign add_302575 = array_index_302253[11:1] + 11'h347;
  assign sel_302577 = $signed({1'h0, add_302473, array_index_302151[0]}) < $signed({1'h0, sel_302475}) ? {add_302473, array_index_302151[0]} : sel_302475;
  assign add_302579 = array_index_302352[11:3] + 9'h0bd;
  assign sel_302582 = $signed({1'h0, add_302477, array_index_302250[2:0]}) < $signed({1'h0, sel_302480}) ? {add_302477, array_index_302250[2:0]} : sel_302480;
  assign add_302584 = array_index_302355[11:3] + 9'h0bd;
  assign sel_302587 = $signed({1'h0, add_302482, array_index_302253[2:0]}) < $signed({1'h0, sel_302485}) ? {add_302482, array_index_302253[2:0]} : sel_302485;
  assign add_302589 = array_index_302454[11:1] + 11'h247;
  assign sel_302592 = $signed({1'h0, add_302487, array_index_302352[0]}) < $signed({1'h0, sel_302490}) ? {add_302487, array_index_302352[0]} : sel_302490;
  assign add_302594 = array_index_302457[11:1] + 11'h247;
  assign sel_302597 = $signed({1'h0, add_302492, array_index_302355[0]}) < $signed({1'h0, sel_302495}) ? {add_302492, array_index_302355[0]} : sel_302495;
  assign add_302622 = array_index_302556[11:0] + 12'h247;
  assign sel_302624 = $signed({1'h0, add_302520}) < $signed({1'h0, sel_302522}) ? add_302520 : sel_302522;
  assign add_302627 = array_index_302559[11:0] + 12'h247;
  assign sel_302629 = $signed({1'h0, add_302525}) < $signed({1'h0, sel_302527}) ? add_302525 : sel_302527;
  assign array_index_302658 = set1_unflattened[8'hc6];
  assign array_index_302661 = set2_unflattened[8'hc6];
  assign add_302665 = array_index_302250[11:1] + 11'h79d;
  assign sel_302667 = $signed({1'h0, add_302563, array_index_302148[0]}) < $signed({1'h0, sel_302565}) ? {add_302563, array_index_302148[0]} : sel_302565;
  assign add_302669 = array_index_302253[11:1] + 11'h79d;
  assign sel_302671 = $signed({1'h0, add_302567, array_index_302151[0]}) < $signed({1'h0, sel_302569}) ? {add_302567, array_index_302151[0]} : sel_302569;
  assign add_302673 = array_index_302352[11:1] + 11'h347;
  assign sel_302675 = $signed({1'h0, add_302571, array_index_302250[0]}) < $signed({1'h0, sel_302573}) ? {add_302571, array_index_302250[0]} : sel_302573;
  assign add_302677 = array_index_302355[11:1] + 11'h347;
  assign sel_302679 = $signed({1'h0, add_302575, array_index_302253[0]}) < $signed({1'h0, sel_302577}) ? {add_302575, array_index_302253[0]} : sel_302577;
  assign add_302681 = array_index_302454[11:3] + 9'h0bd;
  assign sel_302684 = $signed({1'h0, add_302579, array_index_302352[2:0]}) < $signed({1'h0, sel_302582}) ? {add_302579, array_index_302352[2:0]} : sel_302582;
  assign add_302686 = array_index_302457[11:3] + 9'h0bd;
  assign sel_302689 = $signed({1'h0, add_302584, array_index_302355[2:0]}) < $signed({1'h0, sel_302587}) ? {add_302584, array_index_302355[2:0]} : sel_302587;
  assign add_302691 = array_index_302556[11:1] + 11'h247;
  assign sel_302694 = $signed({1'h0, add_302589, array_index_302454[0]}) < $signed({1'h0, sel_302592}) ? {add_302589, array_index_302454[0]} : sel_302592;
  assign add_302696 = array_index_302559[11:1] + 11'h247;
  assign sel_302699 = $signed({1'h0, add_302594, array_index_302457[0]}) < $signed({1'h0, sel_302597}) ? {add_302594, array_index_302457[0]} : sel_302597;
  assign add_302724 = array_index_302658[11:0] + 12'h247;
  assign sel_302726 = $signed({1'h0, add_302622}) < $signed({1'h0, sel_302624}) ? add_302622 : sel_302624;
  assign add_302729 = array_index_302661[11:0] + 12'h247;
  assign sel_302731 = $signed({1'h0, add_302627}) < $signed({1'h0, sel_302629}) ? add_302627 : sel_302629;
  assign array_index_302760 = set1_unflattened[8'h63];
  assign array_index_302763 = set2_unflattened[8'hc7];
  assign add_302767 = array_index_302352[11:1] + 11'h79d;
  assign sel_302769 = $signed({1'h0, add_302665, array_index_302250[0]}) < $signed({1'h0, sel_302667}) ? {add_302665, array_index_302250[0]} : sel_302667;
  assign add_302771 = array_index_302355[11:1] + 11'h79d;
  assign sel_302773 = $signed({1'h0, add_302669, array_index_302253[0]}) < $signed({1'h0, sel_302671}) ? {add_302669, array_index_302253[0]} : sel_302671;
  assign add_302775 = array_index_302454[11:1] + 11'h347;
  assign sel_302777 = $signed({1'h0, add_302673, array_index_302352[0]}) < $signed({1'h0, sel_302675}) ? {add_302673, array_index_302352[0]} : sel_302675;
  assign add_302779 = array_index_302457[11:1] + 11'h347;
  assign sel_302781 = $signed({1'h0, add_302677, array_index_302355[0]}) < $signed({1'h0, sel_302679}) ? {add_302677, array_index_302355[0]} : sel_302679;
  assign add_302783 = array_index_302556[11:3] + 9'h0bd;
  assign sel_302786 = $signed({1'h0, add_302681, array_index_302454[2:0]}) < $signed({1'h0, sel_302684}) ? {add_302681, array_index_302454[2:0]} : sel_302684;
  assign add_302788 = array_index_302559[11:3] + 9'h0bd;
  assign sel_302791 = $signed({1'h0, add_302686, array_index_302457[2:0]}) < $signed({1'h0, sel_302689}) ? {add_302686, array_index_302457[2:0]} : sel_302689;
  assign add_302793 = array_index_302658[11:1] + 11'h247;
  assign sel_302796 = $signed({1'h0, add_302691, array_index_302556[0]}) < $signed({1'h0, sel_302694}) ? {add_302691, array_index_302556[0]} : sel_302694;
  assign add_302798 = array_index_302661[11:1] + 11'h247;
  assign sel_302801 = $signed({1'h0, add_302696, array_index_302559[0]}) < $signed({1'h0, sel_302699}) ? {add_302696, array_index_302559[0]} : sel_302699;
  assign add_302825 = array_index_302760[11:0] + 12'h247;
  assign sel_302827 = $signed({1'h0, add_302724}) < $signed({1'h0, sel_302726}) ? add_302724 : sel_302726;
  assign add_302829 = array_index_302763[11:0] + 12'h247;
  assign sel_302831 = $signed({1'h0, add_302729}) < $signed({1'h0, sel_302731}) ? add_302729 : sel_302731;
  assign add_302865 = array_index_302454[11:1] + 11'h79d;
  assign sel_302867 = $signed({1'h0, add_302767, array_index_302352[0]}) < $signed({1'h0, sel_302769}) ? {add_302767, array_index_302352[0]} : sel_302769;
  assign add_302869 = array_index_302457[11:1] + 11'h79d;
  assign sel_302871 = $signed({1'h0, add_302771, array_index_302355[0]}) < $signed({1'h0, sel_302773}) ? {add_302771, array_index_302355[0]} : sel_302773;
  assign add_302873 = array_index_302556[11:1] + 11'h347;
  assign sel_302875 = $signed({1'h0, add_302775, array_index_302454[0]}) < $signed({1'h0, sel_302777}) ? {add_302775, array_index_302454[0]} : sel_302777;
  assign add_302877 = array_index_302559[11:1] + 11'h347;
  assign sel_302879 = $signed({1'h0, add_302779, array_index_302457[0]}) < $signed({1'h0, sel_302781}) ? {add_302779, array_index_302457[0]} : sel_302781;
  assign add_302881 = array_index_302658[11:3] + 9'h0bd;
  assign sel_302884 = $signed({1'h0, add_302783, array_index_302556[2:0]}) < $signed({1'h0, sel_302786}) ? {add_302783, array_index_302556[2:0]} : sel_302786;
  assign add_302886 = array_index_302661[11:3] + 9'h0bd;
  assign sel_302889 = $signed({1'h0, add_302788, array_index_302559[2:0]}) < $signed({1'h0, sel_302791}) ? {add_302788, array_index_302559[2:0]} : sel_302791;
  assign add_302891 = array_index_302760[11:1] + 11'h247;
  assign sel_302894 = $signed({1'h0, add_302793, array_index_302658[0]}) < $signed({1'h0, sel_302796}) ? {add_302793, array_index_302658[0]} : sel_302796;
  assign add_302896 = array_index_302763[11:1] + 11'h247;
  assign sel_302899 = $signed({1'h0, add_302798, array_index_302661[0]}) < $signed({1'h0, sel_302801}) ? {add_302798, array_index_302661[0]} : sel_302801;
  assign add_302947 = array_index_302556[11:1] + 11'h79d;
  assign sel_302949 = $signed({1'h0, add_302865, array_index_302454[0]}) < $signed({1'h0, sel_302867}) ? {add_302865, array_index_302454[0]} : sel_302867;
  assign add_302951 = array_index_302559[11:1] + 11'h79d;
  assign sel_302953 = $signed({1'h0, add_302869, array_index_302457[0]}) < $signed({1'h0, sel_302871}) ? {add_302869, array_index_302457[0]} : sel_302871;
  assign add_302955 = array_index_302658[11:1] + 11'h347;
  assign sel_302957 = $signed({1'h0, add_302873, array_index_302556[0]}) < $signed({1'h0, sel_302875}) ? {add_302873, array_index_302556[0]} : sel_302875;
  assign add_302959 = array_index_302661[11:1] + 11'h347;
  assign sel_302961 = $signed({1'h0, add_302877, array_index_302559[0]}) < $signed({1'h0, sel_302879}) ? {add_302877, array_index_302559[0]} : sel_302879;
  assign add_302963 = array_index_302760[11:3] + 9'h0bd;
  assign sel_302966 = $signed({1'h0, add_302881, array_index_302658[2:0]}) < $signed({1'h0, sel_302884}) ? {add_302881, array_index_302658[2:0]} : sel_302884;
  assign add_302968 = array_index_302763[11:3] + 9'h0bd;
  assign sel_302971 = $signed({1'h0, add_302886, array_index_302661[2:0]}) < $signed({1'h0, sel_302889}) ? {add_302886, array_index_302661[2:0]} : sel_302889;
  assign concat_302974 = {1'h0, ($signed({1'h0, add_302825}) < $signed({1'h0, sel_302827}) ? add_302825 : sel_302827) == ($signed({1'h0, add_302829}) < $signed({1'h0, sel_302831}) ? add_302829 : sel_302831)};
  assign add_302989 = concat_302974 + 2'h1;
  assign add_303009 = array_index_302658[11:1] + 11'h79d;
  assign sel_303011 = $signed({1'h0, add_302947, array_index_302556[0]}) < $signed({1'h0, sel_302949}) ? {add_302947, array_index_302556[0]} : sel_302949;
  assign add_303013 = array_index_302661[11:1] + 11'h79d;
  assign sel_303015 = $signed({1'h0, add_302951, array_index_302559[0]}) < $signed({1'h0, sel_302953}) ? {add_302951, array_index_302559[0]} : sel_302953;
  assign add_303017 = array_index_302760[11:1] + 11'h347;
  assign sel_303019 = $signed({1'h0, add_302955, array_index_302658[0]}) < $signed({1'h0, sel_302957}) ? {add_302955, array_index_302658[0]} : sel_302957;
  assign add_303021 = array_index_302763[11:1] + 11'h347;
  assign sel_303023 = $signed({1'h0, add_302959, array_index_302661[0]}) < $signed({1'h0, sel_302961}) ? {add_302959, array_index_302661[0]} : sel_302961;
  assign concat_303026 = {1'h0, ($signed({1'h0, add_302891, array_index_302760[0]}) < $signed({1'h0, sel_302894}) ? {add_302891, array_index_302760[0]} : sel_302894) == ($signed({1'h0, add_302896, array_index_302763[0]}) < $signed({1'h0, sel_302899}) ? {add_302896, array_index_302763[0]} : sel_302899) ? add_302989 : concat_302974};
  assign add_303037 = concat_303026 + 3'h1;
  assign add_303051 = array_index_302760[11:1] + 11'h79d;
  assign sel_303053 = $signed({1'h0, add_303009, array_index_302658[0]}) < $signed({1'h0, sel_303011}) ? {add_303009, array_index_302658[0]} : sel_303011;
  assign add_303055 = array_index_302763[11:1] + 11'h79d;
  assign sel_303057 = $signed({1'h0, add_303013, array_index_302661[0]}) < $signed({1'h0, sel_303015}) ? {add_303013, array_index_302661[0]} : sel_303015;
  assign concat_303060 = {1'h0, ($signed({1'h0, add_302963, array_index_302760[2:0]}) < $signed({1'h0, sel_302966}) ? {add_302963, array_index_302760[2:0]} : sel_302966) == ($signed({1'h0, add_302968, array_index_302763[2:0]}) < $signed({1'h0, sel_302971}) ? {add_302968, array_index_302763[2:0]} : sel_302971) ? add_303037 : concat_303026};
  assign add_303067 = concat_303060 + 4'h1;
  assign concat_303076 = {1'h0, ($signed({1'h0, add_303017, array_index_302760[0]}) < $signed({1'h0, sel_303019}) ? {add_303017, array_index_302760[0]} : sel_303019) == ($signed({1'h0, add_303021, array_index_302763[0]}) < $signed({1'h0, sel_303023}) ? {add_303021, array_index_302763[0]} : sel_303023) ? add_303067 : concat_303060};
  assign add_303079 = concat_303076 + 5'h01;
  assign out = {{11'h000, ($signed({1'h0, add_303051, array_index_302760[0]}) < $signed({1'h0, sel_303053}) ? {add_303051, array_index_302760[0]} : sel_303053) == ($signed({1'h0, add_303055, array_index_302763[0]}) < $signed({1'h0, sel_303057}) ? {add_303055, array_index_302763[0]} : sel_303057) ? add_303079 : concat_303076}, {set1_unflattened[199], set1_unflattened[198], set1_unflattened[197], set1_unflattened[196], set1_unflattened[195], set1_unflattened[194], set1_unflattened[193], set1_unflattened[192], set1_unflattened[191], set1_unflattened[190], set1_unflattened[189], set1_unflattened[188], set1_unflattened[187], set1_unflattened[186], set1_unflattened[185], set1_unflattened[184], set1_unflattened[183], set1_unflattened[182], set1_unflattened[181], set1_unflattened[180], set1_unflattened[179], set1_unflattened[178], set1_unflattened[177], set1_unflattened[176], set1_unflattened[175], set1_unflattened[174], set1_unflattened[173], set1_unflattened[172], set1_unflattened[171], set1_unflattened[170], set1_unflattened[169], set1_unflattened[168], set1_unflattened[167], set1_unflattened[166], set1_unflattened[165], set1_unflattened[164], set1_unflattened[163], set1_unflattened[162], set1_unflattened[161], set1_unflattened[160], set1_unflattened[159], set1_unflattened[158], set1_unflattened[157], set1_unflattened[156], set1_unflattened[155], set1_unflattened[154], set1_unflattened[153], set1_unflattened[152], set1_unflattened[151], set1_unflattened[150], set1_unflattened[149], set1_unflattened[148], set1_unflattened[147], set1_unflattened[146], set1_unflattened[145], set1_unflattened[144], set1_unflattened[143], set1_unflattened[142], set1_unflattened[141], set1_unflattened[140], set1_unflattened[139], set1_unflattened[138], set1_unflattened[137], set1_unflattened[136], set1_unflattened[135], set1_unflattened[134], set1_unflattened[133], set1_unflattened[132], set1_unflattened[131], set1_unflattened[130], set1_unflattened[129], set1_unflattened[128], set1_unflattened[127], set1_unflattened[126], set1_unflattened[125], set1_unflattened[124], set1_unflattened[123], set1_unflattened[122], set1_unflattened[121], set1_unflattened[120], set1_unflattened[119], set1_unflattened[118], set1_unflattened[117], set1_unflattened[116], set1_unflattened[115], set1_unflattened[114], set1_unflattened[113], set1_unflattened[112], set1_unflattened[111], set1_unflattened[110], set1_unflattened[109], set1_unflattened[108], set1_unflattened[107], set1_unflattened[106], set1_unflattened[105], set1_unflattened[104], set1_unflattened[103], set1_unflattened[102], set1_unflattened[101], set1_unflattened[100], set1_unflattened[99], set1_unflattened[98], set1_unflattened[97], set1_unflattened[96], set1_unflattened[95], set1_unflattened[94], set1_unflattened[93], set1_unflattened[92], set1_unflattened[91], set1_unflattened[90], set1_unflattened[89], set1_unflattened[88], set1_unflattened[87], set1_unflattened[86], set1_unflattened[85], set1_unflattened[84], set1_unflattened[83], set1_unflattened[82], set1_unflattened[81], set1_unflattened[80], set1_unflattened[79], set1_unflattened[78], set1_unflattened[77], set1_unflattened[76], set1_unflattened[75], set1_unflattened[74], set1_unflattened[73], set1_unflattened[72], set1_unflattened[71], set1_unflattened[70], set1_unflattened[69], set1_unflattened[68], set1_unflattened[67], set1_unflattened[66], set1_unflattened[65], set1_unflattened[64], set1_unflattened[63], set1_unflattened[62], set1_unflattened[61], set1_unflattened[60], set1_unflattened[59], set1_unflattened[58], set1_unflattened[57], set1_unflattened[56], set1_unflattened[55], set1_unflattened[54], set1_unflattened[53], set1_unflattened[52], set1_unflattened[51], set1_unflattened[50], set1_unflattened[49], set1_unflattened[48], set1_unflattened[47], set1_unflattened[46], set1_unflattened[45], set1_unflattened[44], set1_unflattened[43], set1_unflattened[42], set1_unflattened[41], set1_unflattened[40], set1_unflattened[39], set1_unflattened[38], set1_unflattened[37], set1_unflattened[36], set1_unflattened[35], set1_unflattened[34], set1_unflattened[33], set1_unflattened[32], set1_unflattened[31], set1_unflattened[30], set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[199], set2_unflattened[198], set2_unflattened[197], set2_unflattened[196], set2_unflattened[195], set2_unflattened[194], set2_unflattened[193], set2_unflattened[192], set2_unflattened[191], set2_unflattened[190], set2_unflattened[189], set2_unflattened[188], set2_unflattened[187], set2_unflattened[186], set2_unflattened[185], set2_unflattened[184], set2_unflattened[183], set2_unflattened[182], set2_unflattened[181], set2_unflattened[180], set2_unflattened[179], set2_unflattened[178], set2_unflattened[177], set2_unflattened[176], set2_unflattened[175], set2_unflattened[174], set2_unflattened[173], set2_unflattened[172], set2_unflattened[171], set2_unflattened[170], set2_unflattened[169], set2_unflattened[168], set2_unflattened[167], set2_unflattened[166], set2_unflattened[165], set2_unflattened[164], set2_unflattened[163], set2_unflattened[162], set2_unflattened[161], set2_unflattened[160], set2_unflattened[159], set2_unflattened[158], set2_unflattened[157], set2_unflattened[156], set2_unflattened[155], set2_unflattened[154], set2_unflattened[153], set2_unflattened[152], set2_unflattened[151], set2_unflattened[150], set2_unflattened[149], set2_unflattened[148], set2_unflattened[147], set2_unflattened[146], set2_unflattened[145], set2_unflattened[144], set2_unflattened[143], set2_unflattened[142], set2_unflattened[141], set2_unflattened[140], set2_unflattened[139], set2_unflattened[138], set2_unflattened[137], set2_unflattened[136], set2_unflattened[135], set2_unflattened[134], set2_unflattened[133], set2_unflattened[132], set2_unflattened[131], set2_unflattened[130], set2_unflattened[129], set2_unflattened[128], set2_unflattened[127], set2_unflattened[126], set2_unflattened[125], set2_unflattened[124], set2_unflattened[123], set2_unflattened[122], set2_unflattened[121], set2_unflattened[120], set2_unflattened[119], set2_unflattened[118], set2_unflattened[117], set2_unflattened[116], set2_unflattened[115], set2_unflattened[114], set2_unflattened[113], set2_unflattened[112], set2_unflattened[111], set2_unflattened[110], set2_unflattened[109], set2_unflattened[108], set2_unflattened[107], set2_unflattened[106], set2_unflattened[105], set2_unflattened[104], set2_unflattened[103], set2_unflattened[102], set2_unflattened[101], set2_unflattened[100], set2_unflattened[99], set2_unflattened[98], set2_unflattened[97], set2_unflattened[96], set2_unflattened[95], set2_unflattened[94], set2_unflattened[93], set2_unflattened[92], set2_unflattened[91], set2_unflattened[90], set2_unflattened[89], set2_unflattened[88], set2_unflattened[87], set2_unflattened[86], set2_unflattened[85], set2_unflattened[84], set2_unflattened[83], set2_unflattened[82], set2_unflattened[81], set2_unflattened[80], set2_unflattened[79], set2_unflattened[78], set2_unflattened[77], set2_unflattened[76], set2_unflattened[75], set2_unflattened[74], set2_unflattened[73], set2_unflattened[72], set2_unflattened[71], set2_unflattened[70], set2_unflattened[69], set2_unflattened[68], set2_unflattened[67], set2_unflattened[66], set2_unflattened[65], set2_unflattened[64], set2_unflattened[63], set2_unflattened[62], set2_unflattened[61], set2_unflattened[60], set2_unflattened[59], set2_unflattened[58], set2_unflattened[57], set2_unflattened[56], set2_unflattened[55], set2_unflattened[54], set2_unflattened[53], set2_unflattened[52], set2_unflattened[51], set2_unflattened[50], set2_unflattened[49], set2_unflattened[48], set2_unflattened[47], set2_unflattened[46], set2_unflattened[45], set2_unflattened[44], set2_unflattened[43], set2_unflattened[42], set2_unflattened[41], set2_unflattened[40], set2_unflattened[39], set2_unflattened[38], set2_unflattened[37], set2_unflattened[36], set2_unflattened[35], set2_unflattened[34], set2_unflattened[33], set2_unflattened[32], set2_unflattened[31], set2_unflattened[30], set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
