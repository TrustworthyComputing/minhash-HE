module min_hash(
  input wire [799:0] set1,
  input wire [799:0] set2,
  output wire [1615:0] out
);
  // lint_off MULTIPLY
  function automatic [21:0] umul22b_16b_x_6b (input reg [15:0] lhs, input reg [5:0] rhs);
    begin
      umul22b_16b_x_6b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  // lint_off MULTIPLY
  function automatic [22:0] umul23b_16b_x_7b (input reg [15:0] lhs, input reg [6:0] rhs);
    begin
      umul23b_16b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [15:0] set1_unflattened[50];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  assign set1_unflattened[30] = set1[495:480];
  assign set1_unflattened[31] = set1[511:496];
  assign set1_unflattened[32] = set1[527:512];
  assign set1_unflattened[33] = set1[543:528];
  assign set1_unflattened[34] = set1[559:544];
  assign set1_unflattened[35] = set1[575:560];
  assign set1_unflattened[36] = set1[591:576];
  assign set1_unflattened[37] = set1[607:592];
  assign set1_unflattened[38] = set1[623:608];
  assign set1_unflattened[39] = set1[639:624];
  assign set1_unflattened[40] = set1[655:640];
  assign set1_unflattened[41] = set1[671:656];
  assign set1_unflattened[42] = set1[687:672];
  assign set1_unflattened[43] = set1[703:688];
  assign set1_unflattened[44] = set1[719:704];
  assign set1_unflattened[45] = set1[735:720];
  assign set1_unflattened[46] = set1[751:736];
  assign set1_unflattened[47] = set1[767:752];
  assign set1_unflattened[48] = set1[783:768];
  assign set1_unflattened[49] = set1[799:784];
  wire [15:0] set2_unflattened[50];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  assign set2_unflattened[30] = set2[495:480];
  assign set2_unflattened[31] = set2[511:496];
  assign set2_unflattened[32] = set2[527:512];
  assign set2_unflattened[33] = set2[543:528];
  assign set2_unflattened[34] = set2[559:544];
  assign set2_unflattened[35] = set2[575:560];
  assign set2_unflattened[36] = set2[591:576];
  assign set2_unflattened[37] = set2[607:592];
  assign set2_unflattened[38] = set2[623:608];
  assign set2_unflattened[39] = set2[639:624];
  assign set2_unflattened[40] = set2[655:640];
  assign set2_unflattened[41] = set2[671:656];
  assign set2_unflattened[42] = set2[687:672];
  assign set2_unflattened[43] = set2[703:688];
  assign set2_unflattened[44] = set2[719:704];
  assign set2_unflattened[45] = set2[735:720];
  assign set2_unflattened[46] = set2[751:736];
  assign set2_unflattened[47] = set2[767:752];
  assign set2_unflattened[48] = set2[783:768];
  assign set2_unflattened[49] = set2[799:784];
  wire [15:0] array_index_86589;
  wire [15:0] array_index_86591;
  wire [21:0] umul_86593;
  wire [21:0] umul_86594;
  wire [21:0] umul_86603;
  wire [21:0] umul_86604;
  wire [15:0] array_index_86605;
  wire [15:0] array_index_86609;
  wire [21:0] umul_86617;
  wire [15:0] add_86619;
  wire [21:0] umul_86621;
  wire [15:0] add_86623;
  wire [21:0] umul_86643;
  wire [21:0] umul_86644;
  wire [21:0] umul_86645;
  wire [21:0] add_86647;
  wire [21:0] umul_86649;
  wire [21:0] add_86651;
  wire [15:0] array_index_86653;
  wire [31:0] smod_86657;
  wire [15:0] array_index_86658;
  wire [31:0] smod_86662;
  wire [21:0] umul_86675;
  wire [15:0] add_86677;
  wire [21:0] umul_86681;
  wire [15:0] add_86683;
  wire [31:0] smod_86698;
  wire [31:0] smod_86702;
  wire [22:0] umul_86717;
  wire [22:0] umul_86718;
  wire [21:0] umul_86719;
  wire [20:0] add_86721;
  wire [21:0] umul_86723;
  wire [20:0] add_86725;
  wire [21:0] umul_86727;
  wire [21:0] add_86729;
  wire [21:0] umul_86733;
  wire [21:0] add_86735;
  wire [15:0] array_index_86739;
  wire [31:0] smod_86743;
  wire [15:0] array_index_86746;
  wire [31:0] smod_86750;
  wire [21:0] umul_86777;
  wire [15:0] add_86779;
  wire [15:0] sel_86784;
  wire [21:0] umul_86785;
  wire [15:0] add_86787;
  wire [15:0] sel_86792;
  wire [31:0] smod_86804;
  wire [31:0] smod_86808;
  wire [31:0] smod_86812;
  wire [31:0] smod_86818;
  wire [22:0] umul_86835;
  wire [22:0] umul_86836;
  wire [22:0] umul_86837;
  wire [22:0] add_86839;
  wire [22:0] umul_86841;
  wire [22:0] add_86843;
  wire [21:0] umul_86845;
  wire [20:0] add_86847;
  wire [21:0] umul_86851;
  wire [20:0] add_86853;
  wire [21:0] umul_86857;
  wire [21:0] add_86859;
  wire [15:0] sel_86864;
  wire [21:0] umul_86865;
  wire [21:0] add_86867;
  wire [15:0] sel_86872;
  wire [15:0] array_index_86873;
  wire [31:0] smod_86877;
  wire [15:0] array_index_86879;
  wire [31:0] smod_86883;
  wire [21:0] umul_86921;
  wire [15:0] add_86923;
  wire [15:0] sel_86928;
  wire [21:0] umul_86929;
  wire [15:0] add_86931;
  wire [15:0] sel_86936;
  wire [31:0] smod_86946;
  wire [31:0] smod_86950;
  wire [31:0] smod_86954;
  wire [31:0] smod_86960;
  wire [31:0] smod_86966;
  wire [31:0] smod_86971;
  wire [22:0] umul_86987;
  wire [20:0] add_86989;
  wire [22:0] umul_86991;
  wire [20:0] add_86993;
  wire [22:0] umul_86995;
  wire [22:0] add_86997;
  wire [22:0] umul_87001;
  wire [22:0] add_87003;
  wire [21:0] umul_87007;
  wire [20:0] add_87009;
  wire [15:0] sel_87014;
  wire [21:0] umul_87015;
  wire [20:0] add_87017;
  wire [15:0] sel_87022;
  wire [21:0] umul_87023;
  wire [21:0] add_87025;
  wire [15:0] sel_87030;
  wire [21:0] umul_87031;
  wire [21:0] add_87033;
  wire [15:0] sel_87038;
  wire [15:0] array_index_87039;
  wire [31:0] smod_87043;
  wire [15:0] array_index_87045;
  wire [31:0] smod_87049;
  wire [21:0] umul_87095;
  wire [15:0] add_87097;
  wire [15:0] sel_87102;
  wire [21:0] umul_87103;
  wire [15:0] add_87105;
  wire [15:0] sel_87110;
  wire [31:0] smod_87114;
  wire [31:0] smod_87118;
  wire [31:0] smod_87122;
  wire [31:0] smod_87128;
  wire [31:0] smod_87134;
  wire [31:0] smod_87139;
  wire [31:0] smod_87144;
  wire [31:0] smod_87149;
  wire [22:0] umul_87165;
  wire [20:0] add_87167;
  wire [22:0] umul_87171;
  wire [20:0] add_87173;
  wire [22:0] umul_87177;
  wire [22:0] add_87179;
  wire [15:0] sel_87184;
  wire [22:0] umul_87185;
  wire [22:0] add_87187;
  wire [15:0] sel_87192;
  wire [21:0] umul_87193;
  wire [20:0] add_87195;
  wire [15:0] sel_87200;
  wire [21:0] umul_87201;
  wire [20:0] add_87203;
  wire [15:0] sel_87208;
  wire [21:0] umul_87209;
  wire [21:0] add_87211;
  wire [15:0] sel_87216;
  wire [21:0] umul_87217;
  wire [21:0] add_87219;
  wire [15:0] sel_87224;
  wire [15:0] array_index_87225;
  wire [31:0] smod_87229;
  wire [15:0] array_index_87231;
  wire [31:0] smod_87235;
  wire [21:0] umul_87285;
  wire [15:0] add_87287;
  wire [15:0] sel_87292;
  wire [21:0] umul_87293;
  wire [15:0] add_87295;
  wire [15:0] sel_87300;
  wire [31:0] smod_87304;
  wire [31:0] smod_87310;
  wire [31:0] smod_87316;
  wire [31:0] smod_87321;
  wire [31:0] smod_87326;
  wire [31:0] smod_87331;
  wire [31:0] smod_87336;
  wire [31:0] smod_87341;
  wire [22:0] umul_87357;
  wire [20:0] add_87359;
  wire [15:0] sel_87364;
  wire [22:0] umul_87365;
  wire [20:0] add_87367;
  wire [15:0] sel_87372;
  wire [22:0] umul_87373;
  wire [22:0] add_87375;
  wire [15:0] sel_87380;
  wire [22:0] umul_87381;
  wire [22:0] add_87383;
  wire [15:0] sel_87388;
  wire [21:0] umul_87389;
  wire [20:0] add_87391;
  wire [15:0] sel_87396;
  wire [21:0] umul_87397;
  wire [20:0] add_87399;
  wire [15:0] sel_87404;
  wire [21:0] umul_87405;
  wire [21:0] add_87407;
  wire [15:0] sel_87412;
  wire [21:0] umul_87413;
  wire [21:0] add_87415;
  wire [15:0] sel_87420;
  wire [15:0] array_index_87421;
  wire [31:0] smod_87425;
  wire [15:0] array_index_87427;
  wire [31:0] smod_87431;
  wire [21:0] umul_87481;
  wire [15:0] add_87483;
  wire [15:0] sel_87488;
  wire [21:0] umul_87489;
  wire [15:0] add_87491;
  wire [15:0] sel_87496;
  wire [31:0] smod_87500;
  wire [31:0] smod_87505;
  wire [31:0] smod_87510;
  wire [31:0] smod_87515;
  wire [31:0] smod_87520;
  wire [31:0] smod_87525;
  wire [31:0] smod_87530;
  wire [31:0] smod_87535;
  wire [22:0] umul_87551;
  wire [20:0] add_87553;
  wire [15:0] sel_87558;
  wire [22:0] umul_87559;
  wire [20:0] add_87561;
  wire [15:0] sel_87566;
  wire [22:0] umul_87567;
  wire [22:0] add_87569;
  wire [15:0] sel_87574;
  wire [22:0] umul_87575;
  wire [22:0] add_87577;
  wire [15:0] sel_87582;
  wire [21:0] umul_87583;
  wire [20:0] add_87585;
  wire [15:0] sel_87590;
  wire [21:0] umul_87591;
  wire [20:0] add_87593;
  wire [15:0] sel_87598;
  wire [21:0] umul_87599;
  wire [21:0] add_87601;
  wire [15:0] sel_87606;
  wire [21:0] umul_87607;
  wire [21:0] add_87609;
  wire [15:0] sel_87614;
  wire [15:0] array_index_87615;
  wire [31:0] smod_87619;
  wire [15:0] array_index_87621;
  wire [31:0] smod_87625;
  wire [21:0] umul_87675;
  wire [15:0] add_87677;
  wire [15:0] sel_87682;
  wire [21:0] umul_87683;
  wire [15:0] add_87685;
  wire [15:0] sel_87690;
  wire [31:0] smod_87694;
  wire [31:0] smod_87699;
  wire [31:0] smod_87704;
  wire [31:0] smod_87709;
  wire [31:0] smod_87714;
  wire [31:0] smod_87719;
  wire [31:0] smod_87724;
  wire [31:0] smod_87729;
  wire [22:0] umul_87745;
  wire [20:0] add_87747;
  wire [15:0] sel_87752;
  wire [22:0] umul_87753;
  wire [20:0] add_87755;
  wire [15:0] sel_87760;
  wire [22:0] umul_87761;
  wire [22:0] add_87763;
  wire [15:0] sel_87768;
  wire [22:0] umul_87769;
  wire [22:0] add_87771;
  wire [15:0] sel_87776;
  wire [21:0] umul_87777;
  wire [20:0] add_87779;
  wire [15:0] sel_87784;
  wire [21:0] umul_87785;
  wire [20:0] add_87787;
  wire [15:0] sel_87792;
  wire [21:0] umul_87793;
  wire [21:0] add_87795;
  wire [15:0] sel_87800;
  wire [21:0] umul_87801;
  wire [21:0] add_87803;
  wire [15:0] sel_87808;
  wire [15:0] array_index_87809;
  wire [31:0] smod_87813;
  wire [15:0] array_index_87815;
  wire [31:0] smod_87819;
  wire [21:0] umul_87869;
  wire [15:0] add_87871;
  wire [15:0] sel_87876;
  wire [21:0] umul_87877;
  wire [15:0] add_87879;
  wire [15:0] sel_87884;
  wire [31:0] smod_87888;
  wire [31:0] smod_87893;
  wire [31:0] smod_87898;
  wire [31:0] smod_87903;
  wire [31:0] smod_87908;
  wire [31:0] smod_87913;
  wire [31:0] smod_87918;
  wire [31:0] smod_87923;
  wire [22:0] umul_87939;
  wire [20:0] add_87941;
  wire [15:0] sel_87946;
  wire [22:0] umul_87947;
  wire [20:0] add_87949;
  wire [15:0] sel_87954;
  wire [22:0] umul_87955;
  wire [22:0] add_87957;
  wire [15:0] sel_87962;
  wire [22:0] umul_87963;
  wire [22:0] add_87965;
  wire [15:0] sel_87970;
  wire [21:0] umul_87971;
  wire [20:0] add_87973;
  wire [15:0] sel_87978;
  wire [21:0] umul_87979;
  wire [20:0] add_87981;
  wire [15:0] sel_87986;
  wire [21:0] umul_87987;
  wire [21:0] add_87989;
  wire [15:0] sel_87994;
  wire [21:0] umul_87995;
  wire [21:0] add_87997;
  wire [15:0] sel_88002;
  wire [15:0] array_index_88003;
  wire [31:0] smod_88007;
  wire [15:0] array_index_88009;
  wire [31:0] smod_88013;
  wire [21:0] umul_88063;
  wire [15:0] add_88065;
  wire [15:0] sel_88070;
  wire [21:0] umul_88071;
  wire [15:0] add_88073;
  wire [15:0] sel_88078;
  wire [31:0] smod_88082;
  wire [31:0] smod_88087;
  wire [31:0] smod_88092;
  wire [31:0] smod_88097;
  wire [31:0] smod_88102;
  wire [31:0] smod_88107;
  wire [31:0] smod_88112;
  wire [31:0] smod_88117;
  wire [22:0] umul_88133;
  wire [20:0] add_88135;
  wire [15:0] sel_88140;
  wire [22:0] umul_88141;
  wire [20:0] add_88143;
  wire [15:0] sel_88148;
  wire [22:0] umul_88149;
  wire [22:0] add_88151;
  wire [15:0] sel_88156;
  wire [22:0] umul_88157;
  wire [22:0] add_88159;
  wire [15:0] sel_88164;
  wire [21:0] umul_88165;
  wire [20:0] add_88167;
  wire [15:0] sel_88172;
  wire [21:0] umul_88173;
  wire [20:0] add_88175;
  wire [15:0] sel_88180;
  wire [21:0] umul_88181;
  wire [21:0] add_88183;
  wire [15:0] sel_88188;
  wire [21:0] umul_88189;
  wire [21:0] add_88191;
  wire [15:0] sel_88196;
  wire [15:0] array_index_88197;
  wire [31:0] smod_88201;
  wire [15:0] array_index_88203;
  wire [31:0] smod_88207;
  wire [21:0] umul_88257;
  wire [15:0] add_88259;
  wire [15:0] sel_88264;
  wire [21:0] umul_88265;
  wire [15:0] add_88267;
  wire [15:0] sel_88272;
  wire [31:0] smod_88276;
  wire [31:0] smod_88281;
  wire [31:0] smod_88286;
  wire [31:0] smod_88291;
  wire [31:0] smod_88296;
  wire [31:0] smod_88301;
  wire [31:0] smod_88306;
  wire [31:0] smod_88311;
  wire [22:0] umul_88327;
  wire [20:0] add_88329;
  wire [15:0] sel_88334;
  wire [22:0] umul_88335;
  wire [20:0] add_88337;
  wire [15:0] sel_88342;
  wire [22:0] umul_88343;
  wire [22:0] add_88345;
  wire [15:0] sel_88350;
  wire [22:0] umul_88351;
  wire [22:0] add_88353;
  wire [15:0] sel_88358;
  wire [21:0] umul_88359;
  wire [20:0] add_88361;
  wire [15:0] sel_88366;
  wire [21:0] umul_88367;
  wire [20:0] add_88369;
  wire [15:0] sel_88374;
  wire [21:0] umul_88375;
  wire [21:0] add_88377;
  wire [15:0] sel_88382;
  wire [21:0] umul_88383;
  wire [21:0] add_88385;
  wire [15:0] sel_88390;
  wire [15:0] array_index_88391;
  wire [31:0] smod_88395;
  wire [15:0] array_index_88397;
  wire [31:0] smod_88401;
  wire [21:0] umul_88451;
  wire [15:0] add_88453;
  wire [15:0] sel_88458;
  wire [21:0] umul_88459;
  wire [15:0] add_88461;
  wire [15:0] sel_88466;
  wire [31:0] smod_88470;
  wire [31:0] smod_88475;
  wire [31:0] smod_88480;
  wire [31:0] smod_88485;
  wire [31:0] smod_88490;
  wire [31:0] smod_88495;
  wire [31:0] smod_88500;
  wire [31:0] smod_88505;
  wire [22:0] umul_88521;
  wire [20:0] add_88523;
  wire [15:0] sel_88528;
  wire [22:0] umul_88529;
  wire [20:0] add_88531;
  wire [15:0] sel_88536;
  wire [22:0] umul_88537;
  wire [22:0] add_88539;
  wire [15:0] sel_88544;
  wire [22:0] umul_88545;
  wire [22:0] add_88547;
  wire [15:0] sel_88552;
  wire [21:0] umul_88553;
  wire [20:0] add_88555;
  wire [15:0] sel_88560;
  wire [21:0] umul_88561;
  wire [20:0] add_88563;
  wire [15:0] sel_88568;
  wire [21:0] umul_88569;
  wire [21:0] add_88571;
  wire [15:0] sel_88576;
  wire [21:0] umul_88577;
  wire [21:0] add_88579;
  wire [15:0] sel_88584;
  wire [15:0] array_index_88585;
  wire [31:0] smod_88589;
  wire [15:0] array_index_88591;
  wire [31:0] smod_88595;
  wire [21:0] umul_88645;
  wire [15:0] add_88647;
  wire [15:0] sel_88652;
  wire [21:0] umul_88653;
  wire [15:0] add_88655;
  wire [15:0] sel_88660;
  wire [31:0] smod_88664;
  wire [31:0] smod_88669;
  wire [31:0] smod_88674;
  wire [31:0] smod_88679;
  wire [31:0] smod_88684;
  wire [31:0] smod_88689;
  wire [31:0] smod_88694;
  wire [31:0] smod_88699;
  wire [22:0] umul_88715;
  wire [20:0] add_88717;
  wire [15:0] sel_88722;
  wire [22:0] umul_88723;
  wire [20:0] add_88725;
  wire [15:0] sel_88730;
  wire [22:0] umul_88731;
  wire [22:0] add_88733;
  wire [15:0] sel_88738;
  wire [22:0] umul_88739;
  wire [22:0] add_88741;
  wire [15:0] sel_88746;
  wire [21:0] umul_88747;
  wire [20:0] add_88749;
  wire [15:0] sel_88754;
  wire [21:0] umul_88755;
  wire [20:0] add_88757;
  wire [15:0] sel_88762;
  wire [21:0] umul_88763;
  wire [21:0] add_88765;
  wire [15:0] sel_88770;
  wire [21:0] umul_88771;
  wire [21:0] add_88773;
  wire [15:0] sel_88778;
  wire [15:0] array_index_88779;
  wire [31:0] smod_88783;
  wire [15:0] array_index_88785;
  wire [31:0] smod_88789;
  wire [21:0] umul_88839;
  wire [15:0] add_88841;
  wire [15:0] sel_88846;
  wire [21:0] umul_88847;
  wire [15:0] add_88849;
  wire [15:0] sel_88854;
  wire [31:0] smod_88858;
  wire [31:0] smod_88863;
  wire [31:0] smod_88868;
  wire [31:0] smod_88873;
  wire [31:0] smod_88878;
  wire [31:0] smod_88883;
  wire [31:0] smod_88888;
  wire [31:0] smod_88893;
  wire [22:0] umul_88909;
  wire [20:0] add_88911;
  wire [15:0] sel_88916;
  wire [22:0] umul_88917;
  wire [20:0] add_88919;
  wire [15:0] sel_88924;
  wire [22:0] umul_88925;
  wire [22:0] add_88927;
  wire [15:0] sel_88932;
  wire [22:0] umul_88933;
  wire [22:0] add_88935;
  wire [15:0] sel_88940;
  wire [21:0] umul_88941;
  wire [20:0] add_88943;
  wire [15:0] sel_88948;
  wire [21:0] umul_88949;
  wire [20:0] add_88951;
  wire [15:0] sel_88956;
  wire [21:0] umul_88957;
  wire [21:0] add_88959;
  wire [15:0] sel_88964;
  wire [21:0] umul_88965;
  wire [21:0] add_88967;
  wire [15:0] sel_88972;
  wire [15:0] array_index_88973;
  wire [31:0] smod_88977;
  wire [15:0] array_index_88979;
  wire [31:0] smod_88983;
  wire [21:0] umul_89033;
  wire [15:0] add_89035;
  wire [15:0] sel_89040;
  wire [21:0] umul_89041;
  wire [15:0] add_89043;
  wire [15:0] sel_89048;
  wire [31:0] smod_89052;
  wire [31:0] smod_89057;
  wire [31:0] smod_89062;
  wire [31:0] smod_89067;
  wire [31:0] smod_89072;
  wire [31:0] smod_89077;
  wire [31:0] smod_89082;
  wire [31:0] smod_89087;
  wire [22:0] umul_89103;
  wire [20:0] add_89105;
  wire [15:0] sel_89110;
  wire [22:0] umul_89111;
  wire [20:0] add_89113;
  wire [15:0] sel_89118;
  wire [22:0] umul_89119;
  wire [22:0] add_89121;
  wire [15:0] sel_89126;
  wire [22:0] umul_89127;
  wire [22:0] add_89129;
  wire [15:0] sel_89134;
  wire [21:0] umul_89135;
  wire [20:0] add_89137;
  wire [15:0] sel_89142;
  wire [21:0] umul_89143;
  wire [20:0] add_89145;
  wire [15:0] sel_89150;
  wire [21:0] umul_89151;
  wire [21:0] add_89153;
  wire [15:0] sel_89158;
  wire [21:0] umul_89159;
  wire [21:0] add_89161;
  wire [15:0] sel_89166;
  wire [15:0] array_index_89167;
  wire [31:0] smod_89171;
  wire [15:0] array_index_89173;
  wire [31:0] smod_89177;
  wire [21:0] umul_89227;
  wire [15:0] add_89229;
  wire [15:0] sel_89234;
  wire [21:0] umul_89235;
  wire [15:0] add_89237;
  wire [15:0] sel_89242;
  wire [31:0] smod_89246;
  wire [31:0] smod_89251;
  wire [31:0] smod_89256;
  wire [31:0] smod_89261;
  wire [31:0] smod_89266;
  wire [31:0] smod_89271;
  wire [31:0] smod_89276;
  wire [31:0] smod_89281;
  wire [22:0] umul_89297;
  wire [20:0] add_89299;
  wire [15:0] sel_89304;
  wire [22:0] umul_89305;
  wire [20:0] add_89307;
  wire [15:0] sel_89312;
  wire [22:0] umul_89313;
  wire [22:0] add_89315;
  wire [15:0] sel_89320;
  wire [22:0] umul_89321;
  wire [22:0] add_89323;
  wire [15:0] sel_89328;
  wire [21:0] umul_89329;
  wire [20:0] add_89331;
  wire [15:0] sel_89336;
  wire [21:0] umul_89337;
  wire [20:0] add_89339;
  wire [15:0] sel_89344;
  wire [21:0] umul_89345;
  wire [21:0] add_89347;
  wire [15:0] sel_89352;
  wire [21:0] umul_89353;
  wire [21:0] add_89355;
  wire [15:0] sel_89360;
  wire [15:0] array_index_89361;
  wire [31:0] smod_89365;
  wire [15:0] array_index_89367;
  wire [31:0] smod_89371;
  wire [21:0] umul_89421;
  wire [15:0] add_89423;
  wire [15:0] sel_89428;
  wire [21:0] umul_89429;
  wire [15:0] add_89431;
  wire [15:0] sel_89436;
  wire [31:0] smod_89440;
  wire [31:0] smod_89445;
  wire [31:0] smod_89450;
  wire [31:0] smod_89455;
  wire [31:0] smod_89460;
  wire [31:0] smod_89465;
  wire [31:0] smod_89470;
  wire [31:0] smod_89475;
  wire [22:0] umul_89491;
  wire [20:0] add_89493;
  wire [15:0] sel_89498;
  wire [22:0] umul_89499;
  wire [20:0] add_89501;
  wire [15:0] sel_89506;
  wire [22:0] umul_89507;
  wire [22:0] add_89509;
  wire [15:0] sel_89514;
  wire [22:0] umul_89515;
  wire [22:0] add_89517;
  wire [15:0] sel_89522;
  wire [21:0] umul_89523;
  wire [20:0] add_89525;
  wire [15:0] sel_89530;
  wire [21:0] umul_89531;
  wire [20:0] add_89533;
  wire [15:0] sel_89538;
  wire [21:0] umul_89539;
  wire [21:0] add_89541;
  wire [15:0] sel_89546;
  wire [21:0] umul_89547;
  wire [21:0] add_89549;
  wire [15:0] sel_89554;
  wire [15:0] array_index_89555;
  wire [31:0] smod_89559;
  wire [15:0] array_index_89561;
  wire [31:0] smod_89565;
  wire [21:0] umul_89615;
  wire [15:0] add_89617;
  wire [15:0] sel_89622;
  wire [21:0] umul_89623;
  wire [15:0] add_89625;
  wire [15:0] sel_89630;
  wire [31:0] smod_89634;
  wire [31:0] smod_89639;
  wire [31:0] smod_89644;
  wire [31:0] smod_89649;
  wire [31:0] smod_89654;
  wire [31:0] smod_89659;
  wire [31:0] smod_89664;
  wire [31:0] smod_89669;
  wire [22:0] umul_89685;
  wire [20:0] add_89687;
  wire [15:0] sel_89692;
  wire [22:0] umul_89693;
  wire [20:0] add_89695;
  wire [15:0] sel_89700;
  wire [22:0] umul_89701;
  wire [22:0] add_89703;
  wire [15:0] sel_89708;
  wire [22:0] umul_89709;
  wire [22:0] add_89711;
  wire [15:0] sel_89716;
  wire [21:0] umul_89717;
  wire [20:0] add_89719;
  wire [15:0] sel_89724;
  wire [21:0] umul_89725;
  wire [20:0] add_89727;
  wire [15:0] sel_89732;
  wire [21:0] umul_89733;
  wire [21:0] add_89735;
  wire [15:0] sel_89740;
  wire [21:0] umul_89741;
  wire [21:0] add_89743;
  wire [15:0] sel_89748;
  wire [15:0] array_index_89749;
  wire [31:0] smod_89753;
  wire [15:0] array_index_89755;
  wire [31:0] smod_89759;
  wire [21:0] umul_89809;
  wire [15:0] add_89811;
  wire [15:0] sel_89816;
  wire [21:0] umul_89817;
  wire [15:0] add_89819;
  wire [15:0] sel_89824;
  wire [31:0] smod_89828;
  wire [31:0] smod_89833;
  wire [31:0] smod_89838;
  wire [31:0] smod_89843;
  wire [31:0] smod_89848;
  wire [31:0] smod_89853;
  wire [31:0] smod_89858;
  wire [31:0] smod_89863;
  wire [22:0] umul_89879;
  wire [20:0] add_89881;
  wire [15:0] sel_89886;
  wire [22:0] umul_89887;
  wire [20:0] add_89889;
  wire [15:0] sel_89894;
  wire [22:0] umul_89895;
  wire [22:0] add_89897;
  wire [15:0] sel_89902;
  wire [22:0] umul_89903;
  wire [22:0] add_89905;
  wire [15:0] sel_89910;
  wire [21:0] umul_89911;
  wire [20:0] add_89913;
  wire [15:0] sel_89918;
  wire [21:0] umul_89919;
  wire [20:0] add_89921;
  wire [15:0] sel_89926;
  wire [21:0] umul_89927;
  wire [21:0] add_89929;
  wire [15:0] sel_89934;
  wire [21:0] umul_89935;
  wire [21:0] add_89937;
  wire [15:0] sel_89942;
  wire [15:0] array_index_89943;
  wire [31:0] smod_89947;
  wire [15:0] array_index_89949;
  wire [31:0] smod_89953;
  wire [21:0] umul_90003;
  wire [15:0] add_90005;
  wire [15:0] sel_90010;
  wire [21:0] umul_90011;
  wire [15:0] add_90013;
  wire [15:0] sel_90018;
  wire [31:0] smod_90022;
  wire [31:0] smod_90027;
  wire [31:0] smod_90032;
  wire [31:0] smod_90037;
  wire [31:0] smod_90042;
  wire [31:0] smod_90047;
  wire [31:0] smod_90052;
  wire [31:0] smod_90057;
  wire [22:0] umul_90073;
  wire [20:0] add_90075;
  wire [15:0] sel_90080;
  wire [22:0] umul_90081;
  wire [20:0] add_90083;
  wire [15:0] sel_90088;
  wire [22:0] umul_90089;
  wire [22:0] add_90091;
  wire [15:0] sel_90096;
  wire [22:0] umul_90097;
  wire [22:0] add_90099;
  wire [15:0] sel_90104;
  wire [21:0] umul_90105;
  wire [20:0] add_90107;
  wire [15:0] sel_90112;
  wire [21:0] umul_90113;
  wire [20:0] add_90115;
  wire [15:0] sel_90120;
  wire [21:0] umul_90121;
  wire [21:0] add_90123;
  wire [15:0] sel_90128;
  wire [21:0] umul_90129;
  wire [21:0] add_90131;
  wire [15:0] sel_90136;
  wire [15:0] array_index_90137;
  wire [31:0] smod_90141;
  wire [15:0] array_index_90143;
  wire [31:0] smod_90147;
  wire [21:0] umul_90197;
  wire [15:0] add_90199;
  wire [15:0] sel_90204;
  wire [21:0] umul_90205;
  wire [15:0] add_90207;
  wire [15:0] sel_90212;
  wire [31:0] smod_90216;
  wire [31:0] smod_90221;
  wire [31:0] smod_90226;
  wire [31:0] smod_90231;
  wire [31:0] smod_90236;
  wire [31:0] smod_90241;
  wire [31:0] smod_90246;
  wire [31:0] smod_90251;
  wire [22:0] umul_90267;
  wire [20:0] add_90269;
  wire [15:0] sel_90274;
  wire [22:0] umul_90275;
  wire [20:0] add_90277;
  wire [15:0] sel_90282;
  wire [22:0] umul_90283;
  wire [22:0] add_90285;
  wire [15:0] sel_90290;
  wire [22:0] umul_90291;
  wire [22:0] add_90293;
  wire [15:0] sel_90298;
  wire [21:0] umul_90299;
  wire [20:0] add_90301;
  wire [15:0] sel_90306;
  wire [21:0] umul_90307;
  wire [20:0] add_90309;
  wire [15:0] sel_90314;
  wire [21:0] umul_90315;
  wire [21:0] add_90317;
  wire [15:0] sel_90322;
  wire [21:0] umul_90323;
  wire [21:0] add_90325;
  wire [15:0] sel_90330;
  wire [15:0] array_index_90331;
  wire [31:0] smod_90335;
  wire [15:0] array_index_90337;
  wire [31:0] smod_90341;
  wire [21:0] umul_90391;
  wire [15:0] add_90393;
  wire [15:0] sel_90398;
  wire [21:0] umul_90399;
  wire [15:0] add_90401;
  wire [15:0] sel_90406;
  wire [31:0] smod_90410;
  wire [31:0] smod_90415;
  wire [31:0] smod_90420;
  wire [31:0] smod_90425;
  wire [31:0] smod_90430;
  wire [31:0] smod_90435;
  wire [31:0] smod_90440;
  wire [31:0] smod_90445;
  wire [22:0] umul_90461;
  wire [20:0] add_90463;
  wire [15:0] sel_90468;
  wire [22:0] umul_90469;
  wire [20:0] add_90471;
  wire [15:0] sel_90476;
  wire [22:0] umul_90477;
  wire [22:0] add_90479;
  wire [15:0] sel_90484;
  wire [22:0] umul_90485;
  wire [22:0] add_90487;
  wire [15:0] sel_90492;
  wire [21:0] umul_90493;
  wire [20:0] add_90495;
  wire [15:0] sel_90500;
  wire [21:0] umul_90501;
  wire [20:0] add_90503;
  wire [15:0] sel_90508;
  wire [21:0] umul_90509;
  wire [21:0] add_90511;
  wire [15:0] sel_90516;
  wire [21:0] umul_90517;
  wire [21:0] add_90519;
  wire [15:0] sel_90524;
  wire [15:0] array_index_90525;
  wire [31:0] smod_90529;
  wire [15:0] array_index_90531;
  wire [31:0] smod_90535;
  wire [21:0] umul_90585;
  wire [15:0] add_90587;
  wire [15:0] sel_90592;
  wire [21:0] umul_90593;
  wire [15:0] add_90595;
  wire [15:0] sel_90600;
  wire [31:0] smod_90604;
  wire [31:0] smod_90609;
  wire [31:0] smod_90614;
  wire [31:0] smod_90619;
  wire [31:0] smod_90624;
  wire [31:0] smod_90629;
  wire [31:0] smod_90634;
  wire [31:0] smod_90639;
  wire [22:0] umul_90655;
  wire [20:0] add_90657;
  wire [15:0] sel_90662;
  wire [22:0] umul_90663;
  wire [20:0] add_90665;
  wire [15:0] sel_90670;
  wire [22:0] umul_90671;
  wire [22:0] add_90673;
  wire [15:0] sel_90678;
  wire [22:0] umul_90679;
  wire [22:0] add_90681;
  wire [15:0] sel_90686;
  wire [21:0] umul_90687;
  wire [20:0] add_90689;
  wire [15:0] sel_90694;
  wire [21:0] umul_90695;
  wire [20:0] add_90697;
  wire [15:0] sel_90702;
  wire [21:0] umul_90703;
  wire [21:0] add_90705;
  wire [15:0] sel_90710;
  wire [21:0] umul_90711;
  wire [21:0] add_90713;
  wire [15:0] sel_90718;
  wire [15:0] array_index_90719;
  wire [31:0] smod_90723;
  wire [15:0] array_index_90725;
  wire [31:0] smod_90729;
  wire [21:0] umul_90779;
  wire [15:0] add_90781;
  wire [15:0] sel_90786;
  wire [21:0] umul_90787;
  wire [15:0] add_90789;
  wire [15:0] sel_90794;
  wire [31:0] smod_90798;
  wire [31:0] smod_90803;
  wire [31:0] smod_90808;
  wire [31:0] smod_90813;
  wire [31:0] smod_90818;
  wire [31:0] smod_90823;
  wire [31:0] smod_90828;
  wire [31:0] smod_90833;
  wire [22:0] umul_90849;
  wire [20:0] add_90851;
  wire [15:0] sel_90856;
  wire [22:0] umul_90857;
  wire [20:0] add_90859;
  wire [15:0] sel_90864;
  wire [22:0] umul_90865;
  wire [22:0] add_90867;
  wire [15:0] sel_90872;
  wire [22:0] umul_90873;
  wire [22:0] add_90875;
  wire [15:0] sel_90880;
  wire [21:0] umul_90881;
  wire [20:0] add_90883;
  wire [15:0] sel_90888;
  wire [21:0] umul_90889;
  wire [20:0] add_90891;
  wire [15:0] sel_90896;
  wire [21:0] umul_90897;
  wire [21:0] add_90899;
  wire [15:0] sel_90904;
  wire [21:0] umul_90905;
  wire [21:0] add_90907;
  wire [15:0] sel_90912;
  wire [15:0] array_index_90913;
  wire [31:0] smod_90917;
  wire [15:0] array_index_90919;
  wire [31:0] smod_90923;
  wire [21:0] umul_90973;
  wire [15:0] add_90975;
  wire [15:0] sel_90980;
  wire [21:0] umul_90981;
  wire [15:0] add_90983;
  wire [15:0] sel_90988;
  wire [31:0] smod_90992;
  wire [31:0] smod_90997;
  wire [31:0] smod_91002;
  wire [31:0] smod_91007;
  wire [31:0] smod_91012;
  wire [31:0] smod_91017;
  wire [31:0] smod_91022;
  wire [31:0] smod_91027;
  wire [22:0] umul_91043;
  wire [20:0] add_91045;
  wire [15:0] sel_91050;
  wire [22:0] umul_91051;
  wire [20:0] add_91053;
  wire [15:0] sel_91058;
  wire [22:0] umul_91059;
  wire [22:0] add_91061;
  wire [15:0] sel_91066;
  wire [22:0] umul_91067;
  wire [22:0] add_91069;
  wire [15:0] sel_91074;
  wire [21:0] umul_91075;
  wire [20:0] add_91077;
  wire [15:0] sel_91082;
  wire [21:0] umul_91083;
  wire [20:0] add_91085;
  wire [15:0] sel_91090;
  wire [21:0] umul_91091;
  wire [21:0] add_91093;
  wire [15:0] sel_91098;
  wire [21:0] umul_91099;
  wire [21:0] add_91101;
  wire [15:0] sel_91106;
  wire [15:0] array_index_91107;
  wire [31:0] smod_91111;
  wire [15:0] array_index_91113;
  wire [31:0] smod_91117;
  wire [21:0] umul_91167;
  wire [15:0] add_91169;
  wire [15:0] sel_91174;
  wire [21:0] umul_91175;
  wire [15:0] add_91177;
  wire [15:0] sel_91182;
  wire [31:0] smod_91186;
  wire [31:0] smod_91191;
  wire [31:0] smod_91196;
  wire [31:0] smod_91201;
  wire [31:0] smod_91206;
  wire [31:0] smod_91211;
  wire [31:0] smod_91216;
  wire [31:0] smod_91221;
  wire [22:0] umul_91237;
  wire [20:0] add_91239;
  wire [15:0] sel_91244;
  wire [22:0] umul_91245;
  wire [20:0] add_91247;
  wire [15:0] sel_91252;
  wire [22:0] umul_91253;
  wire [22:0] add_91255;
  wire [15:0] sel_91260;
  wire [22:0] umul_91261;
  wire [22:0] add_91263;
  wire [15:0] sel_91268;
  wire [21:0] umul_91269;
  wire [20:0] add_91271;
  wire [15:0] sel_91276;
  wire [21:0] umul_91277;
  wire [20:0] add_91279;
  wire [15:0] sel_91284;
  wire [21:0] umul_91285;
  wire [21:0] add_91287;
  wire [15:0] sel_91292;
  wire [21:0] umul_91293;
  wire [21:0] add_91295;
  wire [15:0] sel_91300;
  wire [15:0] array_index_91301;
  wire [31:0] smod_91305;
  wire [15:0] array_index_91307;
  wire [31:0] smod_91311;
  wire [21:0] umul_91361;
  wire [15:0] add_91363;
  wire [15:0] sel_91368;
  wire [21:0] umul_91369;
  wire [15:0] add_91371;
  wire [15:0] sel_91376;
  wire [31:0] smod_91380;
  wire [31:0] smod_91385;
  wire [31:0] smod_91390;
  wire [31:0] smod_91395;
  wire [31:0] smod_91400;
  wire [31:0] smod_91405;
  wire [31:0] smod_91410;
  wire [31:0] smod_91415;
  wire [22:0] umul_91431;
  wire [20:0] add_91433;
  wire [15:0] sel_91438;
  wire [22:0] umul_91439;
  wire [20:0] add_91441;
  wire [15:0] sel_91446;
  wire [22:0] umul_91447;
  wire [22:0] add_91449;
  wire [15:0] sel_91454;
  wire [22:0] umul_91455;
  wire [22:0] add_91457;
  wire [15:0] sel_91462;
  wire [21:0] umul_91463;
  wire [20:0] add_91465;
  wire [15:0] sel_91470;
  wire [21:0] umul_91471;
  wire [20:0] add_91473;
  wire [15:0] sel_91478;
  wire [21:0] umul_91479;
  wire [21:0] add_91481;
  wire [15:0] sel_91486;
  wire [21:0] umul_91487;
  wire [21:0] add_91489;
  wire [15:0] sel_91494;
  wire [15:0] array_index_91495;
  wire [31:0] smod_91499;
  wire [15:0] array_index_91501;
  wire [31:0] smod_91505;
  wire [21:0] umul_91555;
  wire [15:0] add_91557;
  wire [15:0] sel_91562;
  wire [21:0] umul_91563;
  wire [15:0] add_91565;
  wire [15:0] sel_91570;
  wire [31:0] smod_91574;
  wire [31:0] smod_91579;
  wire [31:0] smod_91584;
  wire [31:0] smod_91589;
  wire [31:0] smod_91594;
  wire [31:0] smod_91599;
  wire [31:0] smod_91604;
  wire [31:0] smod_91609;
  wire [22:0] umul_91625;
  wire [20:0] add_91627;
  wire [15:0] sel_91632;
  wire [22:0] umul_91633;
  wire [20:0] add_91635;
  wire [15:0] sel_91640;
  wire [22:0] umul_91641;
  wire [22:0] add_91643;
  wire [15:0] sel_91648;
  wire [22:0] umul_91649;
  wire [22:0] add_91651;
  wire [15:0] sel_91656;
  wire [21:0] umul_91657;
  wire [20:0] add_91659;
  wire [15:0] sel_91664;
  wire [21:0] umul_91665;
  wire [20:0] add_91667;
  wire [15:0] sel_91672;
  wire [21:0] umul_91673;
  wire [21:0] add_91675;
  wire [15:0] sel_91680;
  wire [21:0] umul_91681;
  wire [21:0] add_91683;
  wire [15:0] sel_91688;
  wire [15:0] array_index_91689;
  wire [31:0] smod_91693;
  wire [15:0] array_index_91695;
  wire [31:0] smod_91699;
  wire [21:0] umul_91749;
  wire [15:0] add_91751;
  wire [15:0] sel_91756;
  wire [21:0] umul_91757;
  wire [15:0] add_91759;
  wire [15:0] sel_91764;
  wire [31:0] smod_91768;
  wire [31:0] smod_91773;
  wire [31:0] smod_91778;
  wire [31:0] smod_91783;
  wire [31:0] smod_91788;
  wire [31:0] smod_91793;
  wire [31:0] smod_91798;
  wire [31:0] smod_91803;
  wire [22:0] umul_91819;
  wire [20:0] add_91821;
  wire [15:0] sel_91826;
  wire [22:0] umul_91827;
  wire [20:0] add_91829;
  wire [15:0] sel_91834;
  wire [22:0] umul_91835;
  wire [22:0] add_91837;
  wire [15:0] sel_91842;
  wire [22:0] umul_91843;
  wire [22:0] add_91845;
  wire [15:0] sel_91850;
  wire [21:0] umul_91851;
  wire [20:0] add_91853;
  wire [15:0] sel_91858;
  wire [21:0] umul_91859;
  wire [20:0] add_91861;
  wire [15:0] sel_91866;
  wire [21:0] umul_91867;
  wire [21:0] add_91869;
  wire [15:0] sel_91874;
  wire [21:0] umul_91875;
  wire [21:0] add_91877;
  wire [15:0] sel_91882;
  wire [15:0] array_index_91883;
  wire [31:0] smod_91887;
  wire [15:0] array_index_91889;
  wire [31:0] smod_91893;
  wire [21:0] umul_91943;
  wire [15:0] add_91945;
  wire [15:0] sel_91950;
  wire [21:0] umul_91951;
  wire [15:0] add_91953;
  wire [15:0] sel_91958;
  wire [31:0] smod_91962;
  wire [31:0] smod_91967;
  wire [31:0] smod_91972;
  wire [31:0] smod_91977;
  wire [31:0] smod_91982;
  wire [31:0] smod_91987;
  wire [31:0] smod_91992;
  wire [31:0] smod_91997;
  wire [22:0] umul_92013;
  wire [20:0] add_92015;
  wire [15:0] sel_92020;
  wire [22:0] umul_92021;
  wire [20:0] add_92023;
  wire [15:0] sel_92028;
  wire [22:0] umul_92029;
  wire [22:0] add_92031;
  wire [15:0] sel_92036;
  wire [22:0] umul_92037;
  wire [22:0] add_92039;
  wire [15:0] sel_92044;
  wire [21:0] umul_92045;
  wire [20:0] add_92047;
  wire [15:0] sel_92052;
  wire [21:0] umul_92053;
  wire [20:0] add_92055;
  wire [15:0] sel_92060;
  wire [21:0] umul_92061;
  wire [21:0] add_92063;
  wire [15:0] sel_92068;
  wire [21:0] umul_92069;
  wire [21:0] add_92071;
  wire [15:0] sel_92076;
  wire [15:0] array_index_92077;
  wire [31:0] smod_92081;
  wire [15:0] array_index_92083;
  wire [31:0] smod_92087;
  wire [21:0] umul_92137;
  wire [15:0] add_92139;
  wire [15:0] sel_92144;
  wire [21:0] umul_92145;
  wire [15:0] add_92147;
  wire [15:0] sel_92152;
  wire [31:0] smod_92156;
  wire [31:0] smod_92161;
  wire [31:0] smod_92166;
  wire [31:0] smod_92171;
  wire [31:0] smod_92176;
  wire [31:0] smod_92181;
  wire [31:0] smod_92186;
  wire [31:0] smod_92191;
  wire [22:0] umul_92207;
  wire [20:0] add_92209;
  wire [15:0] sel_92214;
  wire [22:0] umul_92215;
  wire [20:0] add_92217;
  wire [15:0] sel_92222;
  wire [22:0] umul_92223;
  wire [22:0] add_92225;
  wire [15:0] sel_92230;
  wire [22:0] umul_92231;
  wire [22:0] add_92233;
  wire [15:0] sel_92238;
  wire [21:0] umul_92239;
  wire [20:0] add_92241;
  wire [15:0] sel_92246;
  wire [21:0] umul_92247;
  wire [20:0] add_92249;
  wire [15:0] sel_92254;
  wire [21:0] umul_92255;
  wire [21:0] add_92257;
  wire [15:0] sel_92262;
  wire [21:0] umul_92263;
  wire [21:0] add_92265;
  wire [15:0] sel_92270;
  wire [15:0] array_index_92271;
  wire [31:0] smod_92275;
  wire [15:0] array_index_92277;
  wire [31:0] smod_92281;
  wire [21:0] umul_92331;
  wire [15:0] add_92333;
  wire [15:0] sel_92338;
  wire [21:0] umul_92339;
  wire [15:0] add_92341;
  wire [15:0] sel_92346;
  wire [31:0] smod_92350;
  wire [31:0] smod_92355;
  wire [31:0] smod_92360;
  wire [31:0] smod_92365;
  wire [31:0] smod_92370;
  wire [31:0] smod_92375;
  wire [31:0] smod_92380;
  wire [31:0] smod_92385;
  wire [22:0] umul_92401;
  wire [20:0] add_92403;
  wire [15:0] sel_92408;
  wire [22:0] umul_92409;
  wire [20:0] add_92411;
  wire [15:0] sel_92416;
  wire [22:0] umul_92417;
  wire [22:0] add_92419;
  wire [15:0] sel_92424;
  wire [22:0] umul_92425;
  wire [22:0] add_92427;
  wire [15:0] sel_92432;
  wire [21:0] umul_92433;
  wire [20:0] add_92435;
  wire [15:0] sel_92440;
  wire [21:0] umul_92441;
  wire [20:0] add_92443;
  wire [15:0] sel_92448;
  wire [21:0] umul_92449;
  wire [21:0] add_92451;
  wire [15:0] sel_92456;
  wire [21:0] umul_92457;
  wire [21:0] add_92459;
  wire [15:0] sel_92464;
  wire [15:0] array_index_92465;
  wire [31:0] smod_92469;
  wire [15:0] array_index_92471;
  wire [31:0] smod_92475;
  wire [21:0] umul_92525;
  wire [15:0] add_92527;
  wire [15:0] sel_92532;
  wire [21:0] umul_92533;
  wire [15:0] add_92535;
  wire [15:0] sel_92540;
  wire [31:0] smod_92544;
  wire [31:0] smod_92549;
  wire [31:0] smod_92554;
  wire [31:0] smod_92559;
  wire [31:0] smod_92564;
  wire [31:0] smod_92569;
  wire [31:0] smod_92574;
  wire [31:0] smod_92579;
  wire [22:0] umul_92595;
  wire [20:0] add_92597;
  wire [15:0] sel_92602;
  wire [22:0] umul_92603;
  wire [20:0] add_92605;
  wire [15:0] sel_92610;
  wire [22:0] umul_92611;
  wire [22:0] add_92613;
  wire [15:0] sel_92618;
  wire [22:0] umul_92619;
  wire [22:0] add_92621;
  wire [15:0] sel_92626;
  wire [21:0] umul_92627;
  wire [20:0] add_92629;
  wire [15:0] sel_92634;
  wire [21:0] umul_92635;
  wire [20:0] add_92637;
  wire [15:0] sel_92642;
  wire [21:0] umul_92643;
  wire [21:0] add_92645;
  wire [15:0] sel_92650;
  wire [21:0] umul_92651;
  wire [21:0] add_92653;
  wire [15:0] sel_92658;
  wire [15:0] array_index_92659;
  wire [31:0] smod_92663;
  wire [15:0] array_index_92665;
  wire [31:0] smod_92669;
  wire [21:0] umul_92719;
  wire [15:0] add_92721;
  wire [15:0] sel_92726;
  wire [21:0] umul_92727;
  wire [15:0] add_92729;
  wire [15:0] sel_92734;
  wire [31:0] smod_92738;
  wire [31:0] smod_92743;
  wire [31:0] smod_92748;
  wire [31:0] smod_92753;
  wire [31:0] smod_92758;
  wire [31:0] smod_92763;
  wire [31:0] smod_92768;
  wire [31:0] smod_92773;
  wire [22:0] umul_92789;
  wire [20:0] add_92791;
  wire [15:0] sel_92796;
  wire [22:0] umul_92797;
  wire [20:0] add_92799;
  wire [15:0] sel_92804;
  wire [22:0] umul_92805;
  wire [22:0] add_92807;
  wire [15:0] sel_92812;
  wire [22:0] umul_92813;
  wire [22:0] add_92815;
  wire [15:0] sel_92820;
  wire [21:0] umul_92821;
  wire [20:0] add_92823;
  wire [15:0] sel_92828;
  wire [21:0] umul_92829;
  wire [20:0] add_92831;
  wire [15:0] sel_92836;
  wire [21:0] umul_92837;
  wire [21:0] add_92839;
  wire [15:0] sel_92844;
  wire [21:0] umul_92845;
  wire [21:0] add_92847;
  wire [15:0] sel_92852;
  wire [15:0] array_index_92853;
  wire [31:0] smod_92857;
  wire [15:0] array_index_92859;
  wire [31:0] smod_92863;
  wire [21:0] umul_92913;
  wire [15:0] add_92915;
  wire [15:0] sel_92920;
  wire [21:0] umul_92921;
  wire [15:0] add_92923;
  wire [15:0] sel_92928;
  wire [31:0] smod_92932;
  wire [31:0] smod_92937;
  wire [31:0] smod_92942;
  wire [31:0] smod_92947;
  wire [31:0] smod_92952;
  wire [31:0] smod_92957;
  wire [31:0] smod_92962;
  wire [31:0] smod_92967;
  wire [22:0] umul_92983;
  wire [20:0] add_92985;
  wire [15:0] sel_92990;
  wire [22:0] umul_92991;
  wire [20:0] add_92993;
  wire [15:0] sel_92998;
  wire [22:0] umul_92999;
  wire [22:0] add_93001;
  wire [15:0] sel_93006;
  wire [22:0] umul_93007;
  wire [22:0] add_93009;
  wire [15:0] sel_93014;
  wire [21:0] umul_93015;
  wire [20:0] add_93017;
  wire [15:0] sel_93022;
  wire [21:0] umul_93023;
  wire [20:0] add_93025;
  wire [15:0] sel_93030;
  wire [21:0] umul_93031;
  wire [21:0] add_93033;
  wire [15:0] sel_93038;
  wire [21:0] umul_93039;
  wire [21:0] add_93041;
  wire [15:0] sel_93046;
  wire [15:0] array_index_93047;
  wire [31:0] smod_93051;
  wire [15:0] array_index_93053;
  wire [31:0] smod_93057;
  wire [21:0] umul_93107;
  wire [15:0] add_93109;
  wire [15:0] sel_93114;
  wire [21:0] umul_93115;
  wire [15:0] add_93117;
  wire [15:0] sel_93122;
  wire [31:0] smod_93126;
  wire [31:0] smod_93131;
  wire [31:0] smod_93136;
  wire [31:0] smod_93141;
  wire [31:0] smod_93146;
  wire [31:0] smod_93151;
  wire [31:0] smod_93156;
  wire [31:0] smod_93161;
  wire [22:0] umul_93177;
  wire [20:0] add_93179;
  wire [15:0] sel_93184;
  wire [22:0] umul_93185;
  wire [20:0] add_93187;
  wire [15:0] sel_93192;
  wire [22:0] umul_93193;
  wire [22:0] add_93195;
  wire [15:0] sel_93200;
  wire [22:0] umul_93201;
  wire [22:0] add_93203;
  wire [15:0] sel_93208;
  wire [21:0] umul_93209;
  wire [20:0] add_93211;
  wire [15:0] sel_93216;
  wire [21:0] umul_93217;
  wire [20:0] add_93219;
  wire [15:0] sel_93224;
  wire [21:0] umul_93225;
  wire [21:0] add_93227;
  wire [15:0] sel_93232;
  wire [21:0] umul_93233;
  wire [21:0] add_93235;
  wire [15:0] sel_93240;
  wire [15:0] array_index_93241;
  wire [31:0] smod_93245;
  wire [15:0] array_index_93247;
  wire [31:0] smod_93251;
  wire [21:0] umul_93301;
  wire [15:0] add_93303;
  wire [15:0] sel_93308;
  wire [21:0] umul_93309;
  wire [15:0] add_93311;
  wire [15:0] sel_93316;
  wire [31:0] smod_93320;
  wire [31:0] smod_93325;
  wire [31:0] smod_93330;
  wire [31:0] smod_93335;
  wire [31:0] smod_93340;
  wire [31:0] smod_93345;
  wire [31:0] smod_93350;
  wire [31:0] smod_93355;
  wire [22:0] umul_93371;
  wire [20:0] add_93373;
  wire [15:0] sel_93378;
  wire [22:0] umul_93379;
  wire [20:0] add_93381;
  wire [15:0] sel_93386;
  wire [22:0] umul_93387;
  wire [22:0] add_93389;
  wire [15:0] sel_93394;
  wire [22:0] umul_93395;
  wire [22:0] add_93397;
  wire [15:0] sel_93402;
  wire [21:0] umul_93403;
  wire [20:0] add_93405;
  wire [15:0] sel_93410;
  wire [21:0] umul_93411;
  wire [20:0] add_93413;
  wire [15:0] sel_93418;
  wire [21:0] umul_93419;
  wire [21:0] add_93421;
  wire [15:0] sel_93426;
  wire [21:0] umul_93427;
  wire [21:0] add_93429;
  wire [15:0] sel_93434;
  wire [15:0] array_index_93435;
  wire [31:0] smod_93439;
  wire [15:0] array_index_93441;
  wire [31:0] smod_93445;
  wire [21:0] umul_93495;
  wire [15:0] add_93497;
  wire [15:0] sel_93502;
  wire [21:0] umul_93503;
  wire [15:0] add_93505;
  wire [15:0] sel_93510;
  wire [31:0] smod_93514;
  wire [31:0] smod_93519;
  wire [31:0] smod_93524;
  wire [31:0] smod_93529;
  wire [31:0] smod_93534;
  wire [31:0] smod_93539;
  wire [31:0] smod_93544;
  wire [31:0] smod_93549;
  wire [22:0] umul_93565;
  wire [20:0] add_93567;
  wire [15:0] sel_93572;
  wire [22:0] umul_93573;
  wire [20:0] add_93575;
  wire [15:0] sel_93580;
  wire [22:0] umul_93581;
  wire [22:0] add_93583;
  wire [15:0] sel_93588;
  wire [22:0] umul_93589;
  wire [22:0] add_93591;
  wire [15:0] sel_93596;
  wire [21:0] umul_93597;
  wire [20:0] add_93599;
  wire [15:0] sel_93604;
  wire [21:0] umul_93605;
  wire [20:0] add_93607;
  wire [15:0] sel_93612;
  wire [21:0] umul_93613;
  wire [21:0] add_93615;
  wire [15:0] sel_93620;
  wire [21:0] umul_93621;
  wire [21:0] add_93623;
  wire [15:0] sel_93628;
  wire [15:0] array_index_93629;
  wire [31:0] smod_93633;
  wire [15:0] array_index_93635;
  wire [31:0] smod_93639;
  wire [21:0] umul_93689;
  wire [15:0] add_93691;
  wire [15:0] sel_93696;
  wire [21:0] umul_93697;
  wire [15:0] add_93699;
  wire [15:0] sel_93704;
  wire [31:0] smod_93708;
  wire [31:0] smod_93713;
  wire [31:0] smod_93718;
  wire [31:0] smod_93723;
  wire [31:0] smod_93728;
  wire [31:0] smod_93733;
  wire [31:0] smod_93738;
  wire [31:0] smod_93743;
  wire [22:0] umul_93759;
  wire [20:0] add_93761;
  wire [15:0] sel_93766;
  wire [22:0] umul_93767;
  wire [20:0] add_93769;
  wire [15:0] sel_93774;
  wire [22:0] umul_93775;
  wire [22:0] add_93777;
  wire [15:0] sel_93782;
  wire [22:0] umul_93783;
  wire [22:0] add_93785;
  wire [15:0] sel_93790;
  wire [21:0] umul_93791;
  wire [20:0] add_93793;
  wire [15:0] sel_93798;
  wire [21:0] umul_93799;
  wire [20:0] add_93801;
  wire [15:0] sel_93806;
  wire [21:0] umul_93807;
  wire [21:0] add_93809;
  wire [15:0] sel_93814;
  wire [21:0] umul_93815;
  wire [21:0] add_93817;
  wire [15:0] sel_93822;
  wire [15:0] array_index_93823;
  wire [31:0] smod_93827;
  wire [15:0] array_index_93829;
  wire [31:0] smod_93833;
  wire [21:0] umul_93883;
  wire [15:0] add_93885;
  wire [15:0] sel_93890;
  wire [21:0] umul_93891;
  wire [15:0] add_93893;
  wire [15:0] sel_93898;
  wire [31:0] smod_93902;
  wire [31:0] smod_93907;
  wire [31:0] smod_93912;
  wire [31:0] smod_93917;
  wire [31:0] smod_93922;
  wire [31:0] smod_93927;
  wire [31:0] smod_93932;
  wire [31:0] smod_93937;
  wire [22:0] umul_93953;
  wire [20:0] add_93955;
  wire [15:0] sel_93960;
  wire [22:0] umul_93961;
  wire [20:0] add_93963;
  wire [15:0] sel_93968;
  wire [22:0] umul_93969;
  wire [22:0] add_93971;
  wire [15:0] sel_93976;
  wire [22:0] umul_93977;
  wire [22:0] add_93979;
  wire [15:0] sel_93984;
  wire [21:0] umul_93985;
  wire [20:0] add_93987;
  wire [15:0] sel_93992;
  wire [21:0] umul_93993;
  wire [20:0] add_93995;
  wire [15:0] sel_94000;
  wire [21:0] umul_94001;
  wire [21:0] add_94003;
  wire [15:0] sel_94008;
  wire [21:0] umul_94009;
  wire [21:0] add_94011;
  wire [15:0] sel_94016;
  wire [15:0] array_index_94017;
  wire [31:0] smod_94021;
  wire [15:0] array_index_94023;
  wire [31:0] smod_94027;
  wire [21:0] umul_94077;
  wire [15:0] add_94079;
  wire [15:0] sel_94084;
  wire [21:0] umul_94085;
  wire [15:0] add_94087;
  wire [15:0] sel_94092;
  wire [31:0] smod_94096;
  wire [31:0] smod_94101;
  wire [31:0] smod_94106;
  wire [31:0] smod_94111;
  wire [31:0] smod_94116;
  wire [31:0] smod_94121;
  wire [31:0] smod_94126;
  wire [31:0] smod_94131;
  wire [22:0] umul_94147;
  wire [20:0] add_94149;
  wire [15:0] sel_94154;
  wire [22:0] umul_94155;
  wire [20:0] add_94157;
  wire [15:0] sel_94162;
  wire [22:0] umul_94163;
  wire [22:0] add_94165;
  wire [15:0] sel_94170;
  wire [22:0] umul_94171;
  wire [22:0] add_94173;
  wire [15:0] sel_94178;
  wire [21:0] umul_94179;
  wire [20:0] add_94181;
  wire [15:0] sel_94186;
  wire [21:0] umul_94187;
  wire [20:0] add_94189;
  wire [15:0] sel_94194;
  wire [21:0] umul_94195;
  wire [21:0] add_94197;
  wire [15:0] sel_94202;
  wire [21:0] umul_94203;
  wire [21:0] add_94205;
  wire [15:0] sel_94210;
  wire [15:0] array_index_94211;
  wire [31:0] smod_94215;
  wire [15:0] array_index_94217;
  wire [31:0] smod_94221;
  wire [21:0] umul_94271;
  wire [15:0] add_94273;
  wire [15:0] sel_94278;
  wire [21:0] umul_94279;
  wire [15:0] add_94281;
  wire [15:0] sel_94286;
  wire [31:0] smod_94290;
  wire [31:0] smod_94295;
  wire [31:0] smod_94300;
  wire [31:0] smod_94305;
  wire [31:0] smod_94310;
  wire [31:0] smod_94315;
  wire [31:0] smod_94320;
  wire [31:0] smod_94325;
  wire [22:0] umul_94341;
  wire [20:0] add_94343;
  wire [15:0] sel_94348;
  wire [22:0] umul_94349;
  wire [20:0] add_94351;
  wire [15:0] sel_94356;
  wire [22:0] umul_94357;
  wire [22:0] add_94359;
  wire [15:0] sel_94364;
  wire [22:0] umul_94365;
  wire [22:0] add_94367;
  wire [15:0] sel_94372;
  wire [21:0] umul_94373;
  wire [20:0] add_94375;
  wire [15:0] sel_94380;
  wire [21:0] umul_94381;
  wire [20:0] add_94383;
  wire [15:0] sel_94388;
  wire [21:0] umul_94389;
  wire [21:0] add_94391;
  wire [15:0] sel_94396;
  wire [21:0] umul_94397;
  wire [21:0] add_94399;
  wire [15:0] sel_94404;
  wire [15:0] array_index_94405;
  wire [31:0] smod_94409;
  wire [15:0] array_index_94411;
  wire [31:0] smod_94415;
  wire [21:0] umul_94465;
  wire [15:0] add_94467;
  wire [15:0] sel_94472;
  wire [21:0] umul_94473;
  wire [15:0] add_94475;
  wire [15:0] sel_94480;
  wire [31:0] smod_94484;
  wire [31:0] smod_94489;
  wire [31:0] smod_94494;
  wire [31:0] smod_94499;
  wire [31:0] smod_94504;
  wire [31:0] smod_94509;
  wire [31:0] smod_94514;
  wire [31:0] smod_94519;
  wire [22:0] umul_94535;
  wire [20:0] add_94537;
  wire [15:0] sel_94542;
  wire [22:0] umul_94543;
  wire [20:0] add_94545;
  wire [15:0] sel_94550;
  wire [22:0] umul_94551;
  wire [22:0] add_94553;
  wire [15:0] sel_94558;
  wire [22:0] umul_94559;
  wire [22:0] add_94561;
  wire [15:0] sel_94566;
  wire [21:0] umul_94567;
  wire [20:0] add_94569;
  wire [15:0] sel_94574;
  wire [21:0] umul_94575;
  wire [20:0] add_94577;
  wire [15:0] sel_94582;
  wire [21:0] umul_94583;
  wire [21:0] add_94585;
  wire [15:0] sel_94590;
  wire [21:0] umul_94591;
  wire [21:0] add_94593;
  wire [15:0] sel_94598;
  wire [15:0] array_index_94599;
  wire [31:0] smod_94603;
  wire [15:0] array_index_94605;
  wire [31:0] smod_94609;
  wire [21:0] umul_94659;
  wire [15:0] add_94661;
  wire [15:0] sel_94666;
  wire [21:0] umul_94667;
  wire [15:0] add_94669;
  wire [15:0] sel_94674;
  wire [31:0] smod_94678;
  wire [31:0] smod_94683;
  wire [31:0] smod_94688;
  wire [31:0] smod_94693;
  wire [31:0] smod_94698;
  wire [31:0] smod_94703;
  wire [31:0] smod_94708;
  wire [31:0] smod_94713;
  wire [22:0] umul_94729;
  wire [20:0] add_94731;
  wire [15:0] sel_94736;
  wire [22:0] umul_94737;
  wire [20:0] add_94739;
  wire [15:0] sel_94744;
  wire [22:0] umul_94745;
  wire [22:0] add_94747;
  wire [15:0] sel_94752;
  wire [22:0] umul_94753;
  wire [22:0] add_94755;
  wire [15:0] sel_94760;
  wire [21:0] umul_94761;
  wire [20:0] add_94763;
  wire [15:0] sel_94768;
  wire [21:0] umul_94769;
  wire [20:0] add_94771;
  wire [15:0] sel_94776;
  wire [21:0] umul_94777;
  wire [21:0] add_94779;
  wire [15:0] sel_94784;
  wire [21:0] umul_94785;
  wire [21:0] add_94787;
  wire [15:0] sel_94792;
  wire [15:0] array_index_94793;
  wire [31:0] smod_94797;
  wire [15:0] array_index_94799;
  wire [31:0] smod_94803;
  wire [21:0] umul_94853;
  wire [15:0] add_94855;
  wire [15:0] sel_94860;
  wire [21:0] umul_94861;
  wire [15:0] add_94863;
  wire [15:0] sel_94868;
  wire [31:0] smod_94872;
  wire [31:0] smod_94877;
  wire [31:0] smod_94882;
  wire [31:0] smod_94887;
  wire [31:0] smod_94892;
  wire [31:0] smod_94897;
  wire [31:0] smod_94902;
  wire [31:0] smod_94907;
  wire [22:0] umul_94923;
  wire [20:0] add_94925;
  wire [15:0] sel_94930;
  wire [22:0] umul_94931;
  wire [20:0] add_94933;
  wire [15:0] sel_94938;
  wire [22:0] umul_94939;
  wire [22:0] add_94941;
  wire [15:0] sel_94946;
  wire [22:0] umul_94947;
  wire [22:0] add_94949;
  wire [15:0] sel_94954;
  wire [21:0] umul_94955;
  wire [20:0] add_94957;
  wire [15:0] sel_94962;
  wire [21:0] umul_94963;
  wire [20:0] add_94965;
  wire [15:0] sel_94970;
  wire [21:0] umul_94971;
  wire [21:0] add_94973;
  wire [15:0] sel_94978;
  wire [21:0] umul_94979;
  wire [21:0] add_94981;
  wire [15:0] sel_94986;
  wire [15:0] array_index_94987;
  wire [31:0] smod_94991;
  wire [15:0] array_index_94993;
  wire [31:0] smod_94997;
  wire [21:0] umul_95047;
  wire [15:0] add_95049;
  wire [15:0] sel_95054;
  wire [21:0] umul_95055;
  wire [15:0] add_95057;
  wire [15:0] sel_95062;
  wire [31:0] smod_95066;
  wire [31:0] smod_95071;
  wire [31:0] smod_95076;
  wire [31:0] smod_95081;
  wire [31:0] smod_95086;
  wire [31:0] smod_95091;
  wire [31:0] smod_95096;
  wire [31:0] smod_95101;
  wire [22:0] umul_95117;
  wire [20:0] add_95119;
  wire [15:0] sel_95124;
  wire [22:0] umul_95125;
  wire [20:0] add_95127;
  wire [15:0] sel_95132;
  wire [22:0] umul_95133;
  wire [22:0] add_95135;
  wire [15:0] sel_95140;
  wire [22:0] umul_95141;
  wire [22:0] add_95143;
  wire [15:0] sel_95148;
  wire [21:0] umul_95149;
  wire [20:0] add_95151;
  wire [15:0] sel_95156;
  wire [21:0] umul_95157;
  wire [20:0] add_95159;
  wire [15:0] sel_95164;
  wire [21:0] umul_95165;
  wire [21:0] add_95167;
  wire [15:0] sel_95172;
  wire [21:0] umul_95173;
  wire [21:0] add_95175;
  wire [15:0] sel_95180;
  wire [15:0] array_index_95181;
  wire [31:0] smod_95185;
  wire [15:0] array_index_95187;
  wire [31:0] smod_95191;
  wire [21:0] umul_95241;
  wire [15:0] add_95243;
  wire [15:0] sel_95248;
  wire [21:0] umul_95249;
  wire [15:0] add_95251;
  wire [15:0] sel_95256;
  wire [31:0] smod_95260;
  wire [31:0] smod_95265;
  wire [31:0] smod_95270;
  wire [31:0] smod_95275;
  wire [31:0] smod_95280;
  wire [31:0] smod_95285;
  wire [31:0] smod_95290;
  wire [31:0] smod_95295;
  wire [22:0] umul_95311;
  wire [20:0] add_95313;
  wire [15:0] sel_95318;
  wire [22:0] umul_95319;
  wire [20:0] add_95321;
  wire [15:0] sel_95326;
  wire [22:0] umul_95327;
  wire [22:0] add_95329;
  wire [15:0] sel_95334;
  wire [22:0] umul_95335;
  wire [22:0] add_95337;
  wire [15:0] sel_95342;
  wire [21:0] umul_95343;
  wire [20:0] add_95345;
  wire [15:0] sel_95350;
  wire [21:0] umul_95351;
  wire [20:0] add_95353;
  wire [15:0] sel_95358;
  wire [21:0] umul_95359;
  wire [21:0] add_95361;
  wire [15:0] sel_95366;
  wire [21:0] umul_95367;
  wire [21:0] add_95369;
  wire [15:0] sel_95374;
  wire [15:0] array_index_95375;
  wire [31:0] smod_95379;
  wire [15:0] array_index_95381;
  wire [31:0] smod_95385;
  wire [21:0] umul_95435;
  wire [15:0] add_95437;
  wire [15:0] sel_95442;
  wire [21:0] umul_95443;
  wire [15:0] add_95445;
  wire [15:0] sel_95450;
  wire [31:0] smod_95454;
  wire [31:0] smod_95459;
  wire [31:0] smod_95464;
  wire [31:0] smod_95469;
  wire [31:0] smod_95474;
  wire [31:0] smod_95479;
  wire [31:0] smod_95484;
  wire [31:0] smod_95489;
  wire [22:0] umul_95505;
  wire [20:0] add_95507;
  wire [15:0] sel_95512;
  wire [22:0] umul_95513;
  wire [20:0] add_95515;
  wire [15:0] sel_95520;
  wire [22:0] umul_95521;
  wire [22:0] add_95523;
  wire [15:0] sel_95528;
  wire [22:0] umul_95529;
  wire [22:0] add_95531;
  wire [15:0] sel_95536;
  wire [21:0] umul_95537;
  wire [20:0] add_95539;
  wire [15:0] sel_95544;
  wire [21:0] umul_95545;
  wire [20:0] add_95547;
  wire [15:0] sel_95552;
  wire [21:0] umul_95553;
  wire [21:0] add_95555;
  wire [15:0] sel_95560;
  wire [21:0] umul_95561;
  wire [21:0] add_95563;
  wire [15:0] sel_95568;
  wire [15:0] array_index_95569;
  wire [31:0] smod_95573;
  wire [15:0] array_index_95575;
  wire [31:0] smod_95579;
  wire [21:0] umul_95629;
  wire [15:0] add_95631;
  wire [15:0] sel_95636;
  wire [21:0] umul_95637;
  wire [15:0] add_95639;
  wire [15:0] sel_95644;
  wire [31:0] smod_95648;
  wire [31:0] smod_95653;
  wire [31:0] smod_95658;
  wire [31:0] smod_95663;
  wire [31:0] smod_95668;
  wire [31:0] smod_95673;
  wire [31:0] smod_95678;
  wire [31:0] smod_95683;
  wire [22:0] umul_95697;
  wire [20:0] add_95699;
  wire [15:0] sel_95704;
  wire [22:0] umul_95705;
  wire [20:0] add_95707;
  wire [15:0] sel_95712;
  wire [22:0] umul_95713;
  wire [22:0] add_95715;
  wire [15:0] sel_95720;
  wire [22:0] umul_95721;
  wire [22:0] add_95723;
  wire [15:0] sel_95728;
  wire [21:0] umul_95729;
  wire [20:0] add_95731;
  wire [15:0] sel_95736;
  wire [21:0] umul_95737;
  wire [20:0] add_95739;
  wire [15:0] sel_95744;
  wire [21:0] umul_95745;
  wire [21:0] add_95747;
  wire [15:0] sel_95752;
  wire [21:0] umul_95753;
  wire [21:0] add_95755;
  wire [15:0] sel_95760;
  wire [31:0] smod_95763;
  wire [31:0] smod_95767;
  wire [15:0] add_95818;
  wire [15:0] sel_95823;
  wire [15:0] add_95825;
  wire [15:0] sel_95830;
  wire [31:0] smod_95834;
  wire [31:0] smod_95839;
  wire [31:0] smod_95844;
  wire [31:0] smod_95849;
  wire [31:0] smod_95854;
  wire [31:0] smod_95859;
  wire [31:0] smod_95863;
  wire [31:0] smod_95867;
  wire [22:0] umul_95877;
  wire [20:0] add_95879;
  wire [15:0] sel_95884;
  wire [22:0] umul_95885;
  wire [20:0] add_95887;
  wire [15:0] sel_95892;
  wire [22:0] umul_95893;
  wire [22:0] add_95895;
  wire [15:0] sel_95900;
  wire [22:0] umul_95901;
  wire [22:0] add_95903;
  wire [15:0] sel_95908;
  wire [21:0] umul_95909;
  wire [20:0] add_95911;
  wire [15:0] sel_95916;
  wire [21:0] umul_95917;
  wire [20:0] add_95919;
  wire [15:0] sel_95924;
  wire [21:0] add_95926;
  wire [15:0] sel_95931;
  wire [21:0] add_95933;
  wire [15:0] sel_95938;
  wire [31:0] smod_95939;
  wire [31:0] smod_95941;
  wire [15:0] sel_95990;
  wire [15:0] sel_95994;
  wire [31:0] smod_95998;
  wire [31:0] smod_96003;
  wire [31:0] smod_96008;
  wire [31:0] smod_96013;
  wire [31:0] smod_96017;
  wire [31:0] smod_96021;
  wire [31:0] smod_96023;
  wire [31:0] smod_96025;
  wire [22:0] umul_96031;
  wire [20:0] add_96033;
  wire [15:0] sel_96038;
  wire [22:0] umul_96039;
  wire [20:0] add_96041;
  wire [15:0] sel_96046;
  wire [22:0] umul_96047;
  wire [22:0] add_96049;
  wire [15:0] sel_96054;
  wire [22:0] umul_96055;
  wire [22:0] add_96057;
  wire [15:0] sel_96062;
  wire [20:0] add_96064;
  wire [15:0] sel_96069;
  wire [20:0] add_96071;
  wire [15:0] sel_96076;
  wire [15:0] sel_96080;
  wire [15:0] sel_96084;
  wire [31:0] smod_96128;
  wire [31:0] smod_96133;
  wire [31:0] smod_96137;
  wire [31:0] smod_96141;
  wire [31:0] smod_96143;
  wire [31:0] smod_96145;
  wire [22:0] umul_96151;
  wire [20:0] add_96153;
  wire [15:0] sel_96158;
  wire [22:0] umul_96159;
  wire [20:0] add_96161;
  wire [15:0] sel_96166;
  wire [22:0] add_96168;
  wire [15:0] sel_96173;
  wire [22:0] add_96175;
  wire [15:0] sel_96180;
  wire [15:0] sel_96184;
  wire [15:0] sel_96188;
  wire [1:0] concat_96191;
  wire [1:0] add_96218;
  wire [31:0] smod_96221;
  wire [31:0] smod_96225;
  wire [31:0] smod_96227;
  wire [31:0] smod_96229;
  wire [20:0] add_96236;
  wire [15:0] sel_96241;
  wire [20:0] add_96243;
  wire [15:0] sel_96248;
  wire [15:0] sel_96252;
  wire [15:0] sel_96256;
  wire [2:0] concat_96259;
  wire [2:0] add_96274;
  wire [31:0] smod_96275;
  wire [31:0] smod_96277;
  wire [15:0] sel_96286;
  wire [15:0] sel_96290;
  wire [3:0] concat_96293;
  wire [3:0] add_96300;
  wire [4:0] concat_96307;
  wire [4:0] add_96310;
  assign array_index_86589 = set1_unflattened[6'h00];
  assign array_index_86591 = set2_unflattened[6'h00];
  assign umul_86593 = umul22b_16b_x_6b(array_index_86589, 6'h35);
  assign umul_86594 = umul22b_16b_x_6b(array_index_86591, 6'h35);
  assign umul_86603 = umul22b_16b_x_6b(array_index_86589, 6'h3b);
  assign umul_86604 = umul22b_16b_x_6b(array_index_86591, 6'h3b);
  assign array_index_86605 = set1_unflattened[6'h01];
  assign array_index_86609 = set2_unflattened[6'h01];
  assign umul_86617 = umul22b_16b_x_6b(array_index_86605, 6'h35);
  assign add_86619 = {1'h0, umul_86593[21:7]} + 16'h007d;
  assign umul_86621 = umul22b_16b_x_6b(array_index_86609, 6'h35);
  assign add_86623 = {1'h0, umul_86594[21:7]} + 16'h007d;
  assign umul_86643 = umul22b_16b_x_6b(array_index_86589, 6'h3d);
  assign umul_86644 = umul22b_16b_x_6b(array_index_86591, 6'h3d);
  assign umul_86645 = umul22b_16b_x_6b(array_index_86605, 6'h3b);
  assign add_86647 = {1'h0, umul_86603[21:1]} + 22'h00_1f59;
  assign umul_86649 = umul22b_16b_x_6b(array_index_86609, 6'h3b);
  assign add_86651 = {1'h0, umul_86604[21:1]} + 22'h00_1f59;
  assign array_index_86653 = set1_unflattened[6'h02];
  assign smod_86657 = $unsigned($signed({9'h000, add_86619, umul_86593[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_86658 = set2_unflattened[6'h02];
  assign smod_86662 = $unsigned($signed({9'h000, add_86623, umul_86594[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_86675 = umul22b_16b_x_6b(array_index_86653, 6'h35);
  assign add_86677 = {1'h0, umul_86617[21:7]} + 16'h007d;
  assign umul_86681 = umul22b_16b_x_6b(array_index_86658, 6'h35);
  assign add_86683 = {1'h0, umul_86621[21:7]} + 16'h007d;
  assign smod_86698 = $unsigned($signed({9'h000, add_86647, umul_86603[0]}) % $signed(32'h0000_3ffd));
  assign smod_86702 = $unsigned($signed({9'h000, add_86651, umul_86604[0]}) % $signed(32'h0000_3ffd));
  assign umul_86717 = umul23b_16b_x_7b(array_index_86589, 7'h47);
  assign umul_86718 = umul23b_16b_x_7b(array_index_86591, 7'h47);
  assign umul_86719 = umul22b_16b_x_6b(array_index_86605, 6'h3d);
  assign add_86721 = {1'h0, umul_86643[21:2]} + 21'h00_0fb9;
  assign umul_86723 = umul22b_16b_x_6b(array_index_86609, 6'h3d);
  assign add_86725 = {1'h0, umul_86644[21:2]} + 21'h00_0fb9;
  assign umul_86727 = umul22b_16b_x_6b(array_index_86653, 6'h3b);
  assign add_86729 = {1'h0, umul_86645[21:1]} + 22'h00_1f59;
  assign umul_86733 = umul22b_16b_x_6b(array_index_86658, 6'h3b);
  assign add_86735 = {1'h0, umul_86649[21:1]} + 22'h00_1f59;
  assign array_index_86739 = set1_unflattened[6'h03];
  assign smod_86743 = $unsigned($signed({9'h000, add_86677, umul_86617[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_86746 = set2_unflattened[6'h03];
  assign smod_86750 = $unsigned($signed({9'h000, add_86683, umul_86621[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_86777 = umul22b_16b_x_6b(array_index_86739, 6'h35);
  assign add_86779 = {1'h0, umul_86675[21:7]} + 16'h007d;
  assign sel_86784 = $signed({1'h0, smod_86657[15:0]}) < $signed(17'h0_3ffd) ? smod_86657[15:0] : 16'h3ffd;
  assign umul_86785 = umul22b_16b_x_6b(array_index_86746, 6'h35);
  assign add_86787 = {1'h0, umul_86681[21:7]} + 16'h007d;
  assign sel_86792 = $signed({1'h0, smod_86662[15:0]}) < $signed(17'h0_3ffd) ? smod_86662[15:0] : 16'h3ffd;
  assign smod_86804 = $unsigned($signed({9'h000, add_86721, umul_86643[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_86808 = $unsigned($signed({9'h000, add_86725, umul_86644[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_86812 = $unsigned($signed({9'h000, add_86729, umul_86645[0]}) % $signed(32'h0000_3ffd));
  assign smod_86818 = $unsigned($signed({9'h000, add_86735, umul_86649[0]}) % $signed(32'h0000_3ffd));
  assign umul_86835 = umul23b_16b_x_7b(array_index_86589, 7'h49);
  assign umul_86836 = umul23b_16b_x_7b(array_index_86591, 7'h49);
  assign umul_86837 = umul23b_16b_x_7b(array_index_86605, 7'h47);
  assign add_86839 = {1'h0, umul_86717[22:1]} + 23'h00_1f8b;
  assign umul_86841 = umul23b_16b_x_7b(array_index_86609, 7'h47);
  assign add_86843 = {1'h0, umul_86718[22:1]} + 23'h00_1f8b;
  assign umul_86845 = umul22b_16b_x_6b(array_index_86653, 6'h3d);
  assign add_86847 = {1'h0, umul_86719[21:2]} + 21'h00_0fb9;
  assign umul_86851 = umul22b_16b_x_6b(array_index_86658, 6'h3d);
  assign add_86853 = {1'h0, umul_86723[21:2]} + 21'h00_0fb9;
  assign umul_86857 = umul22b_16b_x_6b(array_index_86739, 6'h3b);
  assign add_86859 = {1'h0, umul_86727[21:1]} + 22'h00_1f59;
  assign sel_86864 = $signed({1'h0, smod_86698[15:0]}) < $signed(17'h0_3ffd) ? smod_86698[15:0] : 16'h3ffd;
  assign umul_86865 = umul22b_16b_x_6b(array_index_86746, 6'h3b);
  assign add_86867 = {1'h0, umul_86733[21:1]} + 22'h00_1f59;
  assign sel_86872 = $signed({1'h0, smod_86702[15:0]}) < $signed(17'h0_3ffd) ? smod_86702[15:0] : 16'h3ffd;
  assign array_index_86873 = set1_unflattened[6'h04];
  assign smod_86877 = $unsigned($signed({9'h000, add_86779, umul_86675[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_86879 = set2_unflattened[6'h04];
  assign smod_86883 = $unsigned($signed({9'h000, add_86787, umul_86681[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_86921 = umul22b_16b_x_6b(array_index_86873, 6'h35);
  assign add_86923 = {1'h0, umul_86777[21:7]} + 16'h007d;
  assign sel_86928 = $signed({1'h0, smod_86743[15:0]}) < $signed({1'h0, sel_86784}) ? smod_86743[15:0] : sel_86784;
  assign umul_86929 = umul22b_16b_x_6b(array_index_86879, 6'h35);
  assign add_86931 = {1'h0, umul_86785[21:7]} + 16'h007d;
  assign sel_86936 = $signed({1'h0, smod_86750[15:0]}) < $signed({1'h0, sel_86792}) ? smod_86750[15:0] : sel_86792;
  assign smod_86946 = $unsigned($signed({8'h00, add_86839, umul_86717[0]}) % $signed(32'h0000_3ffd));
  assign smod_86950 = $unsigned($signed({8'h00, add_86843, umul_86718[0]}) % $signed(32'h0000_3ffd));
  assign smod_86954 = $unsigned($signed({9'h000, add_86847, umul_86719[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_86960 = $unsigned($signed({9'h000, add_86853, umul_86723[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_86966 = $unsigned($signed({9'h000, add_86859, umul_86727[0]}) % $signed(32'h0000_3ffd));
  assign smod_86971 = $unsigned($signed({9'h000, add_86867, umul_86733[0]}) % $signed(32'h0000_3ffd));
  assign umul_86987 = umul23b_16b_x_7b(array_index_86605, 7'h49);
  assign add_86989 = {1'h0, umul_86835[22:3]} + 21'h00_07e9;
  assign umul_86991 = umul23b_16b_x_7b(array_index_86609, 7'h49);
  assign add_86993 = {1'h0, umul_86836[22:3]} + 21'h00_07e9;
  assign umul_86995 = umul23b_16b_x_7b(array_index_86653, 7'h47);
  assign add_86997 = {1'h0, umul_86837[22:1]} + 23'h00_1f8b;
  assign umul_87001 = umul23b_16b_x_7b(array_index_86658, 7'h47);
  assign add_87003 = {1'h0, umul_86841[22:1]} + 23'h00_1f8b;
  assign umul_87007 = umul22b_16b_x_6b(array_index_86739, 6'h3d);
  assign add_87009 = {1'h0, umul_86845[21:2]} + 21'h00_0fb9;
  assign sel_87014 = $signed({1'h0, smod_86804[15:0]}) < $signed(17'h0_3ffd) ? smod_86804[15:0] : 16'h3ffd;
  assign umul_87015 = umul22b_16b_x_6b(array_index_86746, 6'h3d);
  assign add_87017 = {1'h0, umul_86851[21:2]} + 21'h00_0fb9;
  assign sel_87022 = $signed({1'h0, smod_86808[15:0]}) < $signed(17'h0_3ffd) ? smod_86808[15:0] : 16'h3ffd;
  assign umul_87023 = umul22b_16b_x_6b(array_index_86873, 6'h3b);
  assign add_87025 = {1'h0, umul_86857[21:1]} + 22'h00_1f59;
  assign sel_87030 = $signed({1'h0, smod_86812[15:0]}) < $signed({1'h0, sel_86864}) ? smod_86812[15:0] : sel_86864;
  assign umul_87031 = umul22b_16b_x_6b(array_index_86879, 6'h3b);
  assign add_87033 = {1'h0, umul_86865[21:1]} + 22'h00_1f59;
  assign sel_87038 = $signed({1'h0, smod_86818[15:0]}) < $signed({1'h0, sel_86872}) ? smod_86818[15:0] : sel_86872;
  assign array_index_87039 = set1_unflattened[6'h05];
  assign smod_87043 = $unsigned($signed({9'h000, add_86923, umul_86777[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_87045 = set2_unflattened[6'h05];
  assign smod_87049 = $unsigned($signed({9'h000, add_86931, umul_86785[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_87095 = umul22b_16b_x_6b(array_index_87039, 6'h35);
  assign add_87097 = {1'h0, umul_86921[21:7]} + 16'h007d;
  assign sel_87102 = $signed({1'h0, smod_86877[15:0]}) < $signed({1'h0, sel_86928}) ? smod_86877[15:0] : sel_86928;
  assign umul_87103 = umul22b_16b_x_6b(array_index_87045, 6'h35);
  assign add_87105 = {1'h0, umul_86929[21:7]} + 16'h007d;
  assign sel_87110 = $signed({1'h0, smod_86883[15:0]}) < $signed({1'h0, sel_86936}) ? smod_86883[15:0] : sel_86936;
  assign smod_87114 = $unsigned($signed({8'h00, add_86989, umul_86835[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_87118 = $unsigned($signed({8'h00, add_86993, umul_86836[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_87122 = $unsigned($signed({8'h00, add_86997, umul_86837[0]}) % $signed(32'h0000_3ffd));
  assign smod_87128 = $unsigned($signed({8'h00, add_87003, umul_86841[0]}) % $signed(32'h0000_3ffd));
  assign smod_87134 = $unsigned($signed({9'h000, add_87009, umul_86845[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_87139 = $unsigned($signed({9'h000, add_87017, umul_86851[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_87144 = $unsigned($signed({9'h000, add_87025, umul_86857[0]}) % $signed(32'h0000_3ffd));
  assign smod_87149 = $unsigned($signed({9'h000, add_87033, umul_86865[0]}) % $signed(32'h0000_3ffd));
  assign umul_87165 = umul23b_16b_x_7b(array_index_86653, 7'h49);
  assign add_87167 = {1'h0, umul_86987[22:3]} + 21'h00_07e9;
  assign umul_87171 = umul23b_16b_x_7b(array_index_86658, 7'h49);
  assign add_87173 = {1'h0, umul_86991[22:3]} + 21'h00_07e9;
  assign umul_87177 = umul23b_16b_x_7b(array_index_86739, 7'h47);
  assign add_87179 = {1'h0, umul_86995[22:1]} + 23'h00_1f8b;
  assign sel_87184 = $signed({1'h0, smod_86946[15:0]}) < $signed(17'h0_3ffd) ? smod_86946[15:0] : 16'h3ffd;
  assign umul_87185 = umul23b_16b_x_7b(array_index_86746, 7'h47);
  assign add_87187 = {1'h0, umul_87001[22:1]} + 23'h00_1f8b;
  assign sel_87192 = $signed({1'h0, smod_86950[15:0]}) < $signed(17'h0_3ffd) ? smod_86950[15:0] : 16'h3ffd;
  assign umul_87193 = umul22b_16b_x_6b(array_index_86873, 6'h3d);
  assign add_87195 = {1'h0, umul_87007[21:2]} + 21'h00_0fb9;
  assign sel_87200 = $signed({1'h0, smod_86954[15:0]}) < $signed({1'h0, sel_87014}) ? smod_86954[15:0] : sel_87014;
  assign umul_87201 = umul22b_16b_x_6b(array_index_86879, 6'h3d);
  assign add_87203 = {1'h0, umul_87015[21:2]} + 21'h00_0fb9;
  assign sel_87208 = $signed({1'h0, smod_86960[15:0]}) < $signed({1'h0, sel_87022}) ? smod_86960[15:0] : sel_87022;
  assign umul_87209 = umul22b_16b_x_6b(array_index_87039, 6'h3b);
  assign add_87211 = {1'h0, umul_87023[21:1]} + 22'h00_1f59;
  assign sel_87216 = $signed({1'h0, smod_86966[15:0]}) < $signed({1'h0, sel_87030}) ? smod_86966[15:0] : sel_87030;
  assign umul_87217 = umul22b_16b_x_6b(array_index_87045, 6'h3b);
  assign add_87219 = {1'h0, umul_87031[21:1]} + 22'h00_1f59;
  assign sel_87224 = $signed({1'h0, smod_86971[15:0]}) < $signed({1'h0, sel_87038}) ? smod_86971[15:0] : sel_87038;
  assign array_index_87225 = set1_unflattened[6'h06];
  assign smod_87229 = $unsigned($signed({9'h000, add_87097, umul_86921[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_87231 = set2_unflattened[6'h06];
  assign smod_87235 = $unsigned($signed({9'h000, add_87105, umul_86929[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_87285 = umul22b_16b_x_6b(array_index_87225, 6'h35);
  assign add_87287 = {1'h0, umul_87095[21:7]} + 16'h007d;
  assign sel_87292 = $signed({1'h0, smod_87043[15:0]}) < $signed({1'h0, sel_87102}) ? smod_87043[15:0] : sel_87102;
  assign umul_87293 = umul22b_16b_x_6b(array_index_87231, 6'h35);
  assign add_87295 = {1'h0, umul_87103[21:7]} + 16'h007d;
  assign sel_87300 = $signed({1'h0, smod_87049[15:0]}) < $signed({1'h0, sel_87110}) ? smod_87049[15:0] : sel_87110;
  assign smod_87304 = $unsigned($signed({8'h00, add_87167, umul_86987[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_87310 = $unsigned($signed({8'h00, add_87173, umul_86991[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_87316 = $unsigned($signed({8'h00, add_87179, umul_86995[0]}) % $signed(32'h0000_3ffd));
  assign smod_87321 = $unsigned($signed({8'h00, add_87187, umul_87001[0]}) % $signed(32'h0000_3ffd));
  assign smod_87326 = $unsigned($signed({9'h000, add_87195, umul_87007[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_87331 = $unsigned($signed({9'h000, add_87203, umul_87015[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_87336 = $unsigned($signed({9'h000, add_87211, umul_87023[0]}) % $signed(32'h0000_3ffd));
  assign smod_87341 = $unsigned($signed({9'h000, add_87219, umul_87031[0]}) % $signed(32'h0000_3ffd));
  assign umul_87357 = umul23b_16b_x_7b(array_index_86739, 7'h49);
  assign add_87359 = {1'h0, umul_87165[22:3]} + 21'h00_07e9;
  assign sel_87364 = $signed({1'h0, smod_87114[15:0]}) < $signed(17'h0_3ffd) ? smod_87114[15:0] : 16'h3ffd;
  assign umul_87365 = umul23b_16b_x_7b(array_index_86746, 7'h49);
  assign add_87367 = {1'h0, umul_87171[22:3]} + 21'h00_07e9;
  assign sel_87372 = $signed({1'h0, smod_87118[15:0]}) < $signed(17'h0_3ffd) ? smod_87118[15:0] : 16'h3ffd;
  assign umul_87373 = umul23b_16b_x_7b(array_index_86873, 7'h47);
  assign add_87375 = {1'h0, umul_87177[22:1]} + 23'h00_1f8b;
  assign sel_87380 = $signed({1'h0, smod_87122[15:0]}) < $signed({1'h0, sel_87184}) ? smod_87122[15:0] : sel_87184;
  assign umul_87381 = umul23b_16b_x_7b(array_index_86879, 7'h47);
  assign add_87383 = {1'h0, umul_87185[22:1]} + 23'h00_1f8b;
  assign sel_87388 = $signed({1'h0, smod_87128[15:0]}) < $signed({1'h0, sel_87192}) ? smod_87128[15:0] : sel_87192;
  assign umul_87389 = umul22b_16b_x_6b(array_index_87039, 6'h3d);
  assign add_87391 = {1'h0, umul_87193[21:2]} + 21'h00_0fb9;
  assign sel_87396 = $signed({1'h0, smod_87134[15:0]}) < $signed({1'h0, sel_87200}) ? smod_87134[15:0] : sel_87200;
  assign umul_87397 = umul22b_16b_x_6b(array_index_87045, 6'h3d);
  assign add_87399 = {1'h0, umul_87201[21:2]} + 21'h00_0fb9;
  assign sel_87404 = $signed({1'h0, smod_87139[15:0]}) < $signed({1'h0, sel_87208}) ? smod_87139[15:0] : sel_87208;
  assign umul_87405 = umul22b_16b_x_6b(array_index_87225, 6'h3b);
  assign add_87407 = {1'h0, umul_87209[21:1]} + 22'h00_1f59;
  assign sel_87412 = $signed({1'h0, smod_87144[15:0]}) < $signed({1'h0, sel_87216}) ? smod_87144[15:0] : sel_87216;
  assign umul_87413 = umul22b_16b_x_6b(array_index_87231, 6'h3b);
  assign add_87415 = {1'h0, umul_87217[21:1]} + 22'h00_1f59;
  assign sel_87420 = $signed({1'h0, smod_87149[15:0]}) < $signed({1'h0, sel_87224}) ? smod_87149[15:0] : sel_87224;
  assign array_index_87421 = set1_unflattened[6'h07];
  assign smod_87425 = $unsigned($signed({9'h000, add_87287, umul_87095[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_87427 = set2_unflattened[6'h07];
  assign smod_87431 = $unsigned($signed({9'h000, add_87295, umul_87103[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_87481 = umul22b_16b_x_6b(array_index_87421, 6'h35);
  assign add_87483 = {1'h0, umul_87285[21:7]} + 16'h007d;
  assign sel_87488 = $signed({1'h0, smod_87229[15:0]}) < $signed({1'h0, sel_87292}) ? smod_87229[15:0] : sel_87292;
  assign umul_87489 = umul22b_16b_x_6b(array_index_87427, 6'h35);
  assign add_87491 = {1'h0, umul_87293[21:7]} + 16'h007d;
  assign sel_87496 = $signed({1'h0, smod_87235[15:0]}) < $signed({1'h0, sel_87300}) ? smod_87235[15:0] : sel_87300;
  assign smod_87500 = $unsigned($signed({8'h00, add_87359, umul_87165[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_87505 = $unsigned($signed({8'h00, add_87367, umul_87171[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_87510 = $unsigned($signed({8'h00, add_87375, umul_87177[0]}) % $signed(32'h0000_3ffd));
  assign smod_87515 = $unsigned($signed({8'h00, add_87383, umul_87185[0]}) % $signed(32'h0000_3ffd));
  assign smod_87520 = $unsigned($signed({9'h000, add_87391, umul_87193[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_87525 = $unsigned($signed({9'h000, add_87399, umul_87201[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_87530 = $unsigned($signed({9'h000, add_87407, umul_87209[0]}) % $signed(32'h0000_3ffd));
  assign smod_87535 = $unsigned($signed({9'h000, add_87415, umul_87217[0]}) % $signed(32'h0000_3ffd));
  assign umul_87551 = umul23b_16b_x_7b(array_index_86873, 7'h49);
  assign add_87553 = {1'h0, umul_87357[22:3]} + 21'h00_07e9;
  assign sel_87558 = $signed({1'h0, smod_87304[15:0]}) < $signed({1'h0, sel_87364}) ? smod_87304[15:0] : sel_87364;
  assign umul_87559 = umul23b_16b_x_7b(array_index_86879, 7'h49);
  assign add_87561 = {1'h0, umul_87365[22:3]} + 21'h00_07e9;
  assign sel_87566 = $signed({1'h0, smod_87310[15:0]}) < $signed({1'h0, sel_87372}) ? smod_87310[15:0] : sel_87372;
  assign umul_87567 = umul23b_16b_x_7b(array_index_87039, 7'h47);
  assign add_87569 = {1'h0, umul_87373[22:1]} + 23'h00_1f8b;
  assign sel_87574 = $signed({1'h0, smod_87316[15:0]}) < $signed({1'h0, sel_87380}) ? smod_87316[15:0] : sel_87380;
  assign umul_87575 = umul23b_16b_x_7b(array_index_87045, 7'h47);
  assign add_87577 = {1'h0, umul_87381[22:1]} + 23'h00_1f8b;
  assign sel_87582 = $signed({1'h0, smod_87321[15:0]}) < $signed({1'h0, sel_87388}) ? smod_87321[15:0] : sel_87388;
  assign umul_87583 = umul22b_16b_x_6b(array_index_87225, 6'h3d);
  assign add_87585 = {1'h0, umul_87389[21:2]} + 21'h00_0fb9;
  assign sel_87590 = $signed({1'h0, smod_87326[15:0]}) < $signed({1'h0, sel_87396}) ? smod_87326[15:0] : sel_87396;
  assign umul_87591 = umul22b_16b_x_6b(array_index_87231, 6'h3d);
  assign add_87593 = {1'h0, umul_87397[21:2]} + 21'h00_0fb9;
  assign sel_87598 = $signed({1'h0, smod_87331[15:0]}) < $signed({1'h0, sel_87404}) ? smod_87331[15:0] : sel_87404;
  assign umul_87599 = umul22b_16b_x_6b(array_index_87421, 6'h3b);
  assign add_87601 = {1'h0, umul_87405[21:1]} + 22'h00_1f59;
  assign sel_87606 = $signed({1'h0, smod_87336[15:0]}) < $signed({1'h0, sel_87412}) ? smod_87336[15:0] : sel_87412;
  assign umul_87607 = umul22b_16b_x_6b(array_index_87427, 6'h3b);
  assign add_87609 = {1'h0, umul_87413[21:1]} + 22'h00_1f59;
  assign sel_87614 = $signed({1'h0, smod_87341[15:0]}) < $signed({1'h0, sel_87420}) ? smod_87341[15:0] : sel_87420;
  assign array_index_87615 = set1_unflattened[6'h08];
  assign smod_87619 = $unsigned($signed({9'h000, add_87483, umul_87285[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_87621 = set2_unflattened[6'h08];
  assign smod_87625 = $unsigned($signed({9'h000, add_87491, umul_87293[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_87675 = umul22b_16b_x_6b(array_index_87615, 6'h35);
  assign add_87677 = {1'h0, umul_87481[21:7]} + 16'h007d;
  assign sel_87682 = $signed({1'h0, smod_87425[15:0]}) < $signed({1'h0, sel_87488}) ? smod_87425[15:0] : sel_87488;
  assign umul_87683 = umul22b_16b_x_6b(array_index_87621, 6'h35);
  assign add_87685 = {1'h0, umul_87489[21:7]} + 16'h007d;
  assign sel_87690 = $signed({1'h0, smod_87431[15:0]}) < $signed({1'h0, sel_87496}) ? smod_87431[15:0] : sel_87496;
  assign smod_87694 = $unsigned($signed({8'h00, add_87553, umul_87357[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_87699 = $unsigned($signed({8'h00, add_87561, umul_87365[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_87704 = $unsigned($signed({8'h00, add_87569, umul_87373[0]}) % $signed(32'h0000_3ffd));
  assign smod_87709 = $unsigned($signed({8'h00, add_87577, umul_87381[0]}) % $signed(32'h0000_3ffd));
  assign smod_87714 = $unsigned($signed({9'h000, add_87585, umul_87389[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_87719 = $unsigned($signed({9'h000, add_87593, umul_87397[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_87724 = $unsigned($signed({9'h000, add_87601, umul_87405[0]}) % $signed(32'h0000_3ffd));
  assign smod_87729 = $unsigned($signed({9'h000, add_87609, umul_87413[0]}) % $signed(32'h0000_3ffd));
  assign umul_87745 = umul23b_16b_x_7b(array_index_87039, 7'h49);
  assign add_87747 = {1'h0, umul_87551[22:3]} + 21'h00_07e9;
  assign sel_87752 = $signed({1'h0, smod_87500[15:0]}) < $signed({1'h0, sel_87558}) ? smod_87500[15:0] : sel_87558;
  assign umul_87753 = umul23b_16b_x_7b(array_index_87045, 7'h49);
  assign add_87755 = {1'h0, umul_87559[22:3]} + 21'h00_07e9;
  assign sel_87760 = $signed({1'h0, smod_87505[15:0]}) < $signed({1'h0, sel_87566}) ? smod_87505[15:0] : sel_87566;
  assign umul_87761 = umul23b_16b_x_7b(array_index_87225, 7'h47);
  assign add_87763 = {1'h0, umul_87567[22:1]} + 23'h00_1f8b;
  assign sel_87768 = $signed({1'h0, smod_87510[15:0]}) < $signed({1'h0, sel_87574}) ? smod_87510[15:0] : sel_87574;
  assign umul_87769 = umul23b_16b_x_7b(array_index_87231, 7'h47);
  assign add_87771 = {1'h0, umul_87575[22:1]} + 23'h00_1f8b;
  assign sel_87776 = $signed({1'h0, smod_87515[15:0]}) < $signed({1'h0, sel_87582}) ? smod_87515[15:0] : sel_87582;
  assign umul_87777 = umul22b_16b_x_6b(array_index_87421, 6'h3d);
  assign add_87779 = {1'h0, umul_87583[21:2]} + 21'h00_0fb9;
  assign sel_87784 = $signed({1'h0, smod_87520[15:0]}) < $signed({1'h0, sel_87590}) ? smod_87520[15:0] : sel_87590;
  assign umul_87785 = umul22b_16b_x_6b(array_index_87427, 6'h3d);
  assign add_87787 = {1'h0, umul_87591[21:2]} + 21'h00_0fb9;
  assign sel_87792 = $signed({1'h0, smod_87525[15:0]}) < $signed({1'h0, sel_87598}) ? smod_87525[15:0] : sel_87598;
  assign umul_87793 = umul22b_16b_x_6b(array_index_87615, 6'h3b);
  assign add_87795 = {1'h0, umul_87599[21:1]} + 22'h00_1f59;
  assign sel_87800 = $signed({1'h0, smod_87530[15:0]}) < $signed({1'h0, sel_87606}) ? smod_87530[15:0] : sel_87606;
  assign umul_87801 = umul22b_16b_x_6b(array_index_87621, 6'h3b);
  assign add_87803 = {1'h0, umul_87607[21:1]} + 22'h00_1f59;
  assign sel_87808 = $signed({1'h0, smod_87535[15:0]}) < $signed({1'h0, sel_87614}) ? smod_87535[15:0] : sel_87614;
  assign array_index_87809 = set1_unflattened[6'h09];
  assign smod_87813 = $unsigned($signed({9'h000, add_87677, umul_87481[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_87815 = set2_unflattened[6'h09];
  assign smod_87819 = $unsigned($signed({9'h000, add_87685, umul_87489[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_87869 = umul22b_16b_x_6b(array_index_87809, 6'h35);
  assign add_87871 = {1'h0, umul_87675[21:7]} + 16'h007d;
  assign sel_87876 = $signed({1'h0, smod_87619[15:0]}) < $signed({1'h0, sel_87682}) ? smod_87619[15:0] : sel_87682;
  assign umul_87877 = umul22b_16b_x_6b(array_index_87815, 6'h35);
  assign add_87879 = {1'h0, umul_87683[21:7]} + 16'h007d;
  assign sel_87884 = $signed({1'h0, smod_87625[15:0]}) < $signed({1'h0, sel_87690}) ? smod_87625[15:0] : sel_87690;
  assign smod_87888 = $unsigned($signed({8'h00, add_87747, umul_87551[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_87893 = $unsigned($signed({8'h00, add_87755, umul_87559[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_87898 = $unsigned($signed({8'h00, add_87763, umul_87567[0]}) % $signed(32'h0000_3ffd));
  assign smod_87903 = $unsigned($signed({8'h00, add_87771, umul_87575[0]}) % $signed(32'h0000_3ffd));
  assign smod_87908 = $unsigned($signed({9'h000, add_87779, umul_87583[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_87913 = $unsigned($signed({9'h000, add_87787, umul_87591[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_87918 = $unsigned($signed({9'h000, add_87795, umul_87599[0]}) % $signed(32'h0000_3ffd));
  assign smod_87923 = $unsigned($signed({9'h000, add_87803, umul_87607[0]}) % $signed(32'h0000_3ffd));
  assign umul_87939 = umul23b_16b_x_7b(array_index_87225, 7'h49);
  assign add_87941 = {1'h0, umul_87745[22:3]} + 21'h00_07e9;
  assign sel_87946 = $signed({1'h0, smod_87694[15:0]}) < $signed({1'h0, sel_87752}) ? smod_87694[15:0] : sel_87752;
  assign umul_87947 = umul23b_16b_x_7b(array_index_87231, 7'h49);
  assign add_87949 = {1'h0, umul_87753[22:3]} + 21'h00_07e9;
  assign sel_87954 = $signed({1'h0, smod_87699[15:0]}) < $signed({1'h0, sel_87760}) ? smod_87699[15:0] : sel_87760;
  assign umul_87955 = umul23b_16b_x_7b(array_index_87421, 7'h47);
  assign add_87957 = {1'h0, umul_87761[22:1]} + 23'h00_1f8b;
  assign sel_87962 = $signed({1'h0, smod_87704[15:0]}) < $signed({1'h0, sel_87768}) ? smod_87704[15:0] : sel_87768;
  assign umul_87963 = umul23b_16b_x_7b(array_index_87427, 7'h47);
  assign add_87965 = {1'h0, umul_87769[22:1]} + 23'h00_1f8b;
  assign sel_87970 = $signed({1'h0, smod_87709[15:0]}) < $signed({1'h0, sel_87776}) ? smod_87709[15:0] : sel_87776;
  assign umul_87971 = umul22b_16b_x_6b(array_index_87615, 6'h3d);
  assign add_87973 = {1'h0, umul_87777[21:2]} + 21'h00_0fb9;
  assign sel_87978 = $signed({1'h0, smod_87714[15:0]}) < $signed({1'h0, sel_87784}) ? smod_87714[15:0] : sel_87784;
  assign umul_87979 = umul22b_16b_x_6b(array_index_87621, 6'h3d);
  assign add_87981 = {1'h0, umul_87785[21:2]} + 21'h00_0fb9;
  assign sel_87986 = $signed({1'h0, smod_87719[15:0]}) < $signed({1'h0, sel_87792}) ? smod_87719[15:0] : sel_87792;
  assign umul_87987 = umul22b_16b_x_6b(array_index_87809, 6'h3b);
  assign add_87989 = {1'h0, umul_87793[21:1]} + 22'h00_1f59;
  assign sel_87994 = $signed({1'h0, smod_87724[15:0]}) < $signed({1'h0, sel_87800}) ? smod_87724[15:0] : sel_87800;
  assign umul_87995 = umul22b_16b_x_6b(array_index_87815, 6'h3b);
  assign add_87997 = {1'h0, umul_87801[21:1]} + 22'h00_1f59;
  assign sel_88002 = $signed({1'h0, smod_87729[15:0]}) < $signed({1'h0, sel_87808}) ? smod_87729[15:0] : sel_87808;
  assign array_index_88003 = set1_unflattened[6'h0a];
  assign smod_88007 = $unsigned($signed({9'h000, add_87871, umul_87675[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_88009 = set2_unflattened[6'h0a];
  assign smod_88013 = $unsigned($signed({9'h000, add_87879, umul_87683[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_88063 = umul22b_16b_x_6b(array_index_88003, 6'h35);
  assign add_88065 = {1'h0, umul_87869[21:7]} + 16'h007d;
  assign sel_88070 = $signed({1'h0, smod_87813[15:0]}) < $signed({1'h0, sel_87876}) ? smod_87813[15:0] : sel_87876;
  assign umul_88071 = umul22b_16b_x_6b(array_index_88009, 6'h35);
  assign add_88073 = {1'h0, umul_87877[21:7]} + 16'h007d;
  assign sel_88078 = $signed({1'h0, smod_87819[15:0]}) < $signed({1'h0, sel_87884}) ? smod_87819[15:0] : sel_87884;
  assign smod_88082 = $unsigned($signed({8'h00, add_87941, umul_87745[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_88087 = $unsigned($signed({8'h00, add_87949, umul_87753[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_88092 = $unsigned($signed({8'h00, add_87957, umul_87761[0]}) % $signed(32'h0000_3ffd));
  assign smod_88097 = $unsigned($signed({8'h00, add_87965, umul_87769[0]}) % $signed(32'h0000_3ffd));
  assign smod_88102 = $unsigned($signed({9'h000, add_87973, umul_87777[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_88107 = $unsigned($signed({9'h000, add_87981, umul_87785[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_88112 = $unsigned($signed({9'h000, add_87989, umul_87793[0]}) % $signed(32'h0000_3ffd));
  assign smod_88117 = $unsigned($signed({9'h000, add_87997, umul_87801[0]}) % $signed(32'h0000_3ffd));
  assign umul_88133 = umul23b_16b_x_7b(array_index_87421, 7'h49);
  assign add_88135 = {1'h0, umul_87939[22:3]} + 21'h00_07e9;
  assign sel_88140 = $signed({1'h0, smod_87888[15:0]}) < $signed({1'h0, sel_87946}) ? smod_87888[15:0] : sel_87946;
  assign umul_88141 = umul23b_16b_x_7b(array_index_87427, 7'h49);
  assign add_88143 = {1'h0, umul_87947[22:3]} + 21'h00_07e9;
  assign sel_88148 = $signed({1'h0, smod_87893[15:0]}) < $signed({1'h0, sel_87954}) ? smod_87893[15:0] : sel_87954;
  assign umul_88149 = umul23b_16b_x_7b(array_index_87615, 7'h47);
  assign add_88151 = {1'h0, umul_87955[22:1]} + 23'h00_1f8b;
  assign sel_88156 = $signed({1'h0, smod_87898[15:0]}) < $signed({1'h0, sel_87962}) ? smod_87898[15:0] : sel_87962;
  assign umul_88157 = umul23b_16b_x_7b(array_index_87621, 7'h47);
  assign add_88159 = {1'h0, umul_87963[22:1]} + 23'h00_1f8b;
  assign sel_88164 = $signed({1'h0, smod_87903[15:0]}) < $signed({1'h0, sel_87970}) ? smod_87903[15:0] : sel_87970;
  assign umul_88165 = umul22b_16b_x_6b(array_index_87809, 6'h3d);
  assign add_88167 = {1'h0, umul_87971[21:2]} + 21'h00_0fb9;
  assign sel_88172 = $signed({1'h0, smod_87908[15:0]}) < $signed({1'h0, sel_87978}) ? smod_87908[15:0] : sel_87978;
  assign umul_88173 = umul22b_16b_x_6b(array_index_87815, 6'h3d);
  assign add_88175 = {1'h0, umul_87979[21:2]} + 21'h00_0fb9;
  assign sel_88180 = $signed({1'h0, smod_87913[15:0]}) < $signed({1'h0, sel_87986}) ? smod_87913[15:0] : sel_87986;
  assign umul_88181 = umul22b_16b_x_6b(array_index_88003, 6'h3b);
  assign add_88183 = {1'h0, umul_87987[21:1]} + 22'h00_1f59;
  assign sel_88188 = $signed({1'h0, smod_87918[15:0]}) < $signed({1'h0, sel_87994}) ? smod_87918[15:0] : sel_87994;
  assign umul_88189 = umul22b_16b_x_6b(array_index_88009, 6'h3b);
  assign add_88191 = {1'h0, umul_87995[21:1]} + 22'h00_1f59;
  assign sel_88196 = $signed({1'h0, smod_87923[15:0]}) < $signed({1'h0, sel_88002}) ? smod_87923[15:0] : sel_88002;
  assign array_index_88197 = set1_unflattened[6'h0b];
  assign smod_88201 = $unsigned($signed({9'h000, add_88065, umul_87869[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_88203 = set2_unflattened[6'h0b];
  assign smod_88207 = $unsigned($signed({9'h000, add_88073, umul_87877[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_88257 = umul22b_16b_x_6b(array_index_88197, 6'h35);
  assign add_88259 = {1'h0, umul_88063[21:7]} + 16'h007d;
  assign sel_88264 = $signed({1'h0, smod_88007[15:0]}) < $signed({1'h0, sel_88070}) ? smod_88007[15:0] : sel_88070;
  assign umul_88265 = umul22b_16b_x_6b(array_index_88203, 6'h35);
  assign add_88267 = {1'h0, umul_88071[21:7]} + 16'h007d;
  assign sel_88272 = $signed({1'h0, smod_88013[15:0]}) < $signed({1'h0, sel_88078}) ? smod_88013[15:0] : sel_88078;
  assign smod_88276 = $unsigned($signed({8'h00, add_88135, umul_87939[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_88281 = $unsigned($signed({8'h00, add_88143, umul_87947[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_88286 = $unsigned($signed({8'h00, add_88151, umul_87955[0]}) % $signed(32'h0000_3ffd));
  assign smod_88291 = $unsigned($signed({8'h00, add_88159, umul_87963[0]}) % $signed(32'h0000_3ffd));
  assign smod_88296 = $unsigned($signed({9'h000, add_88167, umul_87971[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_88301 = $unsigned($signed({9'h000, add_88175, umul_87979[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_88306 = $unsigned($signed({9'h000, add_88183, umul_87987[0]}) % $signed(32'h0000_3ffd));
  assign smod_88311 = $unsigned($signed({9'h000, add_88191, umul_87995[0]}) % $signed(32'h0000_3ffd));
  assign umul_88327 = umul23b_16b_x_7b(array_index_87615, 7'h49);
  assign add_88329 = {1'h0, umul_88133[22:3]} + 21'h00_07e9;
  assign sel_88334 = $signed({1'h0, smod_88082[15:0]}) < $signed({1'h0, sel_88140}) ? smod_88082[15:0] : sel_88140;
  assign umul_88335 = umul23b_16b_x_7b(array_index_87621, 7'h49);
  assign add_88337 = {1'h0, umul_88141[22:3]} + 21'h00_07e9;
  assign sel_88342 = $signed({1'h0, smod_88087[15:0]}) < $signed({1'h0, sel_88148}) ? smod_88087[15:0] : sel_88148;
  assign umul_88343 = umul23b_16b_x_7b(array_index_87809, 7'h47);
  assign add_88345 = {1'h0, umul_88149[22:1]} + 23'h00_1f8b;
  assign sel_88350 = $signed({1'h0, smod_88092[15:0]}) < $signed({1'h0, sel_88156}) ? smod_88092[15:0] : sel_88156;
  assign umul_88351 = umul23b_16b_x_7b(array_index_87815, 7'h47);
  assign add_88353 = {1'h0, umul_88157[22:1]} + 23'h00_1f8b;
  assign sel_88358 = $signed({1'h0, smod_88097[15:0]}) < $signed({1'h0, sel_88164}) ? smod_88097[15:0] : sel_88164;
  assign umul_88359 = umul22b_16b_x_6b(array_index_88003, 6'h3d);
  assign add_88361 = {1'h0, umul_88165[21:2]} + 21'h00_0fb9;
  assign sel_88366 = $signed({1'h0, smod_88102[15:0]}) < $signed({1'h0, sel_88172}) ? smod_88102[15:0] : sel_88172;
  assign umul_88367 = umul22b_16b_x_6b(array_index_88009, 6'h3d);
  assign add_88369 = {1'h0, umul_88173[21:2]} + 21'h00_0fb9;
  assign sel_88374 = $signed({1'h0, smod_88107[15:0]}) < $signed({1'h0, sel_88180}) ? smod_88107[15:0] : sel_88180;
  assign umul_88375 = umul22b_16b_x_6b(array_index_88197, 6'h3b);
  assign add_88377 = {1'h0, umul_88181[21:1]} + 22'h00_1f59;
  assign sel_88382 = $signed({1'h0, smod_88112[15:0]}) < $signed({1'h0, sel_88188}) ? smod_88112[15:0] : sel_88188;
  assign umul_88383 = umul22b_16b_x_6b(array_index_88203, 6'h3b);
  assign add_88385 = {1'h0, umul_88189[21:1]} + 22'h00_1f59;
  assign sel_88390 = $signed({1'h0, smod_88117[15:0]}) < $signed({1'h0, sel_88196}) ? smod_88117[15:0] : sel_88196;
  assign array_index_88391 = set1_unflattened[6'h0c];
  assign smod_88395 = $unsigned($signed({9'h000, add_88259, umul_88063[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_88397 = set2_unflattened[6'h0c];
  assign smod_88401 = $unsigned($signed({9'h000, add_88267, umul_88071[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_88451 = umul22b_16b_x_6b(array_index_88391, 6'h35);
  assign add_88453 = {1'h0, umul_88257[21:7]} + 16'h007d;
  assign sel_88458 = $signed({1'h0, smod_88201[15:0]}) < $signed({1'h0, sel_88264}) ? smod_88201[15:0] : sel_88264;
  assign umul_88459 = umul22b_16b_x_6b(array_index_88397, 6'h35);
  assign add_88461 = {1'h0, umul_88265[21:7]} + 16'h007d;
  assign sel_88466 = $signed({1'h0, smod_88207[15:0]}) < $signed({1'h0, sel_88272}) ? smod_88207[15:0] : sel_88272;
  assign smod_88470 = $unsigned($signed({8'h00, add_88329, umul_88133[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_88475 = $unsigned($signed({8'h00, add_88337, umul_88141[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_88480 = $unsigned($signed({8'h00, add_88345, umul_88149[0]}) % $signed(32'h0000_3ffd));
  assign smod_88485 = $unsigned($signed({8'h00, add_88353, umul_88157[0]}) % $signed(32'h0000_3ffd));
  assign smod_88490 = $unsigned($signed({9'h000, add_88361, umul_88165[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_88495 = $unsigned($signed({9'h000, add_88369, umul_88173[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_88500 = $unsigned($signed({9'h000, add_88377, umul_88181[0]}) % $signed(32'h0000_3ffd));
  assign smod_88505 = $unsigned($signed({9'h000, add_88385, umul_88189[0]}) % $signed(32'h0000_3ffd));
  assign umul_88521 = umul23b_16b_x_7b(array_index_87809, 7'h49);
  assign add_88523 = {1'h0, umul_88327[22:3]} + 21'h00_07e9;
  assign sel_88528 = $signed({1'h0, smod_88276[15:0]}) < $signed({1'h0, sel_88334}) ? smod_88276[15:0] : sel_88334;
  assign umul_88529 = umul23b_16b_x_7b(array_index_87815, 7'h49);
  assign add_88531 = {1'h0, umul_88335[22:3]} + 21'h00_07e9;
  assign sel_88536 = $signed({1'h0, smod_88281[15:0]}) < $signed({1'h0, sel_88342}) ? smod_88281[15:0] : sel_88342;
  assign umul_88537 = umul23b_16b_x_7b(array_index_88003, 7'h47);
  assign add_88539 = {1'h0, umul_88343[22:1]} + 23'h00_1f8b;
  assign sel_88544 = $signed({1'h0, smod_88286[15:0]}) < $signed({1'h0, sel_88350}) ? smod_88286[15:0] : sel_88350;
  assign umul_88545 = umul23b_16b_x_7b(array_index_88009, 7'h47);
  assign add_88547 = {1'h0, umul_88351[22:1]} + 23'h00_1f8b;
  assign sel_88552 = $signed({1'h0, smod_88291[15:0]}) < $signed({1'h0, sel_88358}) ? smod_88291[15:0] : sel_88358;
  assign umul_88553 = umul22b_16b_x_6b(array_index_88197, 6'h3d);
  assign add_88555 = {1'h0, umul_88359[21:2]} + 21'h00_0fb9;
  assign sel_88560 = $signed({1'h0, smod_88296[15:0]}) < $signed({1'h0, sel_88366}) ? smod_88296[15:0] : sel_88366;
  assign umul_88561 = umul22b_16b_x_6b(array_index_88203, 6'h3d);
  assign add_88563 = {1'h0, umul_88367[21:2]} + 21'h00_0fb9;
  assign sel_88568 = $signed({1'h0, smod_88301[15:0]}) < $signed({1'h0, sel_88374}) ? smod_88301[15:0] : sel_88374;
  assign umul_88569 = umul22b_16b_x_6b(array_index_88391, 6'h3b);
  assign add_88571 = {1'h0, umul_88375[21:1]} + 22'h00_1f59;
  assign sel_88576 = $signed({1'h0, smod_88306[15:0]}) < $signed({1'h0, sel_88382}) ? smod_88306[15:0] : sel_88382;
  assign umul_88577 = umul22b_16b_x_6b(array_index_88397, 6'h3b);
  assign add_88579 = {1'h0, umul_88383[21:1]} + 22'h00_1f59;
  assign sel_88584 = $signed({1'h0, smod_88311[15:0]}) < $signed({1'h0, sel_88390}) ? smod_88311[15:0] : sel_88390;
  assign array_index_88585 = set1_unflattened[6'h0d];
  assign smod_88589 = $unsigned($signed({9'h000, add_88453, umul_88257[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_88591 = set2_unflattened[6'h0d];
  assign smod_88595 = $unsigned($signed({9'h000, add_88461, umul_88265[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_88645 = umul22b_16b_x_6b(array_index_88585, 6'h35);
  assign add_88647 = {1'h0, umul_88451[21:7]} + 16'h007d;
  assign sel_88652 = $signed({1'h0, smod_88395[15:0]}) < $signed({1'h0, sel_88458}) ? smod_88395[15:0] : sel_88458;
  assign umul_88653 = umul22b_16b_x_6b(array_index_88591, 6'h35);
  assign add_88655 = {1'h0, umul_88459[21:7]} + 16'h007d;
  assign sel_88660 = $signed({1'h0, smod_88401[15:0]}) < $signed({1'h0, sel_88466}) ? smod_88401[15:0] : sel_88466;
  assign smod_88664 = $unsigned($signed({8'h00, add_88523, umul_88327[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_88669 = $unsigned($signed({8'h00, add_88531, umul_88335[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_88674 = $unsigned($signed({8'h00, add_88539, umul_88343[0]}) % $signed(32'h0000_3ffd));
  assign smod_88679 = $unsigned($signed({8'h00, add_88547, umul_88351[0]}) % $signed(32'h0000_3ffd));
  assign smod_88684 = $unsigned($signed({9'h000, add_88555, umul_88359[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_88689 = $unsigned($signed({9'h000, add_88563, umul_88367[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_88694 = $unsigned($signed({9'h000, add_88571, umul_88375[0]}) % $signed(32'h0000_3ffd));
  assign smod_88699 = $unsigned($signed({9'h000, add_88579, umul_88383[0]}) % $signed(32'h0000_3ffd));
  assign umul_88715 = umul23b_16b_x_7b(array_index_88003, 7'h49);
  assign add_88717 = {1'h0, umul_88521[22:3]} + 21'h00_07e9;
  assign sel_88722 = $signed({1'h0, smod_88470[15:0]}) < $signed({1'h0, sel_88528}) ? smod_88470[15:0] : sel_88528;
  assign umul_88723 = umul23b_16b_x_7b(array_index_88009, 7'h49);
  assign add_88725 = {1'h0, umul_88529[22:3]} + 21'h00_07e9;
  assign sel_88730 = $signed({1'h0, smod_88475[15:0]}) < $signed({1'h0, sel_88536}) ? smod_88475[15:0] : sel_88536;
  assign umul_88731 = umul23b_16b_x_7b(array_index_88197, 7'h47);
  assign add_88733 = {1'h0, umul_88537[22:1]} + 23'h00_1f8b;
  assign sel_88738 = $signed({1'h0, smod_88480[15:0]}) < $signed({1'h0, sel_88544}) ? smod_88480[15:0] : sel_88544;
  assign umul_88739 = umul23b_16b_x_7b(array_index_88203, 7'h47);
  assign add_88741 = {1'h0, umul_88545[22:1]} + 23'h00_1f8b;
  assign sel_88746 = $signed({1'h0, smod_88485[15:0]}) < $signed({1'h0, sel_88552}) ? smod_88485[15:0] : sel_88552;
  assign umul_88747 = umul22b_16b_x_6b(array_index_88391, 6'h3d);
  assign add_88749 = {1'h0, umul_88553[21:2]} + 21'h00_0fb9;
  assign sel_88754 = $signed({1'h0, smod_88490[15:0]}) < $signed({1'h0, sel_88560}) ? smod_88490[15:0] : sel_88560;
  assign umul_88755 = umul22b_16b_x_6b(array_index_88397, 6'h3d);
  assign add_88757 = {1'h0, umul_88561[21:2]} + 21'h00_0fb9;
  assign sel_88762 = $signed({1'h0, smod_88495[15:0]}) < $signed({1'h0, sel_88568}) ? smod_88495[15:0] : sel_88568;
  assign umul_88763 = umul22b_16b_x_6b(array_index_88585, 6'h3b);
  assign add_88765 = {1'h0, umul_88569[21:1]} + 22'h00_1f59;
  assign sel_88770 = $signed({1'h0, smod_88500[15:0]}) < $signed({1'h0, sel_88576}) ? smod_88500[15:0] : sel_88576;
  assign umul_88771 = umul22b_16b_x_6b(array_index_88591, 6'h3b);
  assign add_88773 = {1'h0, umul_88577[21:1]} + 22'h00_1f59;
  assign sel_88778 = $signed({1'h0, smod_88505[15:0]}) < $signed({1'h0, sel_88584}) ? smod_88505[15:0] : sel_88584;
  assign array_index_88779 = set1_unflattened[6'h0e];
  assign smod_88783 = $unsigned($signed({9'h000, add_88647, umul_88451[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_88785 = set2_unflattened[6'h0e];
  assign smod_88789 = $unsigned($signed({9'h000, add_88655, umul_88459[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_88839 = umul22b_16b_x_6b(array_index_88779, 6'h35);
  assign add_88841 = {1'h0, umul_88645[21:7]} + 16'h007d;
  assign sel_88846 = $signed({1'h0, smod_88589[15:0]}) < $signed({1'h0, sel_88652}) ? smod_88589[15:0] : sel_88652;
  assign umul_88847 = umul22b_16b_x_6b(array_index_88785, 6'h35);
  assign add_88849 = {1'h0, umul_88653[21:7]} + 16'h007d;
  assign sel_88854 = $signed({1'h0, smod_88595[15:0]}) < $signed({1'h0, sel_88660}) ? smod_88595[15:0] : sel_88660;
  assign smod_88858 = $unsigned($signed({8'h00, add_88717, umul_88521[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_88863 = $unsigned($signed({8'h00, add_88725, umul_88529[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_88868 = $unsigned($signed({8'h00, add_88733, umul_88537[0]}) % $signed(32'h0000_3ffd));
  assign smod_88873 = $unsigned($signed({8'h00, add_88741, umul_88545[0]}) % $signed(32'h0000_3ffd));
  assign smod_88878 = $unsigned($signed({9'h000, add_88749, umul_88553[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_88883 = $unsigned($signed({9'h000, add_88757, umul_88561[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_88888 = $unsigned($signed({9'h000, add_88765, umul_88569[0]}) % $signed(32'h0000_3ffd));
  assign smod_88893 = $unsigned($signed({9'h000, add_88773, umul_88577[0]}) % $signed(32'h0000_3ffd));
  assign umul_88909 = umul23b_16b_x_7b(array_index_88197, 7'h49);
  assign add_88911 = {1'h0, umul_88715[22:3]} + 21'h00_07e9;
  assign sel_88916 = $signed({1'h0, smod_88664[15:0]}) < $signed({1'h0, sel_88722}) ? smod_88664[15:0] : sel_88722;
  assign umul_88917 = umul23b_16b_x_7b(array_index_88203, 7'h49);
  assign add_88919 = {1'h0, umul_88723[22:3]} + 21'h00_07e9;
  assign sel_88924 = $signed({1'h0, smod_88669[15:0]}) < $signed({1'h0, sel_88730}) ? smod_88669[15:0] : sel_88730;
  assign umul_88925 = umul23b_16b_x_7b(array_index_88391, 7'h47);
  assign add_88927 = {1'h0, umul_88731[22:1]} + 23'h00_1f8b;
  assign sel_88932 = $signed({1'h0, smod_88674[15:0]}) < $signed({1'h0, sel_88738}) ? smod_88674[15:0] : sel_88738;
  assign umul_88933 = umul23b_16b_x_7b(array_index_88397, 7'h47);
  assign add_88935 = {1'h0, umul_88739[22:1]} + 23'h00_1f8b;
  assign sel_88940 = $signed({1'h0, smod_88679[15:0]}) < $signed({1'h0, sel_88746}) ? smod_88679[15:0] : sel_88746;
  assign umul_88941 = umul22b_16b_x_6b(array_index_88585, 6'h3d);
  assign add_88943 = {1'h0, umul_88747[21:2]} + 21'h00_0fb9;
  assign sel_88948 = $signed({1'h0, smod_88684[15:0]}) < $signed({1'h0, sel_88754}) ? smod_88684[15:0] : sel_88754;
  assign umul_88949 = umul22b_16b_x_6b(array_index_88591, 6'h3d);
  assign add_88951 = {1'h0, umul_88755[21:2]} + 21'h00_0fb9;
  assign sel_88956 = $signed({1'h0, smod_88689[15:0]}) < $signed({1'h0, sel_88762}) ? smod_88689[15:0] : sel_88762;
  assign umul_88957 = umul22b_16b_x_6b(array_index_88779, 6'h3b);
  assign add_88959 = {1'h0, umul_88763[21:1]} + 22'h00_1f59;
  assign sel_88964 = $signed({1'h0, smod_88694[15:0]}) < $signed({1'h0, sel_88770}) ? smod_88694[15:0] : sel_88770;
  assign umul_88965 = umul22b_16b_x_6b(array_index_88785, 6'h3b);
  assign add_88967 = {1'h0, umul_88771[21:1]} + 22'h00_1f59;
  assign sel_88972 = $signed({1'h0, smod_88699[15:0]}) < $signed({1'h0, sel_88778}) ? smod_88699[15:0] : sel_88778;
  assign array_index_88973 = set1_unflattened[6'h0f];
  assign smod_88977 = $unsigned($signed({9'h000, add_88841, umul_88645[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_88979 = set2_unflattened[6'h0f];
  assign smod_88983 = $unsigned($signed({9'h000, add_88849, umul_88653[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_89033 = umul22b_16b_x_6b(array_index_88973, 6'h35);
  assign add_89035 = {1'h0, umul_88839[21:7]} + 16'h007d;
  assign sel_89040 = $signed({1'h0, smod_88783[15:0]}) < $signed({1'h0, sel_88846}) ? smod_88783[15:0] : sel_88846;
  assign umul_89041 = umul22b_16b_x_6b(array_index_88979, 6'h35);
  assign add_89043 = {1'h0, umul_88847[21:7]} + 16'h007d;
  assign sel_89048 = $signed({1'h0, smod_88789[15:0]}) < $signed({1'h0, sel_88854}) ? smod_88789[15:0] : sel_88854;
  assign smod_89052 = $unsigned($signed({8'h00, add_88911, umul_88715[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_89057 = $unsigned($signed({8'h00, add_88919, umul_88723[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_89062 = $unsigned($signed({8'h00, add_88927, umul_88731[0]}) % $signed(32'h0000_3ffd));
  assign smod_89067 = $unsigned($signed({8'h00, add_88935, umul_88739[0]}) % $signed(32'h0000_3ffd));
  assign smod_89072 = $unsigned($signed({9'h000, add_88943, umul_88747[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_89077 = $unsigned($signed({9'h000, add_88951, umul_88755[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_89082 = $unsigned($signed({9'h000, add_88959, umul_88763[0]}) % $signed(32'h0000_3ffd));
  assign smod_89087 = $unsigned($signed({9'h000, add_88967, umul_88771[0]}) % $signed(32'h0000_3ffd));
  assign umul_89103 = umul23b_16b_x_7b(array_index_88391, 7'h49);
  assign add_89105 = {1'h0, umul_88909[22:3]} + 21'h00_07e9;
  assign sel_89110 = $signed({1'h0, smod_88858[15:0]}) < $signed({1'h0, sel_88916}) ? smod_88858[15:0] : sel_88916;
  assign umul_89111 = umul23b_16b_x_7b(array_index_88397, 7'h49);
  assign add_89113 = {1'h0, umul_88917[22:3]} + 21'h00_07e9;
  assign sel_89118 = $signed({1'h0, smod_88863[15:0]}) < $signed({1'h0, sel_88924}) ? smod_88863[15:0] : sel_88924;
  assign umul_89119 = umul23b_16b_x_7b(array_index_88585, 7'h47);
  assign add_89121 = {1'h0, umul_88925[22:1]} + 23'h00_1f8b;
  assign sel_89126 = $signed({1'h0, smod_88868[15:0]}) < $signed({1'h0, sel_88932}) ? smod_88868[15:0] : sel_88932;
  assign umul_89127 = umul23b_16b_x_7b(array_index_88591, 7'h47);
  assign add_89129 = {1'h0, umul_88933[22:1]} + 23'h00_1f8b;
  assign sel_89134 = $signed({1'h0, smod_88873[15:0]}) < $signed({1'h0, sel_88940}) ? smod_88873[15:0] : sel_88940;
  assign umul_89135 = umul22b_16b_x_6b(array_index_88779, 6'h3d);
  assign add_89137 = {1'h0, umul_88941[21:2]} + 21'h00_0fb9;
  assign sel_89142 = $signed({1'h0, smod_88878[15:0]}) < $signed({1'h0, sel_88948}) ? smod_88878[15:0] : sel_88948;
  assign umul_89143 = umul22b_16b_x_6b(array_index_88785, 6'h3d);
  assign add_89145 = {1'h0, umul_88949[21:2]} + 21'h00_0fb9;
  assign sel_89150 = $signed({1'h0, smod_88883[15:0]}) < $signed({1'h0, sel_88956}) ? smod_88883[15:0] : sel_88956;
  assign umul_89151 = umul22b_16b_x_6b(array_index_88973, 6'h3b);
  assign add_89153 = {1'h0, umul_88957[21:1]} + 22'h00_1f59;
  assign sel_89158 = $signed({1'h0, smod_88888[15:0]}) < $signed({1'h0, sel_88964}) ? smod_88888[15:0] : sel_88964;
  assign umul_89159 = umul22b_16b_x_6b(array_index_88979, 6'h3b);
  assign add_89161 = {1'h0, umul_88965[21:1]} + 22'h00_1f59;
  assign sel_89166 = $signed({1'h0, smod_88893[15:0]}) < $signed({1'h0, sel_88972}) ? smod_88893[15:0] : sel_88972;
  assign array_index_89167 = set1_unflattened[6'h10];
  assign smod_89171 = $unsigned($signed({9'h000, add_89035, umul_88839[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_89173 = set2_unflattened[6'h10];
  assign smod_89177 = $unsigned($signed({9'h000, add_89043, umul_88847[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_89227 = umul22b_16b_x_6b(array_index_89167, 6'h35);
  assign add_89229 = {1'h0, umul_89033[21:7]} + 16'h007d;
  assign sel_89234 = $signed({1'h0, smod_88977[15:0]}) < $signed({1'h0, sel_89040}) ? smod_88977[15:0] : sel_89040;
  assign umul_89235 = umul22b_16b_x_6b(array_index_89173, 6'h35);
  assign add_89237 = {1'h0, umul_89041[21:7]} + 16'h007d;
  assign sel_89242 = $signed({1'h0, smod_88983[15:0]}) < $signed({1'h0, sel_89048}) ? smod_88983[15:0] : sel_89048;
  assign smod_89246 = $unsigned($signed({8'h00, add_89105, umul_88909[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_89251 = $unsigned($signed({8'h00, add_89113, umul_88917[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_89256 = $unsigned($signed({8'h00, add_89121, umul_88925[0]}) % $signed(32'h0000_3ffd));
  assign smod_89261 = $unsigned($signed({8'h00, add_89129, umul_88933[0]}) % $signed(32'h0000_3ffd));
  assign smod_89266 = $unsigned($signed({9'h000, add_89137, umul_88941[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_89271 = $unsigned($signed({9'h000, add_89145, umul_88949[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_89276 = $unsigned($signed({9'h000, add_89153, umul_88957[0]}) % $signed(32'h0000_3ffd));
  assign smod_89281 = $unsigned($signed({9'h000, add_89161, umul_88965[0]}) % $signed(32'h0000_3ffd));
  assign umul_89297 = umul23b_16b_x_7b(array_index_88585, 7'h49);
  assign add_89299 = {1'h0, umul_89103[22:3]} + 21'h00_07e9;
  assign sel_89304 = $signed({1'h0, smod_89052[15:0]}) < $signed({1'h0, sel_89110}) ? smod_89052[15:0] : sel_89110;
  assign umul_89305 = umul23b_16b_x_7b(array_index_88591, 7'h49);
  assign add_89307 = {1'h0, umul_89111[22:3]} + 21'h00_07e9;
  assign sel_89312 = $signed({1'h0, smod_89057[15:0]}) < $signed({1'h0, sel_89118}) ? smod_89057[15:0] : sel_89118;
  assign umul_89313 = umul23b_16b_x_7b(array_index_88779, 7'h47);
  assign add_89315 = {1'h0, umul_89119[22:1]} + 23'h00_1f8b;
  assign sel_89320 = $signed({1'h0, smod_89062[15:0]}) < $signed({1'h0, sel_89126}) ? smod_89062[15:0] : sel_89126;
  assign umul_89321 = umul23b_16b_x_7b(array_index_88785, 7'h47);
  assign add_89323 = {1'h0, umul_89127[22:1]} + 23'h00_1f8b;
  assign sel_89328 = $signed({1'h0, smod_89067[15:0]}) < $signed({1'h0, sel_89134}) ? smod_89067[15:0] : sel_89134;
  assign umul_89329 = umul22b_16b_x_6b(array_index_88973, 6'h3d);
  assign add_89331 = {1'h0, umul_89135[21:2]} + 21'h00_0fb9;
  assign sel_89336 = $signed({1'h0, smod_89072[15:0]}) < $signed({1'h0, sel_89142}) ? smod_89072[15:0] : sel_89142;
  assign umul_89337 = umul22b_16b_x_6b(array_index_88979, 6'h3d);
  assign add_89339 = {1'h0, umul_89143[21:2]} + 21'h00_0fb9;
  assign sel_89344 = $signed({1'h0, smod_89077[15:0]}) < $signed({1'h0, sel_89150}) ? smod_89077[15:0] : sel_89150;
  assign umul_89345 = umul22b_16b_x_6b(array_index_89167, 6'h3b);
  assign add_89347 = {1'h0, umul_89151[21:1]} + 22'h00_1f59;
  assign sel_89352 = $signed({1'h0, smod_89082[15:0]}) < $signed({1'h0, sel_89158}) ? smod_89082[15:0] : sel_89158;
  assign umul_89353 = umul22b_16b_x_6b(array_index_89173, 6'h3b);
  assign add_89355 = {1'h0, umul_89159[21:1]} + 22'h00_1f59;
  assign sel_89360 = $signed({1'h0, smod_89087[15:0]}) < $signed({1'h0, sel_89166}) ? smod_89087[15:0] : sel_89166;
  assign array_index_89361 = set1_unflattened[6'h11];
  assign smod_89365 = $unsigned($signed({9'h000, add_89229, umul_89033[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_89367 = set2_unflattened[6'h11];
  assign smod_89371 = $unsigned($signed({9'h000, add_89237, umul_89041[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_89421 = umul22b_16b_x_6b(array_index_89361, 6'h35);
  assign add_89423 = {1'h0, umul_89227[21:7]} + 16'h007d;
  assign sel_89428 = $signed({1'h0, smod_89171[15:0]}) < $signed({1'h0, sel_89234}) ? smod_89171[15:0] : sel_89234;
  assign umul_89429 = umul22b_16b_x_6b(array_index_89367, 6'h35);
  assign add_89431 = {1'h0, umul_89235[21:7]} + 16'h007d;
  assign sel_89436 = $signed({1'h0, smod_89177[15:0]}) < $signed({1'h0, sel_89242}) ? smod_89177[15:0] : sel_89242;
  assign smod_89440 = $unsigned($signed({8'h00, add_89299, umul_89103[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_89445 = $unsigned($signed({8'h00, add_89307, umul_89111[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_89450 = $unsigned($signed({8'h00, add_89315, umul_89119[0]}) % $signed(32'h0000_3ffd));
  assign smod_89455 = $unsigned($signed({8'h00, add_89323, umul_89127[0]}) % $signed(32'h0000_3ffd));
  assign smod_89460 = $unsigned($signed({9'h000, add_89331, umul_89135[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_89465 = $unsigned($signed({9'h000, add_89339, umul_89143[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_89470 = $unsigned($signed({9'h000, add_89347, umul_89151[0]}) % $signed(32'h0000_3ffd));
  assign smod_89475 = $unsigned($signed({9'h000, add_89355, umul_89159[0]}) % $signed(32'h0000_3ffd));
  assign umul_89491 = umul23b_16b_x_7b(array_index_88779, 7'h49);
  assign add_89493 = {1'h0, umul_89297[22:3]} + 21'h00_07e9;
  assign sel_89498 = $signed({1'h0, smod_89246[15:0]}) < $signed({1'h0, sel_89304}) ? smod_89246[15:0] : sel_89304;
  assign umul_89499 = umul23b_16b_x_7b(array_index_88785, 7'h49);
  assign add_89501 = {1'h0, umul_89305[22:3]} + 21'h00_07e9;
  assign sel_89506 = $signed({1'h0, smod_89251[15:0]}) < $signed({1'h0, sel_89312}) ? smod_89251[15:0] : sel_89312;
  assign umul_89507 = umul23b_16b_x_7b(array_index_88973, 7'h47);
  assign add_89509 = {1'h0, umul_89313[22:1]} + 23'h00_1f8b;
  assign sel_89514 = $signed({1'h0, smod_89256[15:0]}) < $signed({1'h0, sel_89320}) ? smod_89256[15:0] : sel_89320;
  assign umul_89515 = umul23b_16b_x_7b(array_index_88979, 7'h47);
  assign add_89517 = {1'h0, umul_89321[22:1]} + 23'h00_1f8b;
  assign sel_89522 = $signed({1'h0, smod_89261[15:0]}) < $signed({1'h0, sel_89328}) ? smod_89261[15:0] : sel_89328;
  assign umul_89523 = umul22b_16b_x_6b(array_index_89167, 6'h3d);
  assign add_89525 = {1'h0, umul_89329[21:2]} + 21'h00_0fb9;
  assign sel_89530 = $signed({1'h0, smod_89266[15:0]}) < $signed({1'h0, sel_89336}) ? smod_89266[15:0] : sel_89336;
  assign umul_89531 = umul22b_16b_x_6b(array_index_89173, 6'h3d);
  assign add_89533 = {1'h0, umul_89337[21:2]} + 21'h00_0fb9;
  assign sel_89538 = $signed({1'h0, smod_89271[15:0]}) < $signed({1'h0, sel_89344}) ? smod_89271[15:0] : sel_89344;
  assign umul_89539 = umul22b_16b_x_6b(array_index_89361, 6'h3b);
  assign add_89541 = {1'h0, umul_89345[21:1]} + 22'h00_1f59;
  assign sel_89546 = $signed({1'h0, smod_89276[15:0]}) < $signed({1'h0, sel_89352}) ? smod_89276[15:0] : sel_89352;
  assign umul_89547 = umul22b_16b_x_6b(array_index_89367, 6'h3b);
  assign add_89549 = {1'h0, umul_89353[21:1]} + 22'h00_1f59;
  assign sel_89554 = $signed({1'h0, smod_89281[15:0]}) < $signed({1'h0, sel_89360}) ? smod_89281[15:0] : sel_89360;
  assign array_index_89555 = set1_unflattened[6'h12];
  assign smod_89559 = $unsigned($signed({9'h000, add_89423, umul_89227[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_89561 = set2_unflattened[6'h12];
  assign smod_89565 = $unsigned($signed({9'h000, add_89431, umul_89235[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_89615 = umul22b_16b_x_6b(array_index_89555, 6'h35);
  assign add_89617 = {1'h0, umul_89421[21:7]} + 16'h007d;
  assign sel_89622 = $signed({1'h0, smod_89365[15:0]}) < $signed({1'h0, sel_89428}) ? smod_89365[15:0] : sel_89428;
  assign umul_89623 = umul22b_16b_x_6b(array_index_89561, 6'h35);
  assign add_89625 = {1'h0, umul_89429[21:7]} + 16'h007d;
  assign sel_89630 = $signed({1'h0, smod_89371[15:0]}) < $signed({1'h0, sel_89436}) ? smod_89371[15:0] : sel_89436;
  assign smod_89634 = $unsigned($signed({8'h00, add_89493, umul_89297[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_89639 = $unsigned($signed({8'h00, add_89501, umul_89305[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_89644 = $unsigned($signed({8'h00, add_89509, umul_89313[0]}) % $signed(32'h0000_3ffd));
  assign smod_89649 = $unsigned($signed({8'h00, add_89517, umul_89321[0]}) % $signed(32'h0000_3ffd));
  assign smod_89654 = $unsigned($signed({9'h000, add_89525, umul_89329[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_89659 = $unsigned($signed({9'h000, add_89533, umul_89337[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_89664 = $unsigned($signed({9'h000, add_89541, umul_89345[0]}) % $signed(32'h0000_3ffd));
  assign smod_89669 = $unsigned($signed({9'h000, add_89549, umul_89353[0]}) % $signed(32'h0000_3ffd));
  assign umul_89685 = umul23b_16b_x_7b(array_index_88973, 7'h49);
  assign add_89687 = {1'h0, umul_89491[22:3]} + 21'h00_07e9;
  assign sel_89692 = $signed({1'h0, smod_89440[15:0]}) < $signed({1'h0, sel_89498}) ? smod_89440[15:0] : sel_89498;
  assign umul_89693 = umul23b_16b_x_7b(array_index_88979, 7'h49);
  assign add_89695 = {1'h0, umul_89499[22:3]} + 21'h00_07e9;
  assign sel_89700 = $signed({1'h0, smod_89445[15:0]}) < $signed({1'h0, sel_89506}) ? smod_89445[15:0] : sel_89506;
  assign umul_89701 = umul23b_16b_x_7b(array_index_89167, 7'h47);
  assign add_89703 = {1'h0, umul_89507[22:1]} + 23'h00_1f8b;
  assign sel_89708 = $signed({1'h0, smod_89450[15:0]}) < $signed({1'h0, sel_89514}) ? smod_89450[15:0] : sel_89514;
  assign umul_89709 = umul23b_16b_x_7b(array_index_89173, 7'h47);
  assign add_89711 = {1'h0, umul_89515[22:1]} + 23'h00_1f8b;
  assign sel_89716 = $signed({1'h0, smod_89455[15:0]}) < $signed({1'h0, sel_89522}) ? smod_89455[15:0] : sel_89522;
  assign umul_89717 = umul22b_16b_x_6b(array_index_89361, 6'h3d);
  assign add_89719 = {1'h0, umul_89523[21:2]} + 21'h00_0fb9;
  assign sel_89724 = $signed({1'h0, smod_89460[15:0]}) < $signed({1'h0, sel_89530}) ? smod_89460[15:0] : sel_89530;
  assign umul_89725 = umul22b_16b_x_6b(array_index_89367, 6'h3d);
  assign add_89727 = {1'h0, umul_89531[21:2]} + 21'h00_0fb9;
  assign sel_89732 = $signed({1'h0, smod_89465[15:0]}) < $signed({1'h0, sel_89538}) ? smod_89465[15:0] : sel_89538;
  assign umul_89733 = umul22b_16b_x_6b(array_index_89555, 6'h3b);
  assign add_89735 = {1'h0, umul_89539[21:1]} + 22'h00_1f59;
  assign sel_89740 = $signed({1'h0, smod_89470[15:0]}) < $signed({1'h0, sel_89546}) ? smod_89470[15:0] : sel_89546;
  assign umul_89741 = umul22b_16b_x_6b(array_index_89561, 6'h3b);
  assign add_89743 = {1'h0, umul_89547[21:1]} + 22'h00_1f59;
  assign sel_89748 = $signed({1'h0, smod_89475[15:0]}) < $signed({1'h0, sel_89554}) ? smod_89475[15:0] : sel_89554;
  assign array_index_89749 = set1_unflattened[6'h13];
  assign smod_89753 = $unsigned($signed({9'h000, add_89617, umul_89421[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_89755 = set2_unflattened[6'h13];
  assign smod_89759 = $unsigned($signed({9'h000, add_89625, umul_89429[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_89809 = umul22b_16b_x_6b(array_index_89749, 6'h35);
  assign add_89811 = {1'h0, umul_89615[21:7]} + 16'h007d;
  assign sel_89816 = $signed({1'h0, smod_89559[15:0]}) < $signed({1'h0, sel_89622}) ? smod_89559[15:0] : sel_89622;
  assign umul_89817 = umul22b_16b_x_6b(array_index_89755, 6'h35);
  assign add_89819 = {1'h0, umul_89623[21:7]} + 16'h007d;
  assign sel_89824 = $signed({1'h0, smod_89565[15:0]}) < $signed({1'h0, sel_89630}) ? smod_89565[15:0] : sel_89630;
  assign smod_89828 = $unsigned($signed({8'h00, add_89687, umul_89491[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_89833 = $unsigned($signed({8'h00, add_89695, umul_89499[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_89838 = $unsigned($signed({8'h00, add_89703, umul_89507[0]}) % $signed(32'h0000_3ffd));
  assign smod_89843 = $unsigned($signed({8'h00, add_89711, umul_89515[0]}) % $signed(32'h0000_3ffd));
  assign smod_89848 = $unsigned($signed({9'h000, add_89719, umul_89523[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_89853 = $unsigned($signed({9'h000, add_89727, umul_89531[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_89858 = $unsigned($signed({9'h000, add_89735, umul_89539[0]}) % $signed(32'h0000_3ffd));
  assign smod_89863 = $unsigned($signed({9'h000, add_89743, umul_89547[0]}) % $signed(32'h0000_3ffd));
  assign umul_89879 = umul23b_16b_x_7b(array_index_89167, 7'h49);
  assign add_89881 = {1'h0, umul_89685[22:3]} + 21'h00_07e9;
  assign sel_89886 = $signed({1'h0, smod_89634[15:0]}) < $signed({1'h0, sel_89692}) ? smod_89634[15:0] : sel_89692;
  assign umul_89887 = umul23b_16b_x_7b(array_index_89173, 7'h49);
  assign add_89889 = {1'h0, umul_89693[22:3]} + 21'h00_07e9;
  assign sel_89894 = $signed({1'h0, smod_89639[15:0]}) < $signed({1'h0, sel_89700}) ? smod_89639[15:0] : sel_89700;
  assign umul_89895 = umul23b_16b_x_7b(array_index_89361, 7'h47);
  assign add_89897 = {1'h0, umul_89701[22:1]} + 23'h00_1f8b;
  assign sel_89902 = $signed({1'h0, smod_89644[15:0]}) < $signed({1'h0, sel_89708}) ? smod_89644[15:0] : sel_89708;
  assign umul_89903 = umul23b_16b_x_7b(array_index_89367, 7'h47);
  assign add_89905 = {1'h0, umul_89709[22:1]} + 23'h00_1f8b;
  assign sel_89910 = $signed({1'h0, smod_89649[15:0]}) < $signed({1'h0, sel_89716}) ? smod_89649[15:0] : sel_89716;
  assign umul_89911 = umul22b_16b_x_6b(array_index_89555, 6'h3d);
  assign add_89913 = {1'h0, umul_89717[21:2]} + 21'h00_0fb9;
  assign sel_89918 = $signed({1'h0, smod_89654[15:0]}) < $signed({1'h0, sel_89724}) ? smod_89654[15:0] : sel_89724;
  assign umul_89919 = umul22b_16b_x_6b(array_index_89561, 6'h3d);
  assign add_89921 = {1'h0, umul_89725[21:2]} + 21'h00_0fb9;
  assign sel_89926 = $signed({1'h0, smod_89659[15:0]}) < $signed({1'h0, sel_89732}) ? smod_89659[15:0] : sel_89732;
  assign umul_89927 = umul22b_16b_x_6b(array_index_89749, 6'h3b);
  assign add_89929 = {1'h0, umul_89733[21:1]} + 22'h00_1f59;
  assign sel_89934 = $signed({1'h0, smod_89664[15:0]}) < $signed({1'h0, sel_89740}) ? smod_89664[15:0] : sel_89740;
  assign umul_89935 = umul22b_16b_x_6b(array_index_89755, 6'h3b);
  assign add_89937 = {1'h0, umul_89741[21:1]} + 22'h00_1f59;
  assign sel_89942 = $signed({1'h0, smod_89669[15:0]}) < $signed({1'h0, sel_89748}) ? smod_89669[15:0] : sel_89748;
  assign array_index_89943 = set1_unflattened[6'h14];
  assign smod_89947 = $unsigned($signed({9'h000, add_89811, umul_89615[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_89949 = set2_unflattened[6'h14];
  assign smod_89953 = $unsigned($signed({9'h000, add_89819, umul_89623[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_90003 = umul22b_16b_x_6b(array_index_89943, 6'h35);
  assign add_90005 = {1'h0, umul_89809[21:7]} + 16'h007d;
  assign sel_90010 = $signed({1'h0, smod_89753[15:0]}) < $signed({1'h0, sel_89816}) ? smod_89753[15:0] : sel_89816;
  assign umul_90011 = umul22b_16b_x_6b(array_index_89949, 6'h35);
  assign add_90013 = {1'h0, umul_89817[21:7]} + 16'h007d;
  assign sel_90018 = $signed({1'h0, smod_89759[15:0]}) < $signed({1'h0, sel_89824}) ? smod_89759[15:0] : sel_89824;
  assign smod_90022 = $unsigned($signed({8'h00, add_89881, umul_89685[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_90027 = $unsigned($signed({8'h00, add_89889, umul_89693[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_90032 = $unsigned($signed({8'h00, add_89897, umul_89701[0]}) % $signed(32'h0000_3ffd));
  assign smod_90037 = $unsigned($signed({8'h00, add_89905, umul_89709[0]}) % $signed(32'h0000_3ffd));
  assign smod_90042 = $unsigned($signed({9'h000, add_89913, umul_89717[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_90047 = $unsigned($signed({9'h000, add_89921, umul_89725[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_90052 = $unsigned($signed({9'h000, add_89929, umul_89733[0]}) % $signed(32'h0000_3ffd));
  assign smod_90057 = $unsigned($signed({9'h000, add_89937, umul_89741[0]}) % $signed(32'h0000_3ffd));
  assign umul_90073 = umul23b_16b_x_7b(array_index_89361, 7'h49);
  assign add_90075 = {1'h0, umul_89879[22:3]} + 21'h00_07e9;
  assign sel_90080 = $signed({1'h0, smod_89828[15:0]}) < $signed({1'h0, sel_89886}) ? smod_89828[15:0] : sel_89886;
  assign umul_90081 = umul23b_16b_x_7b(array_index_89367, 7'h49);
  assign add_90083 = {1'h0, umul_89887[22:3]} + 21'h00_07e9;
  assign sel_90088 = $signed({1'h0, smod_89833[15:0]}) < $signed({1'h0, sel_89894}) ? smod_89833[15:0] : sel_89894;
  assign umul_90089 = umul23b_16b_x_7b(array_index_89555, 7'h47);
  assign add_90091 = {1'h0, umul_89895[22:1]} + 23'h00_1f8b;
  assign sel_90096 = $signed({1'h0, smod_89838[15:0]}) < $signed({1'h0, sel_89902}) ? smod_89838[15:0] : sel_89902;
  assign umul_90097 = umul23b_16b_x_7b(array_index_89561, 7'h47);
  assign add_90099 = {1'h0, umul_89903[22:1]} + 23'h00_1f8b;
  assign sel_90104 = $signed({1'h0, smod_89843[15:0]}) < $signed({1'h0, sel_89910}) ? smod_89843[15:0] : sel_89910;
  assign umul_90105 = umul22b_16b_x_6b(array_index_89749, 6'h3d);
  assign add_90107 = {1'h0, umul_89911[21:2]} + 21'h00_0fb9;
  assign sel_90112 = $signed({1'h0, smod_89848[15:0]}) < $signed({1'h0, sel_89918}) ? smod_89848[15:0] : sel_89918;
  assign umul_90113 = umul22b_16b_x_6b(array_index_89755, 6'h3d);
  assign add_90115 = {1'h0, umul_89919[21:2]} + 21'h00_0fb9;
  assign sel_90120 = $signed({1'h0, smod_89853[15:0]}) < $signed({1'h0, sel_89926}) ? smod_89853[15:0] : sel_89926;
  assign umul_90121 = umul22b_16b_x_6b(array_index_89943, 6'h3b);
  assign add_90123 = {1'h0, umul_89927[21:1]} + 22'h00_1f59;
  assign sel_90128 = $signed({1'h0, smod_89858[15:0]}) < $signed({1'h0, sel_89934}) ? smod_89858[15:0] : sel_89934;
  assign umul_90129 = umul22b_16b_x_6b(array_index_89949, 6'h3b);
  assign add_90131 = {1'h0, umul_89935[21:1]} + 22'h00_1f59;
  assign sel_90136 = $signed({1'h0, smod_89863[15:0]}) < $signed({1'h0, sel_89942}) ? smod_89863[15:0] : sel_89942;
  assign array_index_90137 = set1_unflattened[6'h15];
  assign smod_90141 = $unsigned($signed({9'h000, add_90005, umul_89809[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_90143 = set2_unflattened[6'h15];
  assign smod_90147 = $unsigned($signed({9'h000, add_90013, umul_89817[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_90197 = umul22b_16b_x_6b(array_index_90137, 6'h35);
  assign add_90199 = {1'h0, umul_90003[21:7]} + 16'h007d;
  assign sel_90204 = $signed({1'h0, smod_89947[15:0]}) < $signed({1'h0, sel_90010}) ? smod_89947[15:0] : sel_90010;
  assign umul_90205 = umul22b_16b_x_6b(array_index_90143, 6'h35);
  assign add_90207 = {1'h0, umul_90011[21:7]} + 16'h007d;
  assign sel_90212 = $signed({1'h0, smod_89953[15:0]}) < $signed({1'h0, sel_90018}) ? smod_89953[15:0] : sel_90018;
  assign smod_90216 = $unsigned($signed({8'h00, add_90075, umul_89879[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_90221 = $unsigned($signed({8'h00, add_90083, umul_89887[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_90226 = $unsigned($signed({8'h00, add_90091, umul_89895[0]}) % $signed(32'h0000_3ffd));
  assign smod_90231 = $unsigned($signed({8'h00, add_90099, umul_89903[0]}) % $signed(32'h0000_3ffd));
  assign smod_90236 = $unsigned($signed({9'h000, add_90107, umul_89911[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_90241 = $unsigned($signed({9'h000, add_90115, umul_89919[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_90246 = $unsigned($signed({9'h000, add_90123, umul_89927[0]}) % $signed(32'h0000_3ffd));
  assign smod_90251 = $unsigned($signed({9'h000, add_90131, umul_89935[0]}) % $signed(32'h0000_3ffd));
  assign umul_90267 = umul23b_16b_x_7b(array_index_89555, 7'h49);
  assign add_90269 = {1'h0, umul_90073[22:3]} + 21'h00_07e9;
  assign sel_90274 = $signed({1'h0, smod_90022[15:0]}) < $signed({1'h0, sel_90080}) ? smod_90022[15:0] : sel_90080;
  assign umul_90275 = umul23b_16b_x_7b(array_index_89561, 7'h49);
  assign add_90277 = {1'h0, umul_90081[22:3]} + 21'h00_07e9;
  assign sel_90282 = $signed({1'h0, smod_90027[15:0]}) < $signed({1'h0, sel_90088}) ? smod_90027[15:0] : sel_90088;
  assign umul_90283 = umul23b_16b_x_7b(array_index_89749, 7'h47);
  assign add_90285 = {1'h0, umul_90089[22:1]} + 23'h00_1f8b;
  assign sel_90290 = $signed({1'h0, smod_90032[15:0]}) < $signed({1'h0, sel_90096}) ? smod_90032[15:0] : sel_90096;
  assign umul_90291 = umul23b_16b_x_7b(array_index_89755, 7'h47);
  assign add_90293 = {1'h0, umul_90097[22:1]} + 23'h00_1f8b;
  assign sel_90298 = $signed({1'h0, smod_90037[15:0]}) < $signed({1'h0, sel_90104}) ? smod_90037[15:0] : sel_90104;
  assign umul_90299 = umul22b_16b_x_6b(array_index_89943, 6'h3d);
  assign add_90301 = {1'h0, umul_90105[21:2]} + 21'h00_0fb9;
  assign sel_90306 = $signed({1'h0, smod_90042[15:0]}) < $signed({1'h0, sel_90112}) ? smod_90042[15:0] : sel_90112;
  assign umul_90307 = umul22b_16b_x_6b(array_index_89949, 6'h3d);
  assign add_90309 = {1'h0, umul_90113[21:2]} + 21'h00_0fb9;
  assign sel_90314 = $signed({1'h0, smod_90047[15:0]}) < $signed({1'h0, sel_90120}) ? smod_90047[15:0] : sel_90120;
  assign umul_90315 = umul22b_16b_x_6b(array_index_90137, 6'h3b);
  assign add_90317 = {1'h0, umul_90121[21:1]} + 22'h00_1f59;
  assign sel_90322 = $signed({1'h0, smod_90052[15:0]}) < $signed({1'h0, sel_90128}) ? smod_90052[15:0] : sel_90128;
  assign umul_90323 = umul22b_16b_x_6b(array_index_90143, 6'h3b);
  assign add_90325 = {1'h0, umul_90129[21:1]} + 22'h00_1f59;
  assign sel_90330 = $signed({1'h0, smod_90057[15:0]}) < $signed({1'h0, sel_90136}) ? smod_90057[15:0] : sel_90136;
  assign array_index_90331 = set1_unflattened[6'h16];
  assign smod_90335 = $unsigned($signed({9'h000, add_90199, umul_90003[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_90337 = set2_unflattened[6'h16];
  assign smod_90341 = $unsigned($signed({9'h000, add_90207, umul_90011[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_90391 = umul22b_16b_x_6b(array_index_90331, 6'h35);
  assign add_90393 = {1'h0, umul_90197[21:7]} + 16'h007d;
  assign sel_90398 = $signed({1'h0, smod_90141[15:0]}) < $signed({1'h0, sel_90204}) ? smod_90141[15:0] : sel_90204;
  assign umul_90399 = umul22b_16b_x_6b(array_index_90337, 6'h35);
  assign add_90401 = {1'h0, umul_90205[21:7]} + 16'h007d;
  assign sel_90406 = $signed({1'h0, smod_90147[15:0]}) < $signed({1'h0, sel_90212}) ? smod_90147[15:0] : sel_90212;
  assign smod_90410 = $unsigned($signed({8'h00, add_90269, umul_90073[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_90415 = $unsigned($signed({8'h00, add_90277, umul_90081[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_90420 = $unsigned($signed({8'h00, add_90285, umul_90089[0]}) % $signed(32'h0000_3ffd));
  assign smod_90425 = $unsigned($signed({8'h00, add_90293, umul_90097[0]}) % $signed(32'h0000_3ffd));
  assign smod_90430 = $unsigned($signed({9'h000, add_90301, umul_90105[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_90435 = $unsigned($signed({9'h000, add_90309, umul_90113[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_90440 = $unsigned($signed({9'h000, add_90317, umul_90121[0]}) % $signed(32'h0000_3ffd));
  assign smod_90445 = $unsigned($signed({9'h000, add_90325, umul_90129[0]}) % $signed(32'h0000_3ffd));
  assign umul_90461 = umul23b_16b_x_7b(array_index_89749, 7'h49);
  assign add_90463 = {1'h0, umul_90267[22:3]} + 21'h00_07e9;
  assign sel_90468 = $signed({1'h0, smod_90216[15:0]}) < $signed({1'h0, sel_90274}) ? smod_90216[15:0] : sel_90274;
  assign umul_90469 = umul23b_16b_x_7b(array_index_89755, 7'h49);
  assign add_90471 = {1'h0, umul_90275[22:3]} + 21'h00_07e9;
  assign sel_90476 = $signed({1'h0, smod_90221[15:0]}) < $signed({1'h0, sel_90282}) ? smod_90221[15:0] : sel_90282;
  assign umul_90477 = umul23b_16b_x_7b(array_index_89943, 7'h47);
  assign add_90479 = {1'h0, umul_90283[22:1]} + 23'h00_1f8b;
  assign sel_90484 = $signed({1'h0, smod_90226[15:0]}) < $signed({1'h0, sel_90290}) ? smod_90226[15:0] : sel_90290;
  assign umul_90485 = umul23b_16b_x_7b(array_index_89949, 7'h47);
  assign add_90487 = {1'h0, umul_90291[22:1]} + 23'h00_1f8b;
  assign sel_90492 = $signed({1'h0, smod_90231[15:0]}) < $signed({1'h0, sel_90298}) ? smod_90231[15:0] : sel_90298;
  assign umul_90493 = umul22b_16b_x_6b(array_index_90137, 6'h3d);
  assign add_90495 = {1'h0, umul_90299[21:2]} + 21'h00_0fb9;
  assign sel_90500 = $signed({1'h0, smod_90236[15:0]}) < $signed({1'h0, sel_90306}) ? smod_90236[15:0] : sel_90306;
  assign umul_90501 = umul22b_16b_x_6b(array_index_90143, 6'h3d);
  assign add_90503 = {1'h0, umul_90307[21:2]} + 21'h00_0fb9;
  assign sel_90508 = $signed({1'h0, smod_90241[15:0]}) < $signed({1'h0, sel_90314}) ? smod_90241[15:0] : sel_90314;
  assign umul_90509 = umul22b_16b_x_6b(array_index_90331, 6'h3b);
  assign add_90511 = {1'h0, umul_90315[21:1]} + 22'h00_1f59;
  assign sel_90516 = $signed({1'h0, smod_90246[15:0]}) < $signed({1'h0, sel_90322}) ? smod_90246[15:0] : sel_90322;
  assign umul_90517 = umul22b_16b_x_6b(array_index_90337, 6'h3b);
  assign add_90519 = {1'h0, umul_90323[21:1]} + 22'h00_1f59;
  assign sel_90524 = $signed({1'h0, smod_90251[15:0]}) < $signed({1'h0, sel_90330}) ? smod_90251[15:0] : sel_90330;
  assign array_index_90525 = set1_unflattened[6'h17];
  assign smod_90529 = $unsigned($signed({9'h000, add_90393, umul_90197[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_90531 = set2_unflattened[6'h17];
  assign smod_90535 = $unsigned($signed({9'h000, add_90401, umul_90205[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_90585 = umul22b_16b_x_6b(array_index_90525, 6'h35);
  assign add_90587 = {1'h0, umul_90391[21:7]} + 16'h007d;
  assign sel_90592 = $signed({1'h0, smod_90335[15:0]}) < $signed({1'h0, sel_90398}) ? smod_90335[15:0] : sel_90398;
  assign umul_90593 = umul22b_16b_x_6b(array_index_90531, 6'h35);
  assign add_90595 = {1'h0, umul_90399[21:7]} + 16'h007d;
  assign sel_90600 = $signed({1'h0, smod_90341[15:0]}) < $signed({1'h0, sel_90406}) ? smod_90341[15:0] : sel_90406;
  assign smod_90604 = $unsigned($signed({8'h00, add_90463, umul_90267[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_90609 = $unsigned($signed({8'h00, add_90471, umul_90275[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_90614 = $unsigned($signed({8'h00, add_90479, umul_90283[0]}) % $signed(32'h0000_3ffd));
  assign smod_90619 = $unsigned($signed({8'h00, add_90487, umul_90291[0]}) % $signed(32'h0000_3ffd));
  assign smod_90624 = $unsigned($signed({9'h000, add_90495, umul_90299[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_90629 = $unsigned($signed({9'h000, add_90503, umul_90307[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_90634 = $unsigned($signed({9'h000, add_90511, umul_90315[0]}) % $signed(32'h0000_3ffd));
  assign smod_90639 = $unsigned($signed({9'h000, add_90519, umul_90323[0]}) % $signed(32'h0000_3ffd));
  assign umul_90655 = umul23b_16b_x_7b(array_index_89943, 7'h49);
  assign add_90657 = {1'h0, umul_90461[22:3]} + 21'h00_07e9;
  assign sel_90662 = $signed({1'h0, smod_90410[15:0]}) < $signed({1'h0, sel_90468}) ? smod_90410[15:0] : sel_90468;
  assign umul_90663 = umul23b_16b_x_7b(array_index_89949, 7'h49);
  assign add_90665 = {1'h0, umul_90469[22:3]} + 21'h00_07e9;
  assign sel_90670 = $signed({1'h0, smod_90415[15:0]}) < $signed({1'h0, sel_90476}) ? smod_90415[15:0] : sel_90476;
  assign umul_90671 = umul23b_16b_x_7b(array_index_90137, 7'h47);
  assign add_90673 = {1'h0, umul_90477[22:1]} + 23'h00_1f8b;
  assign sel_90678 = $signed({1'h0, smod_90420[15:0]}) < $signed({1'h0, sel_90484}) ? smod_90420[15:0] : sel_90484;
  assign umul_90679 = umul23b_16b_x_7b(array_index_90143, 7'h47);
  assign add_90681 = {1'h0, umul_90485[22:1]} + 23'h00_1f8b;
  assign sel_90686 = $signed({1'h0, smod_90425[15:0]}) < $signed({1'h0, sel_90492}) ? smod_90425[15:0] : sel_90492;
  assign umul_90687 = umul22b_16b_x_6b(array_index_90331, 6'h3d);
  assign add_90689 = {1'h0, umul_90493[21:2]} + 21'h00_0fb9;
  assign sel_90694 = $signed({1'h0, smod_90430[15:0]}) < $signed({1'h0, sel_90500}) ? smod_90430[15:0] : sel_90500;
  assign umul_90695 = umul22b_16b_x_6b(array_index_90337, 6'h3d);
  assign add_90697 = {1'h0, umul_90501[21:2]} + 21'h00_0fb9;
  assign sel_90702 = $signed({1'h0, smod_90435[15:0]}) < $signed({1'h0, sel_90508}) ? smod_90435[15:0] : sel_90508;
  assign umul_90703 = umul22b_16b_x_6b(array_index_90525, 6'h3b);
  assign add_90705 = {1'h0, umul_90509[21:1]} + 22'h00_1f59;
  assign sel_90710 = $signed({1'h0, smod_90440[15:0]}) < $signed({1'h0, sel_90516}) ? smod_90440[15:0] : sel_90516;
  assign umul_90711 = umul22b_16b_x_6b(array_index_90531, 6'h3b);
  assign add_90713 = {1'h0, umul_90517[21:1]} + 22'h00_1f59;
  assign sel_90718 = $signed({1'h0, smod_90445[15:0]}) < $signed({1'h0, sel_90524}) ? smod_90445[15:0] : sel_90524;
  assign array_index_90719 = set1_unflattened[6'h18];
  assign smod_90723 = $unsigned($signed({9'h000, add_90587, umul_90391[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_90725 = set2_unflattened[6'h18];
  assign smod_90729 = $unsigned($signed({9'h000, add_90595, umul_90399[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_90779 = umul22b_16b_x_6b(array_index_90719, 6'h35);
  assign add_90781 = {1'h0, umul_90585[21:7]} + 16'h007d;
  assign sel_90786 = $signed({1'h0, smod_90529[15:0]}) < $signed({1'h0, sel_90592}) ? smod_90529[15:0] : sel_90592;
  assign umul_90787 = umul22b_16b_x_6b(array_index_90725, 6'h35);
  assign add_90789 = {1'h0, umul_90593[21:7]} + 16'h007d;
  assign sel_90794 = $signed({1'h0, smod_90535[15:0]}) < $signed({1'h0, sel_90600}) ? smod_90535[15:0] : sel_90600;
  assign smod_90798 = $unsigned($signed({8'h00, add_90657, umul_90461[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_90803 = $unsigned($signed({8'h00, add_90665, umul_90469[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_90808 = $unsigned($signed({8'h00, add_90673, umul_90477[0]}) % $signed(32'h0000_3ffd));
  assign smod_90813 = $unsigned($signed({8'h00, add_90681, umul_90485[0]}) % $signed(32'h0000_3ffd));
  assign smod_90818 = $unsigned($signed({9'h000, add_90689, umul_90493[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_90823 = $unsigned($signed({9'h000, add_90697, umul_90501[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_90828 = $unsigned($signed({9'h000, add_90705, umul_90509[0]}) % $signed(32'h0000_3ffd));
  assign smod_90833 = $unsigned($signed({9'h000, add_90713, umul_90517[0]}) % $signed(32'h0000_3ffd));
  assign umul_90849 = umul23b_16b_x_7b(array_index_90137, 7'h49);
  assign add_90851 = {1'h0, umul_90655[22:3]} + 21'h00_07e9;
  assign sel_90856 = $signed({1'h0, smod_90604[15:0]}) < $signed({1'h0, sel_90662}) ? smod_90604[15:0] : sel_90662;
  assign umul_90857 = umul23b_16b_x_7b(array_index_90143, 7'h49);
  assign add_90859 = {1'h0, umul_90663[22:3]} + 21'h00_07e9;
  assign sel_90864 = $signed({1'h0, smod_90609[15:0]}) < $signed({1'h0, sel_90670}) ? smod_90609[15:0] : sel_90670;
  assign umul_90865 = umul23b_16b_x_7b(array_index_90331, 7'h47);
  assign add_90867 = {1'h0, umul_90671[22:1]} + 23'h00_1f8b;
  assign sel_90872 = $signed({1'h0, smod_90614[15:0]}) < $signed({1'h0, sel_90678}) ? smod_90614[15:0] : sel_90678;
  assign umul_90873 = umul23b_16b_x_7b(array_index_90337, 7'h47);
  assign add_90875 = {1'h0, umul_90679[22:1]} + 23'h00_1f8b;
  assign sel_90880 = $signed({1'h0, smod_90619[15:0]}) < $signed({1'h0, sel_90686}) ? smod_90619[15:0] : sel_90686;
  assign umul_90881 = umul22b_16b_x_6b(array_index_90525, 6'h3d);
  assign add_90883 = {1'h0, umul_90687[21:2]} + 21'h00_0fb9;
  assign sel_90888 = $signed({1'h0, smod_90624[15:0]}) < $signed({1'h0, sel_90694}) ? smod_90624[15:0] : sel_90694;
  assign umul_90889 = umul22b_16b_x_6b(array_index_90531, 6'h3d);
  assign add_90891 = {1'h0, umul_90695[21:2]} + 21'h00_0fb9;
  assign sel_90896 = $signed({1'h0, smod_90629[15:0]}) < $signed({1'h0, sel_90702}) ? smod_90629[15:0] : sel_90702;
  assign umul_90897 = umul22b_16b_x_6b(array_index_90719, 6'h3b);
  assign add_90899 = {1'h0, umul_90703[21:1]} + 22'h00_1f59;
  assign sel_90904 = $signed({1'h0, smod_90634[15:0]}) < $signed({1'h0, sel_90710}) ? smod_90634[15:0] : sel_90710;
  assign umul_90905 = umul22b_16b_x_6b(array_index_90725, 6'h3b);
  assign add_90907 = {1'h0, umul_90711[21:1]} + 22'h00_1f59;
  assign sel_90912 = $signed({1'h0, smod_90639[15:0]}) < $signed({1'h0, sel_90718}) ? smod_90639[15:0] : sel_90718;
  assign array_index_90913 = set1_unflattened[6'h19];
  assign smod_90917 = $unsigned($signed({9'h000, add_90781, umul_90585[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_90919 = set2_unflattened[6'h19];
  assign smod_90923 = $unsigned($signed({9'h000, add_90789, umul_90593[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_90973 = umul22b_16b_x_6b(array_index_90913, 6'h35);
  assign add_90975 = {1'h0, umul_90779[21:7]} + 16'h007d;
  assign sel_90980 = $signed({1'h0, smod_90723[15:0]}) < $signed({1'h0, sel_90786}) ? smod_90723[15:0] : sel_90786;
  assign umul_90981 = umul22b_16b_x_6b(array_index_90919, 6'h35);
  assign add_90983 = {1'h0, umul_90787[21:7]} + 16'h007d;
  assign sel_90988 = $signed({1'h0, smod_90729[15:0]}) < $signed({1'h0, sel_90794}) ? smod_90729[15:0] : sel_90794;
  assign smod_90992 = $unsigned($signed({8'h00, add_90851, umul_90655[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_90997 = $unsigned($signed({8'h00, add_90859, umul_90663[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_91002 = $unsigned($signed({8'h00, add_90867, umul_90671[0]}) % $signed(32'h0000_3ffd));
  assign smod_91007 = $unsigned($signed({8'h00, add_90875, umul_90679[0]}) % $signed(32'h0000_3ffd));
  assign smod_91012 = $unsigned($signed({9'h000, add_90883, umul_90687[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91017 = $unsigned($signed({9'h000, add_90891, umul_90695[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91022 = $unsigned($signed({9'h000, add_90899, umul_90703[0]}) % $signed(32'h0000_3ffd));
  assign smod_91027 = $unsigned($signed({9'h000, add_90907, umul_90711[0]}) % $signed(32'h0000_3ffd));
  assign umul_91043 = umul23b_16b_x_7b(array_index_90331, 7'h49);
  assign add_91045 = {1'h0, umul_90849[22:3]} + 21'h00_07e9;
  assign sel_91050 = $signed({1'h0, smod_90798[15:0]}) < $signed({1'h0, sel_90856}) ? smod_90798[15:0] : sel_90856;
  assign umul_91051 = umul23b_16b_x_7b(array_index_90337, 7'h49);
  assign add_91053 = {1'h0, umul_90857[22:3]} + 21'h00_07e9;
  assign sel_91058 = $signed({1'h0, smod_90803[15:0]}) < $signed({1'h0, sel_90864}) ? smod_90803[15:0] : sel_90864;
  assign umul_91059 = umul23b_16b_x_7b(array_index_90525, 7'h47);
  assign add_91061 = {1'h0, umul_90865[22:1]} + 23'h00_1f8b;
  assign sel_91066 = $signed({1'h0, smod_90808[15:0]}) < $signed({1'h0, sel_90872}) ? smod_90808[15:0] : sel_90872;
  assign umul_91067 = umul23b_16b_x_7b(array_index_90531, 7'h47);
  assign add_91069 = {1'h0, umul_90873[22:1]} + 23'h00_1f8b;
  assign sel_91074 = $signed({1'h0, smod_90813[15:0]}) < $signed({1'h0, sel_90880}) ? smod_90813[15:0] : sel_90880;
  assign umul_91075 = umul22b_16b_x_6b(array_index_90719, 6'h3d);
  assign add_91077 = {1'h0, umul_90881[21:2]} + 21'h00_0fb9;
  assign sel_91082 = $signed({1'h0, smod_90818[15:0]}) < $signed({1'h0, sel_90888}) ? smod_90818[15:0] : sel_90888;
  assign umul_91083 = umul22b_16b_x_6b(array_index_90725, 6'h3d);
  assign add_91085 = {1'h0, umul_90889[21:2]} + 21'h00_0fb9;
  assign sel_91090 = $signed({1'h0, smod_90823[15:0]}) < $signed({1'h0, sel_90896}) ? smod_90823[15:0] : sel_90896;
  assign umul_91091 = umul22b_16b_x_6b(array_index_90913, 6'h3b);
  assign add_91093 = {1'h0, umul_90897[21:1]} + 22'h00_1f59;
  assign sel_91098 = $signed({1'h0, smod_90828[15:0]}) < $signed({1'h0, sel_90904}) ? smod_90828[15:0] : sel_90904;
  assign umul_91099 = umul22b_16b_x_6b(array_index_90919, 6'h3b);
  assign add_91101 = {1'h0, umul_90905[21:1]} + 22'h00_1f59;
  assign sel_91106 = $signed({1'h0, smod_90833[15:0]}) < $signed({1'h0, sel_90912}) ? smod_90833[15:0] : sel_90912;
  assign array_index_91107 = set1_unflattened[6'h1a];
  assign smod_91111 = $unsigned($signed({9'h000, add_90975, umul_90779[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_91113 = set2_unflattened[6'h1a];
  assign smod_91117 = $unsigned($signed({9'h000, add_90983, umul_90787[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_91167 = umul22b_16b_x_6b(array_index_91107, 6'h35);
  assign add_91169 = {1'h0, umul_90973[21:7]} + 16'h007d;
  assign sel_91174 = $signed({1'h0, smod_90917[15:0]}) < $signed({1'h0, sel_90980}) ? smod_90917[15:0] : sel_90980;
  assign umul_91175 = umul22b_16b_x_6b(array_index_91113, 6'h35);
  assign add_91177 = {1'h0, umul_90981[21:7]} + 16'h007d;
  assign sel_91182 = $signed({1'h0, smod_90923[15:0]}) < $signed({1'h0, sel_90988}) ? smod_90923[15:0] : sel_90988;
  assign smod_91186 = $unsigned($signed({8'h00, add_91045, umul_90849[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_91191 = $unsigned($signed({8'h00, add_91053, umul_90857[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_91196 = $unsigned($signed({8'h00, add_91061, umul_90865[0]}) % $signed(32'h0000_3ffd));
  assign smod_91201 = $unsigned($signed({8'h00, add_91069, umul_90873[0]}) % $signed(32'h0000_3ffd));
  assign smod_91206 = $unsigned($signed({9'h000, add_91077, umul_90881[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91211 = $unsigned($signed({9'h000, add_91085, umul_90889[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91216 = $unsigned($signed({9'h000, add_91093, umul_90897[0]}) % $signed(32'h0000_3ffd));
  assign smod_91221 = $unsigned($signed({9'h000, add_91101, umul_90905[0]}) % $signed(32'h0000_3ffd));
  assign umul_91237 = umul23b_16b_x_7b(array_index_90525, 7'h49);
  assign add_91239 = {1'h0, umul_91043[22:3]} + 21'h00_07e9;
  assign sel_91244 = $signed({1'h0, smod_90992[15:0]}) < $signed({1'h0, sel_91050}) ? smod_90992[15:0] : sel_91050;
  assign umul_91245 = umul23b_16b_x_7b(array_index_90531, 7'h49);
  assign add_91247 = {1'h0, umul_91051[22:3]} + 21'h00_07e9;
  assign sel_91252 = $signed({1'h0, smod_90997[15:0]}) < $signed({1'h0, sel_91058}) ? smod_90997[15:0] : sel_91058;
  assign umul_91253 = umul23b_16b_x_7b(array_index_90719, 7'h47);
  assign add_91255 = {1'h0, umul_91059[22:1]} + 23'h00_1f8b;
  assign sel_91260 = $signed({1'h0, smod_91002[15:0]}) < $signed({1'h0, sel_91066}) ? smod_91002[15:0] : sel_91066;
  assign umul_91261 = umul23b_16b_x_7b(array_index_90725, 7'h47);
  assign add_91263 = {1'h0, umul_91067[22:1]} + 23'h00_1f8b;
  assign sel_91268 = $signed({1'h0, smod_91007[15:0]}) < $signed({1'h0, sel_91074}) ? smod_91007[15:0] : sel_91074;
  assign umul_91269 = umul22b_16b_x_6b(array_index_90913, 6'h3d);
  assign add_91271 = {1'h0, umul_91075[21:2]} + 21'h00_0fb9;
  assign sel_91276 = $signed({1'h0, smod_91012[15:0]}) < $signed({1'h0, sel_91082}) ? smod_91012[15:0] : sel_91082;
  assign umul_91277 = umul22b_16b_x_6b(array_index_90919, 6'h3d);
  assign add_91279 = {1'h0, umul_91083[21:2]} + 21'h00_0fb9;
  assign sel_91284 = $signed({1'h0, smod_91017[15:0]}) < $signed({1'h0, sel_91090}) ? smod_91017[15:0] : sel_91090;
  assign umul_91285 = umul22b_16b_x_6b(array_index_91107, 6'h3b);
  assign add_91287 = {1'h0, umul_91091[21:1]} + 22'h00_1f59;
  assign sel_91292 = $signed({1'h0, smod_91022[15:0]}) < $signed({1'h0, sel_91098}) ? smod_91022[15:0] : sel_91098;
  assign umul_91293 = umul22b_16b_x_6b(array_index_91113, 6'h3b);
  assign add_91295 = {1'h0, umul_91099[21:1]} + 22'h00_1f59;
  assign sel_91300 = $signed({1'h0, smod_91027[15:0]}) < $signed({1'h0, sel_91106}) ? smod_91027[15:0] : sel_91106;
  assign array_index_91301 = set1_unflattened[6'h1b];
  assign smod_91305 = $unsigned($signed({9'h000, add_91169, umul_90973[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_91307 = set2_unflattened[6'h1b];
  assign smod_91311 = $unsigned($signed({9'h000, add_91177, umul_90981[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_91361 = umul22b_16b_x_6b(array_index_91301, 6'h35);
  assign add_91363 = {1'h0, umul_91167[21:7]} + 16'h007d;
  assign sel_91368 = $signed({1'h0, smod_91111[15:0]}) < $signed({1'h0, sel_91174}) ? smod_91111[15:0] : sel_91174;
  assign umul_91369 = umul22b_16b_x_6b(array_index_91307, 6'h35);
  assign add_91371 = {1'h0, umul_91175[21:7]} + 16'h007d;
  assign sel_91376 = $signed({1'h0, smod_91117[15:0]}) < $signed({1'h0, sel_91182}) ? smod_91117[15:0] : sel_91182;
  assign smod_91380 = $unsigned($signed({8'h00, add_91239, umul_91043[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_91385 = $unsigned($signed({8'h00, add_91247, umul_91051[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_91390 = $unsigned($signed({8'h00, add_91255, umul_91059[0]}) % $signed(32'h0000_3ffd));
  assign smod_91395 = $unsigned($signed({8'h00, add_91263, umul_91067[0]}) % $signed(32'h0000_3ffd));
  assign smod_91400 = $unsigned($signed({9'h000, add_91271, umul_91075[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91405 = $unsigned($signed({9'h000, add_91279, umul_91083[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91410 = $unsigned($signed({9'h000, add_91287, umul_91091[0]}) % $signed(32'h0000_3ffd));
  assign smod_91415 = $unsigned($signed({9'h000, add_91295, umul_91099[0]}) % $signed(32'h0000_3ffd));
  assign umul_91431 = umul23b_16b_x_7b(array_index_90719, 7'h49);
  assign add_91433 = {1'h0, umul_91237[22:3]} + 21'h00_07e9;
  assign sel_91438 = $signed({1'h0, smod_91186[15:0]}) < $signed({1'h0, sel_91244}) ? smod_91186[15:0] : sel_91244;
  assign umul_91439 = umul23b_16b_x_7b(array_index_90725, 7'h49);
  assign add_91441 = {1'h0, umul_91245[22:3]} + 21'h00_07e9;
  assign sel_91446 = $signed({1'h0, smod_91191[15:0]}) < $signed({1'h0, sel_91252}) ? smod_91191[15:0] : sel_91252;
  assign umul_91447 = umul23b_16b_x_7b(array_index_90913, 7'h47);
  assign add_91449 = {1'h0, umul_91253[22:1]} + 23'h00_1f8b;
  assign sel_91454 = $signed({1'h0, smod_91196[15:0]}) < $signed({1'h0, sel_91260}) ? smod_91196[15:0] : sel_91260;
  assign umul_91455 = umul23b_16b_x_7b(array_index_90919, 7'h47);
  assign add_91457 = {1'h0, umul_91261[22:1]} + 23'h00_1f8b;
  assign sel_91462 = $signed({1'h0, smod_91201[15:0]}) < $signed({1'h0, sel_91268}) ? smod_91201[15:0] : sel_91268;
  assign umul_91463 = umul22b_16b_x_6b(array_index_91107, 6'h3d);
  assign add_91465 = {1'h0, umul_91269[21:2]} + 21'h00_0fb9;
  assign sel_91470 = $signed({1'h0, smod_91206[15:0]}) < $signed({1'h0, sel_91276}) ? smod_91206[15:0] : sel_91276;
  assign umul_91471 = umul22b_16b_x_6b(array_index_91113, 6'h3d);
  assign add_91473 = {1'h0, umul_91277[21:2]} + 21'h00_0fb9;
  assign sel_91478 = $signed({1'h0, smod_91211[15:0]}) < $signed({1'h0, sel_91284}) ? smod_91211[15:0] : sel_91284;
  assign umul_91479 = umul22b_16b_x_6b(array_index_91301, 6'h3b);
  assign add_91481 = {1'h0, umul_91285[21:1]} + 22'h00_1f59;
  assign sel_91486 = $signed({1'h0, smod_91216[15:0]}) < $signed({1'h0, sel_91292}) ? smod_91216[15:0] : sel_91292;
  assign umul_91487 = umul22b_16b_x_6b(array_index_91307, 6'h3b);
  assign add_91489 = {1'h0, umul_91293[21:1]} + 22'h00_1f59;
  assign sel_91494 = $signed({1'h0, smod_91221[15:0]}) < $signed({1'h0, sel_91300}) ? smod_91221[15:0] : sel_91300;
  assign array_index_91495 = set1_unflattened[6'h1c];
  assign smod_91499 = $unsigned($signed({9'h000, add_91363, umul_91167[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_91501 = set2_unflattened[6'h1c];
  assign smod_91505 = $unsigned($signed({9'h000, add_91371, umul_91175[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_91555 = umul22b_16b_x_6b(array_index_91495, 6'h35);
  assign add_91557 = {1'h0, umul_91361[21:7]} + 16'h007d;
  assign sel_91562 = $signed({1'h0, smod_91305[15:0]}) < $signed({1'h0, sel_91368}) ? smod_91305[15:0] : sel_91368;
  assign umul_91563 = umul22b_16b_x_6b(array_index_91501, 6'h35);
  assign add_91565 = {1'h0, umul_91369[21:7]} + 16'h007d;
  assign sel_91570 = $signed({1'h0, smod_91311[15:0]}) < $signed({1'h0, sel_91376}) ? smod_91311[15:0] : sel_91376;
  assign smod_91574 = $unsigned($signed({8'h00, add_91433, umul_91237[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_91579 = $unsigned($signed({8'h00, add_91441, umul_91245[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_91584 = $unsigned($signed({8'h00, add_91449, umul_91253[0]}) % $signed(32'h0000_3ffd));
  assign smod_91589 = $unsigned($signed({8'h00, add_91457, umul_91261[0]}) % $signed(32'h0000_3ffd));
  assign smod_91594 = $unsigned($signed({9'h000, add_91465, umul_91269[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91599 = $unsigned($signed({9'h000, add_91473, umul_91277[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91604 = $unsigned($signed({9'h000, add_91481, umul_91285[0]}) % $signed(32'h0000_3ffd));
  assign smod_91609 = $unsigned($signed({9'h000, add_91489, umul_91293[0]}) % $signed(32'h0000_3ffd));
  assign umul_91625 = umul23b_16b_x_7b(array_index_90913, 7'h49);
  assign add_91627 = {1'h0, umul_91431[22:3]} + 21'h00_07e9;
  assign sel_91632 = $signed({1'h0, smod_91380[15:0]}) < $signed({1'h0, sel_91438}) ? smod_91380[15:0] : sel_91438;
  assign umul_91633 = umul23b_16b_x_7b(array_index_90919, 7'h49);
  assign add_91635 = {1'h0, umul_91439[22:3]} + 21'h00_07e9;
  assign sel_91640 = $signed({1'h0, smod_91385[15:0]}) < $signed({1'h0, sel_91446}) ? smod_91385[15:0] : sel_91446;
  assign umul_91641 = umul23b_16b_x_7b(array_index_91107, 7'h47);
  assign add_91643 = {1'h0, umul_91447[22:1]} + 23'h00_1f8b;
  assign sel_91648 = $signed({1'h0, smod_91390[15:0]}) < $signed({1'h0, sel_91454}) ? smod_91390[15:0] : sel_91454;
  assign umul_91649 = umul23b_16b_x_7b(array_index_91113, 7'h47);
  assign add_91651 = {1'h0, umul_91455[22:1]} + 23'h00_1f8b;
  assign sel_91656 = $signed({1'h0, smod_91395[15:0]}) < $signed({1'h0, sel_91462}) ? smod_91395[15:0] : sel_91462;
  assign umul_91657 = umul22b_16b_x_6b(array_index_91301, 6'h3d);
  assign add_91659 = {1'h0, umul_91463[21:2]} + 21'h00_0fb9;
  assign sel_91664 = $signed({1'h0, smod_91400[15:0]}) < $signed({1'h0, sel_91470}) ? smod_91400[15:0] : sel_91470;
  assign umul_91665 = umul22b_16b_x_6b(array_index_91307, 6'h3d);
  assign add_91667 = {1'h0, umul_91471[21:2]} + 21'h00_0fb9;
  assign sel_91672 = $signed({1'h0, smod_91405[15:0]}) < $signed({1'h0, sel_91478}) ? smod_91405[15:0] : sel_91478;
  assign umul_91673 = umul22b_16b_x_6b(array_index_91495, 6'h3b);
  assign add_91675 = {1'h0, umul_91479[21:1]} + 22'h00_1f59;
  assign sel_91680 = $signed({1'h0, smod_91410[15:0]}) < $signed({1'h0, sel_91486}) ? smod_91410[15:0] : sel_91486;
  assign umul_91681 = umul22b_16b_x_6b(array_index_91501, 6'h3b);
  assign add_91683 = {1'h0, umul_91487[21:1]} + 22'h00_1f59;
  assign sel_91688 = $signed({1'h0, smod_91415[15:0]}) < $signed({1'h0, sel_91494}) ? smod_91415[15:0] : sel_91494;
  assign array_index_91689 = set1_unflattened[6'h1d];
  assign smod_91693 = $unsigned($signed({9'h000, add_91557, umul_91361[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_91695 = set2_unflattened[6'h1d];
  assign smod_91699 = $unsigned($signed({9'h000, add_91565, umul_91369[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_91749 = umul22b_16b_x_6b(array_index_91689, 6'h35);
  assign add_91751 = {1'h0, umul_91555[21:7]} + 16'h007d;
  assign sel_91756 = $signed({1'h0, smod_91499[15:0]}) < $signed({1'h0, sel_91562}) ? smod_91499[15:0] : sel_91562;
  assign umul_91757 = umul22b_16b_x_6b(array_index_91695, 6'h35);
  assign add_91759 = {1'h0, umul_91563[21:7]} + 16'h007d;
  assign sel_91764 = $signed({1'h0, smod_91505[15:0]}) < $signed({1'h0, sel_91570}) ? smod_91505[15:0] : sel_91570;
  assign smod_91768 = $unsigned($signed({8'h00, add_91627, umul_91431[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_91773 = $unsigned($signed({8'h00, add_91635, umul_91439[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_91778 = $unsigned($signed({8'h00, add_91643, umul_91447[0]}) % $signed(32'h0000_3ffd));
  assign smod_91783 = $unsigned($signed({8'h00, add_91651, umul_91455[0]}) % $signed(32'h0000_3ffd));
  assign smod_91788 = $unsigned($signed({9'h000, add_91659, umul_91463[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91793 = $unsigned($signed({9'h000, add_91667, umul_91471[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91798 = $unsigned($signed({9'h000, add_91675, umul_91479[0]}) % $signed(32'h0000_3ffd));
  assign smod_91803 = $unsigned($signed({9'h000, add_91683, umul_91487[0]}) % $signed(32'h0000_3ffd));
  assign umul_91819 = umul23b_16b_x_7b(array_index_91107, 7'h49);
  assign add_91821 = {1'h0, umul_91625[22:3]} + 21'h00_07e9;
  assign sel_91826 = $signed({1'h0, smod_91574[15:0]}) < $signed({1'h0, sel_91632}) ? smod_91574[15:0] : sel_91632;
  assign umul_91827 = umul23b_16b_x_7b(array_index_91113, 7'h49);
  assign add_91829 = {1'h0, umul_91633[22:3]} + 21'h00_07e9;
  assign sel_91834 = $signed({1'h0, smod_91579[15:0]}) < $signed({1'h0, sel_91640}) ? smod_91579[15:0] : sel_91640;
  assign umul_91835 = umul23b_16b_x_7b(array_index_91301, 7'h47);
  assign add_91837 = {1'h0, umul_91641[22:1]} + 23'h00_1f8b;
  assign sel_91842 = $signed({1'h0, smod_91584[15:0]}) < $signed({1'h0, sel_91648}) ? smod_91584[15:0] : sel_91648;
  assign umul_91843 = umul23b_16b_x_7b(array_index_91307, 7'h47);
  assign add_91845 = {1'h0, umul_91649[22:1]} + 23'h00_1f8b;
  assign sel_91850 = $signed({1'h0, smod_91589[15:0]}) < $signed({1'h0, sel_91656}) ? smod_91589[15:0] : sel_91656;
  assign umul_91851 = umul22b_16b_x_6b(array_index_91495, 6'h3d);
  assign add_91853 = {1'h0, umul_91657[21:2]} + 21'h00_0fb9;
  assign sel_91858 = $signed({1'h0, smod_91594[15:0]}) < $signed({1'h0, sel_91664}) ? smod_91594[15:0] : sel_91664;
  assign umul_91859 = umul22b_16b_x_6b(array_index_91501, 6'h3d);
  assign add_91861 = {1'h0, umul_91665[21:2]} + 21'h00_0fb9;
  assign sel_91866 = $signed({1'h0, smod_91599[15:0]}) < $signed({1'h0, sel_91672}) ? smod_91599[15:0] : sel_91672;
  assign umul_91867 = umul22b_16b_x_6b(array_index_91689, 6'h3b);
  assign add_91869 = {1'h0, umul_91673[21:1]} + 22'h00_1f59;
  assign sel_91874 = $signed({1'h0, smod_91604[15:0]}) < $signed({1'h0, sel_91680}) ? smod_91604[15:0] : sel_91680;
  assign umul_91875 = umul22b_16b_x_6b(array_index_91695, 6'h3b);
  assign add_91877 = {1'h0, umul_91681[21:1]} + 22'h00_1f59;
  assign sel_91882 = $signed({1'h0, smod_91609[15:0]}) < $signed({1'h0, sel_91688}) ? smod_91609[15:0] : sel_91688;
  assign array_index_91883 = set1_unflattened[6'h1e];
  assign smod_91887 = $unsigned($signed({9'h000, add_91751, umul_91555[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_91889 = set2_unflattened[6'h1e];
  assign smod_91893 = $unsigned($signed({9'h000, add_91759, umul_91563[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_91943 = umul22b_16b_x_6b(array_index_91883, 6'h35);
  assign add_91945 = {1'h0, umul_91749[21:7]} + 16'h007d;
  assign sel_91950 = $signed({1'h0, smod_91693[15:0]}) < $signed({1'h0, sel_91756}) ? smod_91693[15:0] : sel_91756;
  assign umul_91951 = umul22b_16b_x_6b(array_index_91889, 6'h35);
  assign add_91953 = {1'h0, umul_91757[21:7]} + 16'h007d;
  assign sel_91958 = $signed({1'h0, smod_91699[15:0]}) < $signed({1'h0, sel_91764}) ? smod_91699[15:0] : sel_91764;
  assign smod_91962 = $unsigned($signed({8'h00, add_91821, umul_91625[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_91967 = $unsigned($signed({8'h00, add_91829, umul_91633[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_91972 = $unsigned($signed({8'h00, add_91837, umul_91641[0]}) % $signed(32'h0000_3ffd));
  assign smod_91977 = $unsigned($signed({8'h00, add_91845, umul_91649[0]}) % $signed(32'h0000_3ffd));
  assign smod_91982 = $unsigned($signed({9'h000, add_91853, umul_91657[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91987 = $unsigned($signed({9'h000, add_91861, umul_91665[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_91992 = $unsigned($signed({9'h000, add_91869, umul_91673[0]}) % $signed(32'h0000_3ffd));
  assign smod_91997 = $unsigned($signed({9'h000, add_91877, umul_91681[0]}) % $signed(32'h0000_3ffd));
  assign umul_92013 = umul23b_16b_x_7b(array_index_91301, 7'h49);
  assign add_92015 = {1'h0, umul_91819[22:3]} + 21'h00_07e9;
  assign sel_92020 = $signed({1'h0, smod_91768[15:0]}) < $signed({1'h0, sel_91826}) ? smod_91768[15:0] : sel_91826;
  assign umul_92021 = umul23b_16b_x_7b(array_index_91307, 7'h49);
  assign add_92023 = {1'h0, umul_91827[22:3]} + 21'h00_07e9;
  assign sel_92028 = $signed({1'h0, smod_91773[15:0]}) < $signed({1'h0, sel_91834}) ? smod_91773[15:0] : sel_91834;
  assign umul_92029 = umul23b_16b_x_7b(array_index_91495, 7'h47);
  assign add_92031 = {1'h0, umul_91835[22:1]} + 23'h00_1f8b;
  assign sel_92036 = $signed({1'h0, smod_91778[15:0]}) < $signed({1'h0, sel_91842}) ? smod_91778[15:0] : sel_91842;
  assign umul_92037 = umul23b_16b_x_7b(array_index_91501, 7'h47);
  assign add_92039 = {1'h0, umul_91843[22:1]} + 23'h00_1f8b;
  assign sel_92044 = $signed({1'h0, smod_91783[15:0]}) < $signed({1'h0, sel_91850}) ? smod_91783[15:0] : sel_91850;
  assign umul_92045 = umul22b_16b_x_6b(array_index_91689, 6'h3d);
  assign add_92047 = {1'h0, umul_91851[21:2]} + 21'h00_0fb9;
  assign sel_92052 = $signed({1'h0, smod_91788[15:0]}) < $signed({1'h0, sel_91858}) ? smod_91788[15:0] : sel_91858;
  assign umul_92053 = umul22b_16b_x_6b(array_index_91695, 6'h3d);
  assign add_92055 = {1'h0, umul_91859[21:2]} + 21'h00_0fb9;
  assign sel_92060 = $signed({1'h0, smod_91793[15:0]}) < $signed({1'h0, sel_91866}) ? smod_91793[15:0] : sel_91866;
  assign umul_92061 = umul22b_16b_x_6b(array_index_91883, 6'h3b);
  assign add_92063 = {1'h0, umul_91867[21:1]} + 22'h00_1f59;
  assign sel_92068 = $signed({1'h0, smod_91798[15:0]}) < $signed({1'h0, sel_91874}) ? smod_91798[15:0] : sel_91874;
  assign umul_92069 = umul22b_16b_x_6b(array_index_91889, 6'h3b);
  assign add_92071 = {1'h0, umul_91875[21:1]} + 22'h00_1f59;
  assign sel_92076 = $signed({1'h0, smod_91803[15:0]}) < $signed({1'h0, sel_91882}) ? smod_91803[15:0] : sel_91882;
  assign array_index_92077 = set1_unflattened[6'h1f];
  assign smod_92081 = $unsigned($signed({9'h000, add_91945, umul_91749[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_92083 = set2_unflattened[6'h1f];
  assign smod_92087 = $unsigned($signed({9'h000, add_91953, umul_91757[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_92137 = umul22b_16b_x_6b(array_index_92077, 6'h35);
  assign add_92139 = {1'h0, umul_91943[21:7]} + 16'h007d;
  assign sel_92144 = $signed({1'h0, smod_91887[15:0]}) < $signed({1'h0, sel_91950}) ? smod_91887[15:0] : sel_91950;
  assign umul_92145 = umul22b_16b_x_6b(array_index_92083, 6'h35);
  assign add_92147 = {1'h0, umul_91951[21:7]} + 16'h007d;
  assign sel_92152 = $signed({1'h0, smod_91893[15:0]}) < $signed({1'h0, sel_91958}) ? smod_91893[15:0] : sel_91958;
  assign smod_92156 = $unsigned($signed({8'h00, add_92015, umul_91819[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_92161 = $unsigned($signed({8'h00, add_92023, umul_91827[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_92166 = $unsigned($signed({8'h00, add_92031, umul_91835[0]}) % $signed(32'h0000_3ffd));
  assign smod_92171 = $unsigned($signed({8'h00, add_92039, umul_91843[0]}) % $signed(32'h0000_3ffd));
  assign smod_92176 = $unsigned($signed({9'h000, add_92047, umul_91851[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_92181 = $unsigned($signed({9'h000, add_92055, umul_91859[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_92186 = $unsigned($signed({9'h000, add_92063, umul_91867[0]}) % $signed(32'h0000_3ffd));
  assign smod_92191 = $unsigned($signed({9'h000, add_92071, umul_91875[0]}) % $signed(32'h0000_3ffd));
  assign umul_92207 = umul23b_16b_x_7b(array_index_91495, 7'h49);
  assign add_92209 = {1'h0, umul_92013[22:3]} + 21'h00_07e9;
  assign sel_92214 = $signed({1'h0, smod_91962[15:0]}) < $signed({1'h0, sel_92020}) ? smod_91962[15:0] : sel_92020;
  assign umul_92215 = umul23b_16b_x_7b(array_index_91501, 7'h49);
  assign add_92217 = {1'h0, umul_92021[22:3]} + 21'h00_07e9;
  assign sel_92222 = $signed({1'h0, smod_91967[15:0]}) < $signed({1'h0, sel_92028}) ? smod_91967[15:0] : sel_92028;
  assign umul_92223 = umul23b_16b_x_7b(array_index_91689, 7'h47);
  assign add_92225 = {1'h0, umul_92029[22:1]} + 23'h00_1f8b;
  assign sel_92230 = $signed({1'h0, smod_91972[15:0]}) < $signed({1'h0, sel_92036}) ? smod_91972[15:0] : sel_92036;
  assign umul_92231 = umul23b_16b_x_7b(array_index_91695, 7'h47);
  assign add_92233 = {1'h0, umul_92037[22:1]} + 23'h00_1f8b;
  assign sel_92238 = $signed({1'h0, smod_91977[15:0]}) < $signed({1'h0, sel_92044}) ? smod_91977[15:0] : sel_92044;
  assign umul_92239 = umul22b_16b_x_6b(array_index_91883, 6'h3d);
  assign add_92241 = {1'h0, umul_92045[21:2]} + 21'h00_0fb9;
  assign sel_92246 = $signed({1'h0, smod_91982[15:0]}) < $signed({1'h0, sel_92052}) ? smod_91982[15:0] : sel_92052;
  assign umul_92247 = umul22b_16b_x_6b(array_index_91889, 6'h3d);
  assign add_92249 = {1'h0, umul_92053[21:2]} + 21'h00_0fb9;
  assign sel_92254 = $signed({1'h0, smod_91987[15:0]}) < $signed({1'h0, sel_92060}) ? smod_91987[15:0] : sel_92060;
  assign umul_92255 = umul22b_16b_x_6b(array_index_92077, 6'h3b);
  assign add_92257 = {1'h0, umul_92061[21:1]} + 22'h00_1f59;
  assign sel_92262 = $signed({1'h0, smod_91992[15:0]}) < $signed({1'h0, sel_92068}) ? smod_91992[15:0] : sel_92068;
  assign umul_92263 = umul22b_16b_x_6b(array_index_92083, 6'h3b);
  assign add_92265 = {1'h0, umul_92069[21:1]} + 22'h00_1f59;
  assign sel_92270 = $signed({1'h0, smod_91997[15:0]}) < $signed({1'h0, sel_92076}) ? smod_91997[15:0] : sel_92076;
  assign array_index_92271 = set1_unflattened[6'h20];
  assign smod_92275 = $unsigned($signed({9'h000, add_92139, umul_91943[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_92277 = set2_unflattened[6'h20];
  assign smod_92281 = $unsigned($signed({9'h000, add_92147, umul_91951[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_92331 = umul22b_16b_x_6b(array_index_92271, 6'h35);
  assign add_92333 = {1'h0, umul_92137[21:7]} + 16'h007d;
  assign sel_92338 = $signed({1'h0, smod_92081[15:0]}) < $signed({1'h0, sel_92144}) ? smod_92081[15:0] : sel_92144;
  assign umul_92339 = umul22b_16b_x_6b(array_index_92277, 6'h35);
  assign add_92341 = {1'h0, umul_92145[21:7]} + 16'h007d;
  assign sel_92346 = $signed({1'h0, smod_92087[15:0]}) < $signed({1'h0, sel_92152}) ? smod_92087[15:0] : sel_92152;
  assign smod_92350 = $unsigned($signed({8'h00, add_92209, umul_92013[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_92355 = $unsigned($signed({8'h00, add_92217, umul_92021[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_92360 = $unsigned($signed({8'h00, add_92225, umul_92029[0]}) % $signed(32'h0000_3ffd));
  assign smod_92365 = $unsigned($signed({8'h00, add_92233, umul_92037[0]}) % $signed(32'h0000_3ffd));
  assign smod_92370 = $unsigned($signed({9'h000, add_92241, umul_92045[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_92375 = $unsigned($signed({9'h000, add_92249, umul_92053[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_92380 = $unsigned($signed({9'h000, add_92257, umul_92061[0]}) % $signed(32'h0000_3ffd));
  assign smod_92385 = $unsigned($signed({9'h000, add_92265, umul_92069[0]}) % $signed(32'h0000_3ffd));
  assign umul_92401 = umul23b_16b_x_7b(array_index_91689, 7'h49);
  assign add_92403 = {1'h0, umul_92207[22:3]} + 21'h00_07e9;
  assign sel_92408 = $signed({1'h0, smod_92156[15:0]}) < $signed({1'h0, sel_92214}) ? smod_92156[15:0] : sel_92214;
  assign umul_92409 = umul23b_16b_x_7b(array_index_91695, 7'h49);
  assign add_92411 = {1'h0, umul_92215[22:3]} + 21'h00_07e9;
  assign sel_92416 = $signed({1'h0, smod_92161[15:0]}) < $signed({1'h0, sel_92222}) ? smod_92161[15:0] : sel_92222;
  assign umul_92417 = umul23b_16b_x_7b(array_index_91883, 7'h47);
  assign add_92419 = {1'h0, umul_92223[22:1]} + 23'h00_1f8b;
  assign sel_92424 = $signed({1'h0, smod_92166[15:0]}) < $signed({1'h0, sel_92230}) ? smod_92166[15:0] : sel_92230;
  assign umul_92425 = umul23b_16b_x_7b(array_index_91889, 7'h47);
  assign add_92427 = {1'h0, umul_92231[22:1]} + 23'h00_1f8b;
  assign sel_92432 = $signed({1'h0, smod_92171[15:0]}) < $signed({1'h0, sel_92238}) ? smod_92171[15:0] : sel_92238;
  assign umul_92433 = umul22b_16b_x_6b(array_index_92077, 6'h3d);
  assign add_92435 = {1'h0, umul_92239[21:2]} + 21'h00_0fb9;
  assign sel_92440 = $signed({1'h0, smod_92176[15:0]}) < $signed({1'h0, sel_92246}) ? smod_92176[15:0] : sel_92246;
  assign umul_92441 = umul22b_16b_x_6b(array_index_92083, 6'h3d);
  assign add_92443 = {1'h0, umul_92247[21:2]} + 21'h00_0fb9;
  assign sel_92448 = $signed({1'h0, smod_92181[15:0]}) < $signed({1'h0, sel_92254}) ? smod_92181[15:0] : sel_92254;
  assign umul_92449 = umul22b_16b_x_6b(array_index_92271, 6'h3b);
  assign add_92451 = {1'h0, umul_92255[21:1]} + 22'h00_1f59;
  assign sel_92456 = $signed({1'h0, smod_92186[15:0]}) < $signed({1'h0, sel_92262}) ? smod_92186[15:0] : sel_92262;
  assign umul_92457 = umul22b_16b_x_6b(array_index_92277, 6'h3b);
  assign add_92459 = {1'h0, umul_92263[21:1]} + 22'h00_1f59;
  assign sel_92464 = $signed({1'h0, smod_92191[15:0]}) < $signed({1'h0, sel_92270}) ? smod_92191[15:0] : sel_92270;
  assign array_index_92465 = set1_unflattened[6'h21];
  assign smod_92469 = $unsigned($signed({9'h000, add_92333, umul_92137[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_92471 = set2_unflattened[6'h21];
  assign smod_92475 = $unsigned($signed({9'h000, add_92341, umul_92145[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_92525 = umul22b_16b_x_6b(array_index_92465, 6'h35);
  assign add_92527 = {1'h0, umul_92331[21:7]} + 16'h007d;
  assign sel_92532 = $signed({1'h0, smod_92275[15:0]}) < $signed({1'h0, sel_92338}) ? smod_92275[15:0] : sel_92338;
  assign umul_92533 = umul22b_16b_x_6b(array_index_92471, 6'h35);
  assign add_92535 = {1'h0, umul_92339[21:7]} + 16'h007d;
  assign sel_92540 = $signed({1'h0, smod_92281[15:0]}) < $signed({1'h0, sel_92346}) ? smod_92281[15:0] : sel_92346;
  assign smod_92544 = $unsigned($signed({8'h00, add_92403, umul_92207[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_92549 = $unsigned($signed({8'h00, add_92411, umul_92215[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_92554 = $unsigned($signed({8'h00, add_92419, umul_92223[0]}) % $signed(32'h0000_3ffd));
  assign smod_92559 = $unsigned($signed({8'h00, add_92427, umul_92231[0]}) % $signed(32'h0000_3ffd));
  assign smod_92564 = $unsigned($signed({9'h000, add_92435, umul_92239[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_92569 = $unsigned($signed({9'h000, add_92443, umul_92247[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_92574 = $unsigned($signed({9'h000, add_92451, umul_92255[0]}) % $signed(32'h0000_3ffd));
  assign smod_92579 = $unsigned($signed({9'h000, add_92459, umul_92263[0]}) % $signed(32'h0000_3ffd));
  assign umul_92595 = umul23b_16b_x_7b(array_index_91883, 7'h49);
  assign add_92597 = {1'h0, umul_92401[22:3]} + 21'h00_07e9;
  assign sel_92602 = $signed({1'h0, smod_92350[15:0]}) < $signed({1'h0, sel_92408}) ? smod_92350[15:0] : sel_92408;
  assign umul_92603 = umul23b_16b_x_7b(array_index_91889, 7'h49);
  assign add_92605 = {1'h0, umul_92409[22:3]} + 21'h00_07e9;
  assign sel_92610 = $signed({1'h0, smod_92355[15:0]}) < $signed({1'h0, sel_92416}) ? smod_92355[15:0] : sel_92416;
  assign umul_92611 = umul23b_16b_x_7b(array_index_92077, 7'h47);
  assign add_92613 = {1'h0, umul_92417[22:1]} + 23'h00_1f8b;
  assign sel_92618 = $signed({1'h0, smod_92360[15:0]}) < $signed({1'h0, sel_92424}) ? smod_92360[15:0] : sel_92424;
  assign umul_92619 = umul23b_16b_x_7b(array_index_92083, 7'h47);
  assign add_92621 = {1'h0, umul_92425[22:1]} + 23'h00_1f8b;
  assign sel_92626 = $signed({1'h0, smod_92365[15:0]}) < $signed({1'h0, sel_92432}) ? smod_92365[15:0] : sel_92432;
  assign umul_92627 = umul22b_16b_x_6b(array_index_92271, 6'h3d);
  assign add_92629 = {1'h0, umul_92433[21:2]} + 21'h00_0fb9;
  assign sel_92634 = $signed({1'h0, smod_92370[15:0]}) < $signed({1'h0, sel_92440}) ? smod_92370[15:0] : sel_92440;
  assign umul_92635 = umul22b_16b_x_6b(array_index_92277, 6'h3d);
  assign add_92637 = {1'h0, umul_92441[21:2]} + 21'h00_0fb9;
  assign sel_92642 = $signed({1'h0, smod_92375[15:0]}) < $signed({1'h0, sel_92448}) ? smod_92375[15:0] : sel_92448;
  assign umul_92643 = umul22b_16b_x_6b(array_index_92465, 6'h3b);
  assign add_92645 = {1'h0, umul_92449[21:1]} + 22'h00_1f59;
  assign sel_92650 = $signed({1'h0, smod_92380[15:0]}) < $signed({1'h0, sel_92456}) ? smod_92380[15:0] : sel_92456;
  assign umul_92651 = umul22b_16b_x_6b(array_index_92471, 6'h3b);
  assign add_92653 = {1'h0, umul_92457[21:1]} + 22'h00_1f59;
  assign sel_92658 = $signed({1'h0, smod_92385[15:0]}) < $signed({1'h0, sel_92464}) ? smod_92385[15:0] : sel_92464;
  assign array_index_92659 = set1_unflattened[6'h22];
  assign smod_92663 = $unsigned($signed({9'h000, add_92527, umul_92331[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_92665 = set2_unflattened[6'h22];
  assign smod_92669 = $unsigned($signed({9'h000, add_92535, umul_92339[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_92719 = umul22b_16b_x_6b(array_index_92659, 6'h35);
  assign add_92721 = {1'h0, umul_92525[21:7]} + 16'h007d;
  assign sel_92726 = $signed({1'h0, smod_92469[15:0]}) < $signed({1'h0, sel_92532}) ? smod_92469[15:0] : sel_92532;
  assign umul_92727 = umul22b_16b_x_6b(array_index_92665, 6'h35);
  assign add_92729 = {1'h0, umul_92533[21:7]} + 16'h007d;
  assign sel_92734 = $signed({1'h0, smod_92475[15:0]}) < $signed({1'h0, sel_92540}) ? smod_92475[15:0] : sel_92540;
  assign smod_92738 = $unsigned($signed({8'h00, add_92597, umul_92401[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_92743 = $unsigned($signed({8'h00, add_92605, umul_92409[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_92748 = $unsigned($signed({8'h00, add_92613, umul_92417[0]}) % $signed(32'h0000_3ffd));
  assign smod_92753 = $unsigned($signed({8'h00, add_92621, umul_92425[0]}) % $signed(32'h0000_3ffd));
  assign smod_92758 = $unsigned($signed({9'h000, add_92629, umul_92433[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_92763 = $unsigned($signed({9'h000, add_92637, umul_92441[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_92768 = $unsigned($signed({9'h000, add_92645, umul_92449[0]}) % $signed(32'h0000_3ffd));
  assign smod_92773 = $unsigned($signed({9'h000, add_92653, umul_92457[0]}) % $signed(32'h0000_3ffd));
  assign umul_92789 = umul23b_16b_x_7b(array_index_92077, 7'h49);
  assign add_92791 = {1'h0, umul_92595[22:3]} + 21'h00_07e9;
  assign sel_92796 = $signed({1'h0, smod_92544[15:0]}) < $signed({1'h0, sel_92602}) ? smod_92544[15:0] : sel_92602;
  assign umul_92797 = umul23b_16b_x_7b(array_index_92083, 7'h49);
  assign add_92799 = {1'h0, umul_92603[22:3]} + 21'h00_07e9;
  assign sel_92804 = $signed({1'h0, smod_92549[15:0]}) < $signed({1'h0, sel_92610}) ? smod_92549[15:0] : sel_92610;
  assign umul_92805 = umul23b_16b_x_7b(array_index_92271, 7'h47);
  assign add_92807 = {1'h0, umul_92611[22:1]} + 23'h00_1f8b;
  assign sel_92812 = $signed({1'h0, smod_92554[15:0]}) < $signed({1'h0, sel_92618}) ? smod_92554[15:0] : sel_92618;
  assign umul_92813 = umul23b_16b_x_7b(array_index_92277, 7'h47);
  assign add_92815 = {1'h0, umul_92619[22:1]} + 23'h00_1f8b;
  assign sel_92820 = $signed({1'h0, smod_92559[15:0]}) < $signed({1'h0, sel_92626}) ? smod_92559[15:0] : sel_92626;
  assign umul_92821 = umul22b_16b_x_6b(array_index_92465, 6'h3d);
  assign add_92823 = {1'h0, umul_92627[21:2]} + 21'h00_0fb9;
  assign sel_92828 = $signed({1'h0, smod_92564[15:0]}) < $signed({1'h0, sel_92634}) ? smod_92564[15:0] : sel_92634;
  assign umul_92829 = umul22b_16b_x_6b(array_index_92471, 6'h3d);
  assign add_92831 = {1'h0, umul_92635[21:2]} + 21'h00_0fb9;
  assign sel_92836 = $signed({1'h0, smod_92569[15:0]}) < $signed({1'h0, sel_92642}) ? smod_92569[15:0] : sel_92642;
  assign umul_92837 = umul22b_16b_x_6b(array_index_92659, 6'h3b);
  assign add_92839 = {1'h0, umul_92643[21:1]} + 22'h00_1f59;
  assign sel_92844 = $signed({1'h0, smod_92574[15:0]}) < $signed({1'h0, sel_92650}) ? smod_92574[15:0] : sel_92650;
  assign umul_92845 = umul22b_16b_x_6b(array_index_92665, 6'h3b);
  assign add_92847 = {1'h0, umul_92651[21:1]} + 22'h00_1f59;
  assign sel_92852 = $signed({1'h0, smod_92579[15:0]}) < $signed({1'h0, sel_92658}) ? smod_92579[15:0] : sel_92658;
  assign array_index_92853 = set1_unflattened[6'h23];
  assign smod_92857 = $unsigned($signed({9'h000, add_92721, umul_92525[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_92859 = set2_unflattened[6'h23];
  assign smod_92863 = $unsigned($signed({9'h000, add_92729, umul_92533[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_92913 = umul22b_16b_x_6b(array_index_92853, 6'h35);
  assign add_92915 = {1'h0, umul_92719[21:7]} + 16'h007d;
  assign sel_92920 = $signed({1'h0, smod_92663[15:0]}) < $signed({1'h0, sel_92726}) ? smod_92663[15:0] : sel_92726;
  assign umul_92921 = umul22b_16b_x_6b(array_index_92859, 6'h35);
  assign add_92923 = {1'h0, umul_92727[21:7]} + 16'h007d;
  assign sel_92928 = $signed({1'h0, smod_92669[15:0]}) < $signed({1'h0, sel_92734}) ? smod_92669[15:0] : sel_92734;
  assign smod_92932 = $unsigned($signed({8'h00, add_92791, umul_92595[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_92937 = $unsigned($signed({8'h00, add_92799, umul_92603[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_92942 = $unsigned($signed({8'h00, add_92807, umul_92611[0]}) % $signed(32'h0000_3ffd));
  assign smod_92947 = $unsigned($signed({8'h00, add_92815, umul_92619[0]}) % $signed(32'h0000_3ffd));
  assign smod_92952 = $unsigned($signed({9'h000, add_92823, umul_92627[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_92957 = $unsigned($signed({9'h000, add_92831, umul_92635[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_92962 = $unsigned($signed({9'h000, add_92839, umul_92643[0]}) % $signed(32'h0000_3ffd));
  assign smod_92967 = $unsigned($signed({9'h000, add_92847, umul_92651[0]}) % $signed(32'h0000_3ffd));
  assign umul_92983 = umul23b_16b_x_7b(array_index_92271, 7'h49);
  assign add_92985 = {1'h0, umul_92789[22:3]} + 21'h00_07e9;
  assign sel_92990 = $signed({1'h0, smod_92738[15:0]}) < $signed({1'h0, sel_92796}) ? smod_92738[15:0] : sel_92796;
  assign umul_92991 = umul23b_16b_x_7b(array_index_92277, 7'h49);
  assign add_92993 = {1'h0, umul_92797[22:3]} + 21'h00_07e9;
  assign sel_92998 = $signed({1'h0, smod_92743[15:0]}) < $signed({1'h0, sel_92804}) ? smod_92743[15:0] : sel_92804;
  assign umul_92999 = umul23b_16b_x_7b(array_index_92465, 7'h47);
  assign add_93001 = {1'h0, umul_92805[22:1]} + 23'h00_1f8b;
  assign sel_93006 = $signed({1'h0, smod_92748[15:0]}) < $signed({1'h0, sel_92812}) ? smod_92748[15:0] : sel_92812;
  assign umul_93007 = umul23b_16b_x_7b(array_index_92471, 7'h47);
  assign add_93009 = {1'h0, umul_92813[22:1]} + 23'h00_1f8b;
  assign sel_93014 = $signed({1'h0, smod_92753[15:0]}) < $signed({1'h0, sel_92820}) ? smod_92753[15:0] : sel_92820;
  assign umul_93015 = umul22b_16b_x_6b(array_index_92659, 6'h3d);
  assign add_93017 = {1'h0, umul_92821[21:2]} + 21'h00_0fb9;
  assign sel_93022 = $signed({1'h0, smod_92758[15:0]}) < $signed({1'h0, sel_92828}) ? smod_92758[15:0] : sel_92828;
  assign umul_93023 = umul22b_16b_x_6b(array_index_92665, 6'h3d);
  assign add_93025 = {1'h0, umul_92829[21:2]} + 21'h00_0fb9;
  assign sel_93030 = $signed({1'h0, smod_92763[15:0]}) < $signed({1'h0, sel_92836}) ? smod_92763[15:0] : sel_92836;
  assign umul_93031 = umul22b_16b_x_6b(array_index_92853, 6'h3b);
  assign add_93033 = {1'h0, umul_92837[21:1]} + 22'h00_1f59;
  assign sel_93038 = $signed({1'h0, smod_92768[15:0]}) < $signed({1'h0, sel_92844}) ? smod_92768[15:0] : sel_92844;
  assign umul_93039 = umul22b_16b_x_6b(array_index_92859, 6'h3b);
  assign add_93041 = {1'h0, umul_92845[21:1]} + 22'h00_1f59;
  assign sel_93046 = $signed({1'h0, smod_92773[15:0]}) < $signed({1'h0, sel_92852}) ? smod_92773[15:0] : sel_92852;
  assign array_index_93047 = set1_unflattened[6'h24];
  assign smod_93051 = $unsigned($signed({9'h000, add_92915, umul_92719[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_93053 = set2_unflattened[6'h24];
  assign smod_93057 = $unsigned($signed({9'h000, add_92923, umul_92727[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_93107 = umul22b_16b_x_6b(array_index_93047, 6'h35);
  assign add_93109 = {1'h0, umul_92913[21:7]} + 16'h007d;
  assign sel_93114 = $signed({1'h0, smod_92857[15:0]}) < $signed({1'h0, sel_92920}) ? smod_92857[15:0] : sel_92920;
  assign umul_93115 = umul22b_16b_x_6b(array_index_93053, 6'h35);
  assign add_93117 = {1'h0, umul_92921[21:7]} + 16'h007d;
  assign sel_93122 = $signed({1'h0, smod_92863[15:0]}) < $signed({1'h0, sel_92928}) ? smod_92863[15:0] : sel_92928;
  assign smod_93126 = $unsigned($signed({8'h00, add_92985, umul_92789[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_93131 = $unsigned($signed({8'h00, add_92993, umul_92797[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_93136 = $unsigned($signed({8'h00, add_93001, umul_92805[0]}) % $signed(32'h0000_3ffd));
  assign smod_93141 = $unsigned($signed({8'h00, add_93009, umul_92813[0]}) % $signed(32'h0000_3ffd));
  assign smod_93146 = $unsigned($signed({9'h000, add_93017, umul_92821[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_93151 = $unsigned($signed({9'h000, add_93025, umul_92829[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_93156 = $unsigned($signed({9'h000, add_93033, umul_92837[0]}) % $signed(32'h0000_3ffd));
  assign smod_93161 = $unsigned($signed({9'h000, add_93041, umul_92845[0]}) % $signed(32'h0000_3ffd));
  assign umul_93177 = umul23b_16b_x_7b(array_index_92465, 7'h49);
  assign add_93179 = {1'h0, umul_92983[22:3]} + 21'h00_07e9;
  assign sel_93184 = $signed({1'h0, smod_92932[15:0]}) < $signed({1'h0, sel_92990}) ? smod_92932[15:0] : sel_92990;
  assign umul_93185 = umul23b_16b_x_7b(array_index_92471, 7'h49);
  assign add_93187 = {1'h0, umul_92991[22:3]} + 21'h00_07e9;
  assign sel_93192 = $signed({1'h0, smod_92937[15:0]}) < $signed({1'h0, sel_92998}) ? smod_92937[15:0] : sel_92998;
  assign umul_93193 = umul23b_16b_x_7b(array_index_92659, 7'h47);
  assign add_93195 = {1'h0, umul_92999[22:1]} + 23'h00_1f8b;
  assign sel_93200 = $signed({1'h0, smod_92942[15:0]}) < $signed({1'h0, sel_93006}) ? smod_92942[15:0] : sel_93006;
  assign umul_93201 = umul23b_16b_x_7b(array_index_92665, 7'h47);
  assign add_93203 = {1'h0, umul_93007[22:1]} + 23'h00_1f8b;
  assign sel_93208 = $signed({1'h0, smod_92947[15:0]}) < $signed({1'h0, sel_93014}) ? smod_92947[15:0] : sel_93014;
  assign umul_93209 = umul22b_16b_x_6b(array_index_92853, 6'h3d);
  assign add_93211 = {1'h0, umul_93015[21:2]} + 21'h00_0fb9;
  assign sel_93216 = $signed({1'h0, smod_92952[15:0]}) < $signed({1'h0, sel_93022}) ? smod_92952[15:0] : sel_93022;
  assign umul_93217 = umul22b_16b_x_6b(array_index_92859, 6'h3d);
  assign add_93219 = {1'h0, umul_93023[21:2]} + 21'h00_0fb9;
  assign sel_93224 = $signed({1'h0, smod_92957[15:0]}) < $signed({1'h0, sel_93030}) ? smod_92957[15:0] : sel_93030;
  assign umul_93225 = umul22b_16b_x_6b(array_index_93047, 6'h3b);
  assign add_93227 = {1'h0, umul_93031[21:1]} + 22'h00_1f59;
  assign sel_93232 = $signed({1'h0, smod_92962[15:0]}) < $signed({1'h0, sel_93038}) ? smod_92962[15:0] : sel_93038;
  assign umul_93233 = umul22b_16b_x_6b(array_index_93053, 6'h3b);
  assign add_93235 = {1'h0, umul_93039[21:1]} + 22'h00_1f59;
  assign sel_93240 = $signed({1'h0, smod_92967[15:0]}) < $signed({1'h0, sel_93046}) ? smod_92967[15:0] : sel_93046;
  assign array_index_93241 = set1_unflattened[6'h25];
  assign smod_93245 = $unsigned($signed({9'h000, add_93109, umul_92913[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_93247 = set2_unflattened[6'h25];
  assign smod_93251 = $unsigned($signed({9'h000, add_93117, umul_92921[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_93301 = umul22b_16b_x_6b(array_index_93241, 6'h35);
  assign add_93303 = {1'h0, umul_93107[21:7]} + 16'h007d;
  assign sel_93308 = $signed({1'h0, smod_93051[15:0]}) < $signed({1'h0, sel_93114}) ? smod_93051[15:0] : sel_93114;
  assign umul_93309 = umul22b_16b_x_6b(array_index_93247, 6'h35);
  assign add_93311 = {1'h0, umul_93115[21:7]} + 16'h007d;
  assign sel_93316 = $signed({1'h0, smod_93057[15:0]}) < $signed({1'h0, sel_93122}) ? smod_93057[15:0] : sel_93122;
  assign smod_93320 = $unsigned($signed({8'h00, add_93179, umul_92983[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_93325 = $unsigned($signed({8'h00, add_93187, umul_92991[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_93330 = $unsigned($signed({8'h00, add_93195, umul_92999[0]}) % $signed(32'h0000_3ffd));
  assign smod_93335 = $unsigned($signed({8'h00, add_93203, umul_93007[0]}) % $signed(32'h0000_3ffd));
  assign smod_93340 = $unsigned($signed({9'h000, add_93211, umul_93015[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_93345 = $unsigned($signed({9'h000, add_93219, umul_93023[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_93350 = $unsigned($signed({9'h000, add_93227, umul_93031[0]}) % $signed(32'h0000_3ffd));
  assign smod_93355 = $unsigned($signed({9'h000, add_93235, umul_93039[0]}) % $signed(32'h0000_3ffd));
  assign umul_93371 = umul23b_16b_x_7b(array_index_92659, 7'h49);
  assign add_93373 = {1'h0, umul_93177[22:3]} + 21'h00_07e9;
  assign sel_93378 = $signed({1'h0, smod_93126[15:0]}) < $signed({1'h0, sel_93184}) ? smod_93126[15:0] : sel_93184;
  assign umul_93379 = umul23b_16b_x_7b(array_index_92665, 7'h49);
  assign add_93381 = {1'h0, umul_93185[22:3]} + 21'h00_07e9;
  assign sel_93386 = $signed({1'h0, smod_93131[15:0]}) < $signed({1'h0, sel_93192}) ? smod_93131[15:0] : sel_93192;
  assign umul_93387 = umul23b_16b_x_7b(array_index_92853, 7'h47);
  assign add_93389 = {1'h0, umul_93193[22:1]} + 23'h00_1f8b;
  assign sel_93394 = $signed({1'h0, smod_93136[15:0]}) < $signed({1'h0, sel_93200}) ? smod_93136[15:0] : sel_93200;
  assign umul_93395 = umul23b_16b_x_7b(array_index_92859, 7'h47);
  assign add_93397 = {1'h0, umul_93201[22:1]} + 23'h00_1f8b;
  assign sel_93402 = $signed({1'h0, smod_93141[15:0]}) < $signed({1'h0, sel_93208}) ? smod_93141[15:0] : sel_93208;
  assign umul_93403 = umul22b_16b_x_6b(array_index_93047, 6'h3d);
  assign add_93405 = {1'h0, umul_93209[21:2]} + 21'h00_0fb9;
  assign sel_93410 = $signed({1'h0, smod_93146[15:0]}) < $signed({1'h0, sel_93216}) ? smod_93146[15:0] : sel_93216;
  assign umul_93411 = umul22b_16b_x_6b(array_index_93053, 6'h3d);
  assign add_93413 = {1'h0, umul_93217[21:2]} + 21'h00_0fb9;
  assign sel_93418 = $signed({1'h0, smod_93151[15:0]}) < $signed({1'h0, sel_93224}) ? smod_93151[15:0] : sel_93224;
  assign umul_93419 = umul22b_16b_x_6b(array_index_93241, 6'h3b);
  assign add_93421 = {1'h0, umul_93225[21:1]} + 22'h00_1f59;
  assign sel_93426 = $signed({1'h0, smod_93156[15:0]}) < $signed({1'h0, sel_93232}) ? smod_93156[15:0] : sel_93232;
  assign umul_93427 = umul22b_16b_x_6b(array_index_93247, 6'h3b);
  assign add_93429 = {1'h0, umul_93233[21:1]} + 22'h00_1f59;
  assign sel_93434 = $signed({1'h0, smod_93161[15:0]}) < $signed({1'h0, sel_93240}) ? smod_93161[15:0] : sel_93240;
  assign array_index_93435 = set1_unflattened[6'h26];
  assign smod_93439 = $unsigned($signed({9'h000, add_93303, umul_93107[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_93441 = set2_unflattened[6'h26];
  assign smod_93445 = $unsigned($signed({9'h000, add_93311, umul_93115[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_93495 = umul22b_16b_x_6b(array_index_93435, 6'h35);
  assign add_93497 = {1'h0, umul_93301[21:7]} + 16'h007d;
  assign sel_93502 = $signed({1'h0, smod_93245[15:0]}) < $signed({1'h0, sel_93308}) ? smod_93245[15:0] : sel_93308;
  assign umul_93503 = umul22b_16b_x_6b(array_index_93441, 6'h35);
  assign add_93505 = {1'h0, umul_93309[21:7]} + 16'h007d;
  assign sel_93510 = $signed({1'h0, smod_93251[15:0]}) < $signed({1'h0, sel_93316}) ? smod_93251[15:0] : sel_93316;
  assign smod_93514 = $unsigned($signed({8'h00, add_93373, umul_93177[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_93519 = $unsigned($signed({8'h00, add_93381, umul_93185[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_93524 = $unsigned($signed({8'h00, add_93389, umul_93193[0]}) % $signed(32'h0000_3ffd));
  assign smod_93529 = $unsigned($signed({8'h00, add_93397, umul_93201[0]}) % $signed(32'h0000_3ffd));
  assign smod_93534 = $unsigned($signed({9'h000, add_93405, umul_93209[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_93539 = $unsigned($signed({9'h000, add_93413, umul_93217[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_93544 = $unsigned($signed({9'h000, add_93421, umul_93225[0]}) % $signed(32'h0000_3ffd));
  assign smod_93549 = $unsigned($signed({9'h000, add_93429, umul_93233[0]}) % $signed(32'h0000_3ffd));
  assign umul_93565 = umul23b_16b_x_7b(array_index_92853, 7'h49);
  assign add_93567 = {1'h0, umul_93371[22:3]} + 21'h00_07e9;
  assign sel_93572 = $signed({1'h0, smod_93320[15:0]}) < $signed({1'h0, sel_93378}) ? smod_93320[15:0] : sel_93378;
  assign umul_93573 = umul23b_16b_x_7b(array_index_92859, 7'h49);
  assign add_93575 = {1'h0, umul_93379[22:3]} + 21'h00_07e9;
  assign sel_93580 = $signed({1'h0, smod_93325[15:0]}) < $signed({1'h0, sel_93386}) ? smod_93325[15:0] : sel_93386;
  assign umul_93581 = umul23b_16b_x_7b(array_index_93047, 7'h47);
  assign add_93583 = {1'h0, umul_93387[22:1]} + 23'h00_1f8b;
  assign sel_93588 = $signed({1'h0, smod_93330[15:0]}) < $signed({1'h0, sel_93394}) ? smod_93330[15:0] : sel_93394;
  assign umul_93589 = umul23b_16b_x_7b(array_index_93053, 7'h47);
  assign add_93591 = {1'h0, umul_93395[22:1]} + 23'h00_1f8b;
  assign sel_93596 = $signed({1'h0, smod_93335[15:0]}) < $signed({1'h0, sel_93402}) ? smod_93335[15:0] : sel_93402;
  assign umul_93597 = umul22b_16b_x_6b(array_index_93241, 6'h3d);
  assign add_93599 = {1'h0, umul_93403[21:2]} + 21'h00_0fb9;
  assign sel_93604 = $signed({1'h0, smod_93340[15:0]}) < $signed({1'h0, sel_93410}) ? smod_93340[15:0] : sel_93410;
  assign umul_93605 = umul22b_16b_x_6b(array_index_93247, 6'h3d);
  assign add_93607 = {1'h0, umul_93411[21:2]} + 21'h00_0fb9;
  assign sel_93612 = $signed({1'h0, smod_93345[15:0]}) < $signed({1'h0, sel_93418}) ? smod_93345[15:0] : sel_93418;
  assign umul_93613 = umul22b_16b_x_6b(array_index_93435, 6'h3b);
  assign add_93615 = {1'h0, umul_93419[21:1]} + 22'h00_1f59;
  assign sel_93620 = $signed({1'h0, smod_93350[15:0]}) < $signed({1'h0, sel_93426}) ? smod_93350[15:0] : sel_93426;
  assign umul_93621 = umul22b_16b_x_6b(array_index_93441, 6'h3b);
  assign add_93623 = {1'h0, umul_93427[21:1]} + 22'h00_1f59;
  assign sel_93628 = $signed({1'h0, smod_93355[15:0]}) < $signed({1'h0, sel_93434}) ? smod_93355[15:0] : sel_93434;
  assign array_index_93629 = set1_unflattened[6'h27];
  assign smod_93633 = $unsigned($signed({9'h000, add_93497, umul_93301[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_93635 = set2_unflattened[6'h27];
  assign smod_93639 = $unsigned($signed({9'h000, add_93505, umul_93309[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_93689 = umul22b_16b_x_6b(array_index_93629, 6'h35);
  assign add_93691 = {1'h0, umul_93495[21:7]} + 16'h007d;
  assign sel_93696 = $signed({1'h0, smod_93439[15:0]}) < $signed({1'h0, sel_93502}) ? smod_93439[15:0] : sel_93502;
  assign umul_93697 = umul22b_16b_x_6b(array_index_93635, 6'h35);
  assign add_93699 = {1'h0, umul_93503[21:7]} + 16'h007d;
  assign sel_93704 = $signed({1'h0, smod_93445[15:0]}) < $signed({1'h0, sel_93510}) ? smod_93445[15:0] : sel_93510;
  assign smod_93708 = $unsigned($signed({8'h00, add_93567, umul_93371[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_93713 = $unsigned($signed({8'h00, add_93575, umul_93379[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_93718 = $unsigned($signed({8'h00, add_93583, umul_93387[0]}) % $signed(32'h0000_3ffd));
  assign smod_93723 = $unsigned($signed({8'h00, add_93591, umul_93395[0]}) % $signed(32'h0000_3ffd));
  assign smod_93728 = $unsigned($signed({9'h000, add_93599, umul_93403[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_93733 = $unsigned($signed({9'h000, add_93607, umul_93411[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_93738 = $unsigned($signed({9'h000, add_93615, umul_93419[0]}) % $signed(32'h0000_3ffd));
  assign smod_93743 = $unsigned($signed({9'h000, add_93623, umul_93427[0]}) % $signed(32'h0000_3ffd));
  assign umul_93759 = umul23b_16b_x_7b(array_index_93047, 7'h49);
  assign add_93761 = {1'h0, umul_93565[22:3]} + 21'h00_07e9;
  assign sel_93766 = $signed({1'h0, smod_93514[15:0]}) < $signed({1'h0, sel_93572}) ? smod_93514[15:0] : sel_93572;
  assign umul_93767 = umul23b_16b_x_7b(array_index_93053, 7'h49);
  assign add_93769 = {1'h0, umul_93573[22:3]} + 21'h00_07e9;
  assign sel_93774 = $signed({1'h0, smod_93519[15:0]}) < $signed({1'h0, sel_93580}) ? smod_93519[15:0] : sel_93580;
  assign umul_93775 = umul23b_16b_x_7b(array_index_93241, 7'h47);
  assign add_93777 = {1'h0, umul_93581[22:1]} + 23'h00_1f8b;
  assign sel_93782 = $signed({1'h0, smod_93524[15:0]}) < $signed({1'h0, sel_93588}) ? smod_93524[15:0] : sel_93588;
  assign umul_93783 = umul23b_16b_x_7b(array_index_93247, 7'h47);
  assign add_93785 = {1'h0, umul_93589[22:1]} + 23'h00_1f8b;
  assign sel_93790 = $signed({1'h0, smod_93529[15:0]}) < $signed({1'h0, sel_93596}) ? smod_93529[15:0] : sel_93596;
  assign umul_93791 = umul22b_16b_x_6b(array_index_93435, 6'h3d);
  assign add_93793 = {1'h0, umul_93597[21:2]} + 21'h00_0fb9;
  assign sel_93798 = $signed({1'h0, smod_93534[15:0]}) < $signed({1'h0, sel_93604}) ? smod_93534[15:0] : sel_93604;
  assign umul_93799 = umul22b_16b_x_6b(array_index_93441, 6'h3d);
  assign add_93801 = {1'h0, umul_93605[21:2]} + 21'h00_0fb9;
  assign sel_93806 = $signed({1'h0, smod_93539[15:0]}) < $signed({1'h0, sel_93612}) ? smod_93539[15:0] : sel_93612;
  assign umul_93807 = umul22b_16b_x_6b(array_index_93629, 6'h3b);
  assign add_93809 = {1'h0, umul_93613[21:1]} + 22'h00_1f59;
  assign sel_93814 = $signed({1'h0, smod_93544[15:0]}) < $signed({1'h0, sel_93620}) ? smod_93544[15:0] : sel_93620;
  assign umul_93815 = umul22b_16b_x_6b(array_index_93635, 6'h3b);
  assign add_93817 = {1'h0, umul_93621[21:1]} + 22'h00_1f59;
  assign sel_93822 = $signed({1'h0, smod_93549[15:0]}) < $signed({1'h0, sel_93628}) ? smod_93549[15:0] : sel_93628;
  assign array_index_93823 = set1_unflattened[6'h28];
  assign smod_93827 = $unsigned($signed({9'h000, add_93691, umul_93495[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_93829 = set2_unflattened[6'h28];
  assign smod_93833 = $unsigned($signed({9'h000, add_93699, umul_93503[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_93883 = umul22b_16b_x_6b(array_index_93823, 6'h35);
  assign add_93885 = {1'h0, umul_93689[21:7]} + 16'h007d;
  assign sel_93890 = $signed({1'h0, smod_93633[15:0]}) < $signed({1'h0, sel_93696}) ? smod_93633[15:0] : sel_93696;
  assign umul_93891 = umul22b_16b_x_6b(array_index_93829, 6'h35);
  assign add_93893 = {1'h0, umul_93697[21:7]} + 16'h007d;
  assign sel_93898 = $signed({1'h0, smod_93639[15:0]}) < $signed({1'h0, sel_93704}) ? smod_93639[15:0] : sel_93704;
  assign smod_93902 = $unsigned($signed({8'h00, add_93761, umul_93565[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_93907 = $unsigned($signed({8'h00, add_93769, umul_93573[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_93912 = $unsigned($signed({8'h00, add_93777, umul_93581[0]}) % $signed(32'h0000_3ffd));
  assign smod_93917 = $unsigned($signed({8'h00, add_93785, umul_93589[0]}) % $signed(32'h0000_3ffd));
  assign smod_93922 = $unsigned($signed({9'h000, add_93793, umul_93597[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_93927 = $unsigned($signed({9'h000, add_93801, umul_93605[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_93932 = $unsigned($signed({9'h000, add_93809, umul_93613[0]}) % $signed(32'h0000_3ffd));
  assign smod_93937 = $unsigned($signed({9'h000, add_93817, umul_93621[0]}) % $signed(32'h0000_3ffd));
  assign umul_93953 = umul23b_16b_x_7b(array_index_93241, 7'h49);
  assign add_93955 = {1'h0, umul_93759[22:3]} + 21'h00_07e9;
  assign sel_93960 = $signed({1'h0, smod_93708[15:0]}) < $signed({1'h0, sel_93766}) ? smod_93708[15:0] : sel_93766;
  assign umul_93961 = umul23b_16b_x_7b(array_index_93247, 7'h49);
  assign add_93963 = {1'h0, umul_93767[22:3]} + 21'h00_07e9;
  assign sel_93968 = $signed({1'h0, smod_93713[15:0]}) < $signed({1'h0, sel_93774}) ? smod_93713[15:0] : sel_93774;
  assign umul_93969 = umul23b_16b_x_7b(array_index_93435, 7'h47);
  assign add_93971 = {1'h0, umul_93775[22:1]} + 23'h00_1f8b;
  assign sel_93976 = $signed({1'h0, smod_93718[15:0]}) < $signed({1'h0, sel_93782}) ? smod_93718[15:0] : sel_93782;
  assign umul_93977 = umul23b_16b_x_7b(array_index_93441, 7'h47);
  assign add_93979 = {1'h0, umul_93783[22:1]} + 23'h00_1f8b;
  assign sel_93984 = $signed({1'h0, smod_93723[15:0]}) < $signed({1'h0, sel_93790}) ? smod_93723[15:0] : sel_93790;
  assign umul_93985 = umul22b_16b_x_6b(array_index_93629, 6'h3d);
  assign add_93987 = {1'h0, umul_93791[21:2]} + 21'h00_0fb9;
  assign sel_93992 = $signed({1'h0, smod_93728[15:0]}) < $signed({1'h0, sel_93798}) ? smod_93728[15:0] : sel_93798;
  assign umul_93993 = umul22b_16b_x_6b(array_index_93635, 6'h3d);
  assign add_93995 = {1'h0, umul_93799[21:2]} + 21'h00_0fb9;
  assign sel_94000 = $signed({1'h0, smod_93733[15:0]}) < $signed({1'h0, sel_93806}) ? smod_93733[15:0] : sel_93806;
  assign umul_94001 = umul22b_16b_x_6b(array_index_93823, 6'h3b);
  assign add_94003 = {1'h0, umul_93807[21:1]} + 22'h00_1f59;
  assign sel_94008 = $signed({1'h0, smod_93738[15:0]}) < $signed({1'h0, sel_93814}) ? smod_93738[15:0] : sel_93814;
  assign umul_94009 = umul22b_16b_x_6b(array_index_93829, 6'h3b);
  assign add_94011 = {1'h0, umul_93815[21:1]} + 22'h00_1f59;
  assign sel_94016 = $signed({1'h0, smod_93743[15:0]}) < $signed({1'h0, sel_93822}) ? smod_93743[15:0] : sel_93822;
  assign array_index_94017 = set1_unflattened[6'h29];
  assign smod_94021 = $unsigned($signed({9'h000, add_93885, umul_93689[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_94023 = set2_unflattened[6'h29];
  assign smod_94027 = $unsigned($signed({9'h000, add_93893, umul_93697[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_94077 = umul22b_16b_x_6b(array_index_94017, 6'h35);
  assign add_94079 = {1'h0, umul_93883[21:7]} + 16'h007d;
  assign sel_94084 = $signed({1'h0, smod_93827[15:0]}) < $signed({1'h0, sel_93890}) ? smod_93827[15:0] : sel_93890;
  assign umul_94085 = umul22b_16b_x_6b(array_index_94023, 6'h35);
  assign add_94087 = {1'h0, umul_93891[21:7]} + 16'h007d;
  assign sel_94092 = $signed({1'h0, smod_93833[15:0]}) < $signed({1'h0, sel_93898}) ? smod_93833[15:0] : sel_93898;
  assign smod_94096 = $unsigned($signed({8'h00, add_93955, umul_93759[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_94101 = $unsigned($signed({8'h00, add_93963, umul_93767[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_94106 = $unsigned($signed({8'h00, add_93971, umul_93775[0]}) % $signed(32'h0000_3ffd));
  assign smod_94111 = $unsigned($signed({8'h00, add_93979, umul_93783[0]}) % $signed(32'h0000_3ffd));
  assign smod_94116 = $unsigned($signed({9'h000, add_93987, umul_93791[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_94121 = $unsigned($signed({9'h000, add_93995, umul_93799[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_94126 = $unsigned($signed({9'h000, add_94003, umul_93807[0]}) % $signed(32'h0000_3ffd));
  assign smod_94131 = $unsigned($signed({9'h000, add_94011, umul_93815[0]}) % $signed(32'h0000_3ffd));
  assign umul_94147 = umul23b_16b_x_7b(array_index_93435, 7'h49);
  assign add_94149 = {1'h0, umul_93953[22:3]} + 21'h00_07e9;
  assign sel_94154 = $signed({1'h0, smod_93902[15:0]}) < $signed({1'h0, sel_93960}) ? smod_93902[15:0] : sel_93960;
  assign umul_94155 = umul23b_16b_x_7b(array_index_93441, 7'h49);
  assign add_94157 = {1'h0, umul_93961[22:3]} + 21'h00_07e9;
  assign sel_94162 = $signed({1'h0, smod_93907[15:0]}) < $signed({1'h0, sel_93968}) ? smod_93907[15:0] : sel_93968;
  assign umul_94163 = umul23b_16b_x_7b(array_index_93629, 7'h47);
  assign add_94165 = {1'h0, umul_93969[22:1]} + 23'h00_1f8b;
  assign sel_94170 = $signed({1'h0, smod_93912[15:0]}) < $signed({1'h0, sel_93976}) ? smod_93912[15:0] : sel_93976;
  assign umul_94171 = umul23b_16b_x_7b(array_index_93635, 7'h47);
  assign add_94173 = {1'h0, umul_93977[22:1]} + 23'h00_1f8b;
  assign sel_94178 = $signed({1'h0, smod_93917[15:0]}) < $signed({1'h0, sel_93984}) ? smod_93917[15:0] : sel_93984;
  assign umul_94179 = umul22b_16b_x_6b(array_index_93823, 6'h3d);
  assign add_94181 = {1'h0, umul_93985[21:2]} + 21'h00_0fb9;
  assign sel_94186 = $signed({1'h0, smod_93922[15:0]}) < $signed({1'h0, sel_93992}) ? smod_93922[15:0] : sel_93992;
  assign umul_94187 = umul22b_16b_x_6b(array_index_93829, 6'h3d);
  assign add_94189 = {1'h0, umul_93993[21:2]} + 21'h00_0fb9;
  assign sel_94194 = $signed({1'h0, smod_93927[15:0]}) < $signed({1'h0, sel_94000}) ? smod_93927[15:0] : sel_94000;
  assign umul_94195 = umul22b_16b_x_6b(array_index_94017, 6'h3b);
  assign add_94197 = {1'h0, umul_94001[21:1]} + 22'h00_1f59;
  assign sel_94202 = $signed({1'h0, smod_93932[15:0]}) < $signed({1'h0, sel_94008}) ? smod_93932[15:0] : sel_94008;
  assign umul_94203 = umul22b_16b_x_6b(array_index_94023, 6'h3b);
  assign add_94205 = {1'h0, umul_94009[21:1]} + 22'h00_1f59;
  assign sel_94210 = $signed({1'h0, smod_93937[15:0]}) < $signed({1'h0, sel_94016}) ? smod_93937[15:0] : sel_94016;
  assign array_index_94211 = set1_unflattened[6'h2a];
  assign smod_94215 = $unsigned($signed({9'h000, add_94079, umul_93883[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_94217 = set2_unflattened[6'h2a];
  assign smod_94221 = $unsigned($signed({9'h000, add_94087, umul_93891[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_94271 = umul22b_16b_x_6b(array_index_94211, 6'h35);
  assign add_94273 = {1'h0, umul_94077[21:7]} + 16'h007d;
  assign sel_94278 = $signed({1'h0, smod_94021[15:0]}) < $signed({1'h0, sel_94084}) ? smod_94021[15:0] : sel_94084;
  assign umul_94279 = umul22b_16b_x_6b(array_index_94217, 6'h35);
  assign add_94281 = {1'h0, umul_94085[21:7]} + 16'h007d;
  assign sel_94286 = $signed({1'h0, smod_94027[15:0]}) < $signed({1'h0, sel_94092}) ? smod_94027[15:0] : sel_94092;
  assign smod_94290 = $unsigned($signed({8'h00, add_94149, umul_93953[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_94295 = $unsigned($signed({8'h00, add_94157, umul_93961[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_94300 = $unsigned($signed({8'h00, add_94165, umul_93969[0]}) % $signed(32'h0000_3ffd));
  assign smod_94305 = $unsigned($signed({8'h00, add_94173, umul_93977[0]}) % $signed(32'h0000_3ffd));
  assign smod_94310 = $unsigned($signed({9'h000, add_94181, umul_93985[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_94315 = $unsigned($signed({9'h000, add_94189, umul_93993[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_94320 = $unsigned($signed({9'h000, add_94197, umul_94001[0]}) % $signed(32'h0000_3ffd));
  assign smod_94325 = $unsigned($signed({9'h000, add_94205, umul_94009[0]}) % $signed(32'h0000_3ffd));
  assign umul_94341 = umul23b_16b_x_7b(array_index_93629, 7'h49);
  assign add_94343 = {1'h0, umul_94147[22:3]} + 21'h00_07e9;
  assign sel_94348 = $signed({1'h0, smod_94096[15:0]}) < $signed({1'h0, sel_94154}) ? smod_94096[15:0] : sel_94154;
  assign umul_94349 = umul23b_16b_x_7b(array_index_93635, 7'h49);
  assign add_94351 = {1'h0, umul_94155[22:3]} + 21'h00_07e9;
  assign sel_94356 = $signed({1'h0, smod_94101[15:0]}) < $signed({1'h0, sel_94162}) ? smod_94101[15:0] : sel_94162;
  assign umul_94357 = umul23b_16b_x_7b(array_index_93823, 7'h47);
  assign add_94359 = {1'h0, umul_94163[22:1]} + 23'h00_1f8b;
  assign sel_94364 = $signed({1'h0, smod_94106[15:0]}) < $signed({1'h0, sel_94170}) ? smod_94106[15:0] : sel_94170;
  assign umul_94365 = umul23b_16b_x_7b(array_index_93829, 7'h47);
  assign add_94367 = {1'h0, umul_94171[22:1]} + 23'h00_1f8b;
  assign sel_94372 = $signed({1'h0, smod_94111[15:0]}) < $signed({1'h0, sel_94178}) ? smod_94111[15:0] : sel_94178;
  assign umul_94373 = umul22b_16b_x_6b(array_index_94017, 6'h3d);
  assign add_94375 = {1'h0, umul_94179[21:2]} + 21'h00_0fb9;
  assign sel_94380 = $signed({1'h0, smod_94116[15:0]}) < $signed({1'h0, sel_94186}) ? smod_94116[15:0] : sel_94186;
  assign umul_94381 = umul22b_16b_x_6b(array_index_94023, 6'h3d);
  assign add_94383 = {1'h0, umul_94187[21:2]} + 21'h00_0fb9;
  assign sel_94388 = $signed({1'h0, smod_94121[15:0]}) < $signed({1'h0, sel_94194}) ? smod_94121[15:0] : sel_94194;
  assign umul_94389 = umul22b_16b_x_6b(array_index_94211, 6'h3b);
  assign add_94391 = {1'h0, umul_94195[21:1]} + 22'h00_1f59;
  assign sel_94396 = $signed({1'h0, smod_94126[15:0]}) < $signed({1'h0, sel_94202}) ? smod_94126[15:0] : sel_94202;
  assign umul_94397 = umul22b_16b_x_6b(array_index_94217, 6'h3b);
  assign add_94399 = {1'h0, umul_94203[21:1]} + 22'h00_1f59;
  assign sel_94404 = $signed({1'h0, smod_94131[15:0]}) < $signed({1'h0, sel_94210}) ? smod_94131[15:0] : sel_94210;
  assign array_index_94405 = set1_unflattened[6'h2b];
  assign smod_94409 = $unsigned($signed({9'h000, add_94273, umul_94077[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_94411 = set2_unflattened[6'h2b];
  assign smod_94415 = $unsigned($signed({9'h000, add_94281, umul_94085[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_94465 = umul22b_16b_x_6b(array_index_94405, 6'h35);
  assign add_94467 = {1'h0, umul_94271[21:7]} + 16'h007d;
  assign sel_94472 = $signed({1'h0, smod_94215[15:0]}) < $signed({1'h0, sel_94278}) ? smod_94215[15:0] : sel_94278;
  assign umul_94473 = umul22b_16b_x_6b(array_index_94411, 6'h35);
  assign add_94475 = {1'h0, umul_94279[21:7]} + 16'h007d;
  assign sel_94480 = $signed({1'h0, smod_94221[15:0]}) < $signed({1'h0, sel_94286}) ? smod_94221[15:0] : sel_94286;
  assign smod_94484 = $unsigned($signed({8'h00, add_94343, umul_94147[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_94489 = $unsigned($signed({8'h00, add_94351, umul_94155[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_94494 = $unsigned($signed({8'h00, add_94359, umul_94163[0]}) % $signed(32'h0000_3ffd));
  assign smod_94499 = $unsigned($signed({8'h00, add_94367, umul_94171[0]}) % $signed(32'h0000_3ffd));
  assign smod_94504 = $unsigned($signed({9'h000, add_94375, umul_94179[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_94509 = $unsigned($signed({9'h000, add_94383, umul_94187[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_94514 = $unsigned($signed({9'h000, add_94391, umul_94195[0]}) % $signed(32'h0000_3ffd));
  assign smod_94519 = $unsigned($signed({9'h000, add_94399, umul_94203[0]}) % $signed(32'h0000_3ffd));
  assign umul_94535 = umul23b_16b_x_7b(array_index_93823, 7'h49);
  assign add_94537 = {1'h0, umul_94341[22:3]} + 21'h00_07e9;
  assign sel_94542 = $signed({1'h0, smod_94290[15:0]}) < $signed({1'h0, sel_94348}) ? smod_94290[15:0] : sel_94348;
  assign umul_94543 = umul23b_16b_x_7b(array_index_93829, 7'h49);
  assign add_94545 = {1'h0, umul_94349[22:3]} + 21'h00_07e9;
  assign sel_94550 = $signed({1'h0, smod_94295[15:0]}) < $signed({1'h0, sel_94356}) ? smod_94295[15:0] : sel_94356;
  assign umul_94551 = umul23b_16b_x_7b(array_index_94017, 7'h47);
  assign add_94553 = {1'h0, umul_94357[22:1]} + 23'h00_1f8b;
  assign sel_94558 = $signed({1'h0, smod_94300[15:0]}) < $signed({1'h0, sel_94364}) ? smod_94300[15:0] : sel_94364;
  assign umul_94559 = umul23b_16b_x_7b(array_index_94023, 7'h47);
  assign add_94561 = {1'h0, umul_94365[22:1]} + 23'h00_1f8b;
  assign sel_94566 = $signed({1'h0, smod_94305[15:0]}) < $signed({1'h0, sel_94372}) ? smod_94305[15:0] : sel_94372;
  assign umul_94567 = umul22b_16b_x_6b(array_index_94211, 6'h3d);
  assign add_94569 = {1'h0, umul_94373[21:2]} + 21'h00_0fb9;
  assign sel_94574 = $signed({1'h0, smod_94310[15:0]}) < $signed({1'h0, sel_94380}) ? smod_94310[15:0] : sel_94380;
  assign umul_94575 = umul22b_16b_x_6b(array_index_94217, 6'h3d);
  assign add_94577 = {1'h0, umul_94381[21:2]} + 21'h00_0fb9;
  assign sel_94582 = $signed({1'h0, smod_94315[15:0]}) < $signed({1'h0, sel_94388}) ? smod_94315[15:0] : sel_94388;
  assign umul_94583 = umul22b_16b_x_6b(array_index_94405, 6'h3b);
  assign add_94585 = {1'h0, umul_94389[21:1]} + 22'h00_1f59;
  assign sel_94590 = $signed({1'h0, smod_94320[15:0]}) < $signed({1'h0, sel_94396}) ? smod_94320[15:0] : sel_94396;
  assign umul_94591 = umul22b_16b_x_6b(array_index_94411, 6'h3b);
  assign add_94593 = {1'h0, umul_94397[21:1]} + 22'h00_1f59;
  assign sel_94598 = $signed({1'h0, smod_94325[15:0]}) < $signed({1'h0, sel_94404}) ? smod_94325[15:0] : sel_94404;
  assign array_index_94599 = set1_unflattened[6'h2c];
  assign smod_94603 = $unsigned($signed({9'h000, add_94467, umul_94271[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_94605 = set2_unflattened[6'h2c];
  assign smod_94609 = $unsigned($signed({9'h000, add_94475, umul_94279[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_94659 = umul22b_16b_x_6b(array_index_94599, 6'h35);
  assign add_94661 = {1'h0, umul_94465[21:7]} + 16'h007d;
  assign sel_94666 = $signed({1'h0, smod_94409[15:0]}) < $signed({1'h0, sel_94472}) ? smod_94409[15:0] : sel_94472;
  assign umul_94667 = umul22b_16b_x_6b(array_index_94605, 6'h35);
  assign add_94669 = {1'h0, umul_94473[21:7]} + 16'h007d;
  assign sel_94674 = $signed({1'h0, smod_94415[15:0]}) < $signed({1'h0, sel_94480}) ? smod_94415[15:0] : sel_94480;
  assign smod_94678 = $unsigned($signed({8'h00, add_94537, umul_94341[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_94683 = $unsigned($signed({8'h00, add_94545, umul_94349[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_94688 = $unsigned($signed({8'h00, add_94553, umul_94357[0]}) % $signed(32'h0000_3ffd));
  assign smod_94693 = $unsigned($signed({8'h00, add_94561, umul_94365[0]}) % $signed(32'h0000_3ffd));
  assign smod_94698 = $unsigned($signed({9'h000, add_94569, umul_94373[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_94703 = $unsigned($signed({9'h000, add_94577, umul_94381[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_94708 = $unsigned($signed({9'h000, add_94585, umul_94389[0]}) % $signed(32'h0000_3ffd));
  assign smod_94713 = $unsigned($signed({9'h000, add_94593, umul_94397[0]}) % $signed(32'h0000_3ffd));
  assign umul_94729 = umul23b_16b_x_7b(array_index_94017, 7'h49);
  assign add_94731 = {1'h0, umul_94535[22:3]} + 21'h00_07e9;
  assign sel_94736 = $signed({1'h0, smod_94484[15:0]}) < $signed({1'h0, sel_94542}) ? smod_94484[15:0] : sel_94542;
  assign umul_94737 = umul23b_16b_x_7b(array_index_94023, 7'h49);
  assign add_94739 = {1'h0, umul_94543[22:3]} + 21'h00_07e9;
  assign sel_94744 = $signed({1'h0, smod_94489[15:0]}) < $signed({1'h0, sel_94550}) ? smod_94489[15:0] : sel_94550;
  assign umul_94745 = umul23b_16b_x_7b(array_index_94211, 7'h47);
  assign add_94747 = {1'h0, umul_94551[22:1]} + 23'h00_1f8b;
  assign sel_94752 = $signed({1'h0, smod_94494[15:0]}) < $signed({1'h0, sel_94558}) ? smod_94494[15:0] : sel_94558;
  assign umul_94753 = umul23b_16b_x_7b(array_index_94217, 7'h47);
  assign add_94755 = {1'h0, umul_94559[22:1]} + 23'h00_1f8b;
  assign sel_94760 = $signed({1'h0, smod_94499[15:0]}) < $signed({1'h0, sel_94566}) ? smod_94499[15:0] : sel_94566;
  assign umul_94761 = umul22b_16b_x_6b(array_index_94405, 6'h3d);
  assign add_94763 = {1'h0, umul_94567[21:2]} + 21'h00_0fb9;
  assign sel_94768 = $signed({1'h0, smod_94504[15:0]}) < $signed({1'h0, sel_94574}) ? smod_94504[15:0] : sel_94574;
  assign umul_94769 = umul22b_16b_x_6b(array_index_94411, 6'h3d);
  assign add_94771 = {1'h0, umul_94575[21:2]} + 21'h00_0fb9;
  assign sel_94776 = $signed({1'h0, smod_94509[15:0]}) < $signed({1'h0, sel_94582}) ? smod_94509[15:0] : sel_94582;
  assign umul_94777 = umul22b_16b_x_6b(array_index_94599, 6'h3b);
  assign add_94779 = {1'h0, umul_94583[21:1]} + 22'h00_1f59;
  assign sel_94784 = $signed({1'h0, smod_94514[15:0]}) < $signed({1'h0, sel_94590}) ? smod_94514[15:0] : sel_94590;
  assign umul_94785 = umul22b_16b_x_6b(array_index_94605, 6'h3b);
  assign add_94787 = {1'h0, umul_94591[21:1]} + 22'h00_1f59;
  assign sel_94792 = $signed({1'h0, smod_94519[15:0]}) < $signed({1'h0, sel_94598}) ? smod_94519[15:0] : sel_94598;
  assign array_index_94793 = set1_unflattened[6'h2d];
  assign smod_94797 = $unsigned($signed({9'h000, add_94661, umul_94465[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_94799 = set2_unflattened[6'h2d];
  assign smod_94803 = $unsigned($signed({9'h000, add_94669, umul_94473[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_94853 = umul22b_16b_x_6b(array_index_94793, 6'h35);
  assign add_94855 = {1'h0, umul_94659[21:7]} + 16'h007d;
  assign sel_94860 = $signed({1'h0, smod_94603[15:0]}) < $signed({1'h0, sel_94666}) ? smod_94603[15:0] : sel_94666;
  assign umul_94861 = umul22b_16b_x_6b(array_index_94799, 6'h35);
  assign add_94863 = {1'h0, umul_94667[21:7]} + 16'h007d;
  assign sel_94868 = $signed({1'h0, smod_94609[15:0]}) < $signed({1'h0, sel_94674}) ? smod_94609[15:0] : sel_94674;
  assign smod_94872 = $unsigned($signed({8'h00, add_94731, umul_94535[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_94877 = $unsigned($signed({8'h00, add_94739, umul_94543[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_94882 = $unsigned($signed({8'h00, add_94747, umul_94551[0]}) % $signed(32'h0000_3ffd));
  assign smod_94887 = $unsigned($signed({8'h00, add_94755, umul_94559[0]}) % $signed(32'h0000_3ffd));
  assign smod_94892 = $unsigned($signed({9'h000, add_94763, umul_94567[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_94897 = $unsigned($signed({9'h000, add_94771, umul_94575[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_94902 = $unsigned($signed({9'h000, add_94779, umul_94583[0]}) % $signed(32'h0000_3ffd));
  assign smod_94907 = $unsigned($signed({9'h000, add_94787, umul_94591[0]}) % $signed(32'h0000_3ffd));
  assign umul_94923 = umul23b_16b_x_7b(array_index_94211, 7'h49);
  assign add_94925 = {1'h0, umul_94729[22:3]} + 21'h00_07e9;
  assign sel_94930 = $signed({1'h0, smod_94678[15:0]}) < $signed({1'h0, sel_94736}) ? smod_94678[15:0] : sel_94736;
  assign umul_94931 = umul23b_16b_x_7b(array_index_94217, 7'h49);
  assign add_94933 = {1'h0, umul_94737[22:3]} + 21'h00_07e9;
  assign sel_94938 = $signed({1'h0, smod_94683[15:0]}) < $signed({1'h0, sel_94744}) ? smod_94683[15:0] : sel_94744;
  assign umul_94939 = umul23b_16b_x_7b(array_index_94405, 7'h47);
  assign add_94941 = {1'h0, umul_94745[22:1]} + 23'h00_1f8b;
  assign sel_94946 = $signed({1'h0, smod_94688[15:0]}) < $signed({1'h0, sel_94752}) ? smod_94688[15:0] : sel_94752;
  assign umul_94947 = umul23b_16b_x_7b(array_index_94411, 7'h47);
  assign add_94949 = {1'h0, umul_94753[22:1]} + 23'h00_1f8b;
  assign sel_94954 = $signed({1'h0, smod_94693[15:0]}) < $signed({1'h0, sel_94760}) ? smod_94693[15:0] : sel_94760;
  assign umul_94955 = umul22b_16b_x_6b(array_index_94599, 6'h3d);
  assign add_94957 = {1'h0, umul_94761[21:2]} + 21'h00_0fb9;
  assign sel_94962 = $signed({1'h0, smod_94698[15:0]}) < $signed({1'h0, sel_94768}) ? smod_94698[15:0] : sel_94768;
  assign umul_94963 = umul22b_16b_x_6b(array_index_94605, 6'h3d);
  assign add_94965 = {1'h0, umul_94769[21:2]} + 21'h00_0fb9;
  assign sel_94970 = $signed({1'h0, smod_94703[15:0]}) < $signed({1'h0, sel_94776}) ? smod_94703[15:0] : sel_94776;
  assign umul_94971 = umul22b_16b_x_6b(array_index_94793, 6'h3b);
  assign add_94973 = {1'h0, umul_94777[21:1]} + 22'h00_1f59;
  assign sel_94978 = $signed({1'h0, smod_94708[15:0]}) < $signed({1'h0, sel_94784}) ? smod_94708[15:0] : sel_94784;
  assign umul_94979 = umul22b_16b_x_6b(array_index_94799, 6'h3b);
  assign add_94981 = {1'h0, umul_94785[21:1]} + 22'h00_1f59;
  assign sel_94986 = $signed({1'h0, smod_94713[15:0]}) < $signed({1'h0, sel_94792}) ? smod_94713[15:0] : sel_94792;
  assign array_index_94987 = set1_unflattened[6'h2e];
  assign smod_94991 = $unsigned($signed({9'h000, add_94855, umul_94659[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_94993 = set2_unflattened[6'h2e];
  assign smod_94997 = $unsigned($signed({9'h000, add_94863, umul_94667[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_95047 = umul22b_16b_x_6b(array_index_94987, 6'h35);
  assign add_95049 = {1'h0, umul_94853[21:7]} + 16'h007d;
  assign sel_95054 = $signed({1'h0, smod_94797[15:0]}) < $signed({1'h0, sel_94860}) ? smod_94797[15:0] : sel_94860;
  assign umul_95055 = umul22b_16b_x_6b(array_index_94993, 6'h35);
  assign add_95057 = {1'h0, umul_94861[21:7]} + 16'h007d;
  assign sel_95062 = $signed({1'h0, smod_94803[15:0]}) < $signed({1'h0, sel_94868}) ? smod_94803[15:0] : sel_94868;
  assign smod_95066 = $unsigned($signed({8'h00, add_94925, umul_94729[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_95071 = $unsigned($signed({8'h00, add_94933, umul_94737[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_95076 = $unsigned($signed({8'h00, add_94941, umul_94745[0]}) % $signed(32'h0000_3ffd));
  assign smod_95081 = $unsigned($signed({8'h00, add_94949, umul_94753[0]}) % $signed(32'h0000_3ffd));
  assign smod_95086 = $unsigned($signed({9'h000, add_94957, umul_94761[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_95091 = $unsigned($signed({9'h000, add_94965, umul_94769[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_95096 = $unsigned($signed({9'h000, add_94973, umul_94777[0]}) % $signed(32'h0000_3ffd));
  assign smod_95101 = $unsigned($signed({9'h000, add_94981, umul_94785[0]}) % $signed(32'h0000_3ffd));
  assign umul_95117 = umul23b_16b_x_7b(array_index_94405, 7'h49);
  assign add_95119 = {1'h0, umul_94923[22:3]} + 21'h00_07e9;
  assign sel_95124 = $signed({1'h0, smod_94872[15:0]}) < $signed({1'h0, sel_94930}) ? smod_94872[15:0] : sel_94930;
  assign umul_95125 = umul23b_16b_x_7b(array_index_94411, 7'h49);
  assign add_95127 = {1'h0, umul_94931[22:3]} + 21'h00_07e9;
  assign sel_95132 = $signed({1'h0, smod_94877[15:0]}) < $signed({1'h0, sel_94938}) ? smod_94877[15:0] : sel_94938;
  assign umul_95133 = umul23b_16b_x_7b(array_index_94599, 7'h47);
  assign add_95135 = {1'h0, umul_94939[22:1]} + 23'h00_1f8b;
  assign sel_95140 = $signed({1'h0, smod_94882[15:0]}) < $signed({1'h0, sel_94946}) ? smod_94882[15:0] : sel_94946;
  assign umul_95141 = umul23b_16b_x_7b(array_index_94605, 7'h47);
  assign add_95143 = {1'h0, umul_94947[22:1]} + 23'h00_1f8b;
  assign sel_95148 = $signed({1'h0, smod_94887[15:0]}) < $signed({1'h0, sel_94954}) ? smod_94887[15:0] : sel_94954;
  assign umul_95149 = umul22b_16b_x_6b(array_index_94793, 6'h3d);
  assign add_95151 = {1'h0, umul_94955[21:2]} + 21'h00_0fb9;
  assign sel_95156 = $signed({1'h0, smod_94892[15:0]}) < $signed({1'h0, sel_94962}) ? smod_94892[15:0] : sel_94962;
  assign umul_95157 = umul22b_16b_x_6b(array_index_94799, 6'h3d);
  assign add_95159 = {1'h0, umul_94963[21:2]} + 21'h00_0fb9;
  assign sel_95164 = $signed({1'h0, smod_94897[15:0]}) < $signed({1'h0, sel_94970}) ? smod_94897[15:0] : sel_94970;
  assign umul_95165 = umul22b_16b_x_6b(array_index_94987, 6'h3b);
  assign add_95167 = {1'h0, umul_94971[21:1]} + 22'h00_1f59;
  assign sel_95172 = $signed({1'h0, smod_94902[15:0]}) < $signed({1'h0, sel_94978}) ? smod_94902[15:0] : sel_94978;
  assign umul_95173 = umul22b_16b_x_6b(array_index_94993, 6'h3b);
  assign add_95175 = {1'h0, umul_94979[21:1]} + 22'h00_1f59;
  assign sel_95180 = $signed({1'h0, smod_94907[15:0]}) < $signed({1'h0, sel_94986}) ? smod_94907[15:0] : sel_94986;
  assign array_index_95181 = set1_unflattened[6'h2f];
  assign smod_95185 = $unsigned($signed({9'h000, add_95049, umul_94853[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_95187 = set2_unflattened[6'h2f];
  assign smod_95191 = $unsigned($signed({9'h000, add_95057, umul_94861[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_95241 = umul22b_16b_x_6b(array_index_95181, 6'h35);
  assign add_95243 = {1'h0, umul_95047[21:7]} + 16'h007d;
  assign sel_95248 = $signed({1'h0, smod_94991[15:0]}) < $signed({1'h0, sel_95054}) ? smod_94991[15:0] : sel_95054;
  assign umul_95249 = umul22b_16b_x_6b(array_index_95187, 6'h35);
  assign add_95251 = {1'h0, umul_95055[21:7]} + 16'h007d;
  assign sel_95256 = $signed({1'h0, smod_94997[15:0]}) < $signed({1'h0, sel_95062}) ? smod_94997[15:0] : sel_95062;
  assign smod_95260 = $unsigned($signed({8'h00, add_95119, umul_94923[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_95265 = $unsigned($signed({8'h00, add_95127, umul_94931[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_95270 = $unsigned($signed({8'h00, add_95135, umul_94939[0]}) % $signed(32'h0000_3ffd));
  assign smod_95275 = $unsigned($signed({8'h00, add_95143, umul_94947[0]}) % $signed(32'h0000_3ffd));
  assign smod_95280 = $unsigned($signed({9'h000, add_95151, umul_94955[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_95285 = $unsigned($signed({9'h000, add_95159, umul_94963[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_95290 = $unsigned($signed({9'h000, add_95167, umul_94971[0]}) % $signed(32'h0000_3ffd));
  assign smod_95295 = $unsigned($signed({9'h000, add_95175, umul_94979[0]}) % $signed(32'h0000_3ffd));
  assign umul_95311 = umul23b_16b_x_7b(array_index_94599, 7'h49);
  assign add_95313 = {1'h0, umul_95117[22:3]} + 21'h00_07e9;
  assign sel_95318 = $signed({1'h0, smod_95066[15:0]}) < $signed({1'h0, sel_95124}) ? smod_95066[15:0] : sel_95124;
  assign umul_95319 = umul23b_16b_x_7b(array_index_94605, 7'h49);
  assign add_95321 = {1'h0, umul_95125[22:3]} + 21'h00_07e9;
  assign sel_95326 = $signed({1'h0, smod_95071[15:0]}) < $signed({1'h0, sel_95132}) ? smod_95071[15:0] : sel_95132;
  assign umul_95327 = umul23b_16b_x_7b(array_index_94793, 7'h47);
  assign add_95329 = {1'h0, umul_95133[22:1]} + 23'h00_1f8b;
  assign sel_95334 = $signed({1'h0, smod_95076[15:0]}) < $signed({1'h0, sel_95140}) ? smod_95076[15:0] : sel_95140;
  assign umul_95335 = umul23b_16b_x_7b(array_index_94799, 7'h47);
  assign add_95337 = {1'h0, umul_95141[22:1]} + 23'h00_1f8b;
  assign sel_95342 = $signed({1'h0, smod_95081[15:0]}) < $signed({1'h0, sel_95148}) ? smod_95081[15:0] : sel_95148;
  assign umul_95343 = umul22b_16b_x_6b(array_index_94987, 6'h3d);
  assign add_95345 = {1'h0, umul_95149[21:2]} + 21'h00_0fb9;
  assign sel_95350 = $signed({1'h0, smod_95086[15:0]}) < $signed({1'h0, sel_95156}) ? smod_95086[15:0] : sel_95156;
  assign umul_95351 = umul22b_16b_x_6b(array_index_94993, 6'h3d);
  assign add_95353 = {1'h0, umul_95157[21:2]} + 21'h00_0fb9;
  assign sel_95358 = $signed({1'h0, smod_95091[15:0]}) < $signed({1'h0, sel_95164}) ? smod_95091[15:0] : sel_95164;
  assign umul_95359 = umul22b_16b_x_6b(array_index_95181, 6'h3b);
  assign add_95361 = {1'h0, umul_95165[21:1]} + 22'h00_1f59;
  assign sel_95366 = $signed({1'h0, smod_95096[15:0]}) < $signed({1'h0, sel_95172}) ? smod_95096[15:0] : sel_95172;
  assign umul_95367 = umul22b_16b_x_6b(array_index_95187, 6'h3b);
  assign add_95369 = {1'h0, umul_95173[21:1]} + 22'h00_1f59;
  assign sel_95374 = $signed({1'h0, smod_95101[15:0]}) < $signed({1'h0, sel_95180}) ? smod_95101[15:0] : sel_95180;
  assign array_index_95375 = set1_unflattened[6'h30];
  assign smod_95379 = $unsigned($signed({9'h000, add_95243, umul_95047[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_95381 = set2_unflattened[6'h30];
  assign smod_95385 = $unsigned($signed({9'h000, add_95251, umul_95055[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_95435 = umul22b_16b_x_6b(array_index_95375, 6'h35);
  assign add_95437 = {1'h0, umul_95241[21:7]} + 16'h007d;
  assign sel_95442 = $signed({1'h0, smod_95185[15:0]}) < $signed({1'h0, sel_95248}) ? smod_95185[15:0] : sel_95248;
  assign umul_95443 = umul22b_16b_x_6b(array_index_95381, 6'h35);
  assign add_95445 = {1'h0, umul_95249[21:7]} + 16'h007d;
  assign sel_95450 = $signed({1'h0, smod_95191[15:0]}) < $signed({1'h0, sel_95256}) ? smod_95191[15:0] : sel_95256;
  assign smod_95454 = $unsigned($signed({8'h00, add_95313, umul_95117[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_95459 = $unsigned($signed({8'h00, add_95321, umul_95125[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_95464 = $unsigned($signed({8'h00, add_95329, umul_95133[0]}) % $signed(32'h0000_3ffd));
  assign smod_95469 = $unsigned($signed({8'h00, add_95337, umul_95141[0]}) % $signed(32'h0000_3ffd));
  assign smod_95474 = $unsigned($signed({9'h000, add_95345, umul_95149[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_95479 = $unsigned($signed({9'h000, add_95353, umul_95157[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_95484 = $unsigned($signed({9'h000, add_95361, umul_95165[0]}) % $signed(32'h0000_3ffd));
  assign smod_95489 = $unsigned($signed({9'h000, add_95369, umul_95173[0]}) % $signed(32'h0000_3ffd));
  assign umul_95505 = umul23b_16b_x_7b(array_index_94793, 7'h49);
  assign add_95507 = {1'h0, umul_95311[22:3]} + 21'h00_07e9;
  assign sel_95512 = $signed({1'h0, smod_95260[15:0]}) < $signed({1'h0, sel_95318}) ? smod_95260[15:0] : sel_95318;
  assign umul_95513 = umul23b_16b_x_7b(array_index_94799, 7'h49);
  assign add_95515 = {1'h0, umul_95319[22:3]} + 21'h00_07e9;
  assign sel_95520 = $signed({1'h0, smod_95265[15:0]}) < $signed({1'h0, sel_95326}) ? smod_95265[15:0] : sel_95326;
  assign umul_95521 = umul23b_16b_x_7b(array_index_94987, 7'h47);
  assign add_95523 = {1'h0, umul_95327[22:1]} + 23'h00_1f8b;
  assign sel_95528 = $signed({1'h0, smod_95270[15:0]}) < $signed({1'h0, sel_95334}) ? smod_95270[15:0] : sel_95334;
  assign umul_95529 = umul23b_16b_x_7b(array_index_94993, 7'h47);
  assign add_95531 = {1'h0, umul_95335[22:1]} + 23'h00_1f8b;
  assign sel_95536 = $signed({1'h0, smod_95275[15:0]}) < $signed({1'h0, sel_95342}) ? smod_95275[15:0] : sel_95342;
  assign umul_95537 = umul22b_16b_x_6b(array_index_95181, 6'h3d);
  assign add_95539 = {1'h0, umul_95343[21:2]} + 21'h00_0fb9;
  assign sel_95544 = $signed({1'h0, smod_95280[15:0]}) < $signed({1'h0, sel_95350}) ? smod_95280[15:0] : sel_95350;
  assign umul_95545 = umul22b_16b_x_6b(array_index_95187, 6'h3d);
  assign add_95547 = {1'h0, umul_95351[21:2]} + 21'h00_0fb9;
  assign sel_95552 = $signed({1'h0, smod_95285[15:0]}) < $signed({1'h0, sel_95358}) ? smod_95285[15:0] : sel_95358;
  assign umul_95553 = umul22b_16b_x_6b(array_index_95375, 6'h3b);
  assign add_95555 = {1'h0, umul_95359[21:1]} + 22'h00_1f59;
  assign sel_95560 = $signed({1'h0, smod_95290[15:0]}) < $signed({1'h0, sel_95366}) ? smod_95290[15:0] : sel_95366;
  assign umul_95561 = umul22b_16b_x_6b(array_index_95381, 6'h3b);
  assign add_95563 = {1'h0, umul_95367[21:1]} + 22'h00_1f59;
  assign sel_95568 = $signed({1'h0, smod_95295[15:0]}) < $signed({1'h0, sel_95374}) ? smod_95295[15:0] : sel_95374;
  assign array_index_95569 = set1_unflattened[6'h31];
  assign smod_95573 = $unsigned($signed({9'h000, add_95437, umul_95241[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_95575 = set2_unflattened[6'h31];
  assign smod_95579 = $unsigned($signed({9'h000, add_95445, umul_95249[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_95629 = umul22b_16b_x_6b(array_index_95569, 6'h35);
  assign add_95631 = {1'h0, umul_95435[21:7]} + 16'h007d;
  assign sel_95636 = $signed({1'h0, smod_95379[15:0]}) < $signed({1'h0, sel_95442}) ? smod_95379[15:0] : sel_95442;
  assign umul_95637 = umul22b_16b_x_6b(array_index_95575, 6'h35);
  assign add_95639 = {1'h0, umul_95443[21:7]} + 16'h007d;
  assign sel_95644 = $signed({1'h0, smod_95385[15:0]}) < $signed({1'h0, sel_95450}) ? smod_95385[15:0] : sel_95450;
  assign smod_95648 = $unsigned($signed({8'h00, add_95507, umul_95311[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_95653 = $unsigned($signed({8'h00, add_95515, umul_95319[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_95658 = $unsigned($signed({8'h00, add_95523, umul_95327[0]}) % $signed(32'h0000_3ffd));
  assign smod_95663 = $unsigned($signed({8'h00, add_95531, umul_95335[0]}) % $signed(32'h0000_3ffd));
  assign smod_95668 = $unsigned($signed({9'h000, add_95539, umul_95343[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_95673 = $unsigned($signed({9'h000, add_95547, umul_95351[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_95678 = $unsigned($signed({9'h000, add_95555, umul_95359[0]}) % $signed(32'h0000_3ffd));
  assign smod_95683 = $unsigned($signed({9'h000, add_95563, umul_95367[0]}) % $signed(32'h0000_3ffd));
  assign umul_95697 = umul23b_16b_x_7b(array_index_94987, 7'h49);
  assign add_95699 = {1'h0, umul_95505[22:3]} + 21'h00_07e9;
  assign sel_95704 = $signed({1'h0, smod_95454[15:0]}) < $signed({1'h0, sel_95512}) ? smod_95454[15:0] : sel_95512;
  assign umul_95705 = umul23b_16b_x_7b(array_index_94993, 7'h49);
  assign add_95707 = {1'h0, umul_95513[22:3]} + 21'h00_07e9;
  assign sel_95712 = $signed({1'h0, smod_95459[15:0]}) < $signed({1'h0, sel_95520}) ? smod_95459[15:0] : sel_95520;
  assign umul_95713 = umul23b_16b_x_7b(array_index_95181, 7'h47);
  assign add_95715 = {1'h0, umul_95521[22:1]} + 23'h00_1f8b;
  assign sel_95720 = $signed({1'h0, smod_95464[15:0]}) < $signed({1'h0, sel_95528}) ? smod_95464[15:0] : sel_95528;
  assign umul_95721 = umul23b_16b_x_7b(array_index_95187, 7'h47);
  assign add_95723 = {1'h0, umul_95529[22:1]} + 23'h00_1f8b;
  assign sel_95728 = $signed({1'h0, smod_95469[15:0]}) < $signed({1'h0, sel_95536}) ? smod_95469[15:0] : sel_95536;
  assign umul_95729 = umul22b_16b_x_6b(array_index_95375, 6'h3d);
  assign add_95731 = {1'h0, umul_95537[21:2]} + 21'h00_0fb9;
  assign sel_95736 = $signed({1'h0, smod_95474[15:0]}) < $signed({1'h0, sel_95544}) ? smod_95474[15:0] : sel_95544;
  assign umul_95737 = umul22b_16b_x_6b(array_index_95381, 6'h3d);
  assign add_95739 = {1'h0, umul_95545[21:2]} + 21'h00_0fb9;
  assign sel_95744 = $signed({1'h0, smod_95479[15:0]}) < $signed({1'h0, sel_95552}) ? smod_95479[15:0] : sel_95552;
  assign umul_95745 = umul22b_16b_x_6b(array_index_95569, 6'h3b);
  assign add_95747 = {1'h0, umul_95553[21:1]} + 22'h00_1f59;
  assign sel_95752 = $signed({1'h0, smod_95484[15:0]}) < $signed({1'h0, sel_95560}) ? smod_95484[15:0] : sel_95560;
  assign umul_95753 = umul22b_16b_x_6b(array_index_95575, 6'h3b);
  assign add_95755 = {1'h0, umul_95561[21:1]} + 22'h00_1f59;
  assign sel_95760 = $signed({1'h0, smod_95489[15:0]}) < $signed({1'h0, sel_95568}) ? smod_95489[15:0] : sel_95568;
  assign smod_95763 = $unsigned($signed({9'h000, add_95631, umul_95435[6:0]}) % $signed(32'h0000_3ffd));
  assign smod_95767 = $unsigned($signed({9'h000, add_95639, umul_95443[6:0]}) % $signed(32'h0000_3ffd));
  assign add_95818 = {1'h0, umul_95629[21:7]} + 16'h007d;
  assign sel_95823 = $signed({1'h0, smod_95573[15:0]}) < $signed({1'h0, sel_95636}) ? smod_95573[15:0] : sel_95636;
  assign add_95825 = {1'h0, umul_95637[21:7]} + 16'h007d;
  assign sel_95830 = $signed({1'h0, smod_95579[15:0]}) < $signed({1'h0, sel_95644}) ? smod_95579[15:0] : sel_95644;
  assign smod_95834 = $unsigned($signed({8'h00, add_95699, umul_95505[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_95839 = $unsigned($signed({8'h00, add_95707, umul_95513[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_95844 = $unsigned($signed({8'h00, add_95715, umul_95521[0]}) % $signed(32'h0000_3ffd));
  assign smod_95849 = $unsigned($signed({8'h00, add_95723, umul_95529[0]}) % $signed(32'h0000_3ffd));
  assign smod_95854 = $unsigned($signed({9'h000, add_95731, umul_95537[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_95859 = $unsigned($signed({9'h000, add_95739, umul_95545[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_95863 = $unsigned($signed({9'h000, add_95747, umul_95553[0]}) % $signed(32'h0000_3ffd));
  assign smod_95867 = $unsigned($signed({9'h000, add_95755, umul_95561[0]}) % $signed(32'h0000_3ffd));
  assign umul_95877 = umul23b_16b_x_7b(array_index_95181, 7'h49);
  assign add_95879 = {1'h0, umul_95697[22:3]} + 21'h00_07e9;
  assign sel_95884 = $signed({1'h0, smod_95648[15:0]}) < $signed({1'h0, sel_95704}) ? smod_95648[15:0] : sel_95704;
  assign umul_95885 = umul23b_16b_x_7b(array_index_95187, 7'h49);
  assign add_95887 = {1'h0, umul_95705[22:3]} + 21'h00_07e9;
  assign sel_95892 = $signed({1'h0, smod_95653[15:0]}) < $signed({1'h0, sel_95712}) ? smod_95653[15:0] : sel_95712;
  assign umul_95893 = umul23b_16b_x_7b(array_index_95375, 7'h47);
  assign add_95895 = {1'h0, umul_95713[22:1]} + 23'h00_1f8b;
  assign sel_95900 = $signed({1'h0, smod_95658[15:0]}) < $signed({1'h0, sel_95720}) ? smod_95658[15:0] : sel_95720;
  assign umul_95901 = umul23b_16b_x_7b(array_index_95381, 7'h47);
  assign add_95903 = {1'h0, umul_95721[22:1]} + 23'h00_1f8b;
  assign sel_95908 = $signed({1'h0, smod_95663[15:0]}) < $signed({1'h0, sel_95728}) ? smod_95663[15:0] : sel_95728;
  assign umul_95909 = umul22b_16b_x_6b(array_index_95569, 6'h3d);
  assign add_95911 = {1'h0, umul_95729[21:2]} + 21'h00_0fb9;
  assign sel_95916 = $signed({1'h0, smod_95668[15:0]}) < $signed({1'h0, sel_95736}) ? smod_95668[15:0] : sel_95736;
  assign umul_95917 = umul22b_16b_x_6b(array_index_95575, 6'h3d);
  assign add_95919 = {1'h0, umul_95737[21:2]} + 21'h00_0fb9;
  assign sel_95924 = $signed({1'h0, smod_95673[15:0]}) < $signed({1'h0, sel_95744}) ? smod_95673[15:0] : sel_95744;
  assign add_95926 = {1'h0, umul_95745[21:1]} + 22'h00_1f59;
  assign sel_95931 = $signed({1'h0, smod_95678[15:0]}) < $signed({1'h0, sel_95752}) ? smod_95678[15:0] : sel_95752;
  assign add_95933 = {1'h0, umul_95753[21:1]} + 22'h00_1f59;
  assign sel_95938 = $signed({1'h0, smod_95683[15:0]}) < $signed({1'h0, sel_95760}) ? smod_95683[15:0] : sel_95760;
  assign smod_95939 = $unsigned($signed({9'h000, add_95818, umul_95629[6:0]}) % $signed(32'h0000_3ffd));
  assign smod_95941 = $unsigned($signed({9'h000, add_95825, umul_95637[6:0]}) % $signed(32'h0000_3ffd));
  assign sel_95990 = $signed({1'h0, smod_95763[15:0]}) < $signed({1'h0, sel_95823}) ? smod_95763[15:0] : sel_95823;
  assign sel_95994 = $signed({1'h0, smod_95767[15:0]}) < $signed({1'h0, sel_95830}) ? smod_95767[15:0] : sel_95830;
  assign smod_95998 = $unsigned($signed({8'h00, add_95879, umul_95697[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_96003 = $unsigned($signed({8'h00, add_95887, umul_95705[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_96008 = $unsigned($signed({8'h00, add_95895, umul_95713[0]}) % $signed(32'h0000_3ffd));
  assign smod_96013 = $unsigned($signed({8'h00, add_95903, umul_95721[0]}) % $signed(32'h0000_3ffd));
  assign smod_96017 = $unsigned($signed({9'h000, add_95911, umul_95729[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_96021 = $unsigned($signed({9'h000, add_95919, umul_95737[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_96023 = $unsigned($signed({9'h000, add_95926, umul_95745[0]}) % $signed(32'h0000_3ffd));
  assign smod_96025 = $unsigned($signed({9'h000, add_95933, umul_95753[0]}) % $signed(32'h0000_3ffd));
  assign umul_96031 = umul23b_16b_x_7b(array_index_95375, 7'h49);
  assign add_96033 = {1'h0, umul_95877[22:3]} + 21'h00_07e9;
  assign sel_96038 = $signed({1'h0, smod_95834[15:0]}) < $signed({1'h0, sel_95884}) ? smod_95834[15:0] : sel_95884;
  assign umul_96039 = umul23b_16b_x_7b(array_index_95381, 7'h49);
  assign add_96041 = {1'h0, umul_95885[22:3]} + 21'h00_07e9;
  assign sel_96046 = $signed({1'h0, smod_95839[15:0]}) < $signed({1'h0, sel_95892}) ? smod_95839[15:0] : sel_95892;
  assign umul_96047 = umul23b_16b_x_7b(array_index_95569, 7'h47);
  assign add_96049 = {1'h0, umul_95893[22:1]} + 23'h00_1f8b;
  assign sel_96054 = $signed({1'h0, smod_95844[15:0]}) < $signed({1'h0, sel_95900}) ? smod_95844[15:0] : sel_95900;
  assign umul_96055 = umul23b_16b_x_7b(array_index_95575, 7'h47);
  assign add_96057 = {1'h0, umul_95901[22:1]} + 23'h00_1f8b;
  assign sel_96062 = $signed({1'h0, smod_95849[15:0]}) < $signed({1'h0, sel_95908}) ? smod_95849[15:0] : sel_95908;
  assign add_96064 = {1'h0, umul_95909[21:2]} + 21'h00_0fb9;
  assign sel_96069 = $signed({1'h0, smod_95854[15:0]}) < $signed({1'h0, sel_95916}) ? smod_95854[15:0] : sel_95916;
  assign add_96071 = {1'h0, umul_95917[21:2]} + 21'h00_0fb9;
  assign sel_96076 = $signed({1'h0, smod_95859[15:0]}) < $signed({1'h0, sel_95924}) ? smod_95859[15:0] : sel_95924;
  assign sel_96080 = $signed({1'h0, smod_95863[15:0]}) < $signed({1'h0, sel_95931}) ? smod_95863[15:0] : sel_95931;
  assign sel_96084 = $signed({1'h0, smod_95867[15:0]}) < $signed({1'h0, sel_95938}) ? smod_95867[15:0] : sel_95938;
  assign smod_96128 = $unsigned($signed({8'h00, add_96033, umul_95877[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_96133 = $unsigned($signed({8'h00, add_96041, umul_95885[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_96137 = $unsigned($signed({8'h00, add_96049, umul_95893[0]}) % $signed(32'h0000_3ffd));
  assign smod_96141 = $unsigned($signed({8'h00, add_96057, umul_95901[0]}) % $signed(32'h0000_3ffd));
  assign smod_96143 = $unsigned($signed({9'h000, add_96064, umul_95909[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_96145 = $unsigned($signed({9'h000, add_96071, umul_95917[1:0]}) % $signed(32'h0000_3ffd));
  assign umul_96151 = umul23b_16b_x_7b(array_index_95569, 7'h49);
  assign add_96153 = {1'h0, umul_96031[22:3]} + 21'h00_07e9;
  assign sel_96158 = $signed({1'h0, smod_95998[15:0]}) < $signed({1'h0, sel_96038}) ? smod_95998[15:0] : sel_96038;
  assign umul_96159 = umul23b_16b_x_7b(array_index_95575, 7'h49);
  assign add_96161 = {1'h0, umul_96039[22:3]} + 21'h00_07e9;
  assign sel_96166 = $signed({1'h0, smod_96003[15:0]}) < $signed({1'h0, sel_96046}) ? smod_96003[15:0] : sel_96046;
  assign add_96168 = {1'h0, umul_96047[22:1]} + 23'h00_1f8b;
  assign sel_96173 = $signed({1'h0, smod_96008[15:0]}) < $signed({1'h0, sel_96054}) ? smod_96008[15:0] : sel_96054;
  assign add_96175 = {1'h0, umul_96055[22:1]} + 23'h00_1f8b;
  assign sel_96180 = $signed({1'h0, smod_96013[15:0]}) < $signed({1'h0, sel_96062}) ? smod_96013[15:0] : sel_96062;
  assign sel_96184 = $signed({1'h0, smod_96017[15:0]}) < $signed({1'h0, sel_96069}) ? smod_96017[15:0] : sel_96069;
  assign sel_96188 = $signed({1'h0, smod_96021[15:0]}) < $signed({1'h0, sel_96076}) ? smod_96021[15:0] : sel_96076;
  assign concat_96191 = {1'h0, ($signed({1'h0, smod_95939[15:0]}) < $signed({1'h0, sel_95990}) ? smod_95939[15:0] : sel_95990) == ($signed({1'h0, smod_95941[15:0]}) < $signed({1'h0, sel_95994}) ? smod_95941[15:0] : sel_95994)};
  assign add_96218 = concat_96191 + 2'h1;
  assign smod_96221 = $unsigned($signed({8'h00, add_96153, umul_96031[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_96225 = $unsigned($signed({8'h00, add_96161, umul_96039[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_96227 = $unsigned($signed({8'h00, add_96168, umul_96047[0]}) % $signed(32'h0000_3ffd));
  assign smod_96229 = $unsigned($signed({8'h00, add_96175, umul_96055[0]}) % $signed(32'h0000_3ffd));
  assign add_96236 = {1'h0, umul_96151[22:3]} + 21'h00_07e9;
  assign sel_96241 = $signed({1'h0, smod_96128[15:0]}) < $signed({1'h0, sel_96158}) ? smod_96128[15:0] : sel_96158;
  assign add_96243 = {1'h0, umul_96159[22:3]} + 21'h00_07e9;
  assign sel_96248 = $signed({1'h0, smod_96133[15:0]}) < $signed({1'h0, sel_96166}) ? smod_96133[15:0] : sel_96166;
  assign sel_96252 = $signed({1'h0, smod_96137[15:0]}) < $signed({1'h0, sel_96173}) ? smod_96137[15:0] : sel_96173;
  assign sel_96256 = $signed({1'h0, smod_96141[15:0]}) < $signed({1'h0, sel_96180}) ? smod_96141[15:0] : sel_96180;
  assign concat_96259 = {1'h0, ($signed({1'h0, smod_96023[15:0]}) < $signed({1'h0, sel_96080}) ? smod_96023[15:0] : sel_96080) == ($signed({1'h0, smod_96025[15:0]}) < $signed({1'h0, sel_96084}) ? smod_96025[15:0] : sel_96084) ? add_96218 : concat_96191};
  assign add_96274 = concat_96259 + 3'h1;
  assign smod_96275 = $unsigned($signed({8'h00, add_96236, umul_96151[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_96277 = $unsigned($signed({8'h00, add_96243, umul_96159[2:0]}) % $signed(32'h0000_3ffd));
  assign sel_96286 = $signed({1'h0, smod_96221[15:0]}) < $signed({1'h0, sel_96241}) ? smod_96221[15:0] : sel_96241;
  assign sel_96290 = $signed({1'h0, smod_96225[15:0]}) < $signed({1'h0, sel_96248}) ? smod_96225[15:0] : sel_96248;
  assign concat_96293 = {1'h0, ($signed({1'h0, smod_96143[15:0]}) < $signed({1'h0, sel_96184}) ? smod_96143[15:0] : sel_96184) == ($signed({1'h0, smod_96145[15:0]}) < $signed({1'h0, sel_96188}) ? smod_96145[15:0] : sel_96188) ? add_96274 : concat_96259};
  assign add_96300 = concat_96293 + 4'h1;
  assign concat_96307 = {1'h0, ($signed({1'h0, smod_96227[15:0]}) < $signed({1'h0, sel_96252}) ? smod_96227[15:0] : sel_96252) == ($signed({1'h0, smod_96229[15:0]}) < $signed({1'h0, sel_96256}) ? smod_96229[15:0] : sel_96256) ? add_96300 : concat_96293};
  assign add_96310 = concat_96307 + 5'h01;
  assign out = {{11'h000, ($signed({1'h0, smod_96275[15:0]}) < $signed({1'h0, sel_96286}) ? smod_96275[15:0] : sel_96286) == ($signed({1'h0, smod_96277[15:0]}) < $signed({1'h0, sel_96290}) ? smod_96277[15:0] : sel_96290) ? add_96310 : concat_96307}, {set1_unflattened[49], set1_unflattened[48], set1_unflattened[47], set1_unflattened[46], set1_unflattened[45], set1_unflattened[44], set1_unflattened[43], set1_unflattened[42], set1_unflattened[41], set1_unflattened[40], set1_unflattened[39], set1_unflattened[38], set1_unflattened[37], set1_unflattened[36], set1_unflattened[35], set1_unflattened[34], set1_unflattened[33], set1_unflattened[32], set1_unflattened[31], set1_unflattened[30], set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[49], set2_unflattened[48], set2_unflattened[47], set2_unflattened[46], set2_unflattened[45], set2_unflattened[44], set2_unflattened[43], set2_unflattened[42], set2_unflattened[41], set2_unflattened[40], set2_unflattened[39], set2_unflattened[38], set2_unflattened[37], set2_unflattened[36], set2_unflattened[35], set2_unflattened[34], set2_unflattened[33], set2_unflattened[32], set2_unflattened[31], set2_unflattened[30], set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
