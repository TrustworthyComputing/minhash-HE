module min_hash(
  input wire [159:0] set1,
  input wire [159:0] set2,
  output wire [327:0] out
);
  wire [15:0] set1_unflattened[10];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  wire [15:0] set2_unflattened[10];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  wire [15:0] array_index_9993;
  wire [15:0] array_index_9994;
  wire [15:0] array_index_9998;
  wire [1:0] concat_9999;
  wire [1:0] add_10002;
  wire [15:0] array_index_10006;
  wire [2:0] concat_10007;
  wire [2:0] add_10010;
  wire [15:0] array_index_10014;
  wire [3:0] concat_10015;
  wire [3:0] add_10018;
  wire [15:0] array_index_10022;
  wire [4:0] concat_10023;
  wire [4:0] add_10026;
  wire [15:0] array_index_10030;
  wire [5:0] concat_10031;
  wire [5:0] add_10034;
  wire [15:0] array_index_10038;
  wire [6:0] concat_10039;
  wire [6:0] add_10042;
  wire [15:0] array_index_10046;
  wire [7:0] concat_10047;
  wire [7:0] add_10051;
  wire [15:0] array_index_10052;
  wire [7:0] sel_10053;
  wire [7:0] add_10057;
  wire [15:0] array_index_10058;
  wire [7:0] sel_10059;
  wire [7:0] add_10063;
  wire [15:0] array_index_10064;
  wire [7:0] sel_10065;
  wire [7:0] add_10068;
  wire [7:0] sel_10069;
  wire [7:0] add_10072;
  wire [7:0] sel_10073;
  wire [7:0] add_10076;
  wire [7:0] sel_10077;
  wire [7:0] add_10080;
  wire [7:0] sel_10081;
  wire [7:0] add_10084;
  wire [7:0] sel_10085;
  wire [7:0] add_10088;
  wire [7:0] sel_10089;
  wire [7:0] add_10092;
  wire [7:0] sel_10093;
  wire [7:0] add_10096;
  wire [7:0] sel_10097;
  wire [7:0] add_10100;
  wire [7:0] sel_10101;
  wire [7:0] add_10105;
  wire [15:0] array_index_10106;
  wire [7:0] sel_10107;
  wire [7:0] add_10110;
  wire [7:0] sel_10111;
  wire [7:0] add_10114;
  wire [7:0] sel_10115;
  wire [7:0] add_10118;
  wire [7:0] sel_10119;
  wire [7:0] add_10122;
  wire [7:0] sel_10123;
  wire [7:0] add_10126;
  wire [7:0] sel_10127;
  wire [7:0] add_10130;
  wire [7:0] sel_10131;
  wire [7:0] add_10134;
  wire [7:0] sel_10135;
  wire [7:0] add_10138;
  wire [7:0] sel_10139;
  wire [7:0] add_10142;
  wire [7:0] sel_10143;
  wire [7:0] add_10147;
  wire [15:0] array_index_10148;
  wire [7:0] sel_10149;
  wire [7:0] add_10152;
  wire [7:0] sel_10153;
  wire [7:0] add_10156;
  wire [7:0] sel_10157;
  wire [7:0] add_10160;
  wire [7:0] sel_10161;
  wire [7:0] add_10164;
  wire [7:0] sel_10165;
  wire [7:0] add_10168;
  wire [7:0] sel_10169;
  wire [7:0] add_10172;
  wire [7:0] sel_10173;
  wire [7:0] add_10176;
  wire [7:0] sel_10177;
  wire [7:0] add_10180;
  wire [7:0] sel_10181;
  wire [7:0] add_10184;
  wire [7:0] sel_10185;
  wire [7:0] add_10189;
  wire [15:0] array_index_10190;
  wire [7:0] sel_10191;
  wire [7:0] add_10194;
  wire [7:0] sel_10195;
  wire [7:0] add_10198;
  wire [7:0] sel_10199;
  wire [7:0] add_10202;
  wire [7:0] sel_10203;
  wire [7:0] add_10206;
  wire [7:0] sel_10207;
  wire [7:0] add_10210;
  wire [7:0] sel_10211;
  wire [7:0] add_10214;
  wire [7:0] sel_10215;
  wire [7:0] add_10218;
  wire [7:0] sel_10219;
  wire [7:0] add_10222;
  wire [7:0] sel_10223;
  wire [7:0] add_10226;
  wire [7:0] sel_10227;
  wire [7:0] add_10231;
  wire [15:0] array_index_10232;
  wire [7:0] sel_10233;
  wire [7:0] add_10236;
  wire [7:0] sel_10237;
  wire [7:0] add_10240;
  wire [7:0] sel_10241;
  wire [7:0] add_10244;
  wire [7:0] sel_10245;
  wire [7:0] add_10248;
  wire [7:0] sel_10249;
  wire [7:0] add_10252;
  wire [7:0] sel_10253;
  wire [7:0] add_10256;
  wire [7:0] sel_10257;
  wire [7:0] add_10260;
  wire [7:0] sel_10261;
  wire [7:0] add_10264;
  wire [7:0] sel_10265;
  wire [7:0] add_10268;
  wire [7:0] sel_10269;
  wire [7:0] add_10273;
  wire [15:0] array_index_10274;
  wire [7:0] sel_10275;
  wire [7:0] add_10278;
  wire [7:0] sel_10279;
  wire [7:0] add_10282;
  wire [7:0] sel_10283;
  wire [7:0] add_10286;
  wire [7:0] sel_10287;
  wire [7:0] add_10290;
  wire [7:0] sel_10291;
  wire [7:0] add_10294;
  wire [7:0] sel_10295;
  wire [7:0] add_10298;
  wire [7:0] sel_10299;
  wire [7:0] add_10302;
  wire [7:0] sel_10303;
  wire [7:0] add_10306;
  wire [7:0] sel_10307;
  wire [7:0] add_10310;
  wire [7:0] sel_10311;
  wire [7:0] add_10315;
  wire [15:0] array_index_10316;
  wire [7:0] sel_10317;
  wire [7:0] add_10320;
  wire [7:0] sel_10321;
  wire [7:0] add_10324;
  wire [7:0] sel_10325;
  wire [7:0] add_10328;
  wire [7:0] sel_10329;
  wire [7:0] add_10332;
  wire [7:0] sel_10333;
  wire [7:0] add_10336;
  wire [7:0] sel_10337;
  wire [7:0] add_10340;
  wire [7:0] sel_10341;
  wire [7:0] add_10344;
  wire [7:0] sel_10345;
  wire [7:0] add_10348;
  wire [7:0] sel_10349;
  wire [7:0] add_10352;
  wire [7:0] sel_10353;
  wire [7:0] add_10357;
  wire [15:0] array_index_10358;
  wire [7:0] sel_10359;
  wire [7:0] add_10362;
  wire [7:0] sel_10363;
  wire [7:0] add_10366;
  wire [7:0] sel_10367;
  wire [7:0] add_10370;
  wire [7:0] sel_10371;
  wire [7:0] add_10374;
  wire [7:0] sel_10375;
  wire [7:0] add_10378;
  wire [7:0] sel_10379;
  wire [7:0] add_10382;
  wire [7:0] sel_10383;
  wire [7:0] add_10386;
  wire [7:0] sel_10387;
  wire [7:0] add_10390;
  wire [7:0] sel_10391;
  wire [7:0] add_10394;
  wire [7:0] sel_10395;
  wire [7:0] add_10399;
  wire [15:0] array_index_10400;
  wire [7:0] sel_10401;
  wire [7:0] add_10404;
  wire [7:0] sel_10405;
  wire [7:0] add_10408;
  wire [7:0] sel_10409;
  wire [7:0] add_10412;
  wire [7:0] sel_10413;
  wire [7:0] add_10416;
  wire [7:0] sel_10417;
  wire [7:0] add_10420;
  wire [7:0] sel_10421;
  wire [7:0] add_10424;
  wire [7:0] sel_10425;
  wire [7:0] add_10428;
  wire [7:0] sel_10429;
  wire [7:0] add_10432;
  wire [7:0] sel_10433;
  wire [7:0] add_10436;
  wire [7:0] sel_10437;
  wire [7:0] add_10440;
  assign array_index_9993 = set1_unflattened[4'h0];
  assign array_index_9994 = set2_unflattened[4'h0];
  assign array_index_9998 = set2_unflattened[4'h1];
  assign concat_9999 = {1'h0, array_index_9993 == array_index_9994};
  assign add_10002 = concat_9999 + 2'h1;
  assign array_index_10006 = set2_unflattened[4'h2];
  assign concat_10007 = {1'h0, array_index_9993 == array_index_9998 ? add_10002 : concat_9999};
  assign add_10010 = concat_10007 + 3'h1;
  assign array_index_10014 = set2_unflattened[4'h3];
  assign concat_10015 = {1'h0, array_index_9993 == array_index_10006 ? add_10010 : concat_10007};
  assign add_10018 = concat_10015 + 4'h1;
  assign array_index_10022 = set2_unflattened[4'h4];
  assign concat_10023 = {1'h0, array_index_9993 == array_index_10014 ? add_10018 : concat_10015};
  assign add_10026 = concat_10023 + 5'h01;
  assign array_index_10030 = set2_unflattened[4'h5];
  assign concat_10031 = {1'h0, array_index_9993 == array_index_10022 ? add_10026 : concat_10023};
  assign add_10034 = concat_10031 + 6'h01;
  assign array_index_10038 = set2_unflattened[4'h6];
  assign concat_10039 = {1'h0, array_index_9993 == array_index_10030 ? add_10034 : concat_10031};
  assign add_10042 = concat_10039 + 7'h01;
  assign array_index_10046 = set2_unflattened[4'h7];
  assign concat_10047 = {1'h0, array_index_9993 == array_index_10038 ? add_10042 : concat_10039};
  assign add_10051 = concat_10047 + 8'h01;
  assign array_index_10052 = set2_unflattened[4'h8];
  assign sel_10053 = array_index_9993 == array_index_10046 ? add_10051 : concat_10047;
  assign add_10057 = sel_10053 + 8'h01;
  assign array_index_10058 = set2_unflattened[4'h9];
  assign sel_10059 = array_index_9993 == array_index_10052 ? add_10057 : sel_10053;
  assign add_10063 = sel_10059 + 8'h01;
  assign array_index_10064 = set1_unflattened[4'h1];
  assign sel_10065 = array_index_9993 == array_index_10058 ? add_10063 : sel_10059;
  assign add_10068 = sel_10065 + 8'h01;
  assign sel_10069 = array_index_10064 == array_index_9994 ? add_10068 : sel_10065;
  assign add_10072 = sel_10069 + 8'h01;
  assign sel_10073 = array_index_10064 == array_index_9998 ? add_10072 : sel_10069;
  assign add_10076 = sel_10073 + 8'h01;
  assign sel_10077 = array_index_10064 == array_index_10006 ? add_10076 : sel_10073;
  assign add_10080 = sel_10077 + 8'h01;
  assign sel_10081 = array_index_10064 == array_index_10014 ? add_10080 : sel_10077;
  assign add_10084 = sel_10081 + 8'h01;
  assign sel_10085 = array_index_10064 == array_index_10022 ? add_10084 : sel_10081;
  assign add_10088 = sel_10085 + 8'h01;
  assign sel_10089 = array_index_10064 == array_index_10030 ? add_10088 : sel_10085;
  assign add_10092 = sel_10089 + 8'h01;
  assign sel_10093 = array_index_10064 == array_index_10038 ? add_10092 : sel_10089;
  assign add_10096 = sel_10093 + 8'h01;
  assign sel_10097 = array_index_10064 == array_index_10046 ? add_10096 : sel_10093;
  assign add_10100 = sel_10097 + 8'h01;
  assign sel_10101 = array_index_10064 == array_index_10052 ? add_10100 : sel_10097;
  assign add_10105 = sel_10101 + 8'h01;
  assign array_index_10106 = set1_unflattened[4'h2];
  assign sel_10107 = array_index_10064 == array_index_10058 ? add_10105 : sel_10101;
  assign add_10110 = sel_10107 + 8'h01;
  assign sel_10111 = array_index_10106 == array_index_9994 ? add_10110 : sel_10107;
  assign add_10114 = sel_10111 + 8'h01;
  assign sel_10115 = array_index_10106 == array_index_9998 ? add_10114 : sel_10111;
  assign add_10118 = sel_10115 + 8'h01;
  assign sel_10119 = array_index_10106 == array_index_10006 ? add_10118 : sel_10115;
  assign add_10122 = sel_10119 + 8'h01;
  assign sel_10123 = array_index_10106 == array_index_10014 ? add_10122 : sel_10119;
  assign add_10126 = sel_10123 + 8'h01;
  assign sel_10127 = array_index_10106 == array_index_10022 ? add_10126 : sel_10123;
  assign add_10130 = sel_10127 + 8'h01;
  assign sel_10131 = array_index_10106 == array_index_10030 ? add_10130 : sel_10127;
  assign add_10134 = sel_10131 + 8'h01;
  assign sel_10135 = array_index_10106 == array_index_10038 ? add_10134 : sel_10131;
  assign add_10138 = sel_10135 + 8'h01;
  assign sel_10139 = array_index_10106 == array_index_10046 ? add_10138 : sel_10135;
  assign add_10142 = sel_10139 + 8'h01;
  assign sel_10143 = array_index_10106 == array_index_10052 ? add_10142 : sel_10139;
  assign add_10147 = sel_10143 + 8'h01;
  assign array_index_10148 = set1_unflattened[4'h3];
  assign sel_10149 = array_index_10106 == array_index_10058 ? add_10147 : sel_10143;
  assign add_10152 = sel_10149 + 8'h01;
  assign sel_10153 = array_index_10148 == array_index_9994 ? add_10152 : sel_10149;
  assign add_10156 = sel_10153 + 8'h01;
  assign sel_10157 = array_index_10148 == array_index_9998 ? add_10156 : sel_10153;
  assign add_10160 = sel_10157 + 8'h01;
  assign sel_10161 = array_index_10148 == array_index_10006 ? add_10160 : sel_10157;
  assign add_10164 = sel_10161 + 8'h01;
  assign sel_10165 = array_index_10148 == array_index_10014 ? add_10164 : sel_10161;
  assign add_10168 = sel_10165 + 8'h01;
  assign sel_10169 = array_index_10148 == array_index_10022 ? add_10168 : sel_10165;
  assign add_10172 = sel_10169 + 8'h01;
  assign sel_10173 = array_index_10148 == array_index_10030 ? add_10172 : sel_10169;
  assign add_10176 = sel_10173 + 8'h01;
  assign sel_10177 = array_index_10148 == array_index_10038 ? add_10176 : sel_10173;
  assign add_10180 = sel_10177 + 8'h01;
  assign sel_10181 = array_index_10148 == array_index_10046 ? add_10180 : sel_10177;
  assign add_10184 = sel_10181 + 8'h01;
  assign sel_10185 = array_index_10148 == array_index_10052 ? add_10184 : sel_10181;
  assign add_10189 = sel_10185 + 8'h01;
  assign array_index_10190 = set1_unflattened[4'h4];
  assign sel_10191 = array_index_10148 == array_index_10058 ? add_10189 : sel_10185;
  assign add_10194 = sel_10191 + 8'h01;
  assign sel_10195 = array_index_10190 == array_index_9994 ? add_10194 : sel_10191;
  assign add_10198 = sel_10195 + 8'h01;
  assign sel_10199 = array_index_10190 == array_index_9998 ? add_10198 : sel_10195;
  assign add_10202 = sel_10199 + 8'h01;
  assign sel_10203 = array_index_10190 == array_index_10006 ? add_10202 : sel_10199;
  assign add_10206 = sel_10203 + 8'h01;
  assign sel_10207 = array_index_10190 == array_index_10014 ? add_10206 : sel_10203;
  assign add_10210 = sel_10207 + 8'h01;
  assign sel_10211 = array_index_10190 == array_index_10022 ? add_10210 : sel_10207;
  assign add_10214 = sel_10211 + 8'h01;
  assign sel_10215 = array_index_10190 == array_index_10030 ? add_10214 : sel_10211;
  assign add_10218 = sel_10215 + 8'h01;
  assign sel_10219 = array_index_10190 == array_index_10038 ? add_10218 : sel_10215;
  assign add_10222 = sel_10219 + 8'h01;
  assign sel_10223 = array_index_10190 == array_index_10046 ? add_10222 : sel_10219;
  assign add_10226 = sel_10223 + 8'h01;
  assign sel_10227 = array_index_10190 == array_index_10052 ? add_10226 : sel_10223;
  assign add_10231 = sel_10227 + 8'h01;
  assign array_index_10232 = set1_unflattened[4'h5];
  assign sel_10233 = array_index_10190 == array_index_10058 ? add_10231 : sel_10227;
  assign add_10236 = sel_10233 + 8'h01;
  assign sel_10237 = array_index_10232 == array_index_9994 ? add_10236 : sel_10233;
  assign add_10240 = sel_10237 + 8'h01;
  assign sel_10241 = array_index_10232 == array_index_9998 ? add_10240 : sel_10237;
  assign add_10244 = sel_10241 + 8'h01;
  assign sel_10245 = array_index_10232 == array_index_10006 ? add_10244 : sel_10241;
  assign add_10248 = sel_10245 + 8'h01;
  assign sel_10249 = array_index_10232 == array_index_10014 ? add_10248 : sel_10245;
  assign add_10252 = sel_10249 + 8'h01;
  assign sel_10253 = array_index_10232 == array_index_10022 ? add_10252 : sel_10249;
  assign add_10256 = sel_10253 + 8'h01;
  assign sel_10257 = array_index_10232 == array_index_10030 ? add_10256 : sel_10253;
  assign add_10260 = sel_10257 + 8'h01;
  assign sel_10261 = array_index_10232 == array_index_10038 ? add_10260 : sel_10257;
  assign add_10264 = sel_10261 + 8'h01;
  assign sel_10265 = array_index_10232 == array_index_10046 ? add_10264 : sel_10261;
  assign add_10268 = sel_10265 + 8'h01;
  assign sel_10269 = array_index_10232 == array_index_10052 ? add_10268 : sel_10265;
  assign add_10273 = sel_10269 + 8'h01;
  assign array_index_10274 = set1_unflattened[4'h6];
  assign sel_10275 = array_index_10232 == array_index_10058 ? add_10273 : sel_10269;
  assign add_10278 = sel_10275 + 8'h01;
  assign sel_10279 = array_index_10274 == array_index_9994 ? add_10278 : sel_10275;
  assign add_10282 = sel_10279 + 8'h01;
  assign sel_10283 = array_index_10274 == array_index_9998 ? add_10282 : sel_10279;
  assign add_10286 = sel_10283 + 8'h01;
  assign sel_10287 = array_index_10274 == array_index_10006 ? add_10286 : sel_10283;
  assign add_10290 = sel_10287 + 8'h01;
  assign sel_10291 = array_index_10274 == array_index_10014 ? add_10290 : sel_10287;
  assign add_10294 = sel_10291 + 8'h01;
  assign sel_10295 = array_index_10274 == array_index_10022 ? add_10294 : sel_10291;
  assign add_10298 = sel_10295 + 8'h01;
  assign sel_10299 = array_index_10274 == array_index_10030 ? add_10298 : sel_10295;
  assign add_10302 = sel_10299 + 8'h01;
  assign sel_10303 = array_index_10274 == array_index_10038 ? add_10302 : sel_10299;
  assign add_10306 = sel_10303 + 8'h01;
  assign sel_10307 = array_index_10274 == array_index_10046 ? add_10306 : sel_10303;
  assign add_10310 = sel_10307 + 8'h01;
  assign sel_10311 = array_index_10274 == array_index_10052 ? add_10310 : sel_10307;
  assign add_10315 = sel_10311 + 8'h01;
  assign array_index_10316 = set1_unflattened[4'h7];
  assign sel_10317 = array_index_10274 == array_index_10058 ? add_10315 : sel_10311;
  assign add_10320 = sel_10317 + 8'h01;
  assign sel_10321 = array_index_10316 == array_index_9994 ? add_10320 : sel_10317;
  assign add_10324 = sel_10321 + 8'h01;
  assign sel_10325 = array_index_10316 == array_index_9998 ? add_10324 : sel_10321;
  assign add_10328 = sel_10325 + 8'h01;
  assign sel_10329 = array_index_10316 == array_index_10006 ? add_10328 : sel_10325;
  assign add_10332 = sel_10329 + 8'h01;
  assign sel_10333 = array_index_10316 == array_index_10014 ? add_10332 : sel_10329;
  assign add_10336 = sel_10333 + 8'h01;
  assign sel_10337 = array_index_10316 == array_index_10022 ? add_10336 : sel_10333;
  assign add_10340 = sel_10337 + 8'h01;
  assign sel_10341 = array_index_10316 == array_index_10030 ? add_10340 : sel_10337;
  assign add_10344 = sel_10341 + 8'h01;
  assign sel_10345 = array_index_10316 == array_index_10038 ? add_10344 : sel_10341;
  assign add_10348 = sel_10345 + 8'h01;
  assign sel_10349 = array_index_10316 == array_index_10046 ? add_10348 : sel_10345;
  assign add_10352 = sel_10349 + 8'h01;
  assign sel_10353 = array_index_10316 == array_index_10052 ? add_10352 : sel_10349;
  assign add_10357 = sel_10353 + 8'h01;
  assign array_index_10358 = set1_unflattened[4'h8];
  assign sel_10359 = array_index_10316 == array_index_10058 ? add_10357 : sel_10353;
  assign add_10362 = sel_10359 + 8'h01;
  assign sel_10363 = array_index_10358 == array_index_9994 ? add_10362 : sel_10359;
  assign add_10366 = sel_10363 + 8'h01;
  assign sel_10367 = array_index_10358 == array_index_9998 ? add_10366 : sel_10363;
  assign add_10370 = sel_10367 + 8'h01;
  assign sel_10371 = array_index_10358 == array_index_10006 ? add_10370 : sel_10367;
  assign add_10374 = sel_10371 + 8'h01;
  assign sel_10375 = array_index_10358 == array_index_10014 ? add_10374 : sel_10371;
  assign add_10378 = sel_10375 + 8'h01;
  assign sel_10379 = array_index_10358 == array_index_10022 ? add_10378 : sel_10375;
  assign add_10382 = sel_10379 + 8'h01;
  assign sel_10383 = array_index_10358 == array_index_10030 ? add_10382 : sel_10379;
  assign add_10386 = sel_10383 + 8'h01;
  assign sel_10387 = array_index_10358 == array_index_10038 ? add_10386 : sel_10383;
  assign add_10390 = sel_10387 + 8'h01;
  assign sel_10391 = array_index_10358 == array_index_10046 ? add_10390 : sel_10387;
  assign add_10394 = sel_10391 + 8'h01;
  assign sel_10395 = array_index_10358 == array_index_10052 ? add_10394 : sel_10391;
  assign add_10399 = sel_10395 + 8'h01;
  assign array_index_10400 = set1_unflattened[4'h9];
  assign sel_10401 = array_index_10358 == array_index_10058 ? add_10399 : sel_10395;
  assign add_10404 = sel_10401 + 8'h01;
  assign sel_10405 = array_index_10400 == array_index_9994 ? add_10404 : sel_10401;
  assign add_10408 = sel_10405 + 8'h01;
  assign sel_10409 = array_index_10400 == array_index_9998 ? add_10408 : sel_10405;
  assign add_10412 = sel_10409 + 8'h01;
  assign sel_10413 = array_index_10400 == array_index_10006 ? add_10412 : sel_10409;
  assign add_10416 = sel_10413 + 8'h01;
  assign sel_10417 = array_index_10400 == array_index_10014 ? add_10416 : sel_10413;
  assign add_10420 = sel_10417 + 8'h01;
  assign sel_10421 = array_index_10400 == array_index_10022 ? add_10420 : sel_10417;
  assign add_10424 = sel_10421 + 8'h01;
  assign sel_10425 = array_index_10400 == array_index_10030 ? add_10424 : sel_10421;
  assign add_10428 = sel_10425 + 8'h01;
  assign sel_10429 = array_index_10400 == array_index_10038 ? add_10428 : sel_10425;
  assign add_10432 = sel_10429 + 8'h01;
  assign sel_10433 = array_index_10400 == array_index_10046 ? add_10432 : sel_10429;
  assign add_10436 = sel_10433 + 8'h01;
  assign sel_10437 = array_index_10400 == array_index_10052 ? add_10436 : sel_10433;
  assign add_10440 = sel_10437 + 8'h01;
  assign out = {array_index_10400 == array_index_10058 ? add_10440 : sel_10437, {set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
