module min_hash(
  input wire [479:0] set1,
  input wire [479:0] set2,
  output wire [975:0] out
);
  wire [15:0] set1_unflattened[30];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  assign set1_unflattened[10] = set1[175:160];
  assign set1_unflattened[11] = set1[191:176];
  assign set1_unflattened[12] = set1[207:192];
  assign set1_unflattened[13] = set1[223:208];
  assign set1_unflattened[14] = set1[239:224];
  assign set1_unflattened[15] = set1[255:240];
  assign set1_unflattened[16] = set1[271:256];
  assign set1_unflattened[17] = set1[287:272];
  assign set1_unflattened[18] = set1[303:288];
  assign set1_unflattened[19] = set1[319:304];
  assign set1_unflattened[20] = set1[335:320];
  assign set1_unflattened[21] = set1[351:336];
  assign set1_unflattened[22] = set1[367:352];
  assign set1_unflattened[23] = set1[383:368];
  assign set1_unflattened[24] = set1[399:384];
  assign set1_unflattened[25] = set1[415:400];
  assign set1_unflattened[26] = set1[431:416];
  assign set1_unflattened[27] = set1[447:432];
  assign set1_unflattened[28] = set1[463:448];
  assign set1_unflattened[29] = set1[479:464];
  wire [15:0] set2_unflattened[30];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  assign set2_unflattened[10] = set2[175:160];
  assign set2_unflattened[11] = set2[191:176];
  assign set2_unflattened[12] = set2[207:192];
  assign set2_unflattened[13] = set2[223:208];
  assign set2_unflattened[14] = set2[239:224];
  assign set2_unflattened[15] = set2[255:240];
  assign set2_unflattened[16] = set2[271:256];
  assign set2_unflattened[17] = set2[287:272];
  assign set2_unflattened[18] = set2[303:288];
  assign set2_unflattened[19] = set2[319:304];
  assign set2_unflattened[20] = set2[335:320];
  assign set2_unflattened[21] = set2[351:336];
  assign set2_unflattened[22] = set2[367:352];
  assign set2_unflattened[23] = set2[383:368];
  assign set2_unflattened[24] = set2[399:384];
  assign set2_unflattened[25] = set2[415:400];
  assign set2_unflattened[26] = set2[431:416];
  assign set2_unflattened[27] = set2[447:432];
  assign set2_unflattened[28] = set2[463:448];
  assign set2_unflattened[29] = set2[479:464];
  wire [15:0] array_index_52563;
  wire [15:0] array_index_52564;
  wire [11:0] add_52571;
  wire [11:0] add_52574;
  wire [15:0] array_index_52579;
  wire [15:0] array_index_52582;
  wire [10:0] add_52586;
  wire [10:0] add_52589;
  wire [11:0] add_52605;
  wire [11:0] sel_52607;
  wire [11:0] add_52610;
  wire [11:0] sel_52612;
  wire [15:0] array_index_52627;
  wire [15:0] array_index_52630;
  wire [8:0] add_52634;
  wire [8:0] add_52637;
  wire [10:0] add_52640;
  wire [11:0] sel_52643;
  wire [10:0] add_52645;
  wire [11:0] sel_52648;
  wire [11:0] add_52665;
  wire [11:0] sel_52667;
  wire [11:0] add_52670;
  wire [11:0] sel_52672;
  wire [15:0] array_index_52693;
  wire [15:0] array_index_52696;
  wire [10:0] add_52700;
  wire [10:0] add_52702;
  wire [8:0] add_52704;
  wire [11:0] sel_52707;
  wire [8:0] add_52709;
  wire [11:0] sel_52712;
  wire [10:0] add_52714;
  wire [11:0] sel_52717;
  wire [10:0] add_52719;
  wire [11:0] sel_52722;
  wire [11:0] add_52743;
  wire [11:0] sel_52745;
  wire [11:0] add_52748;
  wire [11:0] sel_52750;
  wire [15:0] array_index_52777;
  wire [15:0] array_index_52780;
  wire [10:0] add_52784;
  wire [10:0] add_52786;
  wire [10:0] add_52788;
  wire [11:0] sel_52790;
  wire [10:0] add_52792;
  wire [11:0] sel_52794;
  wire [8:0] add_52796;
  wire [11:0] sel_52799;
  wire [8:0] add_52801;
  wire [11:0] sel_52804;
  wire [10:0] add_52806;
  wire [11:0] sel_52809;
  wire [10:0] add_52811;
  wire [11:0] sel_52814;
  wire [11:0] add_52839;
  wire [11:0] sel_52841;
  wire [11:0] add_52844;
  wire [11:0] sel_52846;
  wire [15:0] array_index_52877;
  wire [15:0] array_index_52880;
  wire [10:0] add_52884;
  wire [11:0] sel_52886;
  wire [10:0] add_52888;
  wire [11:0] sel_52890;
  wire [10:0] add_52892;
  wire [11:0] sel_52894;
  wire [10:0] add_52896;
  wire [11:0] sel_52898;
  wire [8:0] add_52900;
  wire [11:0] sel_52903;
  wire [8:0] add_52905;
  wire [11:0] sel_52908;
  wire [10:0] add_52910;
  wire [11:0] sel_52913;
  wire [10:0] add_52915;
  wire [11:0] sel_52918;
  wire [11:0] add_52943;
  wire [11:0] sel_52945;
  wire [11:0] add_52948;
  wire [11:0] sel_52950;
  wire [15:0] array_index_52979;
  wire [15:0] array_index_52982;
  wire [10:0] add_52986;
  wire [11:0] sel_52988;
  wire [10:0] add_52990;
  wire [11:0] sel_52992;
  wire [10:0] add_52994;
  wire [11:0] sel_52996;
  wire [10:0] add_52998;
  wire [11:0] sel_53000;
  wire [8:0] add_53002;
  wire [11:0] sel_53005;
  wire [8:0] add_53007;
  wire [11:0] sel_53010;
  wire [10:0] add_53012;
  wire [11:0] sel_53015;
  wire [10:0] add_53017;
  wire [11:0] sel_53020;
  wire [11:0] add_53045;
  wire [11:0] sel_53047;
  wire [11:0] add_53050;
  wire [11:0] sel_53052;
  wire [15:0] array_index_53081;
  wire [15:0] array_index_53084;
  wire [10:0] add_53088;
  wire [11:0] sel_53090;
  wire [10:0] add_53092;
  wire [11:0] sel_53094;
  wire [10:0] add_53096;
  wire [11:0] sel_53098;
  wire [10:0] add_53100;
  wire [11:0] sel_53102;
  wire [8:0] add_53104;
  wire [11:0] sel_53107;
  wire [8:0] add_53109;
  wire [11:0] sel_53112;
  wire [10:0] add_53114;
  wire [11:0] sel_53117;
  wire [10:0] add_53119;
  wire [11:0] sel_53122;
  wire [11:0] add_53147;
  wire [11:0] sel_53149;
  wire [11:0] add_53152;
  wire [11:0] sel_53154;
  wire [15:0] array_index_53183;
  wire [15:0] array_index_53186;
  wire [10:0] add_53190;
  wire [11:0] sel_53192;
  wire [10:0] add_53194;
  wire [11:0] sel_53196;
  wire [10:0] add_53198;
  wire [11:0] sel_53200;
  wire [10:0] add_53202;
  wire [11:0] sel_53204;
  wire [8:0] add_53206;
  wire [11:0] sel_53209;
  wire [8:0] add_53211;
  wire [11:0] sel_53214;
  wire [10:0] add_53216;
  wire [11:0] sel_53219;
  wire [10:0] add_53221;
  wire [11:0] sel_53224;
  wire [11:0] add_53249;
  wire [11:0] sel_53251;
  wire [11:0] add_53254;
  wire [11:0] sel_53256;
  wire [15:0] array_index_53285;
  wire [15:0] array_index_53288;
  wire [10:0] add_53292;
  wire [11:0] sel_53294;
  wire [10:0] add_53296;
  wire [11:0] sel_53298;
  wire [10:0] add_53300;
  wire [11:0] sel_53302;
  wire [10:0] add_53304;
  wire [11:0] sel_53306;
  wire [8:0] add_53308;
  wire [11:0] sel_53311;
  wire [8:0] add_53313;
  wire [11:0] sel_53316;
  wire [10:0] add_53318;
  wire [11:0] sel_53321;
  wire [10:0] add_53323;
  wire [11:0] sel_53326;
  wire [11:0] add_53351;
  wire [11:0] sel_53353;
  wire [11:0] add_53356;
  wire [11:0] sel_53358;
  wire [15:0] array_index_53387;
  wire [15:0] array_index_53390;
  wire [10:0] add_53394;
  wire [11:0] sel_53396;
  wire [10:0] add_53398;
  wire [11:0] sel_53400;
  wire [10:0] add_53402;
  wire [11:0] sel_53404;
  wire [10:0] add_53406;
  wire [11:0] sel_53408;
  wire [8:0] add_53410;
  wire [11:0] sel_53413;
  wire [8:0] add_53415;
  wire [11:0] sel_53418;
  wire [10:0] add_53420;
  wire [11:0] sel_53423;
  wire [10:0] add_53425;
  wire [11:0] sel_53428;
  wire [11:0] add_53453;
  wire [11:0] sel_53455;
  wire [11:0] add_53458;
  wire [11:0] sel_53460;
  wire [15:0] array_index_53489;
  wire [15:0] array_index_53492;
  wire [10:0] add_53496;
  wire [11:0] sel_53498;
  wire [10:0] add_53500;
  wire [11:0] sel_53502;
  wire [10:0] add_53504;
  wire [11:0] sel_53506;
  wire [10:0] add_53508;
  wire [11:0] sel_53510;
  wire [8:0] add_53512;
  wire [11:0] sel_53515;
  wire [8:0] add_53517;
  wire [11:0] sel_53520;
  wire [10:0] add_53522;
  wire [11:0] sel_53525;
  wire [10:0] add_53527;
  wire [11:0] sel_53530;
  wire [11:0] add_53555;
  wire [11:0] sel_53557;
  wire [11:0] add_53560;
  wire [11:0] sel_53562;
  wire [15:0] array_index_53591;
  wire [15:0] array_index_53594;
  wire [10:0] add_53598;
  wire [11:0] sel_53600;
  wire [10:0] add_53602;
  wire [11:0] sel_53604;
  wire [10:0] add_53606;
  wire [11:0] sel_53608;
  wire [10:0] add_53610;
  wire [11:0] sel_53612;
  wire [8:0] add_53614;
  wire [11:0] sel_53617;
  wire [8:0] add_53619;
  wire [11:0] sel_53622;
  wire [10:0] add_53624;
  wire [11:0] sel_53627;
  wire [10:0] add_53629;
  wire [11:0] sel_53632;
  wire [11:0] add_53657;
  wire [11:0] sel_53659;
  wire [11:0] add_53662;
  wire [11:0] sel_53664;
  wire [15:0] array_index_53693;
  wire [15:0] array_index_53696;
  wire [10:0] add_53700;
  wire [11:0] sel_53702;
  wire [10:0] add_53704;
  wire [11:0] sel_53706;
  wire [10:0] add_53708;
  wire [11:0] sel_53710;
  wire [10:0] add_53712;
  wire [11:0] sel_53714;
  wire [8:0] add_53716;
  wire [11:0] sel_53719;
  wire [8:0] add_53721;
  wire [11:0] sel_53724;
  wire [10:0] add_53726;
  wire [11:0] sel_53729;
  wire [10:0] add_53731;
  wire [11:0] sel_53734;
  wire [11:0] add_53759;
  wire [11:0] sel_53761;
  wire [11:0] add_53764;
  wire [11:0] sel_53766;
  wire [15:0] array_index_53795;
  wire [15:0] array_index_53798;
  wire [10:0] add_53802;
  wire [11:0] sel_53804;
  wire [10:0] add_53806;
  wire [11:0] sel_53808;
  wire [10:0] add_53810;
  wire [11:0] sel_53812;
  wire [10:0] add_53814;
  wire [11:0] sel_53816;
  wire [8:0] add_53818;
  wire [11:0] sel_53821;
  wire [8:0] add_53823;
  wire [11:0] sel_53826;
  wire [10:0] add_53828;
  wire [11:0] sel_53831;
  wire [10:0] add_53833;
  wire [11:0] sel_53836;
  wire [11:0] add_53861;
  wire [11:0] sel_53863;
  wire [11:0] add_53866;
  wire [11:0] sel_53868;
  wire [15:0] array_index_53897;
  wire [15:0] array_index_53900;
  wire [10:0] add_53904;
  wire [11:0] sel_53906;
  wire [10:0] add_53908;
  wire [11:0] sel_53910;
  wire [10:0] add_53912;
  wire [11:0] sel_53914;
  wire [10:0] add_53916;
  wire [11:0] sel_53918;
  wire [8:0] add_53920;
  wire [11:0] sel_53923;
  wire [8:0] add_53925;
  wire [11:0] sel_53928;
  wire [10:0] add_53930;
  wire [11:0] sel_53933;
  wire [10:0] add_53935;
  wire [11:0] sel_53938;
  wire [11:0] add_53963;
  wire [11:0] sel_53965;
  wire [11:0] add_53968;
  wire [11:0] sel_53970;
  wire [15:0] array_index_53999;
  wire [15:0] array_index_54002;
  wire [10:0] add_54006;
  wire [11:0] sel_54008;
  wire [10:0] add_54010;
  wire [11:0] sel_54012;
  wire [10:0] add_54014;
  wire [11:0] sel_54016;
  wire [10:0] add_54018;
  wire [11:0] sel_54020;
  wire [8:0] add_54022;
  wire [11:0] sel_54025;
  wire [8:0] add_54027;
  wire [11:0] sel_54030;
  wire [10:0] add_54032;
  wire [11:0] sel_54035;
  wire [10:0] add_54037;
  wire [11:0] sel_54040;
  wire [11:0] add_54065;
  wire [11:0] sel_54067;
  wire [11:0] add_54070;
  wire [11:0] sel_54072;
  wire [15:0] array_index_54101;
  wire [15:0] array_index_54104;
  wire [10:0] add_54108;
  wire [11:0] sel_54110;
  wire [10:0] add_54112;
  wire [11:0] sel_54114;
  wire [10:0] add_54116;
  wire [11:0] sel_54118;
  wire [10:0] add_54120;
  wire [11:0] sel_54122;
  wire [8:0] add_54124;
  wire [11:0] sel_54127;
  wire [8:0] add_54129;
  wire [11:0] sel_54132;
  wire [10:0] add_54134;
  wire [11:0] sel_54137;
  wire [10:0] add_54139;
  wire [11:0] sel_54142;
  wire [11:0] add_54167;
  wire [11:0] sel_54169;
  wire [11:0] add_54172;
  wire [11:0] sel_54174;
  wire [15:0] array_index_54203;
  wire [15:0] array_index_54206;
  wire [10:0] add_54210;
  wire [11:0] sel_54212;
  wire [10:0] add_54214;
  wire [11:0] sel_54216;
  wire [10:0] add_54218;
  wire [11:0] sel_54220;
  wire [10:0] add_54222;
  wire [11:0] sel_54224;
  wire [8:0] add_54226;
  wire [11:0] sel_54229;
  wire [8:0] add_54231;
  wire [11:0] sel_54234;
  wire [10:0] add_54236;
  wire [11:0] sel_54239;
  wire [10:0] add_54241;
  wire [11:0] sel_54244;
  wire [11:0] add_54269;
  wire [11:0] sel_54271;
  wire [11:0] add_54274;
  wire [11:0] sel_54276;
  wire [15:0] array_index_54305;
  wire [15:0] array_index_54308;
  wire [10:0] add_54312;
  wire [11:0] sel_54314;
  wire [10:0] add_54316;
  wire [11:0] sel_54318;
  wire [10:0] add_54320;
  wire [11:0] sel_54322;
  wire [10:0] add_54324;
  wire [11:0] sel_54326;
  wire [8:0] add_54328;
  wire [11:0] sel_54331;
  wire [8:0] add_54333;
  wire [11:0] sel_54336;
  wire [10:0] add_54338;
  wire [11:0] sel_54341;
  wire [10:0] add_54343;
  wire [11:0] sel_54346;
  wire [11:0] add_54371;
  wire [11:0] sel_54373;
  wire [11:0] add_54376;
  wire [11:0] sel_54378;
  wire [15:0] array_index_54407;
  wire [15:0] array_index_54410;
  wire [10:0] add_54414;
  wire [11:0] sel_54416;
  wire [10:0] add_54418;
  wire [11:0] sel_54420;
  wire [10:0] add_54422;
  wire [11:0] sel_54424;
  wire [10:0] add_54426;
  wire [11:0] sel_54428;
  wire [8:0] add_54430;
  wire [11:0] sel_54433;
  wire [8:0] add_54435;
  wire [11:0] sel_54438;
  wire [10:0] add_54440;
  wire [11:0] sel_54443;
  wire [10:0] add_54445;
  wire [11:0] sel_54448;
  wire [11:0] add_54473;
  wire [11:0] sel_54475;
  wire [11:0] add_54478;
  wire [11:0] sel_54480;
  wire [15:0] array_index_54509;
  wire [15:0] array_index_54512;
  wire [10:0] add_54516;
  wire [11:0] sel_54518;
  wire [10:0] add_54520;
  wire [11:0] sel_54522;
  wire [10:0] add_54524;
  wire [11:0] sel_54526;
  wire [10:0] add_54528;
  wire [11:0] sel_54530;
  wire [8:0] add_54532;
  wire [11:0] sel_54535;
  wire [8:0] add_54537;
  wire [11:0] sel_54540;
  wire [10:0] add_54542;
  wire [11:0] sel_54545;
  wire [10:0] add_54547;
  wire [11:0] sel_54550;
  wire [11:0] add_54575;
  wire [11:0] sel_54577;
  wire [11:0] add_54580;
  wire [11:0] sel_54582;
  wire [15:0] array_index_54611;
  wire [15:0] array_index_54614;
  wire [10:0] add_54618;
  wire [11:0] sel_54620;
  wire [10:0] add_54622;
  wire [11:0] sel_54624;
  wire [10:0] add_54626;
  wire [11:0] sel_54628;
  wire [10:0] add_54630;
  wire [11:0] sel_54632;
  wire [8:0] add_54634;
  wire [11:0] sel_54637;
  wire [8:0] add_54639;
  wire [11:0] sel_54642;
  wire [10:0] add_54644;
  wire [11:0] sel_54647;
  wire [10:0] add_54649;
  wire [11:0] sel_54652;
  wire [11:0] add_54677;
  wire [11:0] sel_54679;
  wire [11:0] add_54682;
  wire [11:0] sel_54684;
  wire [15:0] array_index_54713;
  wire [15:0] array_index_54716;
  wire [10:0] add_54720;
  wire [11:0] sel_54722;
  wire [10:0] add_54724;
  wire [11:0] sel_54726;
  wire [10:0] add_54728;
  wire [11:0] sel_54730;
  wire [10:0] add_54732;
  wire [11:0] sel_54734;
  wire [8:0] add_54736;
  wire [11:0] sel_54739;
  wire [8:0] add_54741;
  wire [11:0] sel_54744;
  wire [10:0] add_54746;
  wire [11:0] sel_54749;
  wire [10:0] add_54751;
  wire [11:0] sel_54754;
  wire [11:0] add_54779;
  wire [11:0] sel_54781;
  wire [11:0] add_54784;
  wire [11:0] sel_54786;
  wire [15:0] array_index_54815;
  wire [15:0] array_index_54818;
  wire [10:0] add_54822;
  wire [11:0] sel_54824;
  wire [10:0] add_54826;
  wire [11:0] sel_54828;
  wire [10:0] add_54830;
  wire [11:0] sel_54832;
  wire [10:0] add_54834;
  wire [11:0] sel_54836;
  wire [8:0] add_54838;
  wire [11:0] sel_54841;
  wire [8:0] add_54843;
  wire [11:0] sel_54846;
  wire [10:0] add_54848;
  wire [11:0] sel_54851;
  wire [10:0] add_54853;
  wire [11:0] sel_54856;
  wire [11:0] add_54881;
  wire [11:0] sel_54883;
  wire [11:0] add_54886;
  wire [11:0] sel_54888;
  wire [15:0] array_index_54917;
  wire [15:0] array_index_54920;
  wire [10:0] add_54924;
  wire [11:0] sel_54926;
  wire [10:0] add_54928;
  wire [11:0] sel_54930;
  wire [10:0] add_54932;
  wire [11:0] sel_54934;
  wire [10:0] add_54936;
  wire [11:0] sel_54938;
  wire [8:0] add_54940;
  wire [11:0] sel_54943;
  wire [8:0] add_54945;
  wire [11:0] sel_54948;
  wire [10:0] add_54950;
  wire [11:0] sel_54953;
  wire [10:0] add_54955;
  wire [11:0] sel_54958;
  wire [11:0] add_54983;
  wire [11:0] sel_54985;
  wire [11:0] add_54988;
  wire [11:0] sel_54990;
  wire [15:0] array_index_55019;
  wire [15:0] array_index_55022;
  wire [10:0] add_55026;
  wire [11:0] sel_55028;
  wire [10:0] add_55030;
  wire [11:0] sel_55032;
  wire [10:0] add_55034;
  wire [11:0] sel_55036;
  wire [10:0] add_55038;
  wire [11:0] sel_55040;
  wire [8:0] add_55042;
  wire [11:0] sel_55045;
  wire [8:0] add_55047;
  wire [11:0] sel_55050;
  wire [10:0] add_55052;
  wire [11:0] sel_55055;
  wire [10:0] add_55057;
  wire [11:0] sel_55060;
  wire [11:0] add_55085;
  wire [11:0] sel_55087;
  wire [11:0] add_55090;
  wire [11:0] sel_55092;
  wire [15:0] array_index_55121;
  wire [15:0] array_index_55124;
  wire [10:0] add_55128;
  wire [11:0] sel_55130;
  wire [10:0] add_55132;
  wire [11:0] sel_55134;
  wire [10:0] add_55136;
  wire [11:0] sel_55138;
  wire [10:0] add_55140;
  wire [11:0] sel_55142;
  wire [8:0] add_55144;
  wire [11:0] sel_55147;
  wire [8:0] add_55149;
  wire [11:0] sel_55152;
  wire [10:0] add_55154;
  wire [11:0] sel_55157;
  wire [10:0] add_55159;
  wire [11:0] sel_55162;
  wire [11:0] add_55187;
  wire [11:0] sel_55189;
  wire [11:0] add_55192;
  wire [11:0] sel_55194;
  wire [15:0] array_index_55223;
  wire [15:0] array_index_55226;
  wire [10:0] add_55230;
  wire [11:0] sel_55232;
  wire [10:0] add_55234;
  wire [11:0] sel_55236;
  wire [10:0] add_55238;
  wire [11:0] sel_55240;
  wire [10:0] add_55242;
  wire [11:0] sel_55244;
  wire [8:0] add_55246;
  wire [11:0] sel_55249;
  wire [8:0] add_55251;
  wire [11:0] sel_55254;
  wire [10:0] add_55256;
  wire [11:0] sel_55259;
  wire [10:0] add_55261;
  wire [11:0] sel_55264;
  wire [11:0] add_55289;
  wire [11:0] sel_55291;
  wire [11:0] add_55294;
  wire [11:0] sel_55296;
  wire [15:0] array_index_55325;
  wire [15:0] array_index_55328;
  wire [10:0] add_55332;
  wire [11:0] sel_55334;
  wire [10:0] add_55336;
  wire [11:0] sel_55338;
  wire [10:0] add_55340;
  wire [11:0] sel_55342;
  wire [10:0] add_55344;
  wire [11:0] sel_55346;
  wire [8:0] add_55348;
  wire [11:0] sel_55351;
  wire [8:0] add_55353;
  wire [11:0] sel_55356;
  wire [10:0] add_55358;
  wire [11:0] sel_55361;
  wire [10:0] add_55363;
  wire [11:0] sel_55366;
  wire [11:0] add_55390;
  wire [11:0] sel_55392;
  wire [11:0] add_55394;
  wire [11:0] sel_55396;
  wire [10:0] add_55430;
  wire [11:0] sel_55432;
  wire [10:0] add_55434;
  wire [11:0] sel_55436;
  wire [10:0] add_55438;
  wire [11:0] sel_55440;
  wire [10:0] add_55442;
  wire [11:0] sel_55444;
  wire [8:0] add_55446;
  wire [11:0] sel_55449;
  wire [8:0] add_55451;
  wire [11:0] sel_55454;
  wire [10:0] add_55456;
  wire [11:0] sel_55459;
  wire [10:0] add_55461;
  wire [11:0] sel_55464;
  wire [10:0] add_55512;
  wire [11:0] sel_55514;
  wire [10:0] add_55516;
  wire [11:0] sel_55518;
  wire [10:0] add_55520;
  wire [11:0] sel_55522;
  wire [10:0] add_55524;
  wire [11:0] sel_55526;
  wire [8:0] add_55528;
  wire [11:0] sel_55531;
  wire [8:0] add_55533;
  wire [11:0] sel_55536;
  wire [1:0] concat_55539;
  wire [1:0] add_55554;
  wire [10:0] add_55574;
  wire [11:0] sel_55576;
  wire [10:0] add_55578;
  wire [11:0] sel_55580;
  wire [10:0] add_55582;
  wire [11:0] sel_55584;
  wire [10:0] add_55586;
  wire [11:0] sel_55588;
  wire [2:0] concat_55591;
  wire [2:0] add_55602;
  wire [10:0] add_55616;
  wire [11:0] sel_55618;
  wire [10:0] add_55620;
  wire [11:0] sel_55622;
  wire [3:0] concat_55625;
  wire [3:0] add_55632;
  wire [4:0] concat_55641;
  wire [4:0] add_55644;
  assign array_index_52563 = set1_unflattened[5'h00];
  assign array_index_52564 = set2_unflattened[5'h00];
  assign add_52571 = array_index_52563[11:0] + 12'h247;
  assign add_52574 = array_index_52564[11:0] + 12'h247;
  assign array_index_52579 = set1_unflattened[5'h01];
  assign array_index_52582 = set2_unflattened[5'h01];
  assign add_52586 = array_index_52563[11:1] + 11'h247;
  assign add_52589 = array_index_52564[11:1] + 11'h247;
  assign add_52605 = array_index_52579[11:0] + 12'h247;
  assign sel_52607 = $signed({1'h0, add_52571}) < $signed(13'h0fff) ? add_52571 : 12'hfff;
  assign add_52610 = array_index_52582[11:0] + 12'h247;
  assign sel_52612 = $signed({1'h0, add_52574}) < $signed(13'h0fff) ? add_52574 : 12'hfff;
  assign array_index_52627 = set1_unflattened[5'h02];
  assign array_index_52630 = set2_unflattened[5'h02];
  assign add_52634 = array_index_52563[11:3] + 9'h0bd;
  assign add_52637 = array_index_52564[11:3] + 9'h0bd;
  assign add_52640 = array_index_52579[11:1] + 11'h247;
  assign sel_52643 = $signed({1'h0, add_52586, array_index_52563[0]}) < $signed(13'h0fff) ? {add_52586, array_index_52563[0]} : 12'hfff;
  assign add_52645 = array_index_52582[11:1] + 11'h247;
  assign sel_52648 = $signed({1'h0, add_52589, array_index_52564[0]}) < $signed(13'h0fff) ? {add_52589, array_index_52564[0]} : 12'hfff;
  assign add_52665 = array_index_52627[11:0] + 12'h247;
  assign sel_52667 = $signed({1'h0, add_52605}) < $signed({1'h0, sel_52607}) ? add_52605 : sel_52607;
  assign add_52670 = array_index_52630[11:0] + 12'h247;
  assign sel_52672 = $signed({1'h0, add_52610}) < $signed({1'h0, sel_52612}) ? add_52610 : sel_52612;
  assign array_index_52693 = set1_unflattened[5'h03];
  assign array_index_52696 = set2_unflattened[5'h03];
  assign add_52700 = array_index_52563[11:1] + 11'h347;
  assign add_52702 = array_index_52564[11:1] + 11'h347;
  assign add_52704 = array_index_52579[11:3] + 9'h0bd;
  assign sel_52707 = $signed({1'h0, add_52634, array_index_52563[2:0]}) < $signed(13'h0fff) ? {add_52634, array_index_52563[2:0]} : 12'hfff;
  assign add_52709 = array_index_52582[11:3] + 9'h0bd;
  assign sel_52712 = $signed({1'h0, add_52637, array_index_52564[2:0]}) < $signed(13'h0fff) ? {add_52637, array_index_52564[2:0]} : 12'hfff;
  assign add_52714 = array_index_52627[11:1] + 11'h247;
  assign sel_52717 = $signed({1'h0, add_52640, array_index_52579[0]}) < $signed({1'h0, sel_52643}) ? {add_52640, array_index_52579[0]} : sel_52643;
  assign add_52719 = array_index_52630[11:1] + 11'h247;
  assign sel_52722 = $signed({1'h0, add_52645, array_index_52582[0]}) < $signed({1'h0, sel_52648}) ? {add_52645, array_index_52582[0]} : sel_52648;
  assign add_52743 = array_index_52693[11:0] + 12'h247;
  assign sel_52745 = $signed({1'h0, add_52665}) < $signed({1'h0, sel_52667}) ? add_52665 : sel_52667;
  assign add_52748 = array_index_52696[11:0] + 12'h247;
  assign sel_52750 = $signed({1'h0, add_52670}) < $signed({1'h0, sel_52672}) ? add_52670 : sel_52672;
  assign array_index_52777 = set1_unflattened[5'h04];
  assign array_index_52780 = set2_unflattened[5'h04];
  assign add_52784 = array_index_52563[11:1] + 11'h79d;
  assign add_52786 = array_index_52564[11:1] + 11'h79d;
  assign add_52788 = array_index_52579[11:1] + 11'h347;
  assign sel_52790 = $signed({1'h0, add_52700, array_index_52563[0]}) < $signed(13'h0fff) ? {add_52700, array_index_52563[0]} : 12'hfff;
  assign add_52792 = array_index_52582[11:1] + 11'h347;
  assign sel_52794 = $signed({1'h0, add_52702, array_index_52564[0]}) < $signed(13'h0fff) ? {add_52702, array_index_52564[0]} : 12'hfff;
  assign add_52796 = array_index_52627[11:3] + 9'h0bd;
  assign sel_52799 = $signed({1'h0, add_52704, array_index_52579[2:0]}) < $signed({1'h0, sel_52707}) ? {add_52704, array_index_52579[2:0]} : sel_52707;
  assign add_52801 = array_index_52630[11:3] + 9'h0bd;
  assign sel_52804 = $signed({1'h0, add_52709, array_index_52582[2:0]}) < $signed({1'h0, sel_52712}) ? {add_52709, array_index_52582[2:0]} : sel_52712;
  assign add_52806 = array_index_52693[11:1] + 11'h247;
  assign sel_52809 = $signed({1'h0, add_52714, array_index_52627[0]}) < $signed({1'h0, sel_52717}) ? {add_52714, array_index_52627[0]} : sel_52717;
  assign add_52811 = array_index_52696[11:1] + 11'h247;
  assign sel_52814 = $signed({1'h0, add_52719, array_index_52630[0]}) < $signed({1'h0, sel_52722}) ? {add_52719, array_index_52630[0]} : sel_52722;
  assign add_52839 = array_index_52777[11:0] + 12'h247;
  assign sel_52841 = $signed({1'h0, add_52743}) < $signed({1'h0, sel_52745}) ? add_52743 : sel_52745;
  assign add_52844 = array_index_52780[11:0] + 12'h247;
  assign sel_52846 = $signed({1'h0, add_52748}) < $signed({1'h0, sel_52750}) ? add_52748 : sel_52750;
  assign array_index_52877 = set1_unflattened[5'h05];
  assign array_index_52880 = set2_unflattened[5'h05];
  assign add_52884 = array_index_52579[11:1] + 11'h79d;
  assign sel_52886 = $signed({1'h0, add_52784, array_index_52563[0]}) < $signed(13'h0fff) ? {add_52784, array_index_52563[0]} : 12'hfff;
  assign add_52888 = array_index_52582[11:1] + 11'h79d;
  assign sel_52890 = $signed({1'h0, add_52786, array_index_52564[0]}) < $signed(13'h0fff) ? {add_52786, array_index_52564[0]} : 12'hfff;
  assign add_52892 = array_index_52627[11:1] + 11'h347;
  assign sel_52894 = $signed({1'h0, add_52788, array_index_52579[0]}) < $signed({1'h0, sel_52790}) ? {add_52788, array_index_52579[0]} : sel_52790;
  assign add_52896 = array_index_52630[11:1] + 11'h347;
  assign sel_52898 = $signed({1'h0, add_52792, array_index_52582[0]}) < $signed({1'h0, sel_52794}) ? {add_52792, array_index_52582[0]} : sel_52794;
  assign add_52900 = array_index_52693[11:3] + 9'h0bd;
  assign sel_52903 = $signed({1'h0, add_52796, array_index_52627[2:0]}) < $signed({1'h0, sel_52799}) ? {add_52796, array_index_52627[2:0]} : sel_52799;
  assign add_52905 = array_index_52696[11:3] + 9'h0bd;
  assign sel_52908 = $signed({1'h0, add_52801, array_index_52630[2:0]}) < $signed({1'h0, sel_52804}) ? {add_52801, array_index_52630[2:0]} : sel_52804;
  assign add_52910 = array_index_52777[11:1] + 11'h247;
  assign sel_52913 = $signed({1'h0, add_52806, array_index_52693[0]}) < $signed({1'h0, sel_52809}) ? {add_52806, array_index_52693[0]} : sel_52809;
  assign add_52915 = array_index_52780[11:1] + 11'h247;
  assign sel_52918 = $signed({1'h0, add_52811, array_index_52696[0]}) < $signed({1'h0, sel_52814}) ? {add_52811, array_index_52696[0]} : sel_52814;
  assign add_52943 = array_index_52877[11:0] + 12'h247;
  assign sel_52945 = $signed({1'h0, add_52839}) < $signed({1'h0, sel_52841}) ? add_52839 : sel_52841;
  assign add_52948 = array_index_52880[11:0] + 12'h247;
  assign sel_52950 = $signed({1'h0, add_52844}) < $signed({1'h0, sel_52846}) ? add_52844 : sel_52846;
  assign array_index_52979 = set1_unflattened[5'h06];
  assign array_index_52982 = set2_unflattened[5'h06];
  assign add_52986 = array_index_52627[11:1] + 11'h79d;
  assign sel_52988 = $signed({1'h0, add_52884, array_index_52579[0]}) < $signed({1'h0, sel_52886}) ? {add_52884, array_index_52579[0]} : sel_52886;
  assign add_52990 = array_index_52630[11:1] + 11'h79d;
  assign sel_52992 = $signed({1'h0, add_52888, array_index_52582[0]}) < $signed({1'h0, sel_52890}) ? {add_52888, array_index_52582[0]} : sel_52890;
  assign add_52994 = array_index_52693[11:1] + 11'h347;
  assign sel_52996 = $signed({1'h0, add_52892, array_index_52627[0]}) < $signed({1'h0, sel_52894}) ? {add_52892, array_index_52627[0]} : sel_52894;
  assign add_52998 = array_index_52696[11:1] + 11'h347;
  assign sel_53000 = $signed({1'h0, add_52896, array_index_52630[0]}) < $signed({1'h0, sel_52898}) ? {add_52896, array_index_52630[0]} : sel_52898;
  assign add_53002 = array_index_52777[11:3] + 9'h0bd;
  assign sel_53005 = $signed({1'h0, add_52900, array_index_52693[2:0]}) < $signed({1'h0, sel_52903}) ? {add_52900, array_index_52693[2:0]} : sel_52903;
  assign add_53007 = array_index_52780[11:3] + 9'h0bd;
  assign sel_53010 = $signed({1'h0, add_52905, array_index_52696[2:0]}) < $signed({1'h0, sel_52908}) ? {add_52905, array_index_52696[2:0]} : sel_52908;
  assign add_53012 = array_index_52877[11:1] + 11'h247;
  assign sel_53015 = $signed({1'h0, add_52910, array_index_52777[0]}) < $signed({1'h0, sel_52913}) ? {add_52910, array_index_52777[0]} : sel_52913;
  assign add_53017 = array_index_52880[11:1] + 11'h247;
  assign sel_53020 = $signed({1'h0, add_52915, array_index_52780[0]}) < $signed({1'h0, sel_52918}) ? {add_52915, array_index_52780[0]} : sel_52918;
  assign add_53045 = array_index_52979[11:0] + 12'h247;
  assign sel_53047 = $signed({1'h0, add_52943}) < $signed({1'h0, sel_52945}) ? add_52943 : sel_52945;
  assign add_53050 = array_index_52982[11:0] + 12'h247;
  assign sel_53052 = $signed({1'h0, add_52948}) < $signed({1'h0, sel_52950}) ? add_52948 : sel_52950;
  assign array_index_53081 = set1_unflattened[5'h07];
  assign array_index_53084 = set2_unflattened[5'h07];
  assign add_53088 = array_index_52693[11:1] + 11'h79d;
  assign sel_53090 = $signed({1'h0, add_52986, array_index_52627[0]}) < $signed({1'h0, sel_52988}) ? {add_52986, array_index_52627[0]} : sel_52988;
  assign add_53092 = array_index_52696[11:1] + 11'h79d;
  assign sel_53094 = $signed({1'h0, add_52990, array_index_52630[0]}) < $signed({1'h0, sel_52992}) ? {add_52990, array_index_52630[0]} : sel_52992;
  assign add_53096 = array_index_52777[11:1] + 11'h347;
  assign sel_53098 = $signed({1'h0, add_52994, array_index_52693[0]}) < $signed({1'h0, sel_52996}) ? {add_52994, array_index_52693[0]} : sel_52996;
  assign add_53100 = array_index_52780[11:1] + 11'h347;
  assign sel_53102 = $signed({1'h0, add_52998, array_index_52696[0]}) < $signed({1'h0, sel_53000}) ? {add_52998, array_index_52696[0]} : sel_53000;
  assign add_53104 = array_index_52877[11:3] + 9'h0bd;
  assign sel_53107 = $signed({1'h0, add_53002, array_index_52777[2:0]}) < $signed({1'h0, sel_53005}) ? {add_53002, array_index_52777[2:0]} : sel_53005;
  assign add_53109 = array_index_52880[11:3] + 9'h0bd;
  assign sel_53112 = $signed({1'h0, add_53007, array_index_52780[2:0]}) < $signed({1'h0, sel_53010}) ? {add_53007, array_index_52780[2:0]} : sel_53010;
  assign add_53114 = array_index_52979[11:1] + 11'h247;
  assign sel_53117 = $signed({1'h0, add_53012, array_index_52877[0]}) < $signed({1'h0, sel_53015}) ? {add_53012, array_index_52877[0]} : sel_53015;
  assign add_53119 = array_index_52982[11:1] + 11'h247;
  assign sel_53122 = $signed({1'h0, add_53017, array_index_52880[0]}) < $signed({1'h0, sel_53020}) ? {add_53017, array_index_52880[0]} : sel_53020;
  assign add_53147 = array_index_53081[11:0] + 12'h247;
  assign sel_53149 = $signed({1'h0, add_53045}) < $signed({1'h0, sel_53047}) ? add_53045 : sel_53047;
  assign add_53152 = array_index_53084[11:0] + 12'h247;
  assign sel_53154 = $signed({1'h0, add_53050}) < $signed({1'h0, sel_53052}) ? add_53050 : sel_53052;
  assign array_index_53183 = set1_unflattened[5'h08];
  assign array_index_53186 = set2_unflattened[5'h08];
  assign add_53190 = array_index_52777[11:1] + 11'h79d;
  assign sel_53192 = $signed({1'h0, add_53088, array_index_52693[0]}) < $signed({1'h0, sel_53090}) ? {add_53088, array_index_52693[0]} : sel_53090;
  assign add_53194 = array_index_52780[11:1] + 11'h79d;
  assign sel_53196 = $signed({1'h0, add_53092, array_index_52696[0]}) < $signed({1'h0, sel_53094}) ? {add_53092, array_index_52696[0]} : sel_53094;
  assign add_53198 = array_index_52877[11:1] + 11'h347;
  assign sel_53200 = $signed({1'h0, add_53096, array_index_52777[0]}) < $signed({1'h0, sel_53098}) ? {add_53096, array_index_52777[0]} : sel_53098;
  assign add_53202 = array_index_52880[11:1] + 11'h347;
  assign sel_53204 = $signed({1'h0, add_53100, array_index_52780[0]}) < $signed({1'h0, sel_53102}) ? {add_53100, array_index_52780[0]} : sel_53102;
  assign add_53206 = array_index_52979[11:3] + 9'h0bd;
  assign sel_53209 = $signed({1'h0, add_53104, array_index_52877[2:0]}) < $signed({1'h0, sel_53107}) ? {add_53104, array_index_52877[2:0]} : sel_53107;
  assign add_53211 = array_index_52982[11:3] + 9'h0bd;
  assign sel_53214 = $signed({1'h0, add_53109, array_index_52880[2:0]}) < $signed({1'h0, sel_53112}) ? {add_53109, array_index_52880[2:0]} : sel_53112;
  assign add_53216 = array_index_53081[11:1] + 11'h247;
  assign sel_53219 = $signed({1'h0, add_53114, array_index_52979[0]}) < $signed({1'h0, sel_53117}) ? {add_53114, array_index_52979[0]} : sel_53117;
  assign add_53221 = array_index_53084[11:1] + 11'h247;
  assign sel_53224 = $signed({1'h0, add_53119, array_index_52982[0]}) < $signed({1'h0, sel_53122}) ? {add_53119, array_index_52982[0]} : sel_53122;
  assign add_53249 = array_index_53183[11:0] + 12'h247;
  assign sel_53251 = $signed({1'h0, add_53147}) < $signed({1'h0, sel_53149}) ? add_53147 : sel_53149;
  assign add_53254 = array_index_53186[11:0] + 12'h247;
  assign sel_53256 = $signed({1'h0, add_53152}) < $signed({1'h0, sel_53154}) ? add_53152 : sel_53154;
  assign array_index_53285 = set1_unflattened[5'h09];
  assign array_index_53288 = set2_unflattened[5'h09];
  assign add_53292 = array_index_52877[11:1] + 11'h79d;
  assign sel_53294 = $signed({1'h0, add_53190, array_index_52777[0]}) < $signed({1'h0, sel_53192}) ? {add_53190, array_index_52777[0]} : sel_53192;
  assign add_53296 = array_index_52880[11:1] + 11'h79d;
  assign sel_53298 = $signed({1'h0, add_53194, array_index_52780[0]}) < $signed({1'h0, sel_53196}) ? {add_53194, array_index_52780[0]} : sel_53196;
  assign add_53300 = array_index_52979[11:1] + 11'h347;
  assign sel_53302 = $signed({1'h0, add_53198, array_index_52877[0]}) < $signed({1'h0, sel_53200}) ? {add_53198, array_index_52877[0]} : sel_53200;
  assign add_53304 = array_index_52982[11:1] + 11'h347;
  assign sel_53306 = $signed({1'h0, add_53202, array_index_52880[0]}) < $signed({1'h0, sel_53204}) ? {add_53202, array_index_52880[0]} : sel_53204;
  assign add_53308 = array_index_53081[11:3] + 9'h0bd;
  assign sel_53311 = $signed({1'h0, add_53206, array_index_52979[2:0]}) < $signed({1'h0, sel_53209}) ? {add_53206, array_index_52979[2:0]} : sel_53209;
  assign add_53313 = array_index_53084[11:3] + 9'h0bd;
  assign sel_53316 = $signed({1'h0, add_53211, array_index_52982[2:0]}) < $signed({1'h0, sel_53214}) ? {add_53211, array_index_52982[2:0]} : sel_53214;
  assign add_53318 = array_index_53183[11:1] + 11'h247;
  assign sel_53321 = $signed({1'h0, add_53216, array_index_53081[0]}) < $signed({1'h0, sel_53219}) ? {add_53216, array_index_53081[0]} : sel_53219;
  assign add_53323 = array_index_53186[11:1] + 11'h247;
  assign sel_53326 = $signed({1'h0, add_53221, array_index_53084[0]}) < $signed({1'h0, sel_53224}) ? {add_53221, array_index_53084[0]} : sel_53224;
  assign add_53351 = array_index_53285[11:0] + 12'h247;
  assign sel_53353 = $signed({1'h0, add_53249}) < $signed({1'h0, sel_53251}) ? add_53249 : sel_53251;
  assign add_53356 = array_index_53288[11:0] + 12'h247;
  assign sel_53358 = $signed({1'h0, add_53254}) < $signed({1'h0, sel_53256}) ? add_53254 : sel_53256;
  assign array_index_53387 = set1_unflattened[5'h0a];
  assign array_index_53390 = set2_unflattened[5'h0a];
  assign add_53394 = array_index_52979[11:1] + 11'h79d;
  assign sel_53396 = $signed({1'h0, add_53292, array_index_52877[0]}) < $signed({1'h0, sel_53294}) ? {add_53292, array_index_52877[0]} : sel_53294;
  assign add_53398 = array_index_52982[11:1] + 11'h79d;
  assign sel_53400 = $signed({1'h0, add_53296, array_index_52880[0]}) < $signed({1'h0, sel_53298}) ? {add_53296, array_index_52880[0]} : sel_53298;
  assign add_53402 = array_index_53081[11:1] + 11'h347;
  assign sel_53404 = $signed({1'h0, add_53300, array_index_52979[0]}) < $signed({1'h0, sel_53302}) ? {add_53300, array_index_52979[0]} : sel_53302;
  assign add_53406 = array_index_53084[11:1] + 11'h347;
  assign sel_53408 = $signed({1'h0, add_53304, array_index_52982[0]}) < $signed({1'h0, sel_53306}) ? {add_53304, array_index_52982[0]} : sel_53306;
  assign add_53410 = array_index_53183[11:3] + 9'h0bd;
  assign sel_53413 = $signed({1'h0, add_53308, array_index_53081[2:0]}) < $signed({1'h0, sel_53311}) ? {add_53308, array_index_53081[2:0]} : sel_53311;
  assign add_53415 = array_index_53186[11:3] + 9'h0bd;
  assign sel_53418 = $signed({1'h0, add_53313, array_index_53084[2:0]}) < $signed({1'h0, sel_53316}) ? {add_53313, array_index_53084[2:0]} : sel_53316;
  assign add_53420 = array_index_53285[11:1] + 11'h247;
  assign sel_53423 = $signed({1'h0, add_53318, array_index_53183[0]}) < $signed({1'h0, sel_53321}) ? {add_53318, array_index_53183[0]} : sel_53321;
  assign add_53425 = array_index_53288[11:1] + 11'h247;
  assign sel_53428 = $signed({1'h0, add_53323, array_index_53186[0]}) < $signed({1'h0, sel_53326}) ? {add_53323, array_index_53186[0]} : sel_53326;
  assign add_53453 = array_index_53387[11:0] + 12'h247;
  assign sel_53455 = $signed({1'h0, add_53351}) < $signed({1'h0, sel_53353}) ? add_53351 : sel_53353;
  assign add_53458 = array_index_53390[11:0] + 12'h247;
  assign sel_53460 = $signed({1'h0, add_53356}) < $signed({1'h0, sel_53358}) ? add_53356 : sel_53358;
  assign array_index_53489 = set1_unflattened[5'h0b];
  assign array_index_53492 = set2_unflattened[5'h0b];
  assign add_53496 = array_index_53081[11:1] + 11'h79d;
  assign sel_53498 = $signed({1'h0, add_53394, array_index_52979[0]}) < $signed({1'h0, sel_53396}) ? {add_53394, array_index_52979[0]} : sel_53396;
  assign add_53500 = array_index_53084[11:1] + 11'h79d;
  assign sel_53502 = $signed({1'h0, add_53398, array_index_52982[0]}) < $signed({1'h0, sel_53400}) ? {add_53398, array_index_52982[0]} : sel_53400;
  assign add_53504 = array_index_53183[11:1] + 11'h347;
  assign sel_53506 = $signed({1'h0, add_53402, array_index_53081[0]}) < $signed({1'h0, sel_53404}) ? {add_53402, array_index_53081[0]} : sel_53404;
  assign add_53508 = array_index_53186[11:1] + 11'h347;
  assign sel_53510 = $signed({1'h0, add_53406, array_index_53084[0]}) < $signed({1'h0, sel_53408}) ? {add_53406, array_index_53084[0]} : sel_53408;
  assign add_53512 = array_index_53285[11:3] + 9'h0bd;
  assign sel_53515 = $signed({1'h0, add_53410, array_index_53183[2:0]}) < $signed({1'h0, sel_53413}) ? {add_53410, array_index_53183[2:0]} : sel_53413;
  assign add_53517 = array_index_53288[11:3] + 9'h0bd;
  assign sel_53520 = $signed({1'h0, add_53415, array_index_53186[2:0]}) < $signed({1'h0, sel_53418}) ? {add_53415, array_index_53186[2:0]} : sel_53418;
  assign add_53522 = array_index_53387[11:1] + 11'h247;
  assign sel_53525 = $signed({1'h0, add_53420, array_index_53285[0]}) < $signed({1'h0, sel_53423}) ? {add_53420, array_index_53285[0]} : sel_53423;
  assign add_53527 = array_index_53390[11:1] + 11'h247;
  assign sel_53530 = $signed({1'h0, add_53425, array_index_53288[0]}) < $signed({1'h0, sel_53428}) ? {add_53425, array_index_53288[0]} : sel_53428;
  assign add_53555 = array_index_53489[11:0] + 12'h247;
  assign sel_53557 = $signed({1'h0, add_53453}) < $signed({1'h0, sel_53455}) ? add_53453 : sel_53455;
  assign add_53560 = array_index_53492[11:0] + 12'h247;
  assign sel_53562 = $signed({1'h0, add_53458}) < $signed({1'h0, sel_53460}) ? add_53458 : sel_53460;
  assign array_index_53591 = set1_unflattened[5'h0c];
  assign array_index_53594 = set2_unflattened[5'h0c];
  assign add_53598 = array_index_53183[11:1] + 11'h79d;
  assign sel_53600 = $signed({1'h0, add_53496, array_index_53081[0]}) < $signed({1'h0, sel_53498}) ? {add_53496, array_index_53081[0]} : sel_53498;
  assign add_53602 = array_index_53186[11:1] + 11'h79d;
  assign sel_53604 = $signed({1'h0, add_53500, array_index_53084[0]}) < $signed({1'h0, sel_53502}) ? {add_53500, array_index_53084[0]} : sel_53502;
  assign add_53606 = array_index_53285[11:1] + 11'h347;
  assign sel_53608 = $signed({1'h0, add_53504, array_index_53183[0]}) < $signed({1'h0, sel_53506}) ? {add_53504, array_index_53183[0]} : sel_53506;
  assign add_53610 = array_index_53288[11:1] + 11'h347;
  assign sel_53612 = $signed({1'h0, add_53508, array_index_53186[0]}) < $signed({1'h0, sel_53510}) ? {add_53508, array_index_53186[0]} : sel_53510;
  assign add_53614 = array_index_53387[11:3] + 9'h0bd;
  assign sel_53617 = $signed({1'h0, add_53512, array_index_53285[2:0]}) < $signed({1'h0, sel_53515}) ? {add_53512, array_index_53285[2:0]} : sel_53515;
  assign add_53619 = array_index_53390[11:3] + 9'h0bd;
  assign sel_53622 = $signed({1'h0, add_53517, array_index_53288[2:0]}) < $signed({1'h0, sel_53520}) ? {add_53517, array_index_53288[2:0]} : sel_53520;
  assign add_53624 = array_index_53489[11:1] + 11'h247;
  assign sel_53627 = $signed({1'h0, add_53522, array_index_53387[0]}) < $signed({1'h0, sel_53525}) ? {add_53522, array_index_53387[0]} : sel_53525;
  assign add_53629 = array_index_53492[11:1] + 11'h247;
  assign sel_53632 = $signed({1'h0, add_53527, array_index_53390[0]}) < $signed({1'h0, sel_53530}) ? {add_53527, array_index_53390[0]} : sel_53530;
  assign add_53657 = array_index_53591[11:0] + 12'h247;
  assign sel_53659 = $signed({1'h0, add_53555}) < $signed({1'h0, sel_53557}) ? add_53555 : sel_53557;
  assign add_53662 = array_index_53594[11:0] + 12'h247;
  assign sel_53664 = $signed({1'h0, add_53560}) < $signed({1'h0, sel_53562}) ? add_53560 : sel_53562;
  assign array_index_53693 = set1_unflattened[5'h0d];
  assign array_index_53696 = set2_unflattened[5'h0d];
  assign add_53700 = array_index_53285[11:1] + 11'h79d;
  assign sel_53702 = $signed({1'h0, add_53598, array_index_53183[0]}) < $signed({1'h0, sel_53600}) ? {add_53598, array_index_53183[0]} : sel_53600;
  assign add_53704 = array_index_53288[11:1] + 11'h79d;
  assign sel_53706 = $signed({1'h0, add_53602, array_index_53186[0]}) < $signed({1'h0, sel_53604}) ? {add_53602, array_index_53186[0]} : sel_53604;
  assign add_53708 = array_index_53387[11:1] + 11'h347;
  assign sel_53710 = $signed({1'h0, add_53606, array_index_53285[0]}) < $signed({1'h0, sel_53608}) ? {add_53606, array_index_53285[0]} : sel_53608;
  assign add_53712 = array_index_53390[11:1] + 11'h347;
  assign sel_53714 = $signed({1'h0, add_53610, array_index_53288[0]}) < $signed({1'h0, sel_53612}) ? {add_53610, array_index_53288[0]} : sel_53612;
  assign add_53716 = array_index_53489[11:3] + 9'h0bd;
  assign sel_53719 = $signed({1'h0, add_53614, array_index_53387[2:0]}) < $signed({1'h0, sel_53617}) ? {add_53614, array_index_53387[2:0]} : sel_53617;
  assign add_53721 = array_index_53492[11:3] + 9'h0bd;
  assign sel_53724 = $signed({1'h0, add_53619, array_index_53390[2:0]}) < $signed({1'h0, sel_53622}) ? {add_53619, array_index_53390[2:0]} : sel_53622;
  assign add_53726 = array_index_53591[11:1] + 11'h247;
  assign sel_53729 = $signed({1'h0, add_53624, array_index_53489[0]}) < $signed({1'h0, sel_53627}) ? {add_53624, array_index_53489[0]} : sel_53627;
  assign add_53731 = array_index_53594[11:1] + 11'h247;
  assign sel_53734 = $signed({1'h0, add_53629, array_index_53492[0]}) < $signed({1'h0, sel_53632}) ? {add_53629, array_index_53492[0]} : sel_53632;
  assign add_53759 = array_index_53693[11:0] + 12'h247;
  assign sel_53761 = $signed({1'h0, add_53657}) < $signed({1'h0, sel_53659}) ? add_53657 : sel_53659;
  assign add_53764 = array_index_53696[11:0] + 12'h247;
  assign sel_53766 = $signed({1'h0, add_53662}) < $signed({1'h0, sel_53664}) ? add_53662 : sel_53664;
  assign array_index_53795 = set1_unflattened[5'h0e];
  assign array_index_53798 = set2_unflattened[5'h0e];
  assign add_53802 = array_index_53387[11:1] + 11'h79d;
  assign sel_53804 = $signed({1'h0, add_53700, array_index_53285[0]}) < $signed({1'h0, sel_53702}) ? {add_53700, array_index_53285[0]} : sel_53702;
  assign add_53806 = array_index_53390[11:1] + 11'h79d;
  assign sel_53808 = $signed({1'h0, add_53704, array_index_53288[0]}) < $signed({1'h0, sel_53706}) ? {add_53704, array_index_53288[0]} : sel_53706;
  assign add_53810 = array_index_53489[11:1] + 11'h347;
  assign sel_53812 = $signed({1'h0, add_53708, array_index_53387[0]}) < $signed({1'h0, sel_53710}) ? {add_53708, array_index_53387[0]} : sel_53710;
  assign add_53814 = array_index_53492[11:1] + 11'h347;
  assign sel_53816 = $signed({1'h0, add_53712, array_index_53390[0]}) < $signed({1'h0, sel_53714}) ? {add_53712, array_index_53390[0]} : sel_53714;
  assign add_53818 = array_index_53591[11:3] + 9'h0bd;
  assign sel_53821 = $signed({1'h0, add_53716, array_index_53489[2:0]}) < $signed({1'h0, sel_53719}) ? {add_53716, array_index_53489[2:0]} : sel_53719;
  assign add_53823 = array_index_53594[11:3] + 9'h0bd;
  assign sel_53826 = $signed({1'h0, add_53721, array_index_53492[2:0]}) < $signed({1'h0, sel_53724}) ? {add_53721, array_index_53492[2:0]} : sel_53724;
  assign add_53828 = array_index_53693[11:1] + 11'h247;
  assign sel_53831 = $signed({1'h0, add_53726, array_index_53591[0]}) < $signed({1'h0, sel_53729}) ? {add_53726, array_index_53591[0]} : sel_53729;
  assign add_53833 = array_index_53696[11:1] + 11'h247;
  assign sel_53836 = $signed({1'h0, add_53731, array_index_53594[0]}) < $signed({1'h0, sel_53734}) ? {add_53731, array_index_53594[0]} : sel_53734;
  assign add_53861 = array_index_53795[11:0] + 12'h247;
  assign sel_53863 = $signed({1'h0, add_53759}) < $signed({1'h0, sel_53761}) ? add_53759 : sel_53761;
  assign add_53866 = array_index_53798[11:0] + 12'h247;
  assign sel_53868 = $signed({1'h0, add_53764}) < $signed({1'h0, sel_53766}) ? add_53764 : sel_53766;
  assign array_index_53897 = set1_unflattened[5'h0f];
  assign array_index_53900 = set2_unflattened[5'h0f];
  assign add_53904 = array_index_53489[11:1] + 11'h79d;
  assign sel_53906 = $signed({1'h0, add_53802, array_index_53387[0]}) < $signed({1'h0, sel_53804}) ? {add_53802, array_index_53387[0]} : sel_53804;
  assign add_53908 = array_index_53492[11:1] + 11'h79d;
  assign sel_53910 = $signed({1'h0, add_53806, array_index_53390[0]}) < $signed({1'h0, sel_53808}) ? {add_53806, array_index_53390[0]} : sel_53808;
  assign add_53912 = array_index_53591[11:1] + 11'h347;
  assign sel_53914 = $signed({1'h0, add_53810, array_index_53489[0]}) < $signed({1'h0, sel_53812}) ? {add_53810, array_index_53489[0]} : sel_53812;
  assign add_53916 = array_index_53594[11:1] + 11'h347;
  assign sel_53918 = $signed({1'h0, add_53814, array_index_53492[0]}) < $signed({1'h0, sel_53816}) ? {add_53814, array_index_53492[0]} : sel_53816;
  assign add_53920 = array_index_53693[11:3] + 9'h0bd;
  assign sel_53923 = $signed({1'h0, add_53818, array_index_53591[2:0]}) < $signed({1'h0, sel_53821}) ? {add_53818, array_index_53591[2:0]} : sel_53821;
  assign add_53925 = array_index_53696[11:3] + 9'h0bd;
  assign sel_53928 = $signed({1'h0, add_53823, array_index_53594[2:0]}) < $signed({1'h0, sel_53826}) ? {add_53823, array_index_53594[2:0]} : sel_53826;
  assign add_53930 = array_index_53795[11:1] + 11'h247;
  assign sel_53933 = $signed({1'h0, add_53828, array_index_53693[0]}) < $signed({1'h0, sel_53831}) ? {add_53828, array_index_53693[0]} : sel_53831;
  assign add_53935 = array_index_53798[11:1] + 11'h247;
  assign sel_53938 = $signed({1'h0, add_53833, array_index_53696[0]}) < $signed({1'h0, sel_53836}) ? {add_53833, array_index_53696[0]} : sel_53836;
  assign add_53963 = array_index_53897[11:0] + 12'h247;
  assign sel_53965 = $signed({1'h0, add_53861}) < $signed({1'h0, sel_53863}) ? add_53861 : sel_53863;
  assign add_53968 = array_index_53900[11:0] + 12'h247;
  assign sel_53970 = $signed({1'h0, add_53866}) < $signed({1'h0, sel_53868}) ? add_53866 : sel_53868;
  assign array_index_53999 = set1_unflattened[5'h10];
  assign array_index_54002 = set2_unflattened[5'h10];
  assign add_54006 = array_index_53591[11:1] + 11'h79d;
  assign sel_54008 = $signed({1'h0, add_53904, array_index_53489[0]}) < $signed({1'h0, sel_53906}) ? {add_53904, array_index_53489[0]} : sel_53906;
  assign add_54010 = array_index_53594[11:1] + 11'h79d;
  assign sel_54012 = $signed({1'h0, add_53908, array_index_53492[0]}) < $signed({1'h0, sel_53910}) ? {add_53908, array_index_53492[0]} : sel_53910;
  assign add_54014 = array_index_53693[11:1] + 11'h347;
  assign sel_54016 = $signed({1'h0, add_53912, array_index_53591[0]}) < $signed({1'h0, sel_53914}) ? {add_53912, array_index_53591[0]} : sel_53914;
  assign add_54018 = array_index_53696[11:1] + 11'h347;
  assign sel_54020 = $signed({1'h0, add_53916, array_index_53594[0]}) < $signed({1'h0, sel_53918}) ? {add_53916, array_index_53594[0]} : sel_53918;
  assign add_54022 = array_index_53795[11:3] + 9'h0bd;
  assign sel_54025 = $signed({1'h0, add_53920, array_index_53693[2:0]}) < $signed({1'h0, sel_53923}) ? {add_53920, array_index_53693[2:0]} : sel_53923;
  assign add_54027 = array_index_53798[11:3] + 9'h0bd;
  assign sel_54030 = $signed({1'h0, add_53925, array_index_53696[2:0]}) < $signed({1'h0, sel_53928}) ? {add_53925, array_index_53696[2:0]} : sel_53928;
  assign add_54032 = array_index_53897[11:1] + 11'h247;
  assign sel_54035 = $signed({1'h0, add_53930, array_index_53795[0]}) < $signed({1'h0, sel_53933}) ? {add_53930, array_index_53795[0]} : sel_53933;
  assign add_54037 = array_index_53900[11:1] + 11'h247;
  assign sel_54040 = $signed({1'h0, add_53935, array_index_53798[0]}) < $signed({1'h0, sel_53938}) ? {add_53935, array_index_53798[0]} : sel_53938;
  assign add_54065 = array_index_53999[11:0] + 12'h247;
  assign sel_54067 = $signed({1'h0, add_53963}) < $signed({1'h0, sel_53965}) ? add_53963 : sel_53965;
  assign add_54070 = array_index_54002[11:0] + 12'h247;
  assign sel_54072 = $signed({1'h0, add_53968}) < $signed({1'h0, sel_53970}) ? add_53968 : sel_53970;
  assign array_index_54101 = set1_unflattened[5'h11];
  assign array_index_54104 = set2_unflattened[5'h11];
  assign add_54108 = array_index_53693[11:1] + 11'h79d;
  assign sel_54110 = $signed({1'h0, add_54006, array_index_53591[0]}) < $signed({1'h0, sel_54008}) ? {add_54006, array_index_53591[0]} : sel_54008;
  assign add_54112 = array_index_53696[11:1] + 11'h79d;
  assign sel_54114 = $signed({1'h0, add_54010, array_index_53594[0]}) < $signed({1'h0, sel_54012}) ? {add_54010, array_index_53594[0]} : sel_54012;
  assign add_54116 = array_index_53795[11:1] + 11'h347;
  assign sel_54118 = $signed({1'h0, add_54014, array_index_53693[0]}) < $signed({1'h0, sel_54016}) ? {add_54014, array_index_53693[0]} : sel_54016;
  assign add_54120 = array_index_53798[11:1] + 11'h347;
  assign sel_54122 = $signed({1'h0, add_54018, array_index_53696[0]}) < $signed({1'h0, sel_54020}) ? {add_54018, array_index_53696[0]} : sel_54020;
  assign add_54124 = array_index_53897[11:3] + 9'h0bd;
  assign sel_54127 = $signed({1'h0, add_54022, array_index_53795[2:0]}) < $signed({1'h0, sel_54025}) ? {add_54022, array_index_53795[2:0]} : sel_54025;
  assign add_54129 = array_index_53900[11:3] + 9'h0bd;
  assign sel_54132 = $signed({1'h0, add_54027, array_index_53798[2:0]}) < $signed({1'h0, sel_54030}) ? {add_54027, array_index_53798[2:0]} : sel_54030;
  assign add_54134 = array_index_53999[11:1] + 11'h247;
  assign sel_54137 = $signed({1'h0, add_54032, array_index_53897[0]}) < $signed({1'h0, sel_54035}) ? {add_54032, array_index_53897[0]} : sel_54035;
  assign add_54139 = array_index_54002[11:1] + 11'h247;
  assign sel_54142 = $signed({1'h0, add_54037, array_index_53900[0]}) < $signed({1'h0, sel_54040}) ? {add_54037, array_index_53900[0]} : sel_54040;
  assign add_54167 = array_index_54101[11:0] + 12'h247;
  assign sel_54169 = $signed({1'h0, add_54065}) < $signed({1'h0, sel_54067}) ? add_54065 : sel_54067;
  assign add_54172 = array_index_54104[11:0] + 12'h247;
  assign sel_54174 = $signed({1'h0, add_54070}) < $signed({1'h0, sel_54072}) ? add_54070 : sel_54072;
  assign array_index_54203 = set1_unflattened[5'h12];
  assign array_index_54206 = set2_unflattened[5'h12];
  assign add_54210 = array_index_53795[11:1] + 11'h79d;
  assign sel_54212 = $signed({1'h0, add_54108, array_index_53693[0]}) < $signed({1'h0, sel_54110}) ? {add_54108, array_index_53693[0]} : sel_54110;
  assign add_54214 = array_index_53798[11:1] + 11'h79d;
  assign sel_54216 = $signed({1'h0, add_54112, array_index_53696[0]}) < $signed({1'h0, sel_54114}) ? {add_54112, array_index_53696[0]} : sel_54114;
  assign add_54218 = array_index_53897[11:1] + 11'h347;
  assign sel_54220 = $signed({1'h0, add_54116, array_index_53795[0]}) < $signed({1'h0, sel_54118}) ? {add_54116, array_index_53795[0]} : sel_54118;
  assign add_54222 = array_index_53900[11:1] + 11'h347;
  assign sel_54224 = $signed({1'h0, add_54120, array_index_53798[0]}) < $signed({1'h0, sel_54122}) ? {add_54120, array_index_53798[0]} : sel_54122;
  assign add_54226 = array_index_53999[11:3] + 9'h0bd;
  assign sel_54229 = $signed({1'h0, add_54124, array_index_53897[2:0]}) < $signed({1'h0, sel_54127}) ? {add_54124, array_index_53897[2:0]} : sel_54127;
  assign add_54231 = array_index_54002[11:3] + 9'h0bd;
  assign sel_54234 = $signed({1'h0, add_54129, array_index_53900[2:0]}) < $signed({1'h0, sel_54132}) ? {add_54129, array_index_53900[2:0]} : sel_54132;
  assign add_54236 = array_index_54101[11:1] + 11'h247;
  assign sel_54239 = $signed({1'h0, add_54134, array_index_53999[0]}) < $signed({1'h0, sel_54137}) ? {add_54134, array_index_53999[0]} : sel_54137;
  assign add_54241 = array_index_54104[11:1] + 11'h247;
  assign sel_54244 = $signed({1'h0, add_54139, array_index_54002[0]}) < $signed({1'h0, sel_54142}) ? {add_54139, array_index_54002[0]} : sel_54142;
  assign add_54269 = array_index_54203[11:0] + 12'h247;
  assign sel_54271 = $signed({1'h0, add_54167}) < $signed({1'h0, sel_54169}) ? add_54167 : sel_54169;
  assign add_54274 = array_index_54206[11:0] + 12'h247;
  assign sel_54276 = $signed({1'h0, add_54172}) < $signed({1'h0, sel_54174}) ? add_54172 : sel_54174;
  assign array_index_54305 = set1_unflattened[5'h13];
  assign array_index_54308 = set2_unflattened[5'h13];
  assign add_54312 = array_index_53897[11:1] + 11'h79d;
  assign sel_54314 = $signed({1'h0, add_54210, array_index_53795[0]}) < $signed({1'h0, sel_54212}) ? {add_54210, array_index_53795[0]} : sel_54212;
  assign add_54316 = array_index_53900[11:1] + 11'h79d;
  assign sel_54318 = $signed({1'h0, add_54214, array_index_53798[0]}) < $signed({1'h0, sel_54216}) ? {add_54214, array_index_53798[0]} : sel_54216;
  assign add_54320 = array_index_53999[11:1] + 11'h347;
  assign sel_54322 = $signed({1'h0, add_54218, array_index_53897[0]}) < $signed({1'h0, sel_54220}) ? {add_54218, array_index_53897[0]} : sel_54220;
  assign add_54324 = array_index_54002[11:1] + 11'h347;
  assign sel_54326 = $signed({1'h0, add_54222, array_index_53900[0]}) < $signed({1'h0, sel_54224}) ? {add_54222, array_index_53900[0]} : sel_54224;
  assign add_54328 = array_index_54101[11:3] + 9'h0bd;
  assign sel_54331 = $signed({1'h0, add_54226, array_index_53999[2:0]}) < $signed({1'h0, sel_54229}) ? {add_54226, array_index_53999[2:0]} : sel_54229;
  assign add_54333 = array_index_54104[11:3] + 9'h0bd;
  assign sel_54336 = $signed({1'h0, add_54231, array_index_54002[2:0]}) < $signed({1'h0, sel_54234}) ? {add_54231, array_index_54002[2:0]} : sel_54234;
  assign add_54338 = array_index_54203[11:1] + 11'h247;
  assign sel_54341 = $signed({1'h0, add_54236, array_index_54101[0]}) < $signed({1'h0, sel_54239}) ? {add_54236, array_index_54101[0]} : sel_54239;
  assign add_54343 = array_index_54206[11:1] + 11'h247;
  assign sel_54346 = $signed({1'h0, add_54241, array_index_54104[0]}) < $signed({1'h0, sel_54244}) ? {add_54241, array_index_54104[0]} : sel_54244;
  assign add_54371 = array_index_54305[11:0] + 12'h247;
  assign sel_54373 = $signed({1'h0, add_54269}) < $signed({1'h0, sel_54271}) ? add_54269 : sel_54271;
  assign add_54376 = array_index_54308[11:0] + 12'h247;
  assign sel_54378 = $signed({1'h0, add_54274}) < $signed({1'h0, sel_54276}) ? add_54274 : sel_54276;
  assign array_index_54407 = set1_unflattened[5'h14];
  assign array_index_54410 = set2_unflattened[5'h14];
  assign add_54414 = array_index_53999[11:1] + 11'h79d;
  assign sel_54416 = $signed({1'h0, add_54312, array_index_53897[0]}) < $signed({1'h0, sel_54314}) ? {add_54312, array_index_53897[0]} : sel_54314;
  assign add_54418 = array_index_54002[11:1] + 11'h79d;
  assign sel_54420 = $signed({1'h0, add_54316, array_index_53900[0]}) < $signed({1'h0, sel_54318}) ? {add_54316, array_index_53900[0]} : sel_54318;
  assign add_54422 = array_index_54101[11:1] + 11'h347;
  assign sel_54424 = $signed({1'h0, add_54320, array_index_53999[0]}) < $signed({1'h0, sel_54322}) ? {add_54320, array_index_53999[0]} : sel_54322;
  assign add_54426 = array_index_54104[11:1] + 11'h347;
  assign sel_54428 = $signed({1'h0, add_54324, array_index_54002[0]}) < $signed({1'h0, sel_54326}) ? {add_54324, array_index_54002[0]} : sel_54326;
  assign add_54430 = array_index_54203[11:3] + 9'h0bd;
  assign sel_54433 = $signed({1'h0, add_54328, array_index_54101[2:0]}) < $signed({1'h0, sel_54331}) ? {add_54328, array_index_54101[2:0]} : sel_54331;
  assign add_54435 = array_index_54206[11:3] + 9'h0bd;
  assign sel_54438 = $signed({1'h0, add_54333, array_index_54104[2:0]}) < $signed({1'h0, sel_54336}) ? {add_54333, array_index_54104[2:0]} : sel_54336;
  assign add_54440 = array_index_54305[11:1] + 11'h247;
  assign sel_54443 = $signed({1'h0, add_54338, array_index_54203[0]}) < $signed({1'h0, sel_54341}) ? {add_54338, array_index_54203[0]} : sel_54341;
  assign add_54445 = array_index_54308[11:1] + 11'h247;
  assign sel_54448 = $signed({1'h0, add_54343, array_index_54206[0]}) < $signed({1'h0, sel_54346}) ? {add_54343, array_index_54206[0]} : sel_54346;
  assign add_54473 = array_index_54407[11:0] + 12'h247;
  assign sel_54475 = $signed({1'h0, add_54371}) < $signed({1'h0, sel_54373}) ? add_54371 : sel_54373;
  assign add_54478 = array_index_54410[11:0] + 12'h247;
  assign sel_54480 = $signed({1'h0, add_54376}) < $signed({1'h0, sel_54378}) ? add_54376 : sel_54378;
  assign array_index_54509 = set1_unflattened[5'h15];
  assign array_index_54512 = set2_unflattened[5'h15];
  assign add_54516 = array_index_54101[11:1] + 11'h79d;
  assign sel_54518 = $signed({1'h0, add_54414, array_index_53999[0]}) < $signed({1'h0, sel_54416}) ? {add_54414, array_index_53999[0]} : sel_54416;
  assign add_54520 = array_index_54104[11:1] + 11'h79d;
  assign sel_54522 = $signed({1'h0, add_54418, array_index_54002[0]}) < $signed({1'h0, sel_54420}) ? {add_54418, array_index_54002[0]} : sel_54420;
  assign add_54524 = array_index_54203[11:1] + 11'h347;
  assign sel_54526 = $signed({1'h0, add_54422, array_index_54101[0]}) < $signed({1'h0, sel_54424}) ? {add_54422, array_index_54101[0]} : sel_54424;
  assign add_54528 = array_index_54206[11:1] + 11'h347;
  assign sel_54530 = $signed({1'h0, add_54426, array_index_54104[0]}) < $signed({1'h0, sel_54428}) ? {add_54426, array_index_54104[0]} : sel_54428;
  assign add_54532 = array_index_54305[11:3] + 9'h0bd;
  assign sel_54535 = $signed({1'h0, add_54430, array_index_54203[2:0]}) < $signed({1'h0, sel_54433}) ? {add_54430, array_index_54203[2:0]} : sel_54433;
  assign add_54537 = array_index_54308[11:3] + 9'h0bd;
  assign sel_54540 = $signed({1'h0, add_54435, array_index_54206[2:0]}) < $signed({1'h0, sel_54438}) ? {add_54435, array_index_54206[2:0]} : sel_54438;
  assign add_54542 = array_index_54407[11:1] + 11'h247;
  assign sel_54545 = $signed({1'h0, add_54440, array_index_54305[0]}) < $signed({1'h0, sel_54443}) ? {add_54440, array_index_54305[0]} : sel_54443;
  assign add_54547 = array_index_54410[11:1] + 11'h247;
  assign sel_54550 = $signed({1'h0, add_54445, array_index_54308[0]}) < $signed({1'h0, sel_54448}) ? {add_54445, array_index_54308[0]} : sel_54448;
  assign add_54575 = array_index_54509[11:0] + 12'h247;
  assign sel_54577 = $signed({1'h0, add_54473}) < $signed({1'h0, sel_54475}) ? add_54473 : sel_54475;
  assign add_54580 = array_index_54512[11:0] + 12'h247;
  assign sel_54582 = $signed({1'h0, add_54478}) < $signed({1'h0, sel_54480}) ? add_54478 : sel_54480;
  assign array_index_54611 = set1_unflattened[5'h16];
  assign array_index_54614 = set2_unflattened[5'h16];
  assign add_54618 = array_index_54203[11:1] + 11'h79d;
  assign sel_54620 = $signed({1'h0, add_54516, array_index_54101[0]}) < $signed({1'h0, sel_54518}) ? {add_54516, array_index_54101[0]} : sel_54518;
  assign add_54622 = array_index_54206[11:1] + 11'h79d;
  assign sel_54624 = $signed({1'h0, add_54520, array_index_54104[0]}) < $signed({1'h0, sel_54522}) ? {add_54520, array_index_54104[0]} : sel_54522;
  assign add_54626 = array_index_54305[11:1] + 11'h347;
  assign sel_54628 = $signed({1'h0, add_54524, array_index_54203[0]}) < $signed({1'h0, sel_54526}) ? {add_54524, array_index_54203[0]} : sel_54526;
  assign add_54630 = array_index_54308[11:1] + 11'h347;
  assign sel_54632 = $signed({1'h0, add_54528, array_index_54206[0]}) < $signed({1'h0, sel_54530}) ? {add_54528, array_index_54206[0]} : sel_54530;
  assign add_54634 = array_index_54407[11:3] + 9'h0bd;
  assign sel_54637 = $signed({1'h0, add_54532, array_index_54305[2:0]}) < $signed({1'h0, sel_54535}) ? {add_54532, array_index_54305[2:0]} : sel_54535;
  assign add_54639 = array_index_54410[11:3] + 9'h0bd;
  assign sel_54642 = $signed({1'h0, add_54537, array_index_54308[2:0]}) < $signed({1'h0, sel_54540}) ? {add_54537, array_index_54308[2:0]} : sel_54540;
  assign add_54644 = array_index_54509[11:1] + 11'h247;
  assign sel_54647 = $signed({1'h0, add_54542, array_index_54407[0]}) < $signed({1'h0, sel_54545}) ? {add_54542, array_index_54407[0]} : sel_54545;
  assign add_54649 = array_index_54512[11:1] + 11'h247;
  assign sel_54652 = $signed({1'h0, add_54547, array_index_54410[0]}) < $signed({1'h0, sel_54550}) ? {add_54547, array_index_54410[0]} : sel_54550;
  assign add_54677 = array_index_54611[11:0] + 12'h247;
  assign sel_54679 = $signed({1'h0, add_54575}) < $signed({1'h0, sel_54577}) ? add_54575 : sel_54577;
  assign add_54682 = array_index_54614[11:0] + 12'h247;
  assign sel_54684 = $signed({1'h0, add_54580}) < $signed({1'h0, sel_54582}) ? add_54580 : sel_54582;
  assign array_index_54713 = set1_unflattened[5'h17];
  assign array_index_54716 = set2_unflattened[5'h17];
  assign add_54720 = array_index_54305[11:1] + 11'h79d;
  assign sel_54722 = $signed({1'h0, add_54618, array_index_54203[0]}) < $signed({1'h0, sel_54620}) ? {add_54618, array_index_54203[0]} : sel_54620;
  assign add_54724 = array_index_54308[11:1] + 11'h79d;
  assign sel_54726 = $signed({1'h0, add_54622, array_index_54206[0]}) < $signed({1'h0, sel_54624}) ? {add_54622, array_index_54206[0]} : sel_54624;
  assign add_54728 = array_index_54407[11:1] + 11'h347;
  assign sel_54730 = $signed({1'h0, add_54626, array_index_54305[0]}) < $signed({1'h0, sel_54628}) ? {add_54626, array_index_54305[0]} : sel_54628;
  assign add_54732 = array_index_54410[11:1] + 11'h347;
  assign sel_54734 = $signed({1'h0, add_54630, array_index_54308[0]}) < $signed({1'h0, sel_54632}) ? {add_54630, array_index_54308[0]} : sel_54632;
  assign add_54736 = array_index_54509[11:3] + 9'h0bd;
  assign sel_54739 = $signed({1'h0, add_54634, array_index_54407[2:0]}) < $signed({1'h0, sel_54637}) ? {add_54634, array_index_54407[2:0]} : sel_54637;
  assign add_54741 = array_index_54512[11:3] + 9'h0bd;
  assign sel_54744 = $signed({1'h0, add_54639, array_index_54410[2:0]}) < $signed({1'h0, sel_54642}) ? {add_54639, array_index_54410[2:0]} : sel_54642;
  assign add_54746 = array_index_54611[11:1] + 11'h247;
  assign sel_54749 = $signed({1'h0, add_54644, array_index_54509[0]}) < $signed({1'h0, sel_54647}) ? {add_54644, array_index_54509[0]} : sel_54647;
  assign add_54751 = array_index_54614[11:1] + 11'h247;
  assign sel_54754 = $signed({1'h0, add_54649, array_index_54512[0]}) < $signed({1'h0, sel_54652}) ? {add_54649, array_index_54512[0]} : sel_54652;
  assign add_54779 = array_index_54713[11:0] + 12'h247;
  assign sel_54781 = $signed({1'h0, add_54677}) < $signed({1'h0, sel_54679}) ? add_54677 : sel_54679;
  assign add_54784 = array_index_54716[11:0] + 12'h247;
  assign sel_54786 = $signed({1'h0, add_54682}) < $signed({1'h0, sel_54684}) ? add_54682 : sel_54684;
  assign array_index_54815 = set1_unflattened[5'h18];
  assign array_index_54818 = set2_unflattened[5'h18];
  assign add_54822 = array_index_54407[11:1] + 11'h79d;
  assign sel_54824 = $signed({1'h0, add_54720, array_index_54305[0]}) < $signed({1'h0, sel_54722}) ? {add_54720, array_index_54305[0]} : sel_54722;
  assign add_54826 = array_index_54410[11:1] + 11'h79d;
  assign sel_54828 = $signed({1'h0, add_54724, array_index_54308[0]}) < $signed({1'h0, sel_54726}) ? {add_54724, array_index_54308[0]} : sel_54726;
  assign add_54830 = array_index_54509[11:1] + 11'h347;
  assign sel_54832 = $signed({1'h0, add_54728, array_index_54407[0]}) < $signed({1'h0, sel_54730}) ? {add_54728, array_index_54407[0]} : sel_54730;
  assign add_54834 = array_index_54512[11:1] + 11'h347;
  assign sel_54836 = $signed({1'h0, add_54732, array_index_54410[0]}) < $signed({1'h0, sel_54734}) ? {add_54732, array_index_54410[0]} : sel_54734;
  assign add_54838 = array_index_54611[11:3] + 9'h0bd;
  assign sel_54841 = $signed({1'h0, add_54736, array_index_54509[2:0]}) < $signed({1'h0, sel_54739}) ? {add_54736, array_index_54509[2:0]} : sel_54739;
  assign add_54843 = array_index_54614[11:3] + 9'h0bd;
  assign sel_54846 = $signed({1'h0, add_54741, array_index_54512[2:0]}) < $signed({1'h0, sel_54744}) ? {add_54741, array_index_54512[2:0]} : sel_54744;
  assign add_54848 = array_index_54713[11:1] + 11'h247;
  assign sel_54851 = $signed({1'h0, add_54746, array_index_54611[0]}) < $signed({1'h0, sel_54749}) ? {add_54746, array_index_54611[0]} : sel_54749;
  assign add_54853 = array_index_54716[11:1] + 11'h247;
  assign sel_54856 = $signed({1'h0, add_54751, array_index_54614[0]}) < $signed({1'h0, sel_54754}) ? {add_54751, array_index_54614[0]} : sel_54754;
  assign add_54881 = array_index_54815[11:0] + 12'h247;
  assign sel_54883 = $signed({1'h0, add_54779}) < $signed({1'h0, sel_54781}) ? add_54779 : sel_54781;
  assign add_54886 = array_index_54818[11:0] + 12'h247;
  assign sel_54888 = $signed({1'h0, add_54784}) < $signed({1'h0, sel_54786}) ? add_54784 : sel_54786;
  assign array_index_54917 = set1_unflattened[5'h19];
  assign array_index_54920 = set2_unflattened[5'h19];
  assign add_54924 = array_index_54509[11:1] + 11'h79d;
  assign sel_54926 = $signed({1'h0, add_54822, array_index_54407[0]}) < $signed({1'h0, sel_54824}) ? {add_54822, array_index_54407[0]} : sel_54824;
  assign add_54928 = array_index_54512[11:1] + 11'h79d;
  assign sel_54930 = $signed({1'h0, add_54826, array_index_54410[0]}) < $signed({1'h0, sel_54828}) ? {add_54826, array_index_54410[0]} : sel_54828;
  assign add_54932 = array_index_54611[11:1] + 11'h347;
  assign sel_54934 = $signed({1'h0, add_54830, array_index_54509[0]}) < $signed({1'h0, sel_54832}) ? {add_54830, array_index_54509[0]} : sel_54832;
  assign add_54936 = array_index_54614[11:1] + 11'h347;
  assign sel_54938 = $signed({1'h0, add_54834, array_index_54512[0]}) < $signed({1'h0, sel_54836}) ? {add_54834, array_index_54512[0]} : sel_54836;
  assign add_54940 = array_index_54713[11:3] + 9'h0bd;
  assign sel_54943 = $signed({1'h0, add_54838, array_index_54611[2:0]}) < $signed({1'h0, sel_54841}) ? {add_54838, array_index_54611[2:0]} : sel_54841;
  assign add_54945 = array_index_54716[11:3] + 9'h0bd;
  assign sel_54948 = $signed({1'h0, add_54843, array_index_54614[2:0]}) < $signed({1'h0, sel_54846}) ? {add_54843, array_index_54614[2:0]} : sel_54846;
  assign add_54950 = array_index_54815[11:1] + 11'h247;
  assign sel_54953 = $signed({1'h0, add_54848, array_index_54713[0]}) < $signed({1'h0, sel_54851}) ? {add_54848, array_index_54713[0]} : sel_54851;
  assign add_54955 = array_index_54818[11:1] + 11'h247;
  assign sel_54958 = $signed({1'h0, add_54853, array_index_54716[0]}) < $signed({1'h0, sel_54856}) ? {add_54853, array_index_54716[0]} : sel_54856;
  assign add_54983 = array_index_54917[11:0] + 12'h247;
  assign sel_54985 = $signed({1'h0, add_54881}) < $signed({1'h0, sel_54883}) ? add_54881 : sel_54883;
  assign add_54988 = array_index_54920[11:0] + 12'h247;
  assign sel_54990 = $signed({1'h0, add_54886}) < $signed({1'h0, sel_54888}) ? add_54886 : sel_54888;
  assign array_index_55019 = set1_unflattened[5'h1a];
  assign array_index_55022 = set2_unflattened[5'h1a];
  assign add_55026 = array_index_54611[11:1] + 11'h79d;
  assign sel_55028 = $signed({1'h0, add_54924, array_index_54509[0]}) < $signed({1'h0, sel_54926}) ? {add_54924, array_index_54509[0]} : sel_54926;
  assign add_55030 = array_index_54614[11:1] + 11'h79d;
  assign sel_55032 = $signed({1'h0, add_54928, array_index_54512[0]}) < $signed({1'h0, sel_54930}) ? {add_54928, array_index_54512[0]} : sel_54930;
  assign add_55034 = array_index_54713[11:1] + 11'h347;
  assign sel_55036 = $signed({1'h0, add_54932, array_index_54611[0]}) < $signed({1'h0, sel_54934}) ? {add_54932, array_index_54611[0]} : sel_54934;
  assign add_55038 = array_index_54716[11:1] + 11'h347;
  assign sel_55040 = $signed({1'h0, add_54936, array_index_54614[0]}) < $signed({1'h0, sel_54938}) ? {add_54936, array_index_54614[0]} : sel_54938;
  assign add_55042 = array_index_54815[11:3] + 9'h0bd;
  assign sel_55045 = $signed({1'h0, add_54940, array_index_54713[2:0]}) < $signed({1'h0, sel_54943}) ? {add_54940, array_index_54713[2:0]} : sel_54943;
  assign add_55047 = array_index_54818[11:3] + 9'h0bd;
  assign sel_55050 = $signed({1'h0, add_54945, array_index_54716[2:0]}) < $signed({1'h0, sel_54948}) ? {add_54945, array_index_54716[2:0]} : sel_54948;
  assign add_55052 = array_index_54917[11:1] + 11'h247;
  assign sel_55055 = $signed({1'h0, add_54950, array_index_54815[0]}) < $signed({1'h0, sel_54953}) ? {add_54950, array_index_54815[0]} : sel_54953;
  assign add_55057 = array_index_54920[11:1] + 11'h247;
  assign sel_55060 = $signed({1'h0, add_54955, array_index_54818[0]}) < $signed({1'h0, sel_54958}) ? {add_54955, array_index_54818[0]} : sel_54958;
  assign add_55085 = array_index_55019[11:0] + 12'h247;
  assign sel_55087 = $signed({1'h0, add_54983}) < $signed({1'h0, sel_54985}) ? add_54983 : sel_54985;
  assign add_55090 = array_index_55022[11:0] + 12'h247;
  assign sel_55092 = $signed({1'h0, add_54988}) < $signed({1'h0, sel_54990}) ? add_54988 : sel_54990;
  assign array_index_55121 = set1_unflattened[5'h1b];
  assign array_index_55124 = set2_unflattened[5'h1b];
  assign add_55128 = array_index_54713[11:1] + 11'h79d;
  assign sel_55130 = $signed({1'h0, add_55026, array_index_54611[0]}) < $signed({1'h0, sel_55028}) ? {add_55026, array_index_54611[0]} : sel_55028;
  assign add_55132 = array_index_54716[11:1] + 11'h79d;
  assign sel_55134 = $signed({1'h0, add_55030, array_index_54614[0]}) < $signed({1'h0, sel_55032}) ? {add_55030, array_index_54614[0]} : sel_55032;
  assign add_55136 = array_index_54815[11:1] + 11'h347;
  assign sel_55138 = $signed({1'h0, add_55034, array_index_54713[0]}) < $signed({1'h0, sel_55036}) ? {add_55034, array_index_54713[0]} : sel_55036;
  assign add_55140 = array_index_54818[11:1] + 11'h347;
  assign sel_55142 = $signed({1'h0, add_55038, array_index_54716[0]}) < $signed({1'h0, sel_55040}) ? {add_55038, array_index_54716[0]} : sel_55040;
  assign add_55144 = array_index_54917[11:3] + 9'h0bd;
  assign sel_55147 = $signed({1'h0, add_55042, array_index_54815[2:0]}) < $signed({1'h0, sel_55045}) ? {add_55042, array_index_54815[2:0]} : sel_55045;
  assign add_55149 = array_index_54920[11:3] + 9'h0bd;
  assign sel_55152 = $signed({1'h0, add_55047, array_index_54818[2:0]}) < $signed({1'h0, sel_55050}) ? {add_55047, array_index_54818[2:0]} : sel_55050;
  assign add_55154 = array_index_55019[11:1] + 11'h247;
  assign sel_55157 = $signed({1'h0, add_55052, array_index_54917[0]}) < $signed({1'h0, sel_55055}) ? {add_55052, array_index_54917[0]} : sel_55055;
  assign add_55159 = array_index_55022[11:1] + 11'h247;
  assign sel_55162 = $signed({1'h0, add_55057, array_index_54920[0]}) < $signed({1'h0, sel_55060}) ? {add_55057, array_index_54920[0]} : sel_55060;
  assign add_55187 = array_index_55121[11:0] + 12'h247;
  assign sel_55189 = $signed({1'h0, add_55085}) < $signed({1'h0, sel_55087}) ? add_55085 : sel_55087;
  assign add_55192 = array_index_55124[11:0] + 12'h247;
  assign sel_55194 = $signed({1'h0, add_55090}) < $signed({1'h0, sel_55092}) ? add_55090 : sel_55092;
  assign array_index_55223 = set1_unflattened[5'h1c];
  assign array_index_55226 = set2_unflattened[5'h1c];
  assign add_55230 = array_index_54815[11:1] + 11'h79d;
  assign sel_55232 = $signed({1'h0, add_55128, array_index_54713[0]}) < $signed({1'h0, sel_55130}) ? {add_55128, array_index_54713[0]} : sel_55130;
  assign add_55234 = array_index_54818[11:1] + 11'h79d;
  assign sel_55236 = $signed({1'h0, add_55132, array_index_54716[0]}) < $signed({1'h0, sel_55134}) ? {add_55132, array_index_54716[0]} : sel_55134;
  assign add_55238 = array_index_54917[11:1] + 11'h347;
  assign sel_55240 = $signed({1'h0, add_55136, array_index_54815[0]}) < $signed({1'h0, sel_55138}) ? {add_55136, array_index_54815[0]} : sel_55138;
  assign add_55242 = array_index_54920[11:1] + 11'h347;
  assign sel_55244 = $signed({1'h0, add_55140, array_index_54818[0]}) < $signed({1'h0, sel_55142}) ? {add_55140, array_index_54818[0]} : sel_55142;
  assign add_55246 = array_index_55019[11:3] + 9'h0bd;
  assign sel_55249 = $signed({1'h0, add_55144, array_index_54917[2:0]}) < $signed({1'h0, sel_55147}) ? {add_55144, array_index_54917[2:0]} : sel_55147;
  assign add_55251 = array_index_55022[11:3] + 9'h0bd;
  assign sel_55254 = $signed({1'h0, add_55149, array_index_54920[2:0]}) < $signed({1'h0, sel_55152}) ? {add_55149, array_index_54920[2:0]} : sel_55152;
  assign add_55256 = array_index_55121[11:1] + 11'h247;
  assign sel_55259 = $signed({1'h0, add_55154, array_index_55019[0]}) < $signed({1'h0, sel_55157}) ? {add_55154, array_index_55019[0]} : sel_55157;
  assign add_55261 = array_index_55124[11:1] + 11'h247;
  assign sel_55264 = $signed({1'h0, add_55159, array_index_55022[0]}) < $signed({1'h0, sel_55162}) ? {add_55159, array_index_55022[0]} : sel_55162;
  assign add_55289 = array_index_55223[11:0] + 12'h247;
  assign sel_55291 = $signed({1'h0, add_55187}) < $signed({1'h0, sel_55189}) ? add_55187 : sel_55189;
  assign add_55294 = array_index_55226[11:0] + 12'h247;
  assign sel_55296 = $signed({1'h0, add_55192}) < $signed({1'h0, sel_55194}) ? add_55192 : sel_55194;
  assign array_index_55325 = set1_unflattened[5'h1d];
  assign array_index_55328 = set2_unflattened[5'h1d];
  assign add_55332 = array_index_54917[11:1] + 11'h79d;
  assign sel_55334 = $signed({1'h0, add_55230, array_index_54815[0]}) < $signed({1'h0, sel_55232}) ? {add_55230, array_index_54815[0]} : sel_55232;
  assign add_55336 = array_index_54920[11:1] + 11'h79d;
  assign sel_55338 = $signed({1'h0, add_55234, array_index_54818[0]}) < $signed({1'h0, sel_55236}) ? {add_55234, array_index_54818[0]} : sel_55236;
  assign add_55340 = array_index_55019[11:1] + 11'h347;
  assign sel_55342 = $signed({1'h0, add_55238, array_index_54917[0]}) < $signed({1'h0, sel_55240}) ? {add_55238, array_index_54917[0]} : sel_55240;
  assign add_55344 = array_index_55022[11:1] + 11'h347;
  assign sel_55346 = $signed({1'h0, add_55242, array_index_54920[0]}) < $signed({1'h0, sel_55244}) ? {add_55242, array_index_54920[0]} : sel_55244;
  assign add_55348 = array_index_55121[11:3] + 9'h0bd;
  assign sel_55351 = $signed({1'h0, add_55246, array_index_55019[2:0]}) < $signed({1'h0, sel_55249}) ? {add_55246, array_index_55019[2:0]} : sel_55249;
  assign add_55353 = array_index_55124[11:3] + 9'h0bd;
  assign sel_55356 = $signed({1'h0, add_55251, array_index_55022[2:0]}) < $signed({1'h0, sel_55254}) ? {add_55251, array_index_55022[2:0]} : sel_55254;
  assign add_55358 = array_index_55223[11:1] + 11'h247;
  assign sel_55361 = $signed({1'h0, add_55256, array_index_55121[0]}) < $signed({1'h0, sel_55259}) ? {add_55256, array_index_55121[0]} : sel_55259;
  assign add_55363 = array_index_55226[11:1] + 11'h247;
  assign sel_55366 = $signed({1'h0, add_55261, array_index_55124[0]}) < $signed({1'h0, sel_55264}) ? {add_55261, array_index_55124[0]} : sel_55264;
  assign add_55390 = array_index_55325[11:0] + 12'h247;
  assign sel_55392 = $signed({1'h0, add_55289}) < $signed({1'h0, sel_55291}) ? add_55289 : sel_55291;
  assign add_55394 = array_index_55328[11:0] + 12'h247;
  assign sel_55396 = $signed({1'h0, add_55294}) < $signed({1'h0, sel_55296}) ? add_55294 : sel_55296;
  assign add_55430 = array_index_55019[11:1] + 11'h79d;
  assign sel_55432 = $signed({1'h0, add_55332, array_index_54917[0]}) < $signed({1'h0, sel_55334}) ? {add_55332, array_index_54917[0]} : sel_55334;
  assign add_55434 = array_index_55022[11:1] + 11'h79d;
  assign sel_55436 = $signed({1'h0, add_55336, array_index_54920[0]}) < $signed({1'h0, sel_55338}) ? {add_55336, array_index_54920[0]} : sel_55338;
  assign add_55438 = array_index_55121[11:1] + 11'h347;
  assign sel_55440 = $signed({1'h0, add_55340, array_index_55019[0]}) < $signed({1'h0, sel_55342}) ? {add_55340, array_index_55019[0]} : sel_55342;
  assign add_55442 = array_index_55124[11:1] + 11'h347;
  assign sel_55444 = $signed({1'h0, add_55344, array_index_55022[0]}) < $signed({1'h0, sel_55346}) ? {add_55344, array_index_55022[0]} : sel_55346;
  assign add_55446 = array_index_55223[11:3] + 9'h0bd;
  assign sel_55449 = $signed({1'h0, add_55348, array_index_55121[2:0]}) < $signed({1'h0, sel_55351}) ? {add_55348, array_index_55121[2:0]} : sel_55351;
  assign add_55451 = array_index_55226[11:3] + 9'h0bd;
  assign sel_55454 = $signed({1'h0, add_55353, array_index_55124[2:0]}) < $signed({1'h0, sel_55356}) ? {add_55353, array_index_55124[2:0]} : sel_55356;
  assign add_55456 = array_index_55325[11:1] + 11'h247;
  assign sel_55459 = $signed({1'h0, add_55358, array_index_55223[0]}) < $signed({1'h0, sel_55361}) ? {add_55358, array_index_55223[0]} : sel_55361;
  assign add_55461 = array_index_55328[11:1] + 11'h247;
  assign sel_55464 = $signed({1'h0, add_55363, array_index_55226[0]}) < $signed({1'h0, sel_55366}) ? {add_55363, array_index_55226[0]} : sel_55366;
  assign add_55512 = array_index_55121[11:1] + 11'h79d;
  assign sel_55514 = $signed({1'h0, add_55430, array_index_55019[0]}) < $signed({1'h0, sel_55432}) ? {add_55430, array_index_55019[0]} : sel_55432;
  assign add_55516 = array_index_55124[11:1] + 11'h79d;
  assign sel_55518 = $signed({1'h0, add_55434, array_index_55022[0]}) < $signed({1'h0, sel_55436}) ? {add_55434, array_index_55022[0]} : sel_55436;
  assign add_55520 = array_index_55223[11:1] + 11'h347;
  assign sel_55522 = $signed({1'h0, add_55438, array_index_55121[0]}) < $signed({1'h0, sel_55440}) ? {add_55438, array_index_55121[0]} : sel_55440;
  assign add_55524 = array_index_55226[11:1] + 11'h347;
  assign sel_55526 = $signed({1'h0, add_55442, array_index_55124[0]}) < $signed({1'h0, sel_55444}) ? {add_55442, array_index_55124[0]} : sel_55444;
  assign add_55528 = array_index_55325[11:3] + 9'h0bd;
  assign sel_55531 = $signed({1'h0, add_55446, array_index_55223[2:0]}) < $signed({1'h0, sel_55449}) ? {add_55446, array_index_55223[2:0]} : sel_55449;
  assign add_55533 = array_index_55328[11:3] + 9'h0bd;
  assign sel_55536 = $signed({1'h0, add_55451, array_index_55226[2:0]}) < $signed({1'h0, sel_55454}) ? {add_55451, array_index_55226[2:0]} : sel_55454;
  assign concat_55539 = {1'h0, ($signed({1'h0, add_55390}) < $signed({1'h0, sel_55392}) ? add_55390 : sel_55392) == ($signed({1'h0, add_55394}) < $signed({1'h0, sel_55396}) ? add_55394 : sel_55396)};
  assign add_55554 = concat_55539 + 2'h1;
  assign add_55574 = array_index_55223[11:1] + 11'h79d;
  assign sel_55576 = $signed({1'h0, add_55512, array_index_55121[0]}) < $signed({1'h0, sel_55514}) ? {add_55512, array_index_55121[0]} : sel_55514;
  assign add_55578 = array_index_55226[11:1] + 11'h79d;
  assign sel_55580 = $signed({1'h0, add_55516, array_index_55124[0]}) < $signed({1'h0, sel_55518}) ? {add_55516, array_index_55124[0]} : sel_55518;
  assign add_55582 = array_index_55325[11:1] + 11'h347;
  assign sel_55584 = $signed({1'h0, add_55520, array_index_55223[0]}) < $signed({1'h0, sel_55522}) ? {add_55520, array_index_55223[0]} : sel_55522;
  assign add_55586 = array_index_55328[11:1] + 11'h347;
  assign sel_55588 = $signed({1'h0, add_55524, array_index_55226[0]}) < $signed({1'h0, sel_55526}) ? {add_55524, array_index_55226[0]} : sel_55526;
  assign concat_55591 = {1'h0, ($signed({1'h0, add_55456, array_index_55325[0]}) < $signed({1'h0, sel_55459}) ? {add_55456, array_index_55325[0]} : sel_55459) == ($signed({1'h0, add_55461, array_index_55328[0]}) < $signed({1'h0, sel_55464}) ? {add_55461, array_index_55328[0]} : sel_55464) ? add_55554 : concat_55539};
  assign add_55602 = concat_55591 + 3'h1;
  assign add_55616 = array_index_55325[11:1] + 11'h79d;
  assign sel_55618 = $signed({1'h0, add_55574, array_index_55223[0]}) < $signed({1'h0, sel_55576}) ? {add_55574, array_index_55223[0]} : sel_55576;
  assign add_55620 = array_index_55328[11:1] + 11'h79d;
  assign sel_55622 = $signed({1'h0, add_55578, array_index_55226[0]}) < $signed({1'h0, sel_55580}) ? {add_55578, array_index_55226[0]} : sel_55580;
  assign concat_55625 = {1'h0, ($signed({1'h0, add_55528, array_index_55325[2:0]}) < $signed({1'h0, sel_55531}) ? {add_55528, array_index_55325[2:0]} : sel_55531) == ($signed({1'h0, add_55533, array_index_55328[2:0]}) < $signed({1'h0, sel_55536}) ? {add_55533, array_index_55328[2:0]} : sel_55536) ? add_55602 : concat_55591};
  assign add_55632 = concat_55625 + 4'h1;
  assign concat_55641 = {1'h0, ($signed({1'h0, add_55582, array_index_55325[0]}) < $signed({1'h0, sel_55584}) ? {add_55582, array_index_55325[0]} : sel_55584) == ($signed({1'h0, add_55586, array_index_55328[0]}) < $signed({1'h0, sel_55588}) ? {add_55586, array_index_55328[0]} : sel_55588) ? add_55632 : concat_55625};
  assign add_55644 = concat_55641 + 5'h01;
  assign out = {{11'h000, ($signed({1'h0, add_55616, array_index_55325[0]}) < $signed({1'h0, sel_55618}) ? {add_55616, array_index_55325[0]} : sel_55618) == ($signed({1'h0, add_55620, array_index_55328[0]}) < $signed({1'h0, sel_55622}) ? {add_55620, array_index_55328[0]} : sel_55622) ? add_55644 : concat_55641}, {set1_unflattened[29], set1_unflattened[28], set1_unflattened[27], set1_unflattened[26], set1_unflattened[25], set1_unflattened[24], set1_unflattened[23], set1_unflattened[22], set1_unflattened[21], set1_unflattened[20], set1_unflattened[19], set1_unflattened[18], set1_unflattened[17], set1_unflattened[16], set1_unflattened[15], set1_unflattened[14], set1_unflattened[13], set1_unflattened[12], set1_unflattened[11], set1_unflattened[10], set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[29], set2_unflattened[28], set2_unflattened[27], set2_unflattened[26], set2_unflattened[25], set2_unflattened[24], set2_unflattened[23], set2_unflattened[22], set2_unflattened[21], set2_unflattened[20], set2_unflattened[19], set2_unflattened[18], set2_unflattened[17], set2_unflattened[16], set2_unflattened[15], set2_unflattened[14], set2_unflattened[13], set2_unflattened[12], set2_unflattened[11], set2_unflattened[10], set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
