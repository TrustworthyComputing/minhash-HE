module min_hash(
  input wire [159:0] set1,
  input wire [159:0] set2,
  output wire [335:0] out
);
  // lint_off MULTIPLY
  function automatic [21:0] umul22b_16b_x_6b (input reg [15:0] lhs, input reg [5:0] rhs);
    begin
      umul22b_16b_x_6b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  // lint_off MULTIPLY
  function automatic [22:0] umul23b_16b_x_7b (input reg [15:0] lhs, input reg [6:0] rhs);
    begin
      umul23b_16b_x_7b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [15:0] set1_unflattened[10];
  assign set1_unflattened[0] = set1[15:0];
  assign set1_unflattened[1] = set1[31:16];
  assign set1_unflattened[2] = set1[47:32];
  assign set1_unflattened[3] = set1[63:48];
  assign set1_unflattened[4] = set1[79:64];
  assign set1_unflattened[5] = set1[95:80];
  assign set1_unflattened[6] = set1[111:96];
  assign set1_unflattened[7] = set1[127:112];
  assign set1_unflattened[8] = set1[143:128];
  assign set1_unflattened[9] = set1[159:144];
  wire [15:0] set2_unflattened[10];
  assign set2_unflattened[0] = set2[15:0];
  assign set2_unflattened[1] = set2[31:16];
  assign set2_unflattened[2] = set2[47:32];
  assign set2_unflattened[3] = set2[63:48];
  assign set2_unflattened[4] = set2[79:64];
  assign set2_unflattened[5] = set2[95:80];
  assign set2_unflattened[6] = set2[111:96];
  assign set2_unflattened[7] = set2[127:112];
  assign set2_unflattened[8] = set2[143:128];
  assign set2_unflattened[9] = set2[159:144];
  wire [15:0] array_index_18114;
  wire [15:0] array_index_18116;
  wire [21:0] umul_18118;
  wire [21:0] umul_18119;
  wire [21:0] umul_18128;
  wire [21:0] umul_18129;
  wire [15:0] array_index_18130;
  wire [15:0] array_index_18134;
  wire [21:0] umul_18142;
  wire [15:0] add_18144;
  wire [21:0] umul_18146;
  wire [15:0] add_18148;
  wire [21:0] umul_18168;
  wire [21:0] umul_18169;
  wire [21:0] umul_18170;
  wire [21:0] add_18172;
  wire [21:0] umul_18174;
  wire [21:0] add_18176;
  wire [15:0] array_index_18178;
  wire [31:0] smod_18182;
  wire [15:0] array_index_18183;
  wire [31:0] smod_18187;
  wire [21:0] umul_18200;
  wire [15:0] add_18202;
  wire [21:0] umul_18206;
  wire [15:0] add_18208;
  wire [31:0] smod_18223;
  wire [31:0] smod_18227;
  wire [22:0] umul_18242;
  wire [22:0] umul_18243;
  wire [21:0] umul_18244;
  wire [20:0] add_18246;
  wire [21:0] umul_18248;
  wire [20:0] add_18250;
  wire [21:0] umul_18252;
  wire [21:0] add_18254;
  wire [21:0] umul_18258;
  wire [21:0] add_18260;
  wire [15:0] array_index_18264;
  wire [31:0] smod_18268;
  wire [15:0] array_index_18271;
  wire [31:0] smod_18275;
  wire [21:0] umul_18302;
  wire [15:0] add_18304;
  wire [15:0] sel_18309;
  wire [21:0] umul_18310;
  wire [15:0] add_18312;
  wire [15:0] sel_18317;
  wire [31:0] smod_18329;
  wire [31:0] smod_18333;
  wire [31:0] smod_18337;
  wire [31:0] smod_18343;
  wire [22:0] umul_18360;
  wire [22:0] umul_18361;
  wire [22:0] umul_18362;
  wire [22:0] add_18364;
  wire [22:0] umul_18366;
  wire [22:0] add_18368;
  wire [21:0] umul_18370;
  wire [20:0] add_18372;
  wire [21:0] umul_18376;
  wire [20:0] add_18378;
  wire [21:0] umul_18382;
  wire [21:0] add_18384;
  wire [15:0] sel_18389;
  wire [21:0] umul_18390;
  wire [21:0] add_18392;
  wire [15:0] sel_18397;
  wire [15:0] array_index_18398;
  wire [31:0] smod_18402;
  wire [15:0] array_index_18404;
  wire [31:0] smod_18408;
  wire [21:0] umul_18446;
  wire [15:0] add_18448;
  wire [15:0] sel_18453;
  wire [21:0] umul_18454;
  wire [15:0] add_18456;
  wire [15:0] sel_18461;
  wire [31:0] smod_18471;
  wire [31:0] smod_18475;
  wire [31:0] smod_18479;
  wire [31:0] smod_18485;
  wire [31:0] smod_18491;
  wire [31:0] smod_18496;
  wire [22:0] umul_18512;
  wire [20:0] add_18514;
  wire [22:0] umul_18516;
  wire [20:0] add_18518;
  wire [22:0] umul_18520;
  wire [22:0] add_18522;
  wire [22:0] umul_18526;
  wire [22:0] add_18528;
  wire [21:0] umul_18532;
  wire [20:0] add_18534;
  wire [15:0] sel_18539;
  wire [21:0] umul_18540;
  wire [20:0] add_18542;
  wire [15:0] sel_18547;
  wire [21:0] umul_18548;
  wire [21:0] add_18550;
  wire [15:0] sel_18555;
  wire [21:0] umul_18556;
  wire [21:0] add_18558;
  wire [15:0] sel_18563;
  wire [15:0] array_index_18564;
  wire [31:0] smod_18568;
  wire [15:0] array_index_18570;
  wire [31:0] smod_18574;
  wire [21:0] umul_18620;
  wire [15:0] add_18622;
  wire [15:0] sel_18627;
  wire [21:0] umul_18628;
  wire [15:0] add_18630;
  wire [15:0] sel_18635;
  wire [31:0] smod_18639;
  wire [31:0] smod_18643;
  wire [31:0] smod_18647;
  wire [31:0] smod_18653;
  wire [31:0] smod_18659;
  wire [31:0] smod_18664;
  wire [31:0] smod_18669;
  wire [31:0] smod_18674;
  wire [22:0] umul_18690;
  wire [20:0] add_18692;
  wire [22:0] umul_18696;
  wire [20:0] add_18698;
  wire [22:0] umul_18702;
  wire [22:0] add_18704;
  wire [15:0] sel_18709;
  wire [22:0] umul_18710;
  wire [22:0] add_18712;
  wire [15:0] sel_18717;
  wire [21:0] umul_18718;
  wire [20:0] add_18720;
  wire [15:0] sel_18725;
  wire [21:0] umul_18726;
  wire [20:0] add_18728;
  wire [15:0] sel_18733;
  wire [21:0] umul_18734;
  wire [21:0] add_18736;
  wire [15:0] sel_18741;
  wire [21:0] umul_18742;
  wire [21:0] add_18744;
  wire [15:0] sel_18749;
  wire [15:0] array_index_18750;
  wire [31:0] smod_18754;
  wire [15:0] array_index_18756;
  wire [31:0] smod_18760;
  wire [21:0] umul_18810;
  wire [15:0] add_18812;
  wire [15:0] sel_18817;
  wire [21:0] umul_18818;
  wire [15:0] add_18820;
  wire [15:0] sel_18825;
  wire [31:0] smod_18829;
  wire [31:0] smod_18835;
  wire [31:0] smod_18841;
  wire [31:0] smod_18846;
  wire [31:0] smod_18851;
  wire [31:0] smod_18856;
  wire [31:0] smod_18861;
  wire [31:0] smod_18866;
  wire [22:0] umul_18882;
  wire [20:0] add_18884;
  wire [15:0] sel_18889;
  wire [22:0] umul_18890;
  wire [20:0] add_18892;
  wire [15:0] sel_18897;
  wire [22:0] umul_18898;
  wire [22:0] add_18900;
  wire [15:0] sel_18905;
  wire [22:0] umul_18906;
  wire [22:0] add_18908;
  wire [15:0] sel_18913;
  wire [21:0] umul_18914;
  wire [20:0] add_18916;
  wire [15:0] sel_18921;
  wire [21:0] umul_18922;
  wire [20:0] add_18924;
  wire [15:0] sel_18929;
  wire [21:0] umul_18930;
  wire [21:0] add_18932;
  wire [15:0] sel_18937;
  wire [21:0] umul_18938;
  wire [21:0] add_18940;
  wire [15:0] sel_18945;
  wire [15:0] array_index_18946;
  wire [31:0] smod_18950;
  wire [15:0] array_index_18952;
  wire [31:0] smod_18956;
  wire [21:0] umul_19006;
  wire [15:0] add_19008;
  wire [15:0] sel_19013;
  wire [21:0] umul_19014;
  wire [15:0] add_19016;
  wire [15:0] sel_19021;
  wire [31:0] smod_19025;
  wire [31:0] smod_19030;
  wire [31:0] smod_19035;
  wire [31:0] smod_19040;
  wire [31:0] smod_19045;
  wire [31:0] smod_19050;
  wire [31:0] smod_19055;
  wire [31:0] smod_19060;
  wire [22:0] umul_19076;
  wire [20:0] add_19078;
  wire [15:0] sel_19083;
  wire [22:0] umul_19084;
  wire [20:0] add_19086;
  wire [15:0] sel_19091;
  wire [22:0] umul_19092;
  wire [22:0] add_19094;
  wire [15:0] sel_19099;
  wire [22:0] umul_19100;
  wire [22:0] add_19102;
  wire [15:0] sel_19107;
  wire [21:0] umul_19108;
  wire [20:0] add_19110;
  wire [15:0] sel_19115;
  wire [21:0] umul_19116;
  wire [20:0] add_19118;
  wire [15:0] sel_19123;
  wire [21:0] umul_19124;
  wire [21:0] add_19126;
  wire [15:0] sel_19131;
  wire [21:0] umul_19132;
  wire [21:0] add_19134;
  wire [15:0] sel_19139;
  wire [15:0] array_index_19140;
  wire [31:0] smod_19144;
  wire [15:0] array_index_19146;
  wire [31:0] smod_19150;
  wire [21:0] umul_19200;
  wire [15:0] add_19202;
  wire [15:0] sel_19207;
  wire [21:0] umul_19208;
  wire [15:0] add_19210;
  wire [15:0] sel_19215;
  wire [31:0] smod_19219;
  wire [31:0] smod_19224;
  wire [31:0] smod_19229;
  wire [31:0] smod_19234;
  wire [31:0] smod_19239;
  wire [31:0] smod_19244;
  wire [31:0] smod_19249;
  wire [31:0] smod_19254;
  wire [22:0] umul_19270;
  wire [20:0] add_19272;
  wire [15:0] sel_19277;
  wire [22:0] umul_19278;
  wire [20:0] add_19280;
  wire [15:0] sel_19285;
  wire [22:0] umul_19286;
  wire [22:0] add_19288;
  wire [15:0] sel_19293;
  wire [22:0] umul_19294;
  wire [22:0] add_19296;
  wire [15:0] sel_19301;
  wire [21:0] umul_19302;
  wire [20:0] add_19304;
  wire [15:0] sel_19309;
  wire [21:0] umul_19310;
  wire [20:0] add_19312;
  wire [15:0] sel_19317;
  wire [21:0] umul_19318;
  wire [21:0] add_19320;
  wire [15:0] sel_19325;
  wire [21:0] umul_19326;
  wire [21:0] add_19328;
  wire [15:0] sel_19333;
  wire [15:0] array_index_19334;
  wire [31:0] smod_19338;
  wire [15:0] array_index_19340;
  wire [31:0] smod_19344;
  wire [21:0] umul_19394;
  wire [15:0] add_19396;
  wire [15:0] sel_19401;
  wire [21:0] umul_19402;
  wire [15:0] add_19404;
  wire [15:0] sel_19409;
  wire [31:0] smod_19413;
  wire [31:0] smod_19418;
  wire [31:0] smod_19423;
  wire [31:0] smod_19428;
  wire [31:0] smod_19433;
  wire [31:0] smod_19438;
  wire [31:0] smod_19443;
  wire [31:0] smod_19448;
  wire [22:0] umul_19462;
  wire [20:0] add_19464;
  wire [15:0] sel_19469;
  wire [22:0] umul_19470;
  wire [20:0] add_19472;
  wire [15:0] sel_19477;
  wire [22:0] umul_19478;
  wire [22:0] add_19480;
  wire [15:0] sel_19485;
  wire [22:0] umul_19486;
  wire [22:0] add_19488;
  wire [15:0] sel_19493;
  wire [21:0] umul_19494;
  wire [20:0] add_19496;
  wire [15:0] sel_19501;
  wire [21:0] umul_19502;
  wire [20:0] add_19504;
  wire [15:0] sel_19509;
  wire [21:0] umul_19510;
  wire [21:0] add_19512;
  wire [15:0] sel_19517;
  wire [21:0] umul_19518;
  wire [21:0] add_19520;
  wire [15:0] sel_19525;
  wire [31:0] smod_19528;
  wire [31:0] smod_19532;
  wire [15:0] add_19583;
  wire [15:0] sel_19588;
  wire [15:0] add_19590;
  wire [15:0] sel_19595;
  wire [31:0] smod_19599;
  wire [31:0] smod_19604;
  wire [31:0] smod_19609;
  wire [31:0] smod_19614;
  wire [31:0] smod_19619;
  wire [31:0] smod_19624;
  wire [31:0] smod_19628;
  wire [31:0] smod_19632;
  wire [22:0] umul_19642;
  wire [20:0] add_19644;
  wire [15:0] sel_19649;
  wire [22:0] umul_19650;
  wire [20:0] add_19652;
  wire [15:0] sel_19657;
  wire [22:0] umul_19658;
  wire [22:0] add_19660;
  wire [15:0] sel_19665;
  wire [22:0] umul_19666;
  wire [22:0] add_19668;
  wire [15:0] sel_19673;
  wire [21:0] umul_19674;
  wire [20:0] add_19676;
  wire [15:0] sel_19681;
  wire [21:0] umul_19682;
  wire [20:0] add_19684;
  wire [15:0] sel_19689;
  wire [21:0] add_19691;
  wire [15:0] sel_19696;
  wire [21:0] add_19698;
  wire [15:0] sel_19703;
  wire [31:0] smod_19704;
  wire [31:0] smod_19706;
  wire [15:0] sel_19755;
  wire [15:0] sel_19759;
  wire [31:0] smod_19763;
  wire [31:0] smod_19768;
  wire [31:0] smod_19773;
  wire [31:0] smod_19778;
  wire [31:0] smod_19782;
  wire [31:0] smod_19786;
  wire [31:0] smod_19788;
  wire [31:0] smod_19790;
  wire [22:0] umul_19796;
  wire [20:0] add_19798;
  wire [15:0] sel_19803;
  wire [22:0] umul_19804;
  wire [20:0] add_19806;
  wire [15:0] sel_19811;
  wire [22:0] umul_19812;
  wire [22:0] add_19814;
  wire [15:0] sel_19819;
  wire [22:0] umul_19820;
  wire [22:0] add_19822;
  wire [15:0] sel_19827;
  wire [20:0] add_19829;
  wire [15:0] sel_19834;
  wire [20:0] add_19836;
  wire [15:0] sel_19841;
  wire [15:0] sel_19845;
  wire [15:0] sel_19849;
  wire [31:0] smod_19893;
  wire [31:0] smod_19898;
  wire [31:0] smod_19902;
  wire [31:0] smod_19906;
  wire [31:0] smod_19908;
  wire [31:0] smod_19910;
  wire [22:0] umul_19916;
  wire [20:0] add_19918;
  wire [15:0] sel_19923;
  wire [22:0] umul_19924;
  wire [20:0] add_19926;
  wire [15:0] sel_19931;
  wire [22:0] add_19933;
  wire [15:0] sel_19938;
  wire [22:0] add_19940;
  wire [15:0] sel_19945;
  wire [15:0] sel_19949;
  wire [15:0] sel_19953;
  wire [1:0] concat_19956;
  wire [1:0] add_19983;
  wire [31:0] smod_19986;
  wire [31:0] smod_19990;
  wire [31:0] smod_19992;
  wire [31:0] smod_19994;
  wire [20:0] add_20001;
  wire [15:0] sel_20006;
  wire [20:0] add_20008;
  wire [15:0] sel_20013;
  wire [15:0] sel_20017;
  wire [15:0] sel_20021;
  wire [2:0] concat_20024;
  wire [2:0] add_20039;
  wire [31:0] smod_20040;
  wire [31:0] smod_20042;
  wire [15:0] sel_20051;
  wire [15:0] sel_20055;
  wire [3:0] concat_20058;
  wire [3:0] add_20065;
  wire [4:0] concat_20072;
  wire [4:0] add_20075;
  assign array_index_18114 = set1_unflattened[4'h0];
  assign array_index_18116 = set2_unflattened[4'h0];
  assign umul_18118 = umul22b_16b_x_6b(array_index_18114, 6'h35);
  assign umul_18119 = umul22b_16b_x_6b(array_index_18116, 6'h35);
  assign umul_18128 = umul22b_16b_x_6b(array_index_18114, 6'h3b);
  assign umul_18129 = umul22b_16b_x_6b(array_index_18116, 6'h3b);
  assign array_index_18130 = set1_unflattened[4'h1];
  assign array_index_18134 = set2_unflattened[4'h1];
  assign umul_18142 = umul22b_16b_x_6b(array_index_18130, 6'h35);
  assign add_18144 = {1'h0, umul_18118[21:7]} + 16'h007d;
  assign umul_18146 = umul22b_16b_x_6b(array_index_18134, 6'h35);
  assign add_18148 = {1'h0, umul_18119[21:7]} + 16'h007d;
  assign umul_18168 = umul22b_16b_x_6b(array_index_18114, 6'h3d);
  assign umul_18169 = umul22b_16b_x_6b(array_index_18116, 6'h3d);
  assign umul_18170 = umul22b_16b_x_6b(array_index_18130, 6'h3b);
  assign add_18172 = {1'h0, umul_18128[21:1]} + 22'h00_1f59;
  assign umul_18174 = umul22b_16b_x_6b(array_index_18134, 6'h3b);
  assign add_18176 = {1'h0, umul_18129[21:1]} + 22'h00_1f59;
  assign array_index_18178 = set1_unflattened[4'h2];
  assign smod_18182 = $unsigned($signed({9'h000, add_18144, umul_18118[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_18183 = set2_unflattened[4'h2];
  assign smod_18187 = $unsigned($signed({9'h000, add_18148, umul_18119[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_18200 = umul22b_16b_x_6b(array_index_18178, 6'h35);
  assign add_18202 = {1'h0, umul_18142[21:7]} + 16'h007d;
  assign umul_18206 = umul22b_16b_x_6b(array_index_18183, 6'h35);
  assign add_18208 = {1'h0, umul_18146[21:7]} + 16'h007d;
  assign smod_18223 = $unsigned($signed({9'h000, add_18172, umul_18128[0]}) % $signed(32'h0000_3ffd));
  assign smod_18227 = $unsigned($signed({9'h000, add_18176, umul_18129[0]}) % $signed(32'h0000_3ffd));
  assign umul_18242 = umul23b_16b_x_7b(array_index_18114, 7'h47);
  assign umul_18243 = umul23b_16b_x_7b(array_index_18116, 7'h47);
  assign umul_18244 = umul22b_16b_x_6b(array_index_18130, 6'h3d);
  assign add_18246 = {1'h0, umul_18168[21:2]} + 21'h00_0fb9;
  assign umul_18248 = umul22b_16b_x_6b(array_index_18134, 6'h3d);
  assign add_18250 = {1'h0, umul_18169[21:2]} + 21'h00_0fb9;
  assign umul_18252 = umul22b_16b_x_6b(array_index_18178, 6'h3b);
  assign add_18254 = {1'h0, umul_18170[21:1]} + 22'h00_1f59;
  assign umul_18258 = umul22b_16b_x_6b(array_index_18183, 6'h3b);
  assign add_18260 = {1'h0, umul_18174[21:1]} + 22'h00_1f59;
  assign array_index_18264 = set1_unflattened[4'h3];
  assign smod_18268 = $unsigned($signed({9'h000, add_18202, umul_18142[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_18271 = set2_unflattened[4'h3];
  assign smod_18275 = $unsigned($signed({9'h000, add_18208, umul_18146[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_18302 = umul22b_16b_x_6b(array_index_18264, 6'h35);
  assign add_18304 = {1'h0, umul_18200[21:7]} + 16'h007d;
  assign sel_18309 = $signed({1'h0, smod_18182[15:0]}) < $signed(17'h0_3ffd) ? smod_18182[15:0] : 16'h3ffd;
  assign umul_18310 = umul22b_16b_x_6b(array_index_18271, 6'h35);
  assign add_18312 = {1'h0, umul_18206[21:7]} + 16'h007d;
  assign sel_18317 = $signed({1'h0, smod_18187[15:0]}) < $signed(17'h0_3ffd) ? smod_18187[15:0] : 16'h3ffd;
  assign smod_18329 = $unsigned($signed({9'h000, add_18246, umul_18168[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_18333 = $unsigned($signed({9'h000, add_18250, umul_18169[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_18337 = $unsigned($signed({9'h000, add_18254, umul_18170[0]}) % $signed(32'h0000_3ffd));
  assign smod_18343 = $unsigned($signed({9'h000, add_18260, umul_18174[0]}) % $signed(32'h0000_3ffd));
  assign umul_18360 = umul23b_16b_x_7b(array_index_18114, 7'h49);
  assign umul_18361 = umul23b_16b_x_7b(array_index_18116, 7'h49);
  assign umul_18362 = umul23b_16b_x_7b(array_index_18130, 7'h47);
  assign add_18364 = {1'h0, umul_18242[22:1]} + 23'h00_1f8b;
  assign umul_18366 = umul23b_16b_x_7b(array_index_18134, 7'h47);
  assign add_18368 = {1'h0, umul_18243[22:1]} + 23'h00_1f8b;
  assign umul_18370 = umul22b_16b_x_6b(array_index_18178, 6'h3d);
  assign add_18372 = {1'h0, umul_18244[21:2]} + 21'h00_0fb9;
  assign umul_18376 = umul22b_16b_x_6b(array_index_18183, 6'h3d);
  assign add_18378 = {1'h0, umul_18248[21:2]} + 21'h00_0fb9;
  assign umul_18382 = umul22b_16b_x_6b(array_index_18264, 6'h3b);
  assign add_18384 = {1'h0, umul_18252[21:1]} + 22'h00_1f59;
  assign sel_18389 = $signed({1'h0, smod_18223[15:0]}) < $signed(17'h0_3ffd) ? smod_18223[15:0] : 16'h3ffd;
  assign umul_18390 = umul22b_16b_x_6b(array_index_18271, 6'h3b);
  assign add_18392 = {1'h0, umul_18258[21:1]} + 22'h00_1f59;
  assign sel_18397 = $signed({1'h0, smod_18227[15:0]}) < $signed(17'h0_3ffd) ? smod_18227[15:0] : 16'h3ffd;
  assign array_index_18398 = set1_unflattened[4'h4];
  assign smod_18402 = $unsigned($signed({9'h000, add_18304, umul_18200[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_18404 = set2_unflattened[4'h4];
  assign smod_18408 = $unsigned($signed({9'h000, add_18312, umul_18206[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_18446 = umul22b_16b_x_6b(array_index_18398, 6'h35);
  assign add_18448 = {1'h0, umul_18302[21:7]} + 16'h007d;
  assign sel_18453 = $signed({1'h0, smod_18268[15:0]}) < $signed({1'h0, sel_18309}) ? smod_18268[15:0] : sel_18309;
  assign umul_18454 = umul22b_16b_x_6b(array_index_18404, 6'h35);
  assign add_18456 = {1'h0, umul_18310[21:7]} + 16'h007d;
  assign sel_18461 = $signed({1'h0, smod_18275[15:0]}) < $signed({1'h0, sel_18317}) ? smod_18275[15:0] : sel_18317;
  assign smod_18471 = $unsigned($signed({8'h00, add_18364, umul_18242[0]}) % $signed(32'h0000_3ffd));
  assign smod_18475 = $unsigned($signed({8'h00, add_18368, umul_18243[0]}) % $signed(32'h0000_3ffd));
  assign smod_18479 = $unsigned($signed({9'h000, add_18372, umul_18244[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_18485 = $unsigned($signed({9'h000, add_18378, umul_18248[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_18491 = $unsigned($signed({9'h000, add_18384, umul_18252[0]}) % $signed(32'h0000_3ffd));
  assign smod_18496 = $unsigned($signed({9'h000, add_18392, umul_18258[0]}) % $signed(32'h0000_3ffd));
  assign umul_18512 = umul23b_16b_x_7b(array_index_18130, 7'h49);
  assign add_18514 = {1'h0, umul_18360[22:3]} + 21'h00_07e9;
  assign umul_18516 = umul23b_16b_x_7b(array_index_18134, 7'h49);
  assign add_18518 = {1'h0, umul_18361[22:3]} + 21'h00_07e9;
  assign umul_18520 = umul23b_16b_x_7b(array_index_18178, 7'h47);
  assign add_18522 = {1'h0, umul_18362[22:1]} + 23'h00_1f8b;
  assign umul_18526 = umul23b_16b_x_7b(array_index_18183, 7'h47);
  assign add_18528 = {1'h0, umul_18366[22:1]} + 23'h00_1f8b;
  assign umul_18532 = umul22b_16b_x_6b(array_index_18264, 6'h3d);
  assign add_18534 = {1'h0, umul_18370[21:2]} + 21'h00_0fb9;
  assign sel_18539 = $signed({1'h0, smod_18329[15:0]}) < $signed(17'h0_3ffd) ? smod_18329[15:0] : 16'h3ffd;
  assign umul_18540 = umul22b_16b_x_6b(array_index_18271, 6'h3d);
  assign add_18542 = {1'h0, umul_18376[21:2]} + 21'h00_0fb9;
  assign sel_18547 = $signed({1'h0, smod_18333[15:0]}) < $signed(17'h0_3ffd) ? smod_18333[15:0] : 16'h3ffd;
  assign umul_18548 = umul22b_16b_x_6b(array_index_18398, 6'h3b);
  assign add_18550 = {1'h0, umul_18382[21:1]} + 22'h00_1f59;
  assign sel_18555 = $signed({1'h0, smod_18337[15:0]}) < $signed({1'h0, sel_18389}) ? smod_18337[15:0] : sel_18389;
  assign umul_18556 = umul22b_16b_x_6b(array_index_18404, 6'h3b);
  assign add_18558 = {1'h0, umul_18390[21:1]} + 22'h00_1f59;
  assign sel_18563 = $signed({1'h0, smod_18343[15:0]}) < $signed({1'h0, sel_18397}) ? smod_18343[15:0] : sel_18397;
  assign array_index_18564 = set1_unflattened[4'h5];
  assign smod_18568 = $unsigned($signed({9'h000, add_18448, umul_18302[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_18570 = set2_unflattened[4'h5];
  assign smod_18574 = $unsigned($signed({9'h000, add_18456, umul_18310[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_18620 = umul22b_16b_x_6b(array_index_18564, 6'h35);
  assign add_18622 = {1'h0, umul_18446[21:7]} + 16'h007d;
  assign sel_18627 = $signed({1'h0, smod_18402[15:0]}) < $signed({1'h0, sel_18453}) ? smod_18402[15:0] : sel_18453;
  assign umul_18628 = umul22b_16b_x_6b(array_index_18570, 6'h35);
  assign add_18630 = {1'h0, umul_18454[21:7]} + 16'h007d;
  assign sel_18635 = $signed({1'h0, smod_18408[15:0]}) < $signed({1'h0, sel_18461}) ? smod_18408[15:0] : sel_18461;
  assign smod_18639 = $unsigned($signed({8'h00, add_18514, umul_18360[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_18643 = $unsigned($signed({8'h00, add_18518, umul_18361[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_18647 = $unsigned($signed({8'h00, add_18522, umul_18362[0]}) % $signed(32'h0000_3ffd));
  assign smod_18653 = $unsigned($signed({8'h00, add_18528, umul_18366[0]}) % $signed(32'h0000_3ffd));
  assign smod_18659 = $unsigned($signed({9'h000, add_18534, umul_18370[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_18664 = $unsigned($signed({9'h000, add_18542, umul_18376[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_18669 = $unsigned($signed({9'h000, add_18550, umul_18382[0]}) % $signed(32'h0000_3ffd));
  assign smod_18674 = $unsigned($signed({9'h000, add_18558, umul_18390[0]}) % $signed(32'h0000_3ffd));
  assign umul_18690 = umul23b_16b_x_7b(array_index_18178, 7'h49);
  assign add_18692 = {1'h0, umul_18512[22:3]} + 21'h00_07e9;
  assign umul_18696 = umul23b_16b_x_7b(array_index_18183, 7'h49);
  assign add_18698 = {1'h0, umul_18516[22:3]} + 21'h00_07e9;
  assign umul_18702 = umul23b_16b_x_7b(array_index_18264, 7'h47);
  assign add_18704 = {1'h0, umul_18520[22:1]} + 23'h00_1f8b;
  assign sel_18709 = $signed({1'h0, smod_18471[15:0]}) < $signed(17'h0_3ffd) ? smod_18471[15:0] : 16'h3ffd;
  assign umul_18710 = umul23b_16b_x_7b(array_index_18271, 7'h47);
  assign add_18712 = {1'h0, umul_18526[22:1]} + 23'h00_1f8b;
  assign sel_18717 = $signed({1'h0, smod_18475[15:0]}) < $signed(17'h0_3ffd) ? smod_18475[15:0] : 16'h3ffd;
  assign umul_18718 = umul22b_16b_x_6b(array_index_18398, 6'h3d);
  assign add_18720 = {1'h0, umul_18532[21:2]} + 21'h00_0fb9;
  assign sel_18725 = $signed({1'h0, smod_18479[15:0]}) < $signed({1'h0, sel_18539}) ? smod_18479[15:0] : sel_18539;
  assign umul_18726 = umul22b_16b_x_6b(array_index_18404, 6'h3d);
  assign add_18728 = {1'h0, umul_18540[21:2]} + 21'h00_0fb9;
  assign sel_18733 = $signed({1'h0, smod_18485[15:0]}) < $signed({1'h0, sel_18547}) ? smod_18485[15:0] : sel_18547;
  assign umul_18734 = umul22b_16b_x_6b(array_index_18564, 6'h3b);
  assign add_18736 = {1'h0, umul_18548[21:1]} + 22'h00_1f59;
  assign sel_18741 = $signed({1'h0, smod_18491[15:0]}) < $signed({1'h0, sel_18555}) ? smod_18491[15:0] : sel_18555;
  assign umul_18742 = umul22b_16b_x_6b(array_index_18570, 6'h3b);
  assign add_18744 = {1'h0, umul_18556[21:1]} + 22'h00_1f59;
  assign sel_18749 = $signed({1'h0, smod_18496[15:0]}) < $signed({1'h0, sel_18563}) ? smod_18496[15:0] : sel_18563;
  assign array_index_18750 = set1_unflattened[4'h6];
  assign smod_18754 = $unsigned($signed({9'h000, add_18622, umul_18446[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_18756 = set2_unflattened[4'h6];
  assign smod_18760 = $unsigned($signed({9'h000, add_18630, umul_18454[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_18810 = umul22b_16b_x_6b(array_index_18750, 6'h35);
  assign add_18812 = {1'h0, umul_18620[21:7]} + 16'h007d;
  assign sel_18817 = $signed({1'h0, smod_18568[15:0]}) < $signed({1'h0, sel_18627}) ? smod_18568[15:0] : sel_18627;
  assign umul_18818 = umul22b_16b_x_6b(array_index_18756, 6'h35);
  assign add_18820 = {1'h0, umul_18628[21:7]} + 16'h007d;
  assign sel_18825 = $signed({1'h0, smod_18574[15:0]}) < $signed({1'h0, sel_18635}) ? smod_18574[15:0] : sel_18635;
  assign smod_18829 = $unsigned($signed({8'h00, add_18692, umul_18512[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_18835 = $unsigned($signed({8'h00, add_18698, umul_18516[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_18841 = $unsigned($signed({8'h00, add_18704, umul_18520[0]}) % $signed(32'h0000_3ffd));
  assign smod_18846 = $unsigned($signed({8'h00, add_18712, umul_18526[0]}) % $signed(32'h0000_3ffd));
  assign smod_18851 = $unsigned($signed({9'h000, add_18720, umul_18532[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_18856 = $unsigned($signed({9'h000, add_18728, umul_18540[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_18861 = $unsigned($signed({9'h000, add_18736, umul_18548[0]}) % $signed(32'h0000_3ffd));
  assign smod_18866 = $unsigned($signed({9'h000, add_18744, umul_18556[0]}) % $signed(32'h0000_3ffd));
  assign umul_18882 = umul23b_16b_x_7b(array_index_18264, 7'h49);
  assign add_18884 = {1'h0, umul_18690[22:3]} + 21'h00_07e9;
  assign sel_18889 = $signed({1'h0, smod_18639[15:0]}) < $signed(17'h0_3ffd) ? smod_18639[15:0] : 16'h3ffd;
  assign umul_18890 = umul23b_16b_x_7b(array_index_18271, 7'h49);
  assign add_18892 = {1'h0, umul_18696[22:3]} + 21'h00_07e9;
  assign sel_18897 = $signed({1'h0, smod_18643[15:0]}) < $signed(17'h0_3ffd) ? smod_18643[15:0] : 16'h3ffd;
  assign umul_18898 = umul23b_16b_x_7b(array_index_18398, 7'h47);
  assign add_18900 = {1'h0, umul_18702[22:1]} + 23'h00_1f8b;
  assign sel_18905 = $signed({1'h0, smod_18647[15:0]}) < $signed({1'h0, sel_18709}) ? smod_18647[15:0] : sel_18709;
  assign umul_18906 = umul23b_16b_x_7b(array_index_18404, 7'h47);
  assign add_18908 = {1'h0, umul_18710[22:1]} + 23'h00_1f8b;
  assign sel_18913 = $signed({1'h0, smod_18653[15:0]}) < $signed({1'h0, sel_18717}) ? smod_18653[15:0] : sel_18717;
  assign umul_18914 = umul22b_16b_x_6b(array_index_18564, 6'h3d);
  assign add_18916 = {1'h0, umul_18718[21:2]} + 21'h00_0fb9;
  assign sel_18921 = $signed({1'h0, smod_18659[15:0]}) < $signed({1'h0, sel_18725}) ? smod_18659[15:0] : sel_18725;
  assign umul_18922 = umul22b_16b_x_6b(array_index_18570, 6'h3d);
  assign add_18924 = {1'h0, umul_18726[21:2]} + 21'h00_0fb9;
  assign sel_18929 = $signed({1'h0, smod_18664[15:0]}) < $signed({1'h0, sel_18733}) ? smod_18664[15:0] : sel_18733;
  assign umul_18930 = umul22b_16b_x_6b(array_index_18750, 6'h3b);
  assign add_18932 = {1'h0, umul_18734[21:1]} + 22'h00_1f59;
  assign sel_18937 = $signed({1'h0, smod_18669[15:0]}) < $signed({1'h0, sel_18741}) ? smod_18669[15:0] : sel_18741;
  assign umul_18938 = umul22b_16b_x_6b(array_index_18756, 6'h3b);
  assign add_18940 = {1'h0, umul_18742[21:1]} + 22'h00_1f59;
  assign sel_18945 = $signed({1'h0, smod_18674[15:0]}) < $signed({1'h0, sel_18749}) ? smod_18674[15:0] : sel_18749;
  assign array_index_18946 = set1_unflattened[4'h7];
  assign smod_18950 = $unsigned($signed({9'h000, add_18812, umul_18620[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_18952 = set2_unflattened[4'h7];
  assign smod_18956 = $unsigned($signed({9'h000, add_18820, umul_18628[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_19006 = umul22b_16b_x_6b(array_index_18946, 6'h35);
  assign add_19008 = {1'h0, umul_18810[21:7]} + 16'h007d;
  assign sel_19013 = $signed({1'h0, smod_18754[15:0]}) < $signed({1'h0, sel_18817}) ? smod_18754[15:0] : sel_18817;
  assign umul_19014 = umul22b_16b_x_6b(array_index_18952, 6'h35);
  assign add_19016 = {1'h0, umul_18818[21:7]} + 16'h007d;
  assign sel_19021 = $signed({1'h0, smod_18760[15:0]}) < $signed({1'h0, sel_18825}) ? smod_18760[15:0] : sel_18825;
  assign smod_19025 = $unsigned($signed({8'h00, add_18884, umul_18690[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19030 = $unsigned($signed({8'h00, add_18892, umul_18696[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19035 = $unsigned($signed({8'h00, add_18900, umul_18702[0]}) % $signed(32'h0000_3ffd));
  assign smod_19040 = $unsigned($signed({8'h00, add_18908, umul_18710[0]}) % $signed(32'h0000_3ffd));
  assign smod_19045 = $unsigned($signed({9'h000, add_18916, umul_18718[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_19050 = $unsigned($signed({9'h000, add_18924, umul_18726[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_19055 = $unsigned($signed({9'h000, add_18932, umul_18734[0]}) % $signed(32'h0000_3ffd));
  assign smod_19060 = $unsigned($signed({9'h000, add_18940, umul_18742[0]}) % $signed(32'h0000_3ffd));
  assign umul_19076 = umul23b_16b_x_7b(array_index_18398, 7'h49);
  assign add_19078 = {1'h0, umul_18882[22:3]} + 21'h00_07e9;
  assign sel_19083 = $signed({1'h0, smod_18829[15:0]}) < $signed({1'h0, sel_18889}) ? smod_18829[15:0] : sel_18889;
  assign umul_19084 = umul23b_16b_x_7b(array_index_18404, 7'h49);
  assign add_19086 = {1'h0, umul_18890[22:3]} + 21'h00_07e9;
  assign sel_19091 = $signed({1'h0, smod_18835[15:0]}) < $signed({1'h0, sel_18897}) ? smod_18835[15:0] : sel_18897;
  assign umul_19092 = umul23b_16b_x_7b(array_index_18564, 7'h47);
  assign add_19094 = {1'h0, umul_18898[22:1]} + 23'h00_1f8b;
  assign sel_19099 = $signed({1'h0, smod_18841[15:0]}) < $signed({1'h0, sel_18905}) ? smod_18841[15:0] : sel_18905;
  assign umul_19100 = umul23b_16b_x_7b(array_index_18570, 7'h47);
  assign add_19102 = {1'h0, umul_18906[22:1]} + 23'h00_1f8b;
  assign sel_19107 = $signed({1'h0, smod_18846[15:0]}) < $signed({1'h0, sel_18913}) ? smod_18846[15:0] : sel_18913;
  assign umul_19108 = umul22b_16b_x_6b(array_index_18750, 6'h3d);
  assign add_19110 = {1'h0, umul_18914[21:2]} + 21'h00_0fb9;
  assign sel_19115 = $signed({1'h0, smod_18851[15:0]}) < $signed({1'h0, sel_18921}) ? smod_18851[15:0] : sel_18921;
  assign umul_19116 = umul22b_16b_x_6b(array_index_18756, 6'h3d);
  assign add_19118 = {1'h0, umul_18922[21:2]} + 21'h00_0fb9;
  assign sel_19123 = $signed({1'h0, smod_18856[15:0]}) < $signed({1'h0, sel_18929}) ? smod_18856[15:0] : sel_18929;
  assign umul_19124 = umul22b_16b_x_6b(array_index_18946, 6'h3b);
  assign add_19126 = {1'h0, umul_18930[21:1]} + 22'h00_1f59;
  assign sel_19131 = $signed({1'h0, smod_18861[15:0]}) < $signed({1'h0, sel_18937}) ? smod_18861[15:0] : sel_18937;
  assign umul_19132 = umul22b_16b_x_6b(array_index_18952, 6'h3b);
  assign add_19134 = {1'h0, umul_18938[21:1]} + 22'h00_1f59;
  assign sel_19139 = $signed({1'h0, smod_18866[15:0]}) < $signed({1'h0, sel_18945}) ? smod_18866[15:0] : sel_18945;
  assign array_index_19140 = set1_unflattened[4'h8];
  assign smod_19144 = $unsigned($signed({9'h000, add_19008, umul_18810[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_19146 = set2_unflattened[4'h8];
  assign smod_19150 = $unsigned($signed({9'h000, add_19016, umul_18818[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_19200 = umul22b_16b_x_6b(array_index_19140, 6'h35);
  assign add_19202 = {1'h0, umul_19006[21:7]} + 16'h007d;
  assign sel_19207 = $signed({1'h0, smod_18950[15:0]}) < $signed({1'h0, sel_19013}) ? smod_18950[15:0] : sel_19013;
  assign umul_19208 = umul22b_16b_x_6b(array_index_19146, 6'h35);
  assign add_19210 = {1'h0, umul_19014[21:7]} + 16'h007d;
  assign sel_19215 = $signed({1'h0, smod_18956[15:0]}) < $signed({1'h0, sel_19021}) ? smod_18956[15:0] : sel_19021;
  assign smod_19219 = $unsigned($signed({8'h00, add_19078, umul_18882[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19224 = $unsigned($signed({8'h00, add_19086, umul_18890[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19229 = $unsigned($signed({8'h00, add_19094, umul_18898[0]}) % $signed(32'h0000_3ffd));
  assign smod_19234 = $unsigned($signed({8'h00, add_19102, umul_18906[0]}) % $signed(32'h0000_3ffd));
  assign smod_19239 = $unsigned($signed({9'h000, add_19110, umul_18914[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_19244 = $unsigned($signed({9'h000, add_19118, umul_18922[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_19249 = $unsigned($signed({9'h000, add_19126, umul_18930[0]}) % $signed(32'h0000_3ffd));
  assign smod_19254 = $unsigned($signed({9'h000, add_19134, umul_18938[0]}) % $signed(32'h0000_3ffd));
  assign umul_19270 = umul23b_16b_x_7b(array_index_18564, 7'h49);
  assign add_19272 = {1'h0, umul_19076[22:3]} + 21'h00_07e9;
  assign sel_19277 = $signed({1'h0, smod_19025[15:0]}) < $signed({1'h0, sel_19083}) ? smod_19025[15:0] : sel_19083;
  assign umul_19278 = umul23b_16b_x_7b(array_index_18570, 7'h49);
  assign add_19280 = {1'h0, umul_19084[22:3]} + 21'h00_07e9;
  assign sel_19285 = $signed({1'h0, smod_19030[15:0]}) < $signed({1'h0, sel_19091}) ? smod_19030[15:0] : sel_19091;
  assign umul_19286 = umul23b_16b_x_7b(array_index_18750, 7'h47);
  assign add_19288 = {1'h0, umul_19092[22:1]} + 23'h00_1f8b;
  assign sel_19293 = $signed({1'h0, smod_19035[15:0]}) < $signed({1'h0, sel_19099}) ? smod_19035[15:0] : sel_19099;
  assign umul_19294 = umul23b_16b_x_7b(array_index_18756, 7'h47);
  assign add_19296 = {1'h0, umul_19100[22:1]} + 23'h00_1f8b;
  assign sel_19301 = $signed({1'h0, smod_19040[15:0]}) < $signed({1'h0, sel_19107}) ? smod_19040[15:0] : sel_19107;
  assign umul_19302 = umul22b_16b_x_6b(array_index_18946, 6'h3d);
  assign add_19304 = {1'h0, umul_19108[21:2]} + 21'h00_0fb9;
  assign sel_19309 = $signed({1'h0, smod_19045[15:0]}) < $signed({1'h0, sel_19115}) ? smod_19045[15:0] : sel_19115;
  assign umul_19310 = umul22b_16b_x_6b(array_index_18952, 6'h3d);
  assign add_19312 = {1'h0, umul_19116[21:2]} + 21'h00_0fb9;
  assign sel_19317 = $signed({1'h0, smod_19050[15:0]}) < $signed({1'h0, sel_19123}) ? smod_19050[15:0] : sel_19123;
  assign umul_19318 = umul22b_16b_x_6b(array_index_19140, 6'h3b);
  assign add_19320 = {1'h0, umul_19124[21:1]} + 22'h00_1f59;
  assign sel_19325 = $signed({1'h0, smod_19055[15:0]}) < $signed({1'h0, sel_19131}) ? smod_19055[15:0] : sel_19131;
  assign umul_19326 = umul22b_16b_x_6b(array_index_19146, 6'h3b);
  assign add_19328 = {1'h0, umul_19132[21:1]} + 22'h00_1f59;
  assign sel_19333 = $signed({1'h0, smod_19060[15:0]}) < $signed({1'h0, sel_19139}) ? smod_19060[15:0] : sel_19139;
  assign array_index_19334 = set1_unflattened[4'h9];
  assign smod_19338 = $unsigned($signed({9'h000, add_19202, umul_19006[6:0]}) % $signed(32'h0000_3ffd));
  assign array_index_19340 = set2_unflattened[4'h9];
  assign smod_19344 = $unsigned($signed({9'h000, add_19210, umul_19014[6:0]}) % $signed(32'h0000_3ffd));
  assign umul_19394 = umul22b_16b_x_6b(array_index_19334, 6'h35);
  assign add_19396 = {1'h0, umul_19200[21:7]} + 16'h007d;
  assign sel_19401 = $signed({1'h0, smod_19144[15:0]}) < $signed({1'h0, sel_19207}) ? smod_19144[15:0] : sel_19207;
  assign umul_19402 = umul22b_16b_x_6b(array_index_19340, 6'h35);
  assign add_19404 = {1'h0, umul_19208[21:7]} + 16'h007d;
  assign sel_19409 = $signed({1'h0, smod_19150[15:0]}) < $signed({1'h0, sel_19215}) ? smod_19150[15:0] : sel_19215;
  assign smod_19413 = $unsigned($signed({8'h00, add_19272, umul_19076[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19418 = $unsigned($signed({8'h00, add_19280, umul_19084[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19423 = $unsigned($signed({8'h00, add_19288, umul_19092[0]}) % $signed(32'h0000_3ffd));
  assign smod_19428 = $unsigned($signed({8'h00, add_19296, umul_19100[0]}) % $signed(32'h0000_3ffd));
  assign smod_19433 = $unsigned($signed({9'h000, add_19304, umul_19108[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_19438 = $unsigned($signed({9'h000, add_19312, umul_19116[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_19443 = $unsigned($signed({9'h000, add_19320, umul_19124[0]}) % $signed(32'h0000_3ffd));
  assign smod_19448 = $unsigned($signed({9'h000, add_19328, umul_19132[0]}) % $signed(32'h0000_3ffd));
  assign umul_19462 = umul23b_16b_x_7b(array_index_18750, 7'h49);
  assign add_19464 = {1'h0, umul_19270[22:3]} + 21'h00_07e9;
  assign sel_19469 = $signed({1'h0, smod_19219[15:0]}) < $signed({1'h0, sel_19277}) ? smod_19219[15:0] : sel_19277;
  assign umul_19470 = umul23b_16b_x_7b(array_index_18756, 7'h49);
  assign add_19472 = {1'h0, umul_19278[22:3]} + 21'h00_07e9;
  assign sel_19477 = $signed({1'h0, smod_19224[15:0]}) < $signed({1'h0, sel_19285}) ? smod_19224[15:0] : sel_19285;
  assign umul_19478 = umul23b_16b_x_7b(array_index_18946, 7'h47);
  assign add_19480 = {1'h0, umul_19286[22:1]} + 23'h00_1f8b;
  assign sel_19485 = $signed({1'h0, smod_19229[15:0]}) < $signed({1'h0, sel_19293}) ? smod_19229[15:0] : sel_19293;
  assign umul_19486 = umul23b_16b_x_7b(array_index_18952, 7'h47);
  assign add_19488 = {1'h0, umul_19294[22:1]} + 23'h00_1f8b;
  assign sel_19493 = $signed({1'h0, smod_19234[15:0]}) < $signed({1'h0, sel_19301}) ? smod_19234[15:0] : sel_19301;
  assign umul_19494 = umul22b_16b_x_6b(array_index_19140, 6'h3d);
  assign add_19496 = {1'h0, umul_19302[21:2]} + 21'h00_0fb9;
  assign sel_19501 = $signed({1'h0, smod_19239[15:0]}) < $signed({1'h0, sel_19309}) ? smod_19239[15:0] : sel_19309;
  assign umul_19502 = umul22b_16b_x_6b(array_index_19146, 6'h3d);
  assign add_19504 = {1'h0, umul_19310[21:2]} + 21'h00_0fb9;
  assign sel_19509 = $signed({1'h0, smod_19244[15:0]}) < $signed({1'h0, sel_19317}) ? smod_19244[15:0] : sel_19317;
  assign umul_19510 = umul22b_16b_x_6b(array_index_19334, 6'h3b);
  assign add_19512 = {1'h0, umul_19318[21:1]} + 22'h00_1f59;
  assign sel_19517 = $signed({1'h0, smod_19249[15:0]}) < $signed({1'h0, sel_19325}) ? smod_19249[15:0] : sel_19325;
  assign umul_19518 = umul22b_16b_x_6b(array_index_19340, 6'h3b);
  assign add_19520 = {1'h0, umul_19326[21:1]} + 22'h00_1f59;
  assign sel_19525 = $signed({1'h0, smod_19254[15:0]}) < $signed({1'h0, sel_19333}) ? smod_19254[15:0] : sel_19333;
  assign smod_19528 = $unsigned($signed({9'h000, add_19396, umul_19200[6:0]}) % $signed(32'h0000_3ffd));
  assign smod_19532 = $unsigned($signed({9'h000, add_19404, umul_19208[6:0]}) % $signed(32'h0000_3ffd));
  assign add_19583 = {1'h0, umul_19394[21:7]} + 16'h007d;
  assign sel_19588 = $signed({1'h0, smod_19338[15:0]}) < $signed({1'h0, sel_19401}) ? smod_19338[15:0] : sel_19401;
  assign add_19590 = {1'h0, umul_19402[21:7]} + 16'h007d;
  assign sel_19595 = $signed({1'h0, smod_19344[15:0]}) < $signed({1'h0, sel_19409}) ? smod_19344[15:0] : sel_19409;
  assign smod_19599 = $unsigned($signed({8'h00, add_19464, umul_19270[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19604 = $unsigned($signed({8'h00, add_19472, umul_19278[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19609 = $unsigned($signed({8'h00, add_19480, umul_19286[0]}) % $signed(32'h0000_3ffd));
  assign smod_19614 = $unsigned($signed({8'h00, add_19488, umul_19294[0]}) % $signed(32'h0000_3ffd));
  assign smod_19619 = $unsigned($signed({9'h000, add_19496, umul_19302[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_19624 = $unsigned($signed({9'h000, add_19504, umul_19310[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_19628 = $unsigned($signed({9'h000, add_19512, umul_19318[0]}) % $signed(32'h0000_3ffd));
  assign smod_19632 = $unsigned($signed({9'h000, add_19520, umul_19326[0]}) % $signed(32'h0000_3ffd));
  assign umul_19642 = umul23b_16b_x_7b(array_index_18946, 7'h49);
  assign add_19644 = {1'h0, umul_19462[22:3]} + 21'h00_07e9;
  assign sel_19649 = $signed({1'h0, smod_19413[15:0]}) < $signed({1'h0, sel_19469}) ? smod_19413[15:0] : sel_19469;
  assign umul_19650 = umul23b_16b_x_7b(array_index_18952, 7'h49);
  assign add_19652 = {1'h0, umul_19470[22:3]} + 21'h00_07e9;
  assign sel_19657 = $signed({1'h0, smod_19418[15:0]}) < $signed({1'h0, sel_19477}) ? smod_19418[15:0] : sel_19477;
  assign umul_19658 = umul23b_16b_x_7b(array_index_19140, 7'h47);
  assign add_19660 = {1'h0, umul_19478[22:1]} + 23'h00_1f8b;
  assign sel_19665 = $signed({1'h0, smod_19423[15:0]}) < $signed({1'h0, sel_19485}) ? smod_19423[15:0] : sel_19485;
  assign umul_19666 = umul23b_16b_x_7b(array_index_19146, 7'h47);
  assign add_19668 = {1'h0, umul_19486[22:1]} + 23'h00_1f8b;
  assign sel_19673 = $signed({1'h0, smod_19428[15:0]}) < $signed({1'h0, sel_19493}) ? smod_19428[15:0] : sel_19493;
  assign umul_19674 = umul22b_16b_x_6b(array_index_19334, 6'h3d);
  assign add_19676 = {1'h0, umul_19494[21:2]} + 21'h00_0fb9;
  assign sel_19681 = $signed({1'h0, smod_19433[15:0]}) < $signed({1'h0, sel_19501}) ? smod_19433[15:0] : sel_19501;
  assign umul_19682 = umul22b_16b_x_6b(array_index_19340, 6'h3d);
  assign add_19684 = {1'h0, umul_19502[21:2]} + 21'h00_0fb9;
  assign sel_19689 = $signed({1'h0, smod_19438[15:0]}) < $signed({1'h0, sel_19509}) ? smod_19438[15:0] : sel_19509;
  assign add_19691 = {1'h0, umul_19510[21:1]} + 22'h00_1f59;
  assign sel_19696 = $signed({1'h0, smod_19443[15:0]}) < $signed({1'h0, sel_19517}) ? smod_19443[15:0] : sel_19517;
  assign add_19698 = {1'h0, umul_19518[21:1]} + 22'h00_1f59;
  assign sel_19703 = $signed({1'h0, smod_19448[15:0]}) < $signed({1'h0, sel_19525}) ? smod_19448[15:0] : sel_19525;
  assign smod_19704 = $unsigned($signed({9'h000, add_19583, umul_19394[6:0]}) % $signed(32'h0000_3ffd));
  assign smod_19706 = $unsigned($signed({9'h000, add_19590, umul_19402[6:0]}) % $signed(32'h0000_3ffd));
  assign sel_19755 = $signed({1'h0, smod_19528[15:0]}) < $signed({1'h0, sel_19588}) ? smod_19528[15:0] : sel_19588;
  assign sel_19759 = $signed({1'h0, smod_19532[15:0]}) < $signed({1'h0, sel_19595}) ? smod_19532[15:0] : sel_19595;
  assign smod_19763 = $unsigned($signed({8'h00, add_19644, umul_19462[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19768 = $unsigned($signed({8'h00, add_19652, umul_19470[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19773 = $unsigned($signed({8'h00, add_19660, umul_19478[0]}) % $signed(32'h0000_3ffd));
  assign smod_19778 = $unsigned($signed({8'h00, add_19668, umul_19486[0]}) % $signed(32'h0000_3ffd));
  assign smod_19782 = $unsigned($signed({9'h000, add_19676, umul_19494[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_19786 = $unsigned($signed({9'h000, add_19684, umul_19502[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_19788 = $unsigned($signed({9'h000, add_19691, umul_19510[0]}) % $signed(32'h0000_3ffd));
  assign smod_19790 = $unsigned($signed({9'h000, add_19698, umul_19518[0]}) % $signed(32'h0000_3ffd));
  assign umul_19796 = umul23b_16b_x_7b(array_index_19140, 7'h49);
  assign add_19798 = {1'h0, umul_19642[22:3]} + 21'h00_07e9;
  assign sel_19803 = $signed({1'h0, smod_19599[15:0]}) < $signed({1'h0, sel_19649}) ? smod_19599[15:0] : sel_19649;
  assign umul_19804 = umul23b_16b_x_7b(array_index_19146, 7'h49);
  assign add_19806 = {1'h0, umul_19650[22:3]} + 21'h00_07e9;
  assign sel_19811 = $signed({1'h0, smod_19604[15:0]}) < $signed({1'h0, sel_19657}) ? smod_19604[15:0] : sel_19657;
  assign umul_19812 = umul23b_16b_x_7b(array_index_19334, 7'h47);
  assign add_19814 = {1'h0, umul_19658[22:1]} + 23'h00_1f8b;
  assign sel_19819 = $signed({1'h0, smod_19609[15:0]}) < $signed({1'h0, sel_19665}) ? smod_19609[15:0] : sel_19665;
  assign umul_19820 = umul23b_16b_x_7b(array_index_19340, 7'h47);
  assign add_19822 = {1'h0, umul_19666[22:1]} + 23'h00_1f8b;
  assign sel_19827 = $signed({1'h0, smod_19614[15:0]}) < $signed({1'h0, sel_19673}) ? smod_19614[15:0] : sel_19673;
  assign add_19829 = {1'h0, umul_19674[21:2]} + 21'h00_0fb9;
  assign sel_19834 = $signed({1'h0, smod_19619[15:0]}) < $signed({1'h0, sel_19681}) ? smod_19619[15:0] : sel_19681;
  assign add_19836 = {1'h0, umul_19682[21:2]} + 21'h00_0fb9;
  assign sel_19841 = $signed({1'h0, smod_19624[15:0]}) < $signed({1'h0, sel_19689}) ? smod_19624[15:0] : sel_19689;
  assign sel_19845 = $signed({1'h0, smod_19628[15:0]}) < $signed({1'h0, sel_19696}) ? smod_19628[15:0] : sel_19696;
  assign sel_19849 = $signed({1'h0, smod_19632[15:0]}) < $signed({1'h0, sel_19703}) ? smod_19632[15:0] : sel_19703;
  assign smod_19893 = $unsigned($signed({8'h00, add_19798, umul_19642[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19898 = $unsigned($signed({8'h00, add_19806, umul_19650[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19902 = $unsigned($signed({8'h00, add_19814, umul_19658[0]}) % $signed(32'h0000_3ffd));
  assign smod_19906 = $unsigned($signed({8'h00, add_19822, umul_19666[0]}) % $signed(32'h0000_3ffd));
  assign smod_19908 = $unsigned($signed({9'h000, add_19829, umul_19674[1:0]}) % $signed(32'h0000_3ffd));
  assign smod_19910 = $unsigned($signed({9'h000, add_19836, umul_19682[1:0]}) % $signed(32'h0000_3ffd));
  assign umul_19916 = umul23b_16b_x_7b(array_index_19334, 7'h49);
  assign add_19918 = {1'h0, umul_19796[22:3]} + 21'h00_07e9;
  assign sel_19923 = $signed({1'h0, smod_19763[15:0]}) < $signed({1'h0, sel_19803}) ? smod_19763[15:0] : sel_19803;
  assign umul_19924 = umul23b_16b_x_7b(array_index_19340, 7'h49);
  assign add_19926 = {1'h0, umul_19804[22:3]} + 21'h00_07e9;
  assign sel_19931 = $signed({1'h0, smod_19768[15:0]}) < $signed({1'h0, sel_19811}) ? smod_19768[15:0] : sel_19811;
  assign add_19933 = {1'h0, umul_19812[22:1]} + 23'h00_1f8b;
  assign sel_19938 = $signed({1'h0, smod_19773[15:0]}) < $signed({1'h0, sel_19819}) ? smod_19773[15:0] : sel_19819;
  assign add_19940 = {1'h0, umul_19820[22:1]} + 23'h00_1f8b;
  assign sel_19945 = $signed({1'h0, smod_19778[15:0]}) < $signed({1'h0, sel_19827}) ? smod_19778[15:0] : sel_19827;
  assign sel_19949 = $signed({1'h0, smod_19782[15:0]}) < $signed({1'h0, sel_19834}) ? smod_19782[15:0] : sel_19834;
  assign sel_19953 = $signed({1'h0, smod_19786[15:0]}) < $signed({1'h0, sel_19841}) ? smod_19786[15:0] : sel_19841;
  assign concat_19956 = {1'h0, ($signed({1'h0, smod_19704[15:0]}) < $signed({1'h0, sel_19755}) ? smod_19704[15:0] : sel_19755) == ($signed({1'h0, smod_19706[15:0]}) < $signed({1'h0, sel_19759}) ? smod_19706[15:0] : sel_19759)};
  assign add_19983 = concat_19956 + 2'h1;
  assign smod_19986 = $unsigned($signed({8'h00, add_19918, umul_19796[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19990 = $unsigned($signed({8'h00, add_19926, umul_19804[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_19992 = $unsigned($signed({8'h00, add_19933, umul_19812[0]}) % $signed(32'h0000_3ffd));
  assign smod_19994 = $unsigned($signed({8'h00, add_19940, umul_19820[0]}) % $signed(32'h0000_3ffd));
  assign add_20001 = {1'h0, umul_19916[22:3]} + 21'h00_07e9;
  assign sel_20006 = $signed({1'h0, smod_19893[15:0]}) < $signed({1'h0, sel_19923}) ? smod_19893[15:0] : sel_19923;
  assign add_20008 = {1'h0, umul_19924[22:3]} + 21'h00_07e9;
  assign sel_20013 = $signed({1'h0, smod_19898[15:0]}) < $signed({1'h0, sel_19931}) ? smod_19898[15:0] : sel_19931;
  assign sel_20017 = $signed({1'h0, smod_19902[15:0]}) < $signed({1'h0, sel_19938}) ? smod_19902[15:0] : sel_19938;
  assign sel_20021 = $signed({1'h0, smod_19906[15:0]}) < $signed({1'h0, sel_19945}) ? smod_19906[15:0] : sel_19945;
  assign concat_20024 = {1'h0, ($signed({1'h0, smod_19788[15:0]}) < $signed({1'h0, sel_19845}) ? smod_19788[15:0] : sel_19845) == ($signed({1'h0, smod_19790[15:0]}) < $signed({1'h0, sel_19849}) ? smod_19790[15:0] : sel_19849) ? add_19983 : concat_19956};
  assign add_20039 = concat_20024 + 3'h1;
  assign smod_20040 = $unsigned($signed({8'h00, add_20001, umul_19916[2:0]}) % $signed(32'h0000_3ffd));
  assign smod_20042 = $unsigned($signed({8'h00, add_20008, umul_19924[2:0]}) % $signed(32'h0000_3ffd));
  assign sel_20051 = $signed({1'h0, smod_19986[15:0]}) < $signed({1'h0, sel_20006}) ? smod_19986[15:0] : sel_20006;
  assign sel_20055 = $signed({1'h0, smod_19990[15:0]}) < $signed({1'h0, sel_20013}) ? smod_19990[15:0] : sel_20013;
  assign concat_20058 = {1'h0, ($signed({1'h0, smod_19908[15:0]}) < $signed({1'h0, sel_19949}) ? smod_19908[15:0] : sel_19949) == ($signed({1'h0, smod_19910[15:0]}) < $signed({1'h0, sel_19953}) ? smod_19910[15:0] : sel_19953) ? add_20039 : concat_20024};
  assign add_20065 = concat_20058 + 4'h1;
  assign concat_20072 = {1'h0, ($signed({1'h0, smod_19992[15:0]}) < $signed({1'h0, sel_20017}) ? smod_19992[15:0] : sel_20017) == ($signed({1'h0, smod_19994[15:0]}) < $signed({1'h0, sel_20021}) ? smod_19994[15:0] : sel_20021) ? add_20065 : concat_20058};
  assign add_20075 = concat_20072 + 5'h01;
  assign out = {{11'h000, ($signed({1'h0, smod_20040[15:0]}) < $signed({1'h0, sel_20051}) ? smod_20040[15:0] : sel_20051) == ($signed({1'h0, smod_20042[15:0]}) < $signed({1'h0, sel_20055}) ? smod_20042[15:0] : sel_20055) ? add_20075 : concat_20072}, {set1_unflattened[9], set1_unflattened[8], set1_unflattened[7], set1_unflattened[6], set1_unflattened[5], set1_unflattened[4], set1_unflattened[3], set1_unflattened[2], set1_unflattened[1], set1_unflattened[0]}, {set2_unflattened[9], set2_unflattened[8], set2_unflattened[7], set2_unflattened[6], set2_unflattened[5], set2_unflattened[4], set2_unflattened[3], set2_unflattened[2], set2_unflattened[1], set2_unflattened[0]}};
endmodule
